// Benchmark "SKOLEMFORMULA" written by ABC on Wed May 18 01:32:33 2022

module SKOLEMFORMULA ( 
    i0, i1,
    i2  );
  input  i0, i1;
  output i2;
  assign i2 = i0 & i1;
endmodule


