// Benchmark "SKOLEMFORMULA" written by ABC on Fri May 27 13:38:44 2022

module SKOLEMFORMULA ( 
    i0, i1,
    i2, i3  );
  input  i0, i1;
  output i2, i3;
  assign i3 = 1'b1;
  assign i2 = i0;
endmodule


