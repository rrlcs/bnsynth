// Verilog file written by procedure writeCombinationalCircuitInVerilog
//Skolem functions to be generated for i_ variables
module formula ( i_1, i_2, i_3, i_4, i_5, i_6, i_7, i_8, i_9, i_10, i_11, i_12, i_13, i_14, i_15, i_16, i_17, i_18, i_19, i_20, i_21, i_22, i_23, i_24, i_25, i_26, i_27, i_28, i_29, x_30, x_31, x_32, x_33, x_34, x_35, x_36, x_37, x_38, x_39, x_40, x_41, x_42, x_43, x_44, x_45, x_46, x_47, x_48, x_49, x_50, x_51, x_52, x_53, x_54, x_55, x_56, x_57, x_58, x_59, x_60, x_61, x_62, x_63, x_64, x_65, x_66, x_67, x_68, x_69, x_70, x_71, x_72, x_73, x_74, x_75, x_76, x_77, x_78, x_79, x_80, x_81, x_82, x_83, x_84, x_85, x_86, x_87, x_88, x_89, x_90, x_91, x_92, x_93, x_94, x_95, x_96, x_97, x_98, x_99, x_100, x_101, x_102, x_103, x_104, x_105, x_106, x_107, x_108, x_109, x_110, x_111, x_112, x_113, x_114, x_115, x_116, x_117, x_118, x_119, x_120, x_121, x_122, x_123, x_124, x_125, x_126, x_127, x_128, x_129, x_130, x_131, x_132, x_133, x_134, x_135, x_136, x_137, x_138, x_139, x_140, x_141, x_142, x_143, x_144, x_145, x_146, x_147, x_148, x_149, x_150, x_151, x_152, x_153, x_154, x_155, x_156, x_157, x_158, x_159, x_160, x_161, x_162, x_163, x_164, x_165, x_166, x_167, x_168, x_169, x_170, x_171, x_172, x_173, x_174, x_175, x_176, x_177, x_178, x_179, x_180, x_181, x_182, x_183, x_184, x_185, x_186, x_187, x_188, x_189, x_190, x_191, x_192, x_193, x_194, x_195, x_196, x_197, x_198, x_199, x_200, x_201, x_202, x_203, x_204, x_205, x_206, x_207, x_208, x_209, x_210, x_211, x_212, x_213, x_214, x_215, x_216, x_217, x_218, x_219, x_220, x_221, x_222, x_223, x_224, x_225, x_226, x_227, x_228, x_229, x_230, x_231, x_232, x_233, x_234, x_235, x_236, x_237, x_238, x_239, x_240, x_241, x_242, x_243, x_244, x_245, x_246, x_247, x_248, x_249, x_250, x_251, x_252, x_253, x_254, x_255, x_256, x_257, x_258, x_259, x_260, x_261, x_262, x_263, x_264, x_265, x_266, x_267, x_268, x_269, x_270, x_271, x_272, x_273, x_274, x_275, x_276, x_277, x_278, x_279, x_280, x_281, x_282, x_283, x_284, x_285, x_286, x_287, x_288, x_289, x_290, x_291, x_292, x_293, x_294, x_295, x_296, x_297, x_298, x_299, x_300, x_301, x_302, x_303, x_304, x_305, x_306, x_307, x_308, x_309, x_310, x_311, x_312, x_313, x_314, x_315, x_316, x_317, x_318, x_319, x_320, x_321, x_322, x_323, x_324, x_325, x_326, x_327, x_328, x_329, x_330, x_331, x_332, x_333, x_334, x_335, x_336, x_337, x_338, x_339, x_340, x_341, x_342, x_343, x_344, x_345, o_1 );
input i_1;
input i_2;
input i_3;
input i_4;
input i_5;
input i_6;
input i_7;
input i_8;
input i_9;
input i_10;
input i_11;
input i_12;
input i_13;
input i_14;
input i_15;
input i_16;
input i_17;
input i_18;
input i_19;
input i_20;
input i_21;
input i_22;
input i_23;
input i_24;
input i_25;
input i_26;
input i_27;
input i_28;
input i_29;
input x_30;
input x_31;
input x_32;
input x_33;
input x_34;
input x_35;
input x_36;
input x_37;
input x_38;
input x_39;
input x_40;
input x_41;
input x_42;
input x_43;
input x_44;
input x_45;
input x_46;
input x_47;
input x_48;
input x_49;
input x_50;
input x_51;
input x_52;
input x_53;
input x_54;
input x_55;
input x_56;
input x_57;
input x_58;
input x_59;
input x_60;
input x_61;
input x_62;
input x_63;
input x_64;
input x_65;
input x_66;
input x_67;
input x_68;
input x_69;
input x_70;
input x_71;
input x_72;
input x_73;
input x_74;
input x_75;
input x_76;
input x_77;
input x_78;
input x_79;
input x_80;
input x_81;
input x_82;
input x_83;
input x_84;
input x_85;
input x_86;
input x_87;
input x_88;
input x_89;
input x_90;
input x_91;
input x_92;
input x_93;
input x_94;
input x_95;
input x_96;
input x_97;
input x_98;
input x_99;
input x_100;
input x_101;
input x_102;
input x_103;
input x_104;
input x_105;
input x_106;
input x_107;
input x_108;
input x_109;
input x_110;
input x_111;
input x_112;
input x_113;
input x_114;
input x_115;
input x_116;
input x_117;
input x_118;
input x_119;
input x_120;
input x_121;
input x_122;
input x_123;
input x_124;
input x_125;
input x_126;
input x_127;
input x_128;
input x_129;
input x_130;
input x_131;
input x_132;
input x_133;
input x_134;
input x_135;
input x_136;
input x_137;
input x_138;
input x_139;
input x_140;
input x_141;
input x_142;
input x_143;
input x_144;
input x_145;
input x_146;
input x_147;
input x_148;
input x_149;
input x_150;
input x_151;
input x_152;
input x_153;
input x_154;
input x_155;
input x_156;
input x_157;
input x_158;
input x_159;
input x_160;
input x_161;
input x_162;
input x_163;
input x_164;
input x_165;
input x_166;
input x_167;
input x_168;
input x_169;
input x_170;
input x_171;
input x_172;
input x_173;
input x_174;
input x_175;
input x_176;
input x_177;
input x_178;
input x_179;
input x_180;
input x_181;
input x_182;
input x_183;
input x_184;
input x_185;
input x_186;
input x_187;
input x_188;
input x_189;
input x_190;
input x_191;
input x_192;
input x_193;
input x_194;
input x_195;
input x_196;
input x_197;
input x_198;
input x_199;
input x_200;
input x_201;
input x_202;
input x_203;
input x_204;
input x_205;
input x_206;
input x_207;
input x_208;
input x_209;
input x_210;
input x_211;
input x_212;
input x_213;
input x_214;
input x_215;
input x_216;
input x_217;
input x_218;
input x_219;
input x_220;
input x_221;
input x_222;
input x_223;
input x_224;
input x_225;
input x_226;
input x_227;
input x_228;
input x_229;
input x_230;
input x_231;
input x_232;
input x_233;
input x_234;
input x_235;
input x_236;
input x_237;
input x_238;
input x_239;
input x_240;
input x_241;
input x_242;
input x_243;
input x_244;
input x_245;
input x_246;
input x_247;
input x_248;
input x_249;
input x_250;
input x_251;
input x_252;
input x_253;
input x_254;
input x_255;
input x_256;
input x_257;
input x_258;
input x_259;
input x_260;
input x_261;
input x_262;
input x_263;
input x_264;
input x_265;
input x_266;
input x_267;
input x_268;
input x_269;
input x_270;
input x_271;
input x_272;
input x_273;
input x_274;
input x_275;
input x_276;
input x_277;
input x_278;
input x_279;
input x_280;
input x_281;
input x_282;
input x_283;
input x_284;
input x_285;
input x_286;
input x_287;
input x_288;
input x_289;
input x_290;
input x_291;
input x_292;
input x_293;
input x_294;
input x_295;
input x_296;
input x_297;
input x_298;
input x_299;
input x_300;
input x_301;
input x_302;
input x_303;
input x_304;
input x_305;
input x_306;
input x_307;
input x_308;
input x_309;
input x_310;
input x_311;
input x_312;
input x_313;
input x_314;
input x_315;
input x_316;
input x_317;
input x_318;
input x_319;
input x_320;
input x_321;
input x_322;
input x_323;
input x_324;
input x_325;
input x_326;
input x_327;
input x_328;
input x_329;
input x_330;
input x_331;
input x_332;
input x_333;
input x_334;
input x_335;
input x_336;
input x_337;
input x_338;
input x_339;
input x_340;
input x_341;
input x_342;
input x_343;
input x_344;
input x_345;
output o_1;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire n_53;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_58;
wire n_59;
wire n_60;
wire n_61;
wire n_62;
wire n_63;
wire n_64;
wire n_65;
wire n_66;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;
wire n_95;
wire n_96;
wire n_97;
wire n_98;
wire n_99;
wire n_100;
wire n_101;
wire n_102;
wire n_103;
wire n_104;
wire n_105;
wire n_106;
wire n_107;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_112;
wire n_113;
wire n_114;
wire n_115;
wire n_116;
wire n_117;
wire n_118;
wire n_119;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_124;
wire n_125;
wire n_126;
wire n_127;
wire n_128;
wire n_129;
wire n_130;
wire n_131;
wire n_132;
wire n_133;
wire n_134;
wire n_135;
wire n_136;
wire n_137;
wire n_138;
wire n_139;
wire n_140;
wire n_141;
wire n_142;
wire n_143;
wire n_144;
wire n_145;
wire n_146;
wire n_147;
wire n_148;
wire n_149;
wire n_150;
wire n_151;
wire n_152;
wire n_153;
wire n_154;
wire n_155;
wire n_156;
wire n_157;
wire n_158;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_163;
wire n_164;
wire n_165;
wire n_166;
wire n_167;
wire n_168;
wire n_169;
wire n_170;
wire n_171;
wire n_172;
wire n_173;
wire n_174;
wire n_175;
wire n_176;
wire n_177;
wire n_178;
wire n_179;
wire n_180;
wire n_181;
wire n_182;
wire n_183;
wire n_184;
wire n_185;
wire n_186;
wire n_187;
wire n_188;
wire n_189;
wire n_190;
wire n_191;
wire n_192;
wire n_193;
wire n_194;
wire n_195;
wire n_196;
wire n_197;
wire n_198;
wire n_199;
wire n_200;
wire n_201;
wire n_202;
wire n_203;
wire n_204;
wire n_205;
wire n_206;
wire n_207;
wire n_208;
wire n_209;
wire n_210;
wire n_211;
wire n_212;
wire n_213;
wire n_214;
wire n_215;
wire n_216;
wire n_217;
wire n_218;
wire n_219;
wire n_220;
wire n_221;
wire n_222;
wire n_223;
wire n_224;
wire n_225;
wire n_226;
wire n_227;
wire n_228;
wire n_229;
wire n_230;
wire n_231;
wire n_232;
wire n_233;
wire n_234;
wire n_235;
wire n_236;
wire n_237;
wire n_238;
wire n_239;
wire n_240;
wire n_241;
wire n_242;
wire n_243;
wire n_244;
wire n_245;
wire n_246;
wire n_247;
wire n_248;
wire n_249;
wire n_250;
wire n_251;
wire n_252;
wire n_253;
wire n_254;
wire n_255;
wire n_256;
wire n_257;
wire n_258;
wire n_259;
wire n_260;
wire n_261;
wire n_262;
wire n_263;
wire n_264;
wire n_265;
wire n_266;
wire n_267;
wire n_268;
wire n_269;
wire n_270;
wire n_271;
wire n_272;
wire n_273;
wire n_274;
wire n_275;
wire n_276;
wire n_277;
wire n_278;
wire n_279;
wire n_280;
wire n_281;
wire n_282;
wire n_283;
wire n_284;
wire n_285;
wire n_286;
wire n_287;
wire n_288;
wire n_289;
wire n_290;
wire n_291;
wire n_292;
wire n_293;
wire n_294;
wire n_295;
wire n_296;
wire n_297;
wire n_298;
wire n_299;
wire n_300;
wire n_301;
wire n_302;
wire n_303;
wire n_304;
wire n_305;
wire n_306;
wire n_307;
wire n_308;
wire n_309;
wire n_310;
wire n_311;
wire n_312;
wire n_313;
wire n_314;
wire n_315;
wire n_316;
wire n_317;
wire n_318;
wire n_319;
wire n_320;
wire n_321;
wire n_322;
wire n_323;
wire n_324;
wire n_325;
wire n_326;
wire n_327;
wire n_328;
wire n_329;
wire n_330;
wire n_331;
wire n_332;
wire n_333;
wire n_334;
wire n_335;
wire n_336;
wire n_337;
wire n_338;
wire n_339;
wire n_340;
wire n_341;
wire n_342;
wire n_343;
wire n_344;
wire n_345;
wire n_346;
wire n_347;
wire n_348;
wire n_349;
wire n_350;
wire n_351;
wire n_352;
wire n_353;
wire n_354;
wire n_355;
wire n_356;
wire n_357;
wire n_358;
wire n_359;
wire n_360;
wire n_361;
wire n_362;
wire n_363;
wire n_364;
wire n_365;
wire n_366;
wire n_367;
wire n_368;
wire n_369;
wire n_370;
wire n_371;
wire n_372;
wire n_373;
wire n_374;
wire n_375;
wire n_376;
wire n_377;
wire n_378;
wire n_379;
wire n_380;
wire n_381;
wire n_382;
wire n_383;
wire n_384;
wire n_385;
wire n_386;
wire n_387;
wire n_388;
wire n_389;
wire n_390;
wire n_391;
wire n_392;
wire n_393;
wire n_394;
wire n_395;
wire n_396;
wire n_397;
wire n_398;
wire n_399;
wire n_400;
wire n_401;
wire n_402;
wire n_403;
wire n_404;
wire n_405;
wire n_406;
wire n_407;
wire n_408;
wire n_409;
wire n_410;
wire n_411;
wire n_412;
wire n_413;
wire n_414;
wire n_415;
wire n_416;
wire n_417;
wire n_418;
wire n_419;
wire n_420;
wire n_421;
wire n_422;
wire n_423;
wire n_424;
wire n_425;
wire n_426;
wire n_427;
wire n_428;
wire n_429;
wire n_430;
wire n_431;
wire n_432;
wire n_433;
wire n_434;
wire n_435;
wire n_436;
wire n_437;
wire n_438;
wire n_439;
wire n_440;
wire n_441;
wire n_442;
wire n_443;
wire n_444;
wire n_445;
wire n_446;
wire n_447;
wire n_448;
wire n_449;
wire n_450;
wire n_451;
wire n_452;
wire n_453;
wire n_454;
wire n_455;
wire n_456;
wire n_457;
wire n_458;
wire n_459;
wire n_460;
wire n_461;
wire n_462;
wire n_463;
wire n_464;
wire n_465;
wire n_466;
wire n_467;
wire n_468;
wire n_469;
wire n_470;
wire n_471;
wire n_472;
wire n_473;
wire n_474;
wire n_475;
wire n_476;
wire n_477;
wire n_478;
wire n_479;
wire n_480;
wire n_481;
wire n_482;
wire n_483;
wire n_484;
wire n_485;
wire n_486;
wire n_487;
wire n_488;
wire n_489;
wire n_490;
wire n_491;
wire n_492;
wire n_493;
wire n_494;
wire n_495;
wire n_496;
wire n_497;
wire n_498;
wire n_499;
wire n_500;
wire n_501;
wire n_502;
wire n_503;
wire n_504;
wire n_505;
wire n_506;
wire n_507;
wire n_508;
wire n_509;
wire n_510;
wire n_511;
wire n_512;
wire n_513;
wire n_514;
wire n_515;
wire n_516;
wire n_517;
wire n_518;
wire n_519;
wire n_520;
wire n_521;
wire n_522;
wire n_523;
wire n_524;
wire n_525;
wire n_526;
wire n_527;
wire n_528;
wire n_529;
wire n_530;
wire n_531;
wire n_532;
wire n_533;
wire n_534;
wire n_535;
wire n_536;
wire n_537;
wire n_538;
wire n_539;
wire n_540;
wire n_541;
wire n_542;
wire n_543;
wire n_544;
wire n_545;
wire n_546;
wire n_547;
wire n_548;
wire n_549;
wire n_550;
wire n_551;
wire n_552;
wire n_553;
wire n_554;
wire n_555;
wire n_556;
wire n_557;
wire n_558;
wire n_559;
wire n_560;
wire n_561;
wire n_562;
wire n_563;
wire n_564;
wire n_565;
wire n_566;
wire n_567;
wire n_568;
wire n_569;
wire n_570;
wire n_571;
wire n_572;
wire n_573;
wire n_574;
wire n_575;
wire n_576;
wire n_577;
wire n_578;
wire n_579;
wire n_580;
wire n_581;
wire n_582;
wire n_583;
wire n_584;
wire n_585;
wire n_586;
wire n_587;
wire n_588;
wire n_589;
wire n_590;
wire n_591;
wire n_592;
wire n_593;
wire n_594;
wire n_595;
wire n_596;
wire n_597;
wire n_598;
wire n_599;
wire n_600;
wire n_601;
wire n_602;
wire n_603;
wire n_604;
wire n_605;
wire n_606;
wire n_607;
wire n_608;
wire n_609;
wire n_610;
wire n_611;
wire n_612;
wire n_613;
wire n_614;
wire n_615;
wire n_616;
wire n_617;
wire n_618;
wire n_619;
wire n_620;
wire n_621;
wire n_622;
wire n_623;
wire n_624;
wire n_625;
wire n_626;
wire n_627;
wire n_628;
wire n_629;
wire n_630;
wire n_631;
wire n_632;
wire n_633;
wire n_634;
wire n_635;
wire n_636;
wire n_637;
wire n_638;
wire n_639;
wire n_640;
wire n_641;
wire n_642;
wire n_643;
wire n_644;
wire n_645;
wire n_646;
wire n_647;
wire n_648;
wire n_649;
wire n_650;
wire n_651;
wire n_652;
wire n_653;
wire n_654;
wire n_655;
wire n_656;
wire n_657;
wire n_658;
wire n_659;
wire n_660;
wire n_661;
wire n_662;
wire n_663;
wire n_664;
wire n_665;
wire n_666;
wire n_667;
wire n_668;
wire n_669;
wire n_670;
wire n_671;
wire n_672;
wire n_673;
wire n_674;
wire n_675;
wire n_676;
wire n_677;
wire n_678;
wire n_679;
wire n_680;
wire n_681;
wire n_682;
wire n_683;
wire n_684;
wire n_685;
wire n_686;
wire n_687;
wire n_688;
wire n_689;
wire n_690;
wire n_691;
wire n_692;
wire n_693;
wire n_694;
wire n_695;
wire n_696;
wire n_697;
wire n_698;
wire n_699;
wire n_700;
wire n_701;
wire n_702;
wire n_703;
wire n_704;
wire n_705;
wire n_706;
wire n_707;
wire n_708;
wire n_709;
wire n_710;
wire n_711;
wire n_712;
wire n_713;
wire n_714;
wire n_715;
wire n_716;
wire n_717;
wire n_718;
wire n_719;
wire n_720;
wire n_721;
wire n_722;
wire n_723;
wire n_724;
wire n_725;
wire n_726;
wire n_727;
wire n_728;
wire n_729;
wire n_730;
wire n_731;
wire n_732;
wire n_733;
wire n_734;
wire n_735;
wire n_736;
wire n_737;
wire n_738;
wire n_739;
wire n_740;
wire n_741;
wire n_742;
wire n_743;
wire n_744;
wire n_745;
wire n_746;
wire n_747;
wire n_748;
wire n_749;
wire n_750;
wire n_751;
wire n_752;
wire n_753;
wire n_754;
wire n_755;
wire n_756;
wire n_757;
wire n_758;
wire n_759;
wire n_760;
wire n_761;
wire n_762;
wire n_763;
wire n_764;
wire n_765;
wire n_766;
wire n_767;
wire n_768;
wire n_769;
wire n_770;
wire n_771;
wire n_772;
wire n_773;
wire n_774;
wire n_775;
wire n_776;
wire n_777;
wire n_778;
wire n_779;
wire n_780;
wire n_781;
wire n_782;
wire n_783;
wire n_784;
wire n_785;
wire n_786;
wire n_787;
wire n_788;
wire n_789;
wire n_790;
wire n_791;
wire n_792;
wire n_793;
wire n_794;
wire n_795;
wire n_796;
wire n_797;
wire n_798;
wire n_799;
wire n_800;
wire n_801;
wire n_802;
wire n_803;
wire n_804;
wire n_805;
wire n_806;
wire n_807;
wire n_808;
wire n_809;
wire n_810;
wire n_811;
wire n_812;
wire n_813;
wire n_814;
wire n_815;
wire n_816;
wire n_817;
wire n_818;
wire n_819;
wire n_820;
wire n_821;
wire n_822;
wire n_823;
wire n_824;
wire n_825;
wire n_826;
wire n_827;
wire n_828;
wire n_829;
wire n_830;
wire n_831;
wire n_832;
wire n_833;
wire n_834;
wire n_835;
wire n_836;
wire n_837;
wire n_838;
wire n_839;
wire n_840;
wire n_841;
wire n_842;
wire n_843;
wire n_844;
wire n_845;
wire n_846;
wire n_847;
wire n_848;
wire n_849;
wire n_850;
wire n_851;
wire n_852;
wire n_853;
wire n_854;
wire n_855;
wire n_856;
wire n_857;
wire n_858;
wire n_859;
wire n_860;
wire n_861;
wire n_862;
wire n_863;
wire n_864;
wire n_865;
wire n_866;
wire n_867;
wire n_868;
wire n_869;
wire n_870;
wire n_871;
wire n_872;
wire n_873;
wire n_874;
wire n_875;
wire n_876;
wire n_877;
wire n_878;
wire n_879;
wire n_880;
wire n_881;
wire n_882;
wire n_883;
wire n_884;
wire n_885;
wire n_886;
wire n_887;
wire n_888;
wire n_889;
wire n_890;
wire n_891;
wire n_892;
wire n_893;
wire n_894;
wire n_895;
wire n_896;
wire n_897;
wire n_898;
wire n_899;
wire n_900;
wire n_901;
wire n_902;
wire n_903;
wire n_904;
wire n_905;
wire n_906;
wire n_907;
wire n_908;
wire n_909;
wire n_910;
wire n_911;
wire n_912;
wire n_913;
wire n_914;
wire n_915;
wire n_916;
wire n_917;
wire n_918;
wire n_919;
wire n_920;
wire n_921;
wire n_922;
wire n_923;
wire n_924;
wire n_925;
wire n_926;
wire n_927;
wire n_928;
wire n_929;
wire n_930;
wire n_931;
wire n_932;
wire n_933;
wire n_934;
wire n_935;
wire n_936;
wire n_937;
wire n_938;
wire n_939;
wire n_940;
wire n_941;
wire n_942;
wire n_943;
wire n_944;
wire n_945;
wire n_946;
wire n_947;
wire n_948;
wire n_949;
wire n_950;
wire n_951;
wire n_952;
wire n_953;
wire n_954;
wire n_955;
wire n_956;
wire n_957;
wire n_958;
wire n_959;
wire n_960;
wire n_961;
wire n_962;
wire n_963;
wire n_964;
wire n_965;
wire n_966;
wire n_967;
wire n_968;
wire n_969;
wire n_970;
wire n_971;
wire n_972;
wire n_973;
wire n_974;
wire n_975;
wire n_976;
wire n_977;
wire n_978;
wire n_979;
wire n_980;
wire n_981;
wire n_982;
wire n_983;
wire n_984;
wire n_985;
wire n_986;
wire n_987;
wire n_988;
wire n_989;
wire n_990;
wire n_991;
wire n_992;
wire n_993;
wire n_994;
wire n_995;
wire n_996;
wire n_997;
wire n_998;
wire n_999;
wire n_1000;
wire n_1001;
wire n_1002;
wire n_1003;
wire n_1004;
wire n_1005;
wire n_1006;
wire n_1007;
wire n_1008;
wire n_1009;
wire n_1010;
wire n_1011;
wire n_1012;
wire n_1013;
wire n_1014;
wire n_1015;
wire n_1016;
wire n_1017;
wire n_1018;
wire n_1019;
wire n_1020;
wire n_1021;
wire n_1022;
wire n_1023;
wire n_1024;
wire n_1025;
wire n_1026;
wire n_1027;
wire n_1028;
wire n_1029;
wire n_1030;
wire n_1031;
wire n_1032;
wire n_1033;
wire n_1034;
wire n_1035;
wire n_1036;
wire n_1037;
wire n_1038;
wire n_1039;
wire n_1040;
wire n_1041;
wire n_1042;
wire n_1043;
wire n_1044;
wire n_1045;
wire n_1046;
wire n_1047;
wire n_1048;
wire n_1049;
wire n_1050;
wire n_1051;
wire n_1052;
wire n_1053;
wire n_1054;
wire n_1055;
wire n_1056;
wire n_1057;
wire n_1058;
wire n_1059;
wire n_1060;
wire n_1061;
wire n_1062;
wire n_1063;
wire n_1064;
wire n_1065;
wire n_1066;
wire n_1067;
wire n_1068;
wire n_1069;
wire n_1070;
wire n_1071;
wire n_1072;
wire n_1073;
wire n_1074;
wire n_1075;
wire n_1076;
wire n_1077;
wire n_1078;
wire n_1079;
wire n_1080;
wire n_1081;
wire n_1082;
wire n_1083;
wire n_1084;
wire n_1085;
wire n_1086;
wire n_1087;
wire n_1088;
wire n_1089;
wire n_1090;
wire n_1091;
wire n_1092;
wire n_1093;
wire n_1094;
wire n_1095;
wire n_1096;
wire n_1097;
wire n_1098;
wire n_1099;
wire n_1100;
wire n_1101;
wire n_1102;
wire n_1103;
wire n_1104;
wire n_1105;
wire n_1106;
wire n_1107;
wire n_1108;
wire n_1109;
wire n_1110;
wire n_1111;
wire n_1112;
wire n_1113;
wire n_1114;
wire n_1115;
wire n_1116;
wire n_1117;
wire n_1118;
wire n_1119;
wire n_1120;
wire n_1121;
wire n_1122;
wire n_1123;
wire n_1124;
wire n_1125;
wire n_1126;
wire n_1127;
wire n_1128;
wire n_1129;
wire n_1130;
wire n_1131;
wire n_1132;
wire n_1133;
wire n_1134;
wire n_1135;
wire n_1136;
wire n_1137;
wire n_1138;
wire n_1139;
wire n_1140;
wire n_1141;
wire n_1142;
wire n_1143;
wire n_1144;
wire n_1145;
wire n_1146;
wire n_1147;
wire n_1148;
wire n_1149;
wire n_1150;
wire n_1151;
wire n_1152;
wire n_1153;
wire n_1154;
wire n_1155;
wire n_1156;
wire n_1157;
wire n_1158;
wire n_1159;
wire n_1160;
wire n_1161;
wire n_1162;
wire n_1163;
wire n_1164;
wire n_1165;
wire n_1166;
wire n_1167;
wire n_1168;
wire n_1169;
wire n_1170;
wire n_1171;
wire n_1172;
wire n_1173;
wire n_1174;
wire n_1175;
wire n_1176;
wire n_1177;
wire n_1178;
wire n_1179;
wire n_1180;
wire n_1181;
wire n_1182;
wire n_1183;
wire n_1184;
wire n_1185;
wire n_1186;
wire n_1187;
wire n_1188;
wire n_1189;
wire n_1190;
wire n_1191;
wire n_1192;
wire n_1193;
wire n_1194;
wire n_1195;
wire n_1196;
wire n_1197;
wire n_1198;
wire n_1199;
wire n_1200;
wire n_1201;
wire n_1202;
wire n_1203;
wire n_1204;
wire n_1205;
wire n_1206;
wire n_1207;
wire n_1208;
wire n_1209;
wire n_1210;
wire n_1211;
wire n_1212;
wire n_1213;
wire n_1214;
wire n_1215;
wire n_1216;
wire n_1217;
wire n_1218;
wire n_1219;
wire n_1220;
wire n_1221;
wire n_1222;
wire n_1223;
wire n_1224;
wire n_1225;
wire n_1226;
wire n_1227;
wire n_1228;
wire n_1229;
wire n_1230;
wire n_1231;
wire n_1232;
wire n_1233;
wire n_1234;
wire n_1235;
wire n_1236;
wire n_1237;
wire n_1238;
wire n_1239;
wire n_1240;
wire n_1241;
wire n_1242;
wire n_1243;
wire n_1244;
wire n_1245;
wire n_1246;
wire n_1247;
wire n_1248;
wire n_1249;
wire n_1250;
wire n_1251;
wire n_1252;
wire n_1253;
wire n_1254;
wire n_1255;
wire n_1256;
wire n_1257;
wire n_1258;
wire n_1259;
wire n_1260;
wire n_1261;
wire n_1262;
wire n_1263;
wire n_1264;
wire n_1265;
wire n_1266;
wire n_1267;
wire n_1268;
wire n_1269;
wire n_1270;
wire n_1271;
wire n_1272;
wire n_1273;
wire n_1274;
wire n_1275;
wire n_1276;
wire n_1277;
wire n_1278;
wire n_1279;
wire n_1280;
wire n_1281;
wire n_1282;
wire n_1283;
wire n_1284;
wire n_1285;
wire n_1286;
wire n_1287;
wire n_1288;
wire n_1289;
wire n_1290;
wire n_1291;
wire n_1292;
wire n_1293;
wire n_1294;
wire n_1295;
wire n_1296;
wire n_1297;
wire n_1298;
wire n_1299;
wire n_1300;
wire n_1301;
wire n_1302;
wire n_1303;
wire n_1304;
wire n_1305;
wire n_1306;
wire n_1307;
wire n_1308;
wire n_1309;
wire n_1310;
wire n_1311;
wire n_1312;
wire n_1313;
wire n_1314;
wire n_1315;
wire n_1316;
wire n_1317;
wire n_1318;
wire n_1319;
wire n_1320;
wire n_1321;
wire n_1322;
wire n_1323;
wire n_1324;
wire n_1325;
wire n_1326;
wire n_1327;
wire n_1328;
wire n_1329;
wire n_1330;
wire n_1331;
wire n_1332;
wire n_1333;
wire n_1334;
wire n_1335;
wire n_1336;
wire n_1337;
wire n_1338;
wire n_1339;
wire n_1340;
wire n_1341;
wire n_1342;
wire n_1343;
wire n_1344;
wire n_1345;
wire n_1346;
wire n_1347;
wire n_1348;
wire n_1349;
wire n_1350;
wire n_1351;
wire n_1352;
wire n_1353;
wire n_1354;
wire n_1355;
wire n_1356;
wire n_1357;
wire n_1358;
wire n_1359;
wire n_1360;
wire n_1361;
wire n_1362;
wire n_1363;
wire n_1364;
wire n_1365;
wire n_1366;
wire n_1367;
wire n_1368;
wire n_1369;
wire n_1370;
wire n_1371;
wire n_1372;
wire n_1373;
wire n_1374;
wire n_1375;
wire n_1376;
wire n_1377;
wire n_1378;
wire n_1379;
wire n_1380;
wire n_1381;
wire n_1382;
wire n_1383;
wire n_1384;
wire n_1385;
wire n_1386;
wire n_1387;
wire n_1388;
wire n_1389;
wire n_1390;
wire n_1391;
wire n_1392;
wire n_1393;
wire n_1394;
wire n_1395;
wire n_1396;
wire n_1397;
wire n_1398;
wire n_1399;
wire n_1400;
wire n_1401;
wire n_1402;
wire n_1403;
wire n_1404;
wire n_1405;
wire n_1406;
wire n_1407;
wire n_1408;
wire n_1409;
wire n_1410;
wire n_1411;
wire n_1412;
wire n_1413;
wire n_1414;
wire n_1415;
wire n_1416;
wire n_1417;
wire n_1418;
wire n_1419;
wire n_1420;
wire n_1421;
wire n_1422;
wire n_1423;
assign n_1 = ~i_10 & ~i_29;
assign n_2 =  x_93 &  n_1;
assign n_3 =  i_29 &  x_85;
assign n_4 =  x_94 &  n_3;
assign n_5 =  x_93 &  n_4;
assign n_6 = ~x_93 & ~n_4;
assign n_7 = ~n_5 & ~n_6;
assign n_8 =  i_29 &  x_54;
assign n_9 =  n_7 &  n_8;
assign n_10 = ~n_2 & ~n_9;
assign n_11 =  x_93 & ~n_10;
assign n_12 = ~x_93 &  n_10;
assign n_13 = ~n_11 & ~n_12;
assign n_14 =  x_92 &  n_1;
assign n_15 =  x_92 &  n_5;
assign n_16 = ~x_92 & ~n_5;
assign n_17 = ~n_15 & ~n_16;
assign n_18 =  i_29 &  x_52;
assign n_19 =  n_17 &  n_18;
assign n_20 = ~n_14 & ~n_19;
assign n_21 =  x_92 & ~n_20;
assign n_22 = ~x_92 &  n_20;
assign n_23 = ~n_21 & ~n_22;
assign n_24 =  i_29 &  x_89;
assign n_25 =  x_98 &  n_24;
assign n_26 =  x_91 &  n_25;
assign n_27 = ~x_91 & ~n_25;
assign n_28 = ~n_26 & ~n_27;
assign n_29 =  i_29 &  x_73;
assign n_30 =  n_28 &  n_29;
assign n_31 = ~i_7 & ~i_29;
assign n_32 =  x_91 &  n_31;
assign n_33 = ~n_30 & ~n_32;
assign n_34 =  x_91 & ~n_33;
assign n_35 = ~x_91 &  n_33;
assign n_36 = ~n_34 & ~n_35;
assign n_37 =  x_90 &  n_26;
assign n_38 = ~x_90 & ~n_26;
assign n_39 = ~n_37 & ~n_38;
assign n_40 =  n_39 &  n_29;
assign n_41 =  x_90 &  n_31;
assign n_42 = ~n_40 & ~n_41;
assign n_43 =  x_90 & ~n_42;
assign n_44 = ~x_90 &  n_42;
assign n_45 = ~n_43 & ~n_44;
assign n_46 =  x_89 &  n_31;
assign n_47 =  x_73 & ~x_89;
assign n_48 =  x_74 & ~n_47;
assign n_49 =  i_29 & ~n_48;
assign n_50 = ~n_46 & ~n_49;
assign n_51 =  x_89 & ~n_50;
assign n_52 = ~x_89 &  n_50;
assign n_53 = ~n_51 & ~n_52;
assign n_54 =  x_88 &  n_37;
assign n_55 = ~x_88 & ~n_37;
assign n_56 = ~n_54 & ~n_55;
assign n_57 =  n_29 &  n_56;
assign n_58 =  x_88 &  n_31;
assign n_59 = ~n_57 & ~n_58;
assign n_60 =  x_88 & ~n_59;
assign n_61 = ~x_88 &  n_59;
assign n_62 = ~n_60 & ~n_61;
assign n_63 =  x_87 &  n_31;
assign n_64 =  x_87 &  n_54;
assign n_65 = ~x_87 & ~n_54;
assign n_66 = ~n_64 & ~n_65;
assign n_67 =  x_73 &  n_66;
assign n_68 =  i_29 &  n_67;
assign n_69 = ~n_63 & ~n_68;
assign n_70 =  x_87 & ~n_69;
assign n_71 = ~x_87 &  n_69;
assign n_72 = ~n_70 & ~n_71;
assign n_73 =  x_86 &  n_64;
assign n_74 = ~x_86 & ~n_64;
assign n_75 = ~n_73 & ~n_74;
assign n_76 =  n_75 &  n_29;
assign n_77 =  x_86 &  n_31;
assign n_78 = ~n_76 & ~n_77;
assign n_79 =  x_86 & ~n_78;
assign n_80 = ~x_86 &  n_78;
assign n_81 = ~n_79 & ~n_80;
assign n_82 =  x_69 & ~x_85;
assign n_83 = ~x_70 & ~n_82;
assign n_84 =  i_29 & ~n_83;
assign n_85 =  x_85 &  n_1;
assign n_86 = ~n_84 & ~n_85;
assign n_87 =  x_85 & ~n_86;
assign n_88 = ~x_85 &  n_86;
assign n_89 = ~n_87 & ~n_88;
assign n_90 =  i_29 &  x_59;
assign n_91 =  x_83 &  n_90;
assign n_92 =  x_81 &  x_82;
assign n_93 =  n_91 &  n_92;
assign n_94 =  x_80 &  n_93;
assign n_95 =  x_79 &  n_94;
assign n_96 = ~x_58 &  x_60;
assign n_97 = ~n_95 &  n_96;
assign n_98 =  x_78 &  n_97;
assign n_99 =  x_79 &  n_96;
assign n_100 =  n_94 &  n_99;
assign n_101 = ~x_78 &  n_100;
assign n_102 = ~x_62 & ~n_101;
assign n_103 = ~n_98 &  n_102;
assign n_104 =  x_100 & ~n_103;
assign n_105 = ~x_100 &  n_103;
assign n_106 = ~n_104 & ~n_105;
assign n_107 = ~x_80 & ~n_93;
assign n_108 = ~n_94 &  n_96;
assign n_109 = ~n_107 &  n_108;
assign n_110 = ~x_64 & ~n_109;
assign n_111 =  x_102 &  n_110;
assign n_112 =  n_91 &  n_96;
assign n_113 = ~x_82 &  n_112;
assign n_114 = ~n_91 &  n_96;
assign n_115 =  x_82 &  n_114;
assign n_116 = ~x_66 & ~n_115;
assign n_117 = ~n_113 &  n_116;
assign n_118 =  x_104 & ~n_117;
assign n_119 = ~x_104 &  n_117;
assign n_120 = ~n_118 & ~n_119;
assign n_121 = ~x_102 & ~n_110;
assign n_122 = ~n_120 & ~n_121;
assign n_123 = ~n_111 &  n_122;
assign n_124 = ~x_79 & ~n_94;
assign n_125 =  n_97 & ~n_124;
assign n_126 = ~x_63 & ~n_125;
assign n_127 = ~x_101 & ~n_126;
assign n_128 =  x_82 & ~n_93;
assign n_129 =  n_112 &  n_128;
assign n_130 =  x_81 &  n_96;
assign n_131 = ~n_93 &  n_130;
assign n_132 = ~x_65 & ~n_131;
assign n_133 = ~n_129 &  n_132;
assign n_134 = ~x_103 & ~n_133;
assign n_135 = ~x_83 & ~n_90;
assign n_136 =  n_114 & ~n_135;
assign n_137 = ~x_67 & ~n_136;
assign n_138 = ~x_105 & ~n_137;
assign n_139 =  x_105 &  n_137;
assign n_140 = ~n_138 & ~n_139;
assign n_141 = ~n_134 &  n_140;
assign n_142 =  x_103 &  n_133;
assign n_143 = ~i_28 & ~x_111;
assign n_144 =  i_28 &  x_111;
assign n_145 = ~n_143 & ~n_144;
assign n_146 = ~x_58 & ~x_60;
assign n_147 =  n_145 &  n_146;
assign n_148 = ~i_29 & ~x_59;
assign n_149 = ~n_90 &  n_96;
assign n_150 = ~n_148 &  n_149;
assign n_151 = ~x_68 & ~n_150;
assign n_152 = ~n_147 &  n_151;
assign n_153 =  x_106 & ~n_152;
assign n_154 = ~x_106 &  n_152;
assign n_155 = ~n_153 & ~n_154;
assign n_156 = ~n_142 & ~n_155;
assign n_157 =  n_141 &  n_156;
assign n_158 = ~n_127 &  n_157;
assign n_159 =  n_123 &  n_158;
assign n_160 = ~n_106 &  n_159;
assign n_161 =  x_35 &  n_73;
assign n_162 = ~x_35 & ~n_73;
assign n_163 = ~n_161 & ~n_162;
assign n_164 = ~x_98 & ~n_24;
assign n_165 = ~n_25 & ~n_164;
assign n_166 = ~i_29 & ~x_89;
assign n_167 =  x_98 & ~n_166;
assign n_168 =  x_74 & ~n_167;
assign n_169 =  x_88 & ~n_168;
assign n_170 =  n_165 &  n_169;
assign n_171 =  n_28 &  n_170;
assign n_172 =  n_39 &  n_171;
assign n_173 =  n_67 &  n_172;
assign n_174 =  n_75 &  n_173;
assign n_175 =  n_163 &  n_174;
assign n_176 =  x_101 &  n_126;
assign n_177 =  x_33 &  x_78;
assign n_178 =  n_95 &  n_177;
assign n_179 =  x_33 &  n_96;
assign n_180 = ~n_178 &  n_179;
assign n_181 = ~x_33 &  x_78;
assign n_182 =  n_100 &  n_181;
assign n_183 = ~x_61 & ~n_182;
assign n_184 = ~n_180 &  n_183;
assign n_185 = ~x_99 & ~n_184;
assign n_186 =  x_99 &  n_184;
assign n_187 = ~n_185 & ~n_186;
assign n_188 = ~n_176 &  n_187;
assign n_189 =  n_175 &  n_188;
assign n_190 =  n_160 &  n_189;
assign n_191 =  x_32 &  n_190;
assign n_192 = ~x_107 & ~n_191;
assign n_193 =  x_77 & ~n_175;
assign n_194 = ~x_108 & ~n_193;
assign n_195 =  x_97 &  n_15;
assign n_196 =  x_95 &  n_195;
assign n_197 =  x_96 &  n_196;
assign n_198 =  x_45 &  n_197;
assign n_199 = ~x_45 & ~n_197;
assign n_200 = ~n_198 & ~n_199;
assign n_201 = ~x_95 & ~n_195;
assign n_202 = ~n_196 & ~n_201;
assign n_203 =  x_48 &  n_202;
assign n_204 = ~x_96 & ~n_196;
assign n_205 = ~n_197 & ~n_204;
assign n_206 = ~x_97 & ~n_15;
assign n_207 = ~n_195 & ~n_206;
assign n_208 = ~x_94 & ~n_3;
assign n_209 = ~n_4 & ~n_208;
assign n_210 =  x_70 &  n_209;
assign n_211 =  i_29 & ~x_85;
assign n_212 = ~i_29 &  x_85;
assign n_213 = ~n_211 & ~n_212;
assign n_214 =  x_69 &  x_94;
assign n_215 = ~n_213 &  n_214;
assign n_216 = ~n_210 & ~n_215;
assign n_217 =  x_54 &  x_56;
assign n_218 =  x_92 & ~x_108;
assign n_219 =  n_217 &  n_218;
assign n_220 =  x_43 &  x_46;
assign n_221 =  x_50 &  x_52;
assign n_222 =  n_220 &  n_221;
assign n_223 =  n_219 &  n_222;
assign n_224 =  n_7 &  n_223;
assign n_225 = ~n_216 &  n_224;
assign n_226 =  n_207 &  n_225;
assign n_227 =  n_205 &  n_226;
assign n_228 =  n_203 &  n_227;
assign n_229 =  n_200 &  n_228;
assign n_230 = ~n_194 & ~n_229;
assign n_231 =  x_77 & ~n_190;
assign n_232 = ~x_30 & ~x_31;
assign n_233 = ~n_231 &  n_232;
assign n_234 = ~n_230 &  n_233;
assign n_235 = ~n_192 &  n_234;
assign n_236 =  x_84 &  n_235;
assign n_237 = ~x_84 & ~n_235;
assign n_238 = ~n_236 & ~n_237;
assign n_239 =  i_29 & ~n_137;
assign n_240 = ~i_9 & ~i_29;
assign n_241 =  x_83 &  n_240;
assign n_242 = ~n_239 & ~n_241;
assign n_243 =  x_83 & ~n_242;
assign n_244 = ~x_83 &  n_242;
assign n_245 = ~n_243 & ~n_244;
assign n_246 =  i_29 & ~n_117;
assign n_247 =  x_82 &  n_240;
assign n_248 = ~n_246 & ~n_247;
assign n_249 =  x_82 & ~n_248;
assign n_250 = ~x_82 &  n_248;
assign n_251 = ~n_249 & ~n_250;
assign n_252 =  i_29 & ~n_133;
assign n_253 =  x_81 &  n_240;
assign n_254 = ~n_252 & ~n_253;
assign n_255 =  x_81 & ~n_254;
assign n_256 = ~x_81 &  n_254;
assign n_257 = ~n_255 & ~n_256;
assign n_258 =  i_29 & ~n_110;
assign n_259 =  x_80 &  n_240;
assign n_260 = ~n_258 & ~n_259;
assign n_261 =  x_80 & ~n_260;
assign n_262 = ~x_80 &  n_260;
assign n_263 = ~n_261 & ~n_262;
assign n_264 =  i_29 & ~n_126;
assign n_265 =  x_79 &  n_240;
assign n_266 = ~n_264 & ~n_265;
assign n_267 =  x_79 & ~n_266;
assign n_268 = ~x_79 &  n_266;
assign n_269 = ~n_267 & ~n_268;
assign n_270 =  i_29 & ~n_103;
assign n_271 =  x_78 &  n_240;
assign n_272 = ~n_270 & ~n_271;
assign n_273 =  x_78 & ~n_272;
assign n_274 = ~x_78 &  n_272;
assign n_275 = ~n_273 & ~n_274;
assign n_276 =  n_192 &  n_230;
assign n_277 =  x_77 &  n_276;
assign n_278 = ~x_77 & ~n_276;
assign n_279 = ~n_277 & ~n_278;
assign n_280 =  n_233 &  n_276;
assign n_281 =  x_76 &  n_280;
assign n_282 = ~x_76 & ~n_280;
assign n_283 = ~n_281 & ~n_282;
assign n_284 = ~n_233 &  n_276;
assign n_285 = ~i_2 & ~i_25;
assign n_286 =  x_111 &  n_285;
assign n_287 =  i_23 &  i_25;
assign n_288 = ~n_286 & ~n_287;
assign n_289 = ~i_8 & ~i_29;
assign n_290 =  x_112 &  n_289;
assign n_291 =  i_29 &  x_111;
assign n_292 = ~n_290 & ~n_291;
assign n_293 =  n_288 & ~n_292;
assign n_294 = ~n_288 &  n_292;
assign n_295 = ~n_293 & ~n_294;
assign n_296 =  n_284 &  n_295;
assign n_297 =  x_75 &  n_296;
assign n_298 = ~x_75 & ~n_296;
assign n_299 = ~n_297 & ~n_298;
assign n_300 = ~n_284 & ~n_235;
assign n_301 =  n_300 &  n_288;
assign n_302 =  x_74 & ~n_301;
assign n_303 = ~x_74 &  n_301;
assign n_304 = ~n_302 & ~n_303;
assign n_305 = ~n_300 &  n_288;
assign n_306 =  x_73 &  n_305;
assign n_307 = ~x_73 & ~n_305;
assign n_308 = ~n_306 & ~n_307;
assign n_309 = ~n_300 & ~n_288;
assign n_310 =  x_72 &  n_309;
assign n_311 = ~x_72 & ~n_309;
assign n_312 = ~n_310 & ~n_311;
assign n_313 =  x_71 &  n_309;
assign n_314 = ~x_71 & ~n_309;
assign n_315 = ~n_313 & ~n_314;
assign n_316 =  n_300 & ~n_288;
assign n_317 =  x_70 &  n_316;
assign n_318 = ~x_70 & ~n_316;
assign n_319 = ~n_317 & ~n_318;
assign n_320 =  x_69 &  n_309;
assign n_321 = ~x_69 & ~n_309;
assign n_322 = ~n_320 & ~n_321;
assign n_323 = ~n_300 &  n_295;
assign n_324 =  i_29 & ~n_152;
assign n_325 =  x_59 &  n_240;
assign n_326 = ~n_324 & ~n_325;
assign n_327 =  n_323 & ~n_326;
assign n_328 =  x_68 &  n_327;
assign n_329 = ~x_68 & ~n_327;
assign n_330 = ~n_328 & ~n_329;
assign n_331 =  n_323 & ~n_242;
assign n_332 =  x_67 &  n_331;
assign n_333 = ~x_67 & ~n_331;
assign n_334 = ~n_332 & ~n_333;
assign n_335 =  n_323 & ~n_248;
assign n_336 =  x_66 &  n_335;
assign n_337 = ~x_66 & ~n_335;
assign n_338 = ~n_336 & ~n_337;
assign n_339 =  n_323 & ~n_254;
assign n_340 =  x_65 &  n_339;
assign n_341 = ~x_65 & ~n_339;
assign n_342 = ~n_340 & ~n_341;
assign n_343 =  n_323 & ~n_260;
assign n_344 =  x_64 &  n_343;
assign n_345 = ~x_64 & ~n_343;
assign n_346 = ~n_344 & ~n_345;
assign n_347 =  n_323 & ~n_266;
assign n_348 =  x_63 &  n_347;
assign n_349 = ~x_63 & ~n_347;
assign n_350 = ~n_348 & ~n_349;
assign n_351 =  x_132 & ~x_133;
assign n_352 = ~x_131 & ~x_132;
assign n_353 =  x_133 &  n_352;
assign n_354 =  x_131 &  n_351;
assign n_355 = ~n_353 & ~n_354;
assign n_356 = ~x_174 & ~x_186;
assign n_357 =  x_174 &  x_186;
assign n_358 = ~n_356 & ~n_357;
assign n_359 = ~n_355 & ~n_358;
assign n_360 =  x_175 &  n_359;
assign n_361 =  i_29 &  x_182;
assign n_362 =  x_181 &  n_361;
assign n_363 =  x_180 &  n_362;
assign n_364 =  x_179 &  n_363;
assign n_365 =  x_178 &  n_364;
assign n_366 =  x_177 &  n_365;
assign n_367 =  x_176 &  n_366;
assign n_368 = ~x_175 & ~n_367;
assign n_369 = ~n_355 &  n_358;
assign n_370 =  x_175 &  n_367;
assign n_371 =  n_369 & ~n_370;
assign n_372 = ~n_368 &  n_371;
assign n_373 = ~n_360 & ~n_372;
assign n_374 =  n_351 & ~n_373;
assign n_375 = ~i_5 & ~n_351;
assign n_376 =  x_134 &  n_375;
assign n_377 = ~n_374 & ~n_376;
assign n_378 =  x_134 & ~n_377;
assign n_379 = ~x_134 &  n_377;
assign n_380 = ~n_378 & ~n_379;
assign n_381 = ~x_187 &  n_352;
assign n_382 =  x_133 & ~n_381;
assign n_383 =  x_177 &  n_359;
assign n_384 = ~x_177 & ~n_365;
assign n_385 = ~n_366 &  n_369;
assign n_386 = ~n_384 &  n_385;
assign n_387 = ~n_383 & ~n_386;
assign n_388 = ~x_152 &  n_387;
assign n_389 =  x_152 & ~n_387;
assign n_390 = ~n_388 & ~n_389;
assign n_391 =  x_179 &  n_359;
assign n_392 = ~x_179 & ~n_363;
assign n_393 = ~n_364 &  n_369;
assign n_394 = ~n_392 &  n_393;
assign n_395 = ~n_391 & ~n_394;
assign n_396 =  x_154 &  n_395;
assign n_397 = ~i_29 & ~x_182;
assign n_398 = ~n_361 & ~n_397;
assign n_399 =  n_369 & ~n_398;
assign n_400 = ~i_28 & ~x_186;
assign n_401 =  i_28 &  x_186;
assign n_402 = ~n_400 & ~n_401;
assign n_403 =  n_355 & ~n_402;
assign n_404 = ~x_182 &  n_359;
assign n_405 = ~n_403 & ~n_404;
assign n_406 = ~n_399 &  n_405;
assign n_407 =  x_157 & ~n_406;
assign n_408 = ~n_396 & ~n_407;
assign n_409 = ~x_157 &  n_406;
assign n_410 =  x_180 &  n_359;
assign n_411 = ~x_180 & ~n_362;
assign n_412 = ~n_363 & ~n_411;
assign n_413 =  n_369 &  n_412;
assign n_414 = ~n_410 & ~n_413;
assign n_415 =  x_155 & ~n_414;
assign n_416 = ~x_155 &  n_414;
assign n_417 = ~n_415 & ~n_416;
assign n_418 = ~n_409 & ~n_417;
assign n_419 =  n_408 &  n_418;
assign n_420 =  x_178 &  n_359;
assign n_421 = ~x_178 & ~n_364;
assign n_422 = ~n_365 &  n_369;
assign n_423 = ~n_421 &  n_422;
assign n_424 = ~n_420 & ~n_423;
assign n_425 =  x_153 &  n_424;
assign n_426 = ~x_153 & ~n_424;
assign n_427 =  x_181 &  n_359;
assign n_428 = ~x_181 & ~n_361;
assign n_429 = ~n_362 & ~n_428;
assign n_430 =  n_369 &  n_429;
assign n_431 = ~n_427 & ~n_430;
assign n_432 =  x_156 & ~n_431;
assign n_433 = ~x_156 &  n_431;
assign n_434 = ~n_432 & ~n_433;
assign n_435 = ~x_154 & ~n_395;
assign n_436 = ~n_434 & ~n_435;
assign n_437 = ~n_426 &  n_436;
assign n_438 = ~n_425 &  n_437;
assign n_439 =  n_419 &  n_438;
assign n_440 = ~n_390 &  n_439;
assign n_441 =  x_150 &  n_373;
assign n_442 =  x_176 &  n_359;
assign n_443 = ~x_176 & ~n_366;
assign n_444 =  n_369 & ~n_367;
assign n_445 = ~n_443 &  n_444;
assign n_446 = ~n_442 & ~n_445;
assign n_447 = ~x_151 &  n_446;
assign n_448 =  x_151 & ~n_446;
assign n_449 = ~n_447 & ~n_448;
assign n_450 = ~x_150 & ~n_373;
assign n_451 = ~n_449 & ~n_450;
assign n_452 = ~n_441 &  n_451;
assign n_453 =  n_440 &  n_452;
assign n_454 = ~x_186 & ~n_355;
assign n_455 =  i_29 &  x_165;
assign n_456 =  x_164 &  n_455;
assign n_457 =  x_163 &  n_456;
assign n_458 =  x_162 &  n_457;
assign n_459 =  x_161 &  n_458;
assign n_460 =  x_160 &  n_459;
assign n_461 =  x_159 &  n_460;
assign n_462 =  x_158 &  n_461;
assign n_463 = ~x_158 & ~n_461;
assign n_464 = ~n_462 & ~n_463;
assign n_465 =  n_454 &  n_464;
assign n_466 = ~x_159 & ~n_460;
assign n_467 = ~n_461 & ~n_466;
assign n_468 =  n_454 &  n_467;
assign n_469 = ~x_161 & ~n_458;
assign n_470 = ~n_459 & ~n_469;
assign n_471 =  n_454 &  n_470;
assign n_472 = ~x_162 & ~n_457;
assign n_473 = ~n_458 & ~n_472;
assign n_474 =  n_454 &  n_473;
assign n_475 = ~i_29 & ~x_165;
assign n_476 = ~n_455 & ~n_475;
assign n_477 = ~n_355 & ~n_476;
assign n_478 = ~x_186 & ~n_477;
assign n_479 = ~x_164 & ~n_455;
assign n_480 = ~n_456 & ~n_479;
assign n_481 =  n_454 &  n_480;
assign n_482 =  x_160 &  x_163;
assign n_483 =  n_481 &  n_482;
assign n_484 =  n_478 &  n_483;
assign n_485 =  n_474 &  n_484;
assign n_486 =  n_471 &  n_485;
assign n_487 =  n_468 &  n_486;
assign n_488 =  n_465 &  n_487;
assign n_489 =  x_132 &  n_488;
assign n_490 =  n_453 &  n_489;
assign n_491 = ~n_382 & ~n_490;
assign n_492 =  x_133 & ~n_491;
assign n_493 = ~x_133 &  n_491;
assign n_494 = ~n_492 & ~n_493;
assign n_495 =  x_131 & ~x_132;
assign n_496 = ~x_133 &  n_495;
assign n_497 =  x_185 &  n_496;
assign n_498 =  n_351 & ~n_488;
assign n_499 =  i_29 &  x_173;
assign n_500 =  x_172 &  n_499;
assign n_501 =  x_171 &  n_500;
assign n_502 =  x_170 &  n_501;
assign n_503 =  x_169 &  n_502;
assign n_504 =  x_168 &  n_503;
assign n_505 =  x_167 &  n_504;
assign n_506 = ~x_166 & ~n_505;
assign n_507 =  x_166 &  n_505;
assign n_508 =  x_186 & ~n_355;
assign n_509 = ~n_507 &  n_508;
assign n_510 = ~n_506 &  n_509;
assign n_511 = ~x_167 & ~n_504;
assign n_512 = ~n_505 &  n_508;
assign n_513 = ~n_511 &  n_512;
assign n_514 = ~x_168 & ~n_503;
assign n_515 = ~n_504 &  n_508;
assign n_516 = ~n_514 &  n_515;
assign n_517 = ~x_169 & ~n_502;
assign n_518 = ~n_503 &  n_508;
assign n_519 = ~n_517 &  n_518;
assign n_520 = ~x_170 & ~n_501;
assign n_521 = ~n_502 &  n_508;
assign n_522 = ~n_520 &  n_521;
assign n_523 = ~i_29 & ~x_173;
assign n_524 = ~n_499 & ~n_523;
assign n_525 = ~n_355 & ~n_524;
assign n_526 = ~x_172 & ~n_499;
assign n_527 = ~n_500 & ~n_526;
assign n_528 =  x_171 &  x_186;
assign n_529 =  n_527 &  n_528;
assign n_530 = ~n_525 &  n_529;
assign n_531 =  n_522 &  n_530;
assign n_532 =  n_519 &  n_531;
assign n_533 =  n_516 &  n_532;
assign n_534 =  n_513 &  n_533;
assign n_535 =  n_510 &  n_534;
assign n_536 =  n_498 & ~n_535;
assign n_537 = ~n_497 & ~n_536;
assign n_538 =  x_132 & ~n_537;
assign n_539 = ~x_132 &  n_537;
assign n_540 = ~n_538 & ~n_539;
assign n_541 =  n_351 & ~n_453;
assign n_542 = ~x_133 &  x_187;
assign n_543 =  n_352 &  n_542;
assign n_544 = ~x_185 &  n_496;
assign n_545 = ~n_543 & ~n_544;
assign n_546 = ~n_498 &  n_545;
assign n_547 = ~n_541 &  n_546;
assign n_548 =  x_131 & ~n_547;
assign n_549 = ~x_131 &  n_547;
assign n_550 = ~n_548 & ~n_549;
assign n_551 =  i_22 &  i_26;
assign n_552 = ~i_3 & ~i_26;
assign n_553 =  x_187 &  n_552;
assign n_554 = ~n_551 & ~n_553;
assign n_555 =  x_187 & ~n_554;
assign n_556 = ~x_187 &  n_554;
assign n_557 = ~n_555 & ~n_556;
assign n_558 =  x_186 &  n_285;
assign n_559 = ~n_287 & ~n_558;
assign n_560 =  x_186 & ~n_559;
assign n_561 = ~x_186 &  n_559;
assign n_562 = ~n_560 & ~n_561;
assign n_563 =  i_21 &  i_24;
assign n_564 = ~i_1 & ~i_24;
assign n_565 =  x_185 &  n_564;
assign n_566 = ~n_563 & ~n_565;
assign n_567 =  x_185 & ~n_566;
assign n_568 = ~x_185 &  n_566;
assign n_569 = ~n_567 & ~n_568;
assign n_570 = ~i_28 & ~n_353;
assign n_571 =  i_29 & ~n_570;
assign n_572 = ~i_12 & ~i_29;
assign n_573 =  x_184 &  n_572;
assign n_574 = ~n_571 & ~n_573;
assign n_575 =  x_184 & ~n_574;
assign n_576 = ~x_184 &  n_574;
assign n_577 = ~n_575 & ~n_576;
assign n_578 = ~x_131 &  n_402;
assign n_579 =  x_131 &  n_358;
assign n_580 =  i_29 &  n_351;
assign n_581 = ~n_579 &  n_580;
assign n_582 = ~n_578 &  n_581;
assign n_583 = ~i_11 & ~i_29;
assign n_584 =  x_183 &  n_583;
assign n_585 = ~n_582 & ~n_584;
assign n_586 =  x_183 & ~n_585;
assign n_587 = ~x_183 &  n_585;
assign n_588 = ~n_586 & ~n_587;
assign n_589 =  i_29 &  n_406;
assign n_590 =  x_182 &  n_240;
assign n_591 = ~n_589 & ~n_590;
assign n_592 =  x_182 & ~n_591;
assign n_593 = ~x_182 &  n_591;
assign n_594 = ~n_592 & ~n_593;
assign n_595 =  i_29 & ~n_431;
assign n_596 =  x_181 &  n_240;
assign n_597 = ~n_595 & ~n_596;
assign n_598 =  x_181 & ~n_597;
assign n_599 = ~x_181 &  n_597;
assign n_600 = ~n_598 & ~n_599;
assign n_601 =  i_29 & ~n_414;
assign n_602 =  x_180 &  n_240;
assign n_603 = ~n_601 & ~n_602;
assign n_604 =  x_180 & ~n_603;
assign n_605 = ~x_180 &  n_603;
assign n_606 = ~n_604 & ~n_605;
assign n_607 =  i_29 & ~n_395;
assign n_608 =  x_179 &  n_240;
assign n_609 = ~n_607 & ~n_608;
assign n_610 =  x_179 & ~n_609;
assign n_611 = ~x_179 &  n_609;
assign n_612 = ~n_610 & ~n_611;
assign n_613 =  i_29 & ~n_424;
assign n_614 =  x_178 &  n_240;
assign n_615 = ~n_613 & ~n_614;
assign n_616 =  x_178 & ~n_615;
assign n_617 = ~x_178 &  n_615;
assign n_618 = ~n_616 & ~n_617;
assign n_619 =  i_29 & ~n_387;
assign n_620 =  x_177 &  n_240;
assign n_621 = ~n_619 & ~n_620;
assign n_622 =  x_177 & ~n_621;
assign n_623 = ~x_177 &  n_621;
assign n_624 = ~n_622 & ~n_623;
assign n_625 =  i_29 & ~n_446;
assign n_626 =  x_176 &  n_240;
assign n_627 = ~n_625 & ~n_626;
assign n_628 =  x_176 & ~n_627;
assign n_629 = ~x_176 &  n_627;
assign n_630 = ~n_628 & ~n_629;
assign n_631 =  i_29 & ~n_373;
assign n_632 =  x_175 &  n_240;
assign n_633 = ~n_631 & ~n_632;
assign n_634 =  x_175 & ~n_633;
assign n_635 = ~x_175 &  n_633;
assign n_636 = ~n_634 & ~n_635;
assign n_637 =  i_29 &  x_186;
assign n_638 =  x_174 &  n_289;
assign n_639 = ~n_637 & ~n_638;
assign n_640 =  x_174 & ~n_639;
assign n_641 = ~x_174 &  n_639;
assign n_642 = ~n_640 & ~n_641;
assign n_643 = ~n_525 &  n_637;
assign n_644 =  x_173 &  n_1;
assign n_645 = ~n_643 & ~n_644;
assign n_646 =  x_173 & ~n_645;
assign n_647 = ~x_173 &  n_645;
assign n_648 = ~n_646 & ~n_647;
assign n_649 =  n_508 &  n_527;
assign n_650 =  i_29 &  n_649;
assign n_651 =  x_172 &  n_1;
assign n_652 = ~n_650 & ~n_651;
assign n_653 =  x_172 & ~n_652;
assign n_654 = ~x_172 &  n_652;
assign n_655 = ~n_653 & ~n_654;
assign n_656 = ~x_171 & ~n_500;
assign n_657 = ~n_501 & ~n_656;
assign n_658 =  n_508 &  n_657;
assign n_659 =  i_29 &  n_658;
assign n_660 =  x_171 &  n_1;
assign n_661 = ~n_659 & ~n_660;
assign n_662 =  x_171 & ~n_661;
assign n_663 = ~x_171 &  n_661;
assign n_664 = ~n_662 & ~n_663;
assign n_665 =  i_29 &  n_522;
assign n_666 =  x_170 &  n_1;
assign n_667 = ~n_665 & ~n_666;
assign n_668 =  x_170 & ~n_667;
assign n_669 = ~x_170 &  n_667;
assign n_670 = ~n_668 & ~n_669;
assign n_671 =  i_29 &  n_519;
assign n_672 =  x_169 &  n_1;
assign n_673 = ~n_671 & ~n_672;
assign n_674 =  x_169 & ~n_673;
assign n_675 = ~x_169 &  n_673;
assign n_676 = ~n_674 & ~n_675;
assign n_677 =  i_29 &  n_516;
assign n_678 =  x_168 &  n_1;
assign n_679 = ~n_677 & ~n_678;
assign n_680 =  x_168 & ~n_679;
assign n_681 = ~x_168 &  n_679;
assign n_682 = ~n_680 & ~n_681;
assign n_683 =  i_29 &  n_513;
assign n_684 =  x_167 &  n_1;
assign n_685 = ~n_683 & ~n_684;
assign n_686 =  x_167 & ~n_685;
assign n_687 = ~x_167 &  n_685;
assign n_688 = ~n_686 & ~n_687;
assign n_689 =  i_29 &  n_510;
assign n_690 =  x_166 &  n_1;
assign n_691 = ~n_689 & ~n_690;
assign n_692 =  x_166 & ~n_691;
assign n_693 = ~x_166 &  n_691;
assign n_694 = ~n_692 & ~n_693;
assign n_695 =  i_29 &  n_478;
assign n_696 =  x_165 &  n_31;
assign n_697 = ~n_695 & ~n_696;
assign n_698 =  x_165 & ~n_697;
assign n_699 = ~x_165 &  n_697;
assign n_700 = ~n_698 & ~n_699;
assign n_701 =  x_164 &  n_31;
assign n_702 =  i_29 &  n_481;
assign n_703 = ~n_701 & ~n_702;
assign n_704 =  x_164 & ~n_703;
assign n_705 = ~x_164 &  n_703;
assign n_706 = ~n_704 & ~n_705;
assign n_707 = ~x_163 & ~n_456;
assign n_708 = ~n_457 & ~n_707;
assign n_709 =  i_29 &  n_454;
assign n_710 =  n_708 &  n_709;
assign n_711 =  x_163 &  n_31;
assign n_712 = ~n_710 & ~n_711;
assign n_713 =  x_163 & ~n_712;
assign n_714 = ~x_163 &  n_712;
assign n_715 = ~n_713 & ~n_714;
assign n_716 =  x_162 &  n_31;
assign n_717 =  i_29 &  n_474;
assign n_718 = ~n_716 & ~n_717;
assign n_719 =  x_162 & ~n_718;
assign n_720 = ~x_162 &  n_718;
assign n_721 = ~n_719 & ~n_720;
assign n_722 =  x_161 &  n_31;
assign n_723 =  i_29 &  n_471;
assign n_724 = ~n_722 & ~n_723;
assign n_725 =  x_161 & ~n_724;
assign n_726 = ~x_161 &  n_724;
assign n_727 = ~n_725 & ~n_726;
assign n_728 = ~x_160 & ~n_459;
assign n_729 = ~n_460 & ~n_728;
assign n_730 =  n_729 &  n_709;
assign n_731 =  x_160 &  n_31;
assign n_732 = ~n_730 & ~n_731;
assign n_733 =  x_160 & ~n_732;
assign n_734 = ~x_160 &  n_732;
assign n_735 = ~n_733 & ~n_734;
assign n_736 =  x_159 &  n_31;
assign n_737 =  i_29 &  n_468;
assign n_738 = ~n_736 & ~n_737;
assign n_739 =  x_159 & ~n_738;
assign n_740 = ~x_159 &  n_738;
assign n_741 = ~n_739 & ~n_740;
assign n_742 =  x_158 &  n_31;
assign n_743 =  i_29 &  n_465;
assign n_744 = ~n_742 & ~n_743;
assign n_745 =  x_158 & ~n_744;
assign n_746 = ~x_158 &  n_744;
assign n_747 = ~n_745 & ~n_746;
assign n_748 =  i_20 &  i_27;
assign n_749 = ~i_4 & ~i_27;
assign n_750 =  x_157 &  n_749;
assign n_751 = ~n_748 & ~n_750;
assign n_752 =  x_157 & ~n_751;
assign n_753 = ~x_157 &  n_751;
assign n_754 = ~n_752 & ~n_753;
assign n_755 =  i_19 &  i_27;
assign n_756 =  x_156 &  n_749;
assign n_757 = ~n_755 & ~n_756;
assign n_758 =  x_156 & ~n_757;
assign n_759 = ~x_156 &  n_757;
assign n_760 = ~n_758 & ~n_759;
assign n_761 =  i_18 &  i_27;
assign n_762 =  x_155 &  n_749;
assign n_763 = ~n_761 & ~n_762;
assign n_764 =  x_155 & ~n_763;
assign n_765 = ~x_155 &  n_763;
assign n_766 = ~n_764 & ~n_765;
assign n_767 =  i_17 &  i_27;
assign n_768 =  x_154 &  n_749;
assign n_769 = ~n_767 & ~n_768;
assign n_770 =  x_154 & ~n_769;
assign n_771 = ~x_154 &  n_769;
assign n_772 = ~n_770 & ~n_771;
assign n_773 =  i_16 &  i_27;
assign n_774 =  x_153 &  n_749;
assign n_775 = ~n_773 & ~n_774;
assign n_776 =  x_153 & ~n_775;
assign n_777 = ~x_153 &  n_775;
assign n_778 = ~n_776 & ~n_777;
assign n_779 =  i_15 &  i_27;
assign n_780 =  x_152 &  n_749;
assign n_781 = ~n_779 & ~n_780;
assign n_782 =  x_152 & ~n_781;
assign n_783 = ~x_152 &  n_781;
assign n_784 = ~n_782 & ~n_783;
assign n_785 =  i_14 &  i_27;
assign n_786 =  x_151 &  n_749;
assign n_787 = ~n_785 & ~n_786;
assign n_788 =  x_151 & ~n_787;
assign n_789 = ~x_151 &  n_787;
assign n_790 = ~n_788 & ~n_789;
assign n_791 =  i_13 &  i_27;
assign n_792 =  x_150 &  n_749;
assign n_793 = ~n_791 & ~n_792;
assign n_794 =  x_150 & ~n_793;
assign n_795 = ~x_150 &  n_793;
assign n_796 = ~n_794 & ~n_795;
assign n_797 = ~i_6 & ~n_351;
assign n_798 =  x_149 &  n_797;
assign n_799 =  n_508 & ~n_524;
assign n_800 = ~x_186 &  n_354;
assign n_801 = ~n_476 &  n_800;
assign n_802 =  n_351 & ~n_801;
assign n_803 = ~n_799 &  n_802;
assign n_804 = ~n_798 & ~n_803;
assign n_805 =  x_149 & ~n_804;
assign n_806 = ~x_149 &  n_804;
assign n_807 = ~n_805 & ~n_806;
assign n_808 =  n_480 &  n_800;
assign n_809 = ~n_649 & ~n_808;
assign n_810 =  n_351 & ~n_809;
assign n_811 =  x_148 &  n_797;
assign n_812 = ~n_810 & ~n_811;
assign n_813 =  x_148 & ~n_812;
assign n_814 = ~x_148 &  n_812;
assign n_815 = ~n_813 & ~n_814;
assign n_816 =  n_800 &  n_708;
assign n_817 = ~n_816 & ~n_658;
assign n_818 =  n_351 & ~n_817;
assign n_819 =  x_147 &  n_797;
assign n_820 = ~n_818 & ~n_819;
assign n_821 =  x_147 & ~n_820;
assign n_822 = ~x_147 &  n_820;
assign n_823 = ~n_821 & ~n_822;
assign n_824 =  n_473 &  n_800;
assign n_825 = ~n_522 & ~n_824;
assign n_826 =  n_351 & ~n_825;
assign n_827 =  x_146 &  n_797;
assign n_828 = ~n_826 & ~n_827;
assign n_829 =  x_146 & ~n_828;
assign n_830 = ~x_146 &  n_828;
assign n_831 = ~n_829 & ~n_830;
assign n_832 =  n_470 &  n_800;
assign n_833 = ~n_519 & ~n_832;
assign n_834 =  n_351 & ~n_833;
assign n_835 =  x_145 &  n_797;
assign n_836 = ~n_834 & ~n_835;
assign n_837 =  x_145 & ~n_836;
assign n_838 = ~x_145 &  n_836;
assign n_839 = ~n_837 & ~n_838;
assign n_840 =  n_800 &  n_729;
assign n_841 = ~n_516 & ~n_840;
assign n_842 =  n_351 & ~n_841;
assign n_843 =  x_144 &  n_797;
assign n_844 = ~n_842 & ~n_843;
assign n_845 =  x_144 & ~n_844;
assign n_846 = ~x_144 &  n_844;
assign n_847 = ~n_845 & ~n_846;
assign n_848 =  n_467 &  n_800;
assign n_849 = ~n_513 & ~n_848;
assign n_850 =  n_351 & ~n_849;
assign n_851 =  x_143 &  n_797;
assign n_852 = ~n_850 & ~n_851;
assign n_853 =  x_143 & ~n_852;
assign n_854 = ~x_143 &  n_852;
assign n_855 = ~n_853 & ~n_854;
assign n_856 =  n_464 &  n_800;
assign n_857 = ~n_510 & ~n_856;
assign n_858 =  n_351 & ~n_857;
assign n_859 =  x_142 &  n_797;
assign n_860 = ~n_858 & ~n_859;
assign n_861 =  x_142 & ~n_860;
assign n_862 = ~x_142 &  n_860;
assign n_863 = ~n_861 & ~n_862;
assign n_864 =  n_351 &  n_406;
assign n_865 =  x_141 &  n_375;
assign n_866 = ~n_864 & ~n_865;
assign n_867 =  x_141 & ~n_866;
assign n_868 = ~x_141 &  n_866;
assign n_869 = ~n_867 & ~n_868;
assign n_870 =  n_351 & ~n_431;
assign n_871 =  x_140 &  n_375;
assign n_872 = ~n_870 & ~n_871;
assign n_873 =  x_140 & ~n_872;
assign n_874 = ~x_140 &  n_872;
assign n_875 = ~n_873 & ~n_874;
assign n_876 =  n_351 & ~n_414;
assign n_877 =  x_139 &  n_375;
assign n_878 = ~n_876 & ~n_877;
assign n_879 =  x_139 & ~n_878;
assign n_880 = ~x_139 &  n_878;
assign n_881 = ~n_879 & ~n_880;
assign n_882 =  n_351 & ~n_395;
assign n_883 =  x_138 &  n_375;
assign n_884 = ~n_882 & ~n_883;
assign n_885 =  x_138 & ~n_884;
assign n_886 = ~x_138 &  n_884;
assign n_887 = ~n_885 & ~n_886;
assign n_888 =  n_351 & ~n_424;
assign n_889 =  x_137 &  n_375;
assign n_890 = ~n_888 & ~n_889;
assign n_891 =  x_137 & ~n_890;
assign n_892 = ~x_137 &  n_890;
assign n_893 = ~n_891 & ~n_892;
assign n_894 =  n_351 & ~n_387;
assign n_895 =  x_136 &  n_375;
assign n_896 = ~n_894 & ~n_895;
assign n_897 =  x_136 & ~n_896;
assign n_898 = ~x_136 &  n_896;
assign n_899 = ~n_897 & ~n_898;
assign n_900 =  n_351 & ~n_446;
assign n_901 =  x_135 &  n_375;
assign n_902 = ~n_900 & ~n_901;
assign n_903 =  x_135 & ~n_902;
assign n_904 = ~x_135 &  n_902;
assign n_905 = ~n_903 & ~n_904;
assign n_906 =  x_130 &  n_572;
assign n_907 = ~i_28 & ~x_84;
assign n_908 =  i_29 & ~n_907;
assign n_909 = ~n_906 & ~n_908;
assign n_910 =  x_130 & ~n_909;
assign n_911 = ~x_130 &  n_909;
assign n_912 = ~n_910 & ~n_911;
assign n_913 =  x_76 & ~n_145;
assign n_914 = ~x_75 & ~n_913;
assign n_915 =  i_29 & ~n_914;
assign n_916 =  x_129 &  n_583;
assign n_917 = ~n_915 & ~n_916;
assign n_918 =  x_129 & ~n_917;
assign n_919 = ~x_129 &  n_917;
assign n_920 = ~n_918 & ~n_919;
assign n_921 = ~i_6 & ~x_77;
assign n_922 =  x_128 &  n_921;
assign n_923 = ~n_24 & ~n_166;
assign n_924 =  x_42 & ~n_923;
assign n_925 = ~x_72 & ~n_924;
assign n_926 =  x_71 & ~n_213;
assign n_927 = ~n_925 & ~n_926;
assign n_928 =  x_77 & ~n_927;
assign n_929 = ~n_922 & ~n_928;
assign n_930 =  x_128 & ~n_929;
assign n_931 = ~x_128 &  n_929;
assign n_932 = ~n_930 & ~n_931;
assign n_933 =  x_57 &  x_77;
assign n_934 =  n_209 &  n_933;
assign n_935 =  x_127 &  n_921;
assign n_936 =  x_42 &  x_77;
assign n_937 = ~x_41 &  n_936;
assign n_938 =  n_165 &  n_937;
assign n_939 = ~n_935 & ~n_938;
assign n_940 = ~n_934 &  n_939;
assign n_941 =  x_127 & ~n_940;
assign n_942 = ~x_127 &  n_940;
assign n_943 = ~n_941 & ~n_942;
assign n_944 =  x_126 &  n_921;
assign n_945 =  x_55 &  n_7;
assign n_946 = ~x_40 &  x_42;
assign n_947 =  n_28 &  n_946;
assign n_948 = ~n_945 & ~n_947;
assign n_949 =  x_77 & ~n_948;
assign n_950 = ~n_944 & ~n_949;
assign n_951 =  x_126 & ~n_950;
assign n_952 = ~x_126 &  n_950;
assign n_953 = ~n_951 & ~n_952;
assign n_954 =  x_53 &  x_77;
assign n_955 =  n_17 &  n_954;
assign n_956 =  x_125 &  n_921;
assign n_957 = ~x_39 &  n_936;
assign n_958 =  n_39 &  n_957;
assign n_959 = ~n_956 & ~n_958;
assign n_960 = ~n_955 &  n_959;
assign n_961 =  x_125 & ~n_960;
assign n_962 = ~x_125 &  n_960;
assign n_963 = ~n_961 & ~n_962;
assign n_964 =  x_51 &  x_77;
assign n_965 =  n_207 &  n_964;
assign n_966 =  x_124 &  n_921;
assign n_967 = ~x_38 &  n_936;
assign n_968 =  n_56 &  n_967;
assign n_969 = ~n_966 & ~n_968;
assign n_970 = ~n_965 &  n_969;
assign n_971 =  x_124 & ~n_970;
assign n_972 = ~x_124 &  n_970;
assign n_973 = ~n_971 & ~n_972;
assign n_974 = ~x_37 &  n_936;
assign n_975 =  n_66 &  n_974;
assign n_976 =  x_123 &  n_921;
assign n_977 =  x_49 &  x_77;
assign n_978 =  n_202 &  n_977;
assign n_979 = ~n_976 & ~n_978;
assign n_980 = ~n_975 &  n_979;
assign n_981 =  x_123 & ~n_980;
assign n_982 = ~x_123 &  n_980;
assign n_983 = ~n_981 & ~n_982;
assign n_984 =  x_122 &  n_921;
assign n_985 =  x_47 &  n_205;
assign n_986 = ~x_36 &  x_42;
assign n_987 =  n_75 &  n_986;
assign n_988 = ~n_985 & ~n_987;
assign n_989 =  x_77 & ~n_988;
assign n_990 = ~n_984 & ~n_989;
assign n_991 =  x_122 & ~n_990;
assign n_992 = ~x_122 &  n_990;
assign n_993 = ~n_991 & ~n_992;
assign n_994 =  x_121 &  n_921;
assign n_995 =  x_44 &  n_200;
assign n_996 = ~x_34 &  x_42;
assign n_997 =  n_163 &  n_996;
assign n_998 = ~n_995 & ~n_997;
assign n_999 =  x_77 & ~n_998;
assign n_1000 = ~n_994 & ~n_999;
assign n_1001 =  x_121 & ~n_1000;
assign n_1002 = ~x_121 &  n_1000;
assign n_1003 = ~n_1001 & ~n_1002;
assign n_1004 =  x_77 & ~n_152;
assign n_1005 = ~i_5 & ~x_77;
assign n_1006 =  x_120 &  n_1005;
assign n_1007 = ~n_1004 & ~n_1006;
assign n_1008 =  x_120 & ~n_1007;
assign n_1009 = ~x_120 &  n_1007;
assign n_1010 = ~n_1008 & ~n_1009;
assign n_1011 =  x_77 & ~n_137;
assign n_1012 =  x_119 &  n_1005;
assign n_1013 = ~n_1011 & ~n_1012;
assign n_1014 =  x_119 & ~n_1013;
assign n_1015 = ~x_119 &  n_1013;
assign n_1016 = ~n_1014 & ~n_1015;
assign n_1017 =  x_77 & ~n_117;
assign n_1018 =  x_118 &  n_1005;
assign n_1019 = ~n_1017 & ~n_1018;
assign n_1020 =  x_118 & ~n_1019;
assign n_1021 = ~x_118 &  n_1019;
assign n_1022 = ~n_1020 & ~n_1021;
assign n_1023 =  x_77 & ~n_133;
assign n_1024 =  x_117 &  n_1005;
assign n_1025 = ~n_1023 & ~n_1024;
assign n_1026 =  x_117 & ~n_1025;
assign n_1027 = ~x_117 &  n_1025;
assign n_1028 = ~n_1026 & ~n_1027;
assign n_1029 =  x_77 & ~n_110;
assign n_1030 =  x_116 &  n_1005;
assign n_1031 = ~n_1029 & ~n_1030;
assign n_1032 =  x_116 & ~n_1031;
assign n_1033 = ~x_116 &  n_1031;
assign n_1034 = ~n_1032 & ~n_1033;
assign n_1035 =  x_77 & ~n_126;
assign n_1036 =  x_115 &  n_1005;
assign n_1037 = ~n_1035 & ~n_1036;
assign n_1038 =  x_115 & ~n_1037;
assign n_1039 = ~x_115 &  n_1037;
assign n_1040 = ~n_1038 & ~n_1039;
assign n_1041 =  x_114 &  n_1005;
assign n_1042 =  x_77 & ~n_103;
assign n_1043 = ~n_1041 & ~n_1042;
assign n_1044 =  x_114 & ~n_1043;
assign n_1045 = ~x_114 &  n_1043;
assign n_1046 = ~n_1044 & ~n_1045;
assign n_1047 =  x_113 &  n_1005;
assign n_1048 =  x_77 & ~n_184;
assign n_1049 = ~n_1047 & ~n_1048;
assign n_1050 =  x_113 & ~n_1049;
assign n_1051 = ~x_113 &  n_1049;
assign n_1052 = ~n_1050 & ~n_1051;
assign n_1053 =  x_112 & ~n_292;
assign n_1054 = ~x_112 &  n_292;
assign n_1055 = ~n_1053 & ~n_1054;
assign n_1056 =  x_111 & ~n_288;
assign n_1057 = ~x_111 &  n_288;
assign n_1058 = ~n_1056 & ~n_1057;
assign n_1059 =  x_110 &  n_564;
assign n_1060 = ~n_1059 & ~n_563;
assign n_1061 =  x_110 & ~n_1060;
assign n_1062 = ~x_110 &  n_1060;
assign n_1063 = ~n_1061 & ~n_1062;
assign n_1064 =  x_109 &  n_552;
assign n_1065 = ~n_1064 & ~n_551;
assign n_1066 =  x_109 & ~n_1065;
assign n_1067 = ~x_109 &  n_1065;
assign n_1068 = ~n_1066 & ~n_1067;
assign n_1069 =  n_192 & ~n_230;
assign n_1070 =  n_1069 & ~n_233;
assign n_1071 = ~n_1060 &  n_1070;
assign n_1072 =  x_108 &  n_1071;
assign n_1073 = ~x_108 & ~n_1071;
assign n_1074 = ~n_1072 & ~n_1073;
assign n_1075 =  n_1065 &  n_234;
assign n_1076 = ~n_192 & ~n_1075;
assign n_1077 =  x_107 &  n_1076;
assign n_1078 = ~x_107 & ~n_1076;
assign n_1079 = ~n_1077 & ~n_1078;
assign n_1080 =  x_106 &  n_749;
assign n_1081 = ~n_1080 & ~n_748;
assign n_1082 =  x_106 & ~n_1081;
assign n_1083 = ~x_106 &  n_1081;
assign n_1084 = ~n_1082 & ~n_1083;
assign n_1085 =  x_105 &  n_749;
assign n_1086 = ~n_1085 & ~n_755;
assign n_1087 =  x_105 & ~n_1086;
assign n_1088 = ~x_105 &  n_1086;
assign n_1089 = ~n_1087 & ~n_1088;
assign n_1090 =  x_104 &  n_749;
assign n_1091 = ~n_1090 & ~n_761;
assign n_1092 =  x_104 & ~n_1091;
assign n_1093 = ~x_104 &  n_1091;
assign n_1094 = ~n_1092 & ~n_1093;
assign n_1095 =  x_103 &  n_749;
assign n_1096 = ~n_1095 & ~n_767;
assign n_1097 =  x_103 & ~n_1096;
assign n_1098 = ~x_103 &  n_1096;
assign n_1099 = ~n_1097 & ~n_1098;
assign n_1100 =  x_102 &  n_749;
assign n_1101 = ~n_1100 & ~n_773;
assign n_1102 =  x_102 & ~n_1101;
assign n_1103 = ~x_102 &  n_1101;
assign n_1104 = ~n_1102 & ~n_1103;
assign n_1105 =  x_101 &  n_749;
assign n_1106 = ~n_1105 & ~n_779;
assign n_1107 =  x_101 & ~n_1106;
assign n_1108 = ~x_101 &  n_1106;
assign n_1109 = ~n_1107 & ~n_1108;
assign n_1110 =  x_100 &  n_749;
assign n_1111 = ~n_1110 & ~n_785;
assign n_1112 =  x_100 & ~n_1111;
assign n_1113 = ~x_100 &  n_1111;
assign n_1114 = ~n_1112 & ~n_1113;
assign n_1115 =  x_99 &  n_749;
assign n_1116 = ~n_1115 & ~n_791;
assign n_1117 =  x_99 & ~n_1116;
assign n_1118 = ~x_99 &  n_1116;
assign n_1119 = ~n_1117 & ~n_1118;
assign n_1120 = ~n_29 & ~n_31;
assign n_1121 =  n_165 & ~n_1120;
assign n_1122 =  x_98 &  n_1121;
assign n_1123 = ~x_98 & ~n_1121;
assign n_1124 = ~n_1122 & ~n_1123;
assign n_1125 =  x_97 &  n_1;
assign n_1126 =  i_29 &  x_50;
assign n_1127 =  n_207 &  n_1126;
assign n_1128 = ~n_1125 & ~n_1127;
assign n_1129 =  x_97 & ~n_1128;
assign n_1130 = ~x_97 &  n_1128;
assign n_1131 = ~n_1129 & ~n_1130;
assign n_1132 =  x_96 &  n_1;
assign n_1133 =  i_29 &  x_46;
assign n_1134 =  n_205 &  n_1133;
assign n_1135 = ~n_1132 & ~n_1134;
assign n_1136 =  x_96 & ~n_1135;
assign n_1137 = ~x_96 &  n_1135;
assign n_1138 = ~n_1136 & ~n_1137;
assign n_1139 =  i_29 &  n_203;
assign n_1140 =  x_95 &  n_1;
assign n_1141 = ~n_1139 & ~n_1140;
assign n_1142 =  x_95 & ~n_1141;
assign n_1143 = ~x_95 &  n_1141;
assign n_1144 = ~n_1142 & ~n_1143;
assign n_1145 =  x_94 &  n_1;
assign n_1146 =  x_94 & ~n_211;
assign n_1147 =  x_56 & ~n_208;
assign n_1148 = ~n_1146 &  n_1147;
assign n_1149 = ~n_1145 & ~n_1148;
assign n_1150 =  x_94 & ~n_1149;
assign n_1151 = ~x_94 &  n_1149;
assign n_1152 = ~n_1150 & ~n_1151;
assign n_1153 =  n_323 & ~n_272;
assign n_1154 =  x_62 &  n_1153;
assign n_1155 = ~x_62 & ~n_1153;
assign n_1156 = ~n_1154 & ~n_1155;
assign n_1157 =  i_29 & ~n_184;
assign n_1158 =  x_33 &  n_240;
assign n_1159 = ~n_1157 & ~n_1158;
assign n_1160 = ~n_1159 &  n_323;
assign n_1161 =  x_61 &  n_1160;
assign n_1162 = ~x_61 & ~n_1160;
assign n_1163 = ~n_1161 & ~n_1162;
assign n_1164 =  x_60 & ~n_300;
assign n_1165 = ~x_60 &  n_300;
assign n_1166 = ~n_1164 & ~n_1165;
assign n_1167 =  x_59 & ~n_326;
assign n_1168 = ~x_59 &  n_326;
assign n_1169 = ~n_1167 & ~n_1168;
assign n_1170 =  x_58 &  n_323;
assign n_1171 = ~x_58 & ~n_323;
assign n_1172 = ~n_1170 & ~n_1171;
assign n_1173 =  x_57 &  n_309;
assign n_1174 = ~x_57 & ~n_309;
assign n_1175 = ~n_1173 & ~n_1174;
assign n_1176 =  x_56 &  n_309;
assign n_1177 = ~x_56 & ~n_309;
assign n_1178 = ~n_1176 & ~n_1177;
assign n_1179 =  x_55 &  n_309;
assign n_1180 = ~x_55 & ~n_309;
assign n_1181 = ~n_1179 & ~n_1180;
assign n_1182 =  x_54 &  n_309;
assign n_1183 = ~x_54 & ~n_309;
assign n_1184 = ~n_1182 & ~n_1183;
assign n_1185 =  x_53 &  n_309;
assign n_1186 = ~x_53 & ~n_309;
assign n_1187 = ~n_1185 & ~n_1186;
assign n_1188 =  x_52 &  n_309;
assign n_1189 = ~x_52 & ~n_309;
assign n_1190 = ~n_1188 & ~n_1189;
assign n_1191 =  x_51 &  n_309;
assign n_1192 = ~x_51 & ~n_309;
assign n_1193 = ~n_1191 & ~n_1192;
assign n_1194 =  x_50 &  n_309;
assign n_1195 = ~x_50 & ~n_309;
assign n_1196 = ~n_1194 & ~n_1195;
assign n_1197 =  x_49 &  n_309;
assign n_1198 = ~x_49 & ~n_309;
assign n_1199 = ~n_1197 & ~n_1198;
assign n_1200 =  x_48 &  n_309;
assign n_1201 = ~x_48 & ~n_309;
assign n_1202 = ~n_1200 & ~n_1201;
assign n_1203 =  x_47 &  n_309;
assign n_1204 = ~x_47 & ~n_309;
assign n_1205 = ~n_1203 & ~n_1204;
assign n_1206 =  x_46 &  n_309;
assign n_1207 = ~x_46 & ~n_309;
assign n_1208 = ~n_1206 & ~n_1207;
assign n_1209 =  x_45 &  n_1;
assign n_1210 =  i_29 &  x_43;
assign n_1211 =  n_200 &  n_1210;
assign n_1212 = ~n_1209 & ~n_1211;
assign n_1213 =  x_45 & ~n_1212;
assign n_1214 = ~x_45 &  n_1212;
assign n_1215 = ~n_1213 & ~n_1214;
assign n_1216 =  x_44 &  n_309;
assign n_1217 = ~x_44 & ~n_309;
assign n_1218 = ~n_1216 & ~n_1217;
assign n_1219 =  x_43 &  n_309;
assign n_1220 = ~x_43 & ~n_309;
assign n_1221 = ~n_1219 & ~n_1220;
assign n_1222 =  x_42 &  n_284;
assign n_1223 = ~x_42 & ~n_284;
assign n_1224 = ~n_1222 & ~n_1223;
assign n_1225 =  x_41 &  n_309;
assign n_1226 = ~x_41 & ~n_309;
assign n_1227 = ~n_1225 & ~n_1226;
assign n_1228 =  x_40 &  n_309;
assign n_1229 = ~x_40 & ~n_309;
assign n_1230 = ~n_1228 & ~n_1229;
assign n_1231 =  x_39 &  n_309;
assign n_1232 = ~x_39 & ~n_309;
assign n_1233 = ~n_1231 & ~n_1232;
assign n_1234 =  x_38 &  n_309;
assign n_1235 = ~x_38 & ~n_309;
assign n_1236 = ~n_1234 & ~n_1235;
assign n_1237 =  x_37 &  n_309;
assign n_1238 = ~x_37 & ~n_309;
assign n_1239 = ~n_1237 & ~n_1238;
assign n_1240 =  x_36 &  n_309;
assign n_1241 = ~x_36 & ~n_309;
assign n_1242 = ~n_1240 & ~n_1241;
assign n_1243 =  n_163 &  n_29;
assign n_1244 =  x_35 &  n_31;
assign n_1245 = ~n_1243 & ~n_1244;
assign n_1246 =  x_35 & ~n_1245;
assign n_1247 = ~x_35 &  n_1245;
assign n_1248 = ~n_1246 & ~n_1247;
assign n_1249 =  x_34 &  n_309;
assign n_1250 = ~x_34 & ~n_309;
assign n_1251 = ~n_1249 & ~n_1250;
assign n_1252 =  x_33 & ~n_1159;
assign n_1253 = ~x_33 &  n_1159;
assign n_1254 = ~n_1252 & ~n_1253;
assign n_1255 =  x_32 &  n_230;
assign n_1256 = ~x_32 & ~n_230;
assign n_1257 = ~n_1255 & ~n_1256;
assign n_1258 = ~n_1065 &  n_233;
assign n_1259 =  n_1069 &  n_1258;
assign n_1260 =  x_30 &  n_1259;
assign n_1261 = ~x_30 & ~n_1259;
assign n_1262 = ~n_1260 & ~n_1261;
assign n_1263 =  n_1060 &  n_1070;
assign n_1264 =  x_31 &  n_1263;
assign n_1265 = ~x_31 & ~n_1263;
assign n_1266 = ~n_1264 & ~n_1265;
assign n_1267 = ~n_1262 & ~n_1266;
assign n_1268 = ~n_1257 &  n_1267;
assign n_1269 = ~n_1254 &  n_1268;
assign n_1270 = ~n_1251 &  n_1269;
assign n_1271 = ~n_1248 &  n_1270;
assign n_1272 = ~n_1242 &  n_1271;
assign n_1273 = ~n_1239 &  n_1272;
assign n_1274 = ~n_1236 &  n_1273;
assign n_1275 = ~n_1233 &  n_1274;
assign n_1276 = ~n_1230 &  n_1275;
assign n_1277 = ~n_1227 &  n_1276;
assign n_1278 = ~n_1224 &  n_1277;
assign n_1279 = ~n_1221 &  n_1278;
assign n_1280 = ~n_1218 &  n_1279;
assign n_1281 = ~n_1215 &  n_1280;
assign n_1282 = ~n_1208 &  n_1281;
assign n_1283 = ~n_1205 &  n_1282;
assign n_1284 = ~n_1202 &  n_1283;
assign n_1285 = ~n_1199 &  n_1284;
assign n_1286 = ~n_1196 &  n_1285;
assign n_1287 = ~n_1193 &  n_1286;
assign n_1288 = ~n_1190 &  n_1287;
assign n_1289 = ~n_1187 &  n_1288;
assign n_1290 = ~n_1184 &  n_1289;
assign n_1291 = ~n_1181 &  n_1290;
assign n_1292 = ~n_1178 &  n_1291;
assign n_1293 = ~n_1175 &  n_1292;
assign n_1294 = ~n_1172 &  n_1293;
assign n_1295 = ~n_1169 &  n_1294;
assign n_1296 = ~n_1166 &  n_1295;
assign n_1297 = ~n_1163 &  n_1296;
assign n_1298 = ~n_1156 &  n_1297;
assign n_1299 = ~n_1152 &  n_1298;
assign n_1300 = ~n_1144 &  n_1299;
assign n_1301 = ~n_1138 &  n_1300;
assign n_1302 = ~n_1131 &  n_1301;
assign n_1303 = ~n_1124 &  n_1302;
assign n_1304 = ~n_1119 &  n_1303;
assign n_1305 = ~n_1114 &  n_1304;
assign n_1306 = ~n_1109 &  n_1305;
assign n_1307 = ~n_1104 &  n_1306;
assign n_1308 = ~n_1099 &  n_1307;
assign n_1309 = ~n_1094 &  n_1308;
assign n_1310 = ~n_1089 &  n_1309;
assign n_1311 = ~n_1084 &  n_1310;
assign n_1312 = ~n_1079 &  n_1311;
assign n_1313 = ~n_1074 &  n_1312;
assign n_1314 = ~n_1068 &  n_1313;
assign n_1315 = ~n_1063 &  n_1314;
assign n_1316 = ~n_1058 &  n_1315;
assign n_1317 = ~n_1055 &  n_1316;
assign n_1318 = ~n_1052 &  n_1317;
assign n_1319 = ~n_1046 &  n_1318;
assign n_1320 = ~n_1040 &  n_1319;
assign n_1321 = ~n_1034 &  n_1320;
assign n_1322 = ~n_1028 &  n_1321;
assign n_1323 = ~n_1022 &  n_1322;
assign n_1324 = ~n_1016 &  n_1323;
assign n_1325 = ~n_1010 &  n_1324;
assign n_1326 = ~n_1003 &  n_1325;
assign n_1327 = ~n_993 &  n_1326;
assign n_1328 = ~n_983 &  n_1327;
assign n_1329 = ~n_973 &  n_1328;
assign n_1330 = ~n_963 &  n_1329;
assign n_1331 = ~n_953 &  n_1330;
assign n_1332 = ~n_943 &  n_1331;
assign n_1333 = ~n_932 &  n_1332;
assign n_1334 = ~n_920 &  n_1333;
assign n_1335 = ~n_912 &  n_1334;
assign n_1336 = ~n_905 &  n_1335;
assign n_1337 = ~n_899 &  n_1336;
assign n_1338 = ~n_893 &  n_1337;
assign n_1339 = ~n_887 &  n_1338;
assign n_1340 = ~n_881 &  n_1339;
assign n_1341 = ~n_875 &  n_1340;
assign n_1342 = ~n_869 &  n_1341;
assign n_1343 = ~n_863 &  n_1342;
assign n_1344 = ~n_855 &  n_1343;
assign n_1345 = ~n_847 &  n_1344;
assign n_1346 = ~n_839 &  n_1345;
assign n_1347 = ~n_831 &  n_1346;
assign n_1348 = ~n_823 &  n_1347;
assign n_1349 = ~n_815 &  n_1348;
assign n_1350 = ~n_807 &  n_1349;
assign n_1351 = ~n_796 &  n_1350;
assign n_1352 = ~n_790 &  n_1351;
assign n_1353 = ~n_784 &  n_1352;
assign n_1354 = ~n_778 &  n_1353;
assign n_1355 = ~n_772 &  n_1354;
assign n_1356 = ~n_766 &  n_1355;
assign n_1357 = ~n_760 &  n_1356;
assign n_1358 = ~n_754 &  n_1357;
assign n_1359 = ~n_747 &  n_1358;
assign n_1360 = ~n_741 &  n_1359;
assign n_1361 = ~n_735 &  n_1360;
assign n_1362 = ~n_727 &  n_1361;
assign n_1363 = ~n_721 &  n_1362;
assign n_1364 = ~n_715 &  n_1363;
assign n_1365 = ~n_706 &  n_1364;
assign n_1366 = ~n_700 &  n_1365;
assign n_1367 = ~n_694 &  n_1366;
assign n_1368 = ~n_688 &  n_1367;
assign n_1369 = ~n_682 &  n_1368;
assign n_1370 = ~n_676 &  n_1369;
assign n_1371 = ~n_670 &  n_1370;
assign n_1372 = ~n_664 &  n_1371;
assign n_1373 = ~n_655 &  n_1372;
assign n_1374 = ~n_648 &  n_1373;
assign n_1375 = ~n_642 &  n_1374;
assign n_1376 = ~n_636 &  n_1375;
assign n_1377 = ~n_630 &  n_1376;
assign n_1378 = ~n_624 &  n_1377;
assign n_1379 = ~n_618 &  n_1378;
assign n_1380 = ~n_612 &  n_1379;
assign n_1381 = ~n_606 &  n_1380;
assign n_1382 = ~n_600 &  n_1381;
assign n_1383 = ~n_594 &  n_1382;
assign n_1384 = ~n_588 &  n_1383;
assign n_1385 = ~n_577 &  n_1384;
assign n_1386 = ~n_569 &  n_1385;
assign n_1387 = ~n_562 &  n_1386;
assign n_1388 = ~n_557 &  n_1387;
assign n_1389 = ~n_550 &  n_1388;
assign n_1390 = ~n_540 &  n_1389;
assign n_1391 = ~n_494 &  n_1390;
assign n_1392 = ~n_380 &  n_1391;
assign n_1393 = ~n_350 &  n_1392;
assign n_1394 = ~n_346 &  n_1393;
assign n_1395 = ~n_342 &  n_1394;
assign n_1396 = ~n_338 &  n_1395;
assign n_1397 = ~n_334 &  n_1396;
assign n_1398 = ~n_330 &  n_1397;
assign n_1399 = ~n_322 &  n_1398;
assign n_1400 = ~n_319 &  n_1399;
assign n_1401 = ~n_315 &  n_1400;
assign n_1402 = ~n_312 &  n_1401;
assign n_1403 = ~n_308 &  n_1402;
assign n_1404 = ~n_304 &  n_1403;
assign n_1405 = ~n_299 &  n_1404;
assign n_1406 = ~n_283 &  n_1405;
assign n_1407 = ~n_279 &  n_1406;
assign n_1408 = ~n_275 &  n_1407;
assign n_1409 = ~n_269 &  n_1408;
assign n_1410 = ~n_263 &  n_1409;
assign n_1411 = ~n_257 &  n_1410;
assign n_1412 = ~n_251 &  n_1411;
assign n_1413 = ~n_245 &  n_1412;
assign n_1414 = ~n_238 &  n_1413;
assign n_1415 = ~n_89 &  n_1414;
assign n_1416 = ~n_81 &  n_1415;
assign n_1417 = ~n_72 &  n_1416;
assign n_1418 = ~n_62 &  n_1417;
assign n_1419 = ~n_53 &  n_1418;
assign n_1420 = ~n_45 &  n_1419;
assign n_1421 = ~n_36 &  n_1420;
assign n_1422 = ~n_23 &  n_1421;
assign n_1423 = ~n_13 &  n_1422;
assign o_1 = ~n_1423;
endmodule

