// Benchmark "SKOLEMFORMULA" written by ABC on Wed May 18 01:44:36 2022

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4,
    i5, i6, i7, i8, i9  );
  input  i0, i1, i2, i3, i4;
  output i5, i6, i7, i8, i9;
  assign i5 = i0;
  assign i6 = i1;
  assign i7 = i2;
  assign i8 = i3;
  assign i9 = i4;
endmodule


