module formula(v_188,v_190,v_192,v_194,v_196,v_198,v_200,v_202,v_204,v_206,v_208,v_210,v_212,v_214,v_216,v_218,v_220,v_222,v_224,v_226,v_228,v_230,v_232,v_234,v_236,v_238,v_240,v_242,v_244,v_246,v_248,v_250,v_251,v_252,v_253,v_254,v_255,v_256,v_257,v_258,v_259,v_260,v_261,v_262,v_263,v_264,v_265,v_266,v_267,v_268,v_269,v_270,v_271,v_272,v_273,v_274,v_275,v_276,v_277,v_278,v_279,v_280,v_281,v_282,v_191,v_203,v_223,v_231,v_235,v_243,v_7,v_8,v_9,v_12,v_13,v_14,v_15,v_16,v_17,v_18,v_19,v_20,v_21,v_24,v_25,v_26,v_27,v_28,v_29,v_30,v_31,v_32,v_33,v_34,v_35,v_36,v_37,v_38,v_39,v_40,v_41,v_44,v_45,v_46,v_47,v_48,v_49,v_52,v_53,v_56,v_57,v_58,v_59,v_60,v_61,v_73,v_74,o_1);
	input v_188;
	input v_190;
	input v_192;
	input v_194;
	input v_196;
	input v_198;
	input v_200;
	input v_202;
	input v_204;
	input v_206;
	input v_208;
	input v_210;
	input v_212;
	input v_214;
	input v_216;
	input v_218;
	input v_220;
	input v_222;
	input v_224;
	input v_226;
	input v_228;
	input v_230;
	input v_232;
	input v_234;
	input v_236;
	input v_238;
	input v_240;
	input v_242;
	input v_244;
	input v_246;
	input v_248;
	input v_250;
	input v_251;
	input v_252;
	input v_253;
	input v_254;
	input v_255;
	input v_256;
	input v_257;
	input v_258;
	input v_259;
	input v_260;
	input v_261;
	input v_262;
	input v_263;
	input v_264;
	input v_265;
	input v_266;
	input v_267;
	input v_268;
	input v_269;
	input v_270;
	input v_271;
	input v_272;
	input v_273;
	input v_274;
	input v_275;
	input v_276;
	input v_277;
	input v_278;
	input v_279;
	input v_280;
	input v_281;
	input v_282;
	input v_191;
	input v_203;
	input v_223;
	input v_231;
	input v_235;
	input v_243;
	input v_7;
	input v_8;
	input v_9;
	input v_12;
	input v_13;
	input v_14;
	input v_15;
	input v_16;
	input v_17;
	input v_18;
	input v_19;
	input v_20;
	input v_21;
	input v_24;
	input v_25;
	input v_26;
	input v_27;
	input v_28;
	input v_29;
	input v_30;
	input v_31;
	input v_32;
	input v_33;
	input v_34;
	input v_35;
	input v_36;
	input v_37;
	input v_38;
	input v_39;
	input v_40;
	input v_41;
	input v_44;
	input v_45;
	input v_46;
	input v_47;
	input v_48;
	input v_49;
	input v_52;
	input v_53;
	input v_56;
	input v_57;
	input v_58;
	input v_59;
	input v_60;
	input v_61;
	input v_73;
	input v_74;
	wire v_187;
	wire v_189;
	wire v_193;
	wire v_195;
	wire v_197;
	wire v_199;
	wire v_201;
	wire v_205;
	wire v_207;
	wire v_209;
	wire v_211;
	wire v_213;
	wire v_215;
	wire v_217;
	wire v_219;
	wire v_221;
	wire v_225;
	wire v_227;
	wire v_229;
	wire v_233;
	wire v_237;
	wire v_239;
	wire v_241;
	wire v_245;
	wire v_247;
	wire v_249;
	wire v_1;
	wire v_2;
	wire v_3;
	wire v_4;
	wire v_5;
	wire v_6;
	wire v_10;
	wire v_11;
	wire v_22;
	wire v_23;
	wire v_42;
	wire v_43;
	wire v_50;
	wire v_51;
	wire v_54;
	wire v_55;
	wire v_62;
	wire v_63;
	wire v_64;
	wire v_65;
	wire v_66;
	wire v_67;
	wire v_68;
	wire v_69;
	wire v_70;
	wire v_71;
	wire v_72;
	wire v_75;
	wire v_76;
	wire v_77;
	wire v_78;
	wire v_79;
	wire v_80;
	wire v_81;
	wire v_82;
	wire v_83;
	wire v_84;
	wire v_85;
	wire v_86;
	wire v_87;
	wire v_88;
	wire v_89;
	wire v_90;
	wire v_91;
	wire v_92;
	wire v_93;
	wire v_94;
	wire v_95;
	wire v_96;
	wire v_97;
	wire v_98;
	wire v_99;
	wire v_100;
	wire v_101;
	wire v_102;
	wire v_103;
	wire v_104;
	wire v_105;
	wire v_106;
	wire v_107;
	wire v_108;
	wire v_109;
	wire v_110;
	wire v_111;
	wire v_112;
	wire v_113;
	wire v_114;
	wire v_115;
	wire v_116;
	wire v_117;
	wire v_118;
	wire v_119;
	wire v_120;
	wire v_121;
	wire v_122;
	wire v_123;
	wire v_124;
	wire v_125;
	wire v_126;
	wire v_127;
	wire v_128;
	wire v_129;
	wire v_130;
	wire v_131;
	wire v_132;
	wire v_133;
	wire v_134;
	wire v_135;
	wire v_136;
	wire v_137;
	wire v_138;
	wire v_139;
	wire v_140;
	wire v_141;
	wire v_142;
	wire v_143;
	wire v_144;
	wire v_145;
	wire v_146;
	wire v_147;
	wire v_148;
	wire v_149;
	wire v_150;
	wire v_151;
	wire v_152;
	wire v_153;
	wire v_154;
	wire v_155;
	wire v_156;
	wire v_157;
	wire v_158;
	wire v_159;
	wire v_160;
	wire v_161;
	wire v_162;
	wire v_163;
	wire v_164;
	wire v_165;
	wire v_166;
	wire v_167;
	wire v_168;
	wire v_169;
	wire v_170;
	wire v_171;
	wire v_172;
	wire v_173;
	wire v_174;
	wire v_175;
	wire v_176;
	wire v_177;
	wire v_178;
	wire v_179;
	wire v_180;
	wire v_181;
	wire v_182;
	wire v_183;
	wire v_184;
	wire v_185;
	wire v_186;
	wire v_283;
	wire x_1;
	wire x_2;
	wire x_3;
	wire x_4;
	wire x_5;
	wire x_6;
	wire x_7;
	wire x_8;
	wire x_9;
	wire x_10;
	wire x_11;
	wire x_12;
	wire x_13;
	wire x_14;
	wire x_15;
	wire x_16;
	wire x_17;
	wire x_18;
	wire x_19;
	wire x_20;
	wire x_21;
	wire x_22;
	wire x_23;
	wire x_24;
	wire x_25;
	wire x_26;
	wire x_27;
	wire x_28;
	wire x_29;
	wire x_30;
	wire x_31;
	wire x_32;
	wire x_33;
	wire x_34;
	wire x_35;
	wire x_36;
	wire x_37;
	wire x_38;
	wire x_39;
	wire x_40;
	wire x_41;
	wire x_42;
	wire x_43;
	wire x_44;
	wire x_45;
	wire x_46;
	wire x_47;
	wire x_48;
	wire x_49;
	wire x_50;
	wire x_51;
	wire x_52;
	wire x_53;
	wire x_54;
	wire x_55;
	wire x_56;
	wire x_57;
	wire x_58;
	wire x_59;
	wire x_60;
	wire x_61;
	wire x_62;
	wire x_63;
	wire x_64;
	wire x_65;
	wire x_66;
	wire x_67;
	wire x_68;
	wire x_69;
	wire x_70;
	wire x_71;
	wire x_72;
	wire x_73;
	wire x_74;
	wire x_75;
	wire x_76;
	wire x_77;
	wire x_78;
	wire x_79;
	wire x_80;
	wire x_81;
	wire x_82;
	wire x_83;
	wire x_84;
	wire x_85;
	wire x_86;
	wire x_87;
	wire x_88;
	wire x_89;
	wire x_90;
	wire x_91;
	wire x_92;
	wire x_93;
	wire x_94;
	wire x_95;
	wire x_96;
	wire x_97;
	wire x_98;
	wire x_99;
	wire x_100;
	wire x_101;
	wire x_102;
	wire x_103;
	wire x_104;
	wire x_105;
	wire x_106;
	wire x_107;
	wire x_108;
	wire x_109;
	wire x_110;
	wire x_111;
	wire x_112;
	wire x_113;
	wire x_114;
	wire x_115;
	wire x_116;
	wire x_117;
	wire x_118;
	wire x_119;
	wire x_120;
	wire x_121;
	wire x_122;
	wire x_123;
	wire x_124;
	wire x_125;
	wire x_126;
	wire x_127;
	wire x_128;
	wire x_129;
	wire x_130;
	wire x_131;
	wire x_132;
	wire x_133;
	wire x_134;
	wire x_135;
	wire x_136;
	wire x_137;
	wire x_138;
	wire x_139;
	wire x_140;
	wire x_141;
	wire x_142;
	wire x_143;
	wire x_144;
	wire x_145;
	wire x_146;
	wire x_147;
	wire x_148;
	wire x_149;
	wire x_150;
	wire x_151;
	wire x_152;
	wire x_153;
	wire x_154;
	wire x_155;
	wire x_156;
	wire x_157;
	wire x_158;
	wire x_159;
	wire x_160;
	wire x_161;
	wire x_162;
	wire x_163;
	wire x_164;
	wire x_165;
	wire x_166;
	wire x_167;
	wire x_168;
	wire x_169;
	wire x_170;
	wire x_171;
	wire x_172;
	wire x_173;
	wire x_174;
	wire x_175;
	wire x_176;
	wire x_177;
	wire x_178;
	wire x_179;
	wire x_180;
	wire x_181;
	wire x_182;
	wire x_183;
	wire x_184;
	wire x_185;
	wire x_186;
	wire x_187;
	wire x_188;
	wire x_189;
	wire x_190;
	wire x_191;
	wire x_192;
	wire x_193;
	wire x_194;
	wire x_195;
	wire x_196;
	wire x_197;
	wire x_198;
	wire x_199;
	wire x_200;
	wire x_201;
	wire x_202;
	wire x_203;
	wire x_204;
	wire x_205;
	wire x_206;
	wire x_207;
	wire x_208;
	wire x_209;
	wire x_210;
	wire x_211;
	wire x_212;
	wire x_213;
	wire x_214;
	wire x_215;
	wire x_216;
	wire x_217;
	wire x_218;
	wire x_219;
	wire x_220;
	wire x_221;
	wire x_222;
	wire x_223;
	wire x_224;
	wire x_225;
	wire x_226;
	wire x_227;
	wire x_228;
	wire x_229;
	wire x_230;
	wire x_231;
	wire x_232;
	wire x_233;
	wire x_234;
	wire x_235;
	wire x_236;
	wire x_237;
	wire x_238;
	wire x_239;
	wire x_240;
	wire x_241;
	wire x_242;
	wire x_243;
	wire x_244;
	wire x_245;
	wire x_246;
	wire x_247;
	wire x_248;
	wire x_249;
	wire x_250;
	wire x_251;
	wire x_252;
	wire x_253;
	wire x_254;
	wire x_255;
	wire x_256;
	wire x_257;
	wire x_258;
	wire x_259;
	wire x_260;
	wire x_261;
	wire x_262;
	wire x_263;
	wire x_264;
	wire x_265;
	wire x_266;
	wire x_267;
	wire x_268;
	wire x_269;
	wire x_270;
	wire x_271;
	wire x_272;
	wire x_273;
	wire x_274;
	wire x_275;
	wire x_276;
	wire x_277;
	wire x_278;
	wire x_279;
	wire x_280;
	wire x_281;
	wire x_282;
	wire x_283;
	wire x_284;
	wire x_285;
	wire x_286;
	wire x_287;
	wire x_288;
	wire x_289;
	wire x_290;
	wire x_291;
	wire x_292;
	wire x_293;
	wire x_294;
	wire x_295;
	wire x_296;
	wire x_297;
	wire x_298;
	wire x_299;
	wire x_300;
	wire x_301;
	wire x_302;
	wire x_303;
	wire x_304;
	wire x_305;
	wire x_306;
	wire x_307;
	wire x_308;
	wire x_309;
	wire x_310;
	wire x_311;
	wire x_312;
	wire x_313;
	wire x_314;
	wire x_315;
	wire x_316;
	wire x_317;
	wire x_318;
	wire x_319;
	wire x_320;
	wire x_321;
	wire x_322;
	wire x_323;
	wire x_324;
	wire x_325;
	wire x_326;
	wire x_327;
	wire x_328;
	wire x_329;
	wire x_330;
	wire x_331;
	wire x_332;
	wire x_333;
	wire x_334;
	wire x_335;
	wire x_336;
	wire x_337;
	wire x_338;
	wire x_339;
	wire x_340;
	wire x_341;
	wire x_342;
	wire x_343;
	wire x_344;
	wire x_345;
	wire x_346;
	wire x_347;
	wire x_348;
	wire x_349;
	wire x_350;
	wire x_351;
	wire x_352;
	wire x_353;
	wire x_354;
	wire x_355;
	wire x_356;
	wire x_357;
	wire x_358;
	wire x_359;
	wire x_360;
	wire x_361;
	wire x_362;
	wire x_363;
	wire x_364;
	wire x_365;
	wire x_366;
	wire x_367;
	wire x_368;
	wire x_369;
	wire x_370;
	wire x_371;
	wire x_372;
	wire x_373;
	wire x_374;
	wire x_375;
	wire x_376;
	wire x_377;
	wire x_378;
	wire x_379;
	wire x_380;
	wire x_381;
	wire x_382;
	wire x_383;
	wire x_384;
	wire x_385;
	wire x_386;
	wire x_387;
	wire x_388;
	wire x_389;
	wire x_390;
	wire x_391;
	wire x_392;
	wire x_393;
	wire x_394;
	wire x_395;
	wire x_396;
	wire x_397;
	wire x_398;
	wire x_399;
	wire x_400;
	wire x_401;
	wire x_402;
	wire x_403;
	wire x_404;
	wire x_405;
	wire x_406;
	wire x_407;
	wire x_408;
	wire x_409;
	wire x_410;
	wire x_411;
	wire x_412;
	wire x_413;
	wire x_414;
	wire x_415;
	wire x_416;
	wire x_417;
	wire x_418;
	wire x_419;
	wire x_420;
	wire x_421;
	wire x_422;
	wire x_423;
	wire x_424;
	wire x_425;
	wire x_426;
	wire x_427;
	wire x_428;
	wire x_429;
	wire x_430;
	wire x_431;
	wire x_432;
	wire x_433;
	wire x_434;
	wire x_435;
	wire x_436;
	wire x_437;
	wire x_438;
	wire x_439;
	wire x_440;
	wire x_441;
	wire x_442;
	wire x_443;
	wire x_444;
	wire x_445;
	wire x_446;
	wire x_447;
	wire x_448;
	wire x_449;
	wire x_450;
	wire x_451;
	wire x_452;
	wire x_453;
	wire x_454;
	wire x_455;
	wire x_456;
	wire x_457;
	wire x_458;
	wire x_459;
	wire x_460;
	wire x_461;
	wire x_462;
	wire x_463;
	wire x_464;
	wire x_465;
	wire x_466;
	wire x_467;
	wire x_468;
	wire x_469;
	wire x_470;
	wire x_471;
	wire x_472;
	wire x_473;
	output o_1;
	assign v_171 = 0 ;
	assign v_168 = 0 ;
	assign v_166 = 0 ;
	assign v_162 = 0 ;
	assign v_159 = 0 ;
	assign v_156 = 0 ;
	assign v_153 = 0 ;
	assign v_150 = 0 ;
	assign v_147 = 0 ;
	assign v_144 = 0 ;
	assign v_140 = 0 ;
	assign v_137 = 0 ;
	assign v_134 = 0 ;
	assign v_131 = 0 ;
	assign v_127 = 0 ;
	assign v_124 = 0 ;
	assign v_120 = 0 ;
	assign v_117 = 0 ;
	assign v_113 = 0 ;
	assign v_110 = 0 ;
	assign v_106 = 0 ;
	assign v_103 = 0 ;
	assign v_100 = 0 ;
	assign v_97 = 0 ;
	assign v_93 = 0 ;
	assign v_90 = 0 ;
	assign v_86 = 0 ;
	assign v_83 = 0 ;
	assign v_81 = 0 ;
	assign v_77 = 0 ;
	assign v_72 = 0 ;
	assign v_5 = 0 ;
	assign v_1 = 0 ;
	assign v_2 = 1 ;
	assign v_3 = 1 ;
	assign v_4 = 1 ;
	assign v_80 = 1 ;
	assign v_89 = 1 ;
	assign v_96 = 1 ;
	assign v_102 = 1 ;
	assign v_109 = 1 ;
	assign v_116 = 1 ;
	assign v_123 = 1 ;
	assign v_130 = 1 ;
	assign v_136 = 1 ;
	assign v_143 = 1 ;
	assign v_149 = 1 ;
	assign v_155 = 1 ;
	assign v_165 = 1 ;
	assign v_173 = 1 ;
	assign v_174 = 1 ;
	assign v_175 = 1 ;
	assign v_176 = 1 ;
	assign v_177 = 1 ;
	assign v_178 = 1 ;
	assign v_179 = 1 ;
	assign v_180 = 1 ;
	assign v_181 = 1 ;
	assign v_182 = 1 ;
	assign v_183 = 1 ;
	assign v_184 = 1 ;
	assign v_185 = 1 ;
	assign v_186 = 1 ;
	assign v_283 = 1 ;
	assign v_6 = v_252 ;
	assign v_10 = (~v_11 & v_70) ;
	assign v_22 = (~v_23 & v_69) ;
	assign v_42 = (~v_43 & v_68) ;
	assign v_50 = (~v_51 & v_67) ;
	assign v_54 = (~v_55 & v_66) ;
	assign v_62 = (~v_63 & v_65) ;
	assign v_64 = (v_247 & v_248) ;
	assign v_75 = ~v_73 ;
	assign v_78 = v_253 ;
	assign v_82 = v_254 ;
	assign v_84 = v_255 ;
	assign v_87 = v_256 ;
	assign v_91 = v_257 ;
	assign v_94 = v_258 ;
	assign v_98 = v_259 ;
	assign v_101 = v_260 ;
	assign v_104 = v_261 ;
	assign v_107 = v_262 ;
	assign v_111 = v_263 ;
	assign v_114 = v_264 ;
	assign v_118 = v_265 ;
	assign v_121 = v_266 ;
	assign v_125 = v_267 ;
	assign v_128 = v_268 ;
	assign v_132 = v_269 ;
	assign v_135 = v_270 ;
	assign v_138 = v_271 ;
	assign v_141 = v_272 ;
	assign v_145 = v_273 ;
	assign v_148 = v_274 ;
	assign v_151 = v_275 ;
	assign v_154 = v_276 ;
	assign v_157 = v_277 ;
	assign v_160 = v_278 ;
	assign v_163 = v_279 ;
	assign v_167 = v_280 ;
	assign v_169 = v_281 ;
	assign v_172 = v_282 ;
	assign v_11 = (v_82 ^ ~v_70) ;
	assign v_23 = (v_101 ^ ~v_69) ;
	assign v_43 = (v_135 ^ ~v_68) ;
	assign v_51 = (v_148 ^ ~v_67) ;
	assign v_55 = (v_154 ^ ~v_66) ;
	assign v_63 = (v_167 ^ ~v_65) ;
	assign v_65 = (v_243 ^ v_244) ;
	assign v_66 = (v_235 ^ v_236) ;
	assign v_67 = (v_231 ^ v_232) ;
	assign v_68 = (v_223 ^ v_224) ;
	assign v_69 = (v_203 ^ v_204) ;
	assign v_70 = (v_191 ^ v_192) ;
	assign v_71 = (v_6 ^ ~v_7) ;
	assign v_76 = (v_75 ^ v_251) ;
	assign v_79 = (v_78 ^ ~v_9) ;
	assign v_85 = (v_84 ^ ~v_13) ;
	assign v_88 = (v_87 ^ ~v_15) ;
	assign v_92 = (v_91 ^ ~v_17) ;
	assign v_95 = (v_94 ^ ~v_19) ;
	assign v_99 = (v_98 ^ ~v_21) ;
	assign v_105 = (v_104 ^ ~v_25) ;
	assign v_108 = (v_107 ^ ~v_27) ;
	assign v_112 = (v_111 ^ ~v_29) ;
	assign v_115 = (v_114 ^ ~v_31) ;
	assign v_119 = (v_118 ^ ~v_33) ;
	assign v_122 = (v_121 ^ ~v_35) ;
	assign v_126 = (v_125 ^ ~v_37) ;
	assign v_129 = (v_128 ^ ~v_39) ;
	assign v_133 = (v_132 ^ ~v_41) ;
	assign v_139 = (v_138 ^ ~v_45) ;
	assign v_142 = (v_141 ^ ~v_47) ;
	assign v_146 = (v_145 ^ ~v_49) ;
	assign v_152 = (v_151 ^ ~v_53) ;
	assign v_158 = (v_157 ^ ~v_57) ;
	assign v_161 = (v_160 ^ ~v_59) ;
	assign v_164 = (v_163 ^ ~v_61) ;
	assign v_170 = (v_169 ^ v_64) ;
	assign v_187 = (v_71 ^ v_188) ;
	assign v_189 = (v_79 ^ v_190) ;
	assign v_193 = (v_85 ^ v_194) ;
	assign v_195 = (v_88 ^ v_196) ;
	assign v_197 = (v_92 ^ v_198) ;
	assign v_199 = (v_95 ^ v_200) ;
	assign v_201 = (v_99 ^ v_202) ;
	assign v_205 = (v_105 ^ v_206) ;
	assign v_207 = (v_108 ^ v_208) ;
	assign v_209 = (v_112 ^ v_210) ;
	assign v_211 = (v_115 ^ v_212) ;
	assign v_213 = (v_119 ^ v_214) ;
	assign v_215 = (v_122 ^ v_216) ;
	assign v_217 = (v_126 ^ v_218) ;
	assign v_219 = (v_129 ^ v_220) ;
	assign v_221 = (v_133 ^ v_222) ;
	assign v_225 = (v_139 ^ v_226) ;
	assign v_227 = (v_142 ^ v_228) ;
	assign v_229 = (v_146 ^ v_230) ;
	assign v_233 = (v_152 ^ v_234) ;
	assign v_237 = (v_158 ^ v_238) ;
	assign v_239 = (v_161 ^ v_240) ;
	assign v_241 = (v_164 ^ v_242) ;
	assign v_245 = (v_170 ^ v_246) ;
	assign v_247 = (v_172 ^ v_248) ;
	assign v_249 = (v_76 ^ v_250) ;
	assign x_1 = ((v_7 | v_189) | v_8) ;
	assign x_2 = ((v_7 | v_190) | v_8) ;
	assign x_3 = (~v_7 | ~v_8) ;
	assign x_4 = ((~v_7 | ~v_189) | ~v_190) ;
	assign x_5 = (((v_8 | v_189) | ~v_190) | v_9) ;
	assign x_6 = (((v_8 | ~v_189) | v_190) | v_9) ;
	assign x_7 = (~v_8 | ~v_9) ;
	assign x_8 = ((~v_8 | v_189) | v_190) ;
	assign x_9 = ((~v_8 | ~v_189) | ~v_190) ;
	assign x_10 = ((v_9 | v_191) | v_10) ;
	assign x_11 = ((v_9 | v_192) | v_10) ;
	assign x_12 = (~v_9 | ~v_10) ;
	assign x_13 = ((~v_9 | ~v_191) | ~v_192) ;
	assign x_14 = ((v_11 | v_193) | v_12) ;
	assign x_15 = ((v_11 | v_194) | v_12) ;
	assign x_16 = (~v_11 | ~v_12) ;
	assign x_17 = ((~v_11 | ~v_193) | ~v_194) ;
	assign x_18 = (((v_12 | v_193) | ~v_194) | v_13) ;
	assign x_19 = (((v_12 | ~v_193) | v_194) | v_13) ;
	assign x_20 = (~v_12 | ~v_13) ;
	assign x_21 = ((~v_12 | v_193) | v_194) ;
	assign x_22 = ((~v_12 | ~v_193) | ~v_194) ;
	assign x_23 = ((v_13 | v_195) | v_14) ;
	assign x_24 = ((v_13 | v_196) | v_14) ;
	assign x_25 = (~v_13 | ~v_14) ;
	assign x_26 = ((~v_13 | ~v_195) | ~v_196) ;
	assign x_27 = (((v_14 | v_195) | ~v_196) | v_15) ;
	assign x_28 = (((v_14 | ~v_195) | v_196) | v_15) ;
	assign x_29 = (~v_14 | ~v_15) ;
	assign x_30 = ((~v_14 | v_195) | v_196) ;
	assign x_31 = ((~v_14 | ~v_195) | ~v_196) ;
	assign x_32 = ((v_15 | v_197) | v_16) ;
	assign x_33 = ((v_15 | v_198) | v_16) ;
	assign x_34 = (~v_15 | ~v_16) ;
	assign x_35 = ((~v_15 | ~v_197) | ~v_198) ;
	assign x_36 = (((v_16 | v_197) | ~v_198) | v_17) ;
	assign x_37 = (((v_16 | ~v_197) | v_198) | v_17) ;
	assign x_38 = (~v_16 | ~v_17) ;
	assign x_39 = ((~v_16 | v_197) | v_198) ;
	assign x_40 = ((~v_16 | ~v_197) | ~v_198) ;
	assign x_41 = ((v_17 | v_199) | v_18) ;
	assign x_42 = ((v_17 | v_200) | v_18) ;
	assign x_43 = (~v_17 | ~v_18) ;
	assign x_44 = ((~v_17 | ~v_199) | ~v_200) ;
	assign x_45 = (((v_18 | v_199) | ~v_200) | v_19) ;
	assign x_46 = (((v_18 | ~v_199) | v_200) | v_19) ;
	assign x_47 = (~v_18 | ~v_19) ;
	assign x_48 = ((~v_18 | v_199) | v_200) ;
	assign x_49 = ((~v_18 | ~v_199) | ~v_200) ;
	assign x_50 = ((v_19 | v_201) | v_20) ;
	assign x_51 = ((v_19 | v_202) | v_20) ;
	assign x_52 = (~v_19 | ~v_20) ;
	assign x_53 = ((~v_19 | ~v_201) | ~v_202) ;
	assign x_54 = (((v_20 | v_201) | ~v_202) | v_21) ;
	assign x_55 = (((v_20 | ~v_201) | v_202) | v_21) ;
	assign x_56 = (~v_20 | ~v_21) ;
	assign x_57 = ((~v_20 | v_201) | v_202) ;
	assign x_58 = ((~v_20 | ~v_201) | ~v_202) ;
	assign x_59 = ((v_21 | v_203) | v_22) ;
	assign x_60 = ((v_21 | v_204) | v_22) ;
	assign x_61 = (~v_21 | ~v_22) ;
	assign x_62 = ((~v_21 | ~v_203) | ~v_204) ;
	assign x_63 = ((v_23 | v_205) | v_24) ;
	assign x_64 = ((v_23 | v_206) | v_24) ;
	assign x_65 = (~v_23 | ~v_24) ;
	assign x_66 = ((~v_23 | ~v_205) | ~v_206) ;
	assign x_67 = (((v_24 | v_205) | ~v_206) | v_25) ;
	assign x_68 = (((v_24 | ~v_205) | v_206) | v_25) ;
	assign x_69 = (~v_24 | ~v_25) ;
	assign x_70 = ((~v_24 | v_205) | v_206) ;
	assign x_71 = ((~v_24 | ~v_205) | ~v_206) ;
	assign x_72 = ((v_25 | v_207) | v_26) ;
	assign x_73 = ((v_25 | v_208) | v_26) ;
	assign x_74 = (~v_25 | ~v_26) ;
	assign x_75 = ((~v_25 | ~v_207) | ~v_208) ;
	assign x_76 = (((v_26 | v_207) | ~v_208) | v_27) ;
	assign x_77 = (((v_26 | ~v_207) | v_208) | v_27) ;
	assign x_78 = (~v_26 | ~v_27) ;
	assign x_79 = ((~v_26 | v_207) | v_208) ;
	assign x_80 = ((~v_26 | ~v_207) | ~v_208) ;
	assign x_81 = ((v_27 | v_209) | v_28) ;
	assign x_82 = ((v_27 | v_210) | v_28) ;
	assign x_83 = (~v_27 | ~v_28) ;
	assign x_84 = ((~v_27 | ~v_209) | ~v_210) ;
	assign x_85 = (((v_28 | v_209) | ~v_210) | v_29) ;
	assign x_86 = (((v_28 | ~v_209) | v_210) | v_29) ;
	assign x_87 = (~v_28 | ~v_29) ;
	assign x_88 = ((~v_28 | v_209) | v_210) ;
	assign x_89 = ((~v_28 | ~v_209) | ~v_210) ;
	assign x_90 = ((v_29 | v_211) | v_30) ;
	assign x_91 = ((v_29 | v_212) | v_30) ;
	assign x_92 = (~v_29 | ~v_30) ;
	assign x_93 = ((~v_29 | ~v_211) | ~v_212) ;
	assign x_94 = (((v_30 | v_211) | ~v_212) | v_31) ;
	assign x_95 = (((v_30 | ~v_211) | v_212) | v_31) ;
	assign x_96 = (~v_30 | ~v_31) ;
	assign x_97 = ((~v_30 | v_211) | v_212) ;
	assign x_98 = ((~v_30 | ~v_211) | ~v_212) ;
	assign x_99 = ((v_31 | v_213) | v_32) ;
	assign x_100 = ((v_31 | v_214) | v_32) ;
	assign x_101 = (~v_31 | ~v_32) ;
	assign x_102 = ((~v_31 | ~v_213) | ~v_214) ;
	assign x_103 = (((v_32 | v_213) | ~v_214) | v_33) ;
	assign x_104 = (((v_32 | ~v_213) | v_214) | v_33) ;
	assign x_105 = (~v_32 | ~v_33) ;
	assign x_106 = ((~v_32 | v_213) | v_214) ;
	assign x_107 = ((~v_32 | ~v_213) | ~v_214) ;
	assign x_108 = ((v_33 | v_215) | v_34) ;
	assign x_109 = ((v_33 | v_216) | v_34) ;
	assign x_110 = (~v_33 | ~v_34) ;
	assign x_111 = ((~v_33 | ~v_215) | ~v_216) ;
	assign x_112 = (((v_34 | v_215) | ~v_216) | v_35) ;
	assign x_113 = (((v_34 | ~v_215) | v_216) | v_35) ;
	assign x_114 = (~v_34 | ~v_35) ;
	assign x_115 = ((~v_34 | v_215) | v_216) ;
	assign x_116 = ((~v_34 | ~v_215) | ~v_216) ;
	assign x_117 = ((v_35 | v_217) | v_36) ;
	assign x_118 = ((v_35 | v_218) | v_36) ;
	assign x_119 = (~v_35 | ~v_36) ;
	assign x_120 = ((~v_35 | ~v_217) | ~v_218) ;
	assign x_121 = (((v_36 | v_217) | ~v_218) | v_37) ;
	assign x_122 = (((v_36 | ~v_217) | v_218) | v_37) ;
	assign x_123 = (~v_36 | ~v_37) ;
	assign x_124 = ((~v_36 | v_217) | v_218) ;
	assign x_125 = ((~v_36 | ~v_217) | ~v_218) ;
	assign x_126 = ((v_37 | v_219) | v_38) ;
	assign x_127 = ((v_37 | v_220) | v_38) ;
	assign x_128 = (~v_37 | ~v_38) ;
	assign x_129 = ((~v_37 | ~v_219) | ~v_220) ;
	assign x_130 = (((v_38 | v_219) | ~v_220) | v_39) ;
	assign x_131 = (((v_38 | ~v_219) | v_220) | v_39) ;
	assign x_132 = (~v_38 | ~v_39) ;
	assign x_133 = ((~v_38 | v_219) | v_220) ;
	assign x_134 = ((~v_38 | ~v_219) | ~v_220) ;
	assign x_135 = ((v_39 | v_221) | v_40) ;
	assign x_136 = ((v_39 | v_222) | v_40) ;
	assign x_137 = (~v_39 | ~v_40) ;
	assign x_138 = ((~v_39 | ~v_221) | ~v_222) ;
	assign x_139 = (((v_40 | v_221) | ~v_222) | v_41) ;
	assign x_140 = (((v_40 | ~v_221) | v_222) | v_41) ;
	assign x_141 = (~v_40 | ~v_41) ;
	assign x_142 = ((~v_40 | v_221) | v_222) ;
	assign x_143 = ((~v_40 | ~v_221) | ~v_222) ;
	assign x_144 = ((v_41 | v_223) | v_42) ;
	assign x_145 = ((v_41 | v_224) | v_42) ;
	assign x_146 = (~v_41 | ~v_42) ;
	assign x_147 = ((~v_41 | ~v_223) | ~v_224) ;
	assign x_148 = ((v_43 | v_225) | v_44) ;
	assign x_149 = ((v_43 | v_226) | v_44) ;
	assign x_150 = (~v_43 | ~v_44) ;
	assign x_151 = ((~v_43 | ~v_225) | ~v_226) ;
	assign x_152 = (((v_44 | v_225) | ~v_226) | v_45) ;
	assign x_153 = (((v_44 | ~v_225) | v_226) | v_45) ;
	assign x_154 = (~v_44 | ~v_45) ;
	assign x_155 = ((~v_44 | v_225) | v_226) ;
	assign x_156 = ((~v_44 | ~v_225) | ~v_226) ;
	assign x_157 = ((v_45 | v_227) | v_46) ;
	assign x_158 = ((v_45 | v_228) | v_46) ;
	assign x_159 = (~v_45 | ~v_46) ;
	assign x_160 = ((~v_45 | ~v_227) | ~v_228) ;
	assign x_161 = (((v_46 | v_227) | ~v_228) | v_47) ;
	assign x_162 = (((v_46 | ~v_227) | v_228) | v_47) ;
	assign x_163 = (~v_46 | ~v_47) ;
	assign x_164 = ((~v_46 | v_227) | v_228) ;
	assign x_165 = ((~v_46 | ~v_227) | ~v_228) ;
	assign x_166 = ((v_47 | v_229) | v_48) ;
	assign x_167 = ((v_47 | v_230) | v_48) ;
	assign x_168 = (~v_47 | ~v_48) ;
	assign x_169 = ((~v_47 | ~v_229) | ~v_230) ;
	assign x_170 = (((v_48 | v_229) | ~v_230) | v_49) ;
	assign x_171 = (((v_48 | ~v_229) | v_230) | v_49) ;
	assign x_172 = (~v_48 | ~v_49) ;
	assign x_173 = ((~v_48 | v_229) | v_230) ;
	assign x_174 = ((~v_48 | ~v_229) | ~v_230) ;
	assign x_175 = ((v_49 | v_231) | v_50) ;
	assign x_176 = ((v_49 | v_232) | v_50) ;
	assign x_177 = (~v_49 | ~v_50) ;
	assign x_178 = ((~v_49 | ~v_231) | ~v_232) ;
	assign x_179 = ((v_51 | v_233) | v_52) ;
	assign x_180 = ((v_51 | v_234) | v_52) ;
	assign x_181 = (~v_51 | ~v_52) ;
	assign x_182 = ((~v_51 | ~v_233) | ~v_234) ;
	assign x_183 = (((v_52 | v_233) | ~v_234) | v_53) ;
	assign x_184 = (((v_52 | ~v_233) | v_234) | v_53) ;
	assign x_185 = (~v_52 | ~v_53) ;
	assign x_186 = ((~v_52 | v_233) | v_234) ;
	assign x_187 = ((~v_52 | ~v_233) | ~v_234) ;
	assign x_188 = ((v_53 | v_235) | v_54) ;
	assign x_189 = ((v_53 | v_236) | v_54) ;
	assign x_190 = (~v_53 | ~v_54) ;
	assign x_191 = ((~v_53 | ~v_235) | ~v_236) ;
	assign x_192 = ((v_55 | v_237) | v_56) ;
	assign x_193 = ((v_55 | v_238) | v_56) ;
	assign x_194 = (~v_55 | ~v_56) ;
	assign x_195 = ((~v_55 | ~v_237) | ~v_238) ;
	assign x_196 = (((v_56 | v_237) | ~v_238) | v_57) ;
	assign x_197 = (((v_56 | ~v_237) | v_238) | v_57) ;
	assign x_198 = (~v_56 | ~v_57) ;
	assign x_199 = ((~v_56 | v_237) | v_238) ;
	assign x_200 = ((~v_56 | ~v_237) | ~v_238) ;
	assign x_201 = ((v_57 | v_239) | v_58) ;
	assign x_202 = ((v_57 | v_240) | v_58) ;
	assign x_203 = (~v_57 | ~v_58) ;
	assign x_204 = ((~v_57 | ~v_239) | ~v_240) ;
	assign x_205 = (((v_58 | v_239) | ~v_240) | v_59) ;
	assign x_206 = (((v_58 | ~v_239) | v_240) | v_59) ;
	assign x_207 = (~v_58 | ~v_59) ;
	assign x_208 = ((~v_58 | v_239) | v_240) ;
	assign x_209 = ((~v_58 | ~v_239) | ~v_240) ;
	assign x_210 = ((v_59 | v_241) | v_60) ;
	assign x_211 = ((v_59 | v_242) | v_60) ;
	assign x_212 = (~v_59 | ~v_60) ;
	assign x_213 = ((~v_59 | ~v_241) | ~v_242) ;
	assign x_214 = (((v_60 | v_241) | ~v_242) | v_61) ;
	assign x_215 = (((v_60 | ~v_241) | v_242) | v_61) ;
	assign x_216 = (~v_60 | ~v_61) ;
	assign x_217 = ((~v_60 | v_241) | v_242) ;
	assign x_218 = ((~v_60 | ~v_241) | ~v_242) ;
	assign x_219 = ((v_61 | v_243) | v_62) ;
	assign x_220 = ((v_61 | v_244) | v_62) ;
	assign x_221 = (~v_61 | ~v_62) ;
	assign x_222 = ((~v_61 | ~v_243) | ~v_244) ;
	assign x_223 = ((v_63 | v_245) | v_64) ;
	assign x_224 = ((v_63 | v_246) | v_64) ;
	assign x_225 = ((v_63 | v_245) | v_246) ;
	assign x_226 = ((~v_63 | ~v_245) | ~v_246) ;
	assign x_227 = ((~v_63 | ~v_246) | ~v_64) ;
	assign x_228 = ((~v_63 | ~v_245) | ~v_64) ;
	assign x_229 = ((v_73 | v_187) | v_74) ;
	assign x_230 = ((v_73 | v_188) | v_74) ;
	assign x_231 = (~v_73 | ~v_74) ;
	assign x_232 = ((~v_73 | ~v_187) | ~v_188) ;
	assign x_233 = (((v_74 | v_187) | ~v_188) | v_7) ;
	assign x_234 = (((v_74 | ~v_187) | v_188) | v_7) ;
	assign x_235 = (~v_74 | ~v_7) ;
	assign x_236 = ((~v_74 | v_187) | v_188) ;
	assign x_237 = ((~v_74 | ~v_187) | ~v_188) ;
	assign x_238 = (x_2 & x_3) ;
	assign x_239 = (x_1 & x_238) ;
	assign x_240 = (x_4 & x_5) ;
	assign x_241 = (x_6 & x_7) ;
	assign x_242 = (x_240 & x_241) ;
	assign x_243 = (x_239 & x_242) ;
	assign x_244 = (x_9 & x_10) ;
	assign x_245 = (x_8 & x_244) ;
	assign x_246 = (x_11 & x_12) ;
	assign x_247 = (x_13 & x_14) ;
	assign x_248 = (x_246 & x_247) ;
	assign x_249 = (x_245 & x_248) ;
	assign x_250 = (x_243 & x_249) ;
	assign x_251 = (x_16 & x_17) ;
	assign x_252 = (x_15 & x_251) ;
	assign x_253 = (x_18 & x_19) ;
	assign x_254 = (x_20 & x_21) ;
	assign x_255 = (x_253 & x_254) ;
	assign x_256 = (x_252 & x_255) ;
	assign x_257 = (x_22 & x_23) ;
	assign x_258 = (x_24 & x_25) ;
	assign x_259 = (x_257 & x_258) ;
	assign x_260 = (x_26 & x_27) ;
	assign x_261 = (x_28 & x_29) ;
	assign x_262 = (x_260 & x_261) ;
	assign x_263 = (x_259 & x_262) ;
	assign x_264 = (x_256 & x_263) ;
	assign x_265 = (x_250 & x_264) ;
	assign x_266 = (x_31 & x_32) ;
	assign x_267 = (x_30 & x_266) ;
	assign x_268 = (x_33 & x_34) ;
	assign x_269 = (x_35 & x_36) ;
	assign x_270 = (x_268 & x_269) ;
	assign x_271 = (x_267 & x_270) ;
	assign x_272 = (x_37 & x_38) ;
	assign x_273 = (x_39 & x_40) ;
	assign x_274 = (x_272 & x_273) ;
	assign x_275 = (x_41 & x_42) ;
	assign x_276 = (x_43 & x_44) ;
	assign x_277 = (x_275 & x_276) ;
	assign x_278 = (x_274 & x_277) ;
	assign x_279 = (x_271 & x_278) ;
	assign x_280 = (x_46 & x_47) ;
	assign x_281 = (x_45 & x_280) ;
	assign x_282 = (x_48 & x_49) ;
	assign x_283 = (x_50 & x_51) ;
	assign x_284 = (x_282 & x_283) ;
	assign x_285 = (x_281 & x_284) ;
	assign x_286 = (x_52 & x_53) ;
	assign x_287 = (x_54 & x_55) ;
	assign x_288 = (x_286 & x_287) ;
	assign x_289 = (x_56 & x_57) ;
	assign x_290 = (x_58 & x_59) ;
	assign x_291 = (x_289 & x_290) ;
	assign x_292 = (x_288 & x_291) ;
	assign x_293 = (x_285 & x_292) ;
	assign x_294 = (x_279 & x_293) ;
	assign x_295 = (x_265 & x_294) ;
	assign x_296 = (x_61 & x_62) ;
	assign x_297 = (x_60 & x_296) ;
	assign x_298 = (x_63 & x_64) ;
	assign x_299 = (x_65 & x_66) ;
	assign x_300 = (x_298 & x_299) ;
	assign x_301 = (x_297 & x_300) ;
	assign x_302 = (x_68 & x_69) ;
	assign x_303 = (x_67 & x_302) ;
	assign x_304 = (x_70 & x_71) ;
	assign x_305 = (x_72 & x_73) ;
	assign x_306 = (x_304 & x_305) ;
	assign x_307 = (x_303 & x_306) ;
	assign x_308 = (x_301 & x_307) ;
	assign x_309 = (x_75 & x_76) ;
	assign x_310 = (x_74 & x_309) ;
	assign x_311 = (x_77 & x_78) ;
	assign x_312 = (x_79 & x_80) ;
	assign x_313 = (x_311 & x_312) ;
	assign x_314 = (x_310 & x_313) ;
	assign x_315 = (x_81 & x_82) ;
	assign x_316 = (x_83 & x_84) ;
	assign x_317 = (x_315 & x_316) ;
	assign x_318 = (x_85 & x_86) ;
	assign x_319 = (x_87 & x_88) ;
	assign x_320 = (x_318 & x_319) ;
	assign x_321 = (x_317 & x_320) ;
	assign x_322 = (x_314 & x_321) ;
	assign x_323 = (x_308 & x_322) ;
	assign x_324 = (x_90 & x_91) ;
	assign x_325 = (x_89 & x_324) ;
	assign x_326 = (x_92 & x_93) ;
	assign x_327 = (x_94 & x_95) ;
	assign x_328 = (x_326 & x_327) ;
	assign x_329 = (x_325 & x_328) ;
	assign x_330 = (x_96 & x_97) ;
	assign x_331 = (x_98 & x_99) ;
	assign x_332 = (x_330 & x_331) ;
	assign x_333 = (x_100 & x_101) ;
	assign x_334 = (x_102 & x_103) ;
	assign x_335 = (x_333 & x_334) ;
	assign x_336 = (x_332 & x_335) ;
	assign x_337 = (x_329 & x_336) ;
	assign x_338 = (x_105 & x_106) ;
	assign x_339 = (x_104 & x_338) ;
	assign x_340 = (x_107 & x_108) ;
	assign x_341 = (x_109 & x_110) ;
	assign x_342 = (x_340 & x_341) ;
	assign x_343 = (x_339 & x_342) ;
	assign x_344 = (x_111 & x_112) ;
	assign x_345 = (x_113 & x_114) ;
	assign x_346 = (x_344 & x_345) ;
	assign x_347 = (x_115 & x_116) ;
	assign x_348 = (x_117 & x_118) ;
	assign x_349 = (x_347 & x_348) ;
	assign x_350 = (x_346 & x_349) ;
	assign x_351 = (x_343 & x_350) ;
	assign x_352 = (x_337 & x_351) ;
	assign x_353 = (x_323 & x_352) ;
	assign x_354 = (x_295 & x_353) ;
	assign x_355 = (x_120 & x_121) ;
	assign x_356 = (x_119 & x_355) ;
	assign x_357 = (x_122 & x_123) ;
	assign x_358 = (x_124 & x_125) ;
	assign x_359 = (x_357 & x_358) ;
	assign x_360 = (x_356 & x_359) ;
	assign x_361 = (x_127 & x_128) ;
	assign x_362 = (x_126 & x_361) ;
	assign x_363 = (x_129 & x_130) ;
	assign x_364 = (x_131 & x_132) ;
	assign x_365 = (x_363 & x_364) ;
	assign x_366 = (x_362 & x_365) ;
	assign x_367 = (x_360 & x_366) ;
	assign x_368 = (x_134 & x_135) ;
	assign x_369 = (x_133 & x_368) ;
	assign x_370 = (x_136 & x_137) ;
	assign x_371 = (x_138 & x_139) ;
	assign x_372 = (x_370 & x_371) ;
	assign x_373 = (x_369 & x_372) ;
	assign x_374 = (x_140 & x_141) ;
	assign x_375 = (x_142 & x_143) ;
	assign x_376 = (x_374 & x_375) ;
	assign x_377 = (x_144 & x_145) ;
	assign x_378 = (x_146 & x_147) ;
	assign x_379 = (x_377 & x_378) ;
	assign x_380 = (x_376 & x_379) ;
	assign x_381 = (x_373 & x_380) ;
	assign x_382 = (x_367 & x_381) ;
	assign x_383 = (x_149 & x_150) ;
	assign x_384 = (x_148 & x_383) ;
	assign x_385 = (x_151 & x_152) ;
	assign x_386 = (x_153 & x_154) ;
	assign x_387 = (x_385 & x_386) ;
	assign x_388 = (x_384 & x_387) ;
	assign x_389 = (x_155 & x_156) ;
	assign x_390 = (x_157 & x_158) ;
	assign x_391 = (x_389 & x_390) ;
	assign x_392 = (x_159 & x_160) ;
	assign x_393 = (x_161 & x_162) ;
	assign x_394 = (x_392 & x_393) ;
	assign x_395 = (x_391 & x_394) ;
	assign x_396 = (x_388 & x_395) ;
	assign x_397 = (x_164 & x_165) ;
	assign x_398 = (x_163 & x_397) ;
	assign x_399 = (x_166 & x_167) ;
	assign x_400 = (x_168 & x_169) ;
	assign x_401 = (x_399 & x_400) ;
	assign x_402 = (x_398 & x_401) ;
	assign x_403 = (x_170 & x_171) ;
	assign x_404 = (x_172 & x_173) ;
	assign x_405 = (x_403 & x_404) ;
	assign x_406 = (x_174 & x_175) ;
	assign x_407 = (x_176 & x_177) ;
	assign x_408 = (x_406 & x_407) ;
	assign x_409 = (x_405 & x_408) ;
	assign x_410 = (x_402 & x_409) ;
	assign x_411 = (x_396 & x_410) ;
	assign x_412 = (x_382 & x_411) ;
	assign x_413 = (x_179 & x_180) ;
	assign x_414 = (x_178 & x_413) ;
	assign x_415 = (x_181 & x_182) ;
	assign x_416 = (x_183 & x_184) ;
	assign x_417 = (x_415 & x_416) ;
	assign x_418 = (x_414 & x_417) ;
	assign x_419 = (x_185 & x_186) ;
	assign x_420 = (x_187 & x_188) ;
	assign x_421 = (x_419 & x_420) ;
	assign x_422 = (x_189 & x_190) ;
	assign x_423 = (x_191 & x_192) ;
	assign x_424 = (x_422 & x_423) ;
	assign x_425 = (x_421 & x_424) ;
	assign x_426 = (x_418 & x_425) ;
	assign x_427 = (x_194 & x_195) ;
	assign x_428 = (x_193 & x_427) ;
	assign x_429 = (x_196 & x_197) ;
	assign x_430 = (x_198 & x_199) ;
	assign x_431 = (x_429 & x_430) ;
	assign x_432 = (x_428 & x_431) ;
	assign x_433 = (x_200 & x_201) ;
	assign x_434 = (x_202 & x_203) ;
	assign x_435 = (x_433 & x_434) ;
	assign x_436 = (x_204 & x_205) ;
	assign x_437 = (x_206 & x_207) ;
	assign x_438 = (x_436 & x_437) ;
	assign x_439 = (x_435 & x_438) ;
	assign x_440 = (x_432 & x_439) ;
	assign x_441 = (x_426 & x_440) ;
	assign x_442 = (x_209 & x_210) ;
	assign x_443 = (x_208 & x_442) ;
	assign x_444 = (x_211 & x_212) ;
	assign x_445 = (x_213 & x_214) ;
	assign x_446 = (x_444 & x_445) ;
	assign x_447 = (x_443 & x_446) ;
	assign x_448 = (x_215 & x_216) ;
	assign x_449 = (x_217 & x_218) ;
	assign x_450 = (x_448 & x_449) ;
	assign x_451 = (x_219 & x_220) ;
	assign x_452 = (x_221 & x_222) ;
	assign x_453 = (x_451 & x_452) ;
	assign x_454 = (x_450 & x_453) ;
	assign x_455 = (x_447 & x_454) ;
	assign x_456 = (x_224 & x_225) ;
	assign x_457 = (x_223 & x_456) ;
	assign x_458 = (x_226 & x_227) ;
	assign x_459 = (x_228 & x_229) ;
	assign x_460 = (x_458 & x_459) ;
	assign x_461 = (x_457 & x_460) ;
	assign x_462 = (x_230 & x_231) ;
	assign x_463 = (x_232 & x_233) ;
	assign x_464 = (x_462 & x_463) ;
	assign x_465 = (x_234 & x_235) ;
	assign x_466 = (x_236 & x_237) ;
	assign x_467 = (x_465 & x_466) ;
	assign x_468 = (x_464 & x_467) ;
	assign x_469 = (x_461 & x_468) ;
	assign x_470 = (x_455 & x_469) ;
	assign x_471 = (x_441 & x_470) ;
	assign x_472 = (x_412 & x_471) ;
	assign x_473 = (x_354 & x_472) ;
	assign o_1 = x_473 ;
endmodule
