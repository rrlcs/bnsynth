module formula_simplified(i2[11],i2[10],i2[9],i2[8],i2[7],i2[6],i1[11],i1[10],i1[9],i1[8],i1[7],i1[6],a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],o_1);
	input i2;
	i2;
	i2;
	i2;
	i2;
	i2;
	i1;
	i1;
	i1;
	i1;
	i1;
	i1;
	a;
	a;
	a;
	a;
	a;
	a;
	a;
	a;
	a;
	a;
	a;
	a;
	wire n_1;
	wire n_2;
	wire n_3;
	wire n_4;
	wire n_5;
	wire n_6;
	wire n_7;
	wire n_8;
	wire n_9;
	wire n_10;
	wire n_11;
	wire n_12;
	wire n_13;
	wire n_14;
	wire n_15;
	wire n_16;
	wire n_17;
	wire n_18;
	wire n_19;
	wire n_20;
	wire n_21;
	wire n_22;
	wire n_23;
	wire n_24;
	wire n_25;
	wire n_26;
	wire n_27;
	wire n_28;
	wire n_29;
	wire n_30;
	wire n_31;
	wire n_32;
	wire n_33;
	wire n_34;
	wire n_35;
	wire n_36;
	wire n_37;
	wire n_38;
	wire n_39;
	wire n_40;
	wire n_41;
	wire n_42;
	wire n_43;
	wire n_44;
	wire n_45;
	wire n_46;
	wire n_47;
	wire n_48;
	wire n_49;
	wire n_50;
	wire n_51;
	wire n_52;
	wire n_53;
	wire n_54;
	wire n_55;
	wire n_56;
	wire n_57;
	wire n_58;
	wire n_59;
	wire n_60;
	wire n_61;
	wire n_62;
	wire n_63;
	wire n_64;
	wire n_65;
	wire n_66;
	wire n_67;
	wire n_68;
	wire n_69;
	wire n_70;
	wire n_71;
	wire n_72;
	wire n_73;
	wire n_74;
	wire n_75;
	wire n_76;
	wire n_77;
	wire n_78;
	wire n_79;
	wire n_80;
	wire n_81;
	wire n_82;
	wire n_83;
	wire n_84;
	wire n_85;
	wire n_86;
	wire n_87;
	wire n_88;
	wire n_89;
	wire n_90;
	wire n_91;
	wire n_92;
	wire n_93;
	wire n_94;
	wire n_95;
	wire n_96;
	wire n_97;
	wire n_98;
	wire n_99;
	wire n_100;
	wire n_101;
	wire n_102;
	wire n_103;
	wire n_104;
	wire n_105;
	wire n_106;
	wire n_107;
	wire n_108;
	wire n_109;
	wire n_110;
	wire n_111;
	wire n_112;
	wire n_113;
	wire n_114;
	wire n_115;
	wire n_116;
	wire n_117;
	wire n_118;
	wire n_119;
	wire n_120;
	wire n_121;
	wire n_122;
	wire n_123;
	wire n_124;
	wire n_125;
	wire n_126;
	wire n_127;
	wire n_128;
	wire n_129;
	wire n_130;
	wire n_131;
	wire n_132;
	wire n_133;
	wire n_134;
	wire n_135;
	wire n_136;
	wire n_137;
	wire n_138;
	wire n_139;
	wire n_140;
	wire n_141;
	wire n_142;
	wire n_143;
	wire n_144;
	wire n_145;
	wire n_146;
	wire n_147;
	wire n_148;
	wire n_149;
	wire n_150;
	wire n_151;
	wire n_152;
	wire n_153;
	wire n_154;
	wire n_155;
	wire n_156;
	wire n_157;
	wire n_158;
	wire n_159;
	wire n_160;
	wire n_161;
	wire n_162;
	wire n_163;
	wire n_164;
	wire n_165;
	wire n_166;
	wire n_167;
	wire n_168;
	wire n_169;
	wire n_170;
	wire n_171;
	wire n_172;
	wire n_173;
	wire n_174;
	wire n_175;
	wire n_176;
	wire n_177;
	wire n_178;
	wire n_179;
	wire n_180;
	wire n_181;
	wire n_182;
	wire n_183;
	wire n_184;
	wire n_185;
	wire n_186;
	wire n_187;
	wire n_188;
	wire n_189;
	wire n_190;
	wire n_191;
	wire n_192;
	wire n_193;
	wire n_194;
	wire n_195;
	wire n_196;
	wire n_197;
	wire n_198;
	wire n_199;
	wire n_200;
	wire n_201;
	wire n_202;
	wire n_203;
	wire n_204;
	wire n_205;
	wire n_206;
	wire n_207;
	wire n_208;
	wire n_209;
	wire n_210;
	wire n_211;
	wire n_212;
	wire n_213;
	wire n_214;
	wire n_215;
	wire n_216;
	wire n_217;
	wire n_218;
	wire n_219;
	wire n_220;
	wire n_221;
	wire n_222;
	wire n_223;
	wire n_224;
	wire n_225;
	wire n_226;
	wire n_227;
	wire n_228;
	wire n_229;
	wire n_230;
	wire n_231;
	wire n_232;
	wire n_233;
	wire n_234;
	wire n_235;
	wire n_236;
	wire n_237;
	wire n_238;
	wire n_239;
	wire n_240;
	wire n_241;
	wire n_242;
	wire n_243;
	wire n_244;
	wire n_245;
	wire n_246;
	wire n_247;
	wire n_248;
	wire n_249;
	wire n_250;
	wire n_251;
	wire n_252;
	wire n_253;
	wire n_254;
	wire n_255;
	wire n_256;
	wire n_257;
	wire n_258;
	wire n_259;
	wire n_260;
	wire n_261;
	wire n_262;
	wire n_263;
	wire n_264;
	wire n_265;
	wire n_266;
	wire n_267;
	wire n_268;
	wire n_269;
	wire n_270;
	wire n_271;
	wire n_272;
	wire n_273;
	wire n_274;
	wire n_275;
	wire n_276;
	wire n_277;
	wire n_278;
	wire n_279;
	wire n_280;
	output o_1;
	assign n_12 = (i2[8] & i1[11]);
	assign n_18 = (i2[9] & i1[11]);
	assign n_257 = (~i2[9] & ~i2[8]);
	assign n_11 = (i2[9] & i1[10]);
	assign n_8 = (i2[8] & i1[10]);
	assign n_250 = (i1[11] & ~i1[10]);
	assign n_17 = (i2[10] & i1[10]);
	assign n_14 = (i2[10] & i1[11]);
	assign n_15 = (i2[11] & i1[10]);
	assign n_245 = (i2[11] & i1[11]);
	assign n_256 = (i2[11] & ~i2[10]);
	assign n_9 = (i2[7] & i1[11]);
	assign n_5 = (i2[7] & i1[10]);
	assign n_6 = (i2[6] & i1[11]);
	assign n_33 = (i2[6] & i1[10]);
	assign n_255 = (~i2[7] & ~i2[6]);
	assign n_50 = (i2[10] & i1[9]);
	assign n_52 = (i2[11] & i1[9]);
	assign n_46 = (i2[9] & i1[9]);
	assign n_42 = (i2[8] & i1[9]);
	assign n_36 = (i2[7] & i1[9]);
	assign n_4 = (i2[6] & i1[9]);
	assign n_93 = (i2[10] & i1[8]);
	assign n_97 = (i2[11] & i1[8]);
	assign n_89 = (i2[9] & i1[8]);
	assign n_251 = (~i1[9] & ~i1[8]);
	assign n_83 = (i2[8] & i1[8]);
	assign n_79 = (i2[7] & i1[8]);
	assign n_3 = (i2[6] & i1[8]);
	assign n_134 = (i2[10] & i1[7]);
	assign n_138 = (i2[11] & i1[7]);
	assign n_128 = (i2[9] & i1[7]);
	assign n_124 = (i2[8] & i1[7]);
	assign n_120 = (i2[7] & i1[7]);
	assign n_2 = (i2[6] & i1[7]);
	assign n_249 = (~i1[7] & ~i1[6]);
	assign n_179 = (i2[11] & i1[6]);
	assign n_173 = (i2[10] & i1[6]);
	assign n_169 = (i2[9] & i1[6]);
	assign n_165 = (i2[8] & i1[6]);
	assign n_161 = (i2[7] & i1[6]);
	assign n_1 = (i2[6] & i1[6]);
	assign n_13 = (n_11 & n_12);
	assign n_21 = (~n_11 & ~n_12);
	assign n_19 = (n_17 & n_18);
	assign n_55 = (~n_17 & ~n_18);
	assign n_16 = (n_14 & n_15);
	assign n_240 = (~n_14 & ~n_15);
	assign n_247 = (a[11] & n_245);
	assign n_246 = (~a[11] & ~n_245);
	assign n_258 = (n_256 & n_257);
	assign n_10 = (n_8 & n_9);
	assign n_25 = (~n_8 & ~n_9);
	assign n_7 = (n_5 & n_6);
	assign n_29 = (~n_5 & ~n_6);
	assign n_252 = (n_250 & n_251);
	assign n_22 = (~n_21 & ~n_13);
	assign n_20 = (~n_16 & ~n_19);
	assign n_53 = (n_16 & n_19);
	assign n_241 = (~n_16 & ~n_240);
	assign n_248 = (~n_246 & ~n_247);
	assign n_259 = (n_255 & n_258);
	assign n_26 = (~n_25 & ~n_10);
	assign n_30 = (~n_29 & ~n_7);
	assign n_253 = (n_249 & n_252);
	assign n_23 = (~n_20 & n_22);
	assign n_48 = (n_20 & ~n_22);
	assign n_54 = (~n_20 & ~n_53);
	assign n_243 = (a[10] & n_241);
	assign n_242 = (~a[10] & ~n_241);
	assign n_254 = (~n_248 & ~n_253);
	assign n_24 = (~n_13 & ~n_23);
	assign n_49 = (~n_23 & ~n_48);
	assign n_56 = (~n_54 & ~n_55);
	assign n_244 = (~n_242 & ~n_243);
	assign n_260 = (n_254 & ~n_259);
	assign n_27 = (~n_24 & n_26);
	assign n_44 = (n_24 & ~n_26);
	assign n_58 = (~n_49 & ~n_50);
	assign n_51 = (n_49 & n_50);
	assign n_57 = (n_52 & n_56);
	assign n_236 = (~n_52 & ~n_56);
	assign n_261 = (~n_244 & n_260);
	assign n_28 = (~n_10 & ~n_27);
	assign n_45 = (~n_27 & ~n_44);
	assign n_59 = (~n_51 & ~n_58);
	assign n_237 = (~n_57 & ~n_236);
	assign n_31 = (~n_28 & n_30);
	assign n_40 = (n_28 & ~n_30);
	assign n_62 = (~n_45 & ~n_46);
	assign n_47 = (n_45 & n_46);
	assign n_60 = (n_57 & n_59);
	assign n_95 = (~n_57 & ~n_59);
	assign n_239 = (a[9] & ~n_237);
	assign n_238 = (~a[9] & n_237);
	assign n_32 = (~n_7 & ~n_31);
	assign n_41 = (~n_31 & ~n_40);
	assign n_63 = (~n_47 & ~n_62);
	assign n_61 = (~n_51 & ~n_60);
	assign n_96 = (~n_60 & ~n_95);
	assign n_262 = (~n_239 & n_261);
	assign n_37 = (n_32 & ~n_33);
	assign n_34 = (~n_32 & n_33);
	assign n_66 = (~n_41 & ~n_42);
	assign n_43 = (n_41 & n_42);
	assign n_64 = (~n_61 & n_63);
	assign n_91 = (n_61 & ~n_63);
	assign n_98 = (n_96 & n_97);
	assign n_232 = (~n_96 & ~n_97);
	assign n_263 = (~n_238 & n_262);
	assign n_38 = (~n_34 & ~n_37);
	assign n_74 = (~n_4 & ~n_34);
	assign n_35 = (n_4 & n_34);
	assign n_67 = (~n_43 & ~n_66);
	assign n_65 = (~n_47 & ~n_64);
	assign n_92 = (~n_64 & ~n_91);
	assign n_233 = (~n_98 & ~n_232);
	assign n_70 = (~n_36 & ~n_38);
	assign n_39 = (n_36 & n_38);
	assign n_75 = (~n_35 & ~n_74);
	assign n_68 = (~n_65 & n_67);
	assign n_87 = (n_65 & ~n_67);
	assign n_99 = (~n_92 & ~n_93);
	assign n_94 = (n_92 & n_93);
	assign n_235 = (a[8] & ~n_233);
	assign n_234 = (~a[8] & n_233);
	assign n_71 = (~n_39 & ~n_70);
	assign n_69 = (~n_43 & ~n_68);
	assign n_88 = (~n_68 & ~n_87);
	assign n_100 = (~n_94 & ~n_99);
	assign n_264 = (~n_235 & n_263);
	assign n_84 = (n_69 & ~n_71);
	assign n_72 = (~n_69 & n_71);
	assign n_103 = (~n_88 & ~n_89);
	assign n_90 = (n_88 & n_89);
	assign n_101 = (n_98 & n_100);
	assign n_136 = (~n_98 & ~n_100);
	assign n_265 = (~n_234 & n_264);
	assign n_85 = (~n_72 & ~n_84);
	assign n_73 = (~n_39 & ~n_72);
	assign n_104 = (~n_90 & ~n_103);
	assign n_102 = (~n_94 & ~n_101);
	assign n_137 = (~n_101 & ~n_136);
	assign n_107 = (~n_83 & ~n_85);
	assign n_86 = (n_83 & n_85);
	assign n_80 = (n_73 & ~n_75);
	assign n_76 = (~n_73 & n_75);
	assign n_105 = (~n_102 & n_104);
	assign n_132 = (n_102 & ~n_104);
	assign n_139 = (n_137 & n_138);
	assign n_228 = (~n_137 & ~n_138);
	assign n_108 = (~n_86 & ~n_107);
	assign n_81 = (~n_76 & ~n_80);
	assign n_77 = (~n_35 & ~n_76);
	assign n_106 = (~n_90 & ~n_105);
	assign n_133 = (~n_105 & ~n_132);
	assign n_229 = (~n_139 & ~n_228);
	assign n_111 = (~n_79 & ~n_81);
	assign n_82 = (n_79 & n_81);
	assign n_115 = (~n_3 & n_77);
	assign n_78 = (n_3 & ~n_77);
	assign n_129 = (n_106 & ~n_108);
	assign n_109 = (~n_106 & n_108);
	assign n_140 = (~n_133 & ~n_134);
	assign n_135 = (n_133 & n_134);
	assign n_231 = (a[7] & ~n_229);
	assign n_230 = (~a[7] & n_229);
	assign n_112 = (~n_82 & ~n_111);
	assign n_116 = (~n_78 & ~n_115);
	assign n_130 = (~n_109 & ~n_129);
	assign n_110 = (~n_86 & ~n_109);
	assign n_141 = (~n_135 & ~n_140);
	assign n_266 = (~n_231 & n_265);
	assign n_144 = (~n_128 & ~n_130);
	assign n_131 = (n_128 & n_130);
	assign n_125 = (n_110 & ~n_112);
	assign n_113 = (~n_110 & n_112);
	assign n_142 = (n_139 & n_141);
	assign n_177 = (~n_139 & ~n_141);
	assign n_267 = (~n_230 & n_266);
	assign n_145 = (~n_131 & ~n_144);
	assign n_126 = (~n_113 & ~n_125);
	assign n_114 = (~n_82 & ~n_113);
	assign n_143 = (~n_135 & ~n_142);
	assign n_178 = (~n_142 & ~n_177);
	assign n_148 = (~n_124 & ~n_126);
	assign n_127 = (n_124 & n_126);
	assign n_121 = (n_114 & ~n_116);
	assign n_117 = (~n_114 & n_116);
	assign n_174 = (n_143 & ~n_145);
	assign n_146 = (~n_143 & n_145);
	assign n_224 = (~n_178 & ~n_179);
	assign n_180 = (n_178 & n_179);
	assign n_149 = (~n_127 & ~n_148);
	assign n_122 = (~n_117 & ~n_121);
	assign n_118 = (~n_78 & ~n_117);
	assign n_175 = (~n_146 & ~n_174);
	assign n_147 = (~n_131 & ~n_146);
	assign n_225 = (~n_180 & ~n_224);
	assign n_152 = (~n_120 & ~n_122);
	assign n_123 = (n_120 & n_122);
	assign n_156 = (~n_2 & n_118);
	assign n_119 = (n_2 & ~n_118);
	assign n_181 = (~n_173 & ~n_175);
	assign n_176 = (n_173 & n_175);
	assign n_170 = (n_147 & ~n_149);
	assign n_150 = (~n_147 & n_149);
	assign n_227 = (a[6] & ~n_225);
	assign n_226 = (~a[6] & n_225);
	assign n_153 = (~n_123 & ~n_152);
	assign n_157 = (~n_119 & ~n_156);
	assign n_182 = (~n_176 & ~n_181);
	assign n_171 = (~n_150 & ~n_170);
	assign n_151 = (~n_127 & ~n_150);
	assign n_268 = (~n_227 & n_267);
	assign n_220 = (~n_180 & ~n_182);
	assign n_183 = (n_180 & n_182);
	assign n_185 = (~n_169 & ~n_171);
	assign n_172 = (n_169 & n_171);
	assign n_166 = (n_151 & ~n_153);
	assign n_154 = (~n_151 & n_153);
	assign n_269 = (~n_226 & n_268);
	assign n_221 = (~n_183 & ~n_220);
	assign n_184 = (~n_176 & ~n_183);
	assign n_186 = (~n_172 & ~n_185);
	assign n_167 = (~n_154 & ~n_166);
	assign n_155 = (~n_123 & ~n_154);
	assign n_223 = (a[5] & ~n_221);
	assign n_222 = (~a[5] & n_221);
	assign n_216 = (n_184 & ~n_186);
	assign n_187 = (~n_184 & n_186);
	assign n_189 = (~n_165 & ~n_167);
	assign n_168 = (n_165 & n_167);
	assign n_162 = (n_155 & ~n_157);
	assign n_158 = (~n_155 & n_157);
	assign n_270 = (~n_223 & n_269);
	assign n_217 = (~n_187 & ~n_216);
	assign n_188 = (~n_172 & ~n_187);
	assign n_190 = (~n_168 & ~n_189);
	assign n_163 = (~n_158 & ~n_162);
	assign n_159 = (~n_119 & ~n_158);
	assign n_271 = (~n_222 & n_270);
	assign n_219 = (a[4] & ~n_217);
	assign n_218 = (~a[4] & n_217);
	assign n_212 = (n_188 & ~n_190);
	assign n_191 = (~n_188 & n_190);
	assign n_193 = (~n_161 & ~n_163);
	assign n_164 = (n_161 & n_163);
	assign n_197 = (~n_1 & n_159);
	assign n_160 = (n_1 & ~n_159);
	assign n_272 = (~n_219 & n_271);
	assign n_213 = (~n_191 & ~n_212);
	assign n_192 = (~n_168 & ~n_191);
	assign n_194 = (~n_164 & ~n_193);
	assign n_198 = (~n_160 & ~n_197);
	assign n_273 = (~n_218 & n_272);
	assign n_215 = (a[3] & ~n_213);
	assign n_214 = (~a[3] & n_213);
	assign n_208 = (n_192 & ~n_194);
	assign n_195 = (~n_192 & n_194);
	assign n_274 = (~n_215 & n_273);
	assign n_209 = (~n_195 & ~n_208);
	assign n_196 = (~n_164 & ~n_195);
	assign n_275 = (~n_214 & n_274);
	assign n_211 = (a[2] & ~n_209);
	assign n_210 = (~a[2] & n_209);
	assign n_204 = (n_196 & ~n_198);
	assign n_199 = (~n_196 & n_198);
	assign n_276 = (~n_211 & n_275);
	assign n_205 = (~n_199 & ~n_204);
	assign n_200 = (~n_160 & ~n_199);
	assign n_277 = (~n_210 & n_276);
	assign n_207 = (a[1] & ~n_205);
	assign n_206 = (~a[1] & n_205);
	assign n_202 = (a[0] & ~n_200);
	assign n_201 = (~a[0] & n_200);
	assign n_278 = (~n_207 & n_277);
	assign n_203 = (~n_201 & ~n_202);
	assign n_279 = (~n_206 & n_278);
	assign n_280 = (~n_203 & n_279);
	assign o_1 = n_28);
endmodule
