// Benchmark "SKOLEMFORMULA" written by ABC on Wed Jun 30 10:48:25 2021

module SKOLEMFORMULA ( 
    i0, i1,
    i2  );
  input  i0, i1;
  output i2;
  assign i2 = 1'b1;
endmodule


