// skolem function for order file variables
// Generated using findDep.cpp 
module formula (v_1, v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_12, v_13, v_14, v_15, v_16, v_17, v_18, v_19, v_20, v_21, v_22, v_23, v_24, v_25, v_26, v_27, v_28, v_29, v_30, v_31, v_32, v_33, v_34, v_35, v_36, v_37, v_38, v_39, v_40, v_41, v_42, v_43, v_44, v_45, v_46, v_47, v_48, v_49, v_50, v_51, v_52, v_53, v_54, v_55, v_56, v_57, v_58, v_59, v_60, v_61, v_62, v_63, v_64, v_65, v_66, v_67, v_68, v_69, v_70, v_71, v_72, v_73, v_74, v_75, v_76, v_77, v_78, v_79, v_80, v_81, v_82, v_83, v_84, v_85, v_86, v_87, v_88, v_89, v_90, v_91, v_92, v_93, v_94, v_95, v_96, v_97, v_98, v_99, v_100, v_101, v_102, v_103, v_104, v_105, v_106, v_107, v_108, v_109, v_110, v_111, v_112, v_113, v_114, v_115, v_116, v_117, v_118, v_119, v_120, v_121, v_122, v_123, v_124, v_125, v_126, v_127, v_128, v_129, v_130, v_131, v_132, v_133, v_134, v_135, v_136, v_137, v_138, v_139, v_140, v_141, v_142, v_143, v_144, v_145, v_146, v_147, v_148, v_276, o_1);
input v_1;
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_13;
input v_14;
input v_15;
input v_16;
input v_17;
input v_18;
input v_19;
input v_20;
input v_21;
input v_22;
input v_23;
input v_24;
input v_25;
input v_26;
input v_27;
input v_28;
input v_29;
input v_30;
input v_31;
input v_32;
input v_33;
input v_34;
input v_35;
input v_36;
input v_37;
input v_38;
input v_39;
input v_40;
input v_41;
input v_42;
input v_43;
input v_44;
input v_45;
input v_46;
input v_47;
input v_48;
input v_49;
input v_50;
input v_51;
input v_52;
input v_53;
input v_54;
input v_55;
input v_56;
input v_57;
input v_58;
input v_59;
input v_60;
input v_61;
input v_62;
input v_63;
input v_64;
input v_65;
input v_66;
input v_67;
input v_68;
input v_69;
input v_70;
input v_71;
input v_72;
input v_73;
input v_74;
input v_75;
input v_76;
input v_77;
input v_78;
input v_79;
input v_80;
input v_81;
input v_82;
input v_83;
input v_84;
input v_85;
input v_86;
input v_87;
input v_88;
input v_89;
input v_90;
input v_91;
input v_92;
input v_93;
input v_94;
input v_95;
input v_96;
input v_97;
input v_98;
input v_99;
input v_100;
input v_101;
input v_102;
input v_103;
input v_104;
input v_105;
input v_106;
input v_107;
input v_108;
input v_109;
input v_110;
input v_111;
input v_112;
input v_113;
input v_114;
input v_115;
input v_116;
input v_117;
input v_118;
input v_119;
input v_120;
input v_121;
input v_122;
input v_123;
input v_124;
input v_125;
input v_126;
input v_127;
input v_128;
input v_129;
input v_130;
input v_131;
input v_132;
input v_133;
input v_134;
input v_135;
input v_136;
input v_137;
input v_138;
input v_139;
input v_140;
input v_141;
input v_142;
input v_143;
input v_144;
input v_145;
input v_146;
input v_147;
input v_148;
input v_276;
output o_1;
wire v_149;
wire v_150;
wire v_151;
wire v_152;
wire v_153;
wire v_154;
wire v_155;
wire v_156;
wire v_157;
wire v_158;
wire v_159;
wire v_160;
wire v_161;
wire v_162;
wire v_163;
wire v_164;
wire v_165;
wire v_166;
wire v_167;
wire v_168;
wire v_169;
wire v_170;
wire v_171;
wire v_172;
wire v_173;
wire v_174;
wire v_175;
wire v_176;
wire v_177;
wire v_178;
wire v_179;
wire v_180;
wire v_181;
wire v_182;
wire v_183;
wire v_184;
wire v_185;
wire v_186;
wire v_187;
wire v_188;
wire v_189;
wire v_190;
wire v_191;
wire v_192;
wire v_193;
wire v_194;
wire v_195;
wire v_196;
wire v_197;
wire v_198;
wire v_199;
wire v_200;
wire v_201;
wire v_202;
wire v_203;
wire v_204;
wire v_205;
wire v_206;
wire v_207;
wire v_208;
wire v_209;
wire v_210;
wire v_211;
wire v_212;
wire v_213;
wire v_214;
wire v_215;
wire v_216;
wire v_217;
wire v_218;
wire v_219;
wire v_220;
wire v_221;
wire v_222;
wire v_223;
wire v_224;
wire v_225;
wire v_226;
wire v_227;
wire v_228;
wire v_229;
wire v_230;
wire v_231;
wire v_232;
wire v_233;
wire v_234;
wire v_235;
wire v_236;
wire v_237;
wire v_238;
wire v_239;
wire v_240;
wire v_241;
wire v_242;
wire v_243;
wire v_244;
wire v_245;
wire v_246;
wire v_247;
wire v_248;
wire v_249;
wire v_250;
wire v_251;
wire v_252;
wire v_253;
wire v_254;
wire v_255;
wire v_256;
wire v_257;
wire v_258;
wire v_259;
wire v_260;
wire v_261;
wire v_262;
wire v_263;
wire v_264;
wire v_265;
wire v_266;
wire v_267;
wire v_268;
wire v_269;
wire v_270;
wire v_271;
wire v_272;
wire v_273;
wire v_274;
wire v_275;
wire v_277;
wire v_278;
wire v_279;
wire v_280;
wire v_281;
wire v_282;
wire v_283;
wire v_284;
wire v_285;
wire v_286;
wire v_287;
wire v_288;
wire v_289;
wire v_290;
wire v_291;
wire v_292;
wire v_293;
wire v_294;
wire v_295;
wire v_296;
wire v_297;
wire v_298;
wire v_299;
wire v_300;
wire v_301;
wire v_302;
wire v_303;
wire v_304;
wire v_305;
wire v_306;
wire v_307;
wire v_308;
wire v_309;
wire v_310;
wire v_311;
wire v_312;
wire v_313;
wire v_314;
wire v_315;
wire v_316;
wire v_317;
wire v_318;
wire v_319;
wire v_320;
wire v_321;
wire v_322;
wire v_323;
wire v_324;
wire v_325;
wire v_326;
wire v_327;
wire v_328;
wire v_329;
wire v_330;
wire v_331;
wire v_332;
wire v_333;
wire v_334;
wire v_335;
wire v_336;
wire v_337;
wire v_338;
wire v_339;
wire v_340;
wire v_341;
wire v_342;
wire v_343;
wire v_344;
wire v_345;
wire v_346;
wire v_347;
wire v_348;
wire v_349;
wire v_350;
wire v_351;
wire v_352;
wire v_353;
wire v_354;
wire v_355;
wire v_356;
wire v_357;
wire v_358;
wire v_359;
wire v_360;
wire v_361;
wire v_362;
wire v_363;
wire v_364;
wire v_365;
wire v_366;
wire v_367;
wire v_368;
wire v_369;
wire v_370;
wire v_371;
wire v_372;
wire v_373;
wire v_374;
wire v_375;
wire v_376;
wire v_377;
wire v_378;
wire v_379;
wire v_380;
wire v_381;
wire v_382;
wire v_383;
wire v_384;
wire v_385;
wire v_386;
wire v_387;
wire v_388;
wire v_389;
wire v_390;
wire v_391;
wire v_392;
wire v_393;
wire v_394;
wire v_395;
wire v_396;
wire v_397;
wire v_398;
wire v_399;
wire v_400;
wire v_401;
wire v_402;
wire v_403;
wire v_404;
wire v_405;
wire v_406;
wire v_407;
wire v_408;
wire v_409;
wire v_410;
wire v_411;
wire v_412;
wire v_413;
wire v_414;
wire v_415;
wire v_416;
wire v_417;
wire v_418;
wire v_419;
wire v_420;
wire v_421;
wire v_422;
wire v_423;
wire v_424;
wire v_425;
wire v_426;
wire v_427;
wire v_428;
wire v_429;
wire v_430;
wire v_431;
wire v_432;
wire v_433;
wire v_434;
wire v_435;
wire v_436;
wire v_437;
wire v_438;
wire v_439;
wire v_440;
wire v_441;
wire v_442;
wire v_443;
wire v_444;
wire v_445;
wire v_446;
wire v_447;
wire v_448;
wire v_449;
wire v_450;
wire v_451;
wire v_452;
wire v_453;
wire v_454;
wire v_455;
wire v_456;
wire v_457;
wire v_458;
wire v_459;
wire v_460;
wire v_461;
wire v_462;
wire v_463;
wire v_464;
wire v_465;
wire v_466;
wire v_467;
wire v_468;
wire v_469;
wire v_470;
wire v_471;
wire v_472;
wire v_473;
wire v_474;
wire v_475;
wire v_476;
wire v_477;
wire v_478;
wire v_479;
wire v_480;
wire v_481;
wire v_482;
wire v_483;
wire v_484;
wire v_485;
wire v_486;
wire v_487;
wire v_488;
wire v_489;
wire v_490;
wire v_491;
wire v_492;
wire v_493;
wire v_494;
wire v_495;
wire v_496;
wire v_497;
wire v_498;
wire v_499;
wire v_500;
wire v_501;
wire v_502;
wire v_503;
wire v_504;
wire v_505;
wire v_506;
wire v_507;
wire v_508;
wire v_509;
wire v_510;
wire v_511;
wire v_512;
wire v_513;
wire v_514;
wire v_515;
wire v_516;
wire v_517;
wire v_518;
wire v_519;
wire v_520;
wire v_521;
wire v_522;
wire v_523;
wire v_524;
wire v_525;
wire v_526;
wire v_527;
wire v_528;
wire v_529;
wire v_530;
wire v_531;
wire v_532;
wire v_533;
wire v_534;
wire v_535;
wire v_536;
wire v_537;
wire v_538;
wire v_539;
wire v_540;
wire v_541;
wire v_542;
wire v_543;
wire v_544;
wire v_545;
wire v_546;
wire v_547;
wire v_548;
wire v_549;
wire v_550;
wire v_551;
wire v_552;
wire v_553;
wire v_554;
wire v_555;
wire v_556;
wire v_557;
wire v_558;
wire v_559;
wire v_560;
wire v_561;
wire v_562;
wire v_563;
wire v_564;
wire v_565;
wire v_566;
wire v_567;
wire v_568;
wire v_569;
wire v_570;
wire v_571;
wire v_572;
wire v_573;
wire v_574;
wire v_575;
wire v_576;
wire v_577;
wire v_578;
wire v_579;
wire v_580;
wire v_581;
wire v_582;
wire v_583;
wire v_584;
wire v_585;
wire v_586;
wire v_587;
wire v_588;
wire v_589;
wire v_590;
wire v_591;
wire v_592;
wire v_593;
wire v_594;
wire v_595;
wire v_596;
wire v_597;
wire v_598;
wire v_599;
wire v_600;
wire v_601;
wire v_602;
wire v_603;
wire v_604;
wire v_605;
wire v_606;
wire v_607;
wire v_608;
wire v_609;
wire v_610;
wire v_611;
wire v_612;
wire v_613;
wire v_614;
wire v_615;
wire v_616;
wire v_617;
wire v_618;
wire v_619;
wire v_620;
wire v_621;
wire v_622;
wire v_623;
wire v_624;
wire v_625;
wire v_626;
wire v_627;
wire v_628;
wire v_629;
wire v_630;
wire v_631;
wire v_632;
wire v_633;
wire v_634;
wire v_635;
wire v_636;
wire v_637;
wire v_638;
wire v_639;
wire v_640;
wire v_641;
wire v_642;
wire v_643;
wire v_644;
wire v_645;
wire v_646;
wire v_647;
wire v_648;
wire v_649;
wire v_650;
wire v_651;
wire v_652;
wire v_653;
wire v_654;
wire v_655;
wire v_656;
wire v_657;
wire v_658;
wire v_659;
wire v_660;
wire v_661;
wire v_662;
wire v_663;
wire v_664;
wire v_665;
wire v_666;
wire v_667;
wire v_668;
wire v_669;
wire v_670;
wire v_671;
wire v_672;
wire v_673;
wire v_674;
wire v_675;
wire v_676;
wire v_677;
wire v_678;
wire v_679;
wire v_680;
wire v_681;
wire v_682;
wire v_683;
wire v_684;
wire v_685;
wire v_686;
wire v_687;
wire v_688;
wire v_689;
wire v_690;
wire v_691;
wire v_692;
wire v_693;
wire v_694;
wire v_695;
wire v_696;
wire v_697;
wire v_698;
wire v_699;
wire v_700;
wire v_701;
wire v_702;
wire v_703;
wire v_704;
wire v_705;
wire v_706;
wire v_707;
wire v_708;
wire v_709;
wire v_710;
wire v_711;
wire v_712;
wire v_713;
wire v_714;
wire v_715;
wire v_716;
wire v_717;
wire v_718;
wire v_719;
wire v_720;
wire v_721;
wire v_722;
wire v_723;
wire v_724;
wire v_725;
wire v_726;
wire v_727;
wire v_728;
wire v_729;
wire v_730;
wire v_731;
wire v_732;
wire v_733;
wire v_734;
wire v_735;
wire v_736;
wire v_737;
wire v_738;
wire v_739;
wire v_740;
wire v_741;
wire v_742;
wire v_743;
wire v_744;
wire v_745;
wire v_746;
wire v_747;
wire v_748;
wire v_749;
wire v_750;
wire v_751;
wire v_752;
wire v_753;
wire v_754;
wire v_755;
wire v_756;
wire v_757;
wire v_758;
wire v_759;
wire v_760;
wire v_761;
wire v_762;
wire v_763;
wire v_764;
wire v_765;
wire v_766;
wire v_767;
wire v_768;
wire v_769;
wire v_770;
wire v_771;
wire v_772;
wire v_773;
wire v_774;
wire v_775;
wire v_776;
wire v_777;
wire v_778;
wire v_779;
wire v_780;
wire v_781;
wire v_782;
wire v_783;
wire v_784;
wire v_785;
wire v_786;
wire v_787;
wire v_788;
wire v_789;
wire v_790;
wire v_791;
wire v_792;
wire v_793;
wire v_794;
wire v_795;
wire v_796;
wire v_797;
wire v_798;
wire v_799;
wire v_800;
wire v_801;
wire v_802;
wire v_803;
wire v_804;
wire v_805;
wire v_806;
wire v_807;
wire v_808;
wire v_809;
wire v_810;
wire v_811;
wire v_812;
wire v_813;
wire v_814;
wire v_815;
wire v_816;
wire v_817;
wire v_818;
wire v_819;
wire v_820;
wire v_821;
wire v_822;
wire v_823;
wire v_824;
wire v_825;
wire v_826;
wire v_827;
wire v_828;
wire v_829;
wire v_830;
wire v_831;
wire v_832;
wire v_833;
wire v_834;
wire v_835;
wire v_836;
wire v_837;
wire v_838;
wire v_839;
wire v_840;
wire v_841;
wire x_1;
wire x_2;
wire x_3;
assign v_640 = 0;
assign v_631 = 0;
assign v_629 = 0;
assign v_613 = 0;
assign v_279 = 0;
assign v_278 = 0;
assign v_234 = 0;
assign v_233 = 0;
assign v_232 = 0;
assign v_231 = 0;
assign v_230 = 0;
assign v_229 = 0;
assign v_228 = 0;
assign v_227 = 0;
assign v_226 = 0;
assign v_157 = 1;
assign v_277 = 1;
assign v_649 = 1;
assign v_149 = v_806 & v_807;
assign v_150 = v_808 & v_809;
assign v_151 = ~v_24 & ~v_25 & ~v_26 & ~v_27;
assign v_152 = ~v_31 & ~v_32 & ~v_33 & ~v_34;
assign v_153 = v_810 & v_811 & v_812 & v_813 & v_814;
assign v_154 = ~v_11 & v_1;
assign v_155 = ~v_11 & v_2;
assign v_158 = v_13;
assign v_159 = ~v_13 & v_156;
assign v_162 = v_161 & v_154;
assign v_164 = v_12 & v_163;
assign v_165 = ~v_12 & v_154;
assign v_169 = ~v_156 & v_58;
assign v_170 = v_156 & v_3;
assign v_172 = ~v_156 & v_59;
assign v_173 = v_156 & v_4;
assign v_175 = ~v_156 & v_60;
assign v_176 = v_156 & v_5;
assign v_178 = ~v_156 & v_61;
assign v_179 = v_156 & v_6;
assign v_181 = ~v_156 & v_62;
assign v_182 = v_156 & v_7;
assign v_184 = ~v_156 & v_63;
assign v_185 = v_156 & v_8;
assign v_187 = ~v_156 & v_64;
assign v_188 = v_156 & v_9;
assign v_190 = ~v_156 & v_65;
assign v_191 = v_156 & v_10;
assign v_193 = v_13 & v_171;
assign v_194 = ~v_13 & v_3;
assign v_196 = v_13 & v_174;
assign v_197 = ~v_13 & v_4;
assign v_199 = v_13 & v_177;
assign v_200 = ~v_13 & v_5;
assign v_202 = v_13 & v_180;
assign v_203 = ~v_13 & v_6;
assign v_205 = v_13 & v_183;
assign v_206 = ~v_13 & v_7;
assign v_208 = v_13 & v_186;
assign v_209 = ~v_13 & v_8;
assign v_211 = v_13 & v_189;
assign v_212 = ~v_13 & v_9;
assign v_214 = v_13 & v_192;
assign v_215 = ~v_13 & v_10;
assign v_225 = v_815 & v_816;
assign v_235 = ~v_14;
assign v_236 = ~v_15 & v_235;
assign v_237 = v_236;
assign v_238 = ~v_16 & v_237;
assign v_239 = v_238;
assign v_240 = ~v_17 & v_239;
assign v_242 = ~v_18 & v_241;
assign v_243 = v_242;
assign v_244 = ~v_19 & v_243;
assign v_246 = ~v_20 & v_245;
assign v_248 = ~v_21 & v_247;
assign v_249 = v_248;
assign v_250 = ~v_22 & v_249;
assign v_251 = v_250;
assign v_252 = ~v_23 & v_251;
assign v_253 = v_252;
assign v_254 = v_253;
assign v_255 = v_254;
assign v_256 = v_255;
assign v_257 = v_256;
assign v_258 = v_257;
assign v_259 = v_258;
assign v_260 = v_259;
assign v_261 = v_260;
assign v_262 = v_261;
assign v_263 = v_262;
assign v_264 = v_263;
assign v_265 = v_264;
assign v_266 = v_265;
assign v_267 = v_266;
assign v_268 = v_267;
assign v_269 = v_268;
assign v_270 = v_269;
assign v_271 = v_270;
assign v_272 = v_271;
assign v_273 = v_272;
assign v_274 = v_273;
assign v_275 = v_274;
assign v_280 = v_66;
assign v_281 = v_40 & v_12;
assign v_282 = ~v_40 & v_281;
assign v_284 = ~v_40 & v_12;
assign v_285 = v_40 & v_283;
assign v_288 = ~v_40 & v_13;
assign v_289 = ~v_46 & v_13;
assign v_291 = ~v_40 & v_290;
assign v_292 = v_40 & v_288;
assign v_295 = v_14;
assign v_297 = v_15 & v_295;
assign v_298 = v_297;
assign v_300 = v_16 & v_298;
assign v_301 = v_300;
assign v_303 = v_17 & v_301;
assign v_304 = v_303;
assign v_306 = v_18 & v_304;
assign v_307 = v_306;
assign v_309 = v_19 & v_307;
assign v_310 = v_309;
assign v_312 = v_20 & v_310;
assign v_313 = v_312;
assign v_315 = v_21 & v_313;
assign v_316 = v_315;
assign v_318 = v_22 & v_316;
assign v_319 = v_318;
assign v_321 = v_23 & v_319;
assign v_322 = v_321;
assign v_323 = ~v_14 & v_275;
assign v_324 = v_275 & v_296;
assign v_325 = v_275 & v_299;
assign v_326 = v_275 & v_302;
assign v_327 = v_275 & v_305;
assign v_328 = v_275 & v_308;
assign v_329 = v_275 & v_311;
assign v_330 = v_275 & v_314;
assign v_331 = v_275 & v_317;
assign v_332 = v_275 & v_320;
assign v_333 = v_1 & v_323;
assign v_334 = ~v_1 & v_14;
assign v_336 = v_1 & v_324;
assign v_337 = ~v_1 & v_15;
assign v_339 = v_1 & v_325;
assign v_340 = ~v_1 & v_16;
assign v_342 = v_1 & v_326;
assign v_343 = ~v_1 & v_17;
assign v_345 = v_1 & v_327;
assign v_346 = ~v_1 & v_18;
assign v_348 = v_1 & v_328;
assign v_349 = ~v_1 & v_19;
assign v_351 = v_1 & v_329;
assign v_352 = ~v_1 & v_20;
assign v_354 = v_1 & v_330;
assign v_355 = ~v_1 & v_21;
assign v_357 = v_1 & v_331;
assign v_358 = ~v_1 & v_22;
assign v_360 = v_1 & v_332;
assign v_361 = ~v_1 & v_23;
assign v_373 = v_817 & v_818;
assign v_374 = v_24;
assign v_376 = v_25 & v_374;
assign v_377 = v_376;
assign v_379 = v_26 & v_377;
assign v_380 = v_379;
assign v_382 = v_27 & v_380;
assign v_383 = v_382;
assign v_384 = ~v_375 & ~v_378 & v_24 & v_381;
assign v_385 = ~v_384 & ~v_24;
assign v_386 = ~v_384 & v_375;
assign v_387 = ~v_384 & v_378;
assign v_388 = ~v_384 & v_381;
assign v_389 = ~v_38 & v_385;
assign v_390 = v_38 & v_24;
assign v_392 = ~v_38 & v_386;
assign v_393 = v_38 & v_25;
assign v_395 = ~v_38 & v_387;
assign v_396 = v_38 & v_26;
assign v_398 = ~v_38 & v_388;
assign v_399 = v_38 & v_27;
assign v_401 = v_38 & v_24;
assign v_402 = ~v_38 & v_391;
assign v_404 = v_38 & v_25;
assign v_405 = ~v_38 & v_394;
assign v_407 = v_38 & v_26;
assign v_408 = ~v_38 & v_397;
assign v_410 = v_38 & v_27;
assign v_411 = ~v_38 & v_400;
assign v_413 = ~v_38 & v_24;
assign v_414 = v_38 & v_403;
assign v_416 = ~v_38 & v_25;
assign v_417 = v_38 & v_406;
assign v_419 = ~v_38 & v_26;
assign v_420 = v_38 & v_409;
assign v_422 = ~v_38 & v_27;
assign v_423 = v_38 & v_412;
assign v_425 = v_38 & v_24;
assign v_426 = ~v_38 & v_415;
assign v_428 = v_38 & v_25;
assign v_429 = ~v_38 & v_418;
assign v_431 = v_38 & v_26;
assign v_432 = ~v_38 & v_421;
assign v_434 = v_38 & v_27;
assign v_435 = ~v_38 & v_424;
assign v_437 = ~v_38 & v_24;
assign v_438 = v_38 & v_427;
assign v_440 = ~v_38 & v_25;
assign v_441 = v_38 & v_430;
assign v_443 = ~v_38 & v_26;
assign v_444 = v_38 & v_433;
assign v_446 = ~v_38 & v_27;
assign v_447 = v_38 & v_436;
assign v_453 = ~v_449 & ~v_450 & ~v_451 & ~v_452;
assign v_454 = v_38 & v_28;
assign v_455 = v_38 & v_28;
assign v_456 = ~v_38 & v_454;
assign v_458 = v_38 & v_457;
assign v_460 = v_38 & v_28;
assign v_461 = ~v_38 & v_459;
assign v_463 = ~v_38 & v_28;
assign v_464 = v_38 & v_462;
assign v_467 = v_38 & v_29;
assign v_468 = v_85 & v_29;
assign v_470 = v_38 & v_469;
assign v_471 = ~v_38 & v_467;
assign v_473 = ~v_38 & v_29;
assign v_474 = v_38 & v_472;
assign v_476 = v_38 & v_29;
assign v_477 = ~v_38 & v_475;
assign v_479 = ~v_38 & v_29;
assign v_480 = v_38 & v_478;
assign v_483 = v_42 & v_30;
assign v_485 = ~v_45 & v_30;
assign v_486 = v_45 & v_484;
assign v_488 = ~v_39 & v_487;
assign v_489 = v_39 & v_30;
assign v_491 = v_39 & v_30;
assign v_492 = ~v_39 & v_490;
assign v_494 = ~v_39 & v_30;
assign v_495 = v_39 & v_493;
assign v_498 = ~v_38 & v_385;
assign v_499 = v_38 & v_31;
assign v_501 = ~v_38 & v_386;
assign v_502 = v_38 & v_32;
assign v_504 = ~v_38 & v_387;
assign v_505 = v_38 & v_33;
assign v_507 = ~v_38 & v_388;
assign v_508 = v_38 & v_34;
assign v_510 = v_38 & v_31;
assign v_511 = ~v_38 & v_500;
assign v_513 = v_38 & v_32;
assign v_514 = ~v_38 & v_503;
assign v_516 = v_38 & v_33;
assign v_517 = ~v_38 & v_506;
assign v_519 = v_38 & v_34;
assign v_520 = ~v_38 & v_509;
assign v_522 = ~v_38 & v_31;
assign v_523 = v_38 & v_512;
assign v_525 = ~v_38 & v_32;
assign v_526 = v_38 & v_515;
assign v_528 = ~v_38 & v_33;
assign v_529 = v_38 & v_518;
assign v_531 = ~v_38 & v_34;
assign v_532 = v_38 & v_521;
assign v_534 = v_38 & v_31;
assign v_535 = ~v_38 & v_524;
assign v_537 = v_38 & v_32;
assign v_538 = ~v_38 & v_527;
assign v_540 = v_38 & v_33;
assign v_541 = ~v_38 & v_530;
assign v_543 = v_38 & v_34;
assign v_544 = ~v_38 & v_533;
assign v_546 = ~v_38 & v_31;
assign v_547 = v_38 & v_536;
assign v_549 = ~v_38 & v_32;
assign v_550 = v_38 & v_539;
assign v_552 = ~v_38 & v_33;
assign v_553 = v_38 & v_542;
assign v_555 = ~v_38 & v_34;
assign v_556 = v_38 & v_545;
assign v_562 = ~v_558 & ~v_559 & ~v_560 & ~v_561;
assign v_563 = v_85 & v_35;
assign v_564 = v_38 & v_563;
assign v_565 = ~v_38 & v_35;
assign v_567 = ~v_38 & v_35;
assign v_568 = v_38 & v_566;
assign v_570 = v_38 & v_35;
assign v_571 = ~v_38 & v_569;
assign v_573 = v_38 & v_572;
assign v_576 = v_13 & v_156;
assign v_577 = ~v_13 & v_36;
assign v_579 = v_12 & v_161;
assign v_580 = ~v_12 & v_578;
assign v_583 = ~v_41 & v_3;
assign v_585 = v_41 & v_4;
assign v_586 = ~v_41 & v_584;
assign v_588 = ~v_41 & v_5;
assign v_589 = v_41 & v_587;
assign v_591 = v_41 & v_6;
assign v_592 = ~v_41 & v_590;
assign v_594 = ~v_41 & v_7;
assign v_595 = v_41 & v_593;
assign v_597 = v_41 & v_8;
assign v_598 = ~v_41 & v_596;
assign v_600 = ~v_41 & v_9;
assign v_601 = v_41 & v_599;
assign v_603 = v_41 & v_10;
assign v_604 = ~v_41 & v_602;
assign v_606 = ~v_41 & v_605;
assign v_607 = ~v_275 & v_606;
assign v_609 = v_1 & v_608;
assign v_612 = ~v_43 & v_38;
assign v_614 = v_612;
assign v_615 = v_38 & v_614;
assign v_617 = ~v_38 & v_616;
assign v_618 = v_38 & v_617;
assign v_620 = v_38 & v_85;
assign v_621 = ~v_38 & v_619;
assign v_623 = v_38 & v_622;
assign v_625 = ~v_38 & v_624;
assign v_626 = v_38 & v_625;
assign v_630 = ~v_39 & v_45;
assign v_632 = v_630;
assign v_633 = ~v_39 & v_632;
assign v_634 = ~v_39 & v_44;
assign v_635 = v_39 & v_633;
assign v_638 = ~v_11 & v_40;
assign v_639 = v_40 & v_638;
assign v_641 = v_639;
assign v_642 = v_40 & v_641;
assign v_644 = ~v_40 & v_643;
assign v_645 = ~v_40 & v_46;
assign v_646 = v_40 & v_644;
assign v_650 = v_41;
assign v_651 = ~v_41 & v_650;
assign v_652 = v_41 & v_651;
assign v_654 = ~v_41 & v_653;
assign v_655 = v_41 & v_654;
assign v_657 = ~v_41 & v_656;
assign v_658 = v_41 & v_657;
assign v_660 = ~v_41 & v_659;
assign v_661 = ~v_41 & v_660;
assign v_663 = ~v_275 & v_662;
assign v_664 = v_275 & v_41;
assign v_666 = v_1 & v_665;
assign v_667 = ~v_1 & v_41;
assign v_670 = ~v_45 & v_42;
assign v_671 = ~v_42 & v_45;
assign v_673 = ~v_39 & v_672;
assign v_674 = v_39 & v_42;
assign v_676 = v_39 & v_42;
assign v_677 = ~v_39 & v_675;
assign v_679 = ~v_39 & v_42;
assign v_680 = v_39 & v_678;
assign v_683 = ~v_42 & v_43;
assign v_684 = ~v_45 & v_43;
assign v_685 = v_45 & v_683;
assign v_687 = ~v_39 & v_686;
assign v_688 = v_39 & v_43;
assign v_690 = v_39 & v_43;
assign v_691 = ~v_39 & v_689;
assign v_693 = ~v_44 & v_43;
assign v_695 = ~v_39 & v_694;
assign v_696 = v_39 & v_692;
assign v_699 = ~v_43 & v_44;
assign v_700 = v_38 & v_699;
assign v_701 = ~v_38 & v_44;
assign v_703 = ~v_38 & v_44;
assign v_704 = v_38 & v_702;
assign v_706 = ~v_38 & v_705;
assign v_708 = ~v_38 & v_44;
assign v_709 = v_38 & v_707;
assign v_711 = v_38 & v_44;
assign v_712 = ~v_38 & v_710;
assign v_714 = ~v_38 & v_44;
assign v_715 = v_38 & v_713;
assign v_717 = v_38 & v_44;
assign v_718 = ~v_38 & v_716;
assign v_720 = ~v_38 & v_44;
assign v_721 = v_38 & v_719;
assign v_724 = ~v_11 & v_45;
assign v_726 = v_40 & v_725;
assign v_727 = ~v_40 & v_45;
assign v_729 = ~v_40 & v_45;
assign v_730 = v_40 & v_728;
assign v_732 = v_40 & v_45;
assign v_733 = ~v_40 & v_731;
assign v_735 = v_40 & v_734;
assign v_737 = v_45 & v_46;
assign v_738 = ~v_39 & v_737;
assign v_739 = v_39 & v_46;
assign v_741 = ~v_39 & v_740;
assign v_743 = ~v_39 & v_46;
assign v_744 = v_39 & v_742;
assign v_747 = v_819 & v_820 & v_821 & v_822 & v_823;
assign v_748 = v_153 & v_747;
assign v_749 = v_824 & v_825;
assign v_750 = v_826 & v_827;
assign v_751 = ~v_126 & ~v_127 & ~v_128 & ~v_129;
assign v_752 = ~v_133 & ~v_134 & ~v_135 & ~v_136;
assign v_753 = v_828 & v_829 & v_830 & v_831 & v_832;
assign v_764 = v_833 & v_834;
assign v_778 = v_835 & v_836;
assign v_783 = ~v_779 & ~v_780 & ~v_781 & ~v_782;
assign v_791 = ~v_787 & ~v_788 & ~v_789 & ~v_790;
assign v_804 = v_837 & v_838 & v_839 & v_840 & v_841;
assign v_805 = v_753 & v_804;
assign v_806 = ~v_3 & ~v_4 & ~v_5 & ~v_6 & ~v_7;
assign v_807 = ~v_8 & ~v_9 & ~v_10;
assign v_808 = ~v_14 & ~v_15 & ~v_16 & ~v_17 & ~v_18;
assign v_809 = ~v_19 & ~v_20 & ~v_21 & ~v_22 & ~v_23;
assign v_810 = ~v_1 & ~v_2 & ~v_11 & ~v_12 & ~v_13;
assign v_811 = ~v_28 & ~v_29 & ~v_30 & ~v_35 & ~v_36;
assign v_812 = ~v_37 & ~v_38 & ~v_39 & ~v_40 & ~v_42;
assign v_813 = ~v_43 & ~v_44 & ~v_45 & ~v_46 & v_149;
assign v_814 = v_150 & v_151 & v_152 & v_41;
assign v_815 = ~v_217 & ~v_218 & ~v_219 & ~v_220 & ~v_221;
assign v_816 = ~v_222 & ~v_223 & ~v_224;
assign v_817 = ~v_363 & ~v_364 & ~v_365 & ~v_366 & ~v_367;
assign v_818 = ~v_368 & ~v_369 & ~v_370 & ~v_371 & ~v_372;
assign v_819 = ~v_167 & ~v_168 & ~v_280 & ~v_287 & ~v_294;
assign v_820 = ~v_466 & ~v_482 & ~v_497 & ~v_575 & ~v_582;
assign v_821 = ~v_611 & ~v_628 & ~v_637 & ~v_648 & ~v_669;
assign v_822 = ~v_682 & ~v_698 & ~v_723 & ~v_736 & ~v_746;
assign v_823 = v_225 & v_373 & v_453 & v_562;
assign v_824 = ~v_105 & ~v_106 & ~v_107 & ~v_108 & ~v_109;
assign v_825 = ~v_110 & ~v_111 & ~v_112;
assign v_826 = ~v_116 & ~v_117 & ~v_118 & ~v_119 & ~v_120;
assign v_827 = ~v_121 & ~v_122 & ~v_123 & ~v_124 & ~v_125;
assign v_828 = ~v_103 & ~v_104 & ~v_113 & ~v_114 & ~v_115;
assign v_829 = ~v_130 & ~v_131 & ~v_132 & ~v_137 & ~v_138;
assign v_830 = ~v_139 & ~v_140 & ~v_141 & ~v_142 & ~v_144;
assign v_831 = ~v_145 & ~v_146 & ~v_147 & ~v_148 & v_749;
assign v_832 = v_750 & v_751 & v_752 & v_143;
assign v_833 = ~v_756 & ~v_757 & ~v_758 & ~v_759 & ~v_760;
assign v_834 = ~v_761 & ~v_762 & ~v_763;
assign v_835 = ~v_768 & ~v_769 & ~v_770 & ~v_771 & ~v_772;
assign v_836 = ~v_773 & ~v_774 & ~v_775 & ~v_776 & ~v_777;
assign v_837 = ~v_754 & ~v_755 & ~v_765 & ~v_766 & ~v_767;
assign v_838 = ~v_784 & ~v_785 & ~v_786 & ~v_792 & ~v_793;
assign v_839 = ~v_794 & ~v_795 & ~v_796 & ~v_797 & ~v_798;
assign v_840 = ~v_799 & ~v_800 & ~v_801 & ~v_802 & ~v_803;
assign v_841 = v_764 & v_778 & v_783 & v_791;
assign v_156 = v_11 | v_155;
assign v_160 = v_158 | v_159;
assign v_161 = ~v_160 | ~v_48;
assign v_163 = v_162 | ~v_161;
assign v_166 = v_164 | v_165;
assign v_171 = v_169 | v_170;
assign v_174 = v_172 | v_173;
assign v_177 = v_175 | v_176;
assign v_180 = v_178 | v_179;
assign v_183 = v_181 | v_182;
assign v_186 = v_184 | v_185;
assign v_189 = v_187 | v_188;
assign v_192 = v_190 | v_191;
assign v_195 = v_193 | v_194;
assign v_198 = v_196 | v_197;
assign v_201 = v_199 | v_200;
assign v_204 = v_202 | v_203;
assign v_207 = v_205 | v_206;
assign v_210 = v_208 | v_209;
assign v_213 = v_211 | v_212;
assign v_216 = v_214 | v_215;
assign v_241 = v_239 | v_240 | ~v_17;
assign v_245 = v_243 | v_244 | ~v_19;
assign v_247 = v_245 | v_246 | ~v_20;
assign v_283 = v_40 | v_282;
assign v_286 = v_284 | v_285;
assign v_290 = v_46 | v_289;
assign v_293 = v_291 | v_292;
assign v_335 = v_333 | v_334;
assign v_338 = v_336 | v_337;
assign v_341 = v_339 | v_340;
assign v_344 = v_342 | v_343;
assign v_347 = v_345 | v_346;
assign v_350 = v_348 | v_349;
assign v_353 = v_351 | v_352;
assign v_356 = v_354 | v_355;
assign v_359 = v_357 | v_358;
assign v_362 = v_360 | v_361;
assign v_391 = v_389 | v_390;
assign v_394 = v_392 | v_393;
assign v_397 = v_395 | v_396;
assign v_400 = v_398 | v_399;
assign v_403 = v_401 | v_402;
assign v_406 = v_404 | v_405;
assign v_409 = v_407 | v_408;
assign v_412 = v_410 | v_411;
assign v_415 = v_413 | v_414;
assign v_418 = v_416 | v_417;
assign v_421 = v_419 | v_420;
assign v_424 = v_422 | v_423;
assign v_427 = v_425 | v_426;
assign v_430 = v_428 | v_429;
assign v_433 = v_431 | v_432;
assign v_436 = v_434 | v_435;
assign v_439 = v_437 | v_438;
assign v_442 = v_440 | v_441;
assign v_445 = v_443 | v_444;
assign v_448 = v_446 | v_447;
assign v_457 = v_455 | v_456;
assign v_459 = v_458 | ~v_38;
assign v_462 = v_460 | v_461;
assign v_465 = v_463 | v_464;
assign v_469 = v_468 | ~v_85;
assign v_472 = v_470 | v_471;
assign v_475 = v_473 | v_474;
assign v_478 = v_476 | v_477;
assign v_481 = v_479 | v_480;
assign v_484 = v_483 | ~v_42;
assign v_487 = v_485 | v_486;
assign v_490 = v_488 | v_489;
assign v_493 = v_491 | v_492;
assign v_496 = v_494 | v_495;
assign v_500 = v_498 | v_499;
assign v_503 = v_501 | v_502;
assign v_506 = v_504 | v_505;
assign v_509 = v_507 | v_508;
assign v_512 = v_510 | v_511;
assign v_515 = v_513 | v_514;
assign v_518 = v_516 | v_517;
assign v_521 = v_519 | v_520;
assign v_524 = v_522 | v_523;
assign v_527 = v_525 | v_526;
assign v_530 = v_528 | v_529;
assign v_533 = v_531 | v_532;
assign v_536 = v_534 | v_535;
assign v_539 = v_537 | v_538;
assign v_542 = v_540 | v_541;
assign v_545 = v_543 | v_544;
assign v_548 = v_546 | v_547;
assign v_551 = v_549 | v_550;
assign v_554 = v_552 | v_553;
assign v_557 = v_555 | v_556;
assign v_566 = v_564 | v_565;
assign v_569 = v_567 | v_568;
assign v_572 = v_570 | v_571;
assign v_574 = v_573 | ~v_38;
assign v_578 = v_576 | v_577;
assign v_581 = v_579 | v_580;
assign v_584 = v_583 | v_41;
assign v_587 = v_585 | v_586;
assign v_590 = v_588 | v_589;
assign v_593 = v_591 | v_592;
assign v_596 = v_594 | v_595;
assign v_599 = v_597 | v_598;
assign v_602 = v_600 | v_601;
assign v_605 = v_603 | v_604;
assign v_608 = v_607 | v_275;
assign v_610 = v_609 | ~v_1;
assign v_616 = v_615 | ~v_38;
assign v_619 = v_618 | ~v_38;
assign v_622 = v_620 | v_621;
assign v_624 = v_623 | ~v_38;
assign v_627 = v_626 | ~v_38;
assign v_636 = v_634 | v_635;
assign v_643 = v_642 | ~v_40;
assign v_647 = v_645 | v_646;
assign v_653 = v_652 | ~v_41;
assign v_656 = v_655 | ~v_41;
assign v_659 = v_658 | ~v_41;
assign v_662 = v_41 | v_661;
assign v_665 = v_663 | v_664;
assign v_668 = v_666 | v_667;
assign v_672 = v_670 | v_671;
assign v_675 = v_673 | v_674;
assign v_678 = v_676 | v_677;
assign v_681 = v_679 | v_680;
assign v_686 = v_684 | v_685;
assign v_689 = v_687 | v_688;
assign v_692 = v_690 | v_691;
assign v_694 = v_44 | v_693;
assign v_697 = v_695 | v_696;
assign v_702 = v_700 | v_701;
assign v_705 = v_703 | v_704;
assign v_707 = v_38 | v_706;
assign v_710 = v_708 | v_709;
assign v_713 = v_711 | v_712;
assign v_716 = v_714 | v_715;
assign v_719 = v_717 | v_718;
assign v_722 = v_720 | v_721;
assign v_725 = v_11 | v_724;
assign v_728 = v_726 | v_727;
assign v_731 = v_729 | v_730;
assign v_734 = v_732 | v_733;
assign v_740 = v_738 | v_739;
assign v_742 = v_39 | v_741;
assign v_745 = v_743 | v_744;
assign v_167 = v_166 ^ v_47;
assign v_168 = v_160 ^ v_49;
assign v_217 = v_195 ^ v_50;
assign v_218 = v_198 ^ v_51;
assign v_219 = v_201 ^ v_52;
assign v_220 = v_204 ^ v_53;
assign v_221 = v_207 ^ v_54;
assign v_222 = v_210 ^ v_55;
assign v_223 = v_213 ^ v_56;
assign v_224 = v_216 ^ v_57;
assign v_287 = v_286 ^ v_67;
assign v_294 = v_293 ^ v_68;
assign v_296 = v_295 ^ v_15;
assign v_299 = v_298 ^ v_16;
assign v_302 = v_301 ^ v_17;
assign v_305 = v_304 ^ v_18;
assign v_308 = v_307 ^ v_19;
assign v_311 = v_310 ^ v_20;
assign v_314 = v_313 ^ v_21;
assign v_317 = v_316 ^ v_22;
assign v_320 = v_319 ^ v_23;
assign v_363 = v_335 ^ v_69;
assign v_364 = v_338 ^ v_70;
assign v_365 = v_341 ^ v_71;
assign v_366 = v_344 ^ v_72;
assign v_367 = v_347 ^ v_73;
assign v_368 = v_350 ^ v_74;
assign v_369 = v_353 ^ v_75;
assign v_370 = v_356 ^ v_76;
assign v_371 = v_359 ^ v_77;
assign v_372 = v_362 ^ v_78;
assign v_375 = v_374 ^ v_25;
assign v_378 = v_377 ^ v_26;
assign v_381 = v_380 ^ v_27;
assign v_449 = v_439 ^ v_79;
assign v_450 = v_442 ^ v_80;
assign v_451 = v_445 ^ v_81;
assign v_452 = v_448 ^ v_82;
assign v_466 = v_465 ^ v_83;
assign v_482 = v_481 ^ v_84;
assign v_497 = v_496 ^ v_86;
assign v_558 = v_548 ^ v_87;
assign v_559 = v_551 ^ v_88;
assign v_560 = v_554 ^ v_89;
assign v_561 = v_557 ^ v_90;
assign v_575 = v_574 ^ v_91;
assign v_582 = v_581 ^ v_92;
assign v_611 = v_610 ^ v_93;
assign v_628 = v_627 ^ v_94;
assign v_637 = v_636 ^ v_95;
assign v_648 = v_647 ^ v_96;
assign v_669 = v_668 ^ v_97;
assign v_682 = v_681 ^ v_98;
assign v_698 = v_697 ^ v_99;
assign v_723 = v_722 ^ v_100;
assign v_736 = v_735 ^ v_101;
assign v_746 = v_745 ^ v_102;
assign v_754 = v_103 ^ v_47;
assign v_755 = v_104 ^ v_49;
assign v_756 = v_105 ^ v_50;
assign v_757 = v_106 ^ v_51;
assign v_758 = v_107 ^ v_52;
assign v_759 = v_108 ^ v_53;
assign v_760 = v_109 ^ v_54;
assign v_761 = v_110 ^ v_55;
assign v_762 = v_111 ^ v_56;
assign v_763 = v_112 ^ v_57;
assign v_765 = v_113 ^ v_66;
assign v_766 = v_114 ^ v_67;
assign v_767 = v_115 ^ v_68;
assign v_768 = v_116 ^ v_69;
assign v_769 = v_117 ^ v_70;
assign v_770 = v_118 ^ v_71;
assign v_771 = v_119 ^ v_72;
assign v_772 = v_120 ^ v_73;
assign v_773 = v_121 ^ v_74;
assign v_774 = v_122 ^ v_75;
assign v_775 = v_123 ^ v_76;
assign v_776 = v_124 ^ v_77;
assign v_777 = v_125 ^ v_78;
assign v_779 = v_126 ^ v_79;
assign v_780 = v_127 ^ v_80;
assign v_781 = v_128 ^ v_81;
assign v_782 = v_129 ^ v_82;
assign v_784 = v_130 ^ v_83;
assign v_785 = v_131 ^ v_84;
assign v_786 = v_132 ^ v_86;
assign v_787 = v_133 ^ v_87;
assign v_788 = v_134 ^ v_88;
assign v_789 = v_135 ^ v_89;
assign v_790 = v_136 ^ v_90;
assign v_792 = v_137 ^ v_91;
assign v_793 = v_138 ^ v_92;
assign v_794 = v_139 ^ v_93;
assign v_795 = v_140 ^ v_94;
assign v_796 = v_141 ^ v_95;
assign v_797 = v_142 ^ v_96;
assign v_798 = v_143 ^ v_97;
assign v_799 = v_144 ^ v_98;
assign v_800 = v_145 ^ v_99;
assign v_801 = v_146 ^ v_100;
assign v_802 = v_147 ^ v_101;
assign v_803 = v_148 ^ v_102;
assign x_1 = v_275 | ~v_276;
assign x_2 = v_805 | ~v_748;
assign x_3 = x_1 & x_2;
assign o_1 = x_3;
endmodule
