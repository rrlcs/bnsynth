// skolem function for order file variables
// Generated using findDep.cpp 
module kenflashp04 (v_279, v_280, v_281, v_282, v_283, v_284, v_285, v_286, v_287, v_288, v_289, v_290, v_291, v_292, v_293, v_294, v_295, v_296, v_297, v_298, v_299, v_300, v_301, v_302, v_303, v_304, v_305, v_306, v_307, v_308, v_309, v_310, v_311, v_312, v_313, v_314, v_315, v_316, v_317, v_318, v_319, v_320, v_321, v_322, v_323, v_324, v_325, v_326, v_327, v_328, v_329, v_330, v_331, v_332, v_333, v_334, v_335, v_336, v_337, v_338, v_339, v_340, v_341, v_342, v_343, v_216, v_217, v_218, v_219, v_220, v_221, v_222, v_223, v_224, v_225, v_226, v_227, v_228, v_229, v_230, v_231, v_232, v_233, v_234, v_235, v_236, v_237, v_238, v_239, v_240, v_241, v_242, v_243, v_244, v_245, v_246, v_247, v_248, v_249, v_250, v_251, v_252, v_253, v_254, v_255, v_256, v_257, v_258, v_259, v_260, v_261, v_262, v_263, v_264, v_265, v_266, v_267, v_268, v_269, v_270, v_271, v_272, v_273, v_274, v_275, v_276, v_277, v_278, v_5, v_6, v_8, v_10, v_11, v_14, v_16, v_18, v_20, v_25, v_29, v_32, v_33, v_34, v_35, v_37, v_39, v_42, v_44, v_45, v_46, v_48, v_49, v_51, v_53, v_54, v_56, v_59, v_65, v_67, v_68, v_69, v_70, v_71, v_72, v_77, v_79, v_80, v_81, v_82, v_84, v_87, v_89, v_90, v_96, v_98, v_99, v_100, v_101, v_102, v_103, v_104, v_107, v_108, v_113, v_115, v_116, v_118, v_119, v_120, v_123, v_126, v_131, v_132, v_135, v_138, v_139, v_140, v_143, v_144, v_145, v_146, v_148, v_154, v_156, v_166, v_169, v_170, v_173, v_177, v_179, v_181, v_184, v_187, v_191, v_192, v_193, v_198, v_199, v_200, v_202, v_207, v_208, v_210, v_211, v_212, v_213, o_1);
input v_279;
input v_280;
input v_281;
input v_282;
input v_283;
input v_284;
input v_285;
input v_286;
input v_287;
input v_288;
input v_289;
input v_290;
input v_291;
input v_292;
input v_293;
input v_294;
input v_295;
input v_296;
input v_297;
input v_298;
input v_299;
input v_300;
input v_301;
input v_302;
input v_303;
input v_304;
input v_305;
input v_306;
input v_307;
input v_308;
input v_309;
input v_310;
input v_311;
input v_312;
input v_313;
input v_314;
input v_315;
input v_316;
input v_317;
input v_318;
input v_319;
input v_320;
input v_321;
input v_322;
input v_323;
input v_324;
input v_325;
input v_326;
input v_327;
input v_328;
input v_329;
input v_330;
input v_331;
input v_332;
input v_333;
input v_334;
input v_335;
input v_336;
input v_337;
input v_338;
input v_339;
input v_340;
input v_341;
input v_342;
input v_343;
input v_216;
input v_217;
input v_218;
input v_219;
input v_220;
input v_221;
input v_222;
input v_223;
input v_224;
input v_225;
input v_226;
input v_227;
input v_228;
input v_229;
input v_230;
input v_231;
input v_232;
input v_233;
input v_234;
input v_235;
input v_236;
input v_237;
input v_238;
input v_239;
input v_240;
input v_241;
input v_242;
input v_243;
input v_244;
input v_245;
input v_246;
input v_247;
input v_248;
input v_249;
input v_250;
input v_251;
input v_252;
input v_253;
input v_254;
input v_255;
input v_256;
input v_257;
input v_258;
input v_259;
input v_260;
input v_261;
input v_262;
input v_263;
input v_264;
input v_265;
input v_266;
input v_267;
input v_268;
input v_269;
input v_270;
input v_271;
input v_272;
input v_273;
input v_274;
input v_275;
input v_276;
input v_277;
input v_278;
input v_5;
input v_6;
input v_8;
input v_10;
input v_11;
input v_14;
input v_16;
input v_18;
input v_20;
input v_25;
input v_29;
input v_32;
input v_33;
input v_34;
input v_35;
input v_37;
input v_39;
input v_42;
input v_44;
input v_45;
input v_46;
input v_48;
input v_49;
input v_51;
input v_53;
input v_54;
input v_56;
input v_59;
input v_65;
input v_67;
input v_68;
input v_69;
input v_70;
input v_71;
input v_72;
input v_77;
input v_79;
input v_80;
input v_81;
input v_82;
input v_84;
input v_87;
input v_89;
input v_90;
input v_96;
input v_98;
input v_99;
input v_100;
input v_101;
input v_102;
input v_103;
input v_104;
input v_107;
input v_108;
input v_113;
input v_115;
input v_116;
input v_118;
input v_119;
input v_120;
input v_123;
input v_126;
input v_131;
input v_132;
input v_135;
input v_138;
input v_139;
input v_140;
input v_143;
input v_144;
input v_145;
input v_146;
input v_148;
input v_154;
input v_156;
input v_166;
input v_169;
input v_170;
input v_173;
input v_177;
input v_179;
input v_181;
input v_184;
input v_187;
input v_191;
input v_192;
input v_193;
input v_198;
input v_199;
input v_200;
input v_202;
input v_207;
input v_208;
input v_210;
input v_211;
input v_212;
input v_213;
output o_1;
wire v_2;
wire v_3;
wire v_4;
wire v_7;
wire v_9;
wire v_12;
wire v_13;
wire v_15;
wire v_17;
wire v_19;
wire v_21;
wire v_22;
wire v_23;
wire v_24;
wire v_26;
wire v_27;
wire v_28;
wire v_30;
wire v_31;
wire v_36;
wire v_38;
wire v_40;
wire v_41;
wire v_43;
wire v_47;
wire v_50;
wire v_52;
wire v_55;
wire v_57;
wire v_58;
wire v_60;
wire v_61;
wire v_62;
wire v_63;
wire v_64;
wire v_66;
wire v_73;
wire v_74;
wire v_75;
wire v_76;
wire v_78;
wire v_83;
wire v_85;
wire v_86;
wire v_88;
wire v_91;
wire v_92;
wire v_93;
wire v_94;
wire v_95;
wire v_97;
wire v_105;
wire v_106;
wire v_109;
wire v_110;
wire v_111;
wire v_112;
wire v_114;
wire v_117;
wire v_121;
wire v_122;
wire v_124;
wire v_125;
wire v_127;
wire v_128;
wire v_129;
wire v_130;
wire v_133;
wire v_134;
wire v_136;
wire v_137;
wire v_141;
wire v_142;
wire v_147;
wire v_149;
wire v_150;
wire v_151;
wire v_152;
wire v_153;
wire v_155;
wire v_157;
wire v_158;
wire v_159;
wire v_160;
wire v_161;
wire v_162;
wire v_163;
wire v_164;
wire v_165;
wire v_167;
wire v_168;
wire v_171;
wire v_172;
wire v_174;
wire v_175;
wire v_176;
wire v_178;
wire v_180;
wire v_182;
wire v_183;
wire v_185;
wire v_186;
wire v_188;
wire v_189;
wire v_190;
wire v_194;
wire v_195;
wire v_196;
wire v_197;
wire v_201;
wire v_203;
wire v_204;
wire v_205;
wire v_206;
wire v_209;
wire v_214;
wire v_215;
wire v_409;
wire x_1;
wire x_2;
wire x_3;
wire x_4;
wire x_5;
wire x_6;
wire x_7;
wire x_8;
wire x_9;
wire x_10;
wire x_11;
wire x_12;
wire x_13;
wire x_14;
wire x_15;
wire x_16;
wire x_17;
wire x_18;
wire x_19;
wire x_20;
wire x_21;
wire x_22;
wire x_23;
wire x_24;
wire x_25;
wire x_26;
wire x_27;
wire x_28;
wire x_29;
wire x_30;
wire x_31;
wire x_32;
wire x_33;
wire x_34;
wire x_35;
wire x_36;
wire x_37;
wire x_38;
wire x_39;
wire x_40;
wire x_41;
wire x_42;
wire x_43;
wire x_44;
wire x_45;
wire x_46;
wire x_47;
wire x_48;
wire x_49;
wire x_50;
wire x_51;
wire x_52;
wire x_53;
wire x_54;
wire x_55;
wire x_56;
wire x_57;
wire x_58;
wire x_59;
wire x_60;
wire x_61;
wire x_62;
wire x_63;
wire x_64;
wire x_65;
wire x_66;
wire x_67;
wire x_68;
wire x_69;
wire x_70;
wire x_71;
wire x_72;
wire x_73;
wire x_74;
wire x_75;
wire x_76;
wire x_77;
wire x_78;
wire x_79;
wire x_80;
wire x_81;
wire x_82;
wire x_83;
wire x_84;
wire x_85;
wire x_86;
wire x_87;
wire x_88;
wire x_89;
wire x_90;
wire x_91;
wire x_92;
wire x_93;
wire x_94;
wire x_95;
wire x_96;
wire x_97;
wire x_98;
wire x_99;
wire x_100;
wire x_101;
wire x_102;
wire x_103;
wire x_104;
wire x_105;
wire x_106;
wire x_107;
wire x_108;
wire x_109;
wire x_110;
wire x_111;
wire x_112;
wire x_113;
wire x_114;
wire x_115;
wire x_116;
wire x_117;
wire x_118;
wire x_119;
wire x_120;
wire x_121;
wire x_122;
wire x_123;
wire x_124;
wire x_125;
wire x_126;
wire x_127;
wire x_128;
wire x_129;
wire x_130;
wire x_131;
wire x_132;
wire x_133;
wire x_134;
wire x_135;
wire x_136;
wire x_137;
wire x_138;
wire x_139;
wire x_140;
wire x_141;
wire x_142;
wire x_143;
wire x_144;
wire x_145;
wire x_146;
wire x_147;
wire x_148;
wire x_149;
wire x_150;
wire x_151;
wire x_152;
wire x_153;
wire x_154;
wire x_155;
wire x_156;
wire x_157;
wire x_158;
wire x_159;
wire x_160;
wire x_161;
wire x_162;
wire x_163;
wire x_164;
wire x_165;
wire x_166;
wire x_167;
wire x_168;
wire x_169;
wire x_170;
wire x_171;
wire x_172;
wire x_173;
wire x_174;
wire x_175;
wire x_176;
wire x_177;
wire x_178;
wire x_179;
wire x_180;
wire x_181;
wire x_182;
wire x_183;
wire x_184;
wire x_185;
wire x_186;
wire x_187;
wire x_188;
wire x_189;
wire x_190;
wire x_191;
wire x_192;
wire x_193;
wire x_194;
wire x_195;
wire x_196;
wire x_197;
wire x_198;
wire x_199;
wire x_200;
wire x_201;
wire x_202;
wire x_203;
wire x_204;
wire x_205;
wire x_206;
wire x_207;
wire x_208;
wire x_209;
wire x_210;
wire x_211;
wire x_212;
wire x_213;
wire x_214;
wire x_215;
wire x_216;
wire x_217;
wire x_218;
wire x_219;
wire x_220;
wire x_221;
wire x_222;
wire x_223;
wire x_224;
wire x_225;
wire x_226;
wire x_227;
wire x_228;
wire x_229;
wire x_230;
wire x_231;
wire x_232;
wire x_233;
wire x_234;
wire x_235;
wire x_236;
wire x_237;
wire x_238;
wire x_239;
wire x_240;
wire x_241;
wire x_242;
wire x_243;
wire x_244;
wire x_245;
wire x_246;
wire x_247;
wire x_248;
wire x_249;
wire x_250;
wire x_251;
wire x_252;
wire x_253;
wire x_254;
wire x_255;
wire x_256;
wire x_257;
wire x_258;
wire x_259;
wire x_260;
wire x_261;
wire x_262;
wire x_263;
wire x_264;
wire x_265;
wire x_266;
wire x_267;
wire x_268;
wire x_269;
wire x_270;
wire x_271;
wire x_272;
wire x_273;
wire x_274;
wire x_275;
wire x_276;
wire x_277;
wire x_278;
wire x_279;
wire x_280;
wire x_281;
wire x_282;
wire x_283;
wire x_284;
wire x_285;
wire x_286;
wire x_287;
wire x_288;
wire x_289;
wire x_290;
wire x_291;
wire x_292;
wire x_293;
wire x_294;
wire x_295;
wire x_296;
wire x_297;
wire x_298;
wire x_299;
wire x_300;
wire x_301;
wire x_302;
wire x_303;
wire x_304;
wire x_305;
wire x_306;
wire x_307;
wire x_308;
wire x_309;
wire x_310;
wire x_311;
wire x_312;
wire x_313;
wire x_314;
wire x_315;
wire x_316;
wire x_317;
wire x_318;
wire x_319;
wire x_320;
wire x_321;
wire x_322;
wire x_323;
wire x_324;
wire x_325;
wire x_326;
wire x_327;
wire x_328;
wire x_329;
wire x_330;
wire x_331;
wire x_332;
wire x_333;
wire x_334;
wire x_335;
wire x_336;
wire x_337;
wire x_338;
wire x_339;
wire x_340;
wire x_341;
wire x_342;
wire x_343;
wire x_344;
wire x_345;
wire x_346;
wire x_347;
wire x_348;
wire x_349;
wire x_350;
wire x_351;
wire x_352;
wire x_353;
wire x_354;
wire x_355;
wire x_356;
wire x_357;
wire x_358;
wire x_359;
wire x_360;
wire x_361;
wire x_362;
wire x_363;
wire x_364;
wire x_365;
wire x_366;
wire x_367;
wire x_368;
wire x_369;
wire x_370;
wire x_371;
wire x_372;
wire x_373;
wire x_374;
wire x_375;
wire x_376;
wire x_377;
wire x_378;
wire x_379;
wire x_380;
wire x_381;
wire x_382;
wire x_383;
wire x_384;
wire x_385;
wire x_386;
wire x_387;
wire x_388;
wire x_389;
wire x_390;
wire x_391;
wire x_392;
wire x_393;
wire x_394;
wire x_395;
wire x_396;
wire x_397;
wire x_398;
wire x_399;
wire x_400;
wire x_401;
wire x_402;
wire x_403;
wire x_404;
wire x_405;
wire x_406;
wire x_407;
wire x_408;
wire x_409;
wire x_410;
wire x_411;
wire x_412;
wire x_413;
wire x_414;
wire x_415;
wire x_416;
wire x_417;
wire x_418;
wire x_419;
wire x_420;
wire x_421;
wire x_422;
wire x_423;
wire x_424;
wire x_425;
wire x_426;
wire x_427;
wire x_428;
wire x_429;
wire x_430;
wire x_431;
wire x_432;
wire x_433;
wire x_434;
wire x_435;
wire x_436;
wire x_437;
wire x_438;
wire x_439;
wire x_440;
wire x_441;
wire x_442;
wire x_443;
wire x_444;
wire x_445;
wire x_446;
wire x_447;
wire x_448;
wire x_449;
wire x_450;
wire x_451;
wire x_452;
wire x_453;
wire x_454;
wire x_455;
wire x_456;
wire x_457;
wire x_458;
wire x_459;
wire x_460;
wire x_461;
wire x_462;
wire x_463;
wire x_464;
wire x_465;
wire x_466;
wire x_467;
wire x_468;
wire x_469;
wire x_470;
wire x_471;
wire x_472;
wire x_473;
wire x_474;
wire x_475;
wire x_476;
wire x_477;
wire x_478;
wire x_479;
wire x_480;
wire x_481;
wire x_482;
wire x_483;
wire x_484;
wire x_485;
wire x_486;
wire x_487;
wire x_488;
wire x_489;
wire x_490;
wire x_491;
wire x_492;
wire x_493;
wire x_494;
wire x_495;
wire x_496;
wire x_497;
wire x_498;
wire x_499;
wire x_500;
wire x_501;
wire x_502;
wire x_503;
wire x_504;
wire x_505;
wire x_506;
wire x_507;
wire x_508;
wire x_509;
wire x_510;
wire x_511;
wire x_512;
wire x_513;
wire x_514;
wire x_515;
wire x_516;
wire x_517;
wire x_518;
wire x_519;
wire x_520;
wire x_521;
wire x_522;
wire x_523;
wire x_524;
wire x_525;
wire x_526;
wire x_527;
wire x_528;
wire x_529;
wire x_530;
wire x_531;
wire x_532;
wire x_533;
wire x_534;
wire x_535;
wire x_536;
wire x_537;
wire x_538;
wire x_539;
wire x_540;
wire x_541;
wire x_542;
wire x_543;
wire x_544;
wire x_545;
wire x_546;
wire x_547;
wire x_548;
wire x_549;
wire x_550;
wire x_551;
wire x_552;
wire x_553;
wire x_554;
wire x_555;
wire x_556;
wire x_557;
wire x_558;
wire x_559;
wire x_560;
wire x_561;
wire x_562;
wire x_563;
wire x_564;
wire x_565;
wire x_566;
wire x_567;
wire x_568;
wire x_569;
wire x_570;
wire x_571;
wire x_572;
wire x_573;
wire x_574;
wire x_575;
wire x_576;
wire x_577;
wire x_578;
wire x_579;
wire x_580;
wire x_581;
wire x_582;
wire x_583;
wire x_584;
wire x_585;
wire x_586;
wire x_587;
wire x_588;
wire x_589;
wire x_590;
wire x_591;
wire x_592;
wire x_593;
wire x_594;
wire x_595;
wire x_596;
wire x_597;
wire x_598;
wire x_599;
wire x_600;
wire x_601;
wire x_602;
wire x_603;
wire x_604;
wire x_605;
wire x_606;
wire x_607;
wire x_608;
wire x_609;
wire x_610;
wire x_611;
wire x_612;
wire x_613;
wire x_614;
wire x_615;
wire x_616;
wire x_617;
wire x_618;
wire x_619;
wire x_620;
wire x_621;
wire x_622;
wire x_623;
wire x_624;
wire x_625;
wire x_626;
wire x_627;
wire x_628;
wire x_629;
wire x_630;
wire x_631;
wire x_632;
wire x_633;
wire x_634;
wire x_635;
wire x_636;
wire x_637;
wire x_638;
wire x_639;
wire x_640;
wire x_641;
wire x_642;
wire x_643;
wire x_644;
wire x_645;
wire x_646;
wire x_647;
wire x_648;
wire x_649;
wire x_650;
wire x_651;
wire x_652;
wire x_653;
wire x_654;
wire x_655;
wire x_656;
wire x_657;
wire x_658;
wire x_659;
wire x_660;
wire x_661;
wire x_662;
wire x_663;
wire x_664;
wire x_665;
wire x_666;
wire x_667;
wire x_668;
wire x_669;
wire x_670;
wire x_671;
wire x_672;
wire x_673;
wire x_674;
wire x_675;
wire x_676;
wire x_677;
wire x_678;
wire x_679;
wire x_680;
wire x_681;
wire x_682;
wire x_683;
wire x_684;
wire x_685;
wire x_686;
wire x_687;
wire x_688;
wire x_689;
wire x_690;
wire x_691;
wire x_692;
wire x_693;
wire x_694;
wire x_695;
wire x_696;
wire x_697;
wire x_698;
wire x_699;
wire x_700;
wire x_701;
wire x_702;
wire x_703;
wire x_704;
wire x_705;
wire x_706;
wire x_707;
wire x_708;
wire x_709;
wire x_710;
wire x_711;
wire x_712;
wire x_713;
wire x_714;
wire x_715;
wire x_716;
wire x_717;
wire x_718;
wire x_719;
wire x_720;
wire x_721;
wire x_722;
wire x_723;
wire x_724;
wire x_725;
wire x_726;
wire x_727;
wire x_728;
wire x_729;
wire x_730;
wire x_731;
wire x_732;
wire x_733;
wire x_734;
wire x_735;
wire x_736;
wire x_737;
wire x_738;
wire x_739;
wire x_740;
wire x_741;
wire x_742;
wire x_743;
wire x_744;
wire x_745;
wire x_746;
wire x_747;
wire x_748;
wire x_749;
wire x_750;
wire x_751;
wire x_752;
wire x_753;
wire x_754;
wire x_755;
wire x_756;
wire x_757;
wire x_758;
wire x_759;
wire x_760;
wire x_761;
wire x_762;
wire x_763;
wire x_764;
wire x_765;
wire x_766;
wire x_767;
wire x_768;
wire x_769;
wire x_770;
wire x_771;
wire x_772;
wire x_773;
wire x_774;
wire x_775;
wire x_776;
wire x_777;
wire x_778;
wire x_779;
wire x_780;
wire x_781;
wire x_782;
wire x_783;
wire x_784;
wire x_785;
wire x_786;
wire x_787;
wire x_788;
wire x_789;
wire x_790;
wire x_791;
wire x_792;
wire x_793;
wire x_794;
wire x_795;
wire x_796;
wire x_797;
wire x_798;
wire x_799;
wire x_800;
wire x_801;
wire x_802;
wire x_803;
wire x_804;
wire x_805;
wire x_806;
wire x_807;
wire x_808;
wire x_809;
wire x_810;
wire x_811;
wire x_812;
wire x_813;
wire x_814;
wire x_815;
wire x_816;
wire x_817;
wire x_818;
wire x_819;
wire x_820;
wire x_821;
wire x_822;
wire x_823;
wire x_824;
wire x_825;
wire x_826;
wire x_827;
wire x_828;
wire x_829;
wire x_830;
wire x_831;
wire x_832;
wire x_833;
wire x_834;
wire x_835;
wire x_836;
wire x_837;
wire x_838;
wire x_839;
wire x_840;
wire x_841;
wire x_842;
wire x_843;
wire x_844;
wire x_845;
wire x_846;
wire x_847;
wire x_848;
wire x_849;
wire x_850;
wire x_851;
wire x_852;
wire x_853;
wire x_854;
wire x_855;
wire x_856;
wire x_857;
wire x_858;
wire x_859;
wire x_860;
wire x_861;
wire x_862;
wire x_863;
wire x_864;
wire x_865;
wire x_866;
wire x_867;
wire x_868;
wire x_869;
wire x_870;
wire x_871;
wire x_872;
wire x_873;
wire x_874;
wire x_875;
wire x_876;
wire x_877;
wire x_878;
wire x_879;
wire x_880;
wire x_881;
wire x_882;
wire x_883;
wire x_884;
wire x_885;
wire x_886;
wire x_887;
wire x_888;
wire x_889;
wire x_890;
wire x_891;
wire x_892;
wire x_893;
wire x_894;
wire x_895;
wire x_896;
wire x_897;
wire x_898;
wire x_899;
wire x_900;
wire x_901;
wire x_902;
wire x_903;
wire x_904;
wire x_905;
wire x_906;
wire x_907;
wire x_908;
wire x_909;
wire x_910;
wire x_911;
wire x_912;
wire x_913;
wire x_914;
wire x_915;
wire x_916;
wire x_917;
wire x_918;
wire x_919;
wire x_920;
wire x_921;
wire x_922;
wire x_923;
wire x_924;
wire x_925;
wire x_926;
wire x_927;
wire x_928;
wire x_929;
wire x_930;
wire x_931;
wire x_932;
wire x_933;
wire x_934;
wire x_935;
wire x_936;
wire x_937;
wire x_938;
wire x_939;
wire x_940;
wire x_941;
wire x_942;
wire x_943;
wire x_944;
wire x_945;
wire x_946;
wire x_947;
wire x_948;
wire x_949;
wire x_950;
wire x_951;
wire x_952;
wire x_953;
wire x_954;
wire x_955;
wire x_956;
wire x_957;
wire x_958;
wire x_959;
wire x_960;
wire x_961;
wire x_962;
wire x_963;
wire x_964;
wire x_965;
wire x_966;
wire x_967;
wire x_968;
wire x_969;
wire x_970;
wire x_971;
wire x_972;
wire x_973;
wire x_974;
wire x_975;
wire x_976;
wire x_977;
wire x_978;
wire x_979;
wire x_980;
wire x_981;
wire x_982;
wire x_983;
wire x_984;
wire x_985;
wire x_986;
wire x_987;
wire x_988;
wire x_989;
wire x_990;
wire x_991;
wire x_992;
wire x_993;
wire x_994;
wire x_995;
wire x_996;
wire x_997;
wire x_998;
wire x_999;
wire x_1000;
wire x_1001;
wire x_1002;
wire x_1003;
wire x_1004;
wire x_1005;
wire x_1006;
wire x_1007;
wire x_1008;
wire x_1009;
wire x_1010;
wire x_1011;
wire x_1012;
wire x_1013;
wire x_1014;
wire x_1015;
wire x_1016;
wire x_1017;
wire x_1018;
wire x_1019;
wire x_1020;
wire x_1021;
wire x_1022;
wire x_1023;
wire x_1024;
wire x_1025;
wire x_1026;
wire x_1027;
wire x_1028;
wire x_1029;
wire x_1030;
wire x_1031;
wire x_1032;
wire x_1033;
wire x_1034;
wire x_1035;
wire x_1036;
wire x_1037;
wire x_1038;
wire x_1039;
wire x_1040;
wire x_1041;
wire x_1042;
wire x_1043;
wire x_1044;
wire x_1045;
wire x_1046;
wire x_1047;
wire x_1048;
wire x_1049;
wire x_1050;
wire x_1051;
wire x_1052;
wire x_1053;
wire x_1054;
wire x_1055;
wire x_1056;
wire x_1057;
wire x_1058;
wire x_1059;
wire x_1060;
wire x_1061;
wire x_1062;
wire x_1063;
wire x_1064;
wire x_1065;
wire x_1066;
wire x_1067;
wire x_1068;
wire x_1069;
wire x_1070;
wire x_1071;
wire x_1072;
wire x_1073;
wire x_1074;
wire x_1075;
wire x_1076;
wire x_1077;
wire x_1078;
wire x_1079;
wire x_1080;
wire x_1081;
wire x_1082;
wire x_1083;
wire x_1084;
wire x_1085;
wire x_1086;
wire x_1087;
wire x_1088;
wire x_1089;
wire x_1090;
wire x_1091;
wire x_1092;
wire x_1093;
wire x_1094;
wire x_1095;
wire x_1096;
wire x_1097;
wire x_1098;
wire x_1099;
wire x_1100;
wire x_1101;
wire x_1102;
wire x_1103;
wire x_1104;
wire x_1105;
wire x_1106;
wire x_1107;
wire x_1108;
wire x_1109;
wire x_1110;
wire x_1111;
wire x_1112;
wire x_1113;
wire x_1114;
wire x_1115;
wire x_1116;
wire x_1117;
wire x_1118;
wire x_1119;
wire x_1120;
wire x_1121;
wire x_1122;
wire x_1123;
wire x_1124;
wire x_1125;
wire x_1126;
wire x_1127;
wire x_1128;
wire x_1129;
wire x_1130;
wire x_1131;
wire x_1132;
wire x_1133;
wire x_1134;
wire x_1135;
wire x_1136;
wire x_1137;
wire x_1138;
wire x_1139;
wire x_1140;
wire x_1141;
wire x_1142;
wire x_1143;
wire x_1144;
wire x_1145;
wire x_1146;
wire x_1147;
wire x_1148;
wire x_1149;
wire x_1150;
wire x_1151;
wire x_1152;
wire x_1153;
assign v_4 = 0;
assign v_2 = 1;
assign v_3 = 1;
assign v_409 = 1;
assign v_7 = v_8 & v_9;
assign v_9 = ~v_10 & ~v_18 & v_14;
assign v_12 = ~v_287 & ~v_288;
assign v_15 = v_288 & v_289;
assign v_17 = ~v_14 & ~v_287;
assign v_19 = ~v_289 & v_291;
assign v_21 = v_8 & v_14 & v_22;
assign v_22 = ~v_10 & v_18;
assign v_23 = ~v_338 & v_339;
assign v_26 = v_338 & v_27;
assign v_27 = ~v_10 & ~v_14 & ~v_18 & v_8;
assign v_28 = ~v_29 & v_33 & v_46 & v_138;
assign v_31 = ~v_14 & v_22 & v_32;
assign v_36 = ~v_37 & v_38;
assign v_40 = ~v_27 & v_280 & v_41 & v_43;
assign v_41 = v_42 & v_9;
assign v_43 = ~v_296 & ~v_297 & v_340;
assign v_47 = ~v_7 & v_282;
assign v_52 = ~v_338 & v_329 & v_339;
assign v_55 = ~v_56 & ~v_90 & v_58 & v_95;
assign v_57 = ~v_296 & ~v_297;
assign v_58 = ~v_81 & ~v_87 & v_59 & v_69;
assign v_61 = ~v_324 & v_325;
assign v_63 = ~v_261 & v_262;
assign v_64 = v_65 & v_66 & v_67;
assign v_66 = ~v_298 & ~v_333 & v_299 & v_334;
assign v_75 = v_342 & v_76 & v_77 & v_78;
assign v_78 = v_79 & v_80;
assign v_86 = ~v_327 & v_328;
assign v_88 = v_65 & v_89;
assign v_92 = ~v_93 & ~v_94 & v_284 & v_321;
assign v_93 = ~v_292 & ~v_293;
assign v_94 = ~v_314 & v_315;
assign v_95 = v_96 & v_107 & v_115 & v_123;
assign v_97 = v_98 & v_99 & v_100 & v_101;
assign v_106 = ~v_264 & v_265;
assign v_109 = ~v_251 & v_252;
assign v_111 = ~v_256 & v_257;
assign v_112 = ~v_319 & v_320;
assign v_114 = ~v_303 & v_280;
assign v_121 = ~v_249 & ~v_250;
assign v_122 = ~v_312 & ~v_313;
assign v_124 = ~v_314 & ~v_315;
assign v_125 = ~v_251 & ~v_252;
assign v_127 = ~v_216 & ~v_278;
assign v_128 = ~v_279 & ~v_341;
assign v_129 = ~v_249 & v_250;
assign v_130 = ~v_312 & v_313;
assign v_133 = ~v_253 & v_254;
assign v_134 = ~v_316 & v_317;
assign v_136 = ~v_285 & ~v_286;
assign v_137 = ~v_222 & ~v_223;
assign v_142 = ~v_304 & ~v_305 & v_338;
assign v_150 = ~v_62 & ~v_105 & ~v_154 & v_151;
assign v_151 = v_152 & v_153 & v_125 & v_127;
assign v_152 = ~v_260 & ~v_261;
assign v_153 = ~v_263 & ~v_264;
assign v_155 = v_156 & v_160 & v_162 & v_163;
assign v_157 = ~v_268 & v_269;
assign v_158 = ~v_275 & ~v_276 & ~v_277 & v_159;
assign v_159 = ~v_267 & ~v_272 & ~v_273 & ~v_274;
assign v_160 = ~v_249 & ~v_250 & v_137 & v_161;
assign v_161 = ~v_217 & ~v_218 & ~v_219 & ~v_221;
assign v_162 = ~v_257 & ~v_258 & ~v_259 & ~v_266;
assign v_163 = ~v_253 & ~v_254 & ~v_255 & ~v_256;
assign v_164 = v_97 & v_165 & v_176 & v_190;
assign v_165 = v_166 & v_169 & v_170 & v_173;
assign v_167 = ~v_325 & v_262;
assign v_168 = ~v_227 & v_290;
assign v_171 = ~v_308 & v_245;
assign v_172 = ~v_226 & v_289;
assign v_174 = ~v_290 & v_227;
assign v_175 = ~v_245 & v_308;
assign v_176 = v_177 & v_181 & v_184 & v_187;
assign v_178 = ~v_301 & v_238;
assign v_180 = ~v_238 & v_301;
assign v_182 = ~v_261 & v_324;
assign v_183 = ~v_317 & v_254;
assign v_185 = ~v_264 & v_327;
assign v_186 = ~v_262 & v_325;
assign v_188 = ~v_234 & v_297;
assign v_189 = ~v_327 & v_264;
assign v_190 = v_191 & v_79 & v_80 & v_192;
assign v_194 = v_195 & v_206 & v_214 & v_215;
assign v_195 = v_77 & v_196 & v_202 & v_203;
assign v_196 = v_24 & v_197 & v_198 & v_199;
assign v_203 = v_204 & v_50 & v_74 & v_205;
assign v_206 = v_207 & v_210 & v_211 & v_212;
assign v_214 = v_38 & v_141 & v_147 & v_149;
assign v_215 = v_30 & v_73 & v_110 & v_117;
assign v_13 = v_10 ^ ~v_11;
assign v_24 = ~v_258 ^ v_321;
assign v_30 = ~v_266 ^ v_329;
assign v_38 = ~v_275 ^ v_338;
assign v_50 = ~v_259 ^ v_322;
assign v_60 = v_323 ^ v_61;
assign v_62 = v_260 ^ v_63;
assign v_73 = ~v_236 ^ v_299;
assign v_74 = ~v_230 ^ v_293;
assign v_76 = ~v_278 ^ v_341;
assign v_83 = v_301 ^ v_334;
assign v_85 = v_326 ^ v_86;
assign v_91 = v_90 ^ v_246;
assign v_105 = v_263 ^ v_106;
assign v_110 = ~v_242 ^ v_305;
assign v_117 = ~v_248 ^ v_311;
assign v_141 = ~v_274 ^ v_337;
assign v_147 = ~v_277 ^ v_340;
assign v_149 = ~v_218 ^ v_281;
assign v_197 = ~v_272 ^ v_335;
assign v_201 = ~v_217 ^ v_280;
assign v_204 = ~v_276 ^ v_339;
assign v_205 = ~v_269 ^ v_332;
assign v_209 = v_239 ^ v_302;
assign x_1 = ~v_194 | v_342 | v_5 | ~v_164;
assign x_2 = ~v_194 | ~v_342 | ~v_5 | ~v_164;
assign x_3 = v_5 | ~v_343 | ~v_6;
assign x_4 = v_5 | v_343 | ~v_150 | ~v_155;
assign x_5 = v_343 | v_150 | ~v_5;
assign x_6 = v_6 | ~v_5 | ~v_343;
assign x_7 = v_343 | v_155 | ~v_5;
assign x_8 = v_6 | ~v_7 | ~v_28;
assign x_9 = v_6 | v_20 | v_25 | ~v_28;
assign x_10 = v_28 | ~v_6;
assign x_11 = v_7 | ~v_6 | ~v_20;
assign x_12 = v_7 | ~v_6 | ~v_25;
assign x_13 = v_8 | v_287 | ~v_288 | ~v_289;
assign x_14 = v_8 | v_288 | v_290 | ~v_287;
assign x_15 = v_8 | v_288 | v_289 | ~v_287;
assign x_16 = v_289 | ~v_8 | ~v_288;
assign x_17 = ~v_8 | ~v_287 | ~v_289 | ~v_290;
assign x_18 = ~v_8 | ~v_287 | ~v_288;
assign x_19 = v_287 | v_288 | ~v_8;
assign x_20 = v_11 | v_290 | ~v_291;
assign x_21 = v_11 | v_289 | ~v_291 | ~v_12;
assign x_22 = v_291 | ~v_11;
assign x_23 = v_12 | ~v_11 | ~v_290;
assign x_24 = ~v_11 | ~v_289 | ~v_290;
assign x_25 = v_13 | v_289 | ~v_287;
assign x_26 = v_13 | v_289 | ~v_288;
assign x_27 = ~v_13 | ~v_289;
assign x_28 = v_287 | v_288 | ~v_13;
assign x_29 = v_14 | v_17 | ~v_15;
assign x_30 = v_14 | v_17 | ~v_16;
assign x_31 = v_15 | v_16 | ~v_14 | ~v_287;
assign x_32 = v_16 | v_288 | v_289 | ~v_291;
assign x_33 = v_16 | v_288 | v_290 | ~v_289;
assign x_34 = v_16 | v_288 | v_289 | ~v_290;
assign x_35 = ~v_16 | ~v_288;
assign x_36 = ~v_16 | ~v_289 | ~v_290;
assign x_37 = v_289 | v_290 | v_291 | ~v_16;
assign x_38 = v_17 | v_287 | ~v_288 | ~v_289;
assign x_39 = v_17 | v_287 | v_290 | ~v_289;
assign x_40 = v_17 | v_287 | v_288 | v_289 | ~v_290;
assign x_41 = v_289 | ~v_17 | ~v_288;
assign x_42 = v_289 | v_290 | ~v_17;
assign x_43 = v_288 | ~v_17 | ~v_289 | ~v_290;
assign x_44 = v_18 | ~v_288 | ~v_19;
assign x_45 = v_18 | v_288 | v_290 | v_19;
assign x_46 = v_18 | ~v_288 | ~v_290;
assign x_47 = v_18 | v_287 | v_290 | ~v_19;
assign x_48 = v_288 | ~v_18 | ~v_290;
assign x_49 = v_290 | v_19 | ~v_18 | ~v_288;
assign x_50 = v_288 | ~v_18 | ~v_287 | ~v_19;
assign x_51 = v_20 | ~v_258 | ~v_21 | ~v_23;
assign x_52 = v_20 | v_23 | v_24 | ~v_21;
assign x_53 = v_21 | ~v_20;
assign x_54 = v_23 | ~v_20 | ~v_24;
assign x_55 = v_258 | ~v_20 | ~v_23;
assign x_56 = v_25 | v_21 | v_24 | v_26;
assign x_57 = v_25 | v_21 | ~v_258 | ~v_26;
assign x_58 = ~v_25 | ~v_21;
assign x_59 = v_258 | ~v_25 | ~v_26;
assign x_60 = v_26 | ~v_25 | ~v_24;
assign x_61 = v_29 | v_31 | ~v_266 | ~v_26;
assign x_62 = v_29 | v_26 | v_30 | v_31;
assign x_63 = ~v_29 | ~v_31;
assign x_64 = v_266 | ~v_29 | ~v_26;
assign x_65 = v_26 | ~v_29 | ~v_30;
assign x_66 = v_32 | v_287 | v_288 | ~v_290;
assign x_67 = v_32 | v_287 | v_289 | ~v_288;
assign x_68 = v_32 | v_287 | v_288 | ~v_289;
assign x_69 = ~v_32 | ~v_287;
assign x_70 = ~v_32 | ~v_288 | ~v_289;
assign x_71 = v_288 | v_289 | v_290 | ~v_32;
assign x_72 = v_33 | ~v_39 | ~v_40;
assign x_73 = v_33 | v_44 | ~v_34;
assign x_74 = v_33 | ~v_34 | ~v_40;
assign x_75 = v_33 | v_44 | ~v_39;
assign x_76 = v_40 | ~v_33 | ~v_44;
assign x_77 = v_34 | v_39 | ~v_33;
assign x_78 = v_34 | v_21 | v_27 | ~v_36;
assign x_79 = v_34 | v_21 | ~v_27 | ~v_35;
assign x_80 = ~v_34 | ~v_21;
assign x_81 = v_35 | ~v_34 | ~v_27;
assign x_82 = v_27 | v_36 | ~v_34;
assign x_83 = v_35 | v_275 | v_276 | v_339;
assign x_84 = v_35 | v_275 | v_276 | ~v_338;
assign x_85 = v_35 | v_275 | v_338 | ~v_276 | ~v_339;
assign x_86 = ~v_35 | ~v_276 | ~v_338;
assign x_87 = v_339 | ~v_35 | ~v_276;
assign x_88 = ~v_35 | ~v_275;
assign x_89 = v_276 | v_338 | ~v_35 | ~v_339;
assign x_90 = v_37 | v_338 | v_339 | ~v_276;
assign x_91 = v_37 | v_276 | v_338 | ~v_339;
assign x_92 = ~v_37 | ~v_338;
assign x_93 = ~v_37 | ~v_276 | ~v_339;
assign x_94 = v_276 | v_339 | ~v_37;
assign x_95 = v_39 | ~v_275 | ~v_338 | ~v_21;
assign x_96 = v_39 | v_275 | v_276 | v_338 | ~v_21;
assign x_97 = v_338 | ~v_39 | ~v_276;
assign x_98 = v_275 | ~v_39 | ~v_338;
assign x_99 = v_21 | ~v_39;
assign x_100 = v_338 | ~v_39 | ~v_275;
assign x_101 = v_42 | ~v_287 | ~v_288;
assign x_102 = v_42 | ~v_287 | ~v_289 | ~v_290;
assign x_103 = v_287 | ~v_42;
assign x_104 = v_288 | v_290 | ~v_42;
assign x_105 = v_288 | v_289 | ~v_42;
assign x_106 = v_44 | v_280 | v_26 | ~v_217;
assign x_107 = v_44 | ~v_217 | ~v_26 | ~v_45;
assign x_108 = v_44 | v_217 | v_26 | ~v_280;
assign x_109 = v_44 | v_217 | v_45 | ~v_26;
assign x_110 = v_217 | ~v_44 | ~v_26 | ~v_45;
assign x_111 = v_26 | ~v_44 | ~v_217 | ~v_280;
assign x_112 = v_45 | ~v_44 | ~v_217 | ~v_26;
assign x_113 = v_217 | v_280 | v_26 | ~v_44;
assign x_114 = v_45 | v_337 | ~v_304;
assign x_115 = v_45 | v_337 | ~v_305;
assign x_116 = ~v_45 | ~v_337;
assign x_117 = v_304 | v_305 | ~v_45;
assign x_118 = v_46 | v_219 | v_47 | ~v_48 | ~v_55;
assign x_119 = v_46 | ~v_219 | ~v_47 | ~v_48 | ~v_55;
assign x_120 = v_55 | ~v_46;
assign x_121 = v_47 | ~v_46 | ~v_219;
assign x_122 = v_48 | ~v_46;
assign x_123 = v_219 | ~v_46 | ~v_47;
assign x_124 = v_48 | v_49 | ~v_31 | ~v_51;
assign x_125 = v_48 | v_31 | ~v_50 | ~v_51;
assign x_126 = v_51 | ~v_48;
assign x_127 = v_31 | v_50 | ~v_48;
assign x_128 = ~v_48 | ~v_31 | ~v_49;
assign x_129 = v_49 | ~v_266 | ~v_281;
assign x_130 = v_49 | v_281 | v_30;
assign x_131 = v_266 | ~v_49 | ~v_281;
assign x_132 = v_281 | ~v_49 | ~v_30;
assign x_133 = v_51 | v_52 | v_54;
assign x_134 = v_51 | v_54 | ~v_53;
assign x_135 = v_51 | v_21 | v_54;
assign x_136 = ~v_51 | ~v_54;
assign x_137 = v_53 | ~v_51 | ~v_21 | ~v_52;
assign x_138 = v_53 | ~v_268 | ~v_304;
assign x_139 = v_53 | v_268 | v_304 | ~v_269 | ~v_305;
assign x_140 = v_53 | v_268 | v_269 | v_304 | v_305;
assign x_141 = v_304 | ~v_53 | ~v_268;
assign x_142 = v_268 | v_305 | ~v_53 | ~v_269;
assign x_143 = v_268 | ~v_53 | ~v_304;
assign x_144 = v_269 | v_304 | ~v_53 | ~v_305;
assign x_145 = v_54 | v_282 | v_24 | ~v_7;
assign x_146 = v_54 | ~v_258 | ~v_282 | ~v_7;
assign x_147 = v_7 | ~v_54;
assign x_148 = v_258 | ~v_54 | ~v_282;
assign x_149 = v_282 | ~v_54 | ~v_24;
assign x_150 = v_56 | v_335 | ~v_272;
assign x_151 = v_56 | v_272 | v_41 | ~v_335;
assign x_152 = v_56 | v_272 | v_57 | ~v_335;
assign x_153 = ~v_56 | ~v_272 | ~v_335;
assign x_154 = v_272 | v_335 | ~v_56;
assign x_155 = v_272 | ~v_56 | ~v_41 | ~v_57;
assign x_156 = v_59 | v_60 | v_62 | v_64 | v_68;
assign x_157 = v_59 | v_64 | v_68 | ~v_60 | ~v_62;
assign x_158 = ~v_59 | ~v_64;
assign x_159 = v_62 | ~v_59 | ~v_60;
assign x_160 = ~v_59 | ~v_68;
assign x_161 = v_60 | ~v_59 | ~v_62;
assign x_162 = v_65 | v_323 | ~v_324;
assign x_163 = v_65 | v_324 | v_325 | ~v_323;
assign x_164 = ~v_65 | ~v_323 | ~v_324;
assign x_165 = v_324 | ~v_65 | ~v_325;
assign x_166 = v_323 | v_324 | ~v_65;
assign x_167 = v_67 | v_334 | ~v_310;
assign x_168 = v_67 | v_311 | ~v_333;
assign x_169 = v_67 | v_311 | v_334;
assign x_170 = v_67 | ~v_310 | ~v_333;
assign x_171 = v_310 | ~v_67 | ~v_311;
assign x_172 = v_333 | ~v_67 | ~v_334;
assign x_173 = v_68 | v_333 | ~v_270;
assign x_174 = v_68 | v_270 | v_334 | ~v_271;
assign x_175 = v_68 | v_270 | ~v_333;
assign x_176 = v_68 | v_271 | v_333 | ~v_334;
assign x_177 = ~v_68 | ~v_270 | ~v_333;
assign x_178 = v_270 | v_333 | ~v_68 | ~v_271 | ~v_334;
assign x_179 = v_270 | v_271 | v_333 | v_334 | ~v_68;
assign x_180 = v_69 | v_70 | v_71 | ~v_72 | ~v_75;
assign x_181 = v_69 | ~v_70 | ~v_71 | ~v_72 | ~v_75;
assign x_182 = v_75 | ~v_69;
assign x_183 = v_71 | ~v_69 | ~v_70;
assign x_184 = v_72 | ~v_69;
assign x_185 = v_70 | ~v_69 | ~v_71;
assign x_186 = v_70 | ~v_326 | ~v_327;
assign x_187 = v_70 | ~v_326 | ~v_328;
assign x_188 = v_326 | ~v_70;
assign x_189 = v_327 | v_328 | ~v_70;
assign x_190 = v_71 | ~v_263 | ~v_264;
assign x_191 = v_71 | ~v_263 | ~v_265;
assign x_192 = v_263 | ~v_71;
assign x_193 = v_264 | v_265 | ~v_71;
assign x_194 = v_72 | ~v_229 | ~v_73;
assign x_195 = v_72 | ~v_235 | ~v_74;
assign x_196 = v_72 | ~v_229 | ~v_235;
assign x_197 = v_72 | ~v_73 | ~v_74;
assign x_198 = v_235 | v_73 | ~v_72;
assign x_199 = v_229 | v_74 | ~v_72;
assign x_200 = v_77 | v_235 | v_298 | ~v_229 | ~v_292;
assign x_201 = v_77 | v_229 | v_292 | ~v_235 | ~v_298;
assign x_202 = v_77 | v_229 | v_235 | v_292 | v_298;
assign x_203 = v_77 | ~v_229 | ~v_235 | ~v_292 | ~v_298;
assign x_204 = v_292 | ~v_77 | ~v_229;
assign x_205 = v_229 | ~v_77 | ~v_292;
assign x_206 = v_235 | ~v_77 | ~v_298;
assign x_207 = v_298 | ~v_77 | ~v_235;
assign x_208 = v_79 | v_247 | v_310 | ~v_244 | ~v_307;
assign x_209 = v_79 | v_244 | v_307 | ~v_247 | ~v_310;
assign x_210 = v_79 | v_244 | v_247 | v_307 | v_310;
assign x_211 = v_79 | ~v_244 | ~v_247 | ~v_307 | ~v_310;
assign x_212 = v_307 | ~v_79 | ~v_244;
assign x_213 = v_244 | ~v_79 | ~v_307;
assign x_214 = v_247 | ~v_79 | ~v_310;
assign x_215 = v_310 | ~v_79 | ~v_247;
assign x_216 = v_80 | v_253 | v_316 | ~v_220 | ~v_283;
assign x_217 = v_80 | v_220 | v_283 | ~v_253 | ~v_316;
assign x_218 = v_80 | v_220 | v_253 | v_283 | v_316;
assign x_219 = v_80 | ~v_220 | ~v_253 | ~v_283 | ~v_316;
assign x_220 = v_283 | ~v_80 | ~v_220;
assign x_221 = v_220 | ~v_80 | ~v_283;
assign x_222 = v_253 | ~v_80 | ~v_316;
assign x_223 = v_316 | ~v_80 | ~v_253;
assign x_224 = v_81 | v_85 | ~v_285 | ~v_82;
assign x_225 = v_81 | v_285 | ~v_82 | ~v_85;
assign x_226 = v_81 | v_286 | v_85 | ~v_82;
assign x_227 = v_82 | ~v_81;
assign x_228 = ~v_81 | ~v_285 | ~v_85;
assign x_229 = v_285 | v_85 | ~v_81 | ~v_286;
assign x_230 = v_82 | v_300 | ~v_333 | ~v_84;
assign x_231 = v_82 | v_333 | ~v_300 | ~v_84;
assign x_232 = v_82 | v_300 | ~v_83 | ~v_84;
assign x_233 = v_84 | ~v_82;
assign x_234 = ~v_82 | ~v_300 | ~v_333;
assign x_235 = v_300 | v_333 | v_83 | ~v_82;
assign x_236 = v_84 | v_326 | ~v_327;
assign x_237 = v_84 | v_327 | v_328 | ~v_326;
assign x_238 = ~v_84 | ~v_326 | ~v_327;
assign x_239 = v_327 | ~v_84 | ~v_328;
assign x_240 = v_326 | v_327 | ~v_84;
assign x_241 = v_87 | v_285 | v_286 | ~v_88;
assign x_242 = v_87 | v_60 | ~v_285 | ~v_88;
assign x_243 = v_87 | v_285 | ~v_60 | ~v_88;
assign x_244 = v_88 | ~v_87;
assign x_245 = ~v_87 | ~v_285 | ~v_60;
assign x_246 = v_285 | v_60 | ~v_87 | ~v_286;
assign x_247 = v_89 | v_333 | ~v_298;
assign x_248 = v_89 | v_298 | v_334 | ~v_299;
assign x_249 = v_89 | v_298 | ~v_333;
assign x_250 = v_89 | v_299 | v_333 | ~v_334;
assign x_251 = ~v_89 | ~v_298 | ~v_333;
assign x_252 = v_298 | v_333 | ~v_89 | ~v_299 | ~v_334;
assign x_253 = v_298 | v_299 | v_333 | v_334 | ~v_89;
assign x_254 = v_91 | ~v_309 | ~v_92;
assign x_255 = v_91 | v_92 | ~v_283;
assign x_256 = v_283 | v_92 | ~v_91;
assign x_257 = v_309 | ~v_91 | ~v_92;
assign x_258 = v_96 | v_65 | v_102 | ~v_97 | ~v_103;
assign x_259 = v_96 | ~v_65 | ~v_97 | ~v_102 | ~v_103;
assign x_260 = v_103 | ~v_96;
assign x_261 = v_102 | ~v_96 | ~v_65;
assign x_262 = v_97 | ~v_96;
assign x_263 = v_65 | ~v_96 | ~v_102;
assign x_264 = v_98 | v_273 | v_336 | ~v_241 | ~v_304;
assign x_265 = v_98 | v_241 | v_304 | ~v_273 | ~v_336;
assign x_266 = v_98 | v_241 | v_273 | v_304 | v_336;
assign x_267 = v_98 | ~v_241 | ~v_273 | ~v_304 | ~v_336;
assign x_268 = v_304 | ~v_98 | ~v_241;
assign x_269 = v_241 | ~v_98 | ~v_304;
assign x_270 = v_273 | ~v_98 | ~v_336;
assign x_271 = v_336 | ~v_98 | ~v_273;
assign x_272 = v_99 | v_256 | v_319 | ~v_221 | ~v_284;
assign x_273 = v_99 | v_221 | v_284 | ~v_256 | ~v_319;
assign x_274 = v_99 | v_221 | v_256 | v_284 | v_319;
assign x_275 = v_99 | ~v_221 | ~v_256 | ~v_284 | ~v_319;
assign x_276 = v_284 | ~v_99 | ~v_221;
assign x_277 = v_221 | ~v_99 | ~v_284;
assign x_278 = v_256 | ~v_99 | ~v_319;
assign x_279 = v_319 | ~v_99 | ~v_256;
assign x_280 = v_100 | v_243 | v_306 | ~v_222 | ~v_285;
assign x_281 = v_100 | v_222 | v_285 | ~v_243 | ~v_306;
assign x_282 = v_100 | v_222 | v_243 | v_285 | v_306;
assign x_283 = v_100 | ~v_222 | ~v_243 | ~v_285 | ~v_306;
assign x_284 = v_285 | ~v_100 | ~v_222;
assign x_285 = v_222 | ~v_100 | ~v_285;
assign x_286 = v_243 | ~v_100 | ~v_306;
assign x_287 = v_306 | ~v_100 | ~v_243;
assign x_288 = v_101 | v_267 | v_330 | ~v_255 | ~v_318;
assign x_289 = v_101 | v_255 | v_318 | ~v_267 | ~v_330;
assign x_290 = v_101 | v_255 | v_267 | v_318 | v_330;
assign x_291 = v_101 | ~v_255 | ~v_267 | ~v_318 | ~v_330;
assign x_292 = v_318 | ~v_101 | ~v_255;
assign x_293 = v_255 | ~v_101 | ~v_318;
assign x_294 = v_267 | ~v_101 | ~v_330;
assign x_295 = v_330 | ~v_101 | ~v_267;
assign x_296 = v_102 | v_260 | ~v_261;
assign x_297 = v_102 | v_261 | v_262 | ~v_260;
assign x_298 = ~v_102 | ~v_260 | ~v_261;
assign x_299 = v_261 | ~v_102 | ~v_262;
assign x_300 = v_260 | v_261 | ~v_102;
assign x_301 = v_103 | v_85 | v_105 | ~v_84 | ~v_104;
assign x_302 = v_103 | v_84 | v_104 | ~v_85 | ~v_105;
assign x_303 = v_103 | v_84 | v_85 | v_104 | v_105;
assign x_304 = v_103 | ~v_84 | ~v_85 | ~v_104 | ~v_105;
assign x_305 = v_104 | ~v_103 | ~v_84;
assign x_306 = v_84 | ~v_103 | ~v_104;
assign x_307 = v_85 | ~v_103 | ~v_105;
assign x_308 = v_105 | ~v_103 | ~v_85;
assign x_309 = v_104 | v_263 | ~v_264;
assign x_310 = v_104 | v_264 | v_265 | ~v_263;
assign x_311 = ~v_104 | ~v_263 | ~v_264;
assign x_312 = v_264 | ~v_104 | ~v_265;
assign x_313 = v_263 | v_264 | ~v_104;
assign x_314 = v_107 | v_113 | ~v_108 | ~v_111 | ~v_112;
assign x_315 = v_107 | v_111 | v_112 | v_113 | ~v_108;
assign x_316 = ~v_107 | ~v_113;
assign x_317 = v_112 | ~v_107 | ~v_111;
assign x_318 = v_108 | ~v_107;
assign x_319 = v_111 | ~v_107 | ~v_112;
assign x_320 = v_108 | v_94 | v_109 | ~v_241;
assign x_321 = v_108 | ~v_241 | ~v_94 | ~v_109;
assign x_322 = v_108 | v_94 | v_109 | ~v_110;
assign x_323 = v_108 | ~v_94 | ~v_109 | ~v_110;
assign x_324 = v_109 | ~v_108 | ~v_94;
assign x_325 = v_94 | ~v_108 | ~v_109;
assign x_326 = v_241 | v_110 | ~v_108;
assign x_327 = v_113 | v_57 | ~v_114;
assign x_328 = v_113 | v_302 | v_57 | ~v_337;
assign x_329 = ~v_113 | ~v_57;
assign x_330 = v_114 | ~v_113 | ~v_302;
assign x_331 = v_337 | v_114 | ~v_113;
assign x_332 = v_115 | v_116 | ~v_247 | ~v_118;
assign x_333 = v_115 | v_116 | ~v_117 | ~v_118;
assign x_334 = v_118 | ~v_115;
assign x_335 = ~v_115 | ~v_116;
assign x_336 = v_247 | v_117 | ~v_115;
assign x_337 = v_116 | v_237 | ~v_300;
assign x_338 = v_116 | v_237 | v_301 | ~v_238;
assign x_339 = ~v_116 | ~v_237;
assign x_340 = v_300 | ~v_116 | ~v_301;
assign x_341 = v_238 | v_300 | ~v_116;
assign x_342 = v_118 | v_119 | ~v_121 | ~v_122;
assign x_343 = v_118 | v_121 | v_122 | ~v_120;
assign x_344 = v_118 | v_119 | v_121 | v_122;
assign x_345 = v_118 | ~v_120 | ~v_121 | ~v_122;
assign x_346 = v_121 | ~v_118 | ~v_122;
assign x_347 = v_122 | ~v_118 | ~v_121;
assign x_348 = v_120 | ~v_118 | ~v_119;
assign x_349 = v_119 | ~v_323 | ~v_324;
assign x_350 = v_119 | ~v_323 | ~v_325;
assign x_351 = v_323 | ~v_119;
assign x_352 = v_324 | v_325 | ~v_119;
assign x_353 = v_120 | ~v_260 | ~v_261;
assign x_354 = v_120 | ~v_260 | ~v_262;
assign x_355 = v_260 | ~v_120;
assign x_356 = v_261 | v_262 | ~v_120;
assign x_357 = v_123 | v_124 | v_125 | ~v_126 | ~v_131;
assign x_358 = v_123 | ~v_124 | ~v_125 | ~v_126 | ~v_131;
assign x_359 = v_131 | ~v_123;
assign x_360 = v_125 | ~v_123 | ~v_124;
assign x_361 = v_126 | ~v_123;
assign x_362 = v_124 | ~v_123 | ~v_125;
assign x_363 = v_126 | v_127 | v_128 | ~v_129 | ~v_130;
assign x_364 = v_126 | ~v_127 | ~v_128 | ~v_129 | ~v_130;
assign x_365 = v_126 | v_127 | v_128 | v_129 | v_130;
assign x_366 = v_126 | v_129 | v_130 | ~v_127 | ~v_128;
assign x_367 = v_127 | ~v_126 | ~v_128;
assign x_368 = v_128 | ~v_126 | ~v_127;
assign x_369 = v_129 | ~v_126 | ~v_130;
assign x_370 = v_130 | ~v_126 | ~v_129;
assign x_371 = v_131 | v_132 | v_133 | v_134 | ~v_135;
assign x_372 = v_131 | v_132 | ~v_133 | ~v_134 | ~v_135;
assign x_373 = v_135 | ~v_131;
assign x_374 = v_134 | ~v_131 | ~v_133;
assign x_375 = ~v_131 | ~v_132;
assign x_376 = v_133 | ~v_131 | ~v_134;
assign x_377 = v_132 | v_300 | ~v_237;
assign x_378 = v_132 | v_238 | v_300 | ~v_301;
assign x_379 = ~v_132 | ~v_300;
assign x_380 = v_237 | ~v_132 | ~v_238;
assign x_381 = v_237 | v_301 | ~v_132;
assign x_382 = v_135 | v_120 | v_136 | v_137;
assign x_383 = v_135 | ~v_119 | ~v_136 | ~v_137;
assign x_384 = v_135 | v_136 | v_137 | ~v_119;
assign x_385 = v_135 | v_120 | ~v_136 | ~v_137;
assign x_386 = v_136 | ~v_135 | ~v_137;
assign x_387 = v_137 | ~v_135 | ~v_136;
assign x_388 = v_119 | ~v_135 | ~v_120;
assign x_389 = v_138 | v_27 | v_139 | ~v_143;
assign x_390 = v_138 | ~v_27 | ~v_140 | ~v_143;
assign x_391 = v_143 | ~v_138;
assign x_392 = v_27 | ~v_138 | ~v_139;
assign x_393 = v_140 | ~v_138 | ~v_27;
assign x_394 = v_139 | v_337 | ~v_274;
assign x_395 = v_139 | v_274 | v_41 | ~v_337;
assign x_396 = v_139 | v_274 | v_43 | ~v_337;
assign x_397 = ~v_139 | ~v_274 | ~v_337;
assign x_398 = v_274 | v_337 | ~v_139;
assign x_399 = v_274 | ~v_139 | ~v_41 | ~v_43;
assign x_400 = v_140 | v_142 | ~v_141;
assign x_401 = v_140 | ~v_274 | ~v_142;
assign x_402 = v_141 | v_142 | ~v_140;
assign x_403 = v_274 | ~v_140 | ~v_142;
assign x_404 = v_143 | ~v_144 | ~v_145;
assign x_405 = v_143 | ~v_21 | ~v_52 | ~v_145;
assign x_406 = v_145 | ~v_143;
assign x_407 = v_21 | v_144 | ~v_143;
assign x_408 = v_52 | v_144 | ~v_143;
assign x_409 = v_144 | ~v_268 | ~v_331;
assign x_410 = v_144 | v_268 | v_331 | ~v_269 | ~v_332;
assign x_411 = v_144 | v_268 | v_269 | v_331 | v_332;
assign x_412 = v_331 | ~v_144 | ~v_268;
assign x_413 = v_268 | v_332 | ~v_144 | ~v_269;
assign x_414 = v_268 | ~v_144 | ~v_331;
assign x_415 = v_269 | v_331 | ~v_144 | ~v_332;
assign x_416 = v_145 | v_31 | v_146 | ~v_149;
assign x_417 = v_145 | v_146 | ~v_31 | ~v_148;
assign x_418 = ~v_145 | ~v_146;
assign x_419 = v_148 | ~v_145 | ~v_31;
assign x_420 = v_31 | v_149 | ~v_145;
assign x_421 = v_146 | v_338 | v_147;
assign x_422 = v_146 | v_27 | v_147;
assign x_423 = v_146 | v_277 | ~v_338 | ~v_27;
assign x_424 = v_338 | ~v_146 | ~v_147;
assign x_425 = v_27 | ~v_146 | ~v_147;
assign x_426 = ~v_146 | ~v_277 | ~v_338 | ~v_27;
assign x_427 = v_148 | v_218 | v_281 | ~v_50;
assign x_428 = v_148 | v_218 | v_259 | ~v_281;
assign x_429 = ~v_148 | ~v_218;
assign x_430 = ~v_148 | ~v_259 | ~v_281;
assign x_431 = v_281 | v_50 | ~v_148;
assign x_432 = v_154 | v_270 | ~v_268;
assign x_433 = v_154 | v_268 | v_269 | ~v_270;
assign x_434 = v_154 | v_269 | v_270 | ~v_271;
assign x_435 = v_268 | ~v_154 | ~v_269;
assign x_436 = ~v_154 | ~v_268 | ~v_270;
assign x_437 = v_268 | v_270 | v_271 | ~v_154;
assign x_438 = v_156 | v_157 | ~v_158;
assign x_439 = v_156 | v_270 | ~v_271 | ~v_158;
assign x_440 = v_158 | ~v_156;
assign x_441 = ~v_156 | ~v_270 | ~v_157;
assign x_442 = v_271 | ~v_156 | ~v_157;
assign x_443 = v_166 | v_225 | v_288 | v_167 | v_168;
assign x_444 = v_166 | v_167 | v_168 | ~v_225 | ~v_288;
assign x_445 = ~v_166 | ~v_167;
assign x_446 = v_288 | ~v_166 | ~v_225;
assign x_447 = ~v_166 | ~v_168;
assign x_448 = v_225 | ~v_166 | ~v_288;
assign x_449 = v_169 | v_232 | v_295 | ~v_231 | ~v_294;
assign x_450 = v_169 | v_231 | v_294 | ~v_232 | ~v_295;
assign x_451 = v_169 | v_231 | v_232 | v_294 | v_295;
assign x_452 = v_169 | ~v_231 | ~v_232 | ~v_294 | ~v_295;
assign x_453 = v_294 | ~v_169 | ~v_231;
assign x_454 = v_231 | ~v_169 | ~v_294;
assign x_455 = v_232 | ~v_169 | ~v_295;
assign x_456 = v_295 | ~v_169 | ~v_232;
assign x_457 = v_170 | v_240 | v_303 | v_171 | v_172;
assign x_458 = v_170 | v_171 | v_172 | ~v_240 | ~v_303;
assign x_459 = ~v_170 | ~v_171;
assign x_460 = v_303 | ~v_170 | ~v_240;
assign x_461 = ~v_170 | ~v_172;
assign x_462 = v_240 | ~v_170 | ~v_303;
assign x_463 = v_173 | v_260 | v_323 | v_174 | v_175;
assign x_464 = v_173 | v_174 | v_175 | ~v_260 | ~v_323;
assign x_465 = ~v_173 | ~v_174;
assign x_466 = v_323 | ~v_173 | ~v_260;
assign x_467 = ~v_173 | ~v_175;
assign x_468 = v_260 | ~v_173 | ~v_323;
assign x_469 = v_177 | v_317 | v_178 | ~v_179;
assign x_470 = v_177 | v_178 | ~v_254 | ~v_179;
assign x_471 = v_179 | ~v_177;
assign x_472 = ~v_177 | ~v_178;
assign x_473 = v_254 | ~v_177 | ~v_317;
assign x_474 = v_179 | v_180 | ~v_297;
assign x_475 = v_179 | v_234 | v_180;
assign x_476 = ~v_179 | ~v_180;
assign x_477 = v_297 | ~v_179 | ~v_234;
assign x_478 = v_181 | v_263 | v_326 | v_182 | v_183;
assign x_479 = v_181 | v_182 | v_183 | ~v_263 | ~v_326;
assign x_480 = ~v_181 | ~v_182;
assign x_481 = v_326 | ~v_181 | ~v_263;
assign x_482 = ~v_181 | ~v_183;
assign x_483 = v_263 | ~v_181 | ~v_326;
assign x_484 = v_184 | v_250 | v_313 | v_185 | v_186;
assign x_485 = v_184 | v_185 | v_186 | ~v_250 | ~v_313;
assign x_486 = ~v_184 | ~v_185;
assign x_487 = v_313 | ~v_184 | ~v_250;
assign x_488 = ~v_184 | ~v_186;
assign x_489 = v_250 | ~v_184 | ~v_313;
assign x_490 = v_187 | v_246 | v_309 | v_188 | v_189;
assign x_491 = v_187 | v_188 | v_189 | ~v_246 | ~v_309;
assign x_492 = ~v_187 | ~v_188;
assign x_493 = v_309 | ~v_187 | ~v_246;
assign x_494 = ~v_187 | ~v_189;
assign x_495 = v_246 | ~v_187 | ~v_309;
assign x_496 = v_191 | v_271 | v_334 | ~v_270 | ~v_333;
assign x_497 = v_191 | v_270 | v_333 | ~v_271 | ~v_334;
assign x_498 = v_191 | v_270 | v_271 | v_333 | v_334;
assign x_499 = v_191 | ~v_270 | ~v_271 | ~v_333 | ~v_334;
assign x_500 = v_333 | ~v_191 | ~v_270;
assign x_501 = v_270 | ~v_191 | ~v_333;
assign x_502 = v_271 | ~v_191 | ~v_334;
assign x_503 = v_334 | ~v_191 | ~v_271;
assign x_504 = v_192 | ~v_328 | ~v_193;
assign x_505 = v_192 | v_265 | ~v_193;
assign x_506 = v_193 | ~v_192;
assign x_507 = v_328 | ~v_192 | ~v_265;
assign x_508 = v_193 | v_226 | v_251;
assign x_509 = v_193 | ~v_289 | ~v_314;
assign x_510 = v_193 | v_226 | ~v_314;
assign x_511 = v_193 | v_251 | ~v_289;
assign x_512 = v_289 | ~v_193 | ~v_226;
assign x_513 = v_314 | ~v_193 | ~v_251;
assign x_514 = v_198 | v_223 | v_286 | ~v_216 | ~v_279;
assign x_515 = v_198 | v_216 | v_279 | ~v_223 | ~v_286;
assign x_516 = v_198 | v_216 | v_223 | v_279 | v_286;
assign x_517 = v_198 | ~v_216 | ~v_223 | ~v_279 | ~v_286;
assign x_518 = v_279 | ~v_198 | ~v_216;
assign x_519 = v_216 | ~v_198 | ~v_279;
assign x_520 = v_223 | ~v_198 | ~v_286;
assign x_521 = v_286 | ~v_198 | ~v_223;
assign x_522 = v_199 | v_219 | v_282 | ~v_76 | ~v_200;
assign x_523 = v_199 | ~v_219 | ~v_282 | ~v_76 | ~v_200;
assign x_524 = v_200 | ~v_199;
assign x_525 = v_282 | ~v_199 | ~v_219;
assign x_526 = v_76 | ~v_199;
assign x_527 = v_219 | ~v_199 | ~v_282;
assign x_528 = v_200 | ~v_268 | ~v_331 | ~v_201;
assign x_529 = v_200 | v_268 | v_331 | ~v_201;
assign x_530 = v_201 | ~v_200;
assign x_531 = v_331 | ~v_200 | ~v_268;
assign x_532 = v_268 | ~v_200 | ~v_331;
assign x_533 = v_202 | v_252 | v_315 | ~v_233 | ~v_296;
assign x_534 = v_202 | v_233 | v_296 | ~v_252 | ~v_315;
assign x_535 = v_202 | v_233 | v_252 | v_296 | v_315;
assign x_536 = v_202 | ~v_233 | ~v_252 | ~v_296 | ~v_315;
assign x_537 = v_296 | ~v_202 | ~v_233;
assign x_538 = v_233 | ~v_202 | ~v_296;
assign x_539 = v_252 | ~v_202 | ~v_315;
assign x_540 = v_315 | ~v_202 | ~v_252;
assign x_541 = v_207 | v_249 | v_312 | v_209 | ~v_208;
assign x_542 = v_207 | v_209 | ~v_249 | ~v_312 | ~v_208;
assign x_543 = ~v_207 | ~v_209;
assign x_544 = v_312 | ~v_207 | ~v_249;
assign x_545 = v_208 | ~v_207;
assign x_546 = v_249 | ~v_207 | ~v_312;
assign x_547 = v_208 | v_257 | v_320 | ~v_228 | ~v_291;
assign x_548 = v_208 | v_228 | v_291 | ~v_257 | ~v_320;
assign x_549 = v_208 | v_228 | v_257 | v_291 | v_320;
assign x_550 = v_208 | ~v_228 | ~v_257 | ~v_291 | ~v_320;
assign x_551 = v_291 | ~v_208 | ~v_228;
assign x_552 = v_228 | ~v_208 | ~v_291;
assign x_553 = v_257 | ~v_208 | ~v_320;
assign x_554 = v_320 | ~v_208 | ~v_257;
assign x_555 = v_210 | v_287 | ~v_265;
assign x_556 = v_210 | v_328 | ~v_224;
assign x_557 = v_210 | ~v_224 | ~v_265;
assign x_558 = v_210 | v_287 | v_328;
assign x_559 = v_265 | ~v_210 | ~v_328;
assign x_560 = v_224 | ~v_210 | ~v_287;
assign x_561 = v_211 | v_237 | v_261;
assign x_562 = v_211 | ~v_300 | ~v_324;
assign x_563 = v_211 | v_237 | ~v_324;
assign x_564 = v_211 | v_261 | ~v_300;
assign x_565 = v_300 | ~v_211 | ~v_237;
assign x_566 = v_324 | ~v_211 | ~v_261;
assign x_567 = v_212 | ~v_251 | ~v_343 | ~v_213;
assign x_568 = v_212 | v_314 | ~v_343 | ~v_213;
assign x_569 = v_213 | ~v_212;
assign x_570 = v_343 | ~v_212;
assign x_571 = v_251 | ~v_212 | ~v_314;
assign x_572 = v_213 | ~v_237 | ~v_287;
assign x_573 = v_213 | v_224 | v_300;
assign x_574 = v_213 | v_224 | ~v_237;
assign x_575 = v_213 | v_300 | ~v_287;
assign x_576 = v_287 | ~v_213 | ~v_224;
assign x_577 = v_237 | ~v_213 | ~v_300;
assign x_578 = x_1 & x_2;
assign x_579 = x_3 & x_4;
assign x_580 = x_578 & x_579;
assign x_581 = x_5 & x_6;
assign x_582 = x_8 & x_9;
assign x_583 = x_7 & x_582;
assign x_584 = x_581 & x_583;
assign x_585 = x_580 & x_584;
assign x_586 = x_10 & x_11;
assign x_587 = x_12 & x_13;
assign x_588 = x_586 & x_587;
assign x_589 = x_14 & x_15;
assign x_590 = x_17 & x_18;
assign x_591 = x_16 & x_590;
assign x_592 = x_589 & x_591;
assign x_593 = x_588 & x_592;
assign x_594 = x_585 & x_593;
assign x_595 = x_19 & x_20;
assign x_596 = x_21 & x_22;
assign x_597 = x_595 & x_596;
assign x_598 = x_23 & x_24;
assign x_599 = x_26 & x_27;
assign x_600 = x_25 & x_599;
assign x_601 = x_598 & x_600;
assign x_602 = x_597 & x_601;
assign x_603 = x_28 & x_29;
assign x_604 = x_30 & x_31;
assign x_605 = x_603 & x_604;
assign x_606 = x_32 & x_33;
assign x_607 = x_35 & x_36;
assign x_608 = x_34 & x_607;
assign x_609 = x_606 & x_608;
assign x_610 = x_605 & x_609;
assign x_611 = x_602 & x_610;
assign x_612 = x_594 & x_611;
assign x_613 = x_37 & x_38;
assign x_614 = x_39 & x_40;
assign x_615 = x_613 & x_614;
assign x_616 = x_41 & x_42;
assign x_617 = x_44 & x_45;
assign x_618 = x_43 & x_617;
assign x_619 = x_616 & x_618;
assign x_620 = x_615 & x_619;
assign x_621 = x_46 & x_47;
assign x_622 = x_48 & x_49;
assign x_623 = x_621 & x_622;
assign x_624 = x_50 & x_51;
assign x_625 = x_53 & x_54;
assign x_626 = x_52 & x_625;
assign x_627 = x_624 & x_626;
assign x_628 = x_623 & x_627;
assign x_629 = x_620 & x_628;
assign x_630 = x_55 & x_56;
assign x_631 = x_57 & x_58;
assign x_632 = x_630 & x_631;
assign x_633 = x_59 & x_60;
assign x_634 = x_62 & x_63;
assign x_635 = x_61 & x_634;
assign x_636 = x_633 & x_635;
assign x_637 = x_632 & x_636;
assign x_638 = x_64 & x_65;
assign x_639 = x_66 & x_67;
assign x_640 = x_638 & x_639;
assign x_641 = x_68 & x_69;
assign x_642 = x_71 & x_72;
assign x_643 = x_70 & x_642;
assign x_644 = x_641 & x_643;
assign x_645 = x_640 & x_644;
assign x_646 = x_637 & x_645;
assign x_647 = x_629 & x_646;
assign x_648 = x_612 & x_647;
assign x_649 = x_73 & x_74;
assign x_650 = x_75 & x_76;
assign x_651 = x_649 & x_650;
assign x_652 = x_77 & x_78;
assign x_653 = x_80 & x_81;
assign x_654 = x_79 & x_653;
assign x_655 = x_652 & x_654;
assign x_656 = x_651 & x_655;
assign x_657 = x_82 & x_83;
assign x_658 = x_84 & x_85;
assign x_659 = x_657 & x_658;
assign x_660 = x_86 & x_87;
assign x_661 = x_89 & x_90;
assign x_662 = x_88 & x_661;
assign x_663 = x_660 & x_662;
assign x_664 = x_659 & x_663;
assign x_665 = x_656 & x_664;
assign x_666 = x_91 & x_92;
assign x_667 = x_93 & x_94;
assign x_668 = x_666 & x_667;
assign x_669 = x_95 & x_96;
assign x_670 = x_98 & x_99;
assign x_671 = x_97 & x_670;
assign x_672 = x_669 & x_671;
assign x_673 = x_668 & x_672;
assign x_674 = x_100 & x_101;
assign x_675 = x_102 & x_103;
assign x_676 = x_674 & x_675;
assign x_677 = x_104 & x_105;
assign x_678 = x_107 & x_108;
assign x_679 = x_106 & x_678;
assign x_680 = x_677 & x_679;
assign x_681 = x_676 & x_680;
assign x_682 = x_673 & x_681;
assign x_683 = x_665 & x_682;
assign x_684 = x_109 & x_110;
assign x_685 = x_111 & x_112;
assign x_686 = x_684 & x_685;
assign x_687 = x_113 & x_114;
assign x_688 = x_116 & x_117;
assign x_689 = x_115 & x_688;
assign x_690 = x_687 & x_689;
assign x_691 = x_686 & x_690;
assign x_692 = x_118 & x_119;
assign x_693 = x_120 & x_121;
assign x_694 = x_692 & x_693;
assign x_695 = x_122 & x_123;
assign x_696 = x_125 & x_126;
assign x_697 = x_124 & x_696;
assign x_698 = x_695 & x_697;
assign x_699 = x_694 & x_698;
assign x_700 = x_691 & x_699;
assign x_701 = x_127 & x_128;
assign x_702 = x_129 & x_130;
assign x_703 = x_701 & x_702;
assign x_704 = x_131 & x_132;
assign x_705 = x_134 & x_135;
assign x_706 = x_133 & x_705;
assign x_707 = x_704 & x_706;
assign x_708 = x_703 & x_707;
assign x_709 = x_136 & x_137;
assign x_710 = x_138 & x_139;
assign x_711 = x_709 & x_710;
assign x_712 = x_140 & x_141;
assign x_713 = x_143 & x_144;
assign x_714 = x_142 & x_713;
assign x_715 = x_712 & x_714;
assign x_716 = x_711 & x_715;
assign x_717 = x_708 & x_716;
assign x_718 = x_700 & x_717;
assign x_719 = x_683 & x_718;
assign x_720 = x_648 & x_719;
assign x_721 = x_145 & x_146;
assign x_722 = x_147 & x_148;
assign x_723 = x_721 & x_722;
assign x_724 = x_149 & x_150;
assign x_725 = x_152 & x_153;
assign x_726 = x_151 & x_725;
assign x_727 = x_724 & x_726;
assign x_728 = x_723 & x_727;
assign x_729 = x_154 & x_155;
assign x_730 = x_156 & x_157;
assign x_731 = x_729 & x_730;
assign x_732 = x_158 & x_159;
assign x_733 = x_161 & x_162;
assign x_734 = x_160 & x_733;
assign x_735 = x_732 & x_734;
assign x_736 = x_731 & x_735;
assign x_737 = x_728 & x_736;
assign x_738 = x_163 & x_164;
assign x_739 = x_165 & x_166;
assign x_740 = x_738 & x_739;
assign x_741 = x_167 & x_168;
assign x_742 = x_170 & x_171;
assign x_743 = x_169 & x_742;
assign x_744 = x_741 & x_743;
assign x_745 = x_740 & x_744;
assign x_746 = x_172 & x_173;
assign x_747 = x_174 & x_175;
assign x_748 = x_746 & x_747;
assign x_749 = x_176 & x_177;
assign x_750 = x_179 & x_180;
assign x_751 = x_178 & x_750;
assign x_752 = x_749 & x_751;
assign x_753 = x_748 & x_752;
assign x_754 = x_745 & x_753;
assign x_755 = x_737 & x_754;
assign x_756 = x_181 & x_182;
assign x_757 = x_183 & x_184;
assign x_758 = x_756 & x_757;
assign x_759 = x_185 & x_186;
assign x_760 = x_188 & x_189;
assign x_761 = x_187 & x_760;
assign x_762 = x_759 & x_761;
assign x_763 = x_758 & x_762;
assign x_764 = x_190 & x_191;
assign x_765 = x_192 & x_193;
assign x_766 = x_764 & x_765;
assign x_767 = x_194 & x_195;
assign x_768 = x_197 & x_198;
assign x_769 = x_196 & x_768;
assign x_770 = x_767 & x_769;
assign x_771 = x_766 & x_770;
assign x_772 = x_763 & x_771;
assign x_773 = x_199 & x_200;
assign x_774 = x_201 & x_202;
assign x_775 = x_773 & x_774;
assign x_776 = x_203 & x_204;
assign x_777 = x_206 & x_207;
assign x_778 = x_205 & x_777;
assign x_779 = x_776 & x_778;
assign x_780 = x_775 & x_779;
assign x_781 = x_208 & x_209;
assign x_782 = x_210 & x_211;
assign x_783 = x_781 & x_782;
assign x_784 = x_212 & x_213;
assign x_785 = x_215 & x_216;
assign x_786 = x_214 & x_785;
assign x_787 = x_784 & x_786;
assign x_788 = x_783 & x_787;
assign x_789 = x_780 & x_788;
assign x_790 = x_772 & x_789;
assign x_791 = x_755 & x_790;
assign x_792 = x_217 & x_218;
assign x_793 = x_219 & x_220;
assign x_794 = x_792 & x_793;
assign x_795 = x_221 & x_222;
assign x_796 = x_224 & x_225;
assign x_797 = x_223 & x_796;
assign x_798 = x_795 & x_797;
assign x_799 = x_794 & x_798;
assign x_800 = x_226 & x_227;
assign x_801 = x_228 & x_229;
assign x_802 = x_800 & x_801;
assign x_803 = x_230 & x_231;
assign x_804 = x_233 & x_234;
assign x_805 = x_232 & x_804;
assign x_806 = x_803 & x_805;
assign x_807 = x_802 & x_806;
assign x_808 = x_799 & x_807;
assign x_809 = x_235 & x_236;
assign x_810 = x_237 & x_238;
assign x_811 = x_809 & x_810;
assign x_812 = x_239 & x_240;
assign x_813 = x_242 & x_243;
assign x_814 = x_241 & x_813;
assign x_815 = x_812 & x_814;
assign x_816 = x_811 & x_815;
assign x_817 = x_244 & x_245;
assign x_818 = x_246 & x_247;
assign x_819 = x_817 & x_818;
assign x_820 = x_248 & x_249;
assign x_821 = x_251 & x_252;
assign x_822 = x_250 & x_821;
assign x_823 = x_820 & x_822;
assign x_824 = x_819 & x_823;
assign x_825 = x_816 & x_824;
assign x_826 = x_808 & x_825;
assign x_827 = x_253 & x_254;
assign x_828 = x_255 & x_256;
assign x_829 = x_827 & x_828;
assign x_830 = x_257 & x_258;
assign x_831 = x_260 & x_261;
assign x_832 = x_259 & x_831;
assign x_833 = x_830 & x_832;
assign x_834 = x_829 & x_833;
assign x_835 = x_262 & x_263;
assign x_836 = x_264 & x_265;
assign x_837 = x_835 & x_836;
assign x_838 = x_266 & x_267;
assign x_839 = x_269 & x_270;
assign x_840 = x_268 & x_839;
assign x_841 = x_838 & x_840;
assign x_842 = x_837 & x_841;
assign x_843 = x_834 & x_842;
assign x_844 = x_271 & x_272;
assign x_845 = x_273 & x_274;
assign x_846 = x_844 & x_845;
assign x_847 = x_275 & x_276;
assign x_848 = x_278 & x_279;
assign x_849 = x_277 & x_848;
assign x_850 = x_847 & x_849;
assign x_851 = x_846 & x_850;
assign x_852 = x_280 & x_281;
assign x_853 = x_282 & x_283;
assign x_854 = x_852 & x_853;
assign x_855 = x_284 & x_285;
assign x_856 = x_287 & x_288;
assign x_857 = x_286 & x_856;
assign x_858 = x_855 & x_857;
assign x_859 = x_854 & x_858;
assign x_860 = x_851 & x_859;
assign x_861 = x_843 & x_860;
assign x_862 = x_826 & x_861;
assign x_863 = x_791 & x_862;
assign x_864 = x_720 & x_863;
assign x_865 = x_289 & x_290;
assign x_866 = x_291 & x_292;
assign x_867 = x_865 & x_866;
assign x_868 = x_293 & x_294;
assign x_869 = x_296 & x_297;
assign x_870 = x_295 & x_869;
assign x_871 = x_868 & x_870;
assign x_872 = x_867 & x_871;
assign x_873 = x_298 & x_299;
assign x_874 = x_300 & x_301;
assign x_875 = x_873 & x_874;
assign x_876 = x_302 & x_303;
assign x_877 = x_305 & x_306;
assign x_878 = x_304 & x_877;
assign x_879 = x_876 & x_878;
assign x_880 = x_875 & x_879;
assign x_881 = x_872 & x_880;
assign x_882 = x_307 & x_308;
assign x_883 = x_309 & x_310;
assign x_884 = x_882 & x_883;
assign x_885 = x_311 & x_312;
assign x_886 = x_314 & x_315;
assign x_887 = x_313 & x_886;
assign x_888 = x_885 & x_887;
assign x_889 = x_884 & x_888;
assign x_890 = x_316 & x_317;
assign x_891 = x_318 & x_319;
assign x_892 = x_890 & x_891;
assign x_893 = x_320 & x_321;
assign x_894 = x_323 & x_324;
assign x_895 = x_322 & x_894;
assign x_896 = x_893 & x_895;
assign x_897 = x_892 & x_896;
assign x_898 = x_889 & x_897;
assign x_899 = x_881 & x_898;
assign x_900 = x_325 & x_326;
assign x_901 = x_327 & x_328;
assign x_902 = x_900 & x_901;
assign x_903 = x_329 & x_330;
assign x_904 = x_332 & x_333;
assign x_905 = x_331 & x_904;
assign x_906 = x_903 & x_905;
assign x_907 = x_902 & x_906;
assign x_908 = x_334 & x_335;
assign x_909 = x_336 & x_337;
assign x_910 = x_908 & x_909;
assign x_911 = x_338 & x_339;
assign x_912 = x_341 & x_342;
assign x_913 = x_340 & x_912;
assign x_914 = x_911 & x_913;
assign x_915 = x_910 & x_914;
assign x_916 = x_907 & x_915;
assign x_917 = x_343 & x_344;
assign x_918 = x_345 & x_346;
assign x_919 = x_917 & x_918;
assign x_920 = x_347 & x_348;
assign x_921 = x_350 & x_351;
assign x_922 = x_349 & x_921;
assign x_923 = x_920 & x_922;
assign x_924 = x_919 & x_923;
assign x_925 = x_352 & x_353;
assign x_926 = x_354 & x_355;
assign x_927 = x_925 & x_926;
assign x_928 = x_356 & x_357;
assign x_929 = x_359 & x_360;
assign x_930 = x_358 & x_929;
assign x_931 = x_928 & x_930;
assign x_932 = x_927 & x_931;
assign x_933 = x_924 & x_932;
assign x_934 = x_916 & x_933;
assign x_935 = x_899 & x_934;
assign x_936 = x_361 & x_362;
assign x_937 = x_363 & x_364;
assign x_938 = x_936 & x_937;
assign x_939 = x_365 & x_366;
assign x_940 = x_368 & x_369;
assign x_941 = x_367 & x_940;
assign x_942 = x_939 & x_941;
assign x_943 = x_938 & x_942;
assign x_944 = x_370 & x_371;
assign x_945 = x_372 & x_373;
assign x_946 = x_944 & x_945;
assign x_947 = x_374 & x_375;
assign x_948 = x_377 & x_378;
assign x_949 = x_376 & x_948;
assign x_950 = x_947 & x_949;
assign x_951 = x_946 & x_950;
assign x_952 = x_943 & x_951;
assign x_953 = x_379 & x_380;
assign x_954 = x_381 & x_382;
assign x_955 = x_953 & x_954;
assign x_956 = x_383 & x_384;
assign x_957 = x_386 & x_387;
assign x_958 = x_385 & x_957;
assign x_959 = x_956 & x_958;
assign x_960 = x_955 & x_959;
assign x_961 = x_388 & x_389;
assign x_962 = x_390 & x_391;
assign x_963 = x_961 & x_962;
assign x_964 = x_392 & x_393;
assign x_965 = x_395 & x_396;
assign x_966 = x_394 & x_965;
assign x_967 = x_964 & x_966;
assign x_968 = x_963 & x_967;
assign x_969 = x_960 & x_968;
assign x_970 = x_952 & x_969;
assign x_971 = x_397 & x_398;
assign x_972 = x_399 & x_400;
assign x_973 = x_971 & x_972;
assign x_974 = x_401 & x_402;
assign x_975 = x_404 & x_405;
assign x_976 = x_403 & x_975;
assign x_977 = x_974 & x_976;
assign x_978 = x_973 & x_977;
assign x_979 = x_406 & x_407;
assign x_980 = x_408 & x_409;
assign x_981 = x_979 & x_980;
assign x_982 = x_410 & x_411;
assign x_983 = x_413 & x_414;
assign x_984 = x_412 & x_983;
assign x_985 = x_982 & x_984;
assign x_986 = x_981 & x_985;
assign x_987 = x_978 & x_986;
assign x_988 = x_415 & x_416;
assign x_989 = x_417 & x_418;
assign x_990 = x_988 & x_989;
assign x_991 = x_419 & x_420;
assign x_992 = x_422 & x_423;
assign x_993 = x_421 & x_992;
assign x_994 = x_991 & x_993;
assign x_995 = x_990 & x_994;
assign x_996 = x_424 & x_425;
assign x_997 = x_426 & x_427;
assign x_998 = x_996 & x_997;
assign x_999 = x_428 & x_429;
assign x_1000 = x_431 & x_432;
assign x_1001 = x_430 & x_1000;
assign x_1002 = x_999 & x_1001;
assign x_1003 = x_998 & x_1002;
assign x_1004 = x_995 & x_1003;
assign x_1005 = x_987 & x_1004;
assign x_1006 = x_970 & x_1005;
assign x_1007 = x_935 & x_1006;
assign x_1008 = x_433 & x_434;
assign x_1009 = x_435 & x_436;
assign x_1010 = x_1008 & x_1009;
assign x_1011 = x_437 & x_438;
assign x_1012 = x_440 & x_441;
assign x_1013 = x_439 & x_1012;
assign x_1014 = x_1011 & x_1013;
assign x_1015 = x_1010 & x_1014;
assign x_1016 = x_442 & x_443;
assign x_1017 = x_444 & x_445;
assign x_1018 = x_1016 & x_1017;
assign x_1019 = x_446 & x_447;
assign x_1020 = x_449 & x_450;
assign x_1021 = x_448 & x_1020;
assign x_1022 = x_1019 & x_1021;
assign x_1023 = x_1018 & x_1022;
assign x_1024 = x_1015 & x_1023;
assign x_1025 = x_451 & x_452;
assign x_1026 = x_453 & x_454;
assign x_1027 = x_1025 & x_1026;
assign x_1028 = x_455 & x_456;
assign x_1029 = x_458 & x_459;
assign x_1030 = x_457 & x_1029;
assign x_1031 = x_1028 & x_1030;
assign x_1032 = x_1027 & x_1031;
assign x_1033 = x_460 & x_461;
assign x_1034 = x_462 & x_463;
assign x_1035 = x_1033 & x_1034;
assign x_1036 = x_464 & x_465;
assign x_1037 = x_467 & x_468;
assign x_1038 = x_466 & x_1037;
assign x_1039 = x_1036 & x_1038;
assign x_1040 = x_1035 & x_1039;
assign x_1041 = x_1032 & x_1040;
assign x_1042 = x_1024 & x_1041;
assign x_1043 = x_469 & x_470;
assign x_1044 = x_471 & x_472;
assign x_1045 = x_1043 & x_1044;
assign x_1046 = x_473 & x_474;
assign x_1047 = x_476 & x_477;
assign x_1048 = x_475 & x_1047;
assign x_1049 = x_1046 & x_1048;
assign x_1050 = x_1045 & x_1049;
assign x_1051 = x_478 & x_479;
assign x_1052 = x_480 & x_481;
assign x_1053 = x_1051 & x_1052;
assign x_1054 = x_482 & x_483;
assign x_1055 = x_485 & x_486;
assign x_1056 = x_484 & x_1055;
assign x_1057 = x_1054 & x_1056;
assign x_1058 = x_1053 & x_1057;
assign x_1059 = x_1050 & x_1058;
assign x_1060 = x_487 & x_488;
assign x_1061 = x_489 & x_490;
assign x_1062 = x_1060 & x_1061;
assign x_1063 = x_491 & x_492;
assign x_1064 = x_494 & x_495;
assign x_1065 = x_493 & x_1064;
assign x_1066 = x_1063 & x_1065;
assign x_1067 = x_1062 & x_1066;
assign x_1068 = x_496 & x_497;
assign x_1069 = x_498 & x_499;
assign x_1070 = x_1068 & x_1069;
assign x_1071 = x_500 & x_501;
assign x_1072 = x_503 & x_504;
assign x_1073 = x_502 & x_1072;
assign x_1074 = x_1071 & x_1073;
assign x_1075 = x_1070 & x_1074;
assign x_1076 = x_1067 & x_1075;
assign x_1077 = x_1059 & x_1076;
assign x_1078 = x_1042 & x_1077;
assign x_1079 = x_505 & x_506;
assign x_1080 = x_507 & x_508;
assign x_1081 = x_1079 & x_1080;
assign x_1082 = x_509 & x_510;
assign x_1083 = x_512 & x_513;
assign x_1084 = x_511 & x_1083;
assign x_1085 = x_1082 & x_1084;
assign x_1086 = x_1081 & x_1085;
assign x_1087 = x_514 & x_515;
assign x_1088 = x_516 & x_517;
assign x_1089 = x_1087 & x_1088;
assign x_1090 = x_518 & x_519;
assign x_1091 = x_521 & x_522;
assign x_1092 = x_520 & x_1091;
assign x_1093 = x_1090 & x_1092;
assign x_1094 = x_1089 & x_1093;
assign x_1095 = x_1086 & x_1094;
assign x_1096 = x_523 & x_524;
assign x_1097 = x_525 & x_526;
assign x_1098 = x_1096 & x_1097;
assign x_1099 = x_527 & x_528;
assign x_1100 = x_530 & x_531;
assign x_1101 = x_529 & x_1100;
assign x_1102 = x_1099 & x_1101;
assign x_1103 = x_1098 & x_1102;
assign x_1104 = x_532 & x_533;
assign x_1105 = x_534 & x_535;
assign x_1106 = x_1104 & x_1105;
assign x_1107 = x_536 & x_537;
assign x_1108 = x_539 & x_540;
assign x_1109 = x_538 & x_1108;
assign x_1110 = x_1107 & x_1109;
assign x_1111 = x_1106 & x_1110;
assign x_1112 = x_1103 & x_1111;
assign x_1113 = x_1095 & x_1112;
assign x_1114 = x_541 & x_542;
assign x_1115 = x_543 & x_544;
assign x_1116 = x_1114 & x_1115;
assign x_1117 = x_545 & x_546;
assign x_1118 = x_548 & x_549;
assign x_1119 = x_547 & x_1118;
assign x_1120 = x_1117 & x_1119;
assign x_1121 = x_1116 & x_1120;
assign x_1122 = x_550 & x_551;
assign x_1123 = x_552 & x_553;
assign x_1124 = x_1122 & x_1123;
assign x_1125 = x_554 & x_555;
assign x_1126 = x_557 & x_558;
assign x_1127 = x_556 & x_1126;
assign x_1128 = x_1125 & x_1127;
assign x_1129 = x_1124 & x_1128;
assign x_1130 = x_1121 & x_1129;
assign x_1131 = x_559 & x_560;
assign x_1132 = x_561 & x_562;
assign x_1133 = x_1131 & x_1132;
assign x_1134 = x_563 & x_564;
assign x_1135 = x_566 & x_567;
assign x_1136 = x_565 & x_1135;
assign x_1137 = x_1134 & x_1136;
assign x_1138 = x_1133 & x_1137;
assign x_1139 = x_568 & x_569;
assign x_1140 = x_571 & x_572;
assign x_1141 = x_570 & x_1140;
assign x_1142 = x_1139 & x_1141;
assign x_1143 = x_573 & x_574;
assign x_1144 = x_576 & x_577;
assign x_1145 = x_575 & x_1144;
assign x_1146 = x_1143 & x_1145;
assign x_1147 = x_1142 & x_1146;
assign x_1148 = x_1138 & x_1147;
assign x_1149 = x_1130 & x_1148;
assign x_1150 = x_1113 & x_1149;
assign x_1151 = x_1078 & x_1150;
assign x_1152 = x_1007 & x_1151;
assign x_1153 = x_864 & x_1152;
assign o_1 = x_1153;
endmodule
