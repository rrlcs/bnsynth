// Benchmark "SKOLEMFORMULA" written by ABC on Fri May 20 19:43:02 2022

module SKOLEMFORMULA ( 
    i0,
    i1, i2, i3  );
  input  i0;
  output i1, i2, i3;
  assign i1 = 1'b1;
  assign i3 = 1'b1;
  assign i2 = ~i0;
endmodule


