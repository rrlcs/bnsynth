// Benchmark "SKOLEMFORMULA" written by ABC on Fri May 20 19:19:16 2022

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7, i8, i9,
    i10, i11, i12, i13, i14, i15, i16, i17, i18, i19  );
  input  i0, i1, i2, i3, i4, i5, i6, i7, i8, i9;
  output i10, i11, i12, i13, i14, i15, i16, i17, i18, i19;
  assign i10 = i0;
  assign i11 = i1;
  assign i12 = i2;
  assign i13 = i3;
  assign i14 = i4;
  assign i15 = i5;
  assign i16 = i6;
  assign i17 = i7;
  assign i18 = i8;
  assign i19 = i9;
endmodule


