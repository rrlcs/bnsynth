module formula(v_1,v_2,v_3,v_4,v_5,v_6,v_7,v_8,v_25,v_26,v_27,v_28,v_29,v_30,v_31,v_32,v_33,v_34,v_35,v_36,v_37,v_38,v_39,v_40,v_41,v_42,v_43,v_44,v_45,v_46,v_47,v_48,v_49,v_50,v_51,v_52,v_53,v_54,v_55,v_56,v_57,v_58,v_59,v_60,v_61,v_62,v_63,v_64,v_65,v_66,v_67,v_68,v_69,v_70,v_71,v_72,v_73,v_74,v_75,v_76,v_77,v_78,v_79,v_80,v_81,v_82,v_83,v_84,v_85,v_86,v_87,v_88,v_89,v_90,v_9,v_10,v_11,v_12,v_13,v_14,v_15,v_16,v_17,v_18,v_19,v_20,v_21,v_22,v_23,v_24,v_91,v_92,v_93,v_94,v_95,v_96,v_97,v_98,v_99,v_100,v_101,v_102,v_103,v_104,v_105,v_106,v_107,v_108,v_109,v_110,v_111,v_112,v_113,v_114,v_115,v_116,v_117,v_118,v_119,v_120,v_121,v_122,v_123,v_124,v_125,v_126,v_127,v_128,v_129,v_130,v_131,v_132,v_133,v_134,v_135,v_136,v_137,v_138,v_139,v_140,v_141,v_142,v_143,v_144,v_145,v_146,v_147,v_148,v_149,v_150,v_151,v_152,v_153,v_154,v_155,v_156,v_157,v_158,v_159,v_160,v_161,v_162,v_163,v_164,v_165,v_166,v_167,v_168,v_169,v_170,v_171,v_172,v_173,v_174,v_175,v_176,v_177,v_178,v_179,v_180,v_181,v_182,v_183,v_184,v_185,v_186,v_187,v_188,v_189,v_190,v_191,v_192,v_193,v_194,v_195,v_196,v_197,v_198,v_199,v_200,v_201,v_202,v_203,v_204,v_205,v_206,v_207,v_208,v_209,v_210,v_211,v_212,v_213,v_214,v_215,v_216,v_217,v_218,v_219,v_220,v_221,v_222,v_223,v_224,v_225,v_226,v_227,v_228,v_229,v_230,v_231,v_232,v_233,v_234,v_235,v_236,v_237,v_238,v_239,v_240,v_241,v_242,v_243,v_244,v_245,v_246,v_247,v_248,v_249,v_250,v_251,v_252,v_253,v_254,v_255,v_256,v_257,v_258,v_259,v_260,v_261,v_262,v_263,v_264,v_265,v_266,v_267,v_268,v_269,v_270,v_271,v_272,v_273,v_274,v_275,v_276,v_277,v_278,v_279,v_280,v_281,v_282,v_283,v_284,v_285,v_286,v_287,v_288,v_289,v_290,v_291,v_292,v_293,v_294,v_295,v_296,v_297,v_298,v_299,v_300,v_301,v_302,v_303,v_304,v_305,v_306,v_307,v_308,v_309,v_310,v_311,v_312,v_313,v_314,v_315,v_316,v_317,v_318,v_319,v_320,v_321,v_322,v_323,v_324,v_325,v_326,v_327,v_328,v_329,v_330,v_331,v_332,v_333,v_334,v_335,v_336,v_337,v_338,v_339,v_340,v_341,v_342,v_343,v_344,v_345,v_346,v_347,v_348,v_349,v_350,v_351,v_352,v_353,v_354,v_355,v_356,v_357,v_358,v_359,v_360,v_361,v_362,v_363,v_364,v_365,v_366,v_367,v_368,v_369,v_370,v_371,v_372,v_373,v_374,v_375,v_376,v_377,v_378,v_379,v_380,v_381,v_382,v_383,v_384,v_385,v_386,v_387,v_388,v_389,v_390,v_391,v_392,v_393,v_394,v_395,v_396,v_397,v_398,v_399,v_400,v_401,v_402,v_403,v_404,v_405,v_406,v_407,v_408,v_409,v_410,v_411,v_412,v_413,v_414,v_415,v_416,v_417,v_418,v_419,v_420,v_421,v_422,v_423,v_424,v_425,v_426,v_427,v_428,v_429,v_430,v_431,v_432,v_433,v_434,v_435,v_436,v_437,v_438,v_439,v_440,v_441,v_442,v_443,v_444,v_445,v_446,v_447,v_448,v_449,v_450,v_451,v_452,v_453,v_454,v_455,v_456,v_457,v_458,v_459,v_460,v_461,v_462,v_463,v_464,v_465,v_466,v_467,v_468,v_469,v_470,v_471,v_472,v_473,v_474,v_475,v_476,v_477,v_478,v_479,v_480,v_481,v_482,v_483,v_484,v_485,v_486,v_487,v_488,v_489,v_490,v_491,v_492,v_493,v_494,v_495,v_496,v_497,v_498,v_499,v_500,v_501,v_502,v_503,v_504,v_505,v_506,v_507,v_508,v_509,v_510,v_511,v_512,v_513,v_514,v_515,v_516,v_517,v_518,v_519,v_520,v_521,v_522,v_523,v_524,v_525,v_526,v_527,v_528,v_529,v_530,v_531,v_532,v_533,v_534,v_535,v_536,v_537,v_538,v_539,v_540,v_541,v_542,v_543,v_544,v_545,v_546,v_547,v_548,v_549,v_550,v_551,v_552,v_553,v_554,v_555,v_556,v_557,v_558,v_559,v_560,v_561,v_562,v_563,v_564,v_565,v_566,v_567,v_568,v_569,v_570,v_571,v_572,v_573,v_574,v_575,v_576,v_577,v_578,v_579,v_580,v_581,v_582,v_583,v_584,v_585,v_586,v_587,v_588,v_589,v_590,v_591,v_592,v_593,v_594,v_595,v_596,v_597,v_598,v_599,v_600,v_601,v_602,v_603,v_604,v_605,v_606,v_607,v_608,v_609,v_610,v_611,v_612,v_613,v_614,v_615,v_616,v_617,v_618,v_619,v_620,v_621,v_622,v_623,v_624,v_625,v_626,v_627,v_628,v_629,v_630,v_631,v_632,v_633,v_634,v_635,v_636,v_637,v_638,v_639,v_640,v_641,v_642,v_643,v_644,v_645,v_646,v_647,v_648,v_649,v_650,v_651,v_652,v_653,v_654,v_655,v_656,v_657,v_658,v_659,v_660,v_661,v_662,v_663,v_664,v_665,v_666,v_667,v_668,v_669,v_670,v_671,v_672,v_673,v_674,v_675,v_676,v_677,v_678,v_679,v_680,v_681,v_682,v_683,v_684,v_685,v_686,v_687,v_688,v_689,v_690,v_691,v_692,v_693,v_695,v_696,v_697,v_698,v_699,v_700,v_701,v_702,v_703,v_704,v_705,v_706,v_707,v_708,v_709,v_710,v_711,v_712,v_713,v_714,v_715,v_716,v_717,v_718,v_719,v_720,v_721,v_722,v_723,v_724,v_725,v_726,v_727,v_728,v_729,v_730,v_731,v_732,v_733,v_734,v_735,v_736,v_737,v_738,v_739,v_740,v_741,v_742,v_743,v_744,v_745,v_746,v_747,v_748,v_749,v_750,v_751,v_752,v_753,v_754,v_755,v_756,v_757,v_758,v_759,v_760,v_761,v_762,v_763,v_764,v_765,v_766,v_767,v_768,v_769,v_770,v_771,v_772,v_773,v_774,v_775,v_776,v_777,v_778,v_779,v_780,v_781,v_782,v_784,v_785,v_786,v_787,v_788,v_789,v_790,v_791,v_792,v_793,v_794,v_795,v_796,v_797,v_798,v_799,v_800,v_801,v_802,v_803,v_804,v_805,v_807,v_808,v_809,v_810,v_811,v_812,v_813,v_814,v_815,v_816,v_817,v_818,v_819,v_820,v_821,v_822,v_823,v_824,v_825,v_826,v_827,v_828,v_830,v_831,v_832,v_833,v_834,v_835,v_836,v_837,v_839,v_840,v_841,v_842,v_843,v_844,v_845,v_846,v_848,v_849,v_850,v_851,v_852,v_853,v_854,v_855,v_857,v_858,v_859,v_860,v_861,v_862,v_863,v_864,v_866,v_867,v_868,v_869,v_870,v_871,v_872,v_873,v_874,v_875,v_876,v_877,v_878,v_879,v_880,v_881,v_882,v_883,v_884,v_885,v_886,v_887,v_888,v_889,v_890,v_891,v_892,v_893,v_894,v_895,v_896,v_897,v_898,v_899,v_900,v_901,v_902,v_903,v_904,v_905,v_906,v_907,v_909,v_910,v_911,v_912,v_913,v_914,v_915,v_916,v_917,v_918,v_919,v_920,v_921,v_922,v_923,v_924,v_925,v_926,v_927,v_928,v_929,v_930,v_931,v_932,v_933,v_934,v_935,v_936,v_937,v_938,v_939,v_940,v_941,v_942,v_943,v_944,v_945,v_946,v_947,v_948,v_950,v_951,v_952,v_953,v_954,v_955,v_956,v_957,v_959,v_960,v_961,v_962,v_963,v_964,v_965,v_966,v_968,v_969,v_970,v_971,v_972,v_973,v_974,v_975,v_977,v_978,v_979,v_980,v_981,v_982,v_983,v_984,v_986,v_987,v_988,v_989,v_990,v_991,v_992,v_993,v_995,v_996,v_997,v_998,v_999,v_1000,v_1001,v_1002,v_1003,v_1004,v_1005,v_1006,v_1007,v_1008,v_1009,v_1010,v_1011,v_1012,v_1013,v_1014,v_1015,v_1016,v_1017,v_1018,v_1019,v_1020,v_1021,v_1022,v_1023,v_1024,v_1025,v_1026,v_1027,v_1028,v_1029,v_1030,v_1031,v_1032,o_1);
	input v_1;
	input v_2;
	input v_3;
	input v_4;
	input v_5;
	input v_6;
	input v_7;
	input v_8;
	input v_25;
	input v_26;
	input v_27;
	input v_28;
	input v_29;
	input v_30;
	input v_31;
	input v_32;
	input v_33;
	input v_34;
	input v_35;
	input v_36;
	input v_37;
	input v_38;
	input v_39;
	input v_40;
	input v_41;
	input v_42;
	input v_43;
	input v_44;
	input v_45;
	input v_46;
	input v_47;
	input v_48;
	input v_49;
	input v_50;
	input v_51;
	input v_52;
	input v_53;
	input v_54;
	input v_55;
	input v_56;
	input v_57;
	input v_58;
	input v_59;
	input v_60;
	input v_61;
	input v_62;
	input v_63;
	input v_64;
	input v_65;
	input v_66;
	input v_67;
	input v_68;
	input v_69;
	input v_70;
	input v_71;
	input v_72;
	input v_73;
	input v_74;
	input v_75;
	input v_76;
	input v_77;
	input v_78;
	input v_79;
	input v_80;
	input v_81;
	input v_82;
	input v_83;
	input v_84;
	input v_85;
	input v_86;
	input v_87;
	input v_88;
	input v_89;
	input v_90;
	input v_9;
	input v_10;
	input v_11;
	input v_12;
	input v_13;
	input v_14;
	input v_15;
	input v_16;
	input v_17;
	input v_18;
	input v_19;
	input v_20;
	input v_21;
	input v_22;
	input v_23;
	input v_24;
	input v_91;
	input v_92;
	input v_93;
	input v_94;
	input v_95;
	input v_96;
	input v_97;
	input v_98;
	input v_99;
	input v_100;
	input v_101;
	input v_102;
	input v_103;
	input v_104;
	input v_105;
	input v_106;
	input v_107;
	input v_108;
	input v_109;
	input v_110;
	input v_111;
	input v_112;
	input v_113;
	input v_114;
	input v_115;
	input v_116;
	input v_117;
	input v_118;
	input v_119;
	input v_120;
	input v_121;
	input v_122;
	input v_123;
	input v_124;
	input v_125;
	input v_126;
	input v_127;
	input v_128;
	input v_129;
	input v_130;
	input v_131;
	input v_132;
	input v_133;
	input v_134;
	input v_135;
	input v_136;
	input v_137;
	input v_138;
	input v_139;
	input v_140;
	input v_141;
	input v_142;
	input v_143;
	input v_144;
	input v_145;
	input v_146;
	input v_147;
	input v_148;
	input v_149;
	input v_150;
	input v_151;
	input v_152;
	input v_153;
	input v_154;
	input v_155;
	input v_156;
	input v_157;
	input v_158;
	input v_159;
	input v_160;
	input v_161;
	input v_162;
	input v_163;
	input v_164;
	input v_165;
	input v_166;
	input v_167;
	input v_168;
	input v_169;
	input v_170;
	input v_171;
	input v_172;
	input v_173;
	input v_174;
	input v_175;
	input v_176;
	input v_177;
	input v_178;
	input v_179;
	input v_180;
	input v_181;
	input v_182;
	input v_183;
	input v_184;
	input v_185;
	input v_186;
	input v_187;
	input v_188;
	input v_189;
	input v_190;
	input v_191;
	input v_192;
	input v_193;
	input v_194;
	input v_195;
	input v_196;
	input v_197;
	input v_198;
	input v_199;
	input v_200;
	input v_201;
	input v_202;
	input v_203;
	input v_204;
	input v_205;
	input v_206;
	input v_207;
	input v_208;
	input v_209;
	input v_210;
	input v_211;
	input v_212;
	input v_213;
	input v_214;
	input v_215;
	input v_216;
	input v_217;
	input v_218;
	input v_219;
	input v_220;
	input v_221;
	input v_222;
	input v_223;
	input v_224;
	input v_225;
	input v_226;
	input v_227;
	input v_228;
	input v_229;
	input v_230;
	input v_231;
	input v_232;
	input v_233;
	input v_234;
	input v_235;
	input v_236;
	input v_237;
	input v_238;
	input v_239;
	input v_240;
	input v_241;
	input v_242;
	input v_243;
	input v_244;
	input v_245;
	input v_246;
	input v_247;
	input v_248;
	input v_249;
	input v_250;
	input v_251;
	input v_252;
	input v_253;
	input v_254;
	input v_255;
	input v_256;
	input v_257;
	input v_258;
	input v_259;
	input v_260;
	input v_261;
	input v_262;
	input v_263;
	input v_264;
	input v_265;
	input v_266;
	input v_267;
	input v_268;
	input v_269;
	input v_270;
	input v_271;
	input v_272;
	input v_273;
	input v_274;
	input v_275;
	input v_276;
	input v_277;
	input v_278;
	input v_279;
	input v_280;
	input v_281;
	input v_282;
	input v_283;
	input v_284;
	input v_285;
	input v_286;
	input v_287;
	input v_288;
	input v_289;
	input v_290;
	input v_291;
	input v_292;
	input v_293;
	input v_294;
	input v_295;
	input v_296;
	input v_297;
	input v_298;
	input v_299;
	input v_300;
	input v_301;
	input v_302;
	input v_303;
	input v_304;
	input v_305;
	input v_306;
	input v_307;
	input v_308;
	input v_309;
	input v_310;
	input v_311;
	input v_312;
	input v_313;
	input v_314;
	input v_315;
	input v_316;
	input v_317;
	input v_318;
	input v_319;
	input v_320;
	input v_321;
	input v_322;
	input v_323;
	input v_324;
	input v_325;
	input v_326;
	input v_327;
	input v_328;
	input v_329;
	input v_330;
	input v_331;
	input v_332;
	input v_333;
	input v_334;
	input v_335;
	input v_336;
	input v_337;
	input v_338;
	input v_339;
	input v_340;
	input v_341;
	input v_342;
	input v_343;
	input v_344;
	input v_345;
	input v_346;
	input v_347;
	input v_348;
	input v_349;
	input v_350;
	input v_351;
	input v_352;
	input v_353;
	input v_354;
	input v_355;
	input v_356;
	input v_357;
	input v_358;
	input v_359;
	input v_360;
	input v_361;
	input v_362;
	input v_363;
	input v_364;
	input v_365;
	input v_366;
	input v_367;
	input v_368;
	input v_369;
	input v_370;
	input v_371;
	input v_372;
	input v_373;
	input v_374;
	input v_375;
	input v_376;
	input v_377;
	input v_378;
	input v_379;
	input v_380;
	input v_381;
	input v_382;
	input v_383;
	input v_384;
	input v_385;
	input v_386;
	input v_387;
	input v_388;
	input v_389;
	input v_390;
	input v_391;
	input v_392;
	input v_393;
	input v_394;
	input v_395;
	input v_396;
	input v_397;
	input v_398;
	input v_399;
	input v_400;
	input v_401;
	input v_402;
	input v_403;
	input v_404;
	input v_405;
	input v_406;
	input v_407;
	input v_408;
	input v_409;
	input v_410;
	input v_411;
	input v_412;
	input v_413;
	input v_414;
	input v_415;
	input v_416;
	input v_417;
	input v_418;
	input v_419;
	input v_420;
	input v_421;
	input v_422;
	input v_423;
	input v_424;
	input v_425;
	input v_426;
	input v_427;
	input v_428;
	input v_429;
	input v_430;
	input v_431;
	input v_432;
	input v_433;
	input v_434;
	input v_435;
	input v_436;
	input v_437;
	input v_438;
	input v_439;
	input v_440;
	input v_441;
	input v_442;
	input v_443;
	input v_444;
	input v_445;
	input v_446;
	input v_447;
	input v_448;
	input v_449;
	input v_450;
	input v_451;
	input v_452;
	input v_453;
	input v_454;
	input v_455;
	input v_456;
	input v_457;
	input v_458;
	input v_459;
	input v_460;
	input v_461;
	input v_462;
	input v_463;
	input v_464;
	input v_465;
	input v_466;
	input v_467;
	input v_468;
	input v_469;
	input v_470;
	input v_471;
	input v_472;
	input v_473;
	input v_474;
	input v_475;
	input v_476;
	input v_477;
	input v_478;
	input v_479;
	input v_480;
	input v_481;
	input v_482;
	input v_483;
	input v_484;
	input v_485;
	input v_486;
	input v_487;
	input v_488;
	input v_489;
	input v_490;
	input v_491;
	input v_492;
	input v_493;
	input v_494;
	input v_495;
	input v_496;
	input v_497;
	input v_498;
	input v_499;
	input v_500;
	input v_501;
	input v_502;
	input v_503;
	input v_504;
	input v_505;
	input v_506;
	input v_507;
	input v_508;
	input v_509;
	input v_510;
	input v_511;
	input v_512;
	input v_513;
	input v_514;
	input v_515;
	input v_516;
	input v_517;
	input v_518;
	input v_519;
	input v_520;
	input v_521;
	input v_522;
	input v_523;
	input v_524;
	input v_525;
	input v_526;
	input v_527;
	input v_528;
	input v_529;
	input v_530;
	input v_531;
	input v_532;
	input v_533;
	input v_534;
	input v_535;
	input v_536;
	input v_537;
	input v_538;
	input v_539;
	input v_540;
	input v_541;
	input v_542;
	input v_543;
	input v_544;
	input v_545;
	input v_546;
	input v_547;
	input v_548;
	input v_549;
	input v_550;
	input v_551;
	input v_552;
	input v_553;
	input v_554;
	input v_555;
	input v_556;
	input v_557;
	input v_558;
	input v_559;
	input v_560;
	input v_561;
	input v_562;
	input v_563;
	input v_564;
	input v_565;
	input v_566;
	input v_567;
	input v_568;
	input v_569;
	input v_570;
	input v_571;
	input v_572;
	input v_573;
	input v_574;
	input v_575;
	input v_576;
	input v_577;
	input v_578;
	input v_579;
	input v_580;
	input v_581;
	input v_582;
	input v_583;
	input v_584;
	input v_585;
	input v_586;
	input v_587;
	input v_588;
	input v_589;
	input v_590;
	input v_591;
	input v_592;
	input v_593;
	input v_594;
	input v_595;
	input v_596;
	input v_597;
	input v_598;
	input v_599;
	input v_600;
	input v_601;
	input v_602;
	input v_603;
	input v_604;
	input v_605;
	input v_606;
	input v_607;
	input v_608;
	input v_609;
	input v_610;
	input v_611;
	input v_612;
	input v_613;
	input v_614;
	input v_615;
	input v_616;
	input v_617;
	input v_618;
	input v_619;
	input v_620;
	input v_621;
	input v_622;
	input v_623;
	input v_624;
	input v_625;
	input v_626;
	input v_627;
	input v_628;
	input v_629;
	input v_630;
	input v_631;
	input v_632;
	input v_633;
	input v_634;
	input v_635;
	input v_636;
	input v_637;
	input v_638;
	input v_639;
	input v_640;
	input v_641;
	input v_642;
	input v_643;
	input v_644;
	input v_645;
	input v_646;
	input v_647;
	input v_648;
	input v_649;
	input v_650;
	input v_651;
	input v_652;
	input v_653;
	input v_654;
	input v_655;
	input v_656;
	input v_657;
	input v_658;
	input v_659;
	input v_660;
	input v_661;
	input v_662;
	input v_663;
	input v_664;
	input v_665;
	input v_666;
	input v_667;
	input v_668;
	input v_669;
	input v_670;
	input v_671;
	input v_672;
	input v_673;
	input v_674;
	input v_675;
	input v_676;
	input v_677;
	input v_678;
	input v_679;
	input v_680;
	input v_681;
	input v_682;
	input v_683;
	input v_684;
	input v_685;
	input v_686;
	input v_687;
	input v_688;
	input v_689;
	input v_690;
	input v_691;
	input v_692;
	input v_693;
	input v_695;
	input v_696;
	input v_697;
	input v_698;
	input v_699;
	input v_700;
	input v_701;
	input v_702;
	input v_703;
	input v_704;
	input v_705;
	input v_706;
	input v_707;
	input v_708;
	input v_709;
	input v_710;
	input v_711;
	input v_712;
	input v_713;
	input v_714;
	input v_715;
	input v_716;
	input v_717;
	input v_718;
	input v_719;
	input v_720;
	input v_721;
	input v_722;
	input v_723;
	input v_724;
	input v_725;
	input v_726;
	input v_727;
	input v_728;
	input v_729;
	input v_730;
	input v_731;
	input v_732;
	input v_733;
	input v_734;
	input v_735;
	input v_736;
	input v_737;
	input v_738;
	input v_739;
	input v_740;
	input v_741;
	input v_742;
	input v_743;
	input v_744;
	input v_745;
	input v_746;
	input v_747;
	input v_748;
	input v_749;
	input v_750;
	input v_751;
	input v_752;
	input v_753;
	input v_754;
	input v_755;
	input v_756;
	input v_757;
	input v_758;
	input v_759;
	input v_760;
	input v_761;
	input v_762;
	input v_763;
	input v_764;
	input v_765;
	input v_766;
	input v_767;
	input v_768;
	input v_769;
	input v_770;
	input v_771;
	input v_772;
	input v_773;
	input v_774;
	input v_775;
	input v_776;
	input v_777;
	input v_778;
	input v_779;
	input v_780;
	input v_781;
	input v_782;
	input v_784;
	input v_785;
	input v_786;
	input v_787;
	input v_788;
	input v_789;
	input v_790;
	input v_791;
	input v_792;
	input v_793;
	input v_794;
	input v_795;
	input v_796;
	input v_797;
	input v_798;
	input v_799;
	input v_800;
	input v_801;
	input v_802;
	input v_803;
	input v_804;
	input v_805;
	input v_807;
	input v_808;
	input v_809;
	input v_810;
	input v_811;
	input v_812;
	input v_813;
	input v_814;
	input v_815;
	input v_816;
	input v_817;
	input v_818;
	input v_819;
	input v_820;
	input v_821;
	input v_822;
	input v_823;
	input v_824;
	input v_825;
	input v_826;
	input v_827;
	input v_828;
	input v_830;
	input v_831;
	input v_832;
	input v_833;
	input v_834;
	input v_835;
	input v_836;
	input v_837;
	input v_839;
	input v_840;
	input v_841;
	input v_842;
	input v_843;
	input v_844;
	input v_845;
	input v_846;
	input v_848;
	input v_849;
	input v_850;
	input v_851;
	input v_852;
	input v_853;
	input v_854;
	input v_855;
	input v_857;
	input v_858;
	input v_859;
	input v_860;
	input v_861;
	input v_862;
	input v_863;
	input v_864;
	input v_866;
	input v_867;
	input v_868;
	input v_869;
	input v_870;
	input v_871;
	input v_872;
	input v_873;
	input v_874;
	input v_875;
	input v_876;
	input v_877;
	input v_878;
	input v_879;
	input v_880;
	input v_881;
	input v_882;
	input v_883;
	input v_884;
	input v_885;
	input v_886;
	input v_887;
	input v_888;
	input v_889;
	input v_890;
	input v_891;
	input v_892;
	input v_893;
	input v_894;
	input v_895;
	input v_896;
	input v_897;
	input v_898;
	input v_899;
	input v_900;
	input v_901;
	input v_902;
	input v_903;
	input v_904;
	input v_905;
	input v_906;
	input v_907;
	input v_909;
	input v_910;
	input v_911;
	input v_912;
	input v_913;
	input v_914;
	input v_915;
	input v_916;
	input v_917;
	input v_918;
	input v_919;
	input v_920;
	input v_921;
	input v_922;
	input v_923;
	input v_924;
	input v_925;
	input v_926;
	input v_927;
	input v_928;
	input v_929;
	input v_930;
	input v_931;
	input v_932;
	input v_933;
	input v_934;
	input v_935;
	input v_936;
	input v_937;
	input v_938;
	input v_939;
	input v_940;
	input v_941;
	input v_942;
	input v_943;
	input v_944;
	input v_945;
	input v_946;
	input v_947;
	input v_948;
	input v_950;
	input v_951;
	input v_952;
	input v_953;
	input v_954;
	input v_955;
	input v_956;
	input v_957;
	input v_959;
	input v_960;
	input v_961;
	input v_962;
	input v_963;
	input v_964;
	input v_965;
	input v_966;
	input v_968;
	input v_969;
	input v_970;
	input v_971;
	input v_972;
	input v_973;
	input v_974;
	input v_975;
	input v_977;
	input v_978;
	input v_979;
	input v_980;
	input v_981;
	input v_982;
	input v_983;
	input v_984;
	input v_986;
	input v_987;
	input v_988;
	input v_989;
	input v_990;
	input v_991;
	input v_992;
	input v_993;
	input v_995;
	input v_996;
	input v_997;
	input v_998;
	input v_999;
	input v_1000;
	input v_1001;
	input v_1002;
	input v_1003;
	input v_1004;
	input v_1005;
	input v_1006;
	input v_1007;
	input v_1008;
	input v_1009;
	input v_1010;
	input v_1011;
	input v_1012;
	input v_1013;
	input v_1014;
	input v_1015;
	input v_1016;
	input v_1017;
	input v_1018;
	input v_1019;
	input v_1020;
	input v_1021;
	input v_1022;
	input v_1023;
	input v_1024;
	input v_1025;
	input v_1026;
	input v_1027;
	input v_1028;
	input v_1029;
	input v_1030;
	input v_1031;
	input v_1032;
	wire v_694;
	wire v_783;
	wire v_806;
	wire v_829;
	wire v_838;
	wire v_847;
	wire v_856;
	wire v_865;
	wire v_908;
	wire v_949;
	wire v_958;
	wire v_967;
	wire v_976;
	wire v_985;
	wire v_994;
	wire v_1033;
	wire v_1034;
	wire x_1;
	wire x_2;
	wire x_3;
	wire x_4;
	wire x_5;
	wire x_6;
	wire x_7;
	wire x_8;
	wire x_9;
	wire x_10;
	wire x_11;
	wire x_12;
	wire x_13;
	wire x_14;
	wire x_15;
	wire x_16;
	wire x_17;
	wire x_18;
	wire x_19;
	wire x_20;
	wire x_21;
	wire x_22;
	wire x_23;
	wire x_24;
	wire x_25;
	wire x_26;
	wire x_27;
	wire x_28;
	wire x_29;
	wire x_30;
	wire x_31;
	wire x_32;
	wire x_33;
	wire x_34;
	wire x_35;
	wire x_36;
	wire x_37;
	wire x_38;
	wire x_39;
	wire x_40;
	wire x_41;
	wire x_42;
	wire x_43;
	wire x_44;
	wire x_45;
	wire x_46;
	wire x_47;
	wire x_48;
	wire x_49;
	wire x_50;
	wire x_51;
	wire x_52;
	wire x_53;
	wire x_54;
	wire x_55;
	wire x_56;
	wire x_57;
	wire x_58;
	wire x_59;
	wire x_60;
	wire x_61;
	wire x_62;
	wire x_63;
	wire x_64;
	wire x_65;
	wire x_66;
	wire x_67;
	wire x_68;
	wire x_69;
	wire x_70;
	wire x_71;
	wire x_72;
	wire x_73;
	wire x_74;
	wire x_75;
	wire x_76;
	wire x_77;
	wire x_78;
	wire x_79;
	wire x_80;
	wire x_81;
	wire x_82;
	wire x_83;
	wire x_84;
	wire x_85;
	wire x_86;
	wire x_87;
	wire x_88;
	wire x_89;
	wire x_90;
	wire x_91;
	wire x_92;
	wire x_93;
	wire x_94;
	wire x_95;
	wire x_96;
	wire x_97;
	wire x_98;
	wire x_99;
	wire x_100;
	wire x_101;
	wire x_102;
	wire x_103;
	wire x_104;
	wire x_105;
	wire x_106;
	wire x_107;
	wire x_108;
	wire x_109;
	wire x_110;
	wire x_111;
	wire x_112;
	wire x_113;
	wire x_114;
	wire x_115;
	wire x_116;
	wire x_117;
	wire x_118;
	wire x_119;
	wire x_120;
	wire x_121;
	wire x_122;
	wire x_123;
	wire x_124;
	wire x_125;
	wire x_126;
	wire x_127;
	wire x_128;
	wire x_129;
	wire x_130;
	wire x_131;
	wire x_132;
	wire x_133;
	wire x_134;
	wire x_135;
	wire x_136;
	wire x_137;
	wire x_138;
	wire x_139;
	wire x_140;
	wire x_141;
	wire x_142;
	wire x_143;
	wire x_144;
	wire x_145;
	wire x_146;
	wire x_147;
	wire x_148;
	wire x_149;
	wire x_150;
	wire x_151;
	wire x_152;
	wire x_153;
	wire x_154;
	wire x_155;
	wire x_156;
	wire x_157;
	wire x_158;
	wire x_159;
	wire x_160;
	wire x_161;
	wire x_162;
	wire x_163;
	wire x_164;
	wire x_165;
	wire x_166;
	wire x_167;
	wire x_168;
	wire x_169;
	wire x_170;
	wire x_171;
	wire x_172;
	wire x_173;
	wire x_174;
	wire x_175;
	wire x_176;
	wire x_177;
	wire x_178;
	wire x_179;
	wire x_180;
	wire x_181;
	wire x_182;
	wire x_183;
	wire x_184;
	wire x_185;
	wire x_186;
	wire x_187;
	wire x_188;
	wire x_189;
	wire x_190;
	wire x_191;
	wire x_192;
	wire x_193;
	wire x_194;
	wire x_195;
	wire x_196;
	wire x_197;
	wire x_198;
	wire x_199;
	wire x_200;
	wire x_201;
	wire x_202;
	wire x_203;
	wire x_204;
	wire x_205;
	wire x_206;
	wire x_207;
	wire x_208;
	wire x_209;
	wire x_210;
	wire x_211;
	wire x_212;
	wire x_213;
	wire x_214;
	wire x_215;
	wire x_216;
	wire x_217;
	wire x_218;
	wire x_219;
	wire x_220;
	wire x_221;
	wire x_222;
	wire x_223;
	wire x_224;
	wire x_225;
	wire x_226;
	wire x_227;
	wire x_228;
	wire x_229;
	wire x_230;
	wire x_231;
	wire x_232;
	wire x_233;
	wire x_234;
	wire x_235;
	wire x_236;
	wire x_237;
	wire x_238;
	wire x_239;
	wire x_240;
	wire x_241;
	wire x_242;
	wire x_243;
	wire x_244;
	wire x_245;
	wire x_246;
	wire x_247;
	wire x_248;
	wire x_249;
	wire x_250;
	wire x_251;
	wire x_252;
	wire x_253;
	wire x_254;
	wire x_255;
	wire x_256;
	wire x_257;
	wire x_258;
	wire x_259;
	wire x_260;
	wire x_261;
	wire x_262;
	wire x_263;
	wire x_264;
	wire x_265;
	wire x_266;
	wire x_267;
	wire x_268;
	wire x_269;
	wire x_270;
	wire x_271;
	wire x_272;
	wire x_273;
	wire x_274;
	wire x_275;
	wire x_276;
	wire x_277;
	wire x_278;
	wire x_279;
	wire x_280;
	wire x_281;
	wire x_282;
	wire x_283;
	wire x_284;
	wire x_285;
	wire x_286;
	wire x_287;
	wire x_288;
	wire x_289;
	wire x_290;
	wire x_291;
	wire x_292;
	wire x_293;
	wire x_294;
	wire x_295;
	wire x_296;
	wire x_297;
	wire x_298;
	wire x_299;
	wire x_300;
	wire x_301;
	wire x_302;
	wire x_303;
	wire x_304;
	wire x_305;
	wire x_306;
	wire x_307;
	wire x_308;
	wire x_309;
	wire x_310;
	wire x_311;
	wire x_312;
	wire x_313;
	wire x_314;
	wire x_315;
	wire x_316;
	wire x_317;
	wire x_318;
	wire x_319;
	wire x_320;
	wire x_321;
	wire x_322;
	wire x_323;
	wire x_324;
	wire x_325;
	wire x_326;
	wire x_327;
	wire x_328;
	wire x_329;
	wire x_330;
	wire x_331;
	wire x_332;
	wire x_333;
	wire x_334;
	wire x_335;
	wire x_336;
	wire x_337;
	wire x_338;
	wire x_339;
	wire x_340;
	wire x_341;
	wire x_342;
	wire x_343;
	wire x_344;
	wire x_345;
	wire x_346;
	wire x_347;
	wire x_348;
	wire x_349;
	wire x_350;
	wire x_351;
	wire x_352;
	wire x_353;
	wire x_354;
	wire x_355;
	wire x_356;
	wire x_357;
	wire x_358;
	wire x_359;
	wire x_360;
	wire x_361;
	wire x_362;
	wire x_363;
	wire x_364;
	wire x_365;
	wire x_366;
	wire x_367;
	wire x_368;
	wire x_369;
	wire x_370;
	wire x_371;
	wire x_372;
	wire x_373;
	wire x_374;
	wire x_375;
	wire x_376;
	wire x_377;
	wire x_378;
	wire x_379;
	wire x_380;
	wire x_381;
	wire x_382;
	wire x_383;
	wire x_384;
	wire x_385;
	wire x_386;
	wire x_387;
	wire x_388;
	wire x_389;
	wire x_390;
	wire x_391;
	wire x_392;
	wire x_393;
	wire x_394;
	wire x_395;
	wire x_396;
	wire x_397;
	wire x_398;
	wire x_399;
	wire x_400;
	wire x_401;
	wire x_402;
	wire x_403;
	wire x_404;
	wire x_405;
	wire x_406;
	wire x_407;
	wire x_408;
	wire x_409;
	wire x_410;
	wire x_411;
	wire x_412;
	wire x_413;
	wire x_414;
	wire x_415;
	wire x_416;
	wire x_417;
	wire x_418;
	wire x_419;
	wire x_420;
	wire x_421;
	wire x_422;
	wire x_423;
	wire x_424;
	wire x_425;
	wire x_426;
	wire x_427;
	wire x_428;
	wire x_429;
	wire x_430;
	wire x_431;
	wire x_432;
	wire x_433;
	wire x_434;
	wire x_435;
	wire x_436;
	wire x_437;
	wire x_438;
	wire x_439;
	wire x_440;
	wire x_441;
	wire x_442;
	wire x_443;
	wire x_444;
	wire x_445;
	wire x_446;
	wire x_447;
	wire x_448;
	wire x_449;
	wire x_450;
	wire x_451;
	wire x_452;
	wire x_453;
	wire x_454;
	wire x_455;
	wire x_456;
	wire x_457;
	wire x_458;
	wire x_459;
	wire x_460;
	wire x_461;
	wire x_462;
	wire x_463;
	wire x_464;
	wire x_465;
	wire x_466;
	wire x_467;
	wire x_468;
	wire x_469;
	wire x_470;
	wire x_471;
	wire x_472;
	wire x_473;
	wire x_474;
	wire x_475;
	wire x_476;
	wire x_477;
	wire x_478;
	wire x_479;
	wire x_480;
	wire x_481;
	wire x_482;
	wire x_483;
	wire x_484;
	wire x_485;
	wire x_486;
	wire x_487;
	wire x_488;
	wire x_489;
	wire x_490;
	wire x_491;
	wire x_492;
	wire x_493;
	wire x_494;
	wire x_495;
	wire x_496;
	wire x_497;
	wire x_498;
	wire x_499;
	wire x_500;
	wire x_501;
	wire x_502;
	wire x_503;
	wire x_504;
	wire x_505;
	wire x_506;
	wire x_507;
	wire x_508;
	wire x_509;
	wire x_510;
	wire x_511;
	wire x_512;
	wire x_513;
	wire x_514;
	wire x_515;
	wire x_516;
	wire x_517;
	wire x_518;
	wire x_519;
	wire x_520;
	wire x_521;
	wire x_522;
	wire x_523;
	wire x_524;
	wire x_525;
	wire x_526;
	wire x_527;
	wire x_528;
	wire x_529;
	wire x_530;
	wire x_531;
	wire x_532;
	wire x_533;
	wire x_534;
	wire x_535;
	wire x_536;
	wire x_537;
	wire x_538;
	wire x_539;
	wire x_540;
	wire x_541;
	wire x_542;
	wire x_543;
	wire x_544;
	wire x_545;
	wire x_546;
	wire x_547;
	wire x_548;
	wire x_549;
	wire x_550;
	wire x_551;
	wire x_552;
	wire x_553;
	wire x_554;
	wire x_555;
	wire x_556;
	wire x_557;
	wire x_558;
	wire x_559;
	wire x_560;
	wire x_561;
	wire x_562;
	wire x_563;
	wire x_564;
	wire x_565;
	wire x_566;
	wire x_567;
	wire x_568;
	wire x_569;
	wire x_570;
	wire x_571;
	wire x_572;
	wire x_573;
	wire x_574;
	wire x_575;
	wire x_576;
	wire x_577;
	wire x_578;
	wire x_579;
	wire x_580;
	wire x_581;
	wire x_582;
	wire x_583;
	wire x_584;
	wire x_585;
	wire x_586;
	wire x_587;
	wire x_588;
	wire x_589;
	wire x_590;
	wire x_591;
	wire x_592;
	wire x_593;
	wire x_594;
	wire x_595;
	wire x_596;
	wire x_597;
	wire x_598;
	wire x_599;
	wire x_600;
	wire x_601;
	wire x_602;
	wire x_603;
	wire x_604;
	wire x_605;
	wire x_606;
	wire x_607;
	wire x_608;
	wire x_609;
	wire x_610;
	wire x_611;
	wire x_612;
	wire x_613;
	wire x_614;
	wire x_615;
	wire x_616;
	wire x_617;
	wire x_618;
	wire x_619;
	wire x_620;
	wire x_621;
	wire x_622;
	wire x_623;
	wire x_624;
	wire x_625;
	wire x_626;
	wire x_627;
	wire x_628;
	wire x_629;
	wire x_630;
	wire x_631;
	wire x_632;
	wire x_633;
	wire x_634;
	wire x_635;
	wire x_636;
	wire x_637;
	wire x_638;
	wire x_639;
	wire x_640;
	wire x_641;
	wire x_642;
	wire x_643;
	wire x_644;
	wire x_645;
	wire x_646;
	wire x_647;
	wire x_648;
	wire x_649;
	wire x_650;
	wire x_651;
	wire x_652;
	wire x_653;
	wire x_654;
	wire x_655;
	wire x_656;
	wire x_657;
	wire x_658;
	wire x_659;
	wire x_660;
	wire x_661;
	wire x_662;
	wire x_663;
	wire x_664;
	wire x_665;
	wire x_666;
	wire x_667;
	wire x_668;
	wire x_669;
	wire x_670;
	wire x_671;
	wire x_672;
	wire x_673;
	wire x_674;
	wire x_675;
	wire x_676;
	wire x_677;
	wire x_678;
	wire x_679;
	wire x_680;
	wire x_681;
	wire x_682;
	wire x_683;
	wire x_684;
	wire x_685;
	wire x_686;
	wire x_687;
	wire x_688;
	wire x_689;
	wire x_690;
	wire x_691;
	wire x_692;
	wire x_693;
	wire x_694;
	wire x_695;
	wire x_696;
	wire x_697;
	wire x_698;
	wire x_699;
	wire x_700;
	wire x_701;
	wire x_702;
	wire x_703;
	wire x_704;
	wire x_705;
	wire x_706;
	wire x_707;
	wire x_708;
	wire x_709;
	wire x_710;
	wire x_711;
	wire x_712;
	wire x_713;
	wire x_714;
	wire x_715;
	wire x_716;
	wire x_717;
	wire x_718;
	wire x_719;
	wire x_720;
	wire x_721;
	wire x_722;
	wire x_723;
	wire x_724;
	wire x_725;
	wire x_726;
	wire x_727;
	wire x_728;
	wire x_729;
	wire x_730;
	wire x_731;
	wire x_732;
	wire x_733;
	wire x_734;
	wire x_735;
	wire x_736;
	wire x_737;
	wire x_738;
	wire x_739;
	wire x_740;
	wire x_741;
	wire x_742;
	wire x_743;
	wire x_744;
	wire x_745;
	wire x_746;
	wire x_747;
	wire x_748;
	wire x_749;
	wire x_750;
	wire x_751;
	wire x_752;
	wire x_753;
	wire x_754;
	wire x_755;
	wire x_756;
	wire x_757;
	wire x_758;
	wire x_759;
	wire x_760;
	wire x_761;
	wire x_762;
	wire x_763;
	wire x_764;
	wire x_765;
	wire x_766;
	wire x_767;
	wire x_768;
	wire x_769;
	wire x_770;
	wire x_771;
	wire x_772;
	wire x_773;
	wire x_774;
	wire x_775;
	wire x_776;
	wire x_777;
	wire x_778;
	wire x_779;
	wire x_780;
	wire x_781;
	wire x_782;
	wire x_783;
	wire x_784;
	wire x_785;
	wire x_786;
	wire x_787;
	wire x_788;
	wire x_789;
	wire x_790;
	wire x_791;
	wire x_792;
	wire x_793;
	wire x_794;
	wire x_795;
	wire x_796;
	wire x_797;
	wire x_798;
	wire x_799;
	wire x_800;
	wire x_801;
	wire x_802;
	wire x_803;
	wire x_804;
	wire x_805;
	wire x_806;
	wire x_807;
	wire x_808;
	wire x_809;
	wire x_810;
	wire x_811;
	wire x_812;
	wire x_813;
	wire x_814;
	wire x_815;
	wire x_816;
	wire x_817;
	wire x_818;
	wire x_819;
	wire x_820;
	wire x_821;
	wire x_822;
	wire x_823;
	wire x_824;
	wire x_825;
	wire x_826;
	wire x_827;
	wire x_828;
	wire x_829;
	wire x_830;
	wire x_831;
	wire x_832;
	wire x_833;
	wire x_834;
	wire x_835;
	wire x_836;
	wire x_837;
	wire x_838;
	wire x_839;
	wire x_840;
	wire x_841;
	wire x_842;
	wire x_843;
	wire x_844;
	wire x_845;
	wire x_846;
	wire x_847;
	wire x_848;
	wire x_849;
	wire x_850;
	wire x_851;
	wire x_852;
	wire x_853;
	wire x_854;
	wire x_855;
	wire x_856;
	wire x_857;
	wire x_858;
	wire x_859;
	wire x_860;
	wire x_861;
	wire x_862;
	wire x_863;
	wire x_864;
	wire x_865;
	wire x_866;
	wire x_867;
	wire x_868;
	wire x_869;
	wire x_870;
	wire x_871;
	wire x_872;
	wire x_873;
	wire x_874;
	wire x_875;
	wire x_876;
	wire x_877;
	wire x_878;
	wire x_879;
	wire x_880;
	wire x_881;
	wire x_882;
	wire x_883;
	wire x_884;
	wire x_885;
	wire x_886;
	wire x_887;
	wire x_888;
	wire x_889;
	wire x_890;
	wire x_891;
	wire x_892;
	wire x_893;
	wire x_894;
	wire x_895;
	wire x_896;
	wire x_897;
	wire x_898;
	wire x_899;
	wire x_900;
	wire x_901;
	wire x_902;
	wire x_903;
	wire x_904;
	wire x_905;
	wire x_906;
	wire x_907;
	wire x_908;
	wire x_909;
	wire x_910;
	wire x_911;
	wire x_912;
	wire x_913;
	wire x_914;
	wire x_915;
	wire x_916;
	wire x_917;
	wire x_918;
	wire x_919;
	wire x_920;
	wire x_921;
	wire x_922;
	wire x_923;
	wire x_924;
	wire x_925;
	wire x_926;
	wire x_927;
	wire x_928;
	wire x_929;
	wire x_930;
	wire x_931;
	wire x_932;
	wire x_933;
	wire x_934;
	wire x_935;
	wire x_936;
	wire x_937;
	wire x_938;
	wire x_939;
	wire x_940;
	wire x_941;
	wire x_942;
	wire x_943;
	wire x_944;
	wire x_945;
	wire x_946;
	wire x_947;
	wire x_948;
	wire x_949;
	wire x_950;
	wire x_951;
	wire x_952;
	wire x_953;
	wire x_954;
	wire x_955;
	wire x_956;
	wire x_957;
	wire x_958;
	wire x_959;
	wire x_960;
	wire x_961;
	wire x_962;
	wire x_963;
	wire x_964;
	wire x_965;
	wire x_966;
	wire x_967;
	wire x_968;
	wire x_969;
	wire x_970;
	wire x_971;
	wire x_972;
	wire x_973;
	wire x_974;
	wire x_975;
	wire x_976;
	wire x_977;
	wire x_978;
	wire x_979;
	wire x_980;
	wire x_981;
	wire x_982;
	wire x_983;
	wire x_984;
	wire x_985;
	wire x_986;
	wire x_987;
	wire x_988;
	wire x_989;
	wire x_990;
	wire x_991;
	wire x_992;
	wire x_993;
	wire x_994;
	wire x_995;
	wire x_996;
	wire x_997;
	wire x_998;
	wire x_999;
	wire x_1000;
	wire x_1001;
	wire x_1002;
	wire x_1003;
	wire x_1004;
	wire x_1005;
	wire x_1006;
	wire x_1007;
	wire x_1008;
	wire x_1009;
	wire x_1010;
	wire x_1011;
	wire x_1012;
	wire x_1013;
	wire x_1014;
	wire x_1015;
	wire x_1016;
	wire x_1017;
	wire x_1018;
	wire x_1019;
	wire x_1020;
	wire x_1021;
	wire x_1022;
	wire x_1023;
	wire x_1024;
	wire x_1025;
	wire x_1026;
	wire x_1027;
	wire x_1028;
	wire x_1029;
	wire x_1030;
	wire x_1031;
	wire x_1032;
	wire x_1033;
	wire x_1034;
	wire x_1035;
	wire x_1036;
	wire x_1037;
	wire x_1038;
	wire x_1039;
	wire x_1040;
	wire x_1041;
	wire x_1042;
	wire x_1043;
	wire x_1044;
	wire x_1045;
	wire x_1046;
	wire x_1047;
	wire x_1048;
	wire x_1049;
	wire x_1050;
	wire x_1051;
	wire x_1052;
	wire x_1053;
	wire x_1054;
	wire x_1055;
	wire x_1056;
	wire x_1057;
	wire x_1058;
	wire x_1059;
	wire x_1060;
	wire x_1061;
	wire x_1062;
	wire x_1063;
	wire x_1064;
	wire x_1065;
	wire x_1066;
	wire x_1067;
	wire x_1068;
	wire x_1069;
	wire x_1070;
	wire x_1071;
	wire x_1072;
	wire x_1073;
	wire x_1074;
	wire x_1075;
	wire x_1076;
	wire x_1077;
	wire x_1078;
	wire x_1079;
	wire x_1080;
	wire x_1081;
	wire x_1082;
	wire x_1083;
	wire x_1084;
	wire x_1085;
	wire x_1086;
	wire x_1087;
	wire x_1088;
	wire x_1089;
	wire x_1090;
	wire x_1091;
	wire x_1092;
	wire x_1093;
	wire x_1094;
	wire x_1095;
	wire x_1096;
	wire x_1097;
	wire x_1098;
	wire x_1099;
	wire x_1100;
	wire x_1101;
	wire x_1102;
	wire x_1103;
	wire x_1104;
	wire x_1105;
	wire x_1106;
	wire x_1107;
	wire x_1108;
	wire x_1109;
	wire x_1110;
	wire x_1111;
	wire x_1112;
	wire x_1113;
	wire x_1114;
	wire x_1115;
	wire x_1116;
	wire x_1117;
	wire x_1118;
	wire x_1119;
	wire x_1120;
	wire x_1121;
	wire x_1122;
	wire x_1123;
	wire x_1124;
	wire x_1125;
	wire x_1126;
	wire x_1127;
	wire x_1128;
	wire x_1129;
	wire x_1130;
	wire x_1131;
	wire x_1132;
	wire x_1133;
	wire x_1134;
	wire x_1135;
	wire x_1136;
	wire x_1137;
	wire x_1138;
	wire x_1139;
	wire x_1140;
	wire x_1141;
	wire x_1142;
	wire x_1143;
	wire x_1144;
	wire x_1145;
	wire x_1146;
	wire x_1147;
	wire x_1148;
	wire x_1149;
	wire x_1150;
	wire x_1151;
	wire x_1152;
	wire x_1153;
	wire x_1154;
	wire x_1155;
	wire x_1156;
	wire x_1157;
	wire x_1158;
	wire x_1159;
	wire x_1160;
	wire x_1161;
	wire x_1162;
	wire x_1163;
	wire x_1164;
	wire x_1165;
	wire x_1166;
	wire x_1167;
	wire x_1168;
	wire x_1169;
	wire x_1170;
	wire x_1171;
	wire x_1172;
	wire x_1173;
	wire x_1174;
	wire x_1175;
	wire x_1176;
	wire x_1177;
	wire x_1178;
	wire x_1179;
	wire x_1180;
	wire x_1181;
	wire x_1182;
	wire x_1183;
	wire x_1184;
	wire x_1185;
	wire x_1186;
	wire x_1187;
	wire x_1188;
	wire x_1189;
	wire x_1190;
	wire x_1191;
	wire x_1192;
	wire x_1193;
	wire x_1194;
	wire x_1195;
	wire x_1196;
	wire x_1197;
	wire x_1198;
	wire x_1199;
	wire x_1200;
	wire x_1201;
	wire x_1202;
	wire x_1203;
	wire x_1204;
	wire x_1205;
	wire x_1206;
	wire x_1207;
	wire x_1208;
	wire x_1209;
	wire x_1210;
	wire x_1211;
	wire x_1212;
	wire x_1213;
	wire x_1214;
	wire x_1215;
	wire x_1216;
	wire x_1217;
	wire x_1218;
	wire x_1219;
	wire x_1220;
	wire x_1221;
	wire x_1222;
	wire x_1223;
	wire x_1224;
	wire x_1225;
	wire x_1226;
	wire x_1227;
	wire x_1228;
	wire x_1229;
	wire x_1230;
	wire x_1231;
	wire x_1232;
	wire x_1233;
	wire x_1234;
	wire x_1235;
	wire x_1236;
	wire x_1237;
	wire x_1238;
	wire x_1239;
	wire x_1240;
	wire x_1241;
	wire x_1242;
	wire x_1243;
	wire x_1244;
	wire x_1245;
	wire x_1246;
	wire x_1247;
	wire x_1248;
	wire x_1249;
	wire x_1250;
	wire x_1251;
	wire x_1252;
	wire x_1253;
	wire x_1254;
	wire x_1255;
	wire x_1256;
	wire x_1257;
	wire x_1258;
	wire x_1259;
	wire x_1260;
	wire x_1261;
	wire x_1262;
	wire x_1263;
	wire x_1264;
	wire x_1265;
	wire x_1266;
	wire x_1267;
	wire x_1268;
	wire x_1269;
	wire x_1270;
	wire x_1271;
	wire x_1272;
	wire x_1273;
	wire x_1274;
	wire x_1275;
	wire x_1276;
	wire x_1277;
	wire x_1278;
	wire x_1279;
	wire x_1280;
	wire x_1281;
	wire x_1282;
	wire x_1283;
	wire x_1284;
	wire x_1285;
	wire x_1286;
	wire x_1287;
	wire x_1288;
	wire x_1289;
	wire x_1290;
	wire x_1291;
	wire x_1292;
	wire x_1293;
	wire x_1294;
	wire x_1295;
	wire x_1296;
	wire x_1297;
	wire x_1298;
	wire x_1299;
	wire x_1300;
	wire x_1301;
	wire x_1302;
	wire x_1303;
	wire x_1304;
	wire x_1305;
	wire x_1306;
	wire x_1307;
	wire x_1308;
	wire x_1309;
	wire x_1310;
	wire x_1311;
	wire x_1312;
	wire x_1313;
	wire x_1314;
	wire x_1315;
	wire x_1316;
	wire x_1317;
	wire x_1318;
	wire x_1319;
	wire x_1320;
	wire x_1321;
	wire x_1322;
	wire x_1323;
	wire x_1324;
	wire x_1325;
	wire x_1326;
	wire x_1327;
	wire x_1328;
	wire x_1329;
	wire x_1330;
	wire x_1331;
	wire x_1332;
	wire x_1333;
	wire x_1334;
	wire x_1335;
	wire x_1336;
	wire x_1337;
	wire x_1338;
	wire x_1339;
	wire x_1340;
	wire x_1341;
	wire x_1342;
	wire x_1343;
	wire x_1344;
	wire x_1345;
	wire x_1346;
	wire x_1347;
	wire x_1348;
	wire x_1349;
	wire x_1350;
	wire x_1351;
	wire x_1352;
	wire x_1353;
	wire x_1354;
	wire x_1355;
	wire x_1356;
	wire x_1357;
	wire x_1358;
	wire x_1359;
	wire x_1360;
	wire x_1361;
	wire x_1362;
	wire x_1363;
	wire x_1364;
	wire x_1365;
	wire x_1366;
	wire x_1367;
	wire x_1368;
	wire x_1369;
	wire x_1370;
	wire x_1371;
	wire x_1372;
	wire x_1373;
	wire x_1374;
	wire x_1375;
	wire x_1376;
	wire x_1377;
	wire x_1378;
	wire x_1379;
	wire x_1380;
	wire x_1381;
	wire x_1382;
	wire x_1383;
	wire x_1384;
	wire x_1385;
	wire x_1386;
	wire x_1387;
	wire x_1388;
	wire x_1389;
	wire x_1390;
	wire x_1391;
	wire x_1392;
	wire x_1393;
	wire x_1394;
	wire x_1395;
	wire x_1396;
	wire x_1397;
	wire x_1398;
	wire x_1399;
	wire x_1400;
	wire x_1401;
	wire x_1402;
	wire x_1403;
	wire x_1404;
	wire x_1405;
	wire x_1406;
	wire x_1407;
	wire x_1408;
	wire x_1409;
	wire x_1410;
	wire x_1411;
	wire x_1412;
	wire x_1413;
	wire x_1414;
	wire x_1415;
	wire x_1416;
	wire x_1417;
	wire x_1418;
	wire x_1419;
	wire x_1420;
	wire x_1421;
	wire x_1422;
	wire x_1423;
	wire x_1424;
	wire x_1425;
	wire x_1426;
	wire x_1427;
	wire x_1428;
	wire x_1429;
	wire x_1430;
	wire x_1431;
	wire x_1432;
	wire x_1433;
	wire x_1434;
	wire x_1435;
	wire x_1436;
	wire x_1437;
	wire x_1438;
	wire x_1439;
	wire x_1440;
	wire x_1441;
	wire x_1442;
	wire x_1443;
	wire x_1444;
	wire x_1445;
	wire x_1446;
	wire x_1447;
	wire x_1448;
	wire x_1449;
	wire x_1450;
	wire x_1451;
	wire x_1452;
	wire x_1453;
	wire x_1454;
	wire x_1455;
	wire x_1456;
	wire x_1457;
	wire x_1458;
	wire x_1459;
	wire x_1460;
	wire x_1461;
	wire x_1462;
	wire x_1463;
	wire x_1464;
	wire x_1465;
	wire x_1466;
	wire x_1467;
	wire x_1468;
	wire x_1469;
	wire x_1470;
	wire x_1471;
	wire x_1472;
	wire x_1473;
	wire x_1474;
	wire x_1475;
	wire x_1476;
	wire x_1477;
	wire x_1478;
	wire x_1479;
	wire x_1480;
	wire x_1481;
	wire x_1482;
	wire x_1483;
	wire x_1484;
	wire x_1485;
	wire x_1486;
	wire x_1487;
	wire x_1488;
	wire x_1489;
	wire x_1490;
	wire x_1491;
	wire x_1492;
	wire x_1493;
	wire x_1494;
	wire x_1495;
	wire x_1496;
	wire x_1497;
	wire x_1498;
	wire x_1499;
	wire x_1500;
	wire x_1501;
	wire x_1502;
	wire x_1503;
	wire x_1504;
	wire x_1505;
	wire x_1506;
	wire x_1507;
	wire x_1508;
	wire x_1509;
	wire x_1510;
	wire x_1511;
	wire x_1512;
	wire x_1513;
	wire x_1514;
	wire x_1515;
	wire x_1516;
	wire x_1517;
	wire x_1518;
	wire x_1519;
	wire x_1520;
	wire x_1521;
	wire x_1522;
	wire x_1523;
	wire x_1524;
	wire x_1525;
	wire x_1526;
	wire x_1527;
	wire x_1528;
	wire x_1529;
	wire x_1530;
	wire x_1531;
	wire x_1532;
	wire x_1533;
	wire x_1534;
	wire x_1535;
	wire x_1536;
	wire x_1537;
	wire x_1538;
	wire x_1539;
	wire x_1540;
	wire x_1541;
	wire x_1542;
	wire x_1543;
	wire x_1544;
	wire x_1545;
	wire x_1546;
	wire x_1547;
	wire x_1548;
	wire x_1549;
	wire x_1550;
	wire x_1551;
	wire x_1552;
	wire x_1553;
	wire x_1554;
	wire x_1555;
	wire x_1556;
	wire x_1557;
	wire x_1558;
	wire x_1559;
	wire x_1560;
	wire x_1561;
	wire x_1562;
	wire x_1563;
	wire x_1564;
	wire x_1565;
	wire x_1566;
	wire x_1567;
	wire x_1568;
	wire x_1569;
	wire x_1570;
	wire x_1571;
	wire x_1572;
	wire x_1573;
	wire x_1574;
	wire x_1575;
	wire x_1576;
	wire x_1577;
	wire x_1578;
	wire x_1579;
	wire x_1580;
	wire x_1581;
	wire x_1582;
	wire x_1583;
	wire x_1584;
	wire x_1585;
	wire x_1586;
	wire x_1587;
	wire x_1588;
	wire x_1589;
	wire x_1590;
	wire x_1591;
	wire x_1592;
	wire x_1593;
	wire x_1594;
	wire x_1595;
	wire x_1596;
	wire x_1597;
	wire x_1598;
	wire x_1599;
	wire x_1600;
	wire x_1601;
	wire x_1602;
	wire x_1603;
	wire x_1604;
	wire x_1605;
	wire x_1606;
	wire x_1607;
	wire x_1608;
	wire x_1609;
	wire x_1610;
	wire x_1611;
	wire x_1612;
	wire x_1613;
	wire x_1614;
	wire x_1615;
	wire x_1616;
	wire x_1617;
	wire x_1618;
	wire x_1619;
	wire x_1620;
	wire x_1621;
	wire x_1622;
	wire x_1623;
	wire x_1624;
	wire x_1625;
	wire x_1626;
	wire x_1627;
	wire x_1628;
	wire x_1629;
	wire x_1630;
	wire x_1631;
	wire x_1632;
	wire x_1633;
	wire x_1634;
	wire x_1635;
	wire x_1636;
	wire x_1637;
	wire x_1638;
	wire x_1639;
	wire x_1640;
	wire x_1641;
	wire x_1642;
	wire x_1643;
	wire x_1644;
	wire x_1645;
	wire x_1646;
	wire x_1647;
	wire x_1648;
	wire x_1649;
	wire x_1650;
	wire x_1651;
	wire x_1652;
	wire x_1653;
	wire x_1654;
	wire x_1655;
	wire x_1656;
	wire x_1657;
	wire x_1658;
	wire x_1659;
	wire x_1660;
	wire x_1661;
	wire x_1662;
	wire x_1663;
	wire x_1664;
	wire x_1665;
	wire x_1666;
	wire x_1667;
	wire x_1668;
	wire x_1669;
	wire x_1670;
	wire x_1671;
	wire x_1672;
	wire x_1673;
	wire x_1674;
	wire x_1675;
	wire x_1676;
	wire x_1677;
	wire x_1678;
	wire x_1679;
	wire x_1680;
	wire x_1681;
	wire x_1682;
	wire x_1683;
	wire x_1684;
	wire x_1685;
	wire x_1686;
	wire x_1687;
	wire x_1688;
	wire x_1689;
	wire x_1690;
	wire x_1691;
	wire x_1692;
	wire x_1693;
	wire x_1694;
	wire x_1695;
	wire x_1696;
	wire x_1697;
	wire x_1698;
	wire x_1699;
	wire x_1700;
	wire x_1701;
	wire x_1702;
	wire x_1703;
	wire x_1704;
	wire x_1705;
	wire x_1706;
	wire x_1707;
	wire x_1708;
	wire x_1709;
	wire x_1710;
	wire x_1711;
	wire x_1712;
	wire x_1713;
	wire x_1714;
	wire x_1715;
	wire x_1716;
	wire x_1717;
	wire x_1718;
	wire x_1719;
	wire x_1720;
	wire x_1721;
	wire x_1722;
	wire x_1723;
	wire x_1724;
	wire x_1725;
	wire x_1726;
	wire x_1727;
	wire x_1728;
	wire x_1729;
	wire x_1730;
	wire x_1731;
	wire x_1732;
	wire x_1733;
	wire x_1734;
	wire x_1735;
	wire x_1736;
	wire x_1737;
	wire x_1738;
	wire x_1739;
	wire x_1740;
	wire x_1741;
	wire x_1742;
	wire x_1743;
	wire x_1744;
	wire x_1745;
	wire x_1746;
	wire x_1747;
	wire x_1748;
	wire x_1749;
	wire x_1750;
	wire x_1751;
	wire x_1752;
	wire x_1753;
	wire x_1754;
	wire x_1755;
	wire x_1756;
	wire x_1757;
	wire x_1758;
	wire x_1759;
	wire x_1760;
	wire x_1761;
	wire x_1762;
	wire x_1763;
	wire x_1764;
	wire x_1765;
	wire x_1766;
	wire x_1767;
	wire x_1768;
	wire x_1769;
	wire x_1770;
	wire x_1771;
	wire x_1772;
	wire x_1773;
	wire x_1774;
	wire x_1775;
	wire x_1776;
	wire x_1777;
	wire x_1778;
	wire x_1779;
	wire x_1780;
	wire x_1781;
	wire x_1782;
	wire x_1783;
	wire x_1784;
	wire x_1785;
	wire x_1786;
	wire x_1787;
	wire x_1788;
	wire x_1789;
	wire x_1790;
	wire x_1791;
	wire x_1792;
	wire x_1793;
	wire x_1794;
	wire x_1795;
	wire x_1796;
	wire x_1797;
	wire x_1798;
	wire x_1799;
	wire x_1800;
	wire x_1801;
	wire x_1802;
	wire x_1803;
	wire x_1804;
	wire x_1805;
	wire x_1806;
	wire x_1807;
	wire x_1808;
	wire x_1809;
	wire x_1810;
	wire x_1811;
	wire x_1812;
	wire x_1813;
	wire x_1814;
	wire x_1815;
	wire x_1816;
	wire x_1817;
	wire x_1818;
	wire x_1819;
	wire x_1820;
	wire x_1821;
	wire x_1822;
	wire x_1823;
	wire x_1824;
	wire x_1825;
	wire x_1826;
	wire x_1827;
	wire x_1828;
	wire x_1829;
	wire x_1830;
	wire x_1831;
	wire x_1832;
	wire x_1833;
	wire x_1834;
	wire x_1835;
	wire x_1836;
	wire x_1837;
	wire x_1838;
	wire x_1839;
	wire x_1840;
	wire x_1841;
	wire x_1842;
	wire x_1843;
	wire x_1844;
	wire x_1845;
	wire x_1846;
	wire x_1847;
	wire x_1848;
	wire x_1849;
	wire x_1850;
	wire x_1851;
	wire x_1852;
	wire x_1853;
	wire x_1854;
	wire x_1855;
	wire x_1856;
	wire x_1857;
	wire x_1858;
	wire x_1859;
	wire x_1860;
	wire x_1861;
	wire x_1862;
	wire x_1863;
	wire x_1864;
	wire x_1865;
	wire x_1866;
	wire x_1867;
	wire x_1868;
	wire x_1869;
	wire x_1870;
	wire x_1871;
	wire x_1872;
	wire x_1873;
	wire x_1874;
	wire x_1875;
	wire x_1876;
	wire x_1877;
	wire x_1878;
	wire x_1879;
	wire x_1880;
	wire x_1881;
	wire x_1882;
	wire x_1883;
	wire x_1884;
	wire x_1885;
	wire x_1886;
	wire x_1887;
	wire x_1888;
	wire x_1889;
	wire x_1890;
	wire x_1891;
	wire x_1892;
	wire x_1893;
	wire x_1894;
	wire x_1895;
	wire x_1896;
	wire x_1897;
	wire x_1898;
	wire x_1899;
	wire x_1900;
	wire x_1901;
	wire x_1902;
	wire x_1903;
	wire x_1904;
	wire x_1905;
	wire x_1906;
	wire x_1907;
	wire x_1908;
	wire x_1909;
	wire x_1910;
	wire x_1911;
	wire x_1912;
	wire x_1913;
	wire x_1914;
	wire x_1915;
	wire x_1916;
	wire x_1917;
	wire x_1918;
	wire x_1919;
	wire x_1920;
	wire x_1921;
	wire x_1922;
	wire x_1923;
	wire x_1924;
	wire x_1925;
	wire x_1926;
	wire x_1927;
	wire x_1928;
	wire x_1929;
	wire x_1930;
	wire x_1931;
	wire x_1932;
	wire x_1933;
	wire x_1934;
	wire x_1935;
	wire x_1936;
	wire x_1937;
	wire x_1938;
	wire x_1939;
	wire x_1940;
	wire x_1941;
	wire x_1942;
	wire x_1943;
	wire x_1944;
	wire x_1945;
	wire x_1946;
	wire x_1947;
	wire x_1948;
	wire x_1949;
	wire x_1950;
	wire x_1951;
	wire x_1952;
	wire x_1953;
	wire x_1954;
	wire x_1955;
	wire x_1956;
	wire x_1957;
	wire x_1958;
	wire x_1959;
	wire x_1960;
	wire x_1961;
	wire x_1962;
	wire x_1963;
	wire x_1964;
	wire x_1965;
	wire x_1966;
	wire x_1967;
	wire x_1968;
	wire x_1969;
	wire x_1970;
	wire x_1971;
	wire x_1972;
	wire x_1973;
	wire x_1974;
	wire x_1975;
	wire x_1976;
	wire x_1977;
	wire x_1978;
	wire x_1979;
	wire x_1980;
	wire x_1981;
	wire x_1982;
	wire x_1983;
	wire x_1984;
	wire x_1985;
	wire x_1986;
	wire x_1987;
	wire x_1988;
	wire x_1989;
	wire x_1990;
	wire x_1991;
	wire x_1992;
	wire x_1993;
	wire x_1994;
	wire x_1995;
	wire x_1996;
	wire x_1997;
	wire x_1998;
	wire x_1999;
	wire x_2000;
	wire x_2001;
	wire x_2002;
	wire x_2003;
	wire x_2004;
	wire x_2005;
	wire x_2006;
	wire x_2007;
	wire x_2008;
	wire x_2009;
	wire x_2010;
	wire x_2011;
	wire x_2012;
	wire x_2013;
	wire x_2014;
	wire x_2015;
	wire x_2016;
	wire x_2017;
	wire x_2018;
	wire x_2019;
	wire x_2020;
	wire x_2021;
	wire x_2022;
	wire x_2023;
	wire x_2024;
	wire x_2025;
	wire x_2026;
	wire x_2027;
	wire x_2028;
	wire x_2029;
	wire x_2030;
	wire x_2031;
	wire x_2032;
	wire x_2033;
	wire x_2034;
	wire x_2035;
	wire x_2036;
	wire x_2037;
	wire x_2038;
	wire x_2039;
	wire x_2040;
	wire x_2041;
	wire x_2042;
	wire x_2043;
	wire x_2044;
	wire x_2045;
	wire x_2046;
	wire x_2047;
	wire x_2048;
	wire x_2049;
	wire x_2050;
	wire x_2051;
	wire x_2052;
	wire x_2053;
	wire x_2054;
	wire x_2055;
	wire x_2056;
	wire x_2057;
	wire x_2058;
	wire x_2059;
	wire x_2060;
	wire x_2061;
	wire x_2062;
	wire x_2063;
	wire x_2064;
	wire x_2065;
	wire x_2066;
	wire x_2067;
	wire x_2068;
	wire x_2069;
	wire x_2070;
	wire x_2071;
	wire x_2072;
	wire x_2073;
	wire x_2074;
	wire x_2075;
	wire x_2076;
	wire x_2077;
	wire x_2078;
	wire x_2079;
	wire x_2080;
	wire x_2081;
	wire x_2082;
	wire x_2083;
	wire x_2084;
	wire x_2085;
	wire x_2086;
	wire x_2087;
	wire x_2088;
	wire x_2089;
	wire x_2090;
	wire x_2091;
	wire x_2092;
	wire x_2093;
	wire x_2094;
	wire x_2095;
	wire x_2096;
	wire x_2097;
	wire x_2098;
	wire x_2099;
	wire x_2100;
	wire x_2101;
	wire x_2102;
	wire x_2103;
	wire x_2104;
	wire x_2105;
	wire x_2106;
	wire x_2107;
	wire x_2108;
	wire x_2109;
	wire x_2110;
	wire x_2111;
	wire x_2112;
	wire x_2113;
	wire x_2114;
	wire x_2115;
	wire x_2116;
	wire x_2117;
	wire x_2118;
	wire x_2119;
	wire x_2120;
	wire x_2121;
	wire x_2122;
	wire x_2123;
	wire x_2124;
	wire x_2125;
	wire x_2126;
	wire x_2127;
	wire x_2128;
	wire x_2129;
	wire x_2130;
	wire x_2131;
	wire x_2132;
	wire x_2133;
	wire x_2134;
	wire x_2135;
	wire x_2136;
	wire x_2137;
	wire x_2138;
	wire x_2139;
	wire x_2140;
	wire x_2141;
	wire x_2142;
	wire x_2143;
	wire x_2144;
	wire x_2145;
	wire x_2146;
	wire x_2147;
	wire x_2148;
	wire x_2149;
	wire x_2150;
	wire x_2151;
	wire x_2152;
	wire x_2153;
	wire x_2154;
	wire x_2155;
	wire x_2156;
	wire x_2157;
	wire x_2158;
	wire x_2159;
	wire x_2160;
	wire x_2161;
	wire x_2162;
	wire x_2163;
	wire x_2164;
	wire x_2165;
	wire x_2166;
	wire x_2167;
	wire x_2168;
	wire x_2169;
	wire x_2170;
	wire x_2171;
	wire x_2172;
	wire x_2173;
	wire x_2174;
	wire x_2175;
	wire x_2176;
	wire x_2177;
	wire x_2178;
	wire x_2179;
	wire x_2180;
	wire x_2181;
	wire x_2182;
	wire x_2183;
	wire x_2184;
	wire x_2185;
	wire x_2186;
	wire x_2187;
	wire x_2188;
	wire x_2189;
	wire x_2190;
	wire x_2191;
	wire x_2192;
	wire x_2193;
	wire x_2194;
	wire x_2195;
	wire x_2196;
	wire x_2197;
	wire x_2198;
	wire x_2199;
	wire x_2200;
	wire x_2201;
	wire x_2202;
	wire x_2203;
	wire x_2204;
	wire x_2205;
	wire x_2206;
	wire x_2207;
	wire x_2208;
	wire x_2209;
	wire x_2210;
	wire x_2211;
	wire x_2212;
	wire x_2213;
	wire x_2214;
	wire x_2215;
	wire x_2216;
	wire x_2217;
	wire x_2218;
	wire x_2219;
	wire x_2220;
	wire x_2221;
	wire x_2222;
	wire x_2223;
	wire x_2224;
	wire x_2225;
	wire x_2226;
	wire x_2227;
	wire x_2228;
	wire x_2229;
	wire x_2230;
	wire x_2231;
	wire x_2232;
	wire x_2233;
	wire x_2234;
	wire x_2235;
	wire x_2236;
	wire x_2237;
	wire x_2238;
	wire x_2239;
	wire x_2240;
	wire x_2241;
	wire x_2242;
	wire x_2243;
	wire x_2244;
	wire x_2245;
	wire x_2246;
	wire x_2247;
	wire x_2248;
	wire x_2249;
	wire x_2250;
	wire x_2251;
	wire x_2252;
	wire x_2253;
	wire x_2254;
	wire x_2255;
	wire x_2256;
	wire x_2257;
	wire x_2258;
	wire x_2259;
	wire x_2260;
	wire x_2261;
	wire x_2262;
	wire x_2263;
	wire x_2264;
	wire x_2265;
	wire x_2266;
	wire x_2267;
	wire x_2268;
	wire x_2269;
	wire x_2270;
	wire x_2271;
	wire x_2272;
	wire x_2273;
	wire x_2274;
	wire x_2275;
	wire x_2276;
	wire x_2277;
	wire x_2278;
	wire x_2279;
	wire x_2280;
	wire x_2281;
	wire x_2282;
	wire x_2283;
	wire x_2284;
	wire x_2285;
	wire x_2286;
	wire x_2287;
	wire x_2288;
	wire x_2289;
	wire x_2290;
	wire x_2291;
	wire x_2292;
	wire x_2293;
	wire x_2294;
	wire x_2295;
	wire x_2296;
	wire x_2297;
	wire x_2298;
	wire x_2299;
	wire x_2300;
	wire x_2301;
	wire x_2302;
	wire x_2303;
	wire x_2304;
	wire x_2305;
	wire x_2306;
	wire x_2307;
	wire x_2308;
	wire x_2309;
	wire x_2310;
	wire x_2311;
	wire x_2312;
	wire x_2313;
	wire x_2314;
	wire x_2315;
	wire x_2316;
	wire x_2317;
	wire x_2318;
	wire x_2319;
	wire x_2320;
	wire x_2321;
	wire x_2322;
	wire x_2323;
	wire x_2324;
	wire x_2325;
	wire x_2326;
	wire x_2327;
	wire x_2328;
	wire x_2329;
	wire x_2330;
	wire x_2331;
	wire x_2332;
	wire x_2333;
	wire x_2334;
	wire x_2335;
	wire x_2336;
	wire x_2337;
	wire x_2338;
	wire x_2339;
	wire x_2340;
	wire x_2341;
	wire x_2342;
	wire x_2343;
	wire x_2344;
	wire x_2345;
	wire x_2346;
	wire x_2347;
	wire x_2348;
	wire x_2349;
	wire x_2350;
	wire x_2351;
	wire x_2352;
	wire x_2353;
	wire x_2354;
	wire x_2355;
	wire x_2356;
	wire x_2357;
	wire x_2358;
	wire x_2359;
	wire x_2360;
	wire x_2361;
	wire x_2362;
	wire x_2363;
	wire x_2364;
	wire x_2365;
	wire x_2366;
	wire x_2367;
	wire x_2368;
	wire x_2369;
	wire x_2370;
	wire x_2371;
	wire x_2372;
	wire x_2373;
	wire x_2374;
	wire x_2375;
	wire x_2376;
	wire x_2377;
	wire x_2378;
	wire x_2379;
	wire x_2380;
	wire x_2381;
	wire x_2382;
	wire x_2383;
	wire x_2384;
	wire x_2385;
	wire x_2386;
	wire x_2387;
	wire x_2388;
	wire x_2389;
	wire x_2390;
	wire x_2391;
	wire x_2392;
	wire x_2393;
	wire x_2394;
	wire x_2395;
	wire x_2396;
	wire x_2397;
	wire x_2398;
	wire x_2399;
	wire x_2400;
	wire x_2401;
	wire x_2402;
	wire x_2403;
	wire x_2404;
	wire x_2405;
	wire x_2406;
	wire x_2407;
	wire x_2408;
	wire x_2409;
	wire x_2410;
	wire x_2411;
	wire x_2412;
	wire x_2413;
	wire x_2414;
	wire x_2415;
	wire x_2416;
	wire x_2417;
	wire x_2418;
	wire x_2419;
	wire x_2420;
	wire x_2421;
	wire x_2422;
	wire x_2423;
	wire x_2424;
	wire x_2425;
	wire x_2426;
	wire x_2427;
	wire x_2428;
	wire x_2429;
	wire x_2430;
	wire x_2431;
	wire x_2432;
	wire x_2433;
	wire x_2434;
	wire x_2435;
	wire x_2436;
	wire x_2437;
	wire x_2438;
	wire x_2439;
	wire x_2440;
	wire x_2441;
	wire x_2442;
	wire x_2443;
	wire x_2444;
	wire x_2445;
	wire x_2446;
	wire x_2447;
	wire x_2448;
	wire x_2449;
	wire x_2450;
	wire x_2451;
	wire x_2452;
	wire x_2453;
	wire x_2454;
	wire x_2455;
	wire x_2456;
	wire x_2457;
	wire x_2458;
	wire x_2459;
	wire x_2460;
	wire x_2461;
	wire x_2462;
	wire x_2463;
	wire x_2464;
	wire x_2465;
	wire x_2466;
	wire x_2467;
	wire x_2468;
	wire x_2469;
	wire x_2470;
	wire x_2471;
	wire x_2472;
	wire x_2473;
	wire x_2474;
	wire x_2475;
	wire x_2476;
	wire x_2477;
	wire x_2478;
	wire x_2479;
	wire x_2480;
	wire x_2481;
	wire x_2482;
	wire x_2483;
	wire x_2484;
	wire x_2485;
	wire x_2486;
	wire x_2487;
	wire x_2488;
	wire x_2489;
	wire x_2490;
	wire x_2491;
	wire x_2492;
	wire x_2493;
	wire x_2494;
	wire x_2495;
	wire x_2496;
	wire x_2497;
	wire x_2498;
	wire x_2499;
	wire x_2500;
	wire x_2501;
	wire x_2502;
	wire x_2503;
	wire x_2504;
	wire x_2505;
	wire x_2506;
	wire x_2507;
	wire x_2508;
	wire x_2509;
	wire x_2510;
	wire x_2511;
	wire x_2512;
	wire x_2513;
	wire x_2514;
	wire x_2515;
	wire x_2516;
	wire x_2517;
	wire x_2518;
	wire x_2519;
	wire x_2520;
	wire x_2521;
	wire x_2522;
	wire x_2523;
	wire x_2524;
	wire x_2525;
	wire x_2526;
	wire x_2527;
	wire x_2528;
	wire x_2529;
	wire x_2530;
	wire x_2531;
	wire x_2532;
	wire x_2533;
	wire x_2534;
	wire x_2535;
	wire x_2536;
	wire x_2537;
	wire x_2538;
	wire x_2539;
	wire x_2540;
	wire x_2541;
	wire x_2542;
	wire x_2543;
	wire x_2544;
	wire x_2545;
	wire x_2546;
	wire x_2547;
	wire x_2548;
	wire x_2549;
	wire x_2550;
	wire x_2551;
	wire x_2552;
	wire x_2553;
	wire x_2554;
	wire x_2555;
	wire x_2556;
	wire x_2557;
	wire x_2558;
	wire x_2559;
	wire x_2560;
	wire x_2561;
	wire x_2562;
	wire x_2563;
	wire x_2564;
	wire x_2565;
	wire x_2566;
	wire x_2567;
	wire x_2568;
	wire x_2569;
	wire x_2570;
	wire x_2571;
	wire x_2572;
	wire x_2573;
	wire x_2574;
	wire x_2575;
	wire x_2576;
	wire x_2577;
	wire x_2578;
	wire x_2579;
	wire x_2580;
	wire x_2581;
	wire x_2582;
	wire x_2583;
	wire x_2584;
	wire x_2585;
	wire x_2586;
	wire x_2587;
	wire x_2588;
	wire x_2589;
	wire x_2590;
	wire x_2591;
	wire x_2592;
	wire x_2593;
	wire x_2594;
	wire x_2595;
	wire x_2596;
	wire x_2597;
	wire x_2598;
	wire x_2599;
	wire x_2600;
	wire x_2601;
	wire x_2602;
	wire x_2603;
	wire x_2604;
	wire x_2605;
	wire x_2606;
	wire x_2607;
	wire x_2608;
	wire x_2609;
	wire x_2610;
	wire x_2611;
	wire x_2612;
	wire x_2613;
	wire x_2614;
	wire x_2615;
	wire x_2616;
	wire x_2617;
	wire x_2618;
	wire x_2619;
	wire x_2620;
	wire x_2621;
	wire x_2622;
	wire x_2623;
	wire x_2624;
	wire x_2625;
	wire x_2626;
	wire x_2627;
	wire x_2628;
	wire x_2629;
	wire x_2630;
	wire x_2631;
	wire x_2632;
	wire x_2633;
	wire x_2634;
	wire x_2635;
	wire x_2636;
	wire x_2637;
	wire x_2638;
	wire x_2639;
	wire x_2640;
	wire x_2641;
	wire x_2642;
	wire x_2643;
	wire x_2644;
	wire x_2645;
	wire x_2646;
	wire x_2647;
	wire x_2648;
	wire x_2649;
	wire x_2650;
	wire x_2651;
	wire x_2652;
	wire x_2653;
	wire x_2654;
	wire x_2655;
	wire x_2656;
	wire x_2657;
	wire x_2658;
	wire x_2659;
	wire x_2660;
	wire x_2661;
	wire x_2662;
	wire x_2663;
	wire x_2664;
	wire x_2665;
	wire x_2666;
	wire x_2667;
	wire x_2668;
	wire x_2669;
	wire x_2670;
	wire x_2671;
	wire x_2672;
	wire x_2673;
	wire x_2674;
	wire x_2675;
	wire x_2676;
	wire x_2677;
	wire x_2678;
	wire x_2679;
	wire x_2680;
	wire x_2681;
	wire x_2682;
	wire x_2683;
	wire x_2684;
	wire x_2685;
	wire x_2686;
	wire x_2687;
	wire x_2688;
	wire x_2689;
	wire x_2690;
	wire x_2691;
	wire x_2692;
	wire x_2693;
	wire x_2694;
	wire x_2695;
	wire x_2696;
	wire x_2697;
	wire x_2698;
	wire x_2699;
	wire x_2700;
	wire x_2701;
	wire x_2702;
	wire x_2703;
	wire x_2704;
	wire x_2705;
	wire x_2706;
	wire x_2707;
	wire x_2708;
	wire x_2709;
	wire x_2710;
	wire x_2711;
	wire x_2712;
	wire x_2713;
	wire x_2714;
	wire x_2715;
	wire x_2716;
	wire x_2717;
	wire x_2718;
	wire x_2719;
	wire x_2720;
	wire x_2721;
	wire x_2722;
	wire x_2723;
	wire x_2724;
	wire x_2725;
	wire x_2726;
	wire x_2727;
	wire x_2728;
	wire x_2729;
	wire x_2730;
	wire x_2731;
	wire x_2732;
	wire x_2733;
	wire x_2734;
	wire x_2735;
	wire x_2736;
	wire x_2737;
	wire x_2738;
	wire x_2739;
	wire x_2740;
	wire x_2741;
	wire x_2742;
	wire x_2743;
	wire x_2744;
	wire x_2745;
	wire x_2746;
	wire x_2747;
	wire x_2748;
	wire x_2749;
	wire x_2750;
	wire x_2751;
	wire x_2752;
	wire x_2753;
	wire x_2754;
	wire x_2755;
	wire x_2756;
	wire x_2757;
	wire x_2758;
	wire x_2759;
	wire x_2760;
	wire x_2761;
	wire x_2762;
	wire x_2763;
	wire x_2764;
	wire x_2765;
	wire x_2766;
	wire x_2767;
	wire x_2768;
	wire x_2769;
	wire x_2770;
	wire x_2771;
	wire x_2772;
	wire x_2773;
	wire x_2774;
	wire x_2775;
	wire x_2776;
	wire x_2777;
	wire x_2778;
	wire x_2779;
	wire x_2780;
	wire x_2781;
	wire x_2782;
	wire x_2783;
	wire x_2784;
	wire x_2785;
	wire x_2786;
	wire x_2787;
	wire x_2788;
	wire x_2789;
	wire x_2790;
	wire x_2791;
	wire x_2792;
	wire x_2793;
	wire x_2794;
	wire x_2795;
	wire x_2796;
	wire x_2797;
	wire x_2798;
	wire x_2799;
	wire x_2800;
	wire x_2801;
	wire x_2802;
	wire x_2803;
	wire x_2804;
	wire x_2805;
	wire x_2806;
	wire x_2807;
	wire x_2808;
	wire x_2809;
	wire x_2810;
	wire x_2811;
	wire x_2812;
	wire x_2813;
	wire x_2814;
	wire x_2815;
	wire x_2816;
	wire x_2817;
	wire x_2818;
	wire x_2819;
	wire x_2820;
	wire x_2821;
	wire x_2822;
	wire x_2823;
	wire x_2824;
	wire x_2825;
	wire x_2826;
	wire x_2827;
	wire x_2828;
	wire x_2829;
	wire x_2830;
	wire x_2831;
	wire x_2832;
	wire x_2833;
	wire x_2834;
	wire x_2835;
	wire x_2836;
	wire x_2837;
	wire x_2838;
	wire x_2839;
	wire x_2840;
	wire x_2841;
	wire x_2842;
	wire x_2843;
	wire x_2844;
	wire x_2845;
	wire x_2846;
	wire x_2847;
	wire x_2848;
	wire x_2849;
	wire x_2850;
	wire x_2851;
	wire x_2852;
	wire x_2853;
	wire x_2854;
	wire x_2855;
	wire x_2856;
	wire x_2857;
	wire x_2858;
	wire x_2859;
	wire x_2860;
	wire x_2861;
	wire x_2862;
	wire x_2863;
	wire x_2864;
	wire x_2865;
	wire x_2866;
	wire x_2867;
	wire x_2868;
	wire x_2869;
	wire x_2870;
	wire x_2871;
	wire x_2872;
	wire x_2873;
	wire x_2874;
	wire x_2875;
	wire x_2876;
	wire x_2877;
	wire x_2878;
	wire x_2879;
	wire x_2880;
	wire x_2881;
	wire x_2882;
	wire x_2883;
	wire x_2884;
	wire x_2885;
	wire x_2886;
	wire x_2887;
	wire x_2888;
	wire x_2889;
	wire x_2890;
	wire x_2891;
	wire x_2892;
	wire x_2893;
	wire x_2894;
	wire x_2895;
	wire x_2896;
	wire x_2897;
	wire x_2898;
	wire x_2899;
	wire x_2900;
	wire x_2901;
	wire x_2902;
	wire x_2903;
	wire x_2904;
	wire x_2905;
	wire x_2906;
	wire x_2907;
	wire x_2908;
	wire x_2909;
	wire x_2910;
	wire x_2911;
	wire x_2912;
	wire x_2913;
	wire x_2914;
	wire x_2915;
	wire x_2916;
	wire x_2917;
	wire x_2918;
	wire x_2919;
	wire x_2920;
	wire x_2921;
	wire x_2922;
	wire x_2923;
	wire x_2924;
	wire x_2925;
	wire x_2926;
	wire x_2927;
	wire x_2928;
	wire x_2929;
	wire x_2930;
	wire x_2931;
	wire x_2932;
	wire x_2933;
	wire x_2934;
	wire x_2935;
	wire x_2936;
	wire x_2937;
	wire x_2938;
	wire x_2939;
	wire x_2940;
	wire x_2941;
	wire x_2942;
	wire x_2943;
	wire x_2944;
	wire x_2945;
	wire x_2946;
	wire x_2947;
	wire x_2948;
	wire x_2949;
	wire x_2950;
	wire x_2951;
	wire x_2952;
	wire x_2953;
	wire x_2954;
	wire x_2955;
	wire x_2956;
	wire x_2957;
	wire x_2958;
	wire x_2959;
	wire x_2960;
	wire x_2961;
	wire x_2962;
	wire x_2963;
	wire x_2964;
	wire x_2965;
	wire x_2966;
	wire x_2967;
	wire x_2968;
	wire x_2969;
	wire x_2970;
	wire x_2971;
	wire x_2972;
	wire x_2973;
	wire x_2974;
	wire x_2975;
	wire x_2976;
	wire x_2977;
	wire x_2978;
	wire x_2979;
	wire x_2980;
	wire x_2981;
	wire x_2982;
	wire x_2983;
	wire x_2984;
	wire x_2985;
	wire x_2986;
	wire x_2987;
	wire x_2988;
	wire x_2989;
	wire x_2990;
	wire x_2991;
	wire x_2992;
	wire x_2993;
	wire x_2994;
	wire x_2995;
	wire x_2996;
	wire x_2997;
	wire x_2998;
	wire x_2999;
	wire x_3000;
	wire x_3001;
	wire x_3002;
	wire x_3003;
	wire x_3004;
	wire x_3005;
	wire x_3006;
	wire x_3007;
	wire x_3008;
	wire x_3009;
	wire x_3010;
	wire x_3011;
	wire x_3012;
	wire x_3013;
	wire x_3014;
	wire x_3015;
	wire x_3016;
	wire x_3017;
	wire x_3018;
	wire x_3019;
	wire x_3020;
	wire x_3021;
	wire x_3022;
	wire x_3023;
	wire x_3024;
	wire x_3025;
	wire x_3026;
	wire x_3027;
	wire x_3028;
	wire x_3029;
	wire x_3030;
	wire x_3031;
	wire x_3032;
	wire x_3033;
	wire x_3034;
	wire x_3035;
	wire x_3036;
	wire x_3037;
	wire x_3038;
	wire x_3039;
	wire x_3040;
	wire x_3041;
	wire x_3042;
	wire x_3043;
	wire x_3044;
	wire x_3045;
	wire x_3046;
	wire x_3047;
	wire x_3048;
	wire x_3049;
	wire x_3050;
	wire x_3051;
	wire x_3052;
	wire x_3053;
	wire x_3054;
	wire x_3055;
	wire x_3056;
	wire x_3057;
	wire x_3058;
	wire x_3059;
	wire x_3060;
	wire x_3061;
	wire x_3062;
	wire x_3063;
	wire x_3064;
	wire x_3065;
	wire x_3066;
	wire x_3067;
	wire x_3068;
	wire x_3069;
	wire x_3070;
	wire x_3071;
	wire x_3072;
	wire x_3073;
	wire x_3074;
	wire x_3075;
	wire x_3076;
	wire x_3077;
	wire x_3078;
	wire x_3079;
	wire x_3080;
	wire x_3081;
	wire x_3082;
	wire x_3083;
	wire x_3084;
	wire x_3085;
	wire x_3086;
	wire x_3087;
	wire x_3088;
	wire x_3089;
	wire x_3090;
	wire x_3091;
	wire x_3092;
	wire x_3093;
	wire x_3094;
	wire x_3095;
	wire x_3096;
	wire x_3097;
	wire x_3098;
	wire x_3099;
	wire x_3100;
	wire x_3101;
	wire x_3102;
	wire x_3103;
	wire x_3104;
	wire x_3105;
	wire x_3106;
	wire x_3107;
	wire x_3108;
	wire x_3109;
	wire x_3110;
	wire x_3111;
	wire x_3112;
	wire x_3113;
	wire x_3114;
	wire x_3115;
	wire x_3116;
	wire x_3117;
	wire x_3118;
	wire x_3119;
	wire x_3120;
	wire x_3121;
	wire x_3122;
	wire x_3123;
	wire x_3124;
	wire x_3125;
	wire x_3126;
	wire x_3127;
	wire x_3128;
	wire x_3129;
	wire x_3130;
	wire x_3131;
	wire x_3132;
	wire x_3133;
	wire x_3134;
	wire x_3135;
	wire x_3136;
	wire x_3137;
	wire x_3138;
	wire x_3139;
	wire x_3140;
	wire x_3141;
	wire x_3142;
	wire x_3143;
	wire x_3144;
	wire x_3145;
	wire x_3146;
	wire x_3147;
	wire x_3148;
	wire x_3149;
	wire x_3150;
	wire x_3151;
	wire x_3152;
	wire x_3153;
	wire x_3154;
	wire x_3155;
	wire x_3156;
	wire x_3157;
	wire x_3158;
	wire x_3159;
	wire x_3160;
	wire x_3161;
	wire x_3162;
	wire x_3163;
	wire x_3164;
	wire x_3165;
	wire x_3166;
	wire x_3167;
	wire x_3168;
	wire x_3169;
	wire x_3170;
	wire x_3171;
	wire x_3172;
	wire x_3173;
	wire x_3174;
	wire x_3175;
	wire x_3176;
	wire x_3177;
	wire x_3178;
	wire x_3179;
	wire x_3180;
	wire x_3181;
	wire x_3182;
	wire x_3183;
	wire x_3184;
	wire x_3185;
	wire x_3186;
	wire x_3187;
	wire x_3188;
	wire x_3189;
	wire x_3190;
	wire x_3191;
	wire x_3192;
	wire x_3193;
	wire x_3194;
	wire x_3195;
	wire x_3196;
	wire x_3197;
	wire x_3198;
	wire x_3199;
	wire x_3200;
	wire x_3201;
	wire x_3202;
	wire x_3203;
	wire x_3204;
	wire x_3205;
	wire x_3206;
	wire x_3207;
	wire x_3208;
	wire x_3209;
	wire x_3210;
	wire x_3211;
	wire x_3212;
	wire x_3213;
	wire x_3214;
	wire x_3215;
	wire x_3216;
	wire x_3217;
	wire x_3218;
	wire x_3219;
	wire x_3220;
	wire x_3221;
	wire x_3222;
	wire x_3223;
	wire x_3224;
	wire x_3225;
	wire x_3226;
	wire x_3227;
	wire x_3228;
	wire x_3229;
	wire x_3230;
	wire x_3231;
	wire x_3232;
	wire x_3233;
	wire x_3234;
	wire x_3235;
	wire x_3236;
	wire x_3237;
	wire x_3238;
	wire x_3239;
	wire x_3240;
	wire x_3241;
	wire x_3242;
	wire x_3243;
	wire x_3244;
	wire x_3245;
	wire x_3246;
	wire x_3247;
	wire x_3248;
	wire x_3249;
	wire x_3250;
	wire x_3251;
	wire x_3252;
	wire x_3253;
	wire x_3254;
	wire x_3255;
	wire x_3256;
	wire x_3257;
	wire x_3258;
	wire x_3259;
	wire x_3260;
	wire x_3261;
	wire x_3262;
	wire x_3263;
	wire x_3264;
	wire x_3265;
	wire x_3266;
	wire x_3267;
	wire x_3268;
	wire x_3269;
	wire x_3270;
	wire x_3271;
	wire x_3272;
	wire x_3273;
	wire x_3274;
	wire x_3275;
	wire x_3276;
	wire x_3277;
	wire x_3278;
	wire x_3279;
	wire x_3280;
	wire x_3281;
	wire x_3282;
	wire x_3283;
	wire x_3284;
	wire x_3285;
	wire x_3286;
	wire x_3287;
	wire x_3288;
	wire x_3289;
	wire x_3290;
	wire x_3291;
	wire x_3292;
	wire x_3293;
	wire x_3294;
	wire x_3295;
	wire x_3296;
	wire x_3297;
	wire x_3298;
	wire x_3299;
	wire x_3300;
	wire x_3301;
	wire x_3302;
	wire x_3303;
	wire x_3304;
	wire x_3305;
	wire x_3306;
	wire x_3307;
	wire x_3308;
	wire x_3309;
	wire x_3310;
	wire x_3311;
	wire x_3312;
	wire x_3313;
	wire x_3314;
	wire x_3315;
	wire x_3316;
	wire x_3317;
	wire x_3318;
	wire x_3319;
	wire x_3320;
	wire x_3321;
	wire x_3322;
	wire x_3323;
	wire x_3324;
	wire x_3325;
	wire x_3326;
	wire x_3327;
	wire x_3328;
	wire x_3329;
	wire x_3330;
	wire x_3331;
	wire x_3332;
	wire x_3333;
	wire x_3334;
	wire x_3335;
	wire x_3336;
	wire x_3337;
	wire x_3338;
	wire x_3339;
	wire x_3340;
	wire x_3341;
	wire x_3342;
	wire x_3343;
	wire x_3344;
	wire x_3345;
	wire x_3346;
	wire x_3347;
	wire x_3348;
	wire x_3349;
	wire x_3350;
	wire x_3351;
	wire x_3352;
	wire x_3353;
	wire x_3354;
	wire x_3355;
	wire x_3356;
	wire x_3357;
	wire x_3358;
	wire x_3359;
	wire x_3360;
	wire x_3361;
	wire x_3362;
	wire x_3363;
	wire x_3364;
	wire x_3365;
	wire x_3366;
	wire x_3367;
	wire x_3368;
	wire x_3369;
	wire x_3370;
	wire x_3371;
	wire x_3372;
	wire x_3373;
	wire x_3374;
	wire x_3375;
	wire x_3376;
	wire x_3377;
	wire x_3378;
	wire x_3379;
	wire x_3380;
	wire x_3381;
	wire x_3382;
	wire x_3383;
	wire x_3384;
	wire x_3385;
	wire x_3386;
	wire x_3387;
	wire x_3388;
	wire x_3389;
	wire x_3390;
	wire x_3391;
	wire x_3392;
	wire x_3393;
	wire x_3394;
	wire x_3395;
	wire x_3396;
	wire x_3397;
	wire x_3398;
	wire x_3399;
	wire x_3400;
	wire x_3401;
	wire x_3402;
	wire x_3403;
	wire x_3404;
	wire x_3405;
	wire x_3406;
	wire x_3407;
	wire x_3408;
	wire x_3409;
	wire x_3410;
	wire x_3411;
	wire x_3412;
	wire x_3413;
	wire x_3414;
	wire x_3415;
	wire x_3416;
	wire x_3417;
	wire x_3418;
	wire x_3419;
	wire x_3420;
	wire x_3421;
	wire x_3422;
	wire x_3423;
	wire x_3424;
	wire x_3425;
	wire x_3426;
	wire x_3427;
	wire x_3428;
	wire x_3429;
	wire x_3430;
	wire x_3431;
	wire x_3432;
	wire x_3433;
	wire x_3434;
	wire x_3435;
	wire x_3436;
	wire x_3437;
	wire x_3438;
	wire x_3439;
	wire x_3440;
	wire x_3441;
	wire x_3442;
	wire x_3443;
	wire x_3444;
	wire x_3445;
	wire x_3446;
	wire x_3447;
	wire x_3448;
	wire x_3449;
	wire x_3450;
	wire x_3451;
	wire x_3452;
	wire x_3453;
	wire x_3454;
	wire x_3455;
	wire x_3456;
	wire x_3457;
	wire x_3458;
	wire x_3459;
	wire x_3460;
	wire x_3461;
	wire x_3462;
	wire x_3463;
	wire x_3464;
	wire x_3465;
	wire x_3466;
	wire x_3467;
	wire x_3468;
	wire x_3469;
	wire x_3470;
	wire x_3471;
	wire x_3472;
	wire x_3473;
	wire x_3474;
	wire x_3475;
	wire x_3476;
	wire x_3477;
	wire x_3478;
	wire x_3479;
	wire x_3480;
	wire x_3481;
	wire x_3482;
	wire x_3483;
	wire x_3484;
	wire x_3485;
	wire x_3486;
	wire x_3487;
	wire x_3488;
	wire x_3489;
	wire x_3490;
	wire x_3491;
	wire x_3492;
	wire x_3493;
	wire x_3494;
	wire x_3495;
	wire x_3496;
	wire x_3497;
	wire x_3498;
	wire x_3499;
	wire x_3500;
	wire x_3501;
	wire x_3502;
	wire x_3503;
	wire x_3504;
	wire x_3505;
	wire x_3506;
	wire x_3507;
	wire x_3508;
	wire x_3509;
	wire x_3510;
	wire x_3511;
	wire x_3512;
	wire x_3513;
	wire x_3514;
	wire x_3515;
	wire x_3516;
	wire x_3517;
	wire x_3518;
	wire x_3519;
	wire x_3520;
	wire x_3521;
	wire x_3522;
	wire x_3523;
	wire x_3524;
	wire x_3525;
	wire x_3526;
	wire x_3527;
	wire x_3528;
	wire x_3529;
	wire x_3530;
	wire x_3531;
	wire x_3532;
	wire x_3533;
	wire x_3534;
	wire x_3535;
	wire x_3536;
	wire x_3537;
	wire x_3538;
	wire x_3539;
	wire x_3540;
	wire x_3541;
	wire x_3542;
	wire x_3543;
	wire x_3544;
	wire x_3545;
	wire x_3546;
	wire x_3547;
	wire x_3548;
	wire x_3549;
	wire x_3550;
	wire x_3551;
	wire x_3552;
	wire x_3553;
	wire x_3554;
	wire x_3555;
	wire x_3556;
	wire x_3557;
	wire x_3558;
	wire x_3559;
	wire x_3560;
	wire x_3561;
	wire x_3562;
	wire x_3563;
	wire x_3564;
	wire x_3565;
	wire x_3566;
	wire x_3567;
	wire x_3568;
	wire x_3569;
	wire x_3570;
	wire x_3571;
	wire x_3572;
	wire x_3573;
	wire x_3574;
	wire x_3575;
	wire x_3576;
	wire x_3577;
	wire x_3578;
	wire x_3579;
	wire x_3580;
	wire x_3581;
	wire x_3582;
	wire x_3583;
	wire x_3584;
	wire x_3585;
	wire x_3586;
	wire x_3587;
	wire x_3588;
	wire x_3589;
	wire x_3590;
	wire x_3591;
	wire x_3592;
	wire x_3593;
	wire x_3594;
	wire x_3595;
	wire x_3596;
	wire x_3597;
	wire x_3598;
	wire x_3599;
	wire x_3600;
	wire x_3601;
	wire x_3602;
	wire x_3603;
	wire x_3604;
	wire x_3605;
	wire x_3606;
	wire x_3607;
	wire x_3608;
	wire x_3609;
	wire x_3610;
	wire x_3611;
	wire x_3612;
	wire x_3613;
	wire x_3614;
	wire x_3615;
	wire x_3616;
	wire x_3617;
	wire x_3618;
	wire x_3619;
	wire x_3620;
	wire x_3621;
	wire x_3622;
	wire x_3623;
	wire x_3624;
	wire x_3625;
	wire x_3626;
	wire x_3627;
	wire x_3628;
	wire x_3629;
	wire x_3630;
	wire x_3631;
	wire x_3632;
	wire x_3633;
	wire x_3634;
	wire x_3635;
	wire x_3636;
	wire x_3637;
	wire x_3638;
	wire x_3639;
	wire x_3640;
	wire x_3641;
	wire x_3642;
	wire x_3643;
	wire x_3644;
	wire x_3645;
	wire x_3646;
	wire x_3647;
	wire x_3648;
	wire x_3649;
	wire x_3650;
	wire x_3651;
	wire x_3652;
	wire x_3653;
	wire x_3654;
	wire x_3655;
	wire x_3656;
	wire x_3657;
	wire x_3658;
	wire x_3659;
	wire x_3660;
	wire x_3661;
	wire x_3662;
	wire x_3663;
	wire x_3664;
	wire x_3665;
	wire x_3666;
	wire x_3667;
	wire x_3668;
	wire x_3669;
	wire x_3670;
	wire x_3671;
	wire x_3672;
	wire x_3673;
	wire x_3674;
	wire x_3675;
	wire x_3676;
	wire x_3677;
	wire x_3678;
	wire x_3679;
	wire x_3680;
	wire x_3681;
	wire x_3682;
	wire x_3683;
	wire x_3684;
	wire x_3685;
	wire x_3686;
	wire x_3687;
	wire x_3688;
	wire x_3689;
	wire x_3690;
	wire x_3691;
	wire x_3692;
	wire x_3693;
	wire x_3694;
	wire x_3695;
	wire x_3696;
	wire x_3697;
	wire x_3698;
	wire x_3699;
	wire x_3700;
	wire x_3701;
	wire x_3702;
	wire x_3703;
	wire x_3704;
	wire x_3705;
	wire x_3706;
	wire x_3707;
	wire x_3708;
	wire x_3709;
	wire x_3710;
	wire x_3711;
	wire x_3712;
	wire x_3713;
	wire x_3714;
	wire x_3715;
	wire x_3716;
	wire x_3717;
	wire x_3718;
	wire x_3719;
	wire x_3720;
	wire x_3721;
	wire x_3722;
	wire x_3723;
	wire x_3724;
	wire x_3725;
	wire x_3726;
	wire x_3727;
	wire x_3728;
	wire x_3729;
	wire x_3730;
	wire x_3731;
	wire x_3732;
	wire x_3733;
	wire x_3734;
	wire x_3735;
	wire x_3736;
	wire x_3737;
	wire x_3738;
	wire x_3739;
	wire x_3740;
	wire x_3741;
	wire x_3742;
	wire x_3743;
	wire x_3744;
	wire x_3745;
	wire x_3746;
	wire x_3747;
	wire x_3748;
	wire x_3749;
	wire x_3750;
	wire x_3751;
	wire x_3752;
	wire x_3753;
	wire x_3754;
	wire x_3755;
	wire x_3756;
	wire x_3757;
	wire x_3758;
	wire x_3759;
	wire x_3760;
	wire x_3761;
	wire x_3762;
	wire x_3763;
	wire x_3764;
	wire x_3765;
	wire x_3766;
	wire x_3767;
	wire x_3768;
	wire x_3769;
	wire x_3770;
	wire x_3771;
	wire x_3772;
	wire x_3773;
	wire x_3774;
	wire x_3775;
	wire x_3776;
	wire x_3777;
	wire x_3778;
	wire x_3779;
	wire x_3780;
	wire x_3781;
	wire x_3782;
	wire x_3783;
	wire x_3784;
	wire x_3785;
	wire x_3786;
	wire x_3787;
	wire x_3788;
	wire x_3789;
	wire x_3790;
	wire x_3791;
	wire x_3792;
	wire x_3793;
	wire x_3794;
	wire x_3795;
	wire x_3796;
	wire x_3797;
	wire x_3798;
	wire x_3799;
	wire x_3800;
	wire x_3801;
	wire x_3802;
	wire x_3803;
	wire x_3804;
	wire x_3805;
	wire x_3806;
	wire x_3807;
	wire x_3808;
	wire x_3809;
	wire x_3810;
	wire x_3811;
	wire x_3812;
	wire x_3813;
	wire x_3814;
	wire x_3815;
	wire x_3816;
	wire x_3817;
	wire x_3818;
	wire x_3819;
	wire x_3820;
	wire x_3821;
	wire x_3822;
	wire x_3823;
	wire x_3824;
	wire x_3825;
	wire x_3826;
	wire x_3827;
	wire x_3828;
	wire x_3829;
	wire x_3830;
	wire x_3831;
	wire x_3832;
	wire x_3833;
	wire x_3834;
	wire x_3835;
	wire x_3836;
	wire x_3837;
	wire x_3838;
	wire x_3839;
	wire x_3840;
	wire x_3841;
	wire x_3842;
	wire x_3843;
	wire x_3844;
	wire x_3845;
	wire x_3846;
	wire x_3847;
	wire x_3848;
	wire x_3849;
	wire x_3850;
	wire x_3851;
	wire x_3852;
	wire x_3853;
	wire x_3854;
	wire x_3855;
	wire x_3856;
	wire x_3857;
	wire x_3858;
	wire x_3859;
	wire x_3860;
	wire x_3861;
	wire x_3862;
	wire x_3863;
	wire x_3864;
	wire x_3865;
	wire x_3866;
	wire x_3867;
	wire x_3868;
	wire x_3869;
	wire x_3870;
	wire x_3871;
	wire x_3872;
	wire x_3873;
	wire x_3874;
	wire x_3875;
	wire x_3876;
	wire x_3877;
	wire x_3878;
	wire x_3879;
	wire x_3880;
	wire x_3881;
	wire x_3882;
	wire x_3883;
	wire x_3884;
	wire x_3885;
	wire x_3886;
	wire x_3887;
	wire x_3888;
	wire x_3889;
	wire x_3890;
	wire x_3891;
	wire x_3892;
	wire x_3893;
	wire x_3894;
	wire x_3895;
	wire x_3896;
	wire x_3897;
	wire x_3898;
	wire x_3899;
	wire x_3900;
	wire x_3901;
	wire x_3902;
	wire x_3903;
	wire x_3904;
	wire x_3905;
	wire x_3906;
	wire x_3907;
	wire x_3908;
	wire x_3909;
	wire x_3910;
	wire x_3911;
	wire x_3912;
	wire x_3913;
	wire x_3914;
	wire x_3915;
	wire x_3916;
	wire x_3917;
	wire x_3918;
	wire x_3919;
	wire x_3920;
	wire x_3921;
	wire x_3922;
	wire x_3923;
	wire x_3924;
	wire x_3925;
	wire x_3926;
	wire x_3927;
	wire x_3928;
	wire x_3929;
	wire x_3930;
	wire x_3931;
	wire x_3932;
	wire x_3933;
	wire x_3934;
	wire x_3935;
	wire x_3936;
	wire x_3937;
	wire x_3938;
	wire x_3939;
	wire x_3940;
	wire x_3941;
	wire x_3942;
	wire x_3943;
	wire x_3944;
	wire x_3945;
	wire x_3946;
	wire x_3947;
	wire x_3948;
	wire x_3949;
	wire x_3950;
	wire x_3951;
	wire x_3952;
	wire x_3953;
	wire x_3954;
	wire x_3955;
	wire x_3956;
	wire x_3957;
	wire x_3958;
	wire x_3959;
	wire x_3960;
	wire x_3961;
	wire x_3962;
	wire x_3963;
	wire x_3964;
	wire x_3965;
	wire x_3966;
	wire x_3967;
	wire x_3968;
	wire x_3969;
	wire x_3970;
	wire x_3971;
	wire x_3972;
	wire x_3973;
	wire x_3974;
	wire x_3975;
	wire x_3976;
	wire x_3977;
	wire x_3978;
	wire x_3979;
	wire x_3980;
	wire x_3981;
	wire x_3982;
	wire x_3983;
	wire x_3984;
	wire x_3985;
	wire x_3986;
	wire x_3987;
	wire x_3988;
	wire x_3989;
	wire x_3990;
	wire x_3991;
	wire x_3992;
	wire x_3993;
	wire x_3994;
	wire x_3995;
	wire x_3996;
	wire x_3997;
	wire x_3998;
	wire x_3999;
	wire x_4000;
	wire x_4001;
	wire x_4002;
	wire x_4003;
	wire x_4004;
	wire x_4005;
	wire x_4006;
	wire x_4007;
	wire x_4008;
	wire x_4009;
	wire x_4010;
	wire x_4011;
	wire x_4012;
	wire x_4013;
	wire x_4014;
	wire x_4015;
	wire x_4016;
	wire x_4017;
	wire x_4018;
	wire x_4019;
	wire x_4020;
	wire x_4021;
	wire x_4022;
	wire x_4023;
	wire x_4024;
	wire x_4025;
	wire x_4026;
	wire x_4027;
	wire x_4028;
	wire x_4029;
	wire x_4030;
	wire x_4031;
	wire x_4032;
	wire x_4033;
	wire x_4034;
	wire x_4035;
	wire x_4036;
	wire x_4037;
	wire x_4038;
	wire x_4039;
	wire x_4040;
	wire x_4041;
	wire x_4042;
	wire x_4043;
	wire x_4044;
	wire x_4045;
	wire x_4046;
	wire x_4047;
	wire x_4048;
	wire x_4049;
	wire x_4050;
	wire x_4051;
	wire x_4052;
	wire x_4053;
	wire x_4054;
	wire x_4055;
	wire x_4056;
	wire x_4057;
	wire x_4058;
	wire x_4059;
	wire x_4060;
	wire x_4061;
	wire x_4062;
	wire x_4063;
	wire x_4064;
	wire x_4065;
	wire x_4066;
	wire x_4067;
	wire x_4068;
	wire x_4069;
	wire x_4070;
	wire x_4071;
	wire x_4072;
	wire x_4073;
	wire x_4074;
	wire x_4075;
	wire x_4076;
	wire x_4077;
	wire x_4078;
	wire x_4079;
	wire x_4080;
	wire x_4081;
	wire x_4082;
	wire x_4083;
	wire x_4084;
	wire x_4085;
	wire x_4086;
	wire x_4087;
	wire x_4088;
	wire x_4089;
	wire x_4090;
	wire x_4091;
	wire x_4092;
	wire x_4093;
	wire x_4094;
	wire x_4095;
	wire x_4096;
	wire x_4097;
	wire x_4098;
	wire x_4099;
	wire x_4100;
	wire x_4101;
	wire x_4102;
	wire x_4103;
	wire x_4104;
	wire x_4105;
	wire x_4106;
	wire x_4107;
	wire x_4108;
	wire x_4109;
	wire x_4110;
	wire x_4111;
	wire x_4112;
	wire x_4113;
	wire x_4114;
	wire x_4115;
	wire x_4116;
	wire x_4117;
	wire x_4118;
	wire x_4119;
	wire x_4120;
	wire x_4121;
	wire x_4122;
	wire x_4123;
	wire x_4124;
	wire x_4125;
	wire x_4126;
	wire x_4127;
	wire x_4128;
	wire x_4129;
	wire x_4130;
	wire x_4131;
	wire x_4132;
	wire x_4133;
	wire x_4134;
	wire x_4135;
	wire x_4136;
	wire x_4137;
	wire x_4138;
	wire x_4139;
	wire x_4140;
	wire x_4141;
	wire x_4142;
	wire x_4143;
	wire x_4144;
	wire x_4145;
	wire x_4146;
	wire x_4147;
	wire x_4148;
	wire x_4149;
	wire x_4150;
	wire x_4151;
	wire x_4152;
	wire x_4153;
	wire x_4154;
	wire x_4155;
	wire x_4156;
	wire x_4157;
	wire x_4158;
	wire x_4159;
	wire x_4160;
	wire x_4161;
	wire x_4162;
	wire x_4163;
	wire x_4164;
	wire x_4165;
	wire x_4166;
	wire x_4167;
	wire x_4168;
	wire x_4169;
	wire x_4170;
	wire x_4171;
	wire x_4172;
	wire x_4173;
	wire x_4174;
	wire x_4175;
	wire x_4176;
	wire x_4177;
	wire x_4178;
	wire x_4179;
	wire x_4180;
	wire x_4181;
	wire x_4182;
	wire x_4183;
	wire x_4184;
	wire x_4185;
	wire x_4186;
	wire x_4187;
	wire x_4188;
	wire x_4189;
	wire x_4190;
	wire x_4191;
	wire x_4192;
	wire x_4193;
	wire x_4194;
	wire x_4195;
	wire x_4196;
	wire x_4197;
	wire x_4198;
	wire x_4199;
	wire x_4200;
	wire x_4201;
	wire x_4202;
	wire x_4203;
	wire x_4204;
	wire x_4205;
	wire x_4206;
	wire x_4207;
	wire x_4208;
	wire x_4209;
	wire x_4210;
	wire x_4211;
	wire x_4212;
	wire x_4213;
	wire x_4214;
	wire x_4215;
	wire x_4216;
	wire x_4217;
	wire x_4218;
	wire x_4219;
	wire x_4220;
	wire x_4221;
	wire x_4222;
	wire x_4223;
	wire x_4224;
	wire x_4225;
	wire x_4226;
	wire x_4227;
	wire x_4228;
	wire x_4229;
	wire x_4230;
	wire x_4231;
	wire x_4232;
	wire x_4233;
	wire x_4234;
	wire x_4235;
	wire x_4236;
	wire x_4237;
	wire x_4238;
	wire x_4239;
	wire x_4240;
	wire x_4241;
	wire x_4242;
	wire x_4243;
	wire x_4244;
	wire x_4245;
	wire x_4246;
	wire x_4247;
	wire x_4248;
	wire x_4249;
	wire x_4250;
	wire x_4251;
	wire x_4252;
	wire x_4253;
	wire x_4254;
	wire x_4255;
	wire x_4256;
	wire x_4257;
	wire x_4258;
	wire x_4259;
	wire x_4260;
	wire x_4261;
	wire x_4262;
	wire x_4263;
	wire x_4264;
	wire x_4265;
	wire x_4266;
	wire x_4267;
	wire x_4268;
	wire x_4269;
	wire x_4270;
	wire x_4271;
	wire x_4272;
	wire x_4273;
	wire x_4274;
	wire x_4275;
	wire x_4276;
	wire x_4277;
	wire x_4278;
	wire x_4279;
	wire x_4280;
	wire x_4281;
	wire x_4282;
	wire x_4283;
	wire x_4284;
	wire x_4285;
	wire x_4286;
	wire x_4287;
	wire x_4288;
	wire x_4289;
	wire x_4290;
	wire x_4291;
	wire x_4292;
	wire x_4293;
	wire x_4294;
	wire x_4295;
	wire x_4296;
	wire x_4297;
	wire x_4298;
	wire x_4299;
	wire x_4300;
	wire x_4301;
	wire x_4302;
	wire x_4303;
	wire x_4304;
	wire x_4305;
	wire x_4306;
	wire x_4307;
	wire x_4308;
	wire x_4309;
	wire x_4310;
	wire x_4311;
	wire x_4312;
	wire x_4313;
	wire x_4314;
	wire x_4315;
	wire x_4316;
	wire x_4317;
	wire x_4318;
	wire x_4319;
	wire x_4320;
	wire x_4321;
	wire x_4322;
	wire x_4323;
	wire x_4324;
	wire x_4325;
	wire x_4326;
	wire x_4327;
	wire x_4328;
	wire x_4329;
	wire x_4330;
	wire x_4331;
	wire x_4332;
	wire x_4333;
	wire x_4334;
	wire x_4335;
	wire x_4336;
	wire x_4337;
	wire x_4338;
	wire x_4339;
	wire x_4340;
	wire x_4341;
	wire x_4342;
	wire x_4343;
	wire x_4344;
	wire x_4345;
	wire x_4346;
	wire x_4347;
	wire x_4348;
	wire x_4349;
	wire x_4350;
	wire x_4351;
	wire x_4352;
	wire x_4353;
	wire x_4354;
	wire x_4355;
	wire x_4356;
	wire x_4357;
	wire x_4358;
	wire x_4359;
	wire x_4360;
	wire x_4361;
	wire x_4362;
	wire x_4363;
	wire x_4364;
	wire x_4365;
	wire x_4366;
	wire x_4367;
	wire x_4368;
	wire x_4369;
	wire x_4370;
	wire x_4371;
	wire x_4372;
	wire x_4373;
	wire x_4374;
	wire x_4375;
	wire x_4376;
	wire x_4377;
	wire x_4378;
	wire x_4379;
	wire x_4380;
	wire x_4381;
	wire x_4382;
	wire x_4383;
	wire x_4384;
	wire x_4385;
	wire x_4386;
	wire x_4387;
	wire x_4388;
	wire x_4389;
	wire x_4390;
	wire x_4391;
	wire x_4392;
	wire x_4393;
	wire x_4394;
	wire x_4395;
	wire x_4396;
	wire x_4397;
	wire x_4398;
	wire x_4399;
	wire x_4400;
	wire x_4401;
	wire x_4402;
	wire x_4403;
	wire x_4404;
	wire x_4405;
	wire x_4406;
	wire x_4407;
	wire x_4408;
	wire x_4409;
	wire x_4410;
	wire x_4411;
	wire x_4412;
	wire x_4413;
	wire x_4414;
	wire x_4415;
	wire x_4416;
	wire x_4417;
	wire x_4418;
	wire x_4419;
	wire x_4420;
	wire x_4421;
	wire x_4422;
	wire x_4423;
	wire x_4424;
	wire x_4425;
	wire x_4426;
	wire x_4427;
	wire x_4428;
	wire x_4429;
	wire x_4430;
	wire x_4431;
	wire x_4432;
	wire x_4433;
	wire x_4434;
	wire x_4435;
	wire x_4436;
	wire x_4437;
	wire x_4438;
	wire x_4439;
	wire x_4440;
	wire x_4441;
	wire x_4442;
	wire x_4443;
	wire x_4444;
	wire x_4445;
	wire x_4446;
	wire x_4447;
	wire x_4448;
	wire x_4449;
	wire x_4450;
	wire x_4451;
	wire x_4452;
	wire x_4453;
	wire x_4454;
	wire x_4455;
	wire x_4456;
	wire x_4457;
	wire x_4458;
	wire x_4459;
	wire x_4460;
	wire x_4461;
	wire x_4462;
	wire x_4463;
	wire x_4464;
	wire x_4465;
	wire x_4466;
	wire x_4467;
	wire x_4468;
	wire x_4469;
	wire x_4470;
	wire x_4471;
	wire x_4472;
	wire x_4473;
	wire x_4474;
	wire x_4475;
	wire x_4476;
	wire x_4477;
	wire x_4478;
	wire x_4479;
	wire x_4480;
	wire x_4481;
	wire x_4482;
	wire x_4483;
	wire x_4484;
	wire x_4485;
	wire x_4486;
	wire x_4487;
	wire x_4488;
	wire x_4489;
	wire x_4490;
	wire x_4491;
	wire x_4492;
	wire x_4493;
	wire x_4494;
	wire x_4495;
	wire x_4496;
	wire x_4497;
	wire x_4498;
	wire x_4499;
	wire x_4500;
	wire x_4501;
	wire x_4502;
	wire x_4503;
	wire x_4504;
	wire x_4505;
	wire x_4506;
	wire x_4507;
	wire x_4508;
	wire x_4509;
	wire x_4510;
	wire x_4511;
	wire x_4512;
	wire x_4513;
	wire x_4514;
	wire x_4515;
	wire x_4516;
	wire x_4517;
	wire x_4518;
	wire x_4519;
	wire x_4520;
	wire x_4521;
	wire x_4522;
	wire x_4523;
	wire x_4524;
	wire x_4525;
	wire x_4526;
	wire x_4527;
	wire x_4528;
	wire x_4529;
	wire x_4530;
	wire x_4531;
	wire x_4532;
	wire x_4533;
	wire x_4534;
	wire x_4535;
	wire x_4536;
	wire x_4537;
	wire x_4538;
	wire x_4539;
	wire x_4540;
	wire x_4541;
	wire x_4542;
	wire x_4543;
	wire x_4544;
	wire x_4545;
	wire x_4546;
	wire x_4547;
	wire x_4548;
	wire x_4549;
	wire x_4550;
	wire x_4551;
	wire x_4552;
	wire x_4553;
	wire x_4554;
	wire x_4555;
	wire x_4556;
	wire x_4557;
	wire x_4558;
	wire x_4559;
	wire x_4560;
	wire x_4561;
	wire x_4562;
	wire x_4563;
	wire x_4564;
	wire x_4565;
	wire x_4566;
	wire x_4567;
	wire x_4568;
	wire x_4569;
	wire x_4570;
	wire x_4571;
	wire x_4572;
	wire x_4573;
	wire x_4574;
	wire x_4575;
	wire x_4576;
	wire x_4577;
	wire x_4578;
	wire x_4579;
	wire x_4580;
	wire x_4581;
	wire x_4582;
	wire x_4583;
	wire x_4584;
	wire x_4585;
	wire x_4586;
	wire x_4587;
	wire x_4588;
	wire x_4589;
	wire x_4590;
	wire x_4591;
	wire x_4592;
	wire x_4593;
	wire x_4594;
	wire x_4595;
	wire x_4596;
	wire x_4597;
	wire x_4598;
	wire x_4599;
	wire x_4600;
	wire x_4601;
	wire x_4602;
	wire x_4603;
	wire x_4604;
	wire x_4605;
	wire x_4606;
	wire x_4607;
	wire x_4608;
	wire x_4609;
	wire x_4610;
	wire x_4611;
	wire x_4612;
	wire x_4613;
	wire x_4614;
	wire x_4615;
	wire x_4616;
	wire x_4617;
	wire x_4618;
	wire x_4619;
	wire x_4620;
	wire x_4621;
	wire x_4622;
	wire x_4623;
	wire x_4624;
	wire x_4625;
	wire x_4626;
	wire x_4627;
	wire x_4628;
	wire x_4629;
	wire x_4630;
	wire x_4631;
	wire x_4632;
	wire x_4633;
	wire x_4634;
	wire x_4635;
	wire x_4636;
	wire x_4637;
	wire x_4638;
	wire x_4639;
	wire x_4640;
	wire x_4641;
	wire x_4642;
	wire x_4643;
	wire x_4644;
	wire x_4645;
	wire x_4646;
	wire x_4647;
	wire x_4648;
	wire x_4649;
	wire x_4650;
	wire x_4651;
	wire x_4652;
	wire x_4653;
	wire x_4654;
	wire x_4655;
	wire x_4656;
	wire x_4657;
	wire x_4658;
	wire x_4659;
	wire x_4660;
	wire x_4661;
	wire x_4662;
	wire x_4663;
	wire x_4664;
	wire x_4665;
	wire x_4666;
	wire x_4667;
	wire x_4668;
	wire x_4669;
	wire x_4670;
	wire x_4671;
	wire x_4672;
	wire x_4673;
	wire x_4674;
	wire x_4675;
	wire x_4676;
	wire x_4677;
	wire x_4678;
	wire x_4679;
	wire x_4680;
	wire x_4681;
	wire x_4682;
	wire x_4683;
	wire x_4684;
	wire x_4685;
	wire x_4686;
	wire x_4687;
	wire x_4688;
	wire x_4689;
	wire x_4690;
	wire x_4691;
	wire x_4692;
	wire x_4693;
	wire x_4694;
	wire x_4695;
	wire x_4696;
	wire x_4697;
	wire x_4698;
	wire x_4699;
	wire x_4700;
	wire x_4701;
	wire x_4702;
	wire x_4703;
	wire x_4704;
	wire x_4705;
	wire x_4706;
	wire x_4707;
	wire x_4708;
	wire x_4709;
	wire x_4710;
	wire x_4711;
	wire x_4712;
	wire x_4713;
	wire x_4714;
	wire x_4715;
	wire x_4716;
	wire x_4717;
	wire x_4718;
	wire x_4719;
	wire x_4720;
	wire x_4721;
	wire x_4722;
	wire x_4723;
	wire x_4724;
	wire x_4725;
	wire x_4726;
	wire x_4727;
	wire x_4728;
	wire x_4729;
	wire x_4730;
	wire x_4731;
	wire x_4732;
	wire x_4733;
	wire x_4734;
	wire x_4735;
	wire x_4736;
	wire x_4737;
	wire x_4738;
	wire x_4739;
	wire x_4740;
	wire x_4741;
	wire x_4742;
	wire x_4743;
	wire x_4744;
	wire x_4745;
	wire x_4746;
	wire x_4747;
	wire x_4748;
	wire x_4749;
	wire x_4750;
	wire x_4751;
	wire x_4752;
	wire x_4753;
	wire x_4754;
	wire x_4755;
	wire x_4756;
	wire x_4757;
	wire x_4758;
	wire x_4759;
	wire x_4760;
	wire x_4761;
	wire x_4762;
	wire x_4763;
	wire x_4764;
	wire x_4765;
	wire x_4766;
	wire x_4767;
	wire x_4768;
	wire x_4769;
	wire x_4770;
	wire x_4771;
	wire x_4772;
	wire x_4773;
	wire x_4774;
	wire x_4775;
	wire x_4776;
	wire x_4777;
	wire x_4778;
	wire x_4779;
	wire x_4780;
	wire x_4781;
	wire x_4782;
	wire x_4783;
	wire x_4784;
	wire x_4785;
	wire x_4786;
	wire x_4787;
	wire x_4788;
	wire x_4789;
	wire x_4790;
	wire x_4791;
	wire x_4792;
	wire x_4793;
	wire x_4794;
	wire x_4795;
	wire x_4796;
	wire x_4797;
	wire x_4798;
	wire x_4799;
	wire x_4800;
	wire x_4801;
	wire x_4802;
	wire x_4803;
	wire x_4804;
	wire x_4805;
	wire x_4806;
	wire x_4807;
	wire x_4808;
	wire x_4809;
	wire x_4810;
	wire x_4811;
	wire x_4812;
	wire x_4813;
	wire x_4814;
	wire x_4815;
	wire x_4816;
	wire x_4817;
	wire x_4818;
	wire x_4819;
	wire x_4820;
	wire x_4821;
	wire x_4822;
	wire x_4823;
	wire x_4824;
	wire x_4825;
	wire x_4826;
	wire x_4827;
	wire x_4828;
	wire x_4829;
	wire x_4830;
	wire x_4831;
	wire x_4832;
	wire x_4833;
	wire x_4834;
	wire x_4835;
	output o_1;
	assign x_2418 = (v_91 | ~v_21) ;
	assign x_2417 = (v_91 | ~v_22) ;
	assign x_2413 = (v_92 | ~v_14) ;
	assign x_2412 = (v_92 | ~v_15) ;
	assign x_2408 = (v_94 | v_23) ;
	assign x_2407 = (v_94 | v_29) ;
	assign x_2399 = (v_98 | v_41) ;
	assign x_2398 = (v_99 | v_19) ;
	assign x_2394 = (((((((((((((((v_35 | v_36) | v_79) | v_71) | v_70) | v_82) | v_88) | ~v_100) | ~v_99) | ~v_98) | ~v_97) | ~v_96) | ~v_95) | ~v_94) | ~v_93) | v_101) ;
	assign x_2393 = (v_102 | ~v_23) ;
	assign x_2389 = (v_104 | v_23) ;
	assign x_2388 = (v_104 | v_28) ;
	assign x_2380 = (v_108 | v_54) ;
	assign x_2379 = (v_109 | v_19) ;
	assign x_2375 = (v_111 | v_27) ;
	assign x_2374 = (v_112 | ~v_20) ;
	assign x_2370 = (v_114 | v_20) ;
	assign x_2369 = (v_114 | v_68) ;
	assign x_2361 = (v_118 | v_69) ;
	assign x_2360 = (((((((((((((((v_61 | v_76) | v_81) | v_62) | v_77) | v_84) | ~v_118) | ~v_117) | v_90) | ~v_116) | ~v_115) | ~v_114) | ~v_113) | ~v_112) | ~v_111) | v_119) ;
	assign x_2356 = (v_121 | ~v_19) ;
	assign x_2355 = (v_121 | v_38) ;
	assign x_2351 = (v_123 | v_29) ;
	assign x_2350 = (v_124 | ~v_9) ;
	assign x_2342 = (v_128 | v_11) ;
	assign x_2341 = (v_128 | v_42) ;
	assign x_2337 = (v_131 | v_19) ;
	assign x_2336 = (v_131 | v_54) ;
	assign x_2332 = (v_133 | v_52) ;
	assign x_2331 = (v_134 | ~v_9) ;
	assign x_2323 = (((((((((((((((v_50 | v_49) | v_48) | v_46) | v_47) | v_73) | v_80) | ~v_137) | ~v_136) | ~v_135) | ~v_134) | ~v_133) | ~v_132) | ~v_131) | ~v_130) | v_138) ;
	assign x_2322 = (v_139 | v_19) ;
	assign x_2318 = (v_141 | ~v_9) ;
	assign x_2317 = (v_141 | v_66) ;
	assign x_2313 = (v_143 | v_64) ;
	assign x_2312 = (v_144 | ~v_17) ;
	assign x_2304 = (v_148 | ~v_138) ;
	assign x_2303 = (v_148 | ~v_129) ;
	assign x_2299 = (v_150 | v_26) ;
	assign x_2298 = (v_151 | ~v_28) ;
	assign x_2294 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_148) | ~v_120) | v_153) ;
	assign x_2293 = (v_154 | ~v_22) ;
	assign x_2285 = (v_158 | v_14) ;
	assign x_2284 = (v_158 | v_56) ;
	assign x_2280 = (v_161 | ~v_22) ;
	assign x_2279 = (v_161 | v_27) ;
	assign x_2275 = (v_163 | v_68) ;
	assign x_2274 = (v_164 | v_14) ;
	assign x_2266 = (v_168 | v_29) ;
	assign x_2265 = (v_169 | ~v_14) ;
	assign x_2261 = (v_171 | ~v_16) ;
	assign x_2260 = (v_171 | v_39) ;
	assign x_2256 = (v_173 | v_43) ;
	assign x_2255 = (((((((((((((((v_35 | v_37) | v_36) | v_79) | v_71) | v_70) | v_88) | ~v_173) | ~v_172) | ~v_171) | ~v_170) | ~v_169) | ~v_98) | ~v_97) | ~v_168) | v_174) ;
	assign x_2247 = (v_178 | ~v_10) ;
	assign x_2246 = (v_178 | v_39) ;
	assign x_2242 = (v_180 | v_29) ;
	assign x_2241 = (v_181 | v_10) ;
	assign x_2237 = (v_183 | v_51) ;
	assign x_2236 = (v_184 | ~v_13) ;
	assign x_2228 = (v_188 | v_10) ;
	assign x_2227 = (v_188 | v_55) ;
	assign x_2223 = (v_191 | ~v_13) ;
	assign x_2222 = (v_191 | v_27) ;
	assign x_2218 = (v_193 | v_30) ;
	assign x_2217 = (v_194 | v_14) ;
	assign x_2209 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_197) | ~v_175) | v_198) ;
	assign x_2208 = (v_199 | ~v_21) ;
	assign x_2204 = (v_201 | v_12) ;
	assign x_2203 = (v_201 | v_42) ;
	assign x_2199 = (v_204 | ~v_21) ;
	assign x_2198 = (v_204 | v_26) ;
	assign x_2190 = (v_209 | ~v_21) ;
	assign x_2189 = (v_209 | v_27) ;
	assign x_2185 = (v_211 | v_65) ;
	assign x_2184 = (v_212 | v_12) ;
	assign x_2180 = (v_214 | ~v_208) ;
	assign x_2179 = (v_214 | ~v_203) ;
	assign x_2171 = (v_218 | v_52) ;
	assign x_2170 = (v_219 | ~v_24) ;
	assign x_2166 = (v_221 | v_16) ;
	assign x_2165 = (v_221 | v_28) ;
	assign x_2161 = (v_224 | ~v_22) ;
	assign x_2160 = (v_224 | v_65) ;
	assign x_2152 = (v_228 | v_27) ;
	assign x_2151 = (v_229 | v_22) ;
	assign x_2147 = (v_231 | v_25) ;
	assign x_2146 = (v_232 | ~v_22) ;
	assign x_2142 = (v_234 | ~v_24) ;
	assign x_2141 = (v_234 | v_40) ;
	assign x_2133 = (v_238 | ~v_223) ;
	assign x_2132 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_238) | ~v_216) | v_239) ;
	assign x_2124 = (v_243 | v_25) ;
	assign x_2123 = (((((((((((((((v_37 | v_34) | v_79) | v_72) | v_71) | v_70) | v_85) | ~v_243) | ~v_127) | ~v_236) | ~v_234) | ~v_121) | ~v_242) | ~v_241) | ~v_240) | v_244) ;
	assign x_2115 = (v_248 | v_28) ;
	assign x_2114 = (((((((((((((((~v_248 | v_50) | v_75) | v_74) | v_47) | v_73) | v_86) | v_80) | ~v_222) | ~v_247) | ~v_219) | ~v_131) | ~v_130) | ~v_246) | ~v_245) | v_249) ;
	assign x_2110 = (v_251 | v_65) ;
	assign x_2109 = (v_252 | v_23) ;
	assign x_2105 = (((((((((((((((~v_253 | v_76) | v_81) | v_63) | v_60) | v_78) | v_77) | ~v_252) | v_87) | ~v_143) | ~v_227) | ~v_226) | ~v_139) | ~v_251) | ~v_250) | v_254) ;
	assign x_2104 = (v_255 | ~v_254) ;
	assign x_2096 = (v_259 | v_18) ;
	assign x_2095 = (v_259 | v_29) ;
	assign x_2091 = (v_262 | ~v_18) ;
	assign x_2090 = (v_262 | v_26) ;
	assign x_2086 = (v_264 | v_55) ;
	assign x_2085 = (v_265 | v_18) ;
	assign x_2077 = (v_269 | v_30) ;
	assign x_2076 = (v_270 | v_15) ;
	assign x_2072 = (v_272 | ~v_266) ;
	assign x_2071 = (v_272 | ~v_261) ;
	assign x_2067 = (v_275 | ~v_273) ;
	assign x_2066 = (v_275 | ~v_256) ;
	assign x_2058 = (v_279 | v_25) ;
	assign x_2057 = (((((((((((((((v_35 | v_37) | v_34) | v_79) | v_72) | v_71) | v_70) | ~v_279) | ~v_99) | ~v_179) | ~v_176) | ~v_96) | ~v_278) | ~v_277) | ~v_276) | v_280) ;
	assign x_2053 = (v_282 | v_52) ;
	assign x_2052 = (v_283 | v_18) ;
	assign x_2048 = (((((((((((((((~v_284 | v_50) | v_48) | v_75) | v_74) | v_47) | v_73) | v_80) | ~v_109) | ~v_186) | ~v_183) | ~v_106) | ~v_283) | ~v_282) | ~v_281) | v_285) ;
	assign x_2047 = (v_286 | ~v_15) ;
	assign x_2039 = (((((((((((((((~v_289 | v_61) | v_76) | v_81) | v_63) | v_60) | v_78) | v_77) | ~v_118) | ~v_116) | ~v_194) | ~v_190) | ~v_288) | ~v_287) | ~v_286) | v_290) ;
	assign x_2038 = (v_291 | ~v_290) ;
	assign x_2034 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_214) | ~v_238) | v_293) ;
	assign x_2033 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_291) | ~v_148) | v_294) ;
	assign x_2029 = (v_296 | ~v_293) ;
	assign x_2028 = (v_296 | ~v_292) ;
	assign x_2020 = (v_300 | ~v_9) ;
	assign x_2019 = (v_300 | v_38) ;
	assign x_2015 = (v_302 | v_41) ;
	assign x_2014 = (((((((((((((((v_32 | v_37) | v_36) | v_34) | v_71) | v_70) | v_85) | ~v_302) | ~v_301) | ~v_236) | ~v_300) | ~v_299) | ~v_298) | ~v_297) | ~v_234) | v_303) ;
	assign x_2010 = (v_305 | v_51) ;
	assign x_2009 = (v_306 | v_21) ;
	assign x_2001 = (((((((((((((((v_50 | v_49) | v_45) | v_74) | v_47) | v_73) | v_86) | ~v_309) | ~v_222) | ~v_308) | ~v_307) | ~v_306) | ~v_305) | ~v_304) | ~v_219) | v_310) ;
	assign x_2000 = (v_311 | ~v_12) ;
	assign x_1996 = (v_313 | ~v_9) ;
	assign x_1995 = (v_313 | v_64) ;
	assign x_1991 = (v_315 | v_67) ;
	assign x_1990 = (v_316 | v_12) ;
	assign x_1982 = (v_320 | v_25) ;
	assign x_1981 = (v_321 | ~v_13) ;
	assign x_1973 = (v_325 | v_52) ;
	assign x_1972 = (v_326 | v_10) ;
	assign x_1964 = (v_330 | v_27) ;
	assign x_1963 = (v_331 | ~v_13) ;
	assign x_1959 = (v_333 | v_13) ;
	assign x_1958 = (v_333 | v_68) ;
	assign x_1954 = (v_335 | ~v_324) ;
	assign x_1953 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_291) | ~v_335) | v_336) ;
	assign x_1945 = (v_341 | v_11) ;
	assign x_1944 = (v_341 | v_29) ;
	assign x_1940 = (v_344 | v_17) ;
	assign x_1939 = (v_344 | v_55) ;
	assign x_1935 = (v_346 | v_26) ;
	assign x_1934 = (((((((((((((((v_50 | v_49) | v_48) | v_45) | v_74) | v_47) | v_73) | ~v_309) | ~v_109) | ~v_346) | ~v_345) | ~v_305) | ~v_344) | ~v_343) | ~v_106) | v_347) ;
	assign x_1926 = (v_351 | v_30) ;
	assign x_1925 = (((((((((((((((v_61 | v_76) | v_63) | v_62) | v_60) | v_58) | v_77) | ~v_351) | ~v_350) | ~v_118) | ~v_315) | ~v_116) | ~v_313) | ~v_349) | ~v_348) | v_352) ;
	assign x_1921 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_214) | ~v_353) | v_354) ;
	assign x_1920 = (((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_120) | v_355) ;
	assign x_1916 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_318) | ~v_356) | v_357) ;
	assign x_1915 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_238) | ~v_120) | v_358) ;
	assign x_1907 = (v_364 | ~v_363) ;
	assign x_1906 = (v_364 | ~v_362) ;
	assign x_1902 = ((~v_364 | ~v_296) | v_365) ;
	assign x_1901 = (v_366 | ~v_363) ;
	assign x_1897 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_175) | ~v_361) | v_368) ;
	assign x_1896 = (v_369 | ~v_355) ;
	assign x_1888 = (v_373 | ~v_372) ;
	assign x_1887 = (v_373 | ~v_371) ;
	assign x_1883 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_148) | ~v_318) | v_376) ;
	assign x_1882 = (((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_255) | v_377) ;
	assign x_1878 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_291) | ~v_378) | v_379) ;
	assign x_1877 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_291) | ~v_255) | v_380) ;
	assign x_1869 = ((~v_383 | ~v_369) | v_384) ;
	assign x_1868 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_197) | ~v_366) | v_385) ;
	assign x_1864 = (v_387 | ~v_358) ;
	assign x_1863 = (v_387 | ~v_386) ;
	assign x_1859 = (v_388 | ~v_17) ;
	assign x_1858 = (v_388 | ~v_18) ;
	assign x_1850 = ((((v_24 | v_23) | v_22) | v_21) | v_391) ;
	assign x_1849 = ((((v_13 | v_16) | v_15) | v_14) | v_392) ;
	assign x_1845 = (v_395 | ~v_393) ;
	assign x_1844 = (v_395 | ~v_392) ;
	assign x_1840 = ((~v_20 | ~v_42) | v_398) ;
	assign x_1839 = ((v_19 | ~v_40) | v_399) ;
	assign x_1831 = (v_404 | ~v_71) ;
	assign x_1830 = (v_404 | ~v_79) ;
	assign x_1822 = (v_404 | ~v_398) ;
	assign x_1821 = (v_404 | ~v_397) ;
	assign x_1813 = ((~v_24 | ~v_54) | v_411) ;
	assign x_1812 = ((~v_19 | ~v_56) | v_412) ;
	assign x_1808 = (v_413 | ~v_74) ;
	assign x_1807 = (v_413 | ~v_80) ;
	assign x_1803 = (v_413 | ~v_411) ;
	assign x_1802 = (v_413 | ~v_410) ;
	assign x_1794 = ((~v_23 | ~v_30) | v_416) ;
	assign x_1793 = ((~v_20 | ~v_68) | v_417) ;
	assign x_1789 = ((~v_19 | ~v_69) | v_421) ;
	assign x_1788 = (v_422 | ~v_61) ;
	assign x_1784 = (v_422 | ~v_81) ;
	assign x_1783 = (v_422 | ~v_84) ;
	assign x_1775 = (v_422 | ~v_415) ;
	assign x_1774 = (v_422 | ~v_414) ;
	assign x_1770 = ((~v_17 | ~v_29) | v_426) ;
	assign x_1769 = ((v_9 | ~v_40) | v_427) ;
	assign x_1765 = ((~v_11 | ~v_42) | v_431) ;
	assign x_1764 = (v_432 | ~v_33) ;
	assign x_1756 = (v_432 | ~v_430) ;
	assign x_1755 = (v_432 | ~v_429) ;
	assign x_1751 = (v_432 | ~v_425) ;
	assign x_1750 = (v_432 | ~v_424) ;
	assign x_1746 = ((v_11 | ~v_52) | v_436) ;
	assign x_1745 = ((v_9 | ~v_53) | v_437) ;
	assign x_1737 = (v_441 | ~v_50) ;
	assign x_1736 = (v_441 | ~v_73) ;
	assign x_1732 = (v_441 | ~v_438) ;
	assign x_1731 = (v_441 | ~v_437) ;
	assign x_1727 = (v_441 | ~v_433) ;
	assign x_1726 = ((~v_19 | ~v_67) | v_442) ;
	assign x_1718 = (v_450 | ~v_59) ;
	assign x_1717 = (v_450 | ~v_60) ;
	assign x_1713 = (v_450 | ~v_76) ;
	assign x_1712 = (v_450 | ~v_81) ;
	assign x_1708 = (v_450 | ~v_446) ;
	assign x_1707 = (v_450 | ~v_445) ;
	assign x_1699 = ((~v_27 | v_26) | v_455) ;
	assign x_1698 = (v_456 | ~v_455) ;
	assign x_1694 = (v_456 | ~v_451) ;
	assign x_1693 = (v_456 | ~v_423) ;
	assign x_1689 = ((v_14 | ~v_53) | v_460) ;
	assign x_1688 = ((~v_14 | ~v_56) | v_461) ;
	assign x_1680 = (v_463 | ~v_89) ;
	assign x_1679 = (v_463 | ~v_462) ;
	assign x_1671 = ((~v_27 | v_22) | v_464) ;
	assign x_1670 = ((v_16 | ~v_65) | v_465) ;
	assign x_1662 = (v_470 | ~v_76) ;
	assign x_1661 = (v_470 | ~v_77) ;
	assign x_1657 = (v_470 | ~v_90) ;
	assign x_1656 = (v_470 | ~v_468) ;
	assign x_1652 = (v_470 | ~v_465) ;
	assign x_1651 = (v_470 | ~v_464) ;
	assign x_1643 = (v_477 | ~v_36) ;
	assign x_1642 = (v_477 | ~v_37) ;
	assign x_1638 = (v_477 | ~v_88) ;
	assign x_1637 = (v_477 | ~v_476) ;
	assign x_1633 = (v_477 | ~v_472) ;
	assign x_1632 = (v_477 | ~v_401) ;
	assign x_1624 = ((~v_13 | ~v_29) | v_483) ;
	assign x_1623 = ((~v_10 | ~v_42) | v_484) ;
	assign x_1619 = (v_485 | ~v_36) ;
	assign x_1618 = (v_485 | ~v_70) ;
	assign x_1614 = (v_485 | ~v_483) ;
	assign x_1613 = (v_485 | ~v_482) ;
	assign x_1605 = ((v_10 | ~v_52) | v_488) ;
	assign x_1604 = ((~v_14 | ~v_54) | v_489) ;
	assign x_1600 = (v_492 | ~v_47) ;
	assign x_1599 = (v_492 | ~v_48) ;
	assign x_1595 = (v_492 | ~v_83) ;
	assign x_1594 = (v_492 | ~v_440) ;
	assign x_1586 = ((v_14 | ~v_64) | v_493) ;
	assign x_1585 = ((~v_27 | v_13) | v_494) ;
	assign x_1581 = ((~v_10 | ~v_68) | v_498) ;
	assign x_1580 = (v_499 | ~v_59) ;
	assign x_1576 = (v_499 | ~v_76) ;
	assign x_1575 = (v_499 | ~v_81) ;
	assign x_1567 = (v_499 | ~v_445) ;
	assign x_1566 = (v_499 | ~v_444) ;
	assign x_1562 = (v_501 | ~v_453) ;
	assign x_1561 = (v_501 | ~v_452) ;
	assign x_1557 = ((~v_21 | ~v_29) | v_503) ;
	assign x_1556 = ((~v_12 | ~v_42) | v_504) ;
	assign x_1548 = (v_506 | ~v_88) ;
	assign x_1547 = (v_506 | ~v_505) ;
	assign x_1543 = (v_506 | ~v_503) ;
	assign x_1542 = (v_506 | ~v_502) ;
	assign x_1538 = ((v_12 | ~v_52) | v_508) ;
	assign x_1537 = ((~v_21 | ~v_28) | v_509) ;
	assign x_1529 = (v_511 | ~v_440) ;
	assign x_1528 = (v_511 | ~v_89) ;
	assign x_1520 = ((~v_27 | v_21) | v_512) ;
	assign x_1519 = ((~v_21 | ~v_30) | v_513) ;
	assign x_1511 = (v_516 | ~v_81) ;
	assign x_1510 = (v_516 | ~v_515) ;
	assign x_1506 = (v_516 | ~v_445) ;
	assign x_1505 = (v_516 | ~v_444) ;
	assign x_1501 = (((~v_516 | ~v_511) | ~v_506) | v_517) ;
	assign x_1500 = (v_518 | ~v_455) ;
	assign x_1492 = ((v_24 | ~v_53) | v_522) ;
	assign x_1491 = ((~v_22 | ~v_55) | v_523) ;
	assign x_1487 = (v_526 | ~v_49) ;
	assign x_1486 = (v_526 | ~v_50) ;
	assign x_1482 = (v_526 | ~v_86) ;
	assign x_1481 = (v_526 | ~v_525) ;
	assign x_1473 = ((v_22 | ~v_65) | v_527) ;
	assign x_1472 = ((~v_16 | ~v_30) | v_528) ;
	assign x_1468 = ((~v_22 | ~v_68) | v_532) ;
	assign x_1467 = (v_533 | ~v_60) ;
	assign x_1463 = (v_533 | ~v_77) ;
	assign x_1462 = (v_533 | ~v_81) ;
	assign x_1454 = (v_533 | ~v_528) ;
	assign x_1453 = (v_533 | ~v_527) ;
	assign x_1449 = ((v_24 | ~v_40) | v_537) ;
	assign x_1448 = ((~v_22 | ~v_42) | v_538) ;
	assign x_1444 = (v_540 | ~v_37) ;
	assign x_1443 = (v_540 | ~v_70) ;
	assign x_1435 = (v_540 | ~v_537) ;
	assign x_1434 = (v_540 | ~v_536) ;
	assign x_1430 = (v_542 | ~v_455) ;
	assign x_1429 = (v_542 | ~v_454) ;
	assign x_1425 = (v_542 | ~v_519) ;
	assign x_1424 = ((~v_39 | v_23) | v_543) ;
	assign x_1416 = (v_547 | ~v_72) ;
	assign x_1415 = (v_547 | ~v_79) ;
	assign x_1411 = (v_547 | ~v_539) ;
	assign x_1410 = (v_547 | ~v_537) ;
	assign x_1406 = (v_547 | ~v_543) ;
	assign x_1405 = ((~v_26 | v_20) | v_548) ;
	assign x_1397 = (v_552 | ~v_74) ;
	assign x_1396 = (v_552 | ~v_75) ;
	assign x_1392 = (v_552 | ~v_550) ;
	assign x_1391 = (v_552 | ~v_522) ;
	assign x_1387 = (v_552 | ~v_548) ;
	assign x_1386 = ((~v_27 | v_20) | v_553) ;
	assign x_1378 = (v_557 | ~v_77) ;
	assign x_1377 = (v_557 | ~v_78) ;
	assign x_1369 = (v_557 | ~v_554) ;
	assign x_1368 = (v_557 | ~v_553) ;
	assign x_1360 = ((~v_39 | v_15) | v_560) ;
	assign x_1359 = ((~v_15 | ~v_42) | v_561) ;
	assign x_1355 = (v_564 | ~v_35) ;
	assign x_1354 = (v_564 | ~v_36) ;
	assign x_1350 = (v_564 | ~v_82) ;
	assign x_1349 = (v_564 | ~v_563) ;
	assign x_1341 = ((~v_26 | v_18) | v_565) ;
	assign x_1340 = ((v_15 | ~v_52) | v_566) ;
	assign x_1336 = (v_569 | ~v_48) ;
	assign x_1335 = (v_569 | ~v_49) ;
	assign x_1331 = (v_569 | ~v_83) ;
	assign x_1330 = (v_569 | ~v_568) ;
	assign x_1322 = ((~v_27 | v_18) | v_570) ;
	assign x_1321 = ((v_15 | ~v_65) | v_571) ;
	assign x_1317 = (v_574 | ~v_61) ;
	assign x_1316 = (v_574 | ~v_62) ;
	assign x_1312 = (v_574 | ~v_84) ;
	assign x_1311 = (v_574 | ~v_446) ;
	assign x_1303 = (((~v_574 | ~v_569) | ~v_564) | v_575) ;
	assign x_1302 = (v_576 | ~v_455) ;
	assign x_1298 = (v_576 | ~v_500) ;
	assign x_1297 = (v_576 | ~v_575) ;
	assign x_1293 = (v_577 | ~v_452) ;
	assign x_1292 = (v_577 | ~v_451) ;
	assign x_1284 = (v_583 | ~v_37) ;
	assign x_1283 = (v_583 | ~v_70) ;
	assign x_1279 = (v_583 | ~v_582) ;
	assign x_1278 = (v_583 | ~v_402) ;
	assign x_1274 = (v_583 | ~v_581) ;
	assign x_1273 = (v_583 | ~v_580) ;
	assign x_1265 = (v_588 | ~v_48) ;
	assign x_1264 = (v_588 | ~v_50) ;
	assign x_1260 = (v_588 | ~v_80) ;
	assign x_1259 = (v_588 | ~v_412) ;
	assign x_1255 = (v_588 | ~v_586) ;
	assign x_1254 = (v_588 | ~v_585) ;
	assign x_1246 = (v_593 | ~v_61) ;
	assign x_1245 = (v_593 | ~v_63) ;
	assign x_1241 = (v_593 | ~v_81) ;
	assign x_1240 = (v_593 | ~v_421) ;
	assign x_1236 = (v_593 | ~v_591) ;
	assign x_1235 = (v_593 | ~v_590) ;
	assign x_1227 = (v_595 | ~v_578) ;
	assign x_1226 = (v_596 | ~v_455) ;
	assign x_1218 = (v_597 | ~v_453) ;
	assign x_1217 = (v_597 | ~v_452) ;
	assign x_1209 = (((((~v_598 | ~v_597) | ~v_596) | ~v_595) | ~v_542) | v_599) ;
	assign x_1208 = ((~v_25 | v_12) | v_600) ;
	assign x_1204 = ((~v_12 | ~v_29) | v_604) ;
	assign x_1203 = ((~v_9 | ~v_41) | v_605) ;
	assign x_1199 = (v_606 | ~v_37) ;
	assign x_1198 = (v_606 | ~v_70) ;
	assign x_1190 = (v_606 | ~v_601) ;
	assign x_1189 = (v_606 | ~v_600) ;
	assign x_1185 = ((~v_21 | ~v_55) | v_609) ;
	assign x_1184 = ((~v_26 | v_12) | v_610) ;
	assign x_1180 = (v_613 | ~v_47) ;
	assign x_1179 = (v_613 | ~v_49) ;
	assign x_1171 = (v_613 | ~v_610) ;
	assign x_1170 = (v_613 | ~v_609) ;
	assign x_1166 = ((~v_27 | v_12) | v_614) ;
	assign x_1165 = ((v_21 | ~v_65) | v_615) ;
	assign x_1161 = ((~v_12 | ~v_30) | v_619) ;
	assign x_1160 = (v_620 | ~v_58) ;
	assign x_1152 = (v_620 | ~v_618) ;
	assign x_1151 = (v_620 | ~v_617) ;
	assign x_1147 = (v_620 | ~v_530) ;
	assign x_1146 = (v_620 | ~v_529) ;
	assign x_1142 = (v_622 | ~v_453) ;
	assign x_1141 = (v_622 | ~v_452) ;
	assign x_1133 = (v_627 | ~v_34) ;
	assign x_1132 = (v_627 | ~v_35) ;
	assign x_1128 = (v_627 | ~v_72) ;
	assign x_1127 = (v_627 | ~v_605) ;
	assign x_1123 = (v_627 | ~v_472) ;
	assign x_1122 = (v_627 | ~v_624) ;
	assign x_1114 = (v_632 | ~v_47) ;
	assign x_1113 = (v_632 | ~v_48) ;
	assign x_1109 = (v_632 | ~v_75) ;
	assign x_1108 = (v_632 | ~v_612) ;
	assign x_1104 = (v_632 | ~v_629) ;
	assign x_1103 = (v_632 | ~v_460) ;
	assign x_1095 = (v_637 | ~v_60) ;
	assign x_1094 = (v_637 | ~v_61) ;
	assign x_1090 = (v_637 | ~v_78) ;
	assign x_1089 = (v_637 | ~v_618) ;
	assign x_1085 = (v_637 | ~v_634) ;
	assign x_1084 = (v_637 | ~v_633) ;
	assign x_1076 = (v_639 | ~v_594) ;
	assign x_1075 = (v_639 | ~v_638) ;
	assign x_1071 = (v_640 | ~v_452) ;
	assign x_1070 = (v_640 | ~v_594) ;
	assign x_1066 = ((~v_17 | ~v_42) | v_643) ;
	assign x_1065 = ((~v_11 | ~v_29) | v_644) ;
	assign x_1057 = (v_645 | ~v_644) ;
	assign x_1056 = (v_645 | ~v_605) ;
	assign x_1052 = (v_645 | ~v_642) ;
	assign x_1051 = (v_645 | ~v_641) ;
	assign x_1047 = ((~v_11 | ~v_28) | v_648) ;
	assign x_1046 = ((~v_26 | v_11) | v_649) ;
	assign x_1038 = (v_650 | ~v_612) ;
	assign x_1037 = (v_650 | ~v_412) ;
	assign x_1033 = (v_650 | ~v_647) ;
	assign x_1032 = (v_650 | ~v_646) ;
	assign x_1028 = ((~v_27 | v_11) | v_653) ;
	assign x_1027 = ((~v_11 | ~v_30) | v_654) ;
	assign x_1019 = (v_655 | ~v_654) ;
	assign x_1018 = (v_655 | ~v_653) ;
	assign x_1014 = (v_655 | ~v_616) ;
	assign x_1013 = (v_655 | ~v_652) ;
	assign x_1009 = (v_657 | ~v_454) ;
	assign x_1008 = (v_657 | ~v_453) ;
	assign x_1000 = (v_658 | ~v_423) ;
	assign x_999 = (((~v_658 | ~v_657) | ~v_640) | v_659) ;
	assign x_995 = (v_660 | ~v_452) ;
	assign x_994 = (v_660 | ~v_621) ;
	assign x_990 = (v_661 | ~v_453) ;
	assign x_989 = (v_661 | ~v_452) ;
	assign x_981 = (v_662 | ~v_656) ;
	assign x_980 = (v_663 | ~v_455) ;
	assign x_976 = (v_663 | ~v_594) ;
	assign x_975 = (((~v_663 | ~v_662) | ~v_661) | v_664) ;
	assign x_971 = (v_665 | ~v_452) ;
	assign x_970 = (v_665 | ~v_638) ;
	assign x_962 = (v_668 | ~v_667) ;
	assign x_961 = (v_668 | ~v_599) ;
	assign x_957 = (v_670 | ~v_453) ;
	assign x_956 = (v_670 | ~v_452) ;
	assign x_952 = (v_671 | ~v_454) ;
	assign x_951 = (v_671 | ~v_453) ;
	assign x_943 = (v_673 | ~v_452) ;
	assign x_942 = (v_673 | ~v_541) ;
	assign x_938 = (v_674 | ~v_453) ;
	assign x_937 = (v_674 | ~v_452) ;
	assign x_933 = (v_675 | ~v_454) ;
	assign x_932 = (v_675 | ~v_453) ;
	assign x_924 = (v_677 | ~v_500) ;
	assign x_923 = (v_677 | ~v_676) ;
	assign x_915 = (v_679 | ~v_454) ;
	assign x_914 = (v_679 | ~v_453) ;
	assign x_906 = (v_680 | ~v_558) ;
	assign x_905 = (((~v_680 | ~v_679) | ~v_678) | v_681) ;
	assign x_901 = (v_682 | ~v_452) ;
	assign x_900 = (v_682 | ~v_594) ;
	assign x_896 = (v_683 | ~v_453) ;
	assign x_895 = (v_683 | ~v_452) ;
	assign x_887 = (v_684 | ~v_621) ;
	assign x_886 = (v_685 | ~v_455) ;
	assign x_882 = (v_685 | ~v_541) ;
	assign x_881 = (((((~v_685 | ~v_684) | ~v_683) | ~v_682) | ~v_677) | v_686) ;
	assign x_877 = (v_688 | ~v_454) ;
	assign x_876 = (v_688 | ~v_453) ;
	assign x_868 = (v_689 | ~v_541) ;
	assign x_867 = (v_689 | ~v_659) ;
	assign x_863 = (v_692 | ~v_4) ;
	assign x_862 = (v_692 | ~v_5) ;
	assign x_858 = (v_693 | ~v_2) ;
	assign x_857 = (v_693 | ~v_3) ;
	assign x_849 = (v_697 | v_29) ;
	assign x_848 = (v_698 | v_14) ;
	assign x_844 = (v_700 | v_26) ;
	assign x_843 = (v_701 | ~v_14) ;
	assign x_839 = (v_703 | v_14) ;
	assign x_838 = (v_703 | v_55) ;
	assign x_830 = (v_708 | v_14) ;
	assign x_829 = (v_708 | v_68) ;
	assign x_825 = (v_710 | ~v_699) ;
	assign x_824 = (((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_710) | v_711) ;
	assign x_820 = (v_715 | ~v_714) ;
	assign x_819 = (v_715 | ~v_713) ;
	assign x_811 = (v_720 | ~v_717) ;
	assign x_810 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_214) | ~v_720) | v_721) ;
	assign x_806 = (v_725 | ~v_724) ;
	assign x_805 = (v_725 | ~v_723) ;
	assign x_801 = ((~v_725 | ~v_383) | v_726) ;
	assign x_800 = (v_727 | ~v_360) ;
	assign x_792 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_255) | ~v_728) | v_729) ;
	assign x_791 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_148) | ~v_720) | v_730) ;
	assign x_787 = (v_731 | ~v_730) ;
	assign x_786 = (v_731 | ~v_729) ;
	assign x_782 = (v_735 | ~v_719) ;
	assign x_781 = (v_735 | ~v_718) ;
	assign x_773 = (v_737 | ~v_711) ;
	assign x_772 = (((((~v_389 | ~v_388) | ~v_737) | ~v_92) | ~v_91) | v_738) ;
	assign x_764 = (v_743 | ~v_36) ;
	assign x_763 = (v_743 | ~v_37) ;
	assign x_755 = (v_743 | ~v_741) ;
	assign x_754 = (v_743 | ~v_740) ;
	assign x_750 = ((~v_14 | ~v_28) | v_746) ;
	assign x_749 = ((~v_14 | ~v_55) | v_747) ;
	assign x_745 = (v_748 | ~v_49) ;
	assign x_744 = (v_748 | ~v_50) ;
	assign x_736 = (v_748 | ~v_746) ;
	assign x_735 = (v_748 | ~v_745) ;
	assign x_731 = ((~v_14 | ~v_30) | v_751) ;
	assign x_730 = ((~v_14 | ~v_68) | v_752) ;
	assign x_726 = (v_753 | ~v_62) ;
	assign x_725 = (v_753 | ~v_63) ;
	assign x_717 = (v_753 | ~v_751) ;
	assign x_716 = (v_753 | ~v_750) ;
	assign x_712 = (v_755 | ~v_454) ;
	assign x_711 = (v_755 | ~v_453) ;
	assign x_707 = (v_756 | ~v_454) ;
	assign x_706 = (v_756 | ~v_453) ;
	assign x_698 = (v_757 | ~v_451) ;
	assign x_697 = (v_757 | ~v_638) ;
	assign x_693 = (v_758 | ~v_452) ;
	assign x_692 = (v_758 | ~v_575) ;
	assign x_688 = (v_760 | ~v_453) ;
	assign x_687 = (v_760 | ~v_452) ;
	assign x_679 = (v_761 | ~v_621) ;
	assign x_678 = (v_762 | ~v_455) ;
	assign x_674 = (v_762 | ~v_575) ;
	assign x_673 = (v_762 | ~v_656) ;
	assign x_669 = (v_763 | ~v_452) ;
	assign x_668 = (v_763 | ~v_638) ;
	assign x_660 = (v_766 | ~v_455) ;
	assign x_659 = (v_766 | ~v_454) ;
	assign x_655 = (v_766 | ~v_423) ;
	assign x_654 = (v_767 | ~v_455) ;
	assign x_650 = (v_767 | ~v_517) ;
	assign x_649 = (v_767 | ~v_638) ;
	assign x_641 = (v_770 | ~v_686) ;
	assign x_640 = (((((~v_663 | ~v_662) | ~v_661) | ~v_689) | ~v_688) | v_771) ;
	assign x_636 = (v_773 | ~v_453) ;
	assign x_635 = (v_773 | ~v_452) ;
	assign x_631 = (v_774 | ~v_454) ;
	assign x_630 = (v_774 | ~v_453) ;
	assign x_622 = (v_777 | ~v_454) ;
	assign x_621 = (v_777 | ~v_453) ;
	assign x_613 = (v_778 | ~v_621) ;
	assign x_612 = (v_778 | ~v_772) ;
	assign x_604 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_255) | ~v_216) | v_784) ;
	assign x_603 = (v_785 | ~v_295) ;
	assign x_599 = (v_787 | ~v_274) ;
	assign x_598 = (v_787 | ~v_273) ;
	assign x_594 = ((~v_787 | ~v_727) | v_788) ;
	assign x_593 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_275) | ~v_120) | v_789) ;
	assign x_585 = (v_793 | ~v_295) ;
	assign x_584 = (v_793 | ~v_294) ;
	assign x_580 = (v_793 | ~v_792) ;
	assign x_579 = (v_793 | ~v_788) ;
	assign x_575 = (v_795 | ~v_453) ;
	assign x_574 = (v_795 | ~v_452) ;
	assign x_566 = (v_797 | ~v_796) ;
	assign x_565 = (v_797 | ~v_575) ;
	assign x_561 = (v_800 | ~v_455) ;
	assign x_560 = (v_800 | ~v_454) ;
	assign x_556 = (v_800 | ~v_423) ;
	assign x_555 = (v_801 | ~v_455) ;
	assign x_547 = (v_803 | ~v_686) ;
	assign x_546 = ((((((((~v_598 | ~v_597) | ~v_596) | ~v_595) | ~v_542) | ~v_803) | ~v_799) | ~v_395) | v_804) ;
	assign x_542 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_378) | ~v_353) | v_807) ;
	assign x_541 = (v_808 | ~v_382) ;
	assign x_537 = (v_810 | ~v_372) ;
	assign x_536 = (v_810 | ~v_809) ;
	assign x_528 = (v_814 | ~v_376) ;
	assign x_527 = (v_814 | ~v_375) ;
	assign x_523 = (v_816 | ~v_382) ;
	assign x_522 = (v_816 | ~v_381) ;
	assign x_518 = (v_816 | ~v_815) ;
	assign x_517 = (v_816 | ~v_811) ;
	assign x_509 = (((~v_685 | ~v_684) | ~v_683) | v_819) ;
	assign x_508 = (v_820 | ~v_455) ;
	assign x_504 = (v_820 | ~v_819) ;
	assign x_503 = (v_820 | ~v_638) ;
	assign x_499 = (v_823 | ~v_455) ;
	assign x_498 = (v_823 | ~v_454) ;
	assign x_490 = (v_824 | ~v_452) ;
	assign x_489 = (v_824 | ~v_575) ;
	assign x_485 = (v_826 | ~v_771) ;
	assign x_484 = ((((((((~v_685 | ~v_684) | ~v_683) | ~v_682) | ~v_677) | ~v_826) | ~v_822) | ~v_395) | v_827) ;
	assign x_480 = ((~v_735 | ~v_727) | v_830) ;
	assign x_479 = ((~v_810 | ~v_369) | v_831) ;
	assign x_471 = (((((~v_389 | ~v_388) | ~v_832) | ~v_92) | ~v_91) | v_833) ;
	assign x_470 = (v_834 | ~v_779) ;
	assign x_462 = ((~v_791 | ~v_735) | v_839) ;
	assign x_461 = ((~v_731 | ~v_369) | v_840) ;
	assign x_453 = (((((~v_389 | ~v_388) | ~v_841) | ~v_92) | ~v_91) | v_842) ;
	assign x_452 = (v_843 | ~v_802) ;
	assign x_448 = ((((((((~v_768 | ~v_767) | ~v_766) | ~v_765) | ~v_760) | ~v_844) | ~v_843) | ~v_395) | v_845) ;
	assign x_447 = (v_846 | ~v_845) ;
	assign x_443 = ((~v_787 | ~v_369) | v_849) ;
	assign x_442 = (v_850 | ~v_215) ;
	assign x_434 = (v_852 | ~v_599) ;
	assign x_433 = (v_852 | ~v_769) ;
	assign x_429 = (v_855 | ~v_854) ;
	assign x_428 = (v_855 | ~v_851) ;
	assign x_424 = (v_859 | ~v_355) ;
	assign x_423 = (v_859 | ~v_354) ;
	assign x_415 = (v_861 | ~v_667) ;
	assign x_414 = (v_862 | ~v_769) ;
	assign x_410 = (v_864 | ~v_860) ;
	assign x_409 = ((((((((v_7 | v_4) | v_6) | v_8) | v_3) | v_2) | ~v_693) | ~v_692) | ~v_864) ;
	assign x_405 = (v_867 | v_29) ;
	assign x_404 = (v_868 | v_24) ;
	assign x_396 = (v_872 | v_52) ;
	assign x_395 = (v_873 | v_24) ;
	assign x_391 = (((((((((((((((v_50 | v_49) | v_74) | v_86) | v_80) | v_44) | ~v_222) | v_89) | ~v_108) | ~v_107) | ~v_219) | ~v_874) | ~v_873) | ~v_872) | ~v_871) | v_875) ;
	assign x_390 = (v_876 | ~v_24) ;
	assign x_386 = (v_878 | v_24) ;
	assign x_385 = (v_878 | v_30) ;
	assign x_377 = ((~v_814 | ~v_369) | v_883) ;
	assign x_376 = ((~v_791 | ~v_810) | v_884) ;
	assign x_372 = (v_885 | ~v_882) ;
	assign x_371 = (((((~v_389 | ~v_388) | ~v_885) | ~v_92) | ~v_91) | v_886) ;
	assign x_367 = ((~v_25 | v_24) | v_890) ;
	assign x_366 = (v_891 | ~v_31) ;
	assign x_358 = (v_891 | ~v_539) ;
	assign x_357 = (v_891 | ~v_401) ;
	assign x_353 = (v_891 | ~v_888) ;
	assign x_352 = (v_891 | ~v_887) ;
	assign x_348 = ((~v_24 | ~v_55) | v_895) ;
	assign x_347 = (v_896 | ~v_44) ;
	assign x_339 = (v_896 | ~v_411) ;
	assign x_338 = (v_896 | ~v_410) ;
	assign x_334 = (v_896 | ~v_893) ;
	assign x_333 = (v_896 | ~v_892) ;
	assign x_329 = ((~v_24 | ~v_68) | v_900) ;
	assign x_328 = (v_901 | ~v_57) ;
	assign x_320 = (v_901 | ~v_418) ;
	assign x_319 = (v_901 | ~v_530) ;
	assign x_311 = (v_903 | ~v_454) ;
	assign x_310 = (v_903 | ~v_453) ;
	assign x_302 = (v_907 | ~v_906) ;
	assign x_301 = (v_907 | ~v_886) ;
	assign x_297 = (v_910 | v_19) ;
	assign x_296 = (v_910 | v_29) ;
	assign x_292 = (v_912 | v_42) ;
	assign x_291 = (((((((((((((((v_31 | v_35) | v_37) | v_36) | v_34) | v_79) | v_71) | ~v_127) | ~v_99) | ~v_912) | ~v_911) | ~v_121) | ~v_96) | ~v_910) | ~v_909) | v_913) ;
	assign x_283 = (v_917 | v_26) ;
	assign x_282 = (((((((((((((((v_50 | v_49) | v_48) | v_74) | v_47) | v_80) | v_44) | ~v_109) | ~v_917) | ~v_131) | ~v_130) | ~v_106) | ~v_916) | ~v_915) | ~v_914) | v_918) ;
	assign x_278 = (v_920 | v_68) ;
	assign x_277 = (v_921 | ~v_19) ;
	assign x_273 = (((((((((((((((v_61 | v_81) | v_63) | v_62) | v_60) | v_57) | v_77) | ~v_118) | ~v_922) | ~v_143) | ~v_921) | ~v_116) | ~v_139) | ~v_920) | ~v_919) | v_923) ;
	assign x_272 = (v_924 | ~v_923) ;
	assign x_264 = (v_927 | ~v_925) ;
	assign x_263 = (((((~v_389 | ~v_388) | ~v_927) | ~v_92) | ~v_91) | v_928) ;
	assign x_259 = ((~v_19 | ~v_42) | v_932) ;
	assign x_258 = (v_933 | ~v_31) ;
	assign x_254 = (v_933 | ~v_37) ;
	assign x_253 = (v_933 | ~v_71) ;
	assign x_245 = (v_933 | ~v_930) ;
	assign x_244 = (v_933 | ~v_929) ;
	assign x_240 = ((~v_26 | v_19) | v_937) ;
	assign x_239 = (v_938 | ~v_44) ;
	assign x_235 = (v_938 | ~v_50) ;
	assign x_234 = (v_938 | ~v_74) ;
	assign x_226 = (v_938 | ~v_935) ;
	assign x_225 = (v_938 | ~v_934) ;
	assign x_221 = ((v_19 | ~v_65) | v_942) ;
	assign x_220 = (v_943 | ~v_57) ;
	assign x_216 = (v_943 | ~v_63) ;
	assign x_215 = (v_943 | ~v_77) ;
	assign x_207 = (v_943 | ~v_940) ;
	assign x_206 = (v_943 | ~v_939) ;
	assign x_202 = (v_945 | ~v_453) ;
	assign x_201 = (v_945 | ~v_452) ;
	assign x_197 = (((((~v_946 | ~v_904) | ~v_776) | ~v_945) | ~v_395) | v_947) ;
	assign x_196 = (v_948 | ~v_947) ;
	assign x_188 = (v_952 | ~v_730) ;
	assign x_187 = (v_952 | ~v_729) ;
	assign x_183 = (v_954 | ~v_798) ;
	assign x_182 = (v_954 | ~v_779) ;
	assign x_178 = (v_957 | ~v_956) ;
	assign x_177 = (v_957 | ~v_953) ;
	assign x_169 = (v_961 | ~v_784) ;
	assign x_168 = (v_961 | ~v_960) ;
	assign x_160 = (v_966 | ~v_965) ;
	assign x_159 = (v_966 | ~v_962) ;
	assign x_151 = (v_970 | ~v_812) ;
	assign x_150 = (v_970 | ~v_969) ;
	assign x_146 = (v_972 | ~v_798) ;
	assign x_145 = (v_973 | ~v_775) ;
	assign x_141 = (v_975 | ~v_971) ;
	assign x_140 = ((((((((v_7 | v_5) | v_6) | v_8) | v_3) | v_1) | ~v_693) | ~v_692) | ~v_975) ;
	assign x_132 = (v_979 | ~v_978) ;
	assign x_131 = (v_979 | ~v_977) ;
	assign x_127 = (v_982 | ~v_667) ;
	assign x_126 = (v_982 | ~v_825) ;
	assign x_122 = ((((((((v_5 | v_6) | v_8) | v_3) | v_2) | v_1) | ~v_693) | ~v_692) | ~v_984) ;
	assign x_121 = ((~v_364 | ~v_731) | v_986) ;
	assign x_113 = (v_988 | ~v_986) ;
	assign x_112 = (((((~v_389 | ~v_388) | ~v_988) | ~v_92) | ~v_91) | v_989) ;
	assign x_108 = (v_991 | ~v_769) ;
	assign x_107 = ((((((((~v_763 | ~v_762) | ~v_761) | ~v_778) | ~v_777) | ~v_991) | ~v_990) | ~v_395) | v_992) ;
	assign x_103 = (v_995 | v_9) ;
	assign x_102 = (v_995 | v_42) ;
	assign x_94 = (v_1000 | ~v_9) ;
	assign x_93 = (v_1000 | v_52) ;
	assign x_89 = (v_1002 | v_26) ;
	assign x_88 = (v_1003 | v_9) ;
	assign x_84 = (v_1005 | v_65) ;
	assign x_83 = (v_1006 | ~v_9) ;
	assign x_75 = (v_1010 | ~v_1004) ;
	assign x_74 = (v_1010 | ~v_999) ;
	assign x_70 = (v_1012 | ~v_736) ;
	assign x_69 = (v_1012 | ~v_1011) ;
	assign x_65 = ((~v_9 | ~v_29) | v_1016) ;
	assign x_64 = ((~v_25 | v_9) | v_1017) ;
	assign x_56 = (v_1018 | ~v_1017) ;
	assign x_55 = (v_1018 | ~v_605) ;
	assign x_51 = (v_1018 | ~v_428) ;
	assign x_50 = (v_1018 | ~v_427) ;
	assign x_46 = ((~v_26 | v_9) | v_1021) ;
	assign x_45 = ((~v_9 | ~v_28) | v_1022) ;
	assign x_37 = (v_1023 | ~v_50) ;
	assign x_36 = (v_1023 | ~v_612) ;
	assign x_32 = (v_1023 | ~v_608) ;
	assign x_31 = (v_1023 | ~v_437) ;
	assign x_27 = ((~v_9 | ~v_68) | v_1026) ;
	assign x_26 = ((~v_9 | ~v_30) | v_1027) ;
	assign x_18 = (v_1028 | ~v_63) ;
	assign x_17 = (v_1028 | ~v_1026) ;
	assign x_9 = (v_1030 | ~v_455) ;
	assign x_8 = (v_1030 | ~v_454) ;
	assign x_4824 = (x_2417 & x_2418) ;
	assign x_2416 = (v_91 | ~v_23) ;
	assign x_2415 = (v_91 | ~v_24) ;
	assign x_2414 = (v_92 | ~v_13) ;
	assign x_4820 = (x_2412 & x_2413) ;
	assign x_2411 = (v_92 | ~v_16) ;
	assign x_2410 = (v_93 | ~v_23) ;
	assign x_2409 = (v_93 | v_25) ;
	assign x_4815 = (x_2407 & x_2408) ;
	assign x_2406 = (v_95 | v_20) ;
	assign x_2405 = (v_95 | v_42) ;
	assign x_2404 = (v_96 | ~v_19) ;
	assign x_2403 = (v_96 | v_40) ;
	assign x_2402 = (v_97 | ~v_24) ;
	assign x_2401 = (v_97 | v_38) ;
	assign x_2400 = (v_98 | v_24) ;
	assign x_4806 = (x_2398 & x_2399) ;
	assign x_2397 = (v_99 | v_43) ;
	assign x_2396 = (v_100 | ~v_20) ;
	assign x_2395 = (v_100 | v_39) ;
	assign x_4802 = (x_2393 & x_2394) ;
	assign x_2392 = (v_102 | v_26) ;
	assign x_2391 = (v_103 | ~v_20) ;
	assign x_2390 = (v_103 | v_52) ;
	assign x_4797 = (x_2388 & x_2389) ;
	assign x_2387 = (v_105 | v_20) ;
	assign x_2386 = (v_105 | v_55) ;
	assign x_2385 = (v_106 | ~v_19) ;
	assign x_2384 = (v_106 | v_53) ;
	assign x_2383 = (v_107 | ~v_24) ;
	assign x_2382 = (v_107 | v_51) ;
	assign x_2381 = (v_108 | v_24) ;
	assign x_4787 = (x_2379 & x_2380) ;
	assign x_2378 = (v_109 | v_56) ;
	assign x_2377 = (((((((((((((((v_49 | v_48) | v_74) | v_73) | v_83) | v_80) | v_89) | ~v_109) | ~v_108) | ~v_107) | ~v_106) | ~v_105) | ~v_104) | ~v_103) | ~v_102) | v_110) ;
	assign x_2376 = (v_111 | ~v_23) ;
	assign x_4783 = (x_2374 & x_2375) ;
	assign x_2373 = (v_112 | v_65) ;
	assign x_2372 = (v_113 | v_23) ;
	assign x_2371 = (v_113 | v_30) ;
	assign x_4778 = (x_2369 & x_2370) ;
	assign x_2368 = (v_115 | ~v_24) ;
	assign x_2367 = (v_115 | v_64) ;
	assign x_2366 = (v_116 | ~v_19) ;
	assign x_2365 = (v_116 | v_66) ;
	assign x_2364 = (v_117 | v_24) ;
	assign x_2363 = (v_117 | v_67) ;
	assign x_2362 = (v_118 | v_19) ;
	assign x_4769 = (x_2360 & x_2361) ;
	assign x_2359 = (v_120 | ~v_119) ;
	assign x_2358 = (v_120 | ~v_110) ;
	assign x_2357 = (v_120 | ~v_101) ;
	assign x_4765 = (x_2355 & x_2356) ;
	assign x_2354 = (v_122 | ~v_17) ;
	assign x_2353 = (v_122 | v_25) ;
	assign x_2352 = (v_123 | v_17) ;
	assign x_4760 = (x_2350 & x_2351) ;
	assign x_2349 = (v_124 | v_40) ;
	assign x_2348 = (v_125 | v_9) ;
	assign x_2347 = (v_125 | v_43) ;
	assign x_2346 = (v_126 | ~v_11) ;
	assign x_2345 = (v_126 | v_39) ;
	assign x_2344 = (v_127 | v_19) ;
	assign x_2343 = (v_127 | v_41) ;
	assign x_4749 = (x_2341 & x_2342) ;
	assign x_2340 = (((((((((((((((v_33 | v_35) | v_37) | v_36) | v_34) | v_79) | v_70) | ~v_128) | ~v_127) | ~v_126) | ~v_125) | ~v_124) | ~v_123) | ~v_122) | ~v_121) | v_129) ;
	assign x_2339 = (v_130 | ~v_19) ;
	assign x_2338 = (v_130 | v_51) ;
	assign x_4745 = (x_2336 & x_2337) ;
	assign x_2335 = (v_132 | ~v_17) ;
	assign x_2334 = (v_132 | v_26) ;
	assign x_2333 = (v_133 | ~v_11) ;
	assign x_4740 = (x_2331 & x_2332) ;
	assign x_2330 = (v_134 | v_53) ;
	assign x_2329 = (v_135 | v_17) ;
	assign x_2328 = (v_135 | v_28) ;
	assign x_2327 = (v_136 | v_11) ;
	assign x_2326 = (v_136 | v_55) ;
	assign x_2325 = (v_137 | v_9) ;
	assign x_2324 = (v_137 | v_56) ;
	assign x_4731 = (x_2322 & x_2323) ;
	assign x_2321 = (v_139 | v_67) ;
	assign x_2320 = (v_140 | ~v_11) ;
	assign x_2319 = (v_140 | v_65) ;
	assign x_4727 = (x_2317 & x_2318) ;
	assign x_2316 = (v_142 | v_9) ;
	assign x_2315 = (v_142 | v_69) ;
	assign x_2314 = (v_143 | ~v_19) ;
	assign x_4722 = (x_2312 & x_2313) ;
	assign x_2311 = (v_144 | v_27) ;
	assign x_2310 = (v_145 | v_11) ;
	assign x_2309 = (v_145 | v_68) ;
	assign x_2308 = (v_146 | v_17) ;
	assign x_2307 = (v_146 | v_30) ;
	assign x_2306 = (((((((((((((((v_61 | v_76) | v_81) | v_63) | v_62) | v_60) | v_59) | ~v_146) | ~v_145) | ~v_144) | ~v_143) | ~v_142) | ~v_141) | ~v_140) | ~v_139) | v_147) ;
	assign x_2305 = (v_148 | ~v_147) ;
	assign x_4712 = (x_2303 & x_2304) ;
	assign x_2302 = (v_149 | ~v_30) ;
	assign x_2301 = (v_149 | v_28) ;
	assign x_2300 = (v_150 | ~v_25) ;
	assign x_4708 = (x_2298 & x_2299) ;
	assign x_2297 = (v_151 | v_29) ;
	assign x_2296 = (v_152 | ~v_26) ;
	assign x_2295 = (v_152 | v_27) ;
	assign x_4703 = (x_2293 & x_2294) ;
	assign x_2292 = (v_154 | v_26) ;
	assign x_2291 = (v_155 | ~v_16) ;
	assign x_2290 = (v_155 | v_52) ;
	assign x_2289 = (v_156 | v_16) ;
	assign x_2288 = (v_156 | v_55) ;
	assign x_2287 = (v_157 | ~v_14) ;
	assign x_2286 = (v_157 | v_53) ;
	assign x_4694 = (x_2284 & x_2285) ;
	assign x_2283 = (v_159 | v_22) ;
	assign x_2282 = (v_159 | v_28) ;
	assign x_2281 = (((((((((((((((v_50 | v_49) | v_48) | v_74) | v_73) | v_80) | v_89) | ~v_159) | ~v_158) | ~v_157) | ~v_108) | ~v_107) | ~v_156) | ~v_155) | ~v_154) | v_160) ;
	assign x_4690 = (x_2279 & x_2280) ;
	assign x_2278 = (v_162 | ~v_16) ;
	assign x_2277 = (v_162 | v_65) ;
	assign x_2276 = (v_163 | v_16) ;
	assign x_4685 = (x_2274 & x_2275) ;
	assign x_2273 = (v_164 | v_69) ;
	assign x_2272 = (v_165 | ~v_14) ;
	assign x_2271 = (v_165 | v_66) ;
	assign x_2270 = (v_166 | v_22) ;
	assign x_2269 = (v_166 | v_30) ;
	assign x_2268 = (((((((((((((((v_61 | v_76) | v_81) | v_63) | v_62) | v_77) | ~v_166) | ~v_117) | v_90) | ~v_165) | ~v_164) | ~v_115) | ~v_163) | ~v_162) | ~v_161) | v_167) ;
	assign x_2267 = (v_168 | v_22) ;
	assign x_4673 = (x_2265 & x_2266) ;
	assign x_2264 = (v_169 | v_40) ;
	assign x_2263 = (v_170 | v_16) ;
	assign x_2262 = (v_170 | v_42) ;
	assign x_4669 = (x_2260 & x_2261) ;
	assign x_2259 = (v_172 | ~v_22) ;
	assign x_2258 = (v_172 | v_25) ;
	assign x_2257 = (v_173 | v_14) ;
	assign x_4664 = (x_2255 & x_2256) ;
	assign x_2254 = (v_175 | ~v_174) ;
	assign x_2253 = (v_175 | ~v_167) ;
	assign x_2252 = (v_175 | ~v_160) ;
	assign x_2251 = (v_176 | ~v_14) ;
	assign x_2250 = (v_176 | v_38) ;
	assign x_2249 = (v_177 | ~v_13) ;
	assign x_2248 = (v_177 | v_25) ;
	assign x_4655 = (x_2246 & x_2247) ;
	assign x_2245 = (v_179 | v_14) ;
	assign x_2244 = (v_179 | v_41) ;
	assign x_2243 = (v_180 | v_13) ;
	assign x_4651 = (x_2241 & x_2242) ;
	assign x_2240 = (v_181 | v_42) ;
	assign x_2239 = (((((((((((((((v_33 | v_35) | v_36) | v_34) | v_79) | v_70) | v_82) | ~v_181) | ~v_180) | ~v_179) | ~v_178) | ~v_177) | ~v_176) | ~v_125) | ~v_124) | v_182) ;
	assign x_2238 = (v_183 | ~v_14) ;
	assign x_4646 = (x_2236 & x_2237) ;
	assign x_2235 = (v_184 | v_26) ;
	assign x_2234 = (v_185 | ~v_10) ;
	assign x_2233 = (v_185 | v_52) ;
	assign x_2232 = (v_186 | v_14) ;
	assign x_2231 = (v_186 | v_54) ;
	assign x_2230 = (v_187 | v_13) ;
	assign x_2229 = (v_187 | v_28) ;
	assign x_4636 = (x_2227 & x_2228) ;
	assign x_2226 = (((((((((((((((v_49 | v_48) | v_46) | v_47) | v_73) | v_83) | v_80) | ~v_137) | ~v_188) | ~v_187) | ~v_186) | ~v_185) | ~v_184) | ~v_183) | ~v_134) | v_189) ;
	assign x_2225 = (v_190 | ~v_14) ;
	assign x_2224 = (v_190 | v_64) ;
	assign x_4632 = (x_2222 & x_2223) ;
	assign x_2221 = (v_192 | ~v_10) ;
	assign x_2220 = (v_192 | v_65) ;
	assign x_2219 = (v_193 | v_13) ;
	assign x_4627 = (x_2217 & x_2218) ;
	assign x_2216 = (v_194 | v_67) ;
	assign x_2215 = (v_195 | v_10) ;
	assign x_2214 = (v_195 | v_68) ;
	assign x_2213 = (((((((((((((((v_61 | v_76) | v_81) | v_62) | v_60) | v_59) | v_84) | ~v_195) | ~v_194) | ~v_193) | ~v_192) | ~v_191) | ~v_190) | ~v_142) | ~v_141) | v_196) ;
	assign x_2212 = (v_197 | ~v_196) ;
	assign x_2211 = (v_197 | ~v_189) ;
	assign x_2210 = (v_197 | ~v_182) ;
	assign x_4618 = (x_2208 & x_2209) ;
	assign x_2207 = (v_199 | v_25) ;
	assign x_2206 = (v_200 | v_21) ;
	assign x_2205 = (v_200 | v_29) ;
	assign x_4614 = (x_2203 & x_2204) ;
	assign x_2202 = (v_202 | ~v_12) ;
	assign x_2201 = (v_202 | v_39) ;
	assign x_2200 = (((((((((((((((v_33 | v_35) | v_37) | v_36) | v_79) | v_70) | v_88) | ~v_202) | ~v_201) | ~v_125) | ~v_124) | ~v_200) | ~v_199) | ~v_98) | ~v_97) | v_203) ;
	assign x_4609 = (x_2198 & x_2199) ;
	assign x_2197 = (v_205 | ~v_12) ;
	assign x_2196 = (v_205 | v_52) ;
	assign x_2195 = (v_206 | v_21) ;
	assign x_2194 = (v_206 | v_28) ;
	assign x_2193 = (v_207 | v_12) ;
	assign x_2192 = (v_207 | v_55) ;
	assign x_2191 = (((((((((((((((v_50 | v_49) | v_48) | v_46) | v_73) | v_80) | ~v_137) | v_89) | ~v_207) | ~v_134) | ~v_206) | ~v_205) | ~v_204) | ~v_108) | ~v_107) | v_208) ;
	assign x_4598 = (x_2189 & x_2190) ;
	assign x_2188 = (v_210 | v_21) ;
	assign x_2187 = (v_210 | v_30) ;
	assign x_2186 = (v_211 | ~v_12) ;
	assign x_4594 = (x_2184 & x_2185) ;
	assign x_2183 = (v_212 | v_68) ;
	assign x_2182 = (((((((((((((((v_61 | v_76) | v_81) | v_63) | v_62) | v_59) | ~v_212) | ~v_117) | v_90) | ~v_211) | ~v_142) | ~v_141) | ~v_210) | ~v_209) | ~v_115) | v_213) ;
	assign x_2181 = (v_214 | ~v_213) ;
	assign x_4589 = (x_2179 & x_2180) ;
	assign x_2178 = (((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_214) | v_215) ;
	assign x_2177 = (v_216 | ~v_215) ;
	assign x_2176 = (v_216 | ~v_198) ;
	assign x_2175 = (v_216 | ~v_153) ;
	assign x_2174 = (v_217 | ~v_16) ;
	assign x_2173 = (v_217 | v_26) ;
	assign x_2172 = (v_218 | ~v_22) ;
	assign x_4580 = (x_2170 & x_2171) ;
	assign x_2169 = (v_219 | v_53) ;
	assign x_2168 = (v_220 | v_22) ;
	assign x_2167 = (v_220 | v_55) ;
	assign x_4576 = (x_2165 & x_2166) ;
	assign x_2164 = (v_222 | v_24) ;
	assign x_2163 = (v_222 | v_56) ;
	assign x_2162 = (((((((((((((((v_50 | v_49) | v_74) | v_47) | v_73) | v_86) | v_80) | ~v_222) | ~v_221) | ~v_220) | ~v_186) | ~v_183) | ~v_219) | ~v_218) | ~v_217) | v_223) ;
	assign x_4571 = (x_2160 & x_2161) ;
	assign x_2159 = (v_225 | v_16) ;
	assign x_2158 = (v_225 | v_30) ;
	assign x_2157 = (v_226 | ~v_24) ;
	assign x_2156 = (v_226 | v_66) ;
	assign x_2155 = (v_227 | v_24) ;
	assign x_2154 = (v_227 | v_69) ;
	assign x_2153 = (v_228 | ~v_16) ;
	assign x_4561 = (x_2151 & x_2152) ;
	assign x_2150 = (v_229 | v_68) ;
	assign x_2149 = (((((((((((((((v_76 | v_81) | v_63) | v_62) | v_60) | v_77) | ~v_229) | v_87) | ~v_194) | ~v_228) | ~v_190) | ~v_227) | ~v_226) | ~v_225) | ~v_224) | v_230) ;
	assign x_2148 = (v_231 | ~v_16) ;
	assign x_4557 = (x_2146 & x_2147) ;
	assign x_2145 = (v_232 | v_39) ;
	assign x_2144 = (v_233 | v_16) ;
	assign x_2143 = (v_233 | v_29) ;
	assign x_4552 = (x_2141 & x_2142) ;
	assign x_2140 = (v_235 | v_22) ;
	assign x_2139 = (v_235 | v_42) ;
	assign x_2138 = (v_236 | v_24) ;
	assign x_2137 = (v_236 | v_43) ;
	assign x_2136 = (((((((((((((((v_37 | v_36) | v_34) | v_79) | v_71) | v_70) | v_85) | ~v_236) | ~v_235) | ~v_179) | ~v_176) | ~v_234) | ~v_233) | ~v_232) | ~v_231) | v_237) ;
	assign x_2135 = (v_238 | ~v_237) ;
	assign x_2134 = (v_238 | ~v_230) ;
	assign x_4543 = (x_2132 & x_2133) ;
	assign x_2131 = (v_240 | ~v_23) ;
	assign x_2130 = (v_240 | v_39) ;
	assign x_2129 = (v_241 | v_20) ;
	assign x_2128 = (v_241 | v_29) ;
	assign x_2127 = (v_242 | v_23) ;
	assign x_2126 = (v_242 | v_42) ;
	assign x_2125 = (v_243 | ~v_20) ;
	assign x_4535 = (x_2123 & x_2124) ;
	assign x_2122 = (v_245 | ~v_20) ;
	assign x_2121 = (v_245 | v_26) ;
	assign x_2120 = (v_246 | ~v_23) ;
	assign x_2119 = (v_246 | v_52) ;
	assign x_2118 = (v_247 | v_23) ;
	assign x_2117 = (v_247 | v_55) ;
	assign x_2116 = (v_248 | v_20) ;
	assign x_4522 = (x_2114 & x_2115) ;
	assign x_2113 = (v_250 | ~v_20) ;
	assign x_2112 = (v_250 | v_27) ;
	assign x_2111 = (v_251 | ~v_23) ;
	assign x_4518 = (x_2109 & x_2110) ;
	assign x_2108 = (v_252 | v_68) ;
	assign x_2107 = (v_253 | v_20) ;
	assign x_2106 = (v_253 | v_30) ;
	assign x_4513 = (x_2104 & x_2105) ;
	assign x_2103 = (v_255 | ~v_249) ;
	assign x_2102 = (v_255 | ~v_244) ;
	assign x_2101 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_214) | ~v_255) | v_256) ;
	assign x_2100 = (v_257 | ~v_15) ;
	assign x_2099 = (v_257 | v_39) ;
	assign x_2098 = (v_258 | v_15) ;
	assign x_2097 = (v_258 | v_42) ;
	assign x_4504 = (x_2095 & x_2096) ;
	assign x_2094 = (v_260 | ~v_18) ;
	assign x_2093 = (v_260 | v_25) ;
	assign x_2092 = (((((((((((((((v_35 | v_36) | v_34) | v_79) | v_71) | v_70) | v_82) | ~v_260) | ~v_127) | ~v_173) | ~v_259) | ~v_169) | ~v_121) | ~v_258) | ~v_257) | v_261) ;
	assign x_4500 = (x_2090 & x_2091) ;
	assign x_2089 = (v_263 | ~v_15) ;
	assign x_2088 = (v_263 | v_52) ;
	assign x_2087 = (v_264 | v_15) ;
	assign x_4495 = (x_2085 & x_2086) ;
	assign x_2084 = (v_265 | v_28) ;
	assign x_2083 = (((((((((((((((v_49 | v_48) | v_74) | v_47) | v_73) | v_83) | v_80) | ~v_265) | ~v_158) | ~v_157) | ~v_131) | ~v_130) | ~v_264) | ~v_263) | ~v_262) | v_266) ;
	assign x_2082 = (v_267 | ~v_18) ;
	assign x_2081 = (v_267 | v_27) ;
	assign x_2080 = (v_268 | ~v_15) ;
	assign x_2079 = (v_268 | v_65) ;
	assign x_2078 = (v_269 | v_18) ;
	assign x_4485 = (x_2076 & x_2077) ;
	assign x_2075 = (v_270 | v_68) ;
	assign x_2074 = (((((((((((((((v_61 | v_76) | v_81) | v_62) | v_60) | v_77) | v_84) | ~v_143) | ~v_165) | ~v_164) | ~v_139) | ~v_270) | ~v_269) | ~v_268) | ~v_267) | v_271) ;
	assign x_2073 = (v_272 | ~v_271) ;
	assign x_4481 = (x_2071 & x_2072) ;
	assign x_2070 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_197) | ~v_272) | v_273) ;
	assign x_2069 = (((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_148) | v_274) ;
	assign x_2068 = (v_275 | ~v_274) ;
	assign x_4476 = (x_2066 & x_2067) ;
	assign x_2065 = (v_276 | ~v_18) ;
	assign x_2064 = (v_276 | v_39) ;
	assign x_2063 = (v_277 | v_15) ;
	assign x_2062 = (v_277 | v_29) ;
	assign x_2061 = (v_278 | v_18) ;
	assign x_2060 = (v_278 | v_42) ;
	assign x_2059 = (v_279 | ~v_15) ;
	assign x_4467 = (x_2057 & x_2058) ;
	assign x_2056 = (v_281 | ~v_15) ;
	assign x_2055 = (v_281 | v_26) ;
	assign x_2054 = (v_282 | ~v_18) ;
	assign x_4463 = (x_2052 & x_2053) ;
	assign x_2051 = (v_283 | v_55) ;
	assign x_2050 = (v_284 | v_15) ;
	assign x_2049 = (v_284 | v_28) ;
	assign x_4458 = (x_2047 & x_2048) ;
	assign x_2046 = (v_286 | v_27) ;
	assign x_2045 = (v_287 | ~v_18) ;
	assign x_2044 = (v_287 | v_65) ;
	assign x_2043 = (v_288 | v_18) ;
	assign x_2042 = (v_288 | v_68) ;
	assign x_2041 = (v_289 | v_15) ;
	assign x_2040 = (v_289 | v_30) ;
	assign x_4447 = (x_2038 & x_2039) ;
	assign x_2037 = (v_291 | ~v_285) ;
	assign x_2036 = (v_291 | ~v_280) ;
	assign x_2035 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_291) | ~v_275) | v_292) ;
	assign x_4443 = (x_2033 & x_2034) ;
	assign x_2032 = (((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_197) | v_295) ;
	assign x_2031 = (v_296 | ~v_295) ;
	assign x_2030 = (v_296 | ~v_294) ;
	assign x_4438 = (x_2028 & x_2029) ;
	assign x_2027 = (v_296 | ~v_239) ;
	assign x_2026 = (v_297 | ~v_12) ;
	assign x_2025 = (v_297 | v_25) ;
	assign x_2024 = (v_298 | ~v_21) ;
	assign x_2023 = (v_298 | v_39) ;
	assign x_2022 = (v_299 | v_21) ;
	assign x_2021 = (v_299 | v_42) ;
	assign x_4429 = (x_2019 & x_2020) ;
	assign x_2018 = (v_301 | v_12) ;
	assign x_2017 = (v_301 | v_29) ;
	assign x_2016 = (v_302 | v_9) ;
	assign x_4425 = (x_2014 & x_2015) ;
	assign x_2013 = (v_304 | ~v_21) ;
	assign x_2012 = (v_304 | v_52) ;
	assign x_2011 = (v_305 | ~v_9) ;
	assign x_4420 = (x_2009 & x_2010) ;
	assign x_2008 = (v_306 | v_55) ;
	assign x_2007 = (v_307 | ~v_12) ;
	assign x_2006 = (v_307 | v_26) ;
	assign x_2005 = (v_308 | v_12) ;
	assign x_2004 = (v_308 | v_28) ;
	assign x_2003 = (v_309 | v_9) ;
	assign x_2002 = (v_309 | v_54) ;
	assign x_4410 = (x_2000 & x_2001) ;
	assign x_1999 = (v_311 | v_27) ;
	assign x_1998 = (v_312 | ~v_21) ;
	assign x_1997 = (v_312 | v_65) ;
	assign x_4406 = (x_1995 & x_1996) ;
	assign x_1994 = (v_314 | v_21) ;
	assign x_1993 = (v_314 | v_68) ;
	assign x_1992 = (v_315 | v_9) ;
	assign x_4401 = (x_1990 & x_1991) ;
	assign x_1989 = (v_316 | v_30) ;
	assign x_1988 = (((((((((((((((v_76 | v_63) | v_62) | v_60) | v_58) | v_77) | ~v_316) | v_87) | ~v_315) | ~v_314) | ~v_313) | ~v_312) | ~v_311) | ~v_227) | ~v_226) | v_317) ;
	assign x_1987 = (v_318 | ~v_317) ;
	assign x_1986 = (v_318 | ~v_310) ;
	assign x_1985 = (v_318 | ~v_303) ;
	assign x_1984 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_120) | ~v_318) | v_319) ;
	assign x_1983 = (v_320 | ~v_10) ;
	assign x_4392 = (x_1981 & x_1982) ;
	assign x_1980 = (v_321 | v_39) ;
	assign x_1979 = (v_322 | v_10) ;
	assign x_1978 = (v_322 | v_29) ;
	assign x_1977 = (v_323 | v_13) ;
	assign x_1976 = (v_323 | v_42) ;
	assign x_1975 = (((((((((((((((v_32 | v_35) | v_37) | v_34) | v_72) | v_71) | v_70) | ~v_302) | ~v_173) | ~v_323) | ~v_322) | ~v_169) | ~v_321) | ~v_320) | ~v_300) | v_324) ;
	assign x_1974 = (v_325 | ~v_13) ;
	assign x_4384 = (x_1972 & x_1973) ;
	assign x_1971 = (v_326 | v_28) ;
	assign x_1970 = (v_327 | v_13) ;
	assign x_1969 = (v_327 | v_55) ;
	assign x_1968 = (v_328 | ~v_10) ;
	assign x_1967 = (v_328 | v_26) ;
	assign x_1966 = (((((((((((((((v_50 | v_48) | v_45) | v_75) | v_74) | v_47) | v_73) | ~v_309) | ~v_328) | ~v_327) | ~v_158) | ~v_326) | ~v_157) | ~v_325) | ~v_305) | v_329) ;
	assign x_1965 = (v_330 | ~v_10) ;
	assign x_4372 = (x_1963 & x_1964) ;
	assign x_1962 = (v_331 | v_65) ;
	assign x_1961 = (v_332 | v_10) ;
	assign x_1960 = (v_332 | v_30) ;
	assign x_4368 = (x_1958 & x_1959) ;
	assign x_1957 = (((((((((((((((v_61 | v_76) | v_63) | v_60) | v_58) | v_78) | v_77) | ~v_315) | ~v_333) | ~v_332) | ~v_165) | ~v_331) | ~v_330) | ~v_313) | ~v_164) | v_334) ;
	assign x_1956 = (v_335 | ~v_334) ;
	assign x_1955 = (v_335 | ~v_329) ;
	assign x_4363 = (x_1953 & x_1954) ;
	assign x_1952 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_291) | ~v_175) | v_337) ;
	assign x_1951 = (v_338 | ~v_11) ;
	assign x_1950 = (v_338 | v_25) ;
	assign x_1949 = (v_339 | ~v_17) ;
	assign x_1948 = (v_339 | v_39) ;
	assign x_1947 = (v_340 | v_17) ;
	assign x_1946 = (v_340 | v_42) ;
	assign x_4354 = (x_1944 & x_1945) ;
	assign x_1943 = (((((((((((((((v_32 | v_35) | v_37) | v_36) | v_34) | v_71) | v_70) | ~v_341) | ~v_302) | ~v_99) | ~v_300) | ~v_340) | ~v_339) | ~v_338) | ~v_96) | v_342) ;
	assign x_1942 = (v_343 | ~v_17) ;
	assign x_1941 = (v_343 | v_52) ;
	assign x_4350 = (x_1939 & x_1940) ;
	assign x_1938 = (v_345 | v_11) ;
	assign x_1937 = (v_345 | v_28) ;
	assign x_1936 = (v_346 | ~v_11) ;
	assign x_4345 = (x_1934 & x_1935) ;
	assign x_1933 = (v_348 | ~v_17) ;
	assign x_1932 = (v_348 | v_65) ;
	assign x_1931 = (v_349 | v_17) ;
	assign x_1930 = (v_349 | v_68) ;
	assign x_1929 = (v_350 | ~v_11) ;
	assign x_1928 = (v_350 | v_27) ;
	assign x_1927 = (v_351 | v_11) ;
	assign x_4335 = (x_1925 & x_1926) ;
	assign x_1924 = (v_353 | ~v_352) ;
	assign x_1923 = (v_353 | ~v_347) ;
	assign x_1922 = (v_353 | ~v_342) ;
	assign x_4331 = (x_1920 & x_1921) ;
	assign x_1919 = (v_356 | ~v_355) ;
	assign x_1918 = (v_356 | ~v_354) ;
	assign x_1917 = (v_356 | ~v_337) ;
	assign x_4326 = (x_1915 & x_1916) ;
	assign x_1914 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_197) | ~v_353) | v_359) ;
	assign x_1913 = (((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_291) | v_360) ;
	assign x_1912 = (v_361 | ~v_360) ;
	assign x_1911 = (v_361 | ~v_359) ;
	assign x_1910 = (v_361 | ~v_358) ;
	assign x_1909 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_335) | ~v_361) | v_362) ;
	assign x_1908 = (((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_353) | v_363) ;
	assign x_4317 = (x_1906 & x_1907) ;
	assign x_1905 = (v_364 | ~v_357) ;
	assign x_1904 = (v_364 | ~v_336) ;
	assign x_1903 = (v_364 | ~v_319) ;
	assign x_4313 = (x_1901 & x_1902) ;
	assign x_1900 = (v_366 | ~v_336) ;
	assign x_1899 = (v_366 | ~v_319) ;
	assign x_1898 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_214) | ~v_366) | v_367) ;
	assign x_4308 = (x_1896 & x_1897) ;
	assign x_1895 = (v_369 | ~v_354) ;
	assign x_1894 = (v_369 | ~v_337) ;
	assign x_1893 = (v_369 | ~v_368) ;
	assign x_1892 = (v_369 | ~v_367) ;
	assign x_1891 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_238) | ~v_335) | v_370) ;
	assign x_1890 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_255) | ~v_353) | v_371) ;
	assign x_1889 = (((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_318) | v_372) ;
	assign x_4297 = (x_1887 & x_1888) ;
	assign x_1886 = (v_373 | ~v_370) ;
	assign x_1885 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_197) | ~v_373) | v_374) ;
	assign x_1884 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_238) | ~v_272) | v_375) ;
	assign x_4293 = (x_1882 & x_1883) ;
	assign x_1881 = (v_378 | ~v_377) ;
	assign x_1880 = (v_378 | ~v_376) ;
	assign x_1879 = (v_378 | ~v_375) ;
	assign x_4288 = (x_1877 & x_1878) ;
	assign x_1876 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_197) | ~v_318) | v_381) ;
	assign x_1875 = (((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_238) | v_382) ;
	assign x_1874 = (v_383 | ~v_382) ;
	assign x_1873 = (v_383 | ~v_381) ;
	assign x_1872 = (v_383 | ~v_380) ;
	assign x_1871 = (v_383 | ~v_379) ;
	assign x_1870 = (v_383 | ~v_374) ;
	assign x_4279 = (x_1868 & x_1869) ;
	assign x_1867 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_238) | ~v_356) | v_386) ;
	assign x_1866 = (v_387 | ~v_360) ;
	assign x_1865 = (v_387 | ~v_359) ;
	assign x_4275 = (x_1863 & x_1864) ;
	assign x_1862 = (v_387 | ~v_385) ;
	assign x_1861 = (v_387 | ~v_384) ;
	assign x_1860 = (v_387 | ~v_365) ;
	assign x_4270 = (x_1858 & x_1859) ;
	assign x_1857 = (v_388 | ~v_19) ;
	assign x_1856 = (v_388 | ~v_20) ;
	assign x_1855 = (v_389 | ~v_9) ;
	assign x_1854 = (v_389 | ~v_10) ;
	assign x_1853 = (v_389 | ~v_11) ;
	assign x_1852 = (v_389 | ~v_12) ;
	assign x_1851 = (((((~v_389 | ~v_388) | ~v_387) | ~v_92) | ~v_91) | v_390) ;
	assign x_4260 = (x_1849 & x_1850) ;
	assign x_1848 = ((((v_20 | v_19) | v_18) | v_17) | v_393) ;
	assign x_1847 = ((((v_9 | v_12) | v_11) | v_10) | v_394) ;
	assign x_1846 = (v_395 | ~v_394) ;
	assign x_4256 = (x_1844 & x_1845) ;
	assign x_1843 = (v_395 | ~v_391) ;
	assign x_1842 = ((~v_25 | v_23) | v_396) ;
	assign x_1841 = ((~v_23 | ~v_29) | v_397) ;
	assign x_4251 = (x_1839 & x_1840) ;
	assign x_1838 = ((~v_38 | v_24) | v_400) ;
	assign x_1837 = ((~v_24 | ~v_41) | v_401) ;
	assign x_1836 = ((~v_19 | ~v_43) | v_402) ;
	assign x_1835 = ((~v_39 | v_20) | v_403) ;
	assign x_1834 = (v_404 | ~v_35) ;
	assign x_1833 = (v_404 | ~v_36) ;
	assign x_1832 = (v_404 | ~v_70) ;
	assign x_4242 = (x_1830 & x_1831) ;
	assign x_1829 = (v_404 | ~v_82) ;
	assign x_1828 = (v_404 | ~v_88) ;
	assign x_1827 = (v_404 | ~v_403) ;
	assign x_1826 = (v_404 | ~v_402) ;
	assign x_1825 = (v_404 | ~v_401) ;
	assign x_1824 = (v_404 | ~v_400) ;
	assign x_1823 = (v_404 | ~v_399) ;
	assign x_4234 = (x_1821 & x_1822) ;
	assign x_1820 = (v_404 | ~v_396) ;
	assign x_1819 = ((~v_26 | v_23) | v_405) ;
	assign x_1818 = ((v_20 | ~v_52) | v_406) ;
	assign x_1817 = ((~v_23 | ~v_28) | v_407) ;
	assign x_1816 = ((~v_20 | ~v_55) | v_408) ;
	assign x_1815 = ((v_19 | ~v_53) | v_409) ;
	assign x_1814 = ((v_24 | ~v_51) | v_410) ;
	assign x_4220 = (x_1812 & x_1813) ;
	assign x_1811 = (v_413 | ~v_48) ;
	assign x_1810 = (v_413 | ~v_49) ;
	assign x_1809 = (v_413 | ~v_73) ;
	assign x_4216 = (x_1807 & x_1808) ;
	assign x_1806 = (v_413 | ~v_83) ;
	assign x_1805 = (v_413 | ~v_89) ;
	assign x_1804 = (v_413 | ~v_412) ;
	assign x_4211 = (x_1802 & x_1803) ;
	assign x_1801 = (v_413 | ~v_409) ;
	assign x_1800 = (v_413 | ~v_408) ;
	assign x_1799 = (v_413 | ~v_407) ;
	assign x_1798 = (v_413 | ~v_406) ;
	assign x_1797 = (v_413 | ~v_405) ;
	assign x_1796 = ((~v_27 | v_23) | v_414) ;
	assign x_1795 = ((v_20 | ~v_65) | v_415) ;
	assign x_4202 = (x_1793 & x_1794) ;
	assign x_1792 = ((v_24 | ~v_64) | v_418) ;
	assign x_1791 = ((v_19 | ~v_66) | v_419) ;
	assign x_1790 = ((~v_24 | ~v_67) | v_420) ;
	assign x_4198 = (x_1788 & x_1789) ;
	assign x_1787 = (v_422 | ~v_62) ;
	assign x_1786 = (v_422 | ~v_76) ;
	assign x_1785 = (v_422 | ~v_77) ;
	assign x_4193 = (x_1783 & x_1784) ;
	assign x_1782 = (v_422 | ~v_421) ;
	assign x_1781 = (v_422 | ~v_420) ;
	assign x_1780 = (v_422 | ~v_90) ;
	assign x_1779 = (v_422 | ~v_419) ;
	assign x_1778 = (v_422 | ~v_418) ;
	assign x_1777 = (v_422 | ~v_417) ;
	assign x_1776 = (v_422 | ~v_416) ;
	assign x_4183 = (x_1774 & x_1775) ;
	assign x_1773 = (((~v_422 | ~v_413) | ~v_404) | v_423) ;
	assign x_1772 = ((~v_38 | v_19) | v_424) ;
	assign x_1771 = ((~v_25 | v_17) | v_425) ;
	assign x_4179 = (x_1769 & x_1770) ;
	assign x_1768 = ((~v_9 | ~v_43) | v_428) ;
	assign x_1767 = ((~v_39 | v_11) | v_429) ;
	assign x_1766 = ((~v_19 | ~v_41) | v_430) ;
	assign x_4174 = (x_1764 & x_1765) ;
	assign x_1763 = (v_432 | ~v_34) ;
	assign x_1762 = (v_432 | ~v_35) ;
	assign x_1761 = (v_432 | ~v_36) ;
	assign x_1760 = (v_432 | ~v_37) ;
	assign x_1759 = (v_432 | ~v_70) ;
	assign x_1758 = (v_432 | ~v_79) ;
	assign x_1757 = (v_432 | ~v_431) ;
	assign x_4165 = (x_1755 & x_1756) ;
	assign x_1754 = (v_432 | ~v_428) ;
	assign x_1753 = (v_432 | ~v_427) ;
	assign x_1752 = (v_432 | ~v_426) ;
	assign x_4161 = (x_1750 & x_1751) ;
	assign x_1749 = ((v_19 | ~v_51) | v_433) ;
	assign x_1748 = ((~v_19 | ~v_54) | v_434) ;
	assign x_1747 = ((~v_26 | v_17) | v_435) ;
	assign x_4156 = (x_1745 & x_1746) ;
	assign x_1744 = ((~v_17 | ~v_28) | v_438) ;
	assign x_1743 = ((~v_11 | ~v_55) | v_439) ;
	assign x_1742 = ((~v_9 | ~v_56) | v_440) ;
	assign x_1741 = (v_441 | ~v_46) ;
	assign x_1740 = (v_441 | ~v_47) ;
	assign x_1739 = (v_441 | ~v_48) ;
	assign x_1738 = (v_441 | ~v_49) ;
	assign x_4145 = (x_1736 & x_1737) ;
	assign x_1735 = (v_441 | ~v_80) ;
	assign x_1734 = (v_441 | ~v_440) ;
	assign x_1733 = (v_441 | ~v_439) ;
	assign x_4141 = (x_1731 & x_1732) ;
	assign x_1730 = (v_441 | ~v_436) ;
	assign x_1729 = (v_441 | ~v_435) ;
	assign x_1728 = (v_441 | ~v_434) ;
	assign x_4136 = (x_1726 & x_1727) ;
	assign x_1725 = ((v_11 | ~v_65) | v_443) ;
	assign x_1724 = ((v_9 | ~v_66) | v_444) ;
	assign x_1723 = ((~v_9 | ~v_69) | v_445) ;
	assign x_1722 = ((v_19 | ~v_64) | v_446) ;
	assign x_1721 = ((~v_27 | v_17) | v_447) ;
	assign x_1720 = ((~v_11 | ~v_68) | v_448) ;
	assign x_1719 = ((~v_17 | ~v_30) | v_449) ;
	assign x_4127 = (x_1717 & x_1718) ;
	assign x_1716 = (v_450 | ~v_61) ;
	assign x_1715 = (v_450 | ~v_62) ;
	assign x_1714 = (v_450 | ~v_63) ;
	assign x_4123 = (x_1712 & x_1713) ;
	assign x_1711 = (v_450 | ~v_449) ;
	assign x_1710 = (v_450 | ~v_448) ;
	assign x_1709 = (v_450 | ~v_447) ;
	assign x_4118 = (x_1707 & x_1708) ;
	assign x_1706 = (v_450 | ~v_444) ;
	assign x_1705 = (v_450 | ~v_443) ;
	assign x_1704 = (v_450 | ~v_442) ;
	assign x_1703 = (((~v_450 | ~v_441) | ~v_432) | v_451) ;
	assign x_1702 = ((~v_28 | v_30) | v_452) ;
	assign x_1701 = ((~v_26 | v_25) | v_453) ;
	assign x_1700 = ((~v_29 | v_28) | v_454) ;
	assign x_4108 = (x_1698 & x_1699) ;
	assign x_1697 = (v_456 | ~v_454) ;
	assign x_1696 = (v_456 | ~v_453) ;
	assign x_1695 = (v_456 | ~v_452) ;
	assign x_4104 = (x_1693 & x_1694) ;
	assign x_1692 = ((~v_26 | v_22) | v_457) ;
	assign x_1691 = ((v_16 | ~v_52) | v_458) ;
	assign x_1690 = ((~v_16 | ~v_55) | v_459) ;
	assign x_4099 = (x_1688 & x_1689) ;
	assign x_1687 = ((~v_22 | ~v_28) | v_462) ;
	assign x_1686 = (v_463 | ~v_48) ;
	assign x_1685 = (v_463 | ~v_49) ;
	assign x_1684 = (v_463 | ~v_50) ;
	assign x_1683 = (v_463 | ~v_73) ;
	assign x_1682 = (v_463 | ~v_74) ;
	assign x_1681 = (v_463 | ~v_80) ;
	assign x_4090 = (x_1679 & x_1680) ;
	assign x_1678 = (v_463 | ~v_461) ;
	assign x_1677 = (v_463 | ~v_460) ;
	assign x_1676 = (v_463 | ~v_411) ;
	assign x_1675 = (v_463 | ~v_410) ;
	assign x_1674 = (v_463 | ~v_459) ;
	assign x_1673 = (v_463 | ~v_458) ;
	assign x_1672 = (v_463 | ~v_457) ;
	assign x_4082 = (x_1670 & x_1671) ;
	assign x_1669 = ((~v_16 | ~v_68) | v_466) ;
	assign x_1668 = ((~v_14 | ~v_69) | v_467) ;
	assign x_1667 = ((v_14 | ~v_66) | v_468) ;
	assign x_1666 = ((~v_22 | ~v_30) | v_469) ;
	assign x_1665 = (v_470 | ~v_61) ;
	assign x_1664 = (v_470 | ~v_62) ;
	assign x_1663 = (v_470 | ~v_63) ;
	assign x_4070 = (x_1661 & x_1662) ;
	assign x_1660 = (v_470 | ~v_81) ;
	assign x_1659 = (v_470 | ~v_469) ;
	assign x_1658 = (v_470 | ~v_420) ;
	assign x_4066 = (x_1656 & x_1657) ;
	assign x_1655 = (v_470 | ~v_467) ;
	assign x_1654 = (v_470 | ~v_418) ;
	assign x_1653 = (v_470 | ~v_466) ;
	assign x_4061 = (x_1651 & x_1652) ;
	assign x_1650 = ((~v_22 | ~v_29) | v_471) ;
	assign x_1649 = ((v_14 | ~v_40) | v_472) ;
	assign x_1648 = ((~v_16 | ~v_42) | v_473) ;
	assign x_1647 = ((~v_39 | v_16) | v_474) ;
	assign x_1646 = ((~v_25 | v_22) | v_475) ;
	assign x_1645 = ((~v_14 | ~v_43) | v_476) ;
	assign x_1644 = (v_477 | ~v_35) ;
	assign x_4052 = (x_1642 & x_1643) ;
	assign x_1641 = (v_477 | ~v_70) ;
	assign x_1640 = (v_477 | ~v_71) ;
	assign x_1639 = (v_477 | ~v_79) ;
	assign x_4048 = (x_1637 & x_1638) ;
	assign x_1636 = (v_477 | ~v_475) ;
	assign x_1635 = (v_477 | ~v_474) ;
	assign x_1634 = (v_477 | ~v_473) ;
	assign x_4043 = (x_1632 & x_1633) ;
	assign x_1631 = (v_477 | ~v_400) ;
	assign x_1630 = (v_477 | ~v_471) ;
	assign x_1629 = (((~v_477 | ~v_470) | ~v_463) | v_478) ;
	assign x_1628 = ((~v_38 | v_14) | v_479) ;
	assign x_1627 = ((~v_25 | v_13) | v_480) ;
	assign x_1626 = ((~v_39 | v_10) | v_481) ;
	assign x_1625 = ((~v_14 | ~v_41) | v_482) ;
	assign x_4033 = (x_1623 & x_1624) ;
	assign x_1622 = (v_485 | ~v_33) ;
	assign x_1621 = (v_485 | ~v_34) ;
	assign x_1620 = (v_485 | ~v_35) ;
	assign x_4029 = (x_1618 & x_1619) ;
	assign x_1617 = (v_485 | ~v_79) ;
	assign x_1616 = (v_485 | ~v_82) ;
	assign x_1615 = (v_485 | ~v_484) ;
	assign x_4024 = (x_1613 & x_1614) ;
	assign x_1612 = (v_485 | ~v_481) ;
	assign x_1611 = (v_485 | ~v_480) ;
	assign x_1610 = (v_485 | ~v_479) ;
	assign x_1609 = (v_485 | ~v_428) ;
	assign x_1608 = (v_485 | ~v_427) ;
	assign x_1607 = ((v_14 | ~v_51) | v_486) ;
	assign x_1606 = ((~v_26 | v_13) | v_487) ;
	assign x_4015 = (x_1604 & x_1605) ;
	assign x_1603 = ((~v_13 | ~v_28) | v_490) ;
	assign x_1602 = ((~v_10 | ~v_55) | v_491) ;
	assign x_1601 = (v_492 | ~v_46) ;
	assign x_4011 = (x_1599 & x_1600) ;
	assign x_1598 = (v_492 | ~v_49) ;
	assign x_1597 = (v_492 | ~v_73) ;
	assign x_1596 = (v_492 | ~v_80) ;
	assign x_4006 = (x_1594 & x_1595) ;
	assign x_1593 = (v_492 | ~v_491) ;
	assign x_1592 = (v_492 | ~v_490) ;
	assign x_1591 = (v_492 | ~v_489) ;
	assign x_1590 = (v_492 | ~v_488) ;
	assign x_1589 = (v_492 | ~v_487) ;
	assign x_1588 = (v_492 | ~v_486) ;
	assign x_1587 = (v_492 | ~v_437) ;
	assign x_3995 = (x_1585 & x_1586) ;
	assign x_1584 = ((v_10 | ~v_65) | v_495) ;
	assign x_1583 = ((~v_13 | ~v_30) | v_496) ;
	assign x_1582 = ((~v_14 | ~v_67) | v_497) ;
	assign x_3991 = (x_1580 & x_1581) ;
	assign x_1579 = (v_499 | ~v_60) ;
	assign x_1578 = (v_499 | ~v_61) ;
	assign x_1577 = (v_499 | ~v_62) ;
	assign x_3986 = (x_1575 & x_1576) ;
	assign x_1574 = (v_499 | ~v_84) ;
	assign x_1573 = (v_499 | ~v_498) ;
	assign x_1572 = (v_499 | ~v_497) ;
	assign x_1571 = (v_499 | ~v_496) ;
	assign x_1570 = (v_499 | ~v_495) ;
	assign x_1569 = (v_499 | ~v_494) ;
	assign x_1568 = (v_499 | ~v_493) ;
	assign x_3977 = (x_1566 & x_1567) ;
	assign x_1565 = (((~v_499 | ~v_492) | ~v_485) | v_500) ;
	assign x_1564 = (v_501 | ~v_455) ;
	assign x_1563 = (v_501 | ~v_454) ;
	assign x_3973 = (x_1561 & x_1562) ;
	assign x_1560 = (v_501 | ~v_500) ;
	assign x_1559 = (v_501 | ~v_478) ;
	assign x_1558 = ((~v_25 | v_21) | v_502) ;
	assign x_3968 = (x_1556 & x_1557) ;
	assign x_1555 = ((~v_39 | v_12) | v_505) ;
	assign x_1554 = (v_506 | ~v_33) ;
	assign x_1553 = (v_506 | ~v_35) ;
	assign x_1552 = (v_506 | ~v_36) ;
	assign x_1551 = (v_506 | ~v_37) ;
	assign x_1550 = (v_506 | ~v_70) ;
	assign x_1549 = (v_506 | ~v_79) ;
	assign x_3958 = (x_1547 & x_1548) ;
	assign x_1546 = (v_506 | ~v_504) ;
	assign x_1545 = (v_506 | ~v_428) ;
	assign x_1544 = (v_506 | ~v_427) ;
	assign x_3954 = (x_1542 & x_1543) ;
	assign x_1541 = (v_506 | ~v_401) ;
	assign x_1540 = (v_506 | ~v_400) ;
	assign x_1539 = ((~v_26 | v_21) | v_507) ;
	assign x_3949 = (x_1537 & x_1538) ;
	assign x_1536 = ((~v_12 | ~v_55) | v_510) ;
	assign x_1535 = (v_511 | ~v_46) ;
	assign x_1534 = (v_511 | ~v_48) ;
	assign x_1533 = (v_511 | ~v_49) ;
	assign x_1532 = (v_511 | ~v_50) ;
	assign x_1531 = (v_511 | ~v_73) ;
	assign x_1530 = (v_511 | ~v_80) ;
	assign x_3940 = (x_1528 & x_1529) ;
	assign x_1527 = (v_511 | ~v_510) ;
	assign x_1526 = (v_511 | ~v_437) ;
	assign x_1525 = (v_511 | ~v_509) ;
	assign x_1524 = (v_511 | ~v_508) ;
	assign x_1523 = (v_511 | ~v_507) ;
	assign x_1522 = (v_511 | ~v_411) ;
	assign x_1521 = (v_511 | ~v_410) ;
	assign x_3932 = (x_1519 & x_1520) ;
	assign x_1518 = ((v_12 | ~v_65) | v_514) ;
	assign x_1517 = ((~v_12 | ~v_68) | v_515) ;
	assign x_1516 = (v_516 | ~v_59) ;
	assign x_1515 = (v_516 | ~v_61) ;
	assign x_1514 = (v_516 | ~v_62) ;
	assign x_1513 = (v_516 | ~v_63) ;
	assign x_1512 = (v_516 | ~v_76) ;
	assign x_3919 = (x_1510 & x_1511) ;
	assign x_1509 = (v_516 | ~v_420) ;
	assign x_1508 = (v_516 | ~v_90) ;
	assign x_1507 = (v_516 | ~v_514) ;
	assign x_3915 = (x_1505 & x_1506) ;
	assign x_1504 = (v_516 | ~v_513) ;
	assign x_1503 = (v_516 | ~v_512) ;
	assign x_1502 = (v_516 | ~v_418) ;
	assign x_3910 = (x_1500 & x_1501) ;
	assign x_1499 = (v_518 | ~v_454) ;
	assign x_1498 = (v_518 | ~v_453) ;
	assign x_1497 = (v_518 | ~v_452) ;
	assign x_1496 = (v_518 | ~v_517) ;
	assign x_1495 = (((~v_518 | ~v_501) | ~v_456) | v_519) ;
	assign x_1494 = ((~v_26 | v_16) | v_520) ;
	assign x_1493 = ((v_22 | ~v_52) | v_521) ;
	assign x_3901 = (x_1491 & x_1492) ;
	assign x_1490 = ((~v_16 | ~v_28) | v_524) ;
	assign x_1489 = ((~v_24 | ~v_56) | v_525) ;
	assign x_1488 = (v_526 | ~v_47) ;
	assign x_3897 = (x_1486 & x_1487) ;
	assign x_1485 = (v_526 | ~v_73) ;
	assign x_1484 = (v_526 | ~v_74) ;
	assign x_1483 = (v_526 | ~v_80) ;
	assign x_3892 = (x_1481 & x_1482) ;
	assign x_1480 = (v_526 | ~v_524) ;
	assign x_1479 = (v_526 | ~v_523) ;
	assign x_1478 = (v_526 | ~v_489) ;
	assign x_1477 = (v_526 | ~v_486) ;
	assign x_1476 = (v_526 | ~v_522) ;
	assign x_1475 = (v_526 | ~v_521) ;
	assign x_1474 = (v_526 | ~v_520) ;
	assign x_3882 = (x_1472 & x_1473) ;
	assign x_1471 = ((v_24 | ~v_66) | v_529) ;
	assign x_1470 = ((~v_24 | ~v_69) | v_530) ;
	assign x_1469 = ((~v_27 | v_16) | v_531) ;
	assign x_3878 = (x_1467 & x_1468) ;
	assign x_1466 = (v_533 | ~v_62) ;
	assign x_1465 = (v_533 | ~v_63) ;
	assign x_1464 = (v_533 | ~v_76) ;
	assign x_3873 = (x_1462 & x_1463) ;
	assign x_1461 = (v_533 | ~v_532) ;
	assign x_1460 = (v_533 | ~v_87) ;
	assign x_1459 = (v_533 | ~v_497) ;
	assign x_1458 = (v_533 | ~v_531) ;
	assign x_1457 = (v_533 | ~v_493) ;
	assign x_1456 = (v_533 | ~v_530) ;
	assign x_1455 = (v_533 | ~v_529) ;
	assign x_3864 = (x_1453 & x_1454) ;
	assign x_1452 = ((~v_25 | v_16) | v_534) ;
	assign x_1451 = ((~v_39 | v_22) | v_535) ;
	assign x_1450 = ((~v_16 | ~v_29) | v_536) ;
	assign x_3860 = (x_1448 & x_1449) ;
	assign x_1447 = ((~v_24 | ~v_43) | v_539) ;
	assign x_1446 = (v_540 | ~v_34) ;
	assign x_1445 = (v_540 | ~v_36) ;
	assign x_3855 = (x_1443 & x_1444) ;
	assign x_1442 = (v_540 | ~v_71) ;
	assign x_1441 = (v_540 | ~v_79) ;
	assign x_1440 = (v_540 | ~v_85) ;
	assign x_1439 = (v_540 | ~v_539) ;
	assign x_1438 = (v_540 | ~v_538) ;
	assign x_1437 = (v_540 | ~v_482) ;
	assign x_1436 = (v_540 | ~v_479) ;
	assign x_3844 = (x_1434 & x_1435) ;
	assign x_1433 = (v_540 | ~v_535) ;
	assign x_1432 = (v_540 | ~v_534) ;
	assign x_1431 = (((~v_540 | ~v_533) | ~v_526) | v_541) ;
	assign x_3840 = (x_1429 & x_1430) ;
	assign x_1428 = (v_542 | ~v_453) ;
	assign x_1427 = (v_542 | ~v_452) ;
	assign x_1426 = (v_542 | ~v_541) ;
	assign x_3835 = (x_1424 & x_1425) ;
	assign x_1423 = ((~v_20 | ~v_29) | v_544) ;
	assign x_1422 = ((~v_23 | ~v_42) | v_545) ;
	assign x_1421 = ((~v_25 | v_20) | v_546) ;
	assign x_1420 = (v_547 | ~v_34) ;
	assign x_1419 = (v_547 | ~v_37) ;
	assign x_1418 = (v_547 | ~v_70) ;
	assign x_1417 = (v_547 | ~v_71) ;
	assign x_3826 = (x_1415 & x_1416) ;
	assign x_1414 = (v_547 | ~v_85) ;
	assign x_1413 = (v_547 | ~v_546) ;
	assign x_1412 = (v_547 | ~v_430) ;
	assign x_3822 = (x_1410 & x_1411) ;
	assign x_1409 = (v_547 | ~v_424) ;
	assign x_1408 = (v_547 | ~v_545) ;
	assign x_1407 = (v_547 | ~v_544) ;
	assign x_3817 = (x_1405 & x_1406) ;
	assign x_1404 = ((v_23 | ~v_52) | v_549) ;
	assign x_1403 = ((~v_23 | ~v_55) | v_550) ;
	assign x_1402 = ((~v_20 | ~v_28) | v_551) ;
	assign x_1401 = (v_552 | ~v_551) ;
	assign x_1400 = (v_552 | ~v_47) ;
	assign x_1399 = (v_552 | ~v_50) ;
	assign x_1398 = (v_552 | ~v_73) ;
	assign x_3807 = (x_1396 & x_1397) ;
	assign x_1395 = (v_552 | ~v_80) ;
	assign x_1394 = (v_552 | ~v_86) ;
	assign x_1393 = (v_552 | ~v_525) ;
	assign x_3803 = (x_1391 & x_1392) ;
	assign x_1390 = (v_552 | ~v_434) ;
	assign x_1389 = (v_552 | ~v_433) ;
	assign x_1388 = (v_552 | ~v_549) ;
	assign x_3798 = (x_1386 & x_1387) ;
	assign x_1385 = ((v_23 | ~v_65) | v_554) ;
	assign x_1384 = ((~v_23 | ~v_68) | v_555) ;
	assign x_1383 = ((~v_20 | ~v_30) | v_556) ;
	assign x_1382 = (v_557 | ~v_556) ;
	assign x_1381 = (v_557 | ~v_60) ;
	assign x_1380 = (v_557 | ~v_63) ;
	assign x_1379 = (v_557 | ~v_76) ;
	assign x_3789 = (x_1377 & x_1378) ;
	assign x_1376 = (v_557 | ~v_81) ;
	assign x_1375 = (v_557 | ~v_555) ;
	assign x_1374 = (v_557 | ~v_87) ;
	assign x_1373 = (v_557 | ~v_446) ;
	assign x_1372 = (v_557 | ~v_530) ;
	assign x_1371 = (v_557 | ~v_529) ;
	assign x_1370 = (v_557 | ~v_442) ;
	assign x_3781 = (x_1368 & x_1369) ;
	assign x_1367 = (((~v_557 | ~v_552) | ~v_547) | v_558) ;
	assign x_1366 = (v_559 | ~v_455) ;
	assign x_1365 = (v_559 | ~v_454) ;
	assign x_1364 = (v_559 | ~v_453) ;
	assign x_1363 = (v_559 | ~v_452) ;
	assign x_1362 = (v_559 | ~v_517) ;
	assign x_1361 = (v_559 | ~v_558) ;
	assign x_3769 = (x_1359 & x_1360) ;
	assign x_1358 = ((~v_18 | ~v_29) | v_562) ;
	assign x_1357 = ((~v_25 | v_18) | v_563) ;
	assign x_1356 = (v_564 | ~v_34) ;
	assign x_3765 = (x_1354 & x_1355) ;
	assign x_1353 = (v_564 | ~v_70) ;
	assign x_1352 = (v_564 | ~v_71) ;
	assign x_1351 = (v_564 | ~v_79) ;
	assign x_3760 = (x_1349 & x_1350) ;
	assign x_1348 = (v_564 | ~v_430) ;
	assign x_1347 = (v_564 | ~v_476) ;
	assign x_1346 = (v_564 | ~v_562) ;
	assign x_1345 = (v_564 | ~v_472) ;
	assign x_1344 = (v_564 | ~v_424) ;
	assign x_1343 = (v_564 | ~v_561) ;
	assign x_1342 = (v_564 | ~v_560) ;
	assign x_3751 = (x_1340 & x_1341) ;
	assign x_1339 = ((~v_15 | ~v_55) | v_567) ;
	assign x_1338 = ((~v_18 | ~v_28) | v_568) ;
	assign x_1337 = (v_569 | ~v_47) ;
	assign x_3747 = (x_1335 & x_1336) ;
	assign x_1334 = (v_569 | ~v_73) ;
	assign x_1333 = (v_569 | ~v_74) ;
	assign x_1332 = (v_569 | ~v_80) ;
	assign x_3742 = (x_1330 & x_1331) ;
	assign x_1329 = (v_569 | ~v_461) ;
	assign x_1328 = (v_569 | ~v_460) ;
	assign x_1327 = (v_569 | ~v_434) ;
	assign x_1326 = (v_569 | ~v_433) ;
	assign x_1325 = (v_569 | ~v_567) ;
	assign x_1324 = (v_569 | ~v_566) ;
	assign x_1323 = (v_569 | ~v_565) ;
	assign x_3732 = (x_1321 & x_1322) ;
	assign x_1320 = ((~v_18 | ~v_30) | v_572) ;
	assign x_1319 = ((~v_15 | ~v_68) | v_573) ;
	assign x_1318 = (v_574 | ~v_60) ;
	assign x_3728 = (x_1316 & x_1317) ;
	assign x_1315 = (v_574 | ~v_76) ;
	assign x_1314 = (v_574 | ~v_77) ;
	assign x_1313 = (v_574 | ~v_81) ;
	assign x_3723 = (x_1311 & x_1312) ;
	assign x_1310 = (v_574 | ~v_468) ;
	assign x_1309 = (v_574 | ~v_467) ;
	assign x_1308 = (v_574 | ~v_442) ;
	assign x_1307 = (v_574 | ~v_573) ;
	assign x_1306 = (v_574 | ~v_572) ;
	assign x_1305 = (v_574 | ~v_571) ;
	assign x_1304 = (v_574 | ~v_570) ;
	assign x_3714 = (x_1302 & x_1303) ;
	assign x_1301 = (v_576 | ~v_454) ;
	assign x_1300 = (v_576 | ~v_453) ;
	assign x_1299 = (v_576 | ~v_452) ;
	assign x_3710 = (x_1297 & x_1298) ;
	assign x_1296 = (v_577 | ~v_455) ;
	assign x_1295 = (v_577 | ~v_454) ;
	assign x_1294 = (v_577 | ~v_453) ;
	assign x_3705 = (x_1292 & x_1293) ;
	assign x_1291 = (((~v_577 | ~v_576) | ~v_559) | v_578) ;
	assign x_1290 = ((~v_39 | v_18) | v_579) ;
	assign x_1289 = ((~v_15 | ~v_29) | v_580) ;
	assign x_1288 = ((~v_18 | ~v_42) | v_581) ;
	assign x_1287 = ((~v_25 | v_15) | v_582) ;
	assign x_1286 = (v_583 | ~v_34) ;
	assign x_1285 = (v_583 | ~v_35) ;
	assign x_3694 = (x_1283 & x_1284) ;
	assign x_1282 = (v_583 | ~v_71) ;
	assign x_1281 = (v_583 | ~v_72) ;
	assign x_1280 = (v_583 | ~v_79) ;
	assign x_3690 = (x_1278 & x_1279) ;
	assign x_1277 = (v_583 | ~v_482) ;
	assign x_1276 = (v_583 | ~v_479) ;
	assign x_1275 = (v_583 | ~v_399) ;
	assign x_3685 = (x_1273 & x_1274) ;
	assign x_1272 = (v_583 | ~v_579) ;
	assign x_1271 = ((~v_26 | v_15) | v_584) ;
	assign x_1270 = ((v_18 | ~v_52) | v_585) ;
	assign x_1269 = ((~v_18 | ~v_55) | v_586) ;
	assign x_1268 = ((~v_15 | ~v_28) | v_587) ;
	assign x_1267 = (v_588 | ~v_587) ;
	assign x_1266 = (v_588 | ~v_47) ;
	assign x_3676 = (x_1264 & x_1265) ;
	assign x_1263 = (v_588 | ~v_73) ;
	assign x_1262 = (v_588 | ~v_74) ;
	assign x_1261 = (v_588 | ~v_75) ;
	assign x_3672 = (x_1259 & x_1260) ;
	assign x_1258 = (v_588 | ~v_489) ;
	assign x_1257 = (v_588 | ~v_486) ;
	assign x_1256 = (v_588 | ~v_409) ;
	assign x_3667 = (x_1254 & x_1255) ;
	assign x_1253 = (v_588 | ~v_584) ;
	assign x_1252 = ((~v_27 | v_15) | v_589) ;
	assign x_1251 = ((v_18 | ~v_65) | v_590) ;
	assign x_1250 = ((~v_18 | ~v_68) | v_591) ;
	assign x_1249 = ((~v_15 | ~v_30) | v_592) ;
	assign x_1248 = (v_593 | ~v_592) ;
	assign x_1247 = (v_593 | ~v_60) ;
	assign x_3657 = (x_1245 & x_1246) ;
	assign x_1244 = (v_593 | ~v_76) ;
	assign x_1243 = (v_593 | ~v_77) ;
	assign x_1242 = (v_593 | ~v_78) ;
	assign x_3653 = (x_1240 & x_1241) ;
	assign x_1239 = (v_593 | ~v_419) ;
	assign x_1238 = (v_593 | ~v_497) ;
	assign x_1237 = (v_593 | ~v_493) ;
	assign x_3648 = (x_1235 & x_1236) ;
	assign x_1234 = (v_593 | ~v_589) ;
	assign x_1233 = (((~v_593 | ~v_588) | ~v_583) | v_594) ;
	assign x_1232 = (v_595 | ~v_455) ;
	assign x_1231 = (v_595 | ~v_454) ;
	assign x_1230 = (v_595 | ~v_453) ;
	assign x_1229 = (v_595 | ~v_452) ;
	assign x_1228 = (v_595 | ~v_594) ;
	assign x_3639 = (x_1226 & x_1227) ;
	assign x_1225 = (v_596 | ~v_454) ;
	assign x_1224 = (v_596 | ~v_453) ;
	assign x_1223 = (v_596 | ~v_452) ;
	assign x_1222 = (v_596 | ~v_517) ;
	assign x_1221 = (v_596 | ~v_541) ;
	assign x_1220 = (v_597 | ~v_455) ;
	assign x_1219 = (v_597 | ~v_454) ;
	assign x_3631 = (x_1217 & x_1218) ;
	assign x_1216 = (v_597 | ~v_594) ;
	assign x_1215 = (v_597 | ~v_451) ;
	assign x_1214 = (v_598 | ~v_455) ;
	assign x_1213 = (v_598 | ~v_454) ;
	assign x_1212 = (v_598 | ~v_453) ;
	assign x_1211 = (v_598 | ~v_452) ;
	assign x_1210 = (v_598 | ~v_500) ;
	assign x_3616 = (x_1208 & x_1209) ;
	assign x_1207 = ((~v_39 | v_21) | v_601) ;
	assign x_1206 = ((~v_21 | ~v_42) | v_602) ;
	assign x_1205 = ((~v_38 | v_9) | v_603) ;
	assign x_3612 = (x_1203 & x_1204) ;
	assign x_1202 = (v_606 | ~v_32) ;
	assign x_1201 = (v_606 | ~v_34) ;
	assign x_1200 = (v_606 | ~v_36) ;
	assign x_3607 = (x_1198 & x_1199) ;
	assign x_1197 = (v_606 | ~v_71) ;
	assign x_1196 = (v_606 | ~v_85) ;
	assign x_1195 = (v_606 | ~v_605) ;
	assign x_1194 = (v_606 | ~v_604) ;
	assign x_1193 = (v_606 | ~v_539) ;
	assign x_1192 = (v_606 | ~v_603) ;
	assign x_1191 = (v_606 | ~v_602) ;
	assign x_3598 = (x_1189 & x_1190) ;
	assign x_1188 = (v_606 | ~v_537) ;
	assign x_1187 = ((v_21 | ~v_52) | v_607) ;
	assign x_1186 = ((v_9 | ~v_51) | v_608) ;
	assign x_3594 = (x_1184 & x_1185) ;
	assign x_1183 = ((~v_12 | ~v_28) | v_611) ;
	assign x_1182 = ((~v_9 | ~v_54) | v_612) ;
	assign x_1181 = (v_613 | ~v_45) ;
	assign x_3589 = (x_1179 & x_1180) ;
	assign x_1178 = (v_613 | ~v_50) ;
	assign x_1177 = (v_613 | ~v_73) ;
	assign x_1176 = (v_613 | ~v_74) ;
	assign x_1175 = (v_613 | ~v_86) ;
	assign x_1174 = (v_613 | ~v_612) ;
	assign x_1173 = (v_613 | ~v_525) ;
	assign x_1172 = (v_613 | ~v_611) ;
	assign x_3579 = (x_1170 & x_1171) ;
	assign x_1169 = (v_613 | ~v_608) ;
	assign x_1168 = (v_613 | ~v_607) ;
	assign x_1167 = (v_613 | ~v_522) ;
	assign x_3575 = (x_1165 & x_1166) ;
	assign x_1164 = ((v_9 | ~v_64) | v_616) ;
	assign x_1163 = ((~v_21 | ~v_68) | v_617) ;
	assign x_1162 = ((~v_9 | ~v_67) | v_618) ;
	assign x_3570 = (x_1160 & x_1161) ;
	assign x_1159 = (v_620 | ~v_60) ;
	assign x_1158 = (v_620 | ~v_62) ;
	assign x_1157 = (v_620 | ~v_63) ;
	assign x_1156 = (v_620 | ~v_76) ;
	assign x_1155 = (v_620 | ~v_77) ;
	assign x_1154 = (v_620 | ~v_619) ;
	assign x_1153 = (v_620 | ~v_87) ;
	assign x_3561 = (x_1151 & x_1152) ;
	assign x_1150 = (v_620 | ~v_616) ;
	assign x_1149 = (v_620 | ~v_615) ;
	assign x_1148 = (v_620 | ~v_614) ;
	assign x_3557 = (x_1146 & x_1147) ;
	assign x_1145 = (((~v_620 | ~v_613) | ~v_606) | v_621) ;
	assign x_1144 = (v_622 | ~v_455) ;
	assign x_1143 = (v_622 | ~v_454) ;
	assign x_3552 = (x_1141 & x_1142) ;
	assign x_1140 = (v_622 | ~v_423) ;
	assign x_1139 = (v_622 | ~v_621) ;
	assign x_1138 = ((~v_25 | v_10) | v_623) ;
	assign x_1137 = ((~v_39 | v_13) | v_624) ;
	assign x_1136 = ((~v_10 | ~v_29) | v_625) ;
	assign x_1135 = ((~v_13 | ~v_42) | v_626) ;
	assign x_1134 = (v_627 | ~v_32) ;
	assign x_3541 = (x_1132 & x_1133) ;
	assign x_1131 = (v_627 | ~v_37) ;
	assign x_1130 = (v_627 | ~v_70) ;
	assign x_1129 = (v_627 | ~v_71) ;
	assign x_3537 = (x_1127 & x_1128) ;
	assign x_1126 = (v_627 | ~v_476) ;
	assign x_1125 = (v_627 | ~v_626) ;
	assign x_1124 = (v_627 | ~v_625) ;
	assign x_3532 = (x_1122 & x_1123) ;
	assign x_1121 = (v_627 | ~v_623) ;
	assign x_1120 = (v_627 | ~v_603) ;
	assign x_1119 = ((v_13 | ~v_52) | v_628) ;
	assign x_1118 = ((~v_10 | ~v_28) | v_629) ;
	assign x_1117 = ((~v_13 | ~v_55) | v_630) ;
	assign x_1116 = ((~v_26 | v_10) | v_631) ;
	assign x_1115 = (v_632 | ~v_45) ;
	assign x_3523 = (x_1113 & x_1114) ;
	assign x_1112 = (v_632 | ~v_50) ;
	assign x_1111 = (v_632 | ~v_73) ;
	assign x_1110 = (v_632 | ~v_74) ;
	assign x_3519 = (x_1108 & x_1109) ;
	assign x_1107 = (v_632 | ~v_631) ;
	assign x_1106 = (v_632 | ~v_630) ;
	assign x_1105 = (v_632 | ~v_461) ;
	assign x_3514 = (x_1103 & x_1104) ;
	assign x_1102 = (v_632 | ~v_628) ;
	assign x_1101 = (v_632 | ~v_608) ;
	assign x_1100 = ((~v_27 | v_10) | v_633) ;
	assign x_1099 = ((v_13 | ~v_65) | v_634) ;
	assign x_1098 = ((~v_10 | ~v_30) | v_635) ;
	assign x_1097 = ((~v_13 | ~v_68) | v_636) ;
	assign x_1096 = (v_637 | ~v_58) ;
	assign x_3504 = (x_1094 & x_1095) ;
	assign x_1093 = (v_637 | ~v_63) ;
	assign x_1092 = (v_637 | ~v_76) ;
	assign x_1091 = (v_637 | ~v_77) ;
	assign x_3500 = (x_1089 & x_1090) ;
	assign x_1088 = (v_637 | ~v_636) ;
	assign x_1087 = (v_637 | ~v_635) ;
	assign x_1086 = (v_637 | ~v_468) ;
	assign x_3495 = (x_1084 & x_1085) ;
	assign x_1083 = (v_637 | ~v_616) ;
	assign x_1082 = (v_637 | ~v_467) ;
	assign x_1081 = (((~v_637 | ~v_632) | ~v_627) | v_638) ;
	assign x_1080 = (v_639 | ~v_455) ;
	assign x_1079 = (v_639 | ~v_454) ;
	assign x_1078 = (v_639 | ~v_453) ;
	assign x_1077 = (v_639 | ~v_452) ;
	assign x_3486 = (x_1075 & x_1076) ;
	assign x_1074 = (v_640 | ~v_455) ;
	assign x_1073 = (v_640 | ~v_454) ;
	assign x_1072 = (v_640 | ~v_453) ;
	assign x_3482 = (x_1070 & x_1071) ;
	assign x_1069 = (v_640 | ~v_478) ;
	assign x_1068 = ((~v_25 | v_11) | v_641) ;
	assign x_1067 = ((~v_39 | v_17) | v_642) ;
	assign x_3477 = (x_1065 & x_1066) ;
	assign x_1064 = (v_645 | ~v_32) ;
	assign x_1063 = (v_645 | ~v_34) ;
	assign x_1062 = (v_645 | ~v_35) ;
	assign x_1061 = (v_645 | ~v_36) ;
	assign x_1060 = (v_645 | ~v_37) ;
	assign x_1059 = (v_645 | ~v_70) ;
	assign x_1058 = (v_645 | ~v_71) ;
	assign x_3465 = (x_1056 & x_1057) ;
	assign x_1055 = (v_645 | ~v_402) ;
	assign x_1054 = (v_645 | ~v_603) ;
	assign x_1053 = (v_645 | ~v_643) ;
	assign x_3461 = (x_1051 & x_1052) ;
	assign x_1050 = (v_645 | ~v_399) ;
	assign x_1049 = ((v_17 | ~v_52) | v_646) ;
	assign x_1048 = ((~v_17 | ~v_55) | v_647) ;
	assign x_3456 = (x_1046 & x_1047) ;
	assign x_1045 = (v_650 | ~v_45) ;
	assign x_1044 = (v_650 | ~v_47) ;
	assign x_1043 = (v_650 | ~v_48) ;
	assign x_1042 = (v_650 | ~v_49) ;
	assign x_1041 = (v_650 | ~v_50) ;
	assign x_1040 = (v_650 | ~v_73) ;
	assign x_1039 = (v_650 | ~v_74) ;
	assign x_3447 = (x_1037 & x_1038) ;
	assign x_1036 = (v_650 | ~v_649) ;
	assign x_1035 = (v_650 | ~v_648) ;
	assign x_1034 = (v_650 | ~v_608) ;
	assign x_3443 = (x_1032 & x_1033) ;
	assign x_1031 = (v_650 | ~v_409) ;
	assign x_1030 = ((v_17 | ~v_65) | v_651) ;
	assign x_1029 = ((~v_17 | ~v_68) | v_652) ;
	assign x_3438 = (x_1027 & x_1028) ;
	assign x_1026 = (v_655 | ~v_58) ;
	assign x_1025 = (v_655 | ~v_60) ;
	assign x_1024 = (v_655 | ~v_61) ;
	assign x_1023 = (v_655 | ~v_62) ;
	assign x_1022 = (v_655 | ~v_63) ;
	assign x_1021 = (v_655 | ~v_76) ;
	assign x_1020 = (v_655 | ~v_77) ;
	assign x_3428 = (x_1018 & x_1019) ;
	assign x_1017 = (v_655 | ~v_421) ;
	assign x_1016 = (v_655 | ~v_618) ;
	assign x_1015 = (v_655 | ~v_419) ;
	assign x_3424 = (x_1013 & x_1014) ;
	assign x_1012 = (v_655 | ~v_651) ;
	assign x_1011 = (((~v_655 | ~v_650) | ~v_645) | v_656) ;
	assign x_1010 = (v_657 | ~v_455) ;
	assign x_3419 = (x_1008 & x_1009) ;
	assign x_1007 = (v_657 | ~v_452) ;
	assign x_1006 = (v_657 | ~v_517) ;
	assign x_1005 = (v_657 | ~v_656) ;
	assign x_1004 = (v_658 | ~v_455) ;
	assign x_1003 = (v_658 | ~v_454) ;
	assign x_1002 = (v_658 | ~v_453) ;
	assign x_1001 = (v_658 | ~v_452) ;
	assign x_3410 = (x_999 & x_1000) ;
	assign x_998 = (v_660 | ~v_455) ;
	assign x_997 = (v_660 | ~v_454) ;
	assign x_996 = (v_660 | ~v_453) ;
	assign x_3406 = (x_994 & x_995) ;
	assign x_993 = (v_660 | ~v_659) ;
	assign x_992 = (v_661 | ~v_455) ;
	assign x_991 = (v_661 | ~v_454) ;
	assign x_3401 = (x_989 & x_990) ;
	assign x_988 = (v_661 | ~v_541) ;
	assign x_987 = (v_661 | ~v_423) ;
	assign x_986 = (v_662 | ~v_455) ;
	assign x_985 = (v_662 | ~v_454) ;
	assign x_984 = (v_662 | ~v_453) ;
	assign x_983 = (v_662 | ~v_452) ;
	assign x_982 = (v_662 | ~v_500) ;
	assign x_3390 = (x_980 & x_981) ;
	assign x_979 = (v_663 | ~v_454) ;
	assign x_978 = (v_663 | ~v_453) ;
	assign x_977 = (v_663 | ~v_452) ;
	assign x_3386 = (x_975 & x_976) ;
	assign x_974 = (v_665 | ~v_455) ;
	assign x_973 = (v_665 | ~v_454) ;
	assign x_972 = (v_665 | ~v_453) ;
	assign x_3381 = (x_970 & x_971) ;
	assign x_969 = (v_665 | ~v_664) ;
	assign x_968 = (v_666 | ~v_455) ;
	assign x_967 = (v_666 | ~v_454) ;
	assign x_966 = (v_666 | ~v_453) ;
	assign x_965 = (v_666 | ~v_452) ;
	assign x_964 = (v_666 | ~v_656) ;
	assign x_963 = (((((~v_666 | ~v_665) | ~v_660) | ~v_639) | ~v_622) | v_667) ;
	assign x_3372 = (x_961 & x_962) ;
	assign x_960 = (((~v_666 | ~v_639) | ~v_622) | v_669) ;
	assign x_959 = (v_670 | ~v_455) ;
	assign x_958 = (v_670 | ~v_454) ;
	assign x_3368 = (x_956 & x_957) ;
	assign x_955 = (v_670 | ~v_517) ;
	assign x_954 = (v_670 | ~v_669) ;
	assign x_953 = (v_671 | ~v_455) ;
	assign x_3363 = (x_951 & x_952) ;
	assign x_950 = (v_671 | ~v_452) ;
	assign x_949 = (v_671 | ~v_478) ;
	assign x_948 = (v_671 | ~v_664) ;
	assign x_947 = (((((~v_658 | ~v_657) | ~v_640) | ~v_671) | ~v_670) | v_672) ;
	assign x_946 = (v_673 | ~v_455) ;
	assign x_945 = (v_673 | ~v_454) ;
	assign x_944 = (v_673 | ~v_453) ;
	assign x_3353 = (x_942 & x_943) ;
	assign x_941 = (v_673 | ~v_638) ;
	assign x_940 = (v_674 | ~v_455) ;
	assign x_939 = (v_674 | ~v_454) ;
	assign x_3349 = (x_937 & x_938) ;
	assign x_936 = (v_674 | ~v_558) ;
	assign x_935 = (v_674 | ~v_656) ;
	assign x_934 = (v_675 | ~v_455) ;
	assign x_3344 = (x_932 & x_933) ;
	assign x_931 = (v_675 | ~v_452) ;
	assign x_930 = (v_675 | ~v_621) ;
	assign x_929 = (((~v_675 | ~v_674) | ~v_673) | v_676) ;
	assign x_928 = (v_677 | ~v_455) ;
	assign x_927 = (v_677 | ~v_454) ;
	assign x_926 = (v_677 | ~v_453) ;
	assign x_925 = (v_677 | ~v_452) ;
	assign x_3335 = (x_923 & x_924) ;
	assign x_922 = (v_678 | ~v_455) ;
	assign x_921 = (v_678 | ~v_454) ;
	assign x_920 = (v_678 | ~v_453) ;
	assign x_919 = (v_678 | ~v_452) ;
	assign x_918 = (v_678 | ~v_541) ;
	assign x_917 = (v_678 | ~v_575) ;
	assign x_916 = (v_679 | ~v_455) ;
	assign x_3327 = (x_914 & x_915) ;
	assign x_913 = (v_679 | ~v_452) ;
	assign x_912 = (v_679 | ~v_451) ;
	assign x_911 = (v_679 | ~v_621) ;
	assign x_910 = (v_680 | ~v_455) ;
	assign x_909 = (v_680 | ~v_454) ;
	assign x_908 = (v_680 | ~v_453) ;
	assign x_907 = (v_680 | ~v_452) ;
	assign x_3314 = (x_905 & x_906) ;
	assign x_904 = (v_682 | ~v_455) ;
	assign x_903 = (v_682 | ~v_454) ;
	assign x_902 = (v_682 | ~v_453) ;
	assign x_3310 = (x_900 & x_901) ;
	assign x_899 = (v_682 | ~v_681) ;
	assign x_898 = (v_683 | ~v_455) ;
	assign x_897 = (v_683 | ~v_454) ;
	assign x_3305 = (x_895 & x_896) ;
	assign x_894 = (v_683 | ~v_594) ;
	assign x_893 = (v_683 | ~v_558) ;
	assign x_892 = (v_684 | ~v_455) ;
	assign x_891 = (v_684 | ~v_454) ;
	assign x_890 = (v_684 | ~v_453) ;
	assign x_889 = (v_684 | ~v_452) ;
	assign x_888 = (v_684 | ~v_500) ;
	assign x_3296 = (x_886 & x_887) ;
	assign x_885 = (v_685 | ~v_454) ;
	assign x_884 = (v_685 | ~v_453) ;
	assign x_883 = (v_685 | ~v_452) ;
	assign x_3292 = (x_881 & x_882) ;
	assign x_880 = (v_687 | ~v_686) ;
	assign x_879 = (v_687 | ~v_672) ;
	assign x_878 = (v_688 | ~v_455) ;
	assign x_3287 = (x_876 & x_877) ;
	assign x_875 = (v_688 | ~v_452) ;
	assign x_874 = (v_688 | ~v_500) ;
	assign x_873 = (v_688 | ~v_669) ;
	assign x_872 = (v_689 | ~v_455) ;
	assign x_871 = (v_689 | ~v_454) ;
	assign x_870 = (v_689 | ~v_453) ;
	assign x_869 = (v_689 | ~v_452) ;
	assign x_3277 = (x_867 & x_868) ;
	assign x_866 = ((((((((~v_663 | ~v_662) | ~v_661) | ~v_689) | ~v_688) | ~v_687) | ~v_668) | ~v_395) | v_690) ;
	assign x_865 = (v_691 | ~v_690) ;
	assign x_864 = (v_691 | ~v_390) ;
	assign x_3273 = (x_862 & x_863) ;
	assign x_861 = (v_692 | ~v_6) ;
	assign x_860 = (v_692 | ~v_8) ;
	assign x_859 = (v_693 | ~v_1) ;
	assign x_3268 = (x_857 & x_858) ;
	assign x_856 = (v_693 | ~v_7) ;
	assign x_855 = ((((((((v_7 | v_4) | v_6) | v_8) | v_2) | v_1) | ~v_693) | ~v_692) | ~v_691) ;
	assign x_854 = (v_695 | ~v_14) ;
	assign x_853 = (v_695 | v_25) ;
	assign x_852 = (v_696 | ~v_14) ;
	assign x_851 = (v_696 | v_39) ;
	assign x_850 = (v_697 | v_14) ;
	assign x_3259 = (x_848 & x_849) ;
	assign x_847 = (v_698 | v_42) ;
	assign x_846 = (((((((((((((((v_31 | v_35) | v_37) | v_36) | v_34) | v_79) | v_71) | ~v_173) | ~v_169) | ~v_179) | ~v_176) | ~v_698) | ~v_697) | ~v_696) | ~v_695) | v_699) ;
	assign x_845 = (v_700 | ~v_14) ;
	assign x_3255 = (x_843 & x_844) ;
	assign x_842 = (v_701 | v_52) ;
	assign x_841 = (v_702 | v_14) ;
	assign x_840 = (v_702 | v_28) ;
	assign x_3250 = (x_838 & x_839) ;
	assign x_837 = (((((((((((((((v_50 | v_49) | v_48) | v_74) | v_47) | v_80) | v_44) | ~v_703) | ~v_158) | ~v_157) | ~v_186) | ~v_183) | ~v_702) | ~v_701) | ~v_700) | v_704) ;
	assign x_836 = (v_705 | ~v_14) ;
	assign x_835 = (v_705 | v_27) ;
	assign x_834 = (v_706 | ~v_14) ;
	assign x_833 = (v_706 | v_65) ;
	assign x_832 = (v_707 | v_14) ;
	assign x_831 = (v_707 | v_30) ;
	assign x_3239 = (x_829 & x_830) ;
	assign x_828 = (((((((((((((((v_61 | v_81) | v_63) | v_62) | v_60) | v_57) | v_77) | ~v_194) | ~v_708) | ~v_165) | ~v_164) | ~v_190) | ~v_707) | ~v_706) | ~v_705) | v_709) ;
	assign x_827 = (v_710 | ~v_709) ;
	assign x_826 = (v_710 | ~v_704) ;
	assign x_3235 = (x_824 & x_825) ;
	assign x_823 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_175) | ~v_255) | v_712) ;
	assign x_822 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_148) | ~v_335) | v_713) ;
	assign x_821 = (((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_272) | v_714) ;
	assign x_3230 = (x_819 & x_820) ;
	assign x_818 = (v_715 | ~v_712) ;
	assign x_817 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_120) | ~v_715) | v_716) ;
	assign x_816 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_175) | ~v_318) | v_717) ;
	assign x_815 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_272) | ~v_353) | v_718) ;
	assign x_814 = (((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_335) | v_719) ;
	assign x_813 = (v_720 | ~v_719) ;
	assign x_812 = (v_720 | ~v_718) ;
	assign x_3221 = (x_810 & x_811) ;
	assign x_809 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_272) | ~v_120) | v_722) ;
	assign x_808 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_214) | ~v_335) | v_723) ;
	assign x_807 = (((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_175) | v_724) ;
	assign x_3217 = (x_805 & x_806) ;
	assign x_804 = (v_725 | ~v_722) ;
	assign x_803 = (v_725 | ~v_721) ;
	assign x_802 = (v_725 | ~v_716) ;
	assign x_3212 = (x_800 & x_801) ;
	assign x_799 = (v_727 | ~v_359) ;
	assign x_798 = (v_727 | ~v_358) ;
	assign x_797 = (v_727 | ~v_386) ;
	assign x_796 = (v_727 | ~v_385) ;
	assign x_795 = (v_728 | ~v_724) ;
	assign x_794 = (v_728 | ~v_723) ;
	assign x_793 = (v_728 | ~v_722) ;
	assign x_3202 = (x_791 & x_792) ;
	assign x_790 = (v_731 | ~v_714) ;
	assign x_789 = (v_731 | ~v_713) ;
	assign x_788 = (v_731 | ~v_712) ;
	assign x_3198 = (x_786 & x_787) ;
	assign x_785 = ((~v_731 | ~v_727) | v_732) ;
	assign x_784 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_353) | ~v_715) | v_733) ;
	assign x_783 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_318) | ~v_728) | v_734) ;
	assign x_3193 = (x_781 & x_782) ;
	assign x_780 = (v_735 | ~v_717) ;
	assign x_779 = (v_735 | ~v_734) ;
	assign x_778 = (v_735 | ~v_733) ;
	assign x_777 = ((~v_296 | ~v_735) | v_736) ;
	assign x_776 = (v_737 | ~v_736) ;
	assign x_775 = (v_737 | ~v_732) ;
	assign x_774 = (v_737 | ~v_726) ;
	assign x_3184 = (x_772 & x_773) ;
	assign x_771 = ((~v_25 | v_14) | v_739) ;
	assign x_770 = ((~v_39 | v_14) | v_740) ;
	assign x_769 = ((~v_14 | ~v_29) | v_741) ;
	assign x_768 = ((~v_14 | ~v_42) | v_742) ;
	assign x_767 = (v_743 | ~v_31) ;
	assign x_766 = (v_743 | ~v_34) ;
	assign x_765 = (v_743 | ~v_35) ;
	assign x_3176 = (x_763 & x_764) ;
	assign x_762 = (v_743 | ~v_71) ;
	assign x_761 = (v_743 | ~v_79) ;
	assign x_760 = (v_743 | ~v_476) ;
	assign x_759 = (v_743 | ~v_472) ;
	assign x_758 = (v_743 | ~v_482) ;
	assign x_757 = (v_743 | ~v_479) ;
	assign x_756 = (v_743 | ~v_742) ;
	assign x_3164 = (x_754 & x_755) ;
	assign x_753 = (v_743 | ~v_739) ;
	assign x_752 = ((~v_26 | v_14) | v_744) ;
	assign x_751 = ((v_14 | ~v_52) | v_745) ;
	assign x_3160 = (x_749 & x_750) ;
	assign x_748 = (v_748 | ~v_44) ;
	assign x_747 = (v_748 | ~v_47) ;
	assign x_746 = (v_748 | ~v_48) ;
	assign x_3155 = (x_744 & x_745) ;
	assign x_743 = (v_748 | ~v_74) ;
	assign x_742 = (v_748 | ~v_80) ;
	assign x_741 = (v_748 | ~v_747) ;
	assign x_740 = (v_748 | ~v_461) ;
	assign x_739 = (v_748 | ~v_460) ;
	assign x_738 = (v_748 | ~v_489) ;
	assign x_737 = (v_748 | ~v_486) ;
	assign x_3146 = (x_735 & x_736) ;
	assign x_734 = (v_748 | ~v_744) ;
	assign x_733 = ((~v_27 | v_14) | v_749) ;
	assign x_732 = ((v_14 | ~v_65) | v_750) ;
	assign x_3142 = (x_730 & x_731) ;
	assign x_729 = (v_753 | ~v_57) ;
	assign x_728 = (v_753 | ~v_60) ;
	assign x_727 = (v_753 | ~v_61) ;
	assign x_3137 = (x_725 & x_726) ;
	assign x_724 = (v_753 | ~v_77) ;
	assign x_723 = (v_753 | ~v_81) ;
	assign x_722 = (v_753 | ~v_497) ;
	assign x_721 = (v_753 | ~v_752) ;
	assign x_720 = (v_753 | ~v_468) ;
	assign x_719 = (v_753 | ~v_467) ;
	assign x_718 = (v_753 | ~v_493) ;
	assign x_3127 = (x_716 & x_717) ;
	assign x_715 = (v_753 | ~v_749) ;
	assign x_714 = (((~v_753 | ~v_748) | ~v_743) | v_754) ;
	assign x_713 = (v_755 | ~v_455) ;
	assign x_3123 = (x_711 & x_712) ;
	assign x_710 = (v_755 | ~v_452) ;
	assign x_709 = (v_755 | ~v_754) ;
	assign x_708 = (v_756 | ~v_455) ;
	assign x_3118 = (x_706 & x_707) ;
	assign x_705 = (v_756 | ~v_452) ;
	assign x_704 = (v_756 | ~v_478) ;
	assign x_703 = (v_756 | ~v_558) ;
	assign x_702 = (v_757 | ~v_455) ;
	assign x_701 = (v_757 | ~v_454) ;
	assign x_700 = (v_757 | ~v_453) ;
	assign x_699 = (v_757 | ~v_452) ;
	assign x_3109 = (x_697 & x_698) ;
	assign x_696 = (v_758 | ~v_455) ;
	assign x_695 = (v_758 | ~v_454) ;
	assign x_694 = (v_758 | ~v_453) ;
	assign x_3105 = (x_692 & x_693) ;
	assign x_691 = (((~v_758 | ~v_757) | ~v_756) | v_759) ;
	assign x_690 = (v_760 | ~v_455) ;
	assign x_689 = (v_760 | ~v_454) ;
	assign x_3100 = (x_687 & x_688) ;
	assign x_686 = (v_760 | ~v_423) ;
	assign x_685 = (v_760 | ~v_759) ;
	assign x_684 = (v_761 | ~v_455) ;
	assign x_683 = (v_761 | ~v_454) ;
	assign x_682 = (v_761 | ~v_453) ;
	assign x_681 = (v_761 | ~v_452) ;
	assign x_680 = (v_761 | ~v_478) ;
	assign x_3089 = (x_678 & x_679) ;
	assign x_677 = (v_762 | ~v_454) ;
	assign x_676 = (v_762 | ~v_453) ;
	assign x_675 = (v_762 | ~v_452) ;
	assign x_3085 = (x_673 & x_674) ;
	assign x_672 = (v_763 | ~v_455) ;
	assign x_671 = (v_763 | ~v_454) ;
	assign x_670 = (v_763 | ~v_453) ;
	assign x_3080 = (x_668 & x_669) ;
	assign x_667 = (((~v_763 | ~v_762) | ~v_761) | v_764) ;
	assign x_666 = (v_765 | ~v_455) ;
	assign x_665 = (v_765 | ~v_454) ;
	assign x_664 = (v_765 | ~v_453) ;
	assign x_663 = (v_765 | ~v_452) ;
	assign x_662 = (v_765 | ~v_517) ;
	assign x_661 = (v_765 | ~v_764) ;
	assign x_3071 = (x_659 & x_660) ;
	assign x_658 = (v_766 | ~v_453) ;
	assign x_657 = (v_766 | ~v_452) ;
	assign x_656 = (v_766 | ~v_575) ;
	assign x_3067 = (x_654 & x_655) ;
	assign x_653 = (v_767 | ~v_454) ;
	assign x_652 = (v_767 | ~v_453) ;
	assign x_651 = (v_767 | ~v_452) ;
	assign x_3062 = (x_649 & x_650) ;
	assign x_648 = (v_768 | ~v_455) ;
	assign x_647 = (v_768 | ~v_454) ;
	assign x_646 = (v_768 | ~v_453) ;
	assign x_645 = (v_768 | ~v_452) ;
	assign x_644 = (v_768 | ~v_478) ;
	assign x_643 = (((((~v_768 | ~v_767) | ~v_766) | ~v_765) | ~v_760) | v_769) ;
	assign x_642 = (v_770 | ~v_769) ;
	assign x_3052 = (x_640 & x_641) ;
	assign x_639 = (((~v_768 | ~v_767) | ~v_766) | v_772) ;
	assign x_638 = (v_773 | ~v_455) ;
	assign x_637 = (v_773 | ~v_454) ;
	assign x_3048 = (x_635 & x_636) ;
	assign x_634 = (v_773 | ~v_558) ;
	assign x_633 = (v_773 | ~v_772) ;
	assign x_632 = (v_774 | ~v_455) ;
	assign x_3043 = (x_630 & x_631) ;
	assign x_629 = (v_774 | ~v_452) ;
	assign x_628 = (v_774 | ~v_451) ;
	assign x_627 = (v_774 | ~v_764) ;
	assign x_626 = (((((~v_758 | ~v_757) | ~v_756) | ~v_774) | ~v_773) | v_775) ;
	assign x_625 = (v_776 | ~v_775) ;
	assign x_624 = (v_776 | ~v_771) ;
	assign x_623 = (v_777 | ~v_455) ;
	assign x_3034 = (x_621 & x_622) ;
	assign x_620 = (v_777 | ~v_452) ;
	assign x_619 = (v_777 | ~v_656) ;
	assign x_618 = (v_777 | ~v_759) ;
	assign x_617 = (v_778 | ~v_455) ;
	assign x_616 = (v_778 | ~v_454) ;
	assign x_615 = (v_778 | ~v_453) ;
	assign x_614 = (v_778 | ~v_452) ;
	assign x_3026 = (x_612 & x_613) ;
	assign x_611 = (((((~v_763 | ~v_762) | ~v_761) | ~v_778) | ~v_777) | v_779) ;
	assign x_610 = (v_780 | ~v_599) ;
	assign x_609 = (v_780 | ~v_779) ;
	assign x_608 = (((((~v_780 | ~v_776) | ~v_770) | ~v_755) | ~v_395) | v_781) ;
	assign x_607 = (v_782 | ~v_781) ;
	assign x_606 = (v_782 | ~v_738) ;
	assign x_605 = ((((((((v_7 | v_5) | v_4) | v_8) | v_2) | v_1) | ~v_693) | ~v_692) | ~v_782) ;
	assign x_3012 = (x_603 & x_604) ;
	assign x_602 = (v_785 | ~v_294) ;
	assign x_601 = (v_785 | ~v_293) ;
	assign x_600 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_785) | ~v_272) | v_786) ;
	assign x_3008 = (x_598 & x_599) ;
	assign x_597 = (v_787 | ~v_256) ;
	assign x_596 = (v_787 | ~v_786) ;
	assign x_595 = (v_787 | ~v_784) ;
	assign x_3003 = (x_593 & x_594) ;
	assign x_592 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_785) | ~v_175) | v_790) ;
	assign x_591 = (v_791 | ~v_215) ;
	assign x_590 = (v_791 | ~v_790) ;
	assign x_589 = (v_791 | ~v_789) ;
	assign x_588 = (v_791 | ~v_198) ;
	assign x_587 = (v_791 | ~v_153) ;
	assign x_586 = ((~v_791 | ~v_383) | v_792) ;
	assign x_2994 = (x_584 & x_585) ;
	assign x_583 = (v_793 | ~v_293) ;
	assign x_582 = (v_793 | ~v_292) ;
	assign x_581 = (v_793 | ~v_239) ;
	assign x_2990 = (x_579 & x_580) ;
	assign x_578 = (((((~v_389 | ~v_388) | ~v_793) | ~v_92) | ~v_91) | v_794) ;
	assign x_577 = (v_795 | ~v_455) ;
	assign x_576 = (v_795 | ~v_454) ;
	assign x_2985 = (x_574 & x_575) ;
	assign x_573 = (v_795 | ~v_558) ;
	assign x_572 = (v_795 | ~v_519) ;
	assign x_571 = (((~v_598 | ~v_597) | ~v_596) | v_796) ;
	assign x_570 = (v_797 | ~v_455) ;
	assign x_569 = (v_797 | ~v_454) ;
	assign x_568 = (v_797 | ~v_453) ;
	assign x_567 = (v_797 | ~v_452) ;
	assign x_2975 = (x_565 & x_566) ;
	assign x_564 = (((((~v_577 | ~v_576) | ~v_559) | ~v_797) | ~v_795) | v_798) ;
	assign x_563 = (v_799 | ~v_798) ;
	assign x_562 = (v_799 | ~v_771) ;
	assign x_2971 = (x_560 & x_561) ;
	assign x_559 = (v_800 | ~v_453) ;
	assign x_558 = (v_800 | ~v_452) ;
	assign x_557 = (v_800 | ~v_578) ;
	assign x_2966 = (x_555 & x_556) ;
	assign x_554 = (v_801 | ~v_454) ;
	assign x_553 = (v_801 | ~v_453) ;
	assign x_552 = (v_801 | ~v_452) ;
	assign x_551 = (v_801 | ~v_796) ;
	assign x_550 = (v_801 | ~v_478) ;
	assign x_549 = (((((~v_518 | ~v_801) | ~v_800) | ~v_501) | ~v_456) | v_802) ;
	assign x_548 = (v_803 | ~v_802) ;
	assign x_2957 = (x_546 & x_547) ;
	assign x_545 = (v_805 | ~v_804) ;
	assign x_544 = (v_805 | ~v_794) ;
	assign x_543 = ((((((((v_7 | v_5) | v_4) | v_6) | v_2) | v_1) | ~v_693) | ~v_692) | ~v_805) ;
	assign x_2953 = (x_541 & x_542) ;
	assign x_540 = (v_808 | ~v_381) ;
	assign x_539 = (v_808 | ~v_380) ;
	assign x_538 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_808) | ~v_335) | v_809) ;
	assign x_2948 = (x_536 & x_537) ;
	assign x_535 = (v_810 | ~v_807) ;
	assign x_534 = (v_810 | ~v_371) ;
	assign x_533 = (v_810 | ~v_370) ;
	assign x_532 = ((~v_810 | ~v_296) | v_811) ;
	assign x_531 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_148) | ~v_373) | v_812) ;
	assign x_530 = ((((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_272) | ~v_808) | v_813) ;
	assign x_529 = (v_814 | ~v_377) ;
	assign x_2937 = (x_527 & x_528) ;
	assign x_526 = (v_814 | ~v_813) ;
	assign x_525 = (v_814 | ~v_812) ;
	assign x_524 = ((~v_814 | ~v_727) | v_815) ;
	assign x_2933 = (x_522 & x_523) ;
	assign x_521 = (v_816 | ~v_380) ;
	assign x_520 = (v_816 | ~v_379) ;
	assign x_519 = (v_816 | ~v_374) ;
	assign x_2928 = (x_517 & x_518) ;
	assign x_516 = (((((~v_389 | ~v_388) | ~v_816) | ~v_92) | ~v_91) | v_817) ;
	assign x_515 = (v_818 | ~v_455) ;
	assign x_514 = (v_818 | ~v_454) ;
	assign x_513 = (v_818 | ~v_453) ;
	assign x_512 = (v_818 | ~v_452) ;
	assign x_511 = (v_818 | ~v_681) ;
	assign x_510 = (v_818 | ~v_656) ;
	assign x_2919 = (x_508 & x_509) ;
	assign x_507 = (v_820 | ~v_454) ;
	assign x_506 = (v_820 | ~v_453) ;
	assign x_505 = (v_820 | ~v_452) ;
	assign x_2915 = (x_503 & x_504) ;
	assign x_502 = (((((~v_675 | ~v_820) | ~v_818) | ~v_674) | ~v_673) | v_821) ;
	assign x_501 = (v_822 | ~v_821) ;
	assign x_500 = (v_822 | ~v_599) ;
	assign x_2910 = (x_498 & x_499) ;
	assign x_497 = (v_823 | ~v_453) ;
	assign x_496 = (v_823 | ~v_452) ;
	assign x_495 = (v_823 | ~v_451) ;
	assign x_494 = (v_823 | ~v_676) ;
	assign x_493 = (v_824 | ~v_455) ;
	assign x_492 = (v_824 | ~v_454) ;
	assign x_491 = (v_824 | ~v_453) ;
	assign x_2900 = (x_489 & x_490) ;
	assign x_488 = (v_824 | ~v_819) ;
	assign x_487 = (((((~v_680 | ~v_679) | ~v_678) | ~v_824) | ~v_823) | v_825) ;
	assign x_486 = (v_826 | ~v_825) ;
	assign x_2896 = (x_484 & x_485) ;
	assign x_483 = (v_828 | ~v_827) ;
	assign x_482 = (v_828 | ~v_817) ;
	assign x_481 = ((((((((v_7 | v_5) | v_6) | v_8) | v_2) | v_1) | ~v_693) | ~v_692) | ~v_828) ;
	assign x_2891 = (x_479 & x_480) ;
	assign x_478 = (v_832 | ~v_363) ;
	assign x_477 = (v_832 | ~v_362) ;
	assign x_476 = (v_832 | ~v_357) ;
	assign x_475 = (v_832 | ~v_336) ;
	assign x_474 = (v_832 | ~v_319) ;
	assign x_473 = (v_832 | ~v_831) ;
	assign x_472 = (v_832 | ~v_830) ;
	assign x_2882 = (x_470 & x_471) ;
	assign x_469 = (v_834 | ~v_771) ;
	assign x_468 = (v_835 | ~v_821) ;
	assign x_467 = (v_835 | ~v_672) ;
	assign x_466 = ((((((((~v_666 | ~v_665) | ~v_660) | ~v_639) | ~v_622) | ~v_835) | ~v_834) | ~v_395) | v_836) ;
	assign x_465 = (v_837 | ~v_836) ;
	assign x_464 = (v_837 | ~v_833) ;
	assign x_463 = ((((((((v_4 | v_6) | v_8) | v_3) | v_2) | v_1) | ~v_693) | ~v_692) | ~v_837) ;
	assign x_2874 = (x_461 & x_462) ;
	assign x_460 = (v_841 | ~v_724) ;
	assign x_459 = (v_841 | ~v_723) ;
	assign x_458 = (v_841 | ~v_722) ;
	assign x_457 = (v_841 | ~v_721) ;
	assign x_456 = (v_841 | ~v_716) ;
	assign x_455 = (v_841 | ~v_840) ;
	assign x_454 = (v_841 | ~v_839) ;
	assign x_2862 = (x_452 & x_453) ;
	assign x_451 = (v_843 | ~v_779) ;
	assign x_450 = (v_844 | ~v_775) ;
	assign x_449 = (v_844 | ~v_672) ;
	assign x_2858 = (x_447 & x_448) ;
	assign x_446 = (v_846 | ~v_842) ;
	assign x_445 = ((((((((v_7 | v_5) | v_4) | v_8) | v_3) | v_2) | ~v_693) | ~v_692) | ~v_846) ;
	assign x_444 = ((~v_296 | ~v_725) | v_848) ;
	assign x_2853 = (x_442 & x_443) ;
	assign x_441 = (v_850 | ~v_790) ;
	assign x_440 = (v_850 | ~v_789) ;
	assign x_439 = (v_850 | ~v_198) ;
	assign x_438 = (v_850 | ~v_153) ;
	assign x_437 = (v_850 | ~v_849) ;
	assign x_436 = (v_850 | ~v_848) ;
	assign x_435 = (((((~v_389 | ~v_388) | ~v_850) | ~v_92) | ~v_91) | v_851) ;
	assign x_2844 = (x_433 & x_434) ;
	assign x_432 = (v_853 | ~v_798) ;
	assign x_431 = (v_853 | ~v_672) ;
	assign x_430 = ((((((((~v_518 | ~v_801) | ~v_800) | ~v_501) | ~v_456) | ~v_853) | ~v_852) | ~v_395) | v_854) ;
	assign x_2840 = (x_428 & x_429) ;
	assign x_427 = ((((((((v_7 | v_5) | v_4) | v_6) | v_3) | v_2) | ~v_693) | ~v_692) | ~v_855) ;
	assign x_426 = ((~v_791 | ~v_364) | v_857) ;
	assign x_425 = ((~v_725 | ~v_727) | v_858) ;
	assign x_2835 = (x_423 & x_424) ;
	assign x_422 = (v_859 | ~v_337) ;
	assign x_421 = (v_859 | ~v_368) ;
	assign x_420 = (v_859 | ~v_367) ;
	assign x_419 = (v_859 | ~v_858) ;
	assign x_418 = (v_859 | ~v_857) ;
	assign x_417 = (((((~v_389 | ~v_388) | ~v_859) | ~v_92) | ~v_91) | v_860) ;
	assign x_416 = (v_861 | ~v_802) ;
	assign x_2825 = (x_414 & x_415) ;
	assign x_413 = (v_862 | ~v_771) ;
	assign x_412 = ((((((((~v_658 | ~v_657) | ~v_640) | ~v_671) | ~v_670) | ~v_862) | ~v_861) | ~v_395) | v_863) ;
	assign x_411 = (v_864 | ~v_863) ;
	assign x_2821 = (x_409 & x_410) ;
	assign x_408 = (v_866 | ~v_24) ;
	assign x_407 = (v_866 | v_39) ;
	assign x_406 = (v_867 | v_24) ;
	assign x_2816 = (x_404 & x_405) ;
	assign x_403 = (v_868 | v_42) ;
	assign x_402 = (v_869 | ~v_24) ;
	assign x_401 = (v_869 | v_25) ;
	assign x_400 = (((((((((((((((v_31 | v_37) | v_36) | v_79) | v_71) | v_85) | ~v_869) | v_88) | ~v_236) | ~v_98) | ~v_97) | ~v_234) | ~v_868) | ~v_867) | ~v_866) | v_870) ;
	assign x_399 = (v_871 | ~v_24) ;
	assign x_398 = (v_871 | v_26) ;
	assign x_397 = (v_872 | ~v_24) ;
	assign x_2807 = (x_395 & x_396) ;
	assign x_394 = (v_873 | v_28) ;
	assign x_393 = (v_874 | v_24) ;
	assign x_392 = (v_874 | v_55) ;
	assign x_2803 = (x_390 & x_391) ;
	assign x_389 = (v_876 | v_27) ;
	assign x_388 = (v_877 | ~v_24) ;
	assign x_387 = (v_877 | v_65) ;
	assign x_2798 = (x_385 & x_386) ;
	assign x_384 = (v_879 | v_24) ;
	assign x_383 = (v_879 | v_68) ;
	assign x_382 = (((((((((((((((v_81 | v_63) | v_62) | v_57) | v_77) | ~v_117) | v_90) | v_87) | ~v_115) | ~v_227) | ~v_226) | ~v_879) | ~v_878) | ~v_877) | ~v_876) | v_880) ;
	assign x_381 = (v_881 | ~v_880) ;
	assign x_380 = (v_881 | ~v_875) ;
	assign x_379 = (v_881 | ~v_870) ;
	assign x_378 = (((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_881) | v_882) ;
	assign x_2787 = (x_376 & x_377) ;
	assign x_375 = (v_885 | ~v_884) ;
	assign x_374 = (v_885 | ~v_883) ;
	assign x_373 = (v_885 | ~v_726) ;
	assign x_2783 = (x_371 & x_372) ;
	assign x_370 = ((~v_39 | v_24) | v_887) ;
	assign x_369 = ((~v_24 | ~v_29) | v_888) ;
	assign x_368 = ((~v_24 | ~v_42) | v_889) ;
	assign x_2778 = (x_366 & x_367) ;
	assign x_365 = (v_891 | ~v_36) ;
	assign x_364 = (v_891 | ~v_37) ;
	assign x_363 = (v_891 | ~v_71) ;
	assign x_362 = (v_891 | ~v_79) ;
	assign x_361 = (v_891 | ~v_85) ;
	assign x_360 = (v_891 | ~v_890) ;
	assign x_359 = (v_891 | ~v_88) ;
	assign x_2769 = (x_357 & x_358) ;
	assign x_356 = (v_891 | ~v_400) ;
	assign x_355 = (v_891 | ~v_537) ;
	assign x_354 = (v_891 | ~v_889) ;
	assign x_2765 = (x_352 & x_353) ;
	assign x_351 = ((~v_26 | v_24) | v_892) ;
	assign x_350 = ((v_24 | ~v_52) | v_893) ;
	assign x_349 = ((~v_24 | ~v_28) | v_894) ;
	assign x_2760 = (x_347 & x_348) ;
	assign x_346 = (v_896 | ~v_49) ;
	assign x_345 = (v_896 | ~v_50) ;
	assign x_344 = (v_896 | ~v_74) ;
	assign x_343 = (v_896 | ~v_80) ;
	assign x_342 = (v_896 | ~v_86) ;
	assign x_341 = (v_896 | ~v_525) ;
	assign x_340 = (v_896 | ~v_89) ;
	assign x_2750 = (x_338 & x_339) ;
	assign x_337 = (v_896 | ~v_522) ;
	assign x_336 = (v_896 | ~v_895) ;
	assign x_335 = (v_896 | ~v_894) ;
	assign x_2746 = (x_333 & x_334) ;
	assign x_332 = ((~v_27 | v_24) | v_897) ;
	assign x_331 = ((v_24 | ~v_65) | v_898) ;
	assign x_330 = ((~v_24 | ~v_30) | v_899) ;
	assign x_2741 = (x_328 & x_329) ;
	assign x_327 = (v_901 | ~v_62) ;
	assign x_326 = (v_901 | ~v_63) ;
	assign x_325 = (v_901 | ~v_77) ;
	assign x_324 = (v_901 | ~v_81) ;
	assign x_323 = (v_901 | ~v_420) ;
	assign x_322 = (v_901 | ~v_87) ;
	assign x_321 = (v_901 | ~v_90) ;
	assign x_2732 = (x_319 & x_320) ;
	assign x_318 = (v_901 | ~v_529) ;
	assign x_317 = (v_901 | ~v_900) ;
	assign x_316 = (v_901 | ~v_899) ;
	assign x_315 = (v_901 | ~v_898) ;
	assign x_314 = (v_901 | ~v_897) ;
	assign x_313 = (((~v_901 | ~v_896) | ~v_891) | v_902) ;
	assign x_312 = (v_903 | ~v_455) ;
	assign x_2724 = (x_310 & x_311) ;
	assign x_309 = (v_903 | ~v_452) ;
	assign x_308 = (v_903 | ~v_902) ;
	assign x_307 = (v_904 | ~v_825) ;
	assign x_306 = (v_904 | ~v_672) ;
	assign x_305 = (v_905 | ~v_802) ;
	assign x_304 = (v_905 | ~v_821) ;
	assign x_303 = (((((~v_905 | ~v_904) | ~v_770) | ~v_903) | ~v_395) | v_906) ;
	assign x_2711 = (x_301 & x_302) ;
	assign x_300 = ((((((((v_7 | v_5) | v_6) | v_8) | v_3) | v_2) | ~v_693) | ~v_692) | ~v_907) ;
	assign x_299 = (v_909 | ~v_19) ;
	assign x_298 = (v_909 | v_39) ;
	assign x_2707 = (x_296 & x_297) ;
	assign x_295 = (v_911 | ~v_19) ;
	assign x_294 = (v_911 | v_25) ;
	assign x_293 = (v_912 | v_19) ;
	assign x_2702 = (x_291 & x_292) ;
	assign x_290 = (v_914 | ~v_19) ;
	assign x_289 = (v_914 | v_52) ;
	assign x_288 = (v_915 | v_19) ;
	assign x_287 = (v_915 | v_28) ;
	assign x_286 = (v_916 | v_19) ;
	assign x_285 = (v_916 | v_55) ;
	assign x_284 = (v_917 | ~v_19) ;
	assign x_2693 = (x_282 & x_283) ;
	assign x_281 = (v_919 | v_19) ;
	assign x_280 = (v_919 | v_30) ;
	assign x_279 = (v_920 | v_19) ;
	assign x_2689 = (x_277 & x_278) ;
	assign x_276 = (v_921 | v_27) ;
	assign x_275 = (v_922 | ~v_19) ;
	assign x_274 = (v_922 | v_65) ;
	assign x_2684 = (x_272 & x_273) ;
	assign x_271 = (v_924 | ~v_918) ;
	assign x_270 = (v_924 | ~v_913) ;
	assign x_269 = (((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_924) | v_925) ;
	assign x_268 = ((~v_787 | ~v_364) | v_926) ;
	assign x_267 = (v_927 | ~v_926) ;
	assign x_266 = (v_927 | ~v_883) ;
	assign x_265 = (v_927 | ~v_732) ;
	assign x_2674 = (x_263 & x_264) ;
	assign x_262 = ((~v_39 | v_19) | v_929) ;
	assign x_261 = ((~v_19 | ~v_29) | v_930) ;
	assign x_260 = ((~v_25 | v_19) | v_931) ;
	assign x_2670 = (x_258 & x_259) ;
	assign x_257 = (v_933 | ~v_34) ;
	assign x_256 = (v_933 | ~v_35) ;
	assign x_255 = (v_933 | ~v_36) ;
	assign x_2665 = (x_253 & x_254) ;
	assign x_252 = (v_933 | ~v_79) ;
	assign x_251 = (v_933 | ~v_430) ;
	assign x_250 = (v_933 | ~v_402) ;
	assign x_249 = (v_933 | ~v_932) ;
	assign x_248 = (v_933 | ~v_931) ;
	assign x_247 = (v_933 | ~v_424) ;
	assign x_246 = (v_933 | ~v_399) ;
	assign x_2656 = (x_244 & x_245) ;
	assign x_243 = ((v_19 | ~v_52) | v_934) ;
	assign x_242 = ((~v_19 | ~v_28) | v_935) ;
	assign x_241 = ((~v_19 | ~v_55) | v_936) ;
	assign x_2652 = (x_239 & x_240) ;
	assign x_238 = (v_938 | ~v_47) ;
	assign x_237 = (v_938 | ~v_48) ;
	assign x_236 = (v_938 | ~v_49) ;
	assign x_2647 = (x_234 & x_235) ;
	assign x_233 = (v_938 | ~v_80) ;
	assign x_232 = (v_938 | ~v_412) ;
	assign x_231 = (v_938 | ~v_937) ;
	assign x_230 = (v_938 | ~v_434) ;
	assign x_229 = (v_938 | ~v_433) ;
	assign x_228 = (v_938 | ~v_409) ;
	assign x_227 = (v_938 | ~v_936) ;
	assign x_2636 = (x_225 & x_226) ;
	assign x_224 = ((~v_19 | ~v_30) | v_939) ;
	assign x_223 = ((~v_19 | ~v_68) | v_940) ;
	assign x_222 = ((~v_27 | v_19) | v_941) ;
	assign x_2632 = (x_220 & x_221) ;
	assign x_219 = (v_943 | ~v_60) ;
	assign x_218 = (v_943 | ~v_61) ;
	assign x_217 = (v_943 | ~v_62) ;
	assign x_2627 = (x_215 & x_216) ;
	assign x_214 = (v_943 | ~v_81) ;
	assign x_213 = (v_943 | ~v_421) ;
	assign x_212 = (v_943 | ~v_942) ;
	assign x_211 = (v_943 | ~v_446) ;
	assign x_210 = (v_943 | ~v_941) ;
	assign x_209 = (v_943 | ~v_419) ;
	assign x_208 = (v_943 | ~v_442) ;
	assign x_2618 = (x_206 & x_207) ;
	assign x_205 = (((~v_943 | ~v_938) | ~v_933) | v_944) ;
	assign x_204 = (v_945 | ~v_455) ;
	assign x_203 = (v_945 | ~v_454) ;
	assign x_2614 = (x_201 & x_202) ;
	assign x_200 = (v_945 | ~v_944) ;
	assign x_199 = (v_946 | ~v_798) ;
	assign x_198 = (v_946 | ~v_667) ;
	assign x_2609 = (x_196 & x_197) ;
	assign x_195 = (v_948 | ~v_928) ;
	assign x_194 = ((((((((v_7 | v_4) | v_6) | v_8) | v_3) | v_1) | ~v_693) | ~v_692) | ~v_948) ;
	assign x_193 = ((~v_787 | ~v_735) | v_950) ;
	assign x_192 = ((~v_725 | ~v_814) | v_951) ;
	assign x_191 = (v_952 | ~v_714) ;
	assign x_190 = (v_952 | ~v_713) ;
	assign x_189 = (v_952 | ~v_712) ;
	assign x_2599 = (x_187 & x_188) ;
	assign x_186 = (v_952 | ~v_951) ;
	assign x_185 = (v_952 | ~v_950) ;
	assign x_184 = (((((~v_389 | ~v_388) | ~v_952) | ~v_92) | ~v_91) | v_953) ;
	assign x_2595 = (x_182 & x_183) ;
	assign x_181 = (v_955 | ~v_769) ;
	assign x_180 = (v_955 | ~v_825) ;
	assign x_179 = ((((((((~v_758 | ~v_757) | ~v_756) | ~v_774) | ~v_773) | ~v_955) | ~v_954) | ~v_395) | v_956) ;
	assign x_2590 = (x_177 & x_178) ;
	assign x_176 = ((((((((v_7 | v_5) | v_4) | v_8) | v_3) | v_1) | ~v_693) | ~v_692) | ~v_957) ;
	assign x_175 = ((~v_296 | ~v_731) | v_959) ;
	assign x_174 = ((~v_791 | ~v_814) | v_960) ;
	assign x_173 = (v_961 | ~v_274) ;
	assign x_172 = (v_961 | ~v_273) ;
	assign x_171 = (v_961 | ~v_256) ;
	assign x_170 = (v_961 | ~v_786) ;
	assign x_2581 = (x_168 & x_169) ;
	assign x_167 = (v_961 | ~v_959) ;
	assign x_166 = (((((~v_389 | ~v_388) | ~v_961) | ~v_92) | ~v_91) | v_962) ;
	assign x_165 = (v_963 | ~v_599) ;
	assign x_164 = (v_963 | ~v_775) ;
	assign x_163 = (v_964 | ~v_802) ;
	assign x_162 = (v_964 | ~v_825) ;
	assign x_161 = ((((((((~v_577 | ~v_576) | ~v_559) | ~v_797) | ~v_795) | ~v_964) | ~v_963) | ~v_395) | v_965) ;
	assign x_2573 = (x_159 & x_160) ;
	assign x_158 = ((((((((v_7 | v_5) | v_4) | v_6) | v_3) | v_1) | ~v_693) | ~v_692) | ~v_966) ;
	assign x_157 = ((~v_810 | ~v_787) | v_968) ;
	assign x_156 = ((~v_731 | ~v_383) | v_969) ;
	assign x_155 = (v_970 | ~v_377) ;
	assign x_154 = (v_970 | ~v_376) ;
	assign x_153 = (v_970 | ~v_375) ;
	assign x_152 = (v_970 | ~v_813) ;
	assign x_2561 = (x_150 & x_151) ;
	assign x_149 = (v_970 | ~v_968) ;
	assign x_148 = (((((~v_389 | ~v_388) | ~v_970) | ~v_92) | ~v_91) | v_971) ;
	assign x_147 = (v_972 | ~v_821) ;
	assign x_2557 = (x_145 & x_146) ;
	assign x_144 = (v_973 | ~v_686) ;
	assign x_143 = ((((((((~v_680 | ~v_679) | ~v_678) | ~v_824) | ~v_823) | ~v_973) | ~v_972) | ~v_395) | v_974) ;
	assign x_142 = (v_975 | ~v_974) ;
	assign x_2552 = (x_140 & x_141) ;
	assign x_139 = ((~v_735 | ~v_383) | v_977) ;
	assign x_138 = ((~v_364 | ~v_814) | v_978) ;
	assign x_137 = (v_979 | ~v_372) ;
	assign x_136 = (v_979 | ~v_809) ;
	assign x_135 = (v_979 | ~v_807) ;
	assign x_134 = (v_979 | ~v_371) ;
	assign x_133 = (v_979 | ~v_370) ;
	assign x_2543 = (x_131 & x_132) ;
	assign x_130 = (((((~v_389 | ~v_388) | ~v_979) | ~v_92) | ~v_91) | v_980) ;
	assign x_129 = (v_981 | ~v_779) ;
	assign x_128 = (v_981 | ~v_686) ;
	assign x_2539 = (x_126 & x_127) ;
	assign x_125 = ((((((((~v_675 | ~v_820) | ~v_818) | ~v_674) | ~v_673) | ~v_982) | ~v_981) | ~v_395) | v_983) ;
	assign x_124 = (v_984 | ~v_983) ;
	assign x_123 = (v_984 | ~v_980) ;
	assign x_2534 = (x_121 & x_122) ;
	assign x_120 = ((~v_810 | ~v_725) | v_987) ;
	assign x_119 = (v_988 | ~v_719) ;
	assign x_118 = (v_988 | ~v_718) ;
	assign x_117 = (v_988 | ~v_717) ;
	assign x_116 = (v_988 | ~v_734) ;
	assign x_115 = (v_988 | ~v_733) ;
	assign x_114 = (v_988 | ~v_987) ;
	assign x_2524 = (x_112 & x_113) ;
	assign x_111 = (v_990 | ~v_667) ;
	assign x_110 = (v_990 | ~v_775) ;
	assign x_109 = (v_991 | ~v_821) ;
	assign x_2520 = (x_107 & x_108) ;
	assign x_106 = (v_993 | ~v_992) ;
	assign x_105 = (v_993 | ~v_989) ;
	assign x_104 = ((((((((v_5 | v_4) | v_8) | v_3) | v_2) | v_1) | ~v_693) | ~v_692) | ~v_993) ;
	assign x_2515 = (x_102 & x_103) ;
	assign x_101 = (v_996 | ~v_9) ;
	assign x_100 = (v_996 | v_39) ;
	assign x_99 = (v_997 | v_9) ;
	assign x_98 = (v_997 | v_29) ;
	assign x_97 = (v_998 | ~v_9) ;
	assign x_96 = (v_998 | v_25) ;
	assign x_95 = (((((((((((((((v_32 | v_31) | v_33) | v_35) | v_37) | v_36) | v_34) | ~v_998) | ~v_302) | ~v_997) | ~v_996) | ~v_300) | ~v_125) | ~v_124) | ~v_995) | v_999) ;
	assign x_2506 = (x_93 & x_94) ;
	assign x_92 = (v_1001 | v_9) ;
	assign x_91 = (v_1001 | v_55) ;
	assign x_90 = (v_1002 | ~v_9) ;
	assign x_2502 = (x_88 & x_89) ;
	assign x_87 = (v_1003 | v_28) ;
	assign x_86 = (((((((((((((((~v_1003 | v_50) | v_49) | v_48) | v_46) | v_45) | v_47) | v_44) | ~v_309) | ~v_137) | ~v_1002) | ~v_1001) | ~v_305) | ~v_134) | ~v_1000) | v_1004) ;
	assign x_85 = (v_1005 | ~v_9) ;
	assign x_2497 = (x_83 & x_84) ;
	assign x_82 = (v_1006 | v_27) ;
	assign x_81 = (v_1007 | v_9) ;
	assign x_80 = (v_1007 | v_68) ;
	assign x_79 = (v_1008 | v_9) ;
	assign x_78 = (v_1008 | v_30) ;
	assign x_77 = (((((((((((((((~v_1008 | v_61) | v_63) | v_62) | v_60) | v_59) | v_58) | v_57) | ~v_1007) | ~v_315) | ~v_1006) | ~v_313) | ~v_142) | ~v_141) | ~v_1005) | v_1009) ;
	assign x_76 = (v_1010 | ~v_1009) ;
	assign x_2486 = (x_74 & x_75) ;
	assign x_73 = (((((~v_152 | ~v_151) | ~v_150) | ~v_149) | ~v_1010) | v_1011) ;
	assign x_72 = (v_1012 | ~v_884) ;
	assign x_71 = (v_1012 | ~v_926) ;
	assign x_2482 = (x_69 & x_70) ;
	assign x_68 = (((((~v_389 | ~v_388) | ~v_1012) | ~v_92) | ~v_91) | v_1013) ;
	assign x_67 = ((~v_9 | ~v_42) | v_1014) ;
	assign x_66 = ((~v_39 | v_9) | v_1015) ;
	assign x_2477 = (x_64 & x_65) ;
	assign x_63 = (v_1018 | ~v_31) ;
	assign x_62 = (v_1018 | ~v_32) ;
	assign x_61 = (v_1018 | ~v_33) ;
	assign x_60 = (v_1018 | ~v_34) ;
	assign x_59 = (v_1018 | ~v_35) ;
	assign x_58 = (v_1018 | ~v_36) ;
	assign x_57 = (v_1018 | ~v_37) ;
	assign x_2468 = (x_55 & x_56) ;
	assign x_54 = (v_1018 | ~v_1016) ;
	assign x_53 = (v_1018 | ~v_1015) ;
	assign x_52 = (v_1018 | ~v_603) ;
	assign x_2464 = (x_50 & x_51) ;
	assign x_49 = (v_1018 | ~v_1014) ;
	assign x_48 = ((v_9 | ~v_52) | v_1019) ;
	assign x_47 = ((~v_9 | ~v_55) | v_1020) ;
	assign x_2459 = (x_45 & x_46) ;
	assign x_44 = (v_1023 | ~v_1022) ;
	assign x_43 = (v_1023 | ~v_44) ;
	assign x_42 = (v_1023 | ~v_45) ;
	assign x_41 = (v_1023 | ~v_46) ;
	assign x_40 = (v_1023 | ~v_47) ;
	assign x_39 = (v_1023 | ~v_48) ;
	assign x_38 = (v_1023 | ~v_49) ;
	assign x_2449 = (x_36 & x_37) ;
	assign x_35 = (v_1023 | ~v_440) ;
	assign x_34 = (v_1023 | ~v_1021) ;
	assign x_33 = (v_1023 | ~v_1020) ;
	assign x_2445 = (x_31 & x_32) ;
	assign x_30 = (v_1023 | ~v_1019) ;
	assign x_29 = ((v_9 | ~v_65) | v_1024) ;
	assign x_28 = ((~v_27 | v_9) | v_1025) ;
	assign x_2440 = (x_26 & x_27) ;
	assign x_25 = (v_1028 | ~v_1027) ;
	assign x_24 = (v_1028 | ~v_57) ;
	assign x_23 = (v_1028 | ~v_58) ;
	assign x_22 = (v_1028 | ~v_59) ;
	assign x_21 = (v_1028 | ~v_60) ;
	assign x_20 = (v_1028 | ~v_61) ;
	assign x_19 = (v_1028 | ~v_62) ;
	assign x_2431 = (x_17 & x_18) ;
	assign x_16 = (v_1028 | ~v_618) ;
	assign x_15 = (v_1028 | ~v_1025) ;
	assign x_14 = (v_1028 | ~v_616) ;
	assign x_13 = (v_1028 | ~v_445) ;
	assign x_12 = (v_1028 | ~v_444) ;
	assign x_11 = (v_1028 | ~v_1024) ;
	assign x_10 = (((~v_1028 | ~v_1023) | ~v_1018) | v_1029) ;
	assign x_2423 = (x_8 & x_9) ;
	assign x_7 = (v_1030 | ~v_453) ;
	assign x_6 = (v_1030 | ~v_452) ;
	assign x_5 = (v_1030 | ~v_1029) ;
	assign x_4 = (((((~v_905 | ~v_946) | ~v_780) | ~v_1030) | ~v_395) | v_1031) ;
	assign x_3 = (v_1032 | ~v_1031) ;
	assign x_2 = (v_1032 | ~v_1013) ;
	assign x_1 = ((((((((v_5 | v_4) | v_6) | v_3) | v_2) | v_1) | ~v_693) | ~v_692) | ~v_1032) ;
	assign x_4825 = (x_2416 & x_4824) ;
	assign x_4823 = (x_2414 & x_2415) ;
	assign x_4821 = (x_2411 & x_4820) ;
	assign x_4819 = (x_2409 & x_2410) ;
	assign x_4816 = (x_2406 & x_4815) ;
	assign x_4814 = (x_2404 & x_2405) ;
	assign x_4812 = (x_2402 & x_2403) ;
	assign x_4811 = (x_2400 & x_2401) ;
	assign x_4807 = (x_2397 & x_4806) ;
	assign x_4805 = (x_2395 & x_2396) ;
	assign x_4803 = (x_2392 & x_4802) ;
	assign x_4801 = (x_2390 & x_2391) ;
	assign x_4798 = (x_2387 & x_4797) ;
	assign x_4796 = (x_2385 & x_2386) ;
	assign x_4794 = (x_2383 & x_2384) ;
	assign x_4793 = (x_2381 & x_2382) ;
	assign x_4788 = (x_2378 & x_4787) ;
	assign x_4786 = (x_2376 & x_2377) ;
	assign x_4784 = (x_2373 & x_4783) ;
	assign x_4782 = (x_2371 & x_2372) ;
	assign x_4779 = (x_2368 & x_4778) ;
	assign x_4777 = (x_2366 & x_2367) ;
	assign x_4775 = (x_2364 & x_2365) ;
	assign x_4774 = (x_2362 & x_2363) ;
	assign x_4770 = (x_2359 & x_4769) ;
	assign x_4768 = (x_2357 & x_2358) ;
	assign x_4766 = (x_2354 & x_4765) ;
	assign x_4764 = (x_2352 & x_2353) ;
	assign x_4761 = (x_2349 & x_4760) ;
	assign x_4759 = (x_2347 & x_2348) ;
	assign x_4757 = (x_2345 & x_2346) ;
	assign x_4756 = (x_2343 & x_2344) ;
	assign x_4750 = (x_2340 & x_4749) ;
	assign x_4748 = (x_2338 & x_2339) ;
	assign x_4746 = (x_2335 & x_4745) ;
	assign x_4744 = (x_2333 & x_2334) ;
	assign x_4741 = (x_2330 & x_4740) ;
	assign x_4739 = (x_2328 & x_2329) ;
	assign x_4737 = (x_2326 & x_2327) ;
	assign x_4736 = (x_2324 & x_2325) ;
	assign x_4732 = (x_2321 & x_4731) ;
	assign x_4730 = (x_2319 & x_2320) ;
	assign x_4728 = (x_2316 & x_4727) ;
	assign x_4726 = (x_2314 & x_2315) ;
	assign x_4723 = (x_2311 & x_4722) ;
	assign x_4721 = (x_2309 & x_2310) ;
	assign x_4719 = (x_2307 & x_2308) ;
	assign x_4718 = (x_2305 & x_2306) ;
	assign x_4713 = (x_2302 & x_4712) ;
	assign x_4711 = (x_2300 & x_2301) ;
	assign x_4709 = (x_2297 & x_4708) ;
	assign x_4707 = (x_2295 & x_2296) ;
	assign x_4704 = (x_2292 & x_4703) ;
	assign x_4702 = (x_2290 & x_2291) ;
	assign x_4700 = (x_2288 & x_2289) ;
	assign x_4699 = (x_2286 & x_2287) ;
	assign x_4695 = (x_2283 & x_4694) ;
	assign x_4693 = (x_2281 & x_2282) ;
	assign x_4691 = (x_2278 & x_4690) ;
	assign x_4689 = (x_2276 & x_2277) ;
	assign x_4686 = (x_2273 & x_4685) ;
	assign x_4684 = (x_2271 & x_2272) ;
	assign x_4682 = (x_2269 & x_2270) ;
	assign x_4681 = (x_2267 & x_2268) ;
	assign x_4674 = (x_2264 & x_4673) ;
	assign x_4672 = (x_2262 & x_2263) ;
	assign x_4670 = (x_2259 & x_4669) ;
	assign x_4668 = (x_2257 & x_2258) ;
	assign x_4665 = (x_2254 & x_4664) ;
	assign x_4663 = (x_2252 & x_2253) ;
	assign x_4661 = (x_2250 & x_2251) ;
	assign x_4660 = (x_2248 & x_2249) ;
	assign x_4656 = (x_2245 & x_4655) ;
	assign x_4654 = (x_2243 & x_2244) ;
	assign x_4652 = (x_2240 & x_4651) ;
	assign x_4650 = (x_2238 & x_2239) ;
	assign x_4647 = (x_2235 & x_4646) ;
	assign x_4645 = (x_2233 & x_2234) ;
	assign x_4643 = (x_2231 & x_2232) ;
	assign x_4642 = (x_2229 & x_2230) ;
	assign x_4637 = (x_2226 & x_4636) ;
	assign x_4635 = (x_2224 & x_2225) ;
	assign x_4633 = (x_2221 & x_4632) ;
	assign x_4631 = (x_2219 & x_2220) ;
	assign x_4628 = (x_2216 & x_4627) ;
	assign x_4626 = (x_2214 & x_2215) ;
	assign x_4624 = (x_2212 & x_2213) ;
	assign x_4623 = (x_2210 & x_2211) ;
	assign x_4619 = (x_2207 & x_4618) ;
	assign x_4617 = (x_2205 & x_2206) ;
	assign x_4615 = (x_2202 & x_4614) ;
	assign x_4613 = (x_2200 & x_2201) ;
	assign x_4610 = (x_2197 & x_4609) ;
	assign x_4608 = (x_2195 & x_2196) ;
	assign x_4606 = (x_2193 & x_2194) ;
	assign x_4605 = (x_2191 & x_2192) ;
	assign x_4599 = (x_2188 & x_4598) ;
	assign x_4597 = (x_2186 & x_2187) ;
	assign x_4595 = (x_2183 & x_4594) ;
	assign x_4593 = (x_2181 & x_2182) ;
	assign x_4590 = (x_2178 & x_4589) ;
	assign x_4588 = (x_2176 & x_2177) ;
	assign x_4586 = (x_2174 & x_2175) ;
	assign x_4585 = (x_2172 & x_2173) ;
	assign x_4581 = (x_2169 & x_4580) ;
	assign x_4579 = (x_2167 & x_2168) ;
	assign x_4577 = (x_2164 & x_4576) ;
	assign x_4575 = (x_2162 & x_2163) ;
	assign x_4572 = (x_2159 & x_4571) ;
	assign x_4570 = (x_2157 & x_2158) ;
	assign x_4568 = (x_2155 & x_2156) ;
	assign x_4567 = (x_2153 & x_2154) ;
	assign x_4562 = (x_2150 & x_4561) ;
	assign x_4560 = (x_2148 & x_2149) ;
	assign x_4558 = (x_2145 & x_4557) ;
	assign x_4556 = (x_2143 & x_2144) ;
	assign x_4553 = (x_2140 & x_4552) ;
	assign x_4551 = (x_2138 & x_2139) ;
	assign x_4549 = (x_2136 & x_2137) ;
	assign x_4548 = (x_2134 & x_2135) ;
	assign x_4544 = (x_2131 & x_4543) ;
	assign x_4542 = (x_2129 & x_2130) ;
	assign x_4540 = (x_2127 & x_2128) ;
	assign x_4539 = (x_2125 & x_2126) ;
	assign x_4536 = (x_2122 & x_4535) ;
	assign x_4534 = (x_2120 & x_2121) ;
	assign x_4532 = (x_2118 & x_2119) ;
	assign x_4531 = (x_2116 & x_2117) ;
	assign x_4523 = (x_2113 & x_4522) ;
	assign x_4521 = (x_2111 & x_2112) ;
	assign x_4519 = (x_2108 & x_4518) ;
	assign x_4517 = (x_2106 & x_2107) ;
	assign x_4514 = (x_2103 & x_4513) ;
	assign x_4512 = (x_2101 & x_2102) ;
	assign x_4510 = (x_2099 & x_2100) ;
	assign x_4509 = (x_2097 & x_2098) ;
	assign x_4505 = (x_2094 & x_4504) ;
	assign x_4503 = (x_2092 & x_2093) ;
	assign x_4501 = (x_2089 & x_4500) ;
	assign x_4499 = (x_2087 & x_2088) ;
	assign x_4496 = (x_2084 & x_4495) ;
	assign x_4494 = (x_2082 & x_2083) ;
	assign x_4492 = (x_2080 & x_2081) ;
	assign x_4491 = (x_2078 & x_2079) ;
	assign x_4486 = (x_2075 & x_4485) ;
	assign x_4484 = (x_2073 & x_2074) ;
	assign x_4482 = (x_2070 & x_4481) ;
	assign x_4480 = (x_2068 & x_2069) ;
	assign x_4477 = (x_2065 & x_4476) ;
	assign x_4475 = (x_2063 & x_2064) ;
	assign x_4473 = (x_2061 & x_2062) ;
	assign x_4472 = (x_2059 & x_2060) ;
	assign x_4468 = (x_2056 & x_4467) ;
	assign x_4466 = (x_2054 & x_2055) ;
	assign x_4464 = (x_2051 & x_4463) ;
	assign x_4462 = (x_2049 & x_2050) ;
	assign x_4459 = (x_2046 & x_4458) ;
	assign x_4457 = (x_2044 & x_2045) ;
	assign x_4455 = (x_2042 & x_2043) ;
	assign x_4454 = (x_2040 & x_2041) ;
	assign x_4448 = (x_2037 & x_4447) ;
	assign x_4446 = (x_2035 & x_2036) ;
	assign x_4444 = (x_2032 & x_4443) ;
	assign x_4442 = (x_2030 & x_2031) ;
	assign x_4439 = (x_2027 & x_4438) ;
	assign x_4437 = (x_2025 & x_2026) ;
	assign x_4435 = (x_2023 & x_2024) ;
	assign x_4434 = (x_2021 & x_2022) ;
	assign x_4430 = (x_2018 & x_4429) ;
	assign x_4428 = (x_2016 & x_2017) ;
	assign x_4426 = (x_2013 & x_4425) ;
	assign x_4424 = (x_2011 & x_2012) ;
	assign x_4421 = (x_2008 & x_4420) ;
	assign x_4419 = (x_2006 & x_2007) ;
	assign x_4417 = (x_2004 & x_2005) ;
	assign x_4416 = (x_2002 & x_2003) ;
	assign x_4411 = (x_1999 & x_4410) ;
	assign x_4409 = (x_1997 & x_1998) ;
	assign x_4407 = (x_1994 & x_4406) ;
	assign x_4405 = (x_1992 & x_1993) ;
	assign x_4402 = (x_1989 & x_4401) ;
	assign x_4400 = (x_1987 & x_1988) ;
	assign x_4398 = (x_1985 & x_1986) ;
	assign x_4397 = (x_1983 & x_1984) ;
	assign x_4393 = (x_1980 & x_4392) ;
	assign x_4391 = (x_1978 & x_1979) ;
	assign x_4389 = (x_1976 & x_1977) ;
	assign x_4388 = (x_1974 & x_1975) ;
	assign x_4385 = (x_1971 & x_4384) ;
	assign x_4383 = (x_1969 & x_1970) ;
	assign x_4381 = (x_1967 & x_1968) ;
	assign x_4380 = (x_1965 & x_1966) ;
	assign x_4373 = (x_1962 & x_4372) ;
	assign x_4371 = (x_1960 & x_1961) ;
	assign x_4369 = (x_1957 & x_4368) ;
	assign x_4367 = (x_1955 & x_1956) ;
	assign x_4364 = (x_1952 & x_4363) ;
	assign x_4362 = (x_1950 & x_1951) ;
	assign x_4360 = (x_1948 & x_1949) ;
	assign x_4359 = (x_1946 & x_1947) ;
	assign x_4355 = (x_1943 & x_4354) ;
	assign x_4353 = (x_1941 & x_1942) ;
	assign x_4351 = (x_1938 & x_4350) ;
	assign x_4349 = (x_1936 & x_1937) ;
	assign x_4346 = (x_1933 & x_4345) ;
	assign x_4344 = (x_1931 & x_1932) ;
	assign x_4342 = (x_1929 & x_1930) ;
	assign x_4341 = (x_1927 & x_1928) ;
	assign x_4336 = (x_1924 & x_4335) ;
	assign x_4334 = (x_1922 & x_1923) ;
	assign x_4332 = (x_1919 & x_4331) ;
	assign x_4330 = (x_1917 & x_1918) ;
	assign x_4327 = (x_1914 & x_4326) ;
	assign x_4325 = (x_1912 & x_1913) ;
	assign x_4323 = (x_1910 & x_1911) ;
	assign x_4322 = (x_1908 & x_1909) ;
	assign x_4318 = (x_1905 & x_4317) ;
	assign x_4316 = (x_1903 & x_1904) ;
	assign x_4314 = (x_1900 & x_4313) ;
	assign x_4312 = (x_1898 & x_1899) ;
	assign x_4309 = (x_1895 & x_4308) ;
	assign x_4307 = (x_1893 & x_1894) ;
	assign x_4305 = (x_1891 & x_1892) ;
	assign x_4304 = (x_1889 & x_1890) ;
	assign x_4298 = (x_1886 & x_4297) ;
	assign x_4296 = (x_1884 & x_1885) ;
	assign x_4294 = (x_1881 & x_4293) ;
	assign x_4292 = (x_1879 & x_1880) ;
	assign x_4289 = (x_1876 & x_4288) ;
	assign x_4287 = (x_1874 & x_1875) ;
	assign x_4285 = (x_1872 & x_1873) ;
	assign x_4284 = (x_1870 & x_1871) ;
	assign x_4280 = (x_1867 & x_4279) ;
	assign x_4278 = (x_1865 & x_1866) ;
	assign x_4276 = (x_1862 & x_4275) ;
	assign x_4274 = (x_1860 & x_1861) ;
	assign x_4271 = (x_1857 & x_4270) ;
	assign x_4269 = (x_1855 & x_1856) ;
	assign x_4267 = (x_1853 & x_1854) ;
	assign x_4266 = (x_1851 & x_1852) ;
	assign x_4261 = (x_1848 & x_4260) ;
	assign x_4259 = (x_1846 & x_1847) ;
	assign x_4257 = (x_1843 & x_4256) ;
	assign x_4255 = (x_1841 & x_1842) ;
	assign x_4252 = (x_1838 & x_4251) ;
	assign x_4250 = (x_1836 & x_1837) ;
	assign x_4248 = (x_1834 & x_1835) ;
	assign x_4247 = (x_1832 & x_1833) ;
	assign x_4243 = (x_1829 & x_4242) ;
	assign x_4241 = (x_1827 & x_1828) ;
	assign x_4239 = (x_1825 & x_1826) ;
	assign x_4238 = (x_1823 & x_1824) ;
	assign x_4235 = (x_1820 & x_4234) ;
	assign x_4233 = (x_1818 & x_1819) ;
	assign x_4231 = (x_1816 & x_1817) ;
	assign x_4230 = (x_1814 & x_1815) ;
	assign x_4221 = (x_1811 & x_4220) ;
	assign x_4219 = (x_1809 & x_1810) ;
	assign x_4217 = (x_1806 & x_4216) ;
	assign x_4215 = (x_1804 & x_1805) ;
	assign x_4212 = (x_1801 & x_4211) ;
	assign x_4210 = (x_1799 & x_1800) ;
	assign x_4208 = (x_1797 & x_1798) ;
	assign x_4207 = (x_1795 & x_1796) ;
	assign x_4203 = (x_1792 & x_4202) ;
	assign x_4201 = (x_1790 & x_1791) ;
	assign x_4199 = (x_1787 & x_4198) ;
	assign x_4197 = (x_1785 & x_1786) ;
	assign x_4194 = (x_1782 & x_4193) ;
	assign x_4192 = (x_1780 & x_1781) ;
	assign x_4190 = (x_1778 & x_1779) ;
	assign x_4189 = (x_1776 & x_1777) ;
	assign x_4184 = (x_1773 & x_4183) ;
	assign x_4182 = (x_1771 & x_1772) ;
	assign x_4180 = (x_1768 & x_4179) ;
	assign x_4178 = (x_1766 & x_1767) ;
	assign x_4175 = (x_1763 & x_4174) ;
	assign x_4173 = (x_1761 & x_1762) ;
	assign x_4171 = (x_1759 & x_1760) ;
	assign x_4170 = (x_1757 & x_1758) ;
	assign x_4166 = (x_1754 & x_4165) ;
	assign x_4164 = (x_1752 & x_1753) ;
	assign x_4162 = (x_1749 & x_4161) ;
	assign x_4160 = (x_1747 & x_1748) ;
	assign x_4157 = (x_1744 & x_4156) ;
	assign x_4155 = (x_1742 & x_1743) ;
	assign x_4153 = (x_1740 & x_1741) ;
	assign x_4152 = (x_1738 & x_1739) ;
	assign x_4146 = (x_1735 & x_4145) ;
	assign x_4144 = (x_1733 & x_1734) ;
	assign x_4142 = (x_1730 & x_4141) ;
	assign x_4140 = (x_1728 & x_1729) ;
	assign x_4137 = (x_1725 & x_4136) ;
	assign x_4135 = (x_1723 & x_1724) ;
	assign x_4133 = (x_1721 & x_1722) ;
	assign x_4132 = (x_1719 & x_1720) ;
	assign x_4128 = (x_1716 & x_4127) ;
	assign x_4126 = (x_1714 & x_1715) ;
	assign x_4124 = (x_1711 & x_4123) ;
	assign x_4122 = (x_1709 & x_1710) ;
	assign x_4119 = (x_1706 & x_4118) ;
	assign x_4117 = (x_1704 & x_1705) ;
	assign x_4115 = (x_1702 & x_1703) ;
	assign x_4114 = (x_1700 & x_1701) ;
	assign x_4109 = (x_1697 & x_4108) ;
	assign x_4107 = (x_1695 & x_1696) ;
	assign x_4105 = (x_1692 & x_4104) ;
	assign x_4103 = (x_1690 & x_1691) ;
	assign x_4100 = (x_1687 & x_4099) ;
	assign x_4098 = (x_1685 & x_1686) ;
	assign x_4096 = (x_1683 & x_1684) ;
	assign x_4095 = (x_1681 & x_1682) ;
	assign x_4091 = (x_1678 & x_4090) ;
	assign x_4089 = (x_1676 & x_1677) ;
	assign x_4087 = (x_1674 & x_1675) ;
	assign x_4086 = (x_1672 & x_1673) ;
	assign x_4083 = (x_1669 & x_4082) ;
	assign x_4081 = (x_1667 & x_1668) ;
	assign x_4079 = (x_1665 & x_1666) ;
	assign x_4078 = (x_1663 & x_1664) ;
	assign x_4071 = (x_1660 & x_4070) ;
	assign x_4069 = (x_1658 & x_1659) ;
	assign x_4067 = (x_1655 & x_4066) ;
	assign x_4065 = (x_1653 & x_1654) ;
	assign x_4062 = (x_1650 & x_4061) ;
	assign x_4060 = (x_1648 & x_1649) ;
	assign x_4058 = (x_1646 & x_1647) ;
	assign x_4057 = (x_1644 & x_1645) ;
	assign x_4053 = (x_1641 & x_4052) ;
	assign x_4051 = (x_1639 & x_1640) ;
	assign x_4049 = (x_1636 & x_4048) ;
	assign x_4047 = (x_1634 & x_1635) ;
	assign x_4044 = (x_1631 & x_4043) ;
	assign x_4042 = (x_1629 & x_1630) ;
	assign x_4040 = (x_1627 & x_1628) ;
	assign x_4039 = (x_1625 & x_1626) ;
	assign x_4034 = (x_1622 & x_4033) ;
	assign x_4032 = (x_1620 & x_1621) ;
	assign x_4030 = (x_1617 & x_4029) ;
	assign x_4028 = (x_1615 & x_1616) ;
	assign x_4025 = (x_1612 & x_4024) ;
	assign x_4023 = (x_1610 & x_1611) ;
	assign x_4021 = (x_1608 & x_1609) ;
	assign x_4020 = (x_1606 & x_1607) ;
	assign x_4016 = (x_1603 & x_4015) ;
	assign x_4014 = (x_1601 & x_1602) ;
	assign x_4012 = (x_1598 & x_4011) ;
	assign x_4010 = (x_1596 & x_1597) ;
	assign x_4007 = (x_1593 & x_4006) ;
	assign x_4005 = (x_1591 & x_1592) ;
	assign x_4003 = (x_1589 & x_1590) ;
	assign x_4002 = (x_1587 & x_1588) ;
	assign x_3996 = (x_1584 & x_3995) ;
	assign x_3994 = (x_1582 & x_1583) ;
	assign x_3992 = (x_1579 & x_3991) ;
	assign x_3990 = (x_1577 & x_1578) ;
	assign x_3987 = (x_1574 & x_3986) ;
	assign x_3985 = (x_1572 & x_1573) ;
	assign x_3983 = (x_1570 & x_1571) ;
	assign x_3982 = (x_1568 & x_1569) ;
	assign x_3978 = (x_1565 & x_3977) ;
	assign x_3976 = (x_1563 & x_1564) ;
	assign x_3974 = (x_1560 & x_3973) ;
	assign x_3972 = (x_1558 & x_1559) ;
	assign x_3969 = (x_1555 & x_3968) ;
	assign x_3967 = (x_1553 & x_1554) ;
	assign x_3965 = (x_1551 & x_1552) ;
	assign x_3964 = (x_1549 & x_1550) ;
	assign x_3959 = (x_1546 & x_3958) ;
	assign x_3957 = (x_1544 & x_1545) ;
	assign x_3955 = (x_1541 & x_3954) ;
	assign x_3953 = (x_1539 & x_1540) ;
	assign x_3950 = (x_1536 & x_3949) ;
	assign x_3948 = (x_1534 & x_1535) ;
	assign x_3946 = (x_1532 & x_1533) ;
	assign x_3945 = (x_1530 & x_1531) ;
	assign x_3941 = (x_1527 & x_3940) ;
	assign x_3939 = (x_1525 & x_1526) ;
	assign x_3937 = (x_1523 & x_1524) ;
	assign x_3936 = (x_1521 & x_1522) ;
	assign x_3933 = (x_1518 & x_3932) ;
	assign x_3931 = (x_1516 & x_1517) ;
	assign x_3929 = (x_1514 & x_1515) ;
	assign x_3928 = (x_1512 & x_1513) ;
	assign x_3920 = (x_1509 & x_3919) ;
	assign x_3918 = (x_1507 & x_1508) ;
	assign x_3916 = (x_1504 & x_3915) ;
	assign x_3914 = (x_1502 & x_1503) ;
	assign x_3911 = (x_1499 & x_3910) ;
	assign x_3909 = (x_1497 & x_1498) ;
	assign x_3907 = (x_1495 & x_1496) ;
	assign x_3906 = (x_1493 & x_1494) ;
	assign x_3902 = (x_1490 & x_3901) ;
	assign x_3900 = (x_1488 & x_1489) ;
	assign x_3898 = (x_1485 & x_3897) ;
	assign x_3896 = (x_1483 & x_1484) ;
	assign x_3893 = (x_1480 & x_3892) ;
	assign x_3891 = (x_1478 & x_1479) ;
	assign x_3889 = (x_1476 & x_1477) ;
	assign x_3888 = (x_1474 & x_1475) ;
	assign x_3883 = (x_1471 & x_3882) ;
	assign x_3881 = (x_1469 & x_1470) ;
	assign x_3879 = (x_1466 & x_3878) ;
	assign x_3877 = (x_1464 & x_1465) ;
	assign x_3874 = (x_1461 & x_3873) ;
	assign x_3872 = (x_1459 & x_1460) ;
	assign x_3870 = (x_1457 & x_1458) ;
	assign x_3869 = (x_1455 & x_1456) ;
	assign x_3865 = (x_1452 & x_3864) ;
	assign x_3863 = (x_1450 & x_1451) ;
	assign x_3861 = (x_1447 & x_3860) ;
	assign x_3859 = (x_1445 & x_1446) ;
	assign x_3856 = (x_1442 & x_3855) ;
	assign x_3854 = (x_1440 & x_1441) ;
	assign x_3852 = (x_1438 & x_1439) ;
	assign x_3851 = (x_1436 & x_1437) ;
	assign x_3845 = (x_1433 & x_3844) ;
	assign x_3843 = (x_1431 & x_1432) ;
	assign x_3841 = (x_1428 & x_3840) ;
	assign x_3839 = (x_1426 & x_1427) ;
	assign x_3836 = (x_1423 & x_3835) ;
	assign x_3834 = (x_1421 & x_1422) ;
	assign x_3832 = (x_1419 & x_1420) ;
	assign x_3831 = (x_1417 & x_1418) ;
	assign x_3827 = (x_1414 & x_3826) ;
	assign x_3825 = (x_1412 & x_1413) ;
	assign x_3823 = (x_1409 & x_3822) ;
	assign x_3821 = (x_1407 & x_1408) ;
	assign x_3818 = (x_1404 & x_3817) ;
	assign x_3816 = (x_1402 & x_1403) ;
	assign x_3814 = (x_1400 & x_1401) ;
	assign x_3813 = (x_1398 & x_1399) ;
	assign x_3808 = (x_1395 & x_3807) ;
	assign x_3806 = (x_1393 & x_1394) ;
	assign x_3804 = (x_1390 & x_3803) ;
	assign x_3802 = (x_1388 & x_1389) ;
	assign x_3799 = (x_1385 & x_3798) ;
	assign x_3797 = (x_1383 & x_1384) ;
	assign x_3795 = (x_1381 & x_1382) ;
	assign x_3794 = (x_1379 & x_1380) ;
	assign x_3790 = (x_1376 & x_3789) ;
	assign x_3788 = (x_1374 & x_1375) ;
	assign x_3786 = (x_1372 & x_1373) ;
	assign x_3785 = (x_1370 & x_1371) ;
	assign x_3782 = (x_1367 & x_3781) ;
	assign x_3780 = (x_1365 & x_1366) ;
	assign x_3778 = (x_1363 & x_1364) ;
	assign x_3777 = (x_1361 & x_1362) ;
	assign x_3770 = (x_1358 & x_3769) ;
	assign x_3768 = (x_1356 & x_1357) ;
	assign x_3766 = (x_1353 & x_3765) ;
	assign x_3764 = (x_1351 & x_1352) ;
	assign x_3761 = (x_1348 & x_3760) ;
	assign x_3759 = (x_1346 & x_1347) ;
	assign x_3757 = (x_1344 & x_1345) ;
	assign x_3756 = (x_1342 & x_1343) ;
	assign x_3752 = (x_1339 & x_3751) ;
	assign x_3750 = (x_1337 & x_1338) ;
	assign x_3748 = (x_1334 & x_3747) ;
	assign x_3746 = (x_1332 & x_1333) ;
	assign x_3743 = (x_1329 & x_3742) ;
	assign x_3741 = (x_1327 & x_1328) ;
	assign x_3739 = (x_1325 & x_1326) ;
	assign x_3738 = (x_1323 & x_1324) ;
	assign x_3733 = (x_1320 & x_3732) ;
	assign x_3731 = (x_1318 & x_1319) ;
	assign x_3729 = (x_1315 & x_3728) ;
	assign x_3727 = (x_1313 & x_1314) ;
	assign x_3724 = (x_1310 & x_3723) ;
	assign x_3722 = (x_1308 & x_1309) ;
	assign x_3720 = (x_1306 & x_1307) ;
	assign x_3719 = (x_1304 & x_1305) ;
	assign x_3715 = (x_1301 & x_3714) ;
	assign x_3713 = (x_1299 & x_1300) ;
	assign x_3711 = (x_1296 & x_3710) ;
	assign x_3709 = (x_1294 & x_1295) ;
	assign x_3706 = (x_1291 & x_3705) ;
	assign x_3704 = (x_1289 & x_1290) ;
	assign x_3702 = (x_1287 & x_1288) ;
	assign x_3701 = (x_1285 & x_1286) ;
	assign x_3695 = (x_1282 & x_3694) ;
	assign x_3693 = (x_1280 & x_1281) ;
	assign x_3691 = (x_1277 & x_3690) ;
	assign x_3689 = (x_1275 & x_1276) ;
	assign x_3686 = (x_1272 & x_3685) ;
	assign x_3684 = (x_1270 & x_1271) ;
	assign x_3682 = (x_1268 & x_1269) ;
	assign x_3681 = (x_1266 & x_1267) ;
	assign x_3677 = (x_1263 & x_3676) ;
	assign x_3675 = (x_1261 & x_1262) ;
	assign x_3673 = (x_1258 & x_3672) ;
	assign x_3671 = (x_1256 & x_1257) ;
	assign x_3668 = (x_1253 & x_3667) ;
	assign x_3666 = (x_1251 & x_1252) ;
	assign x_3664 = (x_1249 & x_1250) ;
	assign x_3663 = (x_1247 & x_1248) ;
	assign x_3658 = (x_1244 & x_3657) ;
	assign x_3656 = (x_1242 & x_1243) ;
	assign x_3654 = (x_1239 & x_3653) ;
	assign x_3652 = (x_1237 & x_1238) ;
	assign x_3649 = (x_1234 & x_3648) ;
	assign x_3647 = (x_1232 & x_1233) ;
	assign x_3645 = (x_1230 & x_1231) ;
	assign x_3644 = (x_1228 & x_1229) ;
	assign x_3640 = (x_1225 & x_3639) ;
	assign x_3638 = (x_1223 & x_1224) ;
	assign x_3636 = (x_1221 & x_1222) ;
	assign x_3635 = (x_1219 & x_1220) ;
	assign x_3632 = (x_1216 & x_3631) ;
	assign x_3630 = (x_1214 & x_1215) ;
	assign x_3628 = (x_1212 & x_1213) ;
	assign x_3627 = (x_1210 & x_1211) ;
	assign x_3617 = (x_1207 & x_3616) ;
	assign x_3615 = (x_1205 & x_1206) ;
	assign x_3613 = (x_1202 & x_3612) ;
	assign x_3611 = (x_1200 & x_1201) ;
	assign x_3608 = (x_1197 & x_3607) ;
	assign x_3606 = (x_1195 & x_1196) ;
	assign x_3604 = (x_1193 & x_1194) ;
	assign x_3603 = (x_1191 & x_1192) ;
	assign x_3599 = (x_1188 & x_3598) ;
	assign x_3597 = (x_1186 & x_1187) ;
	assign x_3595 = (x_1183 & x_3594) ;
	assign x_3593 = (x_1181 & x_1182) ;
	assign x_3590 = (x_1178 & x_3589) ;
	assign x_3588 = (x_1176 & x_1177) ;
	assign x_3586 = (x_1174 & x_1175) ;
	assign x_3585 = (x_1172 & x_1173) ;
	assign x_3580 = (x_1169 & x_3579) ;
	assign x_3578 = (x_1167 & x_1168) ;
	assign x_3576 = (x_1164 & x_3575) ;
	assign x_3574 = (x_1162 & x_1163) ;
	assign x_3571 = (x_1159 & x_3570) ;
	assign x_3569 = (x_1157 & x_1158) ;
	assign x_3567 = (x_1155 & x_1156) ;
	assign x_3566 = (x_1153 & x_1154) ;
	assign x_3562 = (x_1150 & x_3561) ;
	assign x_3560 = (x_1148 & x_1149) ;
	assign x_3558 = (x_1145 & x_3557) ;
	assign x_3556 = (x_1143 & x_1144) ;
	assign x_3553 = (x_1140 & x_3552) ;
	assign x_3551 = (x_1138 & x_1139) ;
	assign x_3549 = (x_1136 & x_1137) ;
	assign x_3548 = (x_1134 & x_1135) ;
	assign x_3542 = (x_1131 & x_3541) ;
	assign x_3540 = (x_1129 & x_1130) ;
	assign x_3538 = (x_1126 & x_3537) ;
	assign x_3536 = (x_1124 & x_1125) ;
	assign x_3533 = (x_1121 & x_3532) ;
	assign x_3531 = (x_1119 & x_1120) ;
	assign x_3529 = (x_1117 & x_1118) ;
	assign x_3528 = (x_1115 & x_1116) ;
	assign x_3524 = (x_1112 & x_3523) ;
	assign x_3522 = (x_1110 & x_1111) ;
	assign x_3520 = (x_1107 & x_3519) ;
	assign x_3518 = (x_1105 & x_1106) ;
	assign x_3515 = (x_1102 & x_3514) ;
	assign x_3513 = (x_1100 & x_1101) ;
	assign x_3511 = (x_1098 & x_1099) ;
	assign x_3510 = (x_1096 & x_1097) ;
	assign x_3505 = (x_1093 & x_3504) ;
	assign x_3503 = (x_1091 & x_1092) ;
	assign x_3501 = (x_1088 & x_3500) ;
	assign x_3499 = (x_1086 & x_1087) ;
	assign x_3496 = (x_1083 & x_3495) ;
	assign x_3494 = (x_1081 & x_1082) ;
	assign x_3492 = (x_1079 & x_1080) ;
	assign x_3491 = (x_1077 & x_1078) ;
	assign x_3487 = (x_1074 & x_3486) ;
	assign x_3485 = (x_1072 & x_1073) ;
	assign x_3483 = (x_1069 & x_3482) ;
	assign x_3481 = (x_1067 & x_1068) ;
	assign x_3478 = (x_1064 & x_3477) ;
	assign x_3476 = (x_1062 & x_1063) ;
	assign x_3474 = (x_1060 & x_1061) ;
	assign x_3473 = (x_1058 & x_1059) ;
	assign x_3466 = (x_1055 & x_3465) ;
	assign x_3464 = (x_1053 & x_1054) ;
	assign x_3462 = (x_1050 & x_3461) ;
	assign x_3460 = (x_1048 & x_1049) ;
	assign x_3457 = (x_1045 & x_3456) ;
	assign x_3455 = (x_1043 & x_1044) ;
	assign x_3453 = (x_1041 & x_1042) ;
	assign x_3452 = (x_1039 & x_1040) ;
	assign x_3448 = (x_1036 & x_3447) ;
	assign x_3446 = (x_1034 & x_1035) ;
	assign x_3444 = (x_1031 & x_3443) ;
	assign x_3442 = (x_1029 & x_1030) ;
	assign x_3439 = (x_1026 & x_3438) ;
	assign x_3437 = (x_1024 & x_1025) ;
	assign x_3435 = (x_1022 & x_1023) ;
	assign x_3434 = (x_1020 & x_1021) ;
	assign x_3429 = (x_1017 & x_3428) ;
	assign x_3427 = (x_1015 & x_1016) ;
	assign x_3425 = (x_1012 & x_3424) ;
	assign x_3423 = (x_1010 & x_1011) ;
	assign x_3420 = (x_1007 & x_3419) ;
	assign x_3418 = (x_1005 & x_1006) ;
	assign x_3416 = (x_1003 & x_1004) ;
	assign x_3415 = (x_1001 & x_1002) ;
	assign x_3411 = (x_998 & x_3410) ;
	assign x_3409 = (x_996 & x_997) ;
	assign x_3407 = (x_993 & x_3406) ;
	assign x_3405 = (x_991 & x_992) ;
	assign x_3402 = (x_988 & x_3401) ;
	assign x_3400 = (x_986 & x_987) ;
	assign x_3398 = (x_984 & x_985) ;
	assign x_3397 = (x_982 & x_983) ;
	assign x_3391 = (x_979 & x_3390) ;
	assign x_3389 = (x_977 & x_978) ;
	assign x_3387 = (x_974 & x_3386) ;
	assign x_3385 = (x_972 & x_973) ;
	assign x_3382 = (x_969 & x_3381) ;
	assign x_3380 = (x_967 & x_968) ;
	assign x_3378 = (x_965 & x_966) ;
	assign x_3377 = (x_963 & x_964) ;
	assign x_3373 = (x_960 & x_3372) ;
	assign x_3371 = (x_958 & x_959) ;
	assign x_3369 = (x_955 & x_3368) ;
	assign x_3367 = (x_953 & x_954) ;
	assign x_3364 = (x_950 & x_3363) ;
	assign x_3362 = (x_948 & x_949) ;
	assign x_3360 = (x_946 & x_947) ;
	assign x_3359 = (x_944 & x_945) ;
	assign x_3354 = (x_941 & x_3353) ;
	assign x_3352 = (x_939 & x_940) ;
	assign x_3350 = (x_936 & x_3349) ;
	assign x_3348 = (x_934 & x_935) ;
	assign x_3345 = (x_931 & x_3344) ;
	assign x_3343 = (x_929 & x_930) ;
	assign x_3341 = (x_927 & x_928) ;
	assign x_3340 = (x_925 & x_926) ;
	assign x_3336 = (x_922 & x_3335) ;
	assign x_3334 = (x_920 & x_921) ;
	assign x_3332 = (x_918 & x_919) ;
	assign x_3331 = (x_916 & x_917) ;
	assign x_3328 = (x_913 & x_3327) ;
	assign x_3326 = (x_911 & x_912) ;
	assign x_3324 = (x_909 & x_910) ;
	assign x_3323 = (x_907 & x_908) ;
	assign x_3315 = (x_904 & x_3314) ;
	assign x_3313 = (x_902 & x_903) ;
	assign x_3311 = (x_899 & x_3310) ;
	assign x_3309 = (x_897 & x_898) ;
	assign x_3306 = (x_894 & x_3305) ;
	assign x_3304 = (x_892 & x_893) ;
	assign x_3302 = (x_890 & x_891) ;
	assign x_3301 = (x_888 & x_889) ;
	assign x_3297 = (x_885 & x_3296) ;
	assign x_3295 = (x_883 & x_884) ;
	assign x_3293 = (x_880 & x_3292) ;
	assign x_3291 = (x_878 & x_879) ;
	assign x_3288 = (x_875 & x_3287) ;
	assign x_3286 = (x_873 & x_874) ;
	assign x_3284 = (x_871 & x_872) ;
	assign x_3283 = (x_869 & x_870) ;
	assign x_3278 = (x_866 & x_3277) ;
	assign x_3276 = (x_864 & x_865) ;
	assign x_3274 = (x_861 & x_3273) ;
	assign x_3272 = (x_859 & x_860) ;
	assign x_3269 = (x_856 & x_3268) ;
	assign x_3267 = (x_854 & x_855) ;
	assign x_3265 = (x_852 & x_853) ;
	assign x_3264 = (x_850 & x_851) ;
	assign x_3260 = (x_847 & x_3259) ;
	assign x_3258 = (x_845 & x_846) ;
	assign x_3256 = (x_842 & x_3255) ;
	assign x_3254 = (x_840 & x_841) ;
	assign x_3251 = (x_837 & x_3250) ;
	assign x_3249 = (x_835 & x_836) ;
	assign x_3247 = (x_833 & x_834) ;
	assign x_3246 = (x_831 & x_832) ;
	assign x_3240 = (x_828 & x_3239) ;
	assign x_3238 = (x_826 & x_827) ;
	assign x_3236 = (x_823 & x_3235) ;
	assign x_3234 = (x_821 & x_822) ;
	assign x_3231 = (x_818 & x_3230) ;
	assign x_3229 = (x_816 & x_817) ;
	assign x_3227 = (x_814 & x_815) ;
	assign x_3226 = (x_812 & x_813) ;
	assign x_3222 = (x_809 & x_3221) ;
	assign x_3220 = (x_807 & x_808) ;
	assign x_3218 = (x_804 & x_3217) ;
	assign x_3216 = (x_802 & x_803) ;
	assign x_3213 = (x_799 & x_3212) ;
	assign x_3211 = (x_797 & x_798) ;
	assign x_3209 = (x_795 & x_796) ;
	assign x_3208 = (x_793 & x_794) ;
	assign x_3203 = (x_790 & x_3202) ;
	assign x_3201 = (x_788 & x_789) ;
	assign x_3199 = (x_785 & x_3198) ;
	assign x_3197 = (x_783 & x_784) ;
	assign x_3194 = (x_780 & x_3193) ;
	assign x_3192 = (x_778 & x_779) ;
	assign x_3190 = (x_776 & x_777) ;
	assign x_3189 = (x_774 & x_775) ;
	assign x_3185 = (x_771 & x_3184) ;
	assign x_3183 = (x_769 & x_770) ;
	assign x_3181 = (x_767 & x_768) ;
	assign x_3180 = (x_765 & x_766) ;
	assign x_3177 = (x_762 & x_3176) ;
	assign x_3175 = (x_760 & x_761) ;
	assign x_3173 = (x_758 & x_759) ;
	assign x_3172 = (x_756 & x_757) ;
	assign x_3165 = (x_753 & x_3164) ;
	assign x_3163 = (x_751 & x_752) ;
	assign x_3161 = (x_748 & x_3160) ;
	assign x_3159 = (x_746 & x_747) ;
	assign x_3156 = (x_743 & x_3155) ;
	assign x_3154 = (x_741 & x_742) ;
	assign x_3152 = (x_739 & x_740) ;
	assign x_3151 = (x_737 & x_738) ;
	assign x_3147 = (x_734 & x_3146) ;
	assign x_3145 = (x_732 & x_733) ;
	assign x_3143 = (x_729 & x_3142) ;
	assign x_3141 = (x_727 & x_728) ;
	assign x_3138 = (x_724 & x_3137) ;
	assign x_3136 = (x_722 & x_723) ;
	assign x_3134 = (x_720 & x_721) ;
	assign x_3133 = (x_718 & x_719) ;
	assign x_3128 = (x_715 & x_3127) ;
	assign x_3126 = (x_713 & x_714) ;
	assign x_3124 = (x_710 & x_3123) ;
	assign x_3122 = (x_708 & x_709) ;
	assign x_3119 = (x_705 & x_3118) ;
	assign x_3117 = (x_703 & x_704) ;
	assign x_3115 = (x_701 & x_702) ;
	assign x_3114 = (x_699 & x_700) ;
	assign x_3110 = (x_696 & x_3109) ;
	assign x_3108 = (x_694 & x_695) ;
	assign x_3106 = (x_691 & x_3105) ;
	assign x_3104 = (x_689 & x_690) ;
	assign x_3101 = (x_686 & x_3100) ;
	assign x_3099 = (x_684 & x_685) ;
	assign x_3097 = (x_682 & x_683) ;
	assign x_3096 = (x_680 & x_681) ;
	assign x_3090 = (x_677 & x_3089) ;
	assign x_3088 = (x_675 & x_676) ;
	assign x_3086 = (x_672 & x_3085) ;
	assign x_3084 = (x_670 & x_671) ;
	assign x_3081 = (x_667 & x_3080) ;
	assign x_3079 = (x_665 & x_666) ;
	assign x_3077 = (x_663 & x_664) ;
	assign x_3076 = (x_661 & x_662) ;
	assign x_3072 = (x_658 & x_3071) ;
	assign x_3070 = (x_656 & x_657) ;
	assign x_3068 = (x_653 & x_3067) ;
	assign x_3066 = (x_651 & x_652) ;
	assign x_3063 = (x_648 & x_3062) ;
	assign x_3061 = (x_646 & x_647) ;
	assign x_3059 = (x_644 & x_645) ;
	assign x_3058 = (x_642 & x_643) ;
	assign x_3053 = (x_639 & x_3052) ;
	assign x_3051 = (x_637 & x_638) ;
	assign x_3049 = (x_634 & x_3048) ;
	assign x_3047 = (x_632 & x_633) ;
	assign x_3044 = (x_629 & x_3043) ;
	assign x_3042 = (x_627 & x_628) ;
	assign x_3040 = (x_625 & x_626) ;
	assign x_3039 = (x_623 & x_624) ;
	assign x_3035 = (x_620 & x_3034) ;
	assign x_3033 = (x_618 & x_619) ;
	assign x_3031 = (x_616 & x_617) ;
	assign x_3030 = (x_614 & x_615) ;
	assign x_3027 = (x_611 & x_3026) ;
	assign x_3025 = (x_609 & x_610) ;
	assign x_3023 = (x_607 & x_608) ;
	assign x_3022 = (x_605 & x_606) ;
	assign x_3013 = (x_602 & x_3012) ;
	assign x_3011 = (x_600 & x_601) ;
	assign x_3009 = (x_597 & x_3008) ;
	assign x_3007 = (x_595 & x_596) ;
	assign x_3004 = (x_592 & x_3003) ;
	assign x_3002 = (x_590 & x_591) ;
	assign x_3000 = (x_588 & x_589) ;
	assign x_2999 = (x_586 & x_587) ;
	assign x_2995 = (x_583 & x_2994) ;
	assign x_2993 = (x_581 & x_582) ;
	assign x_2991 = (x_578 & x_2990) ;
	assign x_2989 = (x_576 & x_577) ;
	assign x_2986 = (x_573 & x_2985) ;
	assign x_2984 = (x_571 & x_572) ;
	assign x_2982 = (x_569 & x_570) ;
	assign x_2981 = (x_567 & x_568) ;
	assign x_2976 = (x_564 & x_2975) ;
	assign x_2974 = (x_562 & x_563) ;
	assign x_2972 = (x_559 & x_2971) ;
	assign x_2970 = (x_557 & x_558) ;
	assign x_2967 = (x_554 & x_2966) ;
	assign x_2965 = (x_552 & x_553) ;
	assign x_2963 = (x_550 & x_551) ;
	assign x_2962 = (x_548 & x_549) ;
	assign x_2958 = (x_545 & x_2957) ;
	assign x_2956 = (x_543 & x_544) ;
	assign x_2954 = (x_540 & x_2953) ;
	assign x_2952 = (x_538 & x_539) ;
	assign x_2949 = (x_535 & x_2948) ;
	assign x_2947 = (x_533 & x_534) ;
	assign x_2945 = (x_531 & x_532) ;
	assign x_2944 = (x_529 & x_530) ;
	assign x_2938 = (x_526 & x_2937) ;
	assign x_2936 = (x_524 & x_525) ;
	assign x_2934 = (x_521 & x_2933) ;
	assign x_2932 = (x_519 & x_520) ;
	assign x_2929 = (x_516 & x_2928) ;
	assign x_2927 = (x_514 & x_515) ;
	assign x_2925 = (x_512 & x_513) ;
	assign x_2924 = (x_510 & x_511) ;
	assign x_2920 = (x_507 & x_2919) ;
	assign x_2918 = (x_505 & x_506) ;
	assign x_2916 = (x_502 & x_2915) ;
	assign x_2914 = (x_500 & x_501) ;
	assign x_2911 = (x_497 & x_2910) ;
	assign x_2909 = (x_495 & x_496) ;
	assign x_2907 = (x_493 & x_494) ;
	assign x_2906 = (x_491 & x_492) ;
	assign x_2901 = (x_488 & x_2900) ;
	assign x_2899 = (x_486 & x_487) ;
	assign x_2897 = (x_483 & x_2896) ;
	assign x_2895 = (x_481 & x_482) ;
	assign x_2892 = (x_478 & x_2891) ;
	assign x_2890 = (x_476 & x_477) ;
	assign x_2888 = (x_474 & x_475) ;
	assign x_2887 = (x_472 & x_473) ;
	assign x_2883 = (x_469 & x_2882) ;
	assign x_2881 = (x_467 & x_468) ;
	assign x_2879 = (x_465 & x_466) ;
	assign x_2878 = (x_463 & x_464) ;
	assign x_2875 = (x_460 & x_2874) ;
	assign x_2873 = (x_458 & x_459) ;
	assign x_2871 = (x_456 & x_457) ;
	assign x_2870 = (x_454 & x_455) ;
	assign x_2863 = (x_451 & x_2862) ;
	assign x_2861 = (x_449 & x_450) ;
	assign x_2859 = (x_446 & x_2858) ;
	assign x_2857 = (x_444 & x_445) ;
	assign x_2854 = (x_441 & x_2853) ;
	assign x_2852 = (x_439 & x_440) ;
	assign x_2850 = (x_437 & x_438) ;
	assign x_2849 = (x_435 & x_436) ;
	assign x_2845 = (x_432 & x_2844) ;
	assign x_2843 = (x_430 & x_431) ;
	assign x_2841 = (x_427 & x_2840) ;
	assign x_2839 = (x_425 & x_426) ;
	assign x_2836 = (x_422 & x_2835) ;
	assign x_2834 = (x_420 & x_421) ;
	assign x_2832 = (x_418 & x_419) ;
	assign x_2831 = (x_416 & x_417) ;
	assign x_2826 = (x_413 & x_2825) ;
	assign x_2824 = (x_411 & x_412) ;
	assign x_2822 = (x_408 & x_2821) ;
	assign x_2820 = (x_406 & x_407) ;
	assign x_2817 = (x_403 & x_2816) ;
	assign x_2815 = (x_401 & x_402) ;
	assign x_2813 = (x_399 & x_400) ;
	assign x_2812 = (x_397 & x_398) ;
	assign x_2808 = (x_394 & x_2807) ;
	assign x_2806 = (x_392 & x_393) ;
	assign x_2804 = (x_389 & x_2803) ;
	assign x_2802 = (x_387 & x_388) ;
	assign x_2799 = (x_384 & x_2798) ;
	assign x_2797 = (x_382 & x_383) ;
	assign x_2795 = (x_380 & x_381) ;
	assign x_2794 = (x_378 & x_379) ;
	assign x_2788 = (x_375 & x_2787) ;
	assign x_2786 = (x_373 & x_374) ;
	assign x_2784 = (x_370 & x_2783) ;
	assign x_2782 = (x_368 & x_369) ;
	assign x_2779 = (x_365 & x_2778) ;
	assign x_2777 = (x_363 & x_364) ;
	assign x_2775 = (x_361 & x_362) ;
	assign x_2774 = (x_359 & x_360) ;
	assign x_2770 = (x_356 & x_2769) ;
	assign x_2768 = (x_354 & x_355) ;
	assign x_2766 = (x_351 & x_2765) ;
	assign x_2764 = (x_349 & x_350) ;
	assign x_2761 = (x_346 & x_2760) ;
	assign x_2759 = (x_344 & x_345) ;
	assign x_2757 = (x_342 & x_343) ;
	assign x_2756 = (x_340 & x_341) ;
	assign x_2751 = (x_337 & x_2750) ;
	assign x_2749 = (x_335 & x_336) ;
	assign x_2747 = (x_332 & x_2746) ;
	assign x_2745 = (x_330 & x_331) ;
	assign x_2742 = (x_327 & x_2741) ;
	assign x_2740 = (x_325 & x_326) ;
	assign x_2738 = (x_323 & x_324) ;
	assign x_2737 = (x_321 & x_322) ;
	assign x_2733 = (x_318 & x_2732) ;
	assign x_2731 = (x_316 & x_317) ;
	assign x_2729 = (x_314 & x_315) ;
	assign x_2728 = (x_312 & x_313) ;
	assign x_2725 = (x_309 & x_2724) ;
	assign x_2723 = (x_307 & x_308) ;
	assign x_2721 = (x_305 & x_306) ;
	assign x_2720 = (x_303 & x_304) ;
	assign x_2712 = (x_300 & x_2711) ;
	assign x_2710 = (x_298 & x_299) ;
	assign x_2708 = (x_295 & x_2707) ;
	assign x_2706 = (x_293 & x_294) ;
	assign x_2703 = (x_290 & x_2702) ;
	assign x_2701 = (x_288 & x_289) ;
	assign x_2699 = (x_286 & x_287) ;
	assign x_2698 = (x_284 & x_285) ;
	assign x_2694 = (x_281 & x_2693) ;
	assign x_2692 = (x_279 & x_280) ;
	assign x_2690 = (x_276 & x_2689) ;
	assign x_2688 = (x_274 & x_275) ;
	assign x_2685 = (x_271 & x_2684) ;
	assign x_2683 = (x_269 & x_270) ;
	assign x_2681 = (x_267 & x_268) ;
	assign x_2680 = (x_265 & x_266) ;
	assign x_2675 = (x_262 & x_2674) ;
	assign x_2673 = (x_260 & x_261) ;
	assign x_2671 = (x_257 & x_2670) ;
	assign x_2669 = (x_255 & x_256) ;
	assign x_2666 = (x_252 & x_2665) ;
	assign x_2664 = (x_250 & x_251) ;
	assign x_2662 = (x_248 & x_249) ;
	assign x_2661 = (x_246 & x_247) ;
	assign x_2657 = (x_243 & x_2656) ;
	assign x_2655 = (x_241 & x_242) ;
	assign x_2653 = (x_238 & x_2652) ;
	assign x_2651 = (x_236 & x_237) ;
	assign x_2648 = (x_233 & x_2647) ;
	assign x_2646 = (x_231 & x_232) ;
	assign x_2644 = (x_229 & x_230) ;
	assign x_2643 = (x_227 & x_228) ;
	assign x_2637 = (x_224 & x_2636) ;
	assign x_2635 = (x_222 & x_223) ;
	assign x_2633 = (x_219 & x_2632) ;
	assign x_2631 = (x_217 & x_218) ;
	assign x_2628 = (x_214 & x_2627) ;
	assign x_2626 = (x_212 & x_213) ;
	assign x_2624 = (x_210 & x_211) ;
	assign x_2623 = (x_208 & x_209) ;
	assign x_2619 = (x_205 & x_2618) ;
	assign x_2617 = (x_203 & x_204) ;
	assign x_2615 = (x_200 & x_2614) ;
	assign x_2613 = (x_198 & x_199) ;
	assign x_2610 = (x_195 & x_2609) ;
	assign x_2608 = (x_193 & x_194) ;
	assign x_2606 = (x_191 & x_192) ;
	assign x_2605 = (x_189 & x_190) ;
	assign x_2600 = (x_186 & x_2599) ;
	assign x_2598 = (x_184 & x_185) ;
	assign x_2596 = (x_181 & x_2595) ;
	assign x_2594 = (x_179 & x_180) ;
	assign x_2591 = (x_176 & x_2590) ;
	assign x_2589 = (x_174 & x_175) ;
	assign x_2587 = (x_172 & x_173) ;
	assign x_2586 = (x_170 & x_171) ;
	assign x_2582 = (x_167 & x_2581) ;
	assign x_2580 = (x_165 & x_166) ;
	assign x_2578 = (x_163 & x_164) ;
	assign x_2577 = (x_161 & x_162) ;
	assign x_2574 = (x_158 & x_2573) ;
	assign x_2572 = (x_156 & x_157) ;
	assign x_2570 = (x_154 & x_155) ;
	assign x_2569 = (x_152 & x_153) ;
	assign x_2562 = (x_149 & x_2561) ;
	assign x_2560 = (x_147 & x_148) ;
	assign x_2558 = (x_144 & x_2557) ;
	assign x_2556 = (x_142 & x_143) ;
	assign x_2553 = (x_139 & x_2552) ;
	assign x_2551 = (x_137 & x_138) ;
	assign x_2549 = (x_135 & x_136) ;
	assign x_2548 = (x_133 & x_134) ;
	assign x_2544 = (x_130 & x_2543) ;
	assign x_2542 = (x_128 & x_129) ;
	assign x_2540 = (x_125 & x_2539) ;
	assign x_2538 = (x_123 & x_124) ;
	assign x_2535 = (x_120 & x_2534) ;
	assign x_2533 = (x_118 & x_119) ;
	assign x_2531 = (x_116 & x_117) ;
	assign x_2530 = (x_114 & x_115) ;
	assign x_2525 = (x_111 & x_2524) ;
	assign x_2523 = (x_109 & x_110) ;
	assign x_2521 = (x_106 & x_2520) ;
	assign x_2519 = (x_104 & x_105) ;
	assign x_2516 = (x_101 & x_2515) ;
	assign x_2514 = (x_99 & x_100) ;
	assign x_2512 = (x_97 & x_98) ;
	assign x_2511 = (x_95 & x_96) ;
	assign x_2507 = (x_92 & x_2506) ;
	assign x_2505 = (x_90 & x_91) ;
	assign x_2503 = (x_87 & x_2502) ;
	assign x_2501 = (x_85 & x_86) ;
	assign x_2498 = (x_82 & x_2497) ;
	assign x_2496 = (x_80 & x_81) ;
	assign x_2494 = (x_78 & x_79) ;
	assign x_2493 = (x_76 & x_77) ;
	assign x_2487 = (x_73 & x_2486) ;
	assign x_2485 = (x_71 & x_72) ;
	assign x_2483 = (x_68 & x_2482) ;
	assign x_2481 = (x_66 & x_67) ;
	assign x_2478 = (x_63 & x_2477) ;
	assign x_2476 = (x_61 & x_62) ;
	assign x_2474 = (x_59 & x_60) ;
	assign x_2473 = (x_57 & x_58) ;
	assign x_2469 = (x_54 & x_2468) ;
	assign x_2467 = (x_52 & x_53) ;
	assign x_2465 = (x_49 & x_2464) ;
	assign x_2463 = (x_47 & x_48) ;
	assign x_2460 = (x_44 & x_2459) ;
	assign x_2458 = (x_42 & x_43) ;
	assign x_2456 = (x_40 & x_41) ;
	assign x_2455 = (x_38 & x_39) ;
	assign x_2450 = (x_35 & x_2449) ;
	assign x_2448 = (x_33 & x_34) ;
	assign x_2446 = (x_30 & x_2445) ;
	assign x_2444 = (x_28 & x_29) ;
	assign x_2441 = (x_25 & x_2440) ;
	assign x_2439 = (x_23 & x_24) ;
	assign x_2437 = (x_21 & x_22) ;
	assign x_2436 = (x_19 & x_20) ;
	assign x_2432 = (x_16 & x_2431) ;
	assign x_2430 = (x_14 & x_15) ;
	assign x_2428 = (x_12 & x_13) ;
	assign x_2427 = (x_10 & x_11) ;
	assign x_2424 = (x_7 & x_2423) ;
	assign x_2422 = (x_5 & x_6) ;
	assign x_2420 = (x_3 & x_4) ;
	assign x_2419 = (x_1 & x_2) ;
	assign x_4826 = (x_4823 & x_4825) ;
	assign x_4822 = (x_4819 & x_4821) ;
	assign x_4817 = (x_4814 & x_4816) ;
	assign x_4813 = (x_4811 & x_4812) ;
	assign x_4808 = (x_4805 & x_4807) ;
	assign x_4804 = (x_4801 & x_4803) ;
	assign x_4799 = (x_4796 & x_4798) ;
	assign x_4795 = (x_4793 & x_4794) ;
	assign x_4789 = (x_4786 & x_4788) ;
	assign x_4785 = (x_4782 & x_4784) ;
	assign x_4780 = (x_4777 & x_4779) ;
	assign x_4776 = (x_4774 & x_4775) ;
	assign x_4771 = (x_4768 & x_4770) ;
	assign x_4767 = (x_4764 & x_4766) ;
	assign x_4762 = (x_4759 & x_4761) ;
	assign x_4758 = (x_4756 & x_4757) ;
	assign x_4751 = (x_4748 & x_4750) ;
	assign x_4747 = (x_4744 & x_4746) ;
	assign x_4742 = (x_4739 & x_4741) ;
	assign x_4738 = (x_4736 & x_4737) ;
	assign x_4733 = (x_4730 & x_4732) ;
	assign x_4729 = (x_4726 & x_4728) ;
	assign x_4724 = (x_4721 & x_4723) ;
	assign x_4720 = (x_4718 & x_4719) ;
	assign x_4714 = (x_4711 & x_4713) ;
	assign x_4710 = (x_4707 & x_4709) ;
	assign x_4705 = (x_4702 & x_4704) ;
	assign x_4701 = (x_4699 & x_4700) ;
	assign x_4696 = (x_4693 & x_4695) ;
	assign x_4692 = (x_4689 & x_4691) ;
	assign x_4687 = (x_4684 & x_4686) ;
	assign x_4683 = (x_4681 & x_4682) ;
	assign x_4675 = (x_4672 & x_4674) ;
	assign x_4671 = (x_4668 & x_4670) ;
	assign x_4666 = (x_4663 & x_4665) ;
	assign x_4662 = (x_4660 & x_4661) ;
	assign x_4657 = (x_4654 & x_4656) ;
	assign x_4653 = (x_4650 & x_4652) ;
	assign x_4648 = (x_4645 & x_4647) ;
	assign x_4644 = (x_4642 & x_4643) ;
	assign x_4638 = (x_4635 & x_4637) ;
	assign x_4634 = (x_4631 & x_4633) ;
	assign x_4629 = (x_4626 & x_4628) ;
	assign x_4625 = (x_4623 & x_4624) ;
	assign x_4620 = (x_4617 & x_4619) ;
	assign x_4616 = (x_4613 & x_4615) ;
	assign x_4611 = (x_4608 & x_4610) ;
	assign x_4607 = (x_4605 & x_4606) ;
	assign x_4600 = (x_4597 & x_4599) ;
	assign x_4596 = (x_4593 & x_4595) ;
	assign x_4591 = (x_4588 & x_4590) ;
	assign x_4587 = (x_4585 & x_4586) ;
	assign x_4582 = (x_4579 & x_4581) ;
	assign x_4578 = (x_4575 & x_4577) ;
	assign x_4573 = (x_4570 & x_4572) ;
	assign x_4569 = (x_4567 & x_4568) ;
	assign x_4563 = (x_4560 & x_4562) ;
	assign x_4559 = (x_4556 & x_4558) ;
	assign x_4554 = (x_4551 & x_4553) ;
	assign x_4550 = (x_4548 & x_4549) ;
	assign x_4545 = (x_4542 & x_4544) ;
	assign x_4541 = (x_4539 & x_4540) ;
	assign x_4537 = (x_4534 & x_4536) ;
	assign x_4533 = (x_4531 & x_4532) ;
	assign x_4524 = (x_4521 & x_4523) ;
	assign x_4520 = (x_4517 & x_4519) ;
	assign x_4515 = (x_4512 & x_4514) ;
	assign x_4511 = (x_4509 & x_4510) ;
	assign x_4506 = (x_4503 & x_4505) ;
	assign x_4502 = (x_4499 & x_4501) ;
	assign x_4497 = (x_4494 & x_4496) ;
	assign x_4493 = (x_4491 & x_4492) ;
	assign x_4487 = (x_4484 & x_4486) ;
	assign x_4483 = (x_4480 & x_4482) ;
	assign x_4478 = (x_4475 & x_4477) ;
	assign x_4474 = (x_4472 & x_4473) ;
	assign x_4469 = (x_4466 & x_4468) ;
	assign x_4465 = (x_4462 & x_4464) ;
	assign x_4460 = (x_4457 & x_4459) ;
	assign x_4456 = (x_4454 & x_4455) ;
	assign x_4449 = (x_4446 & x_4448) ;
	assign x_4445 = (x_4442 & x_4444) ;
	assign x_4440 = (x_4437 & x_4439) ;
	assign x_4436 = (x_4434 & x_4435) ;
	assign x_4431 = (x_4428 & x_4430) ;
	assign x_4427 = (x_4424 & x_4426) ;
	assign x_4422 = (x_4419 & x_4421) ;
	assign x_4418 = (x_4416 & x_4417) ;
	assign x_4412 = (x_4409 & x_4411) ;
	assign x_4408 = (x_4405 & x_4407) ;
	assign x_4403 = (x_4400 & x_4402) ;
	assign x_4399 = (x_4397 & x_4398) ;
	assign x_4394 = (x_4391 & x_4393) ;
	assign x_4390 = (x_4388 & x_4389) ;
	assign x_4386 = (x_4383 & x_4385) ;
	assign x_4382 = (x_4380 & x_4381) ;
	assign x_4374 = (x_4371 & x_4373) ;
	assign x_4370 = (x_4367 & x_4369) ;
	assign x_4365 = (x_4362 & x_4364) ;
	assign x_4361 = (x_4359 & x_4360) ;
	assign x_4356 = (x_4353 & x_4355) ;
	assign x_4352 = (x_4349 & x_4351) ;
	assign x_4347 = (x_4344 & x_4346) ;
	assign x_4343 = (x_4341 & x_4342) ;
	assign x_4337 = (x_4334 & x_4336) ;
	assign x_4333 = (x_4330 & x_4332) ;
	assign x_4328 = (x_4325 & x_4327) ;
	assign x_4324 = (x_4322 & x_4323) ;
	assign x_4319 = (x_4316 & x_4318) ;
	assign x_4315 = (x_4312 & x_4314) ;
	assign x_4310 = (x_4307 & x_4309) ;
	assign x_4306 = (x_4304 & x_4305) ;
	assign x_4299 = (x_4296 & x_4298) ;
	assign x_4295 = (x_4292 & x_4294) ;
	assign x_4290 = (x_4287 & x_4289) ;
	assign x_4286 = (x_4284 & x_4285) ;
	assign x_4281 = (x_4278 & x_4280) ;
	assign x_4277 = (x_4274 & x_4276) ;
	assign x_4272 = (x_4269 & x_4271) ;
	assign x_4268 = (x_4266 & x_4267) ;
	assign x_4262 = (x_4259 & x_4261) ;
	assign x_4258 = (x_4255 & x_4257) ;
	assign x_4253 = (x_4250 & x_4252) ;
	assign x_4249 = (x_4247 & x_4248) ;
	assign x_4244 = (x_4241 & x_4243) ;
	assign x_4240 = (x_4238 & x_4239) ;
	assign x_4236 = (x_4233 & x_4235) ;
	assign x_4232 = (x_4230 & x_4231) ;
	assign x_4222 = (x_4219 & x_4221) ;
	assign x_4218 = (x_4215 & x_4217) ;
	assign x_4213 = (x_4210 & x_4212) ;
	assign x_4209 = (x_4207 & x_4208) ;
	assign x_4204 = (x_4201 & x_4203) ;
	assign x_4200 = (x_4197 & x_4199) ;
	assign x_4195 = (x_4192 & x_4194) ;
	assign x_4191 = (x_4189 & x_4190) ;
	assign x_4185 = (x_4182 & x_4184) ;
	assign x_4181 = (x_4178 & x_4180) ;
	assign x_4176 = (x_4173 & x_4175) ;
	assign x_4172 = (x_4170 & x_4171) ;
	assign x_4167 = (x_4164 & x_4166) ;
	assign x_4163 = (x_4160 & x_4162) ;
	assign x_4158 = (x_4155 & x_4157) ;
	assign x_4154 = (x_4152 & x_4153) ;
	assign x_4147 = (x_4144 & x_4146) ;
	assign x_4143 = (x_4140 & x_4142) ;
	assign x_4138 = (x_4135 & x_4137) ;
	assign x_4134 = (x_4132 & x_4133) ;
	assign x_4129 = (x_4126 & x_4128) ;
	assign x_4125 = (x_4122 & x_4124) ;
	assign x_4120 = (x_4117 & x_4119) ;
	assign x_4116 = (x_4114 & x_4115) ;
	assign x_4110 = (x_4107 & x_4109) ;
	assign x_4106 = (x_4103 & x_4105) ;
	assign x_4101 = (x_4098 & x_4100) ;
	assign x_4097 = (x_4095 & x_4096) ;
	assign x_4092 = (x_4089 & x_4091) ;
	assign x_4088 = (x_4086 & x_4087) ;
	assign x_4084 = (x_4081 & x_4083) ;
	assign x_4080 = (x_4078 & x_4079) ;
	assign x_4072 = (x_4069 & x_4071) ;
	assign x_4068 = (x_4065 & x_4067) ;
	assign x_4063 = (x_4060 & x_4062) ;
	assign x_4059 = (x_4057 & x_4058) ;
	assign x_4054 = (x_4051 & x_4053) ;
	assign x_4050 = (x_4047 & x_4049) ;
	assign x_4045 = (x_4042 & x_4044) ;
	assign x_4041 = (x_4039 & x_4040) ;
	assign x_4035 = (x_4032 & x_4034) ;
	assign x_4031 = (x_4028 & x_4030) ;
	assign x_4026 = (x_4023 & x_4025) ;
	assign x_4022 = (x_4020 & x_4021) ;
	assign x_4017 = (x_4014 & x_4016) ;
	assign x_4013 = (x_4010 & x_4012) ;
	assign x_4008 = (x_4005 & x_4007) ;
	assign x_4004 = (x_4002 & x_4003) ;
	assign x_3997 = (x_3994 & x_3996) ;
	assign x_3993 = (x_3990 & x_3992) ;
	assign x_3988 = (x_3985 & x_3987) ;
	assign x_3984 = (x_3982 & x_3983) ;
	assign x_3979 = (x_3976 & x_3978) ;
	assign x_3975 = (x_3972 & x_3974) ;
	assign x_3970 = (x_3967 & x_3969) ;
	assign x_3966 = (x_3964 & x_3965) ;
	assign x_3960 = (x_3957 & x_3959) ;
	assign x_3956 = (x_3953 & x_3955) ;
	assign x_3951 = (x_3948 & x_3950) ;
	assign x_3947 = (x_3945 & x_3946) ;
	assign x_3942 = (x_3939 & x_3941) ;
	assign x_3938 = (x_3936 & x_3937) ;
	assign x_3934 = (x_3931 & x_3933) ;
	assign x_3930 = (x_3928 & x_3929) ;
	assign x_3921 = (x_3918 & x_3920) ;
	assign x_3917 = (x_3914 & x_3916) ;
	assign x_3912 = (x_3909 & x_3911) ;
	assign x_3908 = (x_3906 & x_3907) ;
	assign x_3903 = (x_3900 & x_3902) ;
	assign x_3899 = (x_3896 & x_3898) ;
	assign x_3894 = (x_3891 & x_3893) ;
	assign x_3890 = (x_3888 & x_3889) ;
	assign x_3884 = (x_3881 & x_3883) ;
	assign x_3880 = (x_3877 & x_3879) ;
	assign x_3875 = (x_3872 & x_3874) ;
	assign x_3871 = (x_3869 & x_3870) ;
	assign x_3866 = (x_3863 & x_3865) ;
	assign x_3862 = (x_3859 & x_3861) ;
	assign x_3857 = (x_3854 & x_3856) ;
	assign x_3853 = (x_3851 & x_3852) ;
	assign x_3846 = (x_3843 & x_3845) ;
	assign x_3842 = (x_3839 & x_3841) ;
	assign x_3837 = (x_3834 & x_3836) ;
	assign x_3833 = (x_3831 & x_3832) ;
	assign x_3828 = (x_3825 & x_3827) ;
	assign x_3824 = (x_3821 & x_3823) ;
	assign x_3819 = (x_3816 & x_3818) ;
	assign x_3815 = (x_3813 & x_3814) ;
	assign x_3809 = (x_3806 & x_3808) ;
	assign x_3805 = (x_3802 & x_3804) ;
	assign x_3800 = (x_3797 & x_3799) ;
	assign x_3796 = (x_3794 & x_3795) ;
	assign x_3791 = (x_3788 & x_3790) ;
	assign x_3787 = (x_3785 & x_3786) ;
	assign x_3783 = (x_3780 & x_3782) ;
	assign x_3779 = (x_3777 & x_3778) ;
	assign x_3771 = (x_3768 & x_3770) ;
	assign x_3767 = (x_3764 & x_3766) ;
	assign x_3762 = (x_3759 & x_3761) ;
	assign x_3758 = (x_3756 & x_3757) ;
	assign x_3753 = (x_3750 & x_3752) ;
	assign x_3749 = (x_3746 & x_3748) ;
	assign x_3744 = (x_3741 & x_3743) ;
	assign x_3740 = (x_3738 & x_3739) ;
	assign x_3734 = (x_3731 & x_3733) ;
	assign x_3730 = (x_3727 & x_3729) ;
	assign x_3725 = (x_3722 & x_3724) ;
	assign x_3721 = (x_3719 & x_3720) ;
	assign x_3716 = (x_3713 & x_3715) ;
	assign x_3712 = (x_3709 & x_3711) ;
	assign x_3707 = (x_3704 & x_3706) ;
	assign x_3703 = (x_3701 & x_3702) ;
	assign x_3696 = (x_3693 & x_3695) ;
	assign x_3692 = (x_3689 & x_3691) ;
	assign x_3687 = (x_3684 & x_3686) ;
	assign x_3683 = (x_3681 & x_3682) ;
	assign x_3678 = (x_3675 & x_3677) ;
	assign x_3674 = (x_3671 & x_3673) ;
	assign x_3669 = (x_3666 & x_3668) ;
	assign x_3665 = (x_3663 & x_3664) ;
	assign x_3659 = (x_3656 & x_3658) ;
	assign x_3655 = (x_3652 & x_3654) ;
	assign x_3650 = (x_3647 & x_3649) ;
	assign x_3646 = (x_3644 & x_3645) ;
	assign x_3641 = (x_3638 & x_3640) ;
	assign x_3637 = (x_3635 & x_3636) ;
	assign x_3633 = (x_3630 & x_3632) ;
	assign x_3629 = (x_3627 & x_3628) ;
	assign x_3618 = (x_3615 & x_3617) ;
	assign x_3614 = (x_3611 & x_3613) ;
	assign x_3609 = (x_3606 & x_3608) ;
	assign x_3605 = (x_3603 & x_3604) ;
	assign x_3600 = (x_3597 & x_3599) ;
	assign x_3596 = (x_3593 & x_3595) ;
	assign x_3591 = (x_3588 & x_3590) ;
	assign x_3587 = (x_3585 & x_3586) ;
	assign x_3581 = (x_3578 & x_3580) ;
	assign x_3577 = (x_3574 & x_3576) ;
	assign x_3572 = (x_3569 & x_3571) ;
	assign x_3568 = (x_3566 & x_3567) ;
	assign x_3563 = (x_3560 & x_3562) ;
	assign x_3559 = (x_3556 & x_3558) ;
	assign x_3554 = (x_3551 & x_3553) ;
	assign x_3550 = (x_3548 & x_3549) ;
	assign x_3543 = (x_3540 & x_3542) ;
	assign x_3539 = (x_3536 & x_3538) ;
	assign x_3534 = (x_3531 & x_3533) ;
	assign x_3530 = (x_3528 & x_3529) ;
	assign x_3525 = (x_3522 & x_3524) ;
	assign x_3521 = (x_3518 & x_3520) ;
	assign x_3516 = (x_3513 & x_3515) ;
	assign x_3512 = (x_3510 & x_3511) ;
	assign x_3506 = (x_3503 & x_3505) ;
	assign x_3502 = (x_3499 & x_3501) ;
	assign x_3497 = (x_3494 & x_3496) ;
	assign x_3493 = (x_3491 & x_3492) ;
	assign x_3488 = (x_3485 & x_3487) ;
	assign x_3484 = (x_3481 & x_3483) ;
	assign x_3479 = (x_3476 & x_3478) ;
	assign x_3475 = (x_3473 & x_3474) ;
	assign x_3467 = (x_3464 & x_3466) ;
	assign x_3463 = (x_3460 & x_3462) ;
	assign x_3458 = (x_3455 & x_3457) ;
	assign x_3454 = (x_3452 & x_3453) ;
	assign x_3449 = (x_3446 & x_3448) ;
	assign x_3445 = (x_3442 & x_3444) ;
	assign x_3440 = (x_3437 & x_3439) ;
	assign x_3436 = (x_3434 & x_3435) ;
	assign x_3430 = (x_3427 & x_3429) ;
	assign x_3426 = (x_3423 & x_3425) ;
	assign x_3421 = (x_3418 & x_3420) ;
	assign x_3417 = (x_3415 & x_3416) ;
	assign x_3412 = (x_3409 & x_3411) ;
	assign x_3408 = (x_3405 & x_3407) ;
	assign x_3403 = (x_3400 & x_3402) ;
	assign x_3399 = (x_3397 & x_3398) ;
	assign x_3392 = (x_3389 & x_3391) ;
	assign x_3388 = (x_3385 & x_3387) ;
	assign x_3383 = (x_3380 & x_3382) ;
	assign x_3379 = (x_3377 & x_3378) ;
	assign x_3374 = (x_3371 & x_3373) ;
	assign x_3370 = (x_3367 & x_3369) ;
	assign x_3365 = (x_3362 & x_3364) ;
	assign x_3361 = (x_3359 & x_3360) ;
	assign x_3355 = (x_3352 & x_3354) ;
	assign x_3351 = (x_3348 & x_3350) ;
	assign x_3346 = (x_3343 & x_3345) ;
	assign x_3342 = (x_3340 & x_3341) ;
	assign x_3337 = (x_3334 & x_3336) ;
	assign x_3333 = (x_3331 & x_3332) ;
	assign x_3329 = (x_3326 & x_3328) ;
	assign x_3325 = (x_3323 & x_3324) ;
	assign x_3316 = (x_3313 & x_3315) ;
	assign x_3312 = (x_3309 & x_3311) ;
	assign x_3307 = (x_3304 & x_3306) ;
	assign x_3303 = (x_3301 & x_3302) ;
	assign x_3298 = (x_3295 & x_3297) ;
	assign x_3294 = (x_3291 & x_3293) ;
	assign x_3289 = (x_3286 & x_3288) ;
	assign x_3285 = (x_3283 & x_3284) ;
	assign x_3279 = (x_3276 & x_3278) ;
	assign x_3275 = (x_3272 & x_3274) ;
	assign x_3270 = (x_3267 & x_3269) ;
	assign x_3266 = (x_3264 & x_3265) ;
	assign x_3261 = (x_3258 & x_3260) ;
	assign x_3257 = (x_3254 & x_3256) ;
	assign x_3252 = (x_3249 & x_3251) ;
	assign x_3248 = (x_3246 & x_3247) ;
	assign x_3241 = (x_3238 & x_3240) ;
	assign x_3237 = (x_3234 & x_3236) ;
	assign x_3232 = (x_3229 & x_3231) ;
	assign x_3228 = (x_3226 & x_3227) ;
	assign x_3223 = (x_3220 & x_3222) ;
	assign x_3219 = (x_3216 & x_3218) ;
	assign x_3214 = (x_3211 & x_3213) ;
	assign x_3210 = (x_3208 & x_3209) ;
	assign x_3204 = (x_3201 & x_3203) ;
	assign x_3200 = (x_3197 & x_3199) ;
	assign x_3195 = (x_3192 & x_3194) ;
	assign x_3191 = (x_3189 & x_3190) ;
	assign x_3186 = (x_3183 & x_3185) ;
	assign x_3182 = (x_3180 & x_3181) ;
	assign x_3178 = (x_3175 & x_3177) ;
	assign x_3174 = (x_3172 & x_3173) ;
	assign x_3166 = (x_3163 & x_3165) ;
	assign x_3162 = (x_3159 & x_3161) ;
	assign x_3157 = (x_3154 & x_3156) ;
	assign x_3153 = (x_3151 & x_3152) ;
	assign x_3148 = (x_3145 & x_3147) ;
	assign x_3144 = (x_3141 & x_3143) ;
	assign x_3139 = (x_3136 & x_3138) ;
	assign x_3135 = (x_3133 & x_3134) ;
	assign x_3129 = (x_3126 & x_3128) ;
	assign x_3125 = (x_3122 & x_3124) ;
	assign x_3120 = (x_3117 & x_3119) ;
	assign x_3116 = (x_3114 & x_3115) ;
	assign x_3111 = (x_3108 & x_3110) ;
	assign x_3107 = (x_3104 & x_3106) ;
	assign x_3102 = (x_3099 & x_3101) ;
	assign x_3098 = (x_3096 & x_3097) ;
	assign x_3091 = (x_3088 & x_3090) ;
	assign x_3087 = (x_3084 & x_3086) ;
	assign x_3082 = (x_3079 & x_3081) ;
	assign x_3078 = (x_3076 & x_3077) ;
	assign x_3073 = (x_3070 & x_3072) ;
	assign x_3069 = (x_3066 & x_3068) ;
	assign x_3064 = (x_3061 & x_3063) ;
	assign x_3060 = (x_3058 & x_3059) ;
	assign x_3054 = (x_3051 & x_3053) ;
	assign x_3050 = (x_3047 & x_3049) ;
	assign x_3045 = (x_3042 & x_3044) ;
	assign x_3041 = (x_3039 & x_3040) ;
	assign x_3036 = (x_3033 & x_3035) ;
	assign x_3032 = (x_3030 & x_3031) ;
	assign x_3028 = (x_3025 & x_3027) ;
	assign x_3024 = (x_3022 & x_3023) ;
	assign x_3014 = (x_3011 & x_3013) ;
	assign x_3010 = (x_3007 & x_3009) ;
	assign x_3005 = (x_3002 & x_3004) ;
	assign x_3001 = (x_2999 & x_3000) ;
	assign x_2996 = (x_2993 & x_2995) ;
	assign x_2992 = (x_2989 & x_2991) ;
	assign x_2987 = (x_2984 & x_2986) ;
	assign x_2983 = (x_2981 & x_2982) ;
	assign x_2977 = (x_2974 & x_2976) ;
	assign x_2973 = (x_2970 & x_2972) ;
	assign x_2968 = (x_2965 & x_2967) ;
	assign x_2964 = (x_2962 & x_2963) ;
	assign x_2959 = (x_2956 & x_2958) ;
	assign x_2955 = (x_2952 & x_2954) ;
	assign x_2950 = (x_2947 & x_2949) ;
	assign x_2946 = (x_2944 & x_2945) ;
	assign x_2939 = (x_2936 & x_2938) ;
	assign x_2935 = (x_2932 & x_2934) ;
	assign x_2930 = (x_2927 & x_2929) ;
	assign x_2926 = (x_2924 & x_2925) ;
	assign x_2921 = (x_2918 & x_2920) ;
	assign x_2917 = (x_2914 & x_2916) ;
	assign x_2912 = (x_2909 & x_2911) ;
	assign x_2908 = (x_2906 & x_2907) ;
	assign x_2902 = (x_2899 & x_2901) ;
	assign x_2898 = (x_2895 & x_2897) ;
	assign x_2893 = (x_2890 & x_2892) ;
	assign x_2889 = (x_2887 & x_2888) ;
	assign x_2884 = (x_2881 & x_2883) ;
	assign x_2880 = (x_2878 & x_2879) ;
	assign x_2876 = (x_2873 & x_2875) ;
	assign x_2872 = (x_2870 & x_2871) ;
	assign x_2864 = (x_2861 & x_2863) ;
	assign x_2860 = (x_2857 & x_2859) ;
	assign x_2855 = (x_2852 & x_2854) ;
	assign x_2851 = (x_2849 & x_2850) ;
	assign x_2846 = (x_2843 & x_2845) ;
	assign x_2842 = (x_2839 & x_2841) ;
	assign x_2837 = (x_2834 & x_2836) ;
	assign x_2833 = (x_2831 & x_2832) ;
	assign x_2827 = (x_2824 & x_2826) ;
	assign x_2823 = (x_2820 & x_2822) ;
	assign x_2818 = (x_2815 & x_2817) ;
	assign x_2814 = (x_2812 & x_2813) ;
	assign x_2809 = (x_2806 & x_2808) ;
	assign x_2805 = (x_2802 & x_2804) ;
	assign x_2800 = (x_2797 & x_2799) ;
	assign x_2796 = (x_2794 & x_2795) ;
	assign x_2789 = (x_2786 & x_2788) ;
	assign x_2785 = (x_2782 & x_2784) ;
	assign x_2780 = (x_2777 & x_2779) ;
	assign x_2776 = (x_2774 & x_2775) ;
	assign x_2771 = (x_2768 & x_2770) ;
	assign x_2767 = (x_2764 & x_2766) ;
	assign x_2762 = (x_2759 & x_2761) ;
	assign x_2758 = (x_2756 & x_2757) ;
	assign x_2752 = (x_2749 & x_2751) ;
	assign x_2748 = (x_2745 & x_2747) ;
	assign x_2743 = (x_2740 & x_2742) ;
	assign x_2739 = (x_2737 & x_2738) ;
	assign x_2734 = (x_2731 & x_2733) ;
	assign x_2730 = (x_2728 & x_2729) ;
	assign x_2726 = (x_2723 & x_2725) ;
	assign x_2722 = (x_2720 & x_2721) ;
	assign x_2713 = (x_2710 & x_2712) ;
	assign x_2709 = (x_2706 & x_2708) ;
	assign x_2704 = (x_2701 & x_2703) ;
	assign x_2700 = (x_2698 & x_2699) ;
	assign x_2695 = (x_2692 & x_2694) ;
	assign x_2691 = (x_2688 & x_2690) ;
	assign x_2686 = (x_2683 & x_2685) ;
	assign x_2682 = (x_2680 & x_2681) ;
	assign x_2676 = (x_2673 & x_2675) ;
	assign x_2672 = (x_2669 & x_2671) ;
	assign x_2667 = (x_2664 & x_2666) ;
	assign x_2663 = (x_2661 & x_2662) ;
	assign x_2658 = (x_2655 & x_2657) ;
	assign x_2654 = (x_2651 & x_2653) ;
	assign x_2649 = (x_2646 & x_2648) ;
	assign x_2645 = (x_2643 & x_2644) ;
	assign x_2638 = (x_2635 & x_2637) ;
	assign x_2634 = (x_2631 & x_2633) ;
	assign x_2629 = (x_2626 & x_2628) ;
	assign x_2625 = (x_2623 & x_2624) ;
	assign x_2620 = (x_2617 & x_2619) ;
	assign x_2616 = (x_2613 & x_2615) ;
	assign x_2611 = (x_2608 & x_2610) ;
	assign x_2607 = (x_2605 & x_2606) ;
	assign x_2601 = (x_2598 & x_2600) ;
	assign x_2597 = (x_2594 & x_2596) ;
	assign x_2592 = (x_2589 & x_2591) ;
	assign x_2588 = (x_2586 & x_2587) ;
	assign x_2583 = (x_2580 & x_2582) ;
	assign x_2579 = (x_2577 & x_2578) ;
	assign x_2575 = (x_2572 & x_2574) ;
	assign x_2571 = (x_2569 & x_2570) ;
	assign x_2563 = (x_2560 & x_2562) ;
	assign x_2559 = (x_2556 & x_2558) ;
	assign x_2554 = (x_2551 & x_2553) ;
	assign x_2550 = (x_2548 & x_2549) ;
	assign x_2545 = (x_2542 & x_2544) ;
	assign x_2541 = (x_2538 & x_2540) ;
	assign x_2536 = (x_2533 & x_2535) ;
	assign x_2532 = (x_2530 & x_2531) ;
	assign x_2526 = (x_2523 & x_2525) ;
	assign x_2522 = (x_2519 & x_2521) ;
	assign x_2517 = (x_2514 & x_2516) ;
	assign x_2513 = (x_2511 & x_2512) ;
	assign x_2508 = (x_2505 & x_2507) ;
	assign x_2504 = (x_2501 & x_2503) ;
	assign x_2499 = (x_2496 & x_2498) ;
	assign x_2495 = (x_2493 & x_2494) ;
	assign x_2488 = (x_2485 & x_2487) ;
	assign x_2484 = (x_2481 & x_2483) ;
	assign x_2479 = (x_2476 & x_2478) ;
	assign x_2475 = (x_2473 & x_2474) ;
	assign x_2470 = (x_2467 & x_2469) ;
	assign x_2466 = (x_2463 & x_2465) ;
	assign x_2461 = (x_2458 & x_2460) ;
	assign x_2457 = (x_2455 & x_2456) ;
	assign x_2451 = (x_2448 & x_2450) ;
	assign x_2447 = (x_2444 & x_2446) ;
	assign x_2442 = (x_2439 & x_2441) ;
	assign x_2438 = (x_2436 & x_2437) ;
	assign x_2433 = (x_2430 & x_2432) ;
	assign x_2429 = (x_2427 & x_2428) ;
	assign x_2425 = (x_2422 & x_2424) ;
	assign x_2421 = (x_2419 & x_2420) ;
	assign x_4827 = (x_4822 & x_4826) ;
	assign x_4818 = (x_4813 & x_4817) ;
	assign x_4809 = (x_4804 & x_4808) ;
	assign x_4800 = (x_4795 & x_4799) ;
	assign x_4790 = (x_4785 & x_4789) ;
	assign x_4781 = (x_4776 & x_4780) ;
	assign x_4772 = (x_4767 & x_4771) ;
	assign x_4763 = (x_4758 & x_4762) ;
	assign x_4752 = (x_4747 & x_4751) ;
	assign x_4743 = (x_4738 & x_4742) ;
	assign x_4734 = (x_4729 & x_4733) ;
	assign x_4725 = (x_4720 & x_4724) ;
	assign x_4715 = (x_4710 & x_4714) ;
	assign x_4706 = (x_4701 & x_4705) ;
	assign x_4697 = (x_4692 & x_4696) ;
	assign x_4688 = (x_4683 & x_4687) ;
	assign x_4676 = (x_4671 & x_4675) ;
	assign x_4667 = (x_4662 & x_4666) ;
	assign x_4658 = (x_4653 & x_4657) ;
	assign x_4649 = (x_4644 & x_4648) ;
	assign x_4639 = (x_4634 & x_4638) ;
	assign x_4630 = (x_4625 & x_4629) ;
	assign x_4621 = (x_4616 & x_4620) ;
	assign x_4612 = (x_4607 & x_4611) ;
	assign x_4601 = (x_4596 & x_4600) ;
	assign x_4592 = (x_4587 & x_4591) ;
	assign x_4583 = (x_4578 & x_4582) ;
	assign x_4574 = (x_4569 & x_4573) ;
	assign x_4564 = (x_4559 & x_4563) ;
	assign x_4555 = (x_4550 & x_4554) ;
	assign x_4546 = (x_4541 & x_4545) ;
	assign x_4538 = (x_4533 & x_4537) ;
	assign x_4525 = (x_4520 & x_4524) ;
	assign x_4516 = (x_4511 & x_4515) ;
	assign x_4507 = (x_4502 & x_4506) ;
	assign x_4498 = (x_4493 & x_4497) ;
	assign x_4488 = (x_4483 & x_4487) ;
	assign x_4479 = (x_4474 & x_4478) ;
	assign x_4470 = (x_4465 & x_4469) ;
	assign x_4461 = (x_4456 & x_4460) ;
	assign x_4450 = (x_4445 & x_4449) ;
	assign x_4441 = (x_4436 & x_4440) ;
	assign x_4432 = (x_4427 & x_4431) ;
	assign x_4423 = (x_4418 & x_4422) ;
	assign x_4413 = (x_4408 & x_4412) ;
	assign x_4404 = (x_4399 & x_4403) ;
	assign x_4395 = (x_4390 & x_4394) ;
	assign x_4387 = (x_4382 & x_4386) ;
	assign x_4375 = (x_4370 & x_4374) ;
	assign x_4366 = (x_4361 & x_4365) ;
	assign x_4357 = (x_4352 & x_4356) ;
	assign x_4348 = (x_4343 & x_4347) ;
	assign x_4338 = (x_4333 & x_4337) ;
	assign x_4329 = (x_4324 & x_4328) ;
	assign x_4320 = (x_4315 & x_4319) ;
	assign x_4311 = (x_4306 & x_4310) ;
	assign x_4300 = (x_4295 & x_4299) ;
	assign x_4291 = (x_4286 & x_4290) ;
	assign x_4282 = (x_4277 & x_4281) ;
	assign x_4273 = (x_4268 & x_4272) ;
	assign x_4263 = (x_4258 & x_4262) ;
	assign x_4254 = (x_4249 & x_4253) ;
	assign x_4245 = (x_4240 & x_4244) ;
	assign x_4237 = (x_4232 & x_4236) ;
	assign x_4223 = (x_4218 & x_4222) ;
	assign x_4214 = (x_4209 & x_4213) ;
	assign x_4205 = (x_4200 & x_4204) ;
	assign x_4196 = (x_4191 & x_4195) ;
	assign x_4186 = (x_4181 & x_4185) ;
	assign x_4177 = (x_4172 & x_4176) ;
	assign x_4168 = (x_4163 & x_4167) ;
	assign x_4159 = (x_4154 & x_4158) ;
	assign x_4148 = (x_4143 & x_4147) ;
	assign x_4139 = (x_4134 & x_4138) ;
	assign x_4130 = (x_4125 & x_4129) ;
	assign x_4121 = (x_4116 & x_4120) ;
	assign x_4111 = (x_4106 & x_4110) ;
	assign x_4102 = (x_4097 & x_4101) ;
	assign x_4093 = (x_4088 & x_4092) ;
	assign x_4085 = (x_4080 & x_4084) ;
	assign x_4073 = (x_4068 & x_4072) ;
	assign x_4064 = (x_4059 & x_4063) ;
	assign x_4055 = (x_4050 & x_4054) ;
	assign x_4046 = (x_4041 & x_4045) ;
	assign x_4036 = (x_4031 & x_4035) ;
	assign x_4027 = (x_4022 & x_4026) ;
	assign x_4018 = (x_4013 & x_4017) ;
	assign x_4009 = (x_4004 & x_4008) ;
	assign x_3998 = (x_3993 & x_3997) ;
	assign x_3989 = (x_3984 & x_3988) ;
	assign x_3980 = (x_3975 & x_3979) ;
	assign x_3971 = (x_3966 & x_3970) ;
	assign x_3961 = (x_3956 & x_3960) ;
	assign x_3952 = (x_3947 & x_3951) ;
	assign x_3943 = (x_3938 & x_3942) ;
	assign x_3935 = (x_3930 & x_3934) ;
	assign x_3922 = (x_3917 & x_3921) ;
	assign x_3913 = (x_3908 & x_3912) ;
	assign x_3904 = (x_3899 & x_3903) ;
	assign x_3895 = (x_3890 & x_3894) ;
	assign x_3885 = (x_3880 & x_3884) ;
	assign x_3876 = (x_3871 & x_3875) ;
	assign x_3867 = (x_3862 & x_3866) ;
	assign x_3858 = (x_3853 & x_3857) ;
	assign x_3847 = (x_3842 & x_3846) ;
	assign x_3838 = (x_3833 & x_3837) ;
	assign x_3829 = (x_3824 & x_3828) ;
	assign x_3820 = (x_3815 & x_3819) ;
	assign x_3810 = (x_3805 & x_3809) ;
	assign x_3801 = (x_3796 & x_3800) ;
	assign x_3792 = (x_3787 & x_3791) ;
	assign x_3784 = (x_3779 & x_3783) ;
	assign x_3772 = (x_3767 & x_3771) ;
	assign x_3763 = (x_3758 & x_3762) ;
	assign x_3754 = (x_3749 & x_3753) ;
	assign x_3745 = (x_3740 & x_3744) ;
	assign x_3735 = (x_3730 & x_3734) ;
	assign x_3726 = (x_3721 & x_3725) ;
	assign x_3717 = (x_3712 & x_3716) ;
	assign x_3708 = (x_3703 & x_3707) ;
	assign x_3697 = (x_3692 & x_3696) ;
	assign x_3688 = (x_3683 & x_3687) ;
	assign x_3679 = (x_3674 & x_3678) ;
	assign x_3670 = (x_3665 & x_3669) ;
	assign x_3660 = (x_3655 & x_3659) ;
	assign x_3651 = (x_3646 & x_3650) ;
	assign x_3642 = (x_3637 & x_3641) ;
	assign x_3634 = (x_3629 & x_3633) ;
	assign x_3619 = (x_3614 & x_3618) ;
	assign x_3610 = (x_3605 & x_3609) ;
	assign x_3601 = (x_3596 & x_3600) ;
	assign x_3592 = (x_3587 & x_3591) ;
	assign x_3582 = (x_3577 & x_3581) ;
	assign x_3573 = (x_3568 & x_3572) ;
	assign x_3564 = (x_3559 & x_3563) ;
	assign x_3555 = (x_3550 & x_3554) ;
	assign x_3544 = (x_3539 & x_3543) ;
	assign x_3535 = (x_3530 & x_3534) ;
	assign x_3526 = (x_3521 & x_3525) ;
	assign x_3517 = (x_3512 & x_3516) ;
	assign x_3507 = (x_3502 & x_3506) ;
	assign x_3498 = (x_3493 & x_3497) ;
	assign x_3489 = (x_3484 & x_3488) ;
	assign x_3480 = (x_3475 & x_3479) ;
	assign x_3468 = (x_3463 & x_3467) ;
	assign x_3459 = (x_3454 & x_3458) ;
	assign x_3450 = (x_3445 & x_3449) ;
	assign x_3441 = (x_3436 & x_3440) ;
	assign x_3431 = (x_3426 & x_3430) ;
	assign x_3422 = (x_3417 & x_3421) ;
	assign x_3413 = (x_3408 & x_3412) ;
	assign x_3404 = (x_3399 & x_3403) ;
	assign x_3393 = (x_3388 & x_3392) ;
	assign x_3384 = (x_3379 & x_3383) ;
	assign x_3375 = (x_3370 & x_3374) ;
	assign x_3366 = (x_3361 & x_3365) ;
	assign x_3356 = (x_3351 & x_3355) ;
	assign x_3347 = (x_3342 & x_3346) ;
	assign x_3338 = (x_3333 & x_3337) ;
	assign x_3330 = (x_3325 & x_3329) ;
	assign x_3317 = (x_3312 & x_3316) ;
	assign x_3308 = (x_3303 & x_3307) ;
	assign x_3299 = (x_3294 & x_3298) ;
	assign x_3290 = (x_3285 & x_3289) ;
	assign x_3280 = (x_3275 & x_3279) ;
	assign x_3271 = (x_3266 & x_3270) ;
	assign x_3262 = (x_3257 & x_3261) ;
	assign x_3253 = (x_3248 & x_3252) ;
	assign x_3242 = (x_3237 & x_3241) ;
	assign x_3233 = (x_3228 & x_3232) ;
	assign x_3224 = (x_3219 & x_3223) ;
	assign x_3215 = (x_3210 & x_3214) ;
	assign x_3205 = (x_3200 & x_3204) ;
	assign x_3196 = (x_3191 & x_3195) ;
	assign x_3187 = (x_3182 & x_3186) ;
	assign x_3179 = (x_3174 & x_3178) ;
	assign x_3167 = (x_3162 & x_3166) ;
	assign x_3158 = (x_3153 & x_3157) ;
	assign x_3149 = (x_3144 & x_3148) ;
	assign x_3140 = (x_3135 & x_3139) ;
	assign x_3130 = (x_3125 & x_3129) ;
	assign x_3121 = (x_3116 & x_3120) ;
	assign x_3112 = (x_3107 & x_3111) ;
	assign x_3103 = (x_3098 & x_3102) ;
	assign x_3092 = (x_3087 & x_3091) ;
	assign x_3083 = (x_3078 & x_3082) ;
	assign x_3074 = (x_3069 & x_3073) ;
	assign x_3065 = (x_3060 & x_3064) ;
	assign x_3055 = (x_3050 & x_3054) ;
	assign x_3046 = (x_3041 & x_3045) ;
	assign x_3037 = (x_3032 & x_3036) ;
	assign x_3029 = (x_3024 & x_3028) ;
	assign x_3015 = (x_3010 & x_3014) ;
	assign x_3006 = (x_3001 & x_3005) ;
	assign x_2997 = (x_2992 & x_2996) ;
	assign x_2988 = (x_2983 & x_2987) ;
	assign x_2978 = (x_2973 & x_2977) ;
	assign x_2969 = (x_2964 & x_2968) ;
	assign x_2960 = (x_2955 & x_2959) ;
	assign x_2951 = (x_2946 & x_2950) ;
	assign x_2940 = (x_2935 & x_2939) ;
	assign x_2931 = (x_2926 & x_2930) ;
	assign x_2922 = (x_2917 & x_2921) ;
	assign x_2913 = (x_2908 & x_2912) ;
	assign x_2903 = (x_2898 & x_2902) ;
	assign x_2894 = (x_2889 & x_2893) ;
	assign x_2885 = (x_2880 & x_2884) ;
	assign x_2877 = (x_2872 & x_2876) ;
	assign x_2865 = (x_2860 & x_2864) ;
	assign x_2856 = (x_2851 & x_2855) ;
	assign x_2847 = (x_2842 & x_2846) ;
	assign x_2838 = (x_2833 & x_2837) ;
	assign x_2828 = (x_2823 & x_2827) ;
	assign x_2819 = (x_2814 & x_2818) ;
	assign x_2810 = (x_2805 & x_2809) ;
	assign x_2801 = (x_2796 & x_2800) ;
	assign x_2790 = (x_2785 & x_2789) ;
	assign x_2781 = (x_2776 & x_2780) ;
	assign x_2772 = (x_2767 & x_2771) ;
	assign x_2763 = (x_2758 & x_2762) ;
	assign x_2753 = (x_2748 & x_2752) ;
	assign x_2744 = (x_2739 & x_2743) ;
	assign x_2735 = (x_2730 & x_2734) ;
	assign x_2727 = (x_2722 & x_2726) ;
	assign x_2714 = (x_2709 & x_2713) ;
	assign x_2705 = (x_2700 & x_2704) ;
	assign x_2696 = (x_2691 & x_2695) ;
	assign x_2687 = (x_2682 & x_2686) ;
	assign x_2677 = (x_2672 & x_2676) ;
	assign x_2668 = (x_2663 & x_2667) ;
	assign x_2659 = (x_2654 & x_2658) ;
	assign x_2650 = (x_2645 & x_2649) ;
	assign x_2639 = (x_2634 & x_2638) ;
	assign x_2630 = (x_2625 & x_2629) ;
	assign x_2621 = (x_2616 & x_2620) ;
	assign x_2612 = (x_2607 & x_2611) ;
	assign x_2602 = (x_2597 & x_2601) ;
	assign x_2593 = (x_2588 & x_2592) ;
	assign x_2584 = (x_2579 & x_2583) ;
	assign x_2576 = (x_2571 & x_2575) ;
	assign x_2564 = (x_2559 & x_2563) ;
	assign x_2555 = (x_2550 & x_2554) ;
	assign x_2546 = (x_2541 & x_2545) ;
	assign x_2537 = (x_2532 & x_2536) ;
	assign x_2527 = (x_2522 & x_2526) ;
	assign x_2518 = (x_2513 & x_2517) ;
	assign x_2509 = (x_2504 & x_2508) ;
	assign x_2500 = (x_2495 & x_2499) ;
	assign x_2489 = (x_2484 & x_2488) ;
	assign x_2480 = (x_2475 & x_2479) ;
	assign x_2471 = (x_2466 & x_2470) ;
	assign x_2462 = (x_2457 & x_2461) ;
	assign x_2452 = (x_2447 & x_2451) ;
	assign x_2443 = (x_2438 & x_2442) ;
	assign x_2434 = (x_2429 & x_2433) ;
	assign x_2426 = (x_2421 & x_2425) ;
	assign x_4828 = (x_4818 & x_4827) ;
	assign x_4810 = (x_4800 & x_4809) ;
	assign x_4791 = (x_4781 & x_4790) ;
	assign x_4773 = (x_4763 & x_4772) ;
	assign x_4753 = (x_4743 & x_4752) ;
	assign x_4735 = (x_4725 & x_4734) ;
	assign x_4716 = (x_4706 & x_4715) ;
	assign x_4698 = (x_4688 & x_4697) ;
	assign x_4677 = (x_4667 & x_4676) ;
	assign x_4659 = (x_4649 & x_4658) ;
	assign x_4640 = (x_4630 & x_4639) ;
	assign x_4622 = (x_4612 & x_4621) ;
	assign x_4602 = (x_4592 & x_4601) ;
	assign x_4584 = (x_4574 & x_4583) ;
	assign x_4565 = (x_4555 & x_4564) ;
	assign x_4547 = (x_4538 & x_4546) ;
	assign x_4526 = (x_4516 & x_4525) ;
	assign x_4508 = (x_4498 & x_4507) ;
	assign x_4489 = (x_4479 & x_4488) ;
	assign x_4471 = (x_4461 & x_4470) ;
	assign x_4451 = (x_4441 & x_4450) ;
	assign x_4433 = (x_4423 & x_4432) ;
	assign x_4414 = (x_4404 & x_4413) ;
	assign x_4396 = (x_4387 & x_4395) ;
	assign x_4376 = (x_4366 & x_4375) ;
	assign x_4358 = (x_4348 & x_4357) ;
	assign x_4339 = (x_4329 & x_4338) ;
	assign x_4321 = (x_4311 & x_4320) ;
	assign x_4301 = (x_4291 & x_4300) ;
	assign x_4283 = (x_4273 & x_4282) ;
	assign x_4264 = (x_4254 & x_4263) ;
	assign x_4246 = (x_4237 & x_4245) ;
	assign x_4224 = (x_4214 & x_4223) ;
	assign x_4206 = (x_4196 & x_4205) ;
	assign x_4187 = (x_4177 & x_4186) ;
	assign x_4169 = (x_4159 & x_4168) ;
	assign x_4149 = (x_4139 & x_4148) ;
	assign x_4131 = (x_4121 & x_4130) ;
	assign x_4112 = (x_4102 & x_4111) ;
	assign x_4094 = (x_4085 & x_4093) ;
	assign x_4074 = (x_4064 & x_4073) ;
	assign x_4056 = (x_4046 & x_4055) ;
	assign x_4037 = (x_4027 & x_4036) ;
	assign x_4019 = (x_4009 & x_4018) ;
	assign x_3999 = (x_3989 & x_3998) ;
	assign x_3981 = (x_3971 & x_3980) ;
	assign x_3962 = (x_3952 & x_3961) ;
	assign x_3944 = (x_3935 & x_3943) ;
	assign x_3923 = (x_3913 & x_3922) ;
	assign x_3905 = (x_3895 & x_3904) ;
	assign x_3886 = (x_3876 & x_3885) ;
	assign x_3868 = (x_3858 & x_3867) ;
	assign x_3848 = (x_3838 & x_3847) ;
	assign x_3830 = (x_3820 & x_3829) ;
	assign x_3811 = (x_3801 & x_3810) ;
	assign x_3793 = (x_3784 & x_3792) ;
	assign x_3773 = (x_3763 & x_3772) ;
	assign x_3755 = (x_3745 & x_3754) ;
	assign x_3736 = (x_3726 & x_3735) ;
	assign x_3718 = (x_3708 & x_3717) ;
	assign x_3698 = (x_3688 & x_3697) ;
	assign x_3680 = (x_3670 & x_3679) ;
	assign x_3661 = (x_3651 & x_3660) ;
	assign x_3643 = (x_3634 & x_3642) ;
	assign x_3620 = (x_3610 & x_3619) ;
	assign x_3602 = (x_3592 & x_3601) ;
	assign x_3583 = (x_3573 & x_3582) ;
	assign x_3565 = (x_3555 & x_3564) ;
	assign x_3545 = (x_3535 & x_3544) ;
	assign x_3527 = (x_3517 & x_3526) ;
	assign x_3508 = (x_3498 & x_3507) ;
	assign x_3490 = (x_3480 & x_3489) ;
	assign x_3469 = (x_3459 & x_3468) ;
	assign x_3451 = (x_3441 & x_3450) ;
	assign x_3432 = (x_3422 & x_3431) ;
	assign x_3414 = (x_3404 & x_3413) ;
	assign x_3394 = (x_3384 & x_3393) ;
	assign x_3376 = (x_3366 & x_3375) ;
	assign x_3357 = (x_3347 & x_3356) ;
	assign x_3339 = (x_3330 & x_3338) ;
	assign x_3318 = (x_3308 & x_3317) ;
	assign x_3300 = (x_3290 & x_3299) ;
	assign x_3281 = (x_3271 & x_3280) ;
	assign x_3263 = (x_3253 & x_3262) ;
	assign x_3243 = (x_3233 & x_3242) ;
	assign x_3225 = (x_3215 & x_3224) ;
	assign x_3206 = (x_3196 & x_3205) ;
	assign x_3188 = (x_3179 & x_3187) ;
	assign x_3168 = (x_3158 & x_3167) ;
	assign x_3150 = (x_3140 & x_3149) ;
	assign x_3131 = (x_3121 & x_3130) ;
	assign x_3113 = (x_3103 & x_3112) ;
	assign x_3093 = (x_3083 & x_3092) ;
	assign x_3075 = (x_3065 & x_3074) ;
	assign x_3056 = (x_3046 & x_3055) ;
	assign x_3038 = (x_3029 & x_3037) ;
	assign x_3016 = (x_3006 & x_3015) ;
	assign x_2998 = (x_2988 & x_2997) ;
	assign x_2979 = (x_2969 & x_2978) ;
	assign x_2961 = (x_2951 & x_2960) ;
	assign x_2941 = (x_2931 & x_2940) ;
	assign x_2923 = (x_2913 & x_2922) ;
	assign x_2904 = (x_2894 & x_2903) ;
	assign x_2886 = (x_2877 & x_2885) ;
	assign x_2866 = (x_2856 & x_2865) ;
	assign x_2848 = (x_2838 & x_2847) ;
	assign x_2829 = (x_2819 & x_2828) ;
	assign x_2811 = (x_2801 & x_2810) ;
	assign x_2791 = (x_2781 & x_2790) ;
	assign x_2773 = (x_2763 & x_2772) ;
	assign x_2754 = (x_2744 & x_2753) ;
	assign x_2736 = (x_2727 & x_2735) ;
	assign x_2715 = (x_2705 & x_2714) ;
	assign x_2697 = (x_2687 & x_2696) ;
	assign x_2678 = (x_2668 & x_2677) ;
	assign x_2660 = (x_2650 & x_2659) ;
	assign x_2640 = (x_2630 & x_2639) ;
	assign x_2622 = (x_2612 & x_2621) ;
	assign x_2603 = (x_2593 & x_2602) ;
	assign x_2585 = (x_2576 & x_2584) ;
	assign x_2565 = (x_2555 & x_2564) ;
	assign x_2547 = (x_2537 & x_2546) ;
	assign x_2528 = (x_2518 & x_2527) ;
	assign x_2510 = (x_2500 & x_2509) ;
	assign x_2490 = (x_2480 & x_2489) ;
	assign x_2472 = (x_2462 & x_2471) ;
	assign x_2453 = (x_2443 & x_2452) ;
	assign x_2435 = (x_2426 & x_2434) ;
	assign x_4829 = (x_4810 & x_4828) ;
	assign x_4792 = (x_4773 & x_4791) ;
	assign x_4754 = (x_4735 & x_4753) ;
	assign x_4717 = (x_4698 & x_4716) ;
	assign x_4678 = (x_4659 & x_4677) ;
	assign x_4641 = (x_4622 & x_4640) ;
	assign x_4603 = (x_4584 & x_4602) ;
	assign x_4566 = (x_4547 & x_4565) ;
	assign x_4527 = (x_4508 & x_4526) ;
	assign x_4490 = (x_4471 & x_4489) ;
	assign x_4452 = (x_4433 & x_4451) ;
	assign x_4415 = (x_4396 & x_4414) ;
	assign x_4377 = (x_4358 & x_4376) ;
	assign x_4340 = (x_4321 & x_4339) ;
	assign x_4302 = (x_4283 & x_4301) ;
	assign x_4265 = (x_4246 & x_4264) ;
	assign x_4225 = (x_4206 & x_4224) ;
	assign x_4188 = (x_4169 & x_4187) ;
	assign x_4150 = (x_4131 & x_4149) ;
	assign x_4113 = (x_4094 & x_4112) ;
	assign x_4075 = (x_4056 & x_4074) ;
	assign x_4038 = (x_4019 & x_4037) ;
	assign x_4000 = (x_3981 & x_3999) ;
	assign x_3963 = (x_3944 & x_3962) ;
	assign x_3924 = (x_3905 & x_3923) ;
	assign x_3887 = (x_3868 & x_3886) ;
	assign x_3849 = (x_3830 & x_3848) ;
	assign x_3812 = (x_3793 & x_3811) ;
	assign x_3774 = (x_3755 & x_3773) ;
	assign x_3737 = (x_3718 & x_3736) ;
	assign x_3699 = (x_3680 & x_3698) ;
	assign x_3662 = (x_3643 & x_3661) ;
	assign x_3621 = (x_3602 & x_3620) ;
	assign x_3584 = (x_3565 & x_3583) ;
	assign x_3546 = (x_3527 & x_3545) ;
	assign x_3509 = (x_3490 & x_3508) ;
	assign x_3470 = (x_3451 & x_3469) ;
	assign x_3433 = (x_3414 & x_3432) ;
	assign x_3395 = (x_3376 & x_3394) ;
	assign x_3358 = (x_3339 & x_3357) ;
	assign x_3319 = (x_3300 & x_3318) ;
	assign x_3282 = (x_3263 & x_3281) ;
	assign x_3244 = (x_3225 & x_3243) ;
	assign x_3207 = (x_3188 & x_3206) ;
	assign x_3169 = (x_3150 & x_3168) ;
	assign x_3132 = (x_3113 & x_3131) ;
	assign x_3094 = (x_3075 & x_3093) ;
	assign x_3057 = (x_3038 & x_3056) ;
	assign x_3017 = (x_2998 & x_3016) ;
	assign x_2980 = (x_2961 & x_2979) ;
	assign x_2942 = (x_2923 & x_2941) ;
	assign x_2905 = (x_2886 & x_2904) ;
	assign x_2867 = (x_2848 & x_2866) ;
	assign x_2830 = (x_2811 & x_2829) ;
	assign x_2792 = (x_2773 & x_2791) ;
	assign x_2755 = (x_2736 & x_2754) ;
	assign x_2716 = (x_2697 & x_2715) ;
	assign x_2679 = (x_2660 & x_2678) ;
	assign x_2641 = (x_2622 & x_2640) ;
	assign x_2604 = (x_2585 & x_2603) ;
	assign x_2566 = (x_2547 & x_2565) ;
	assign x_2529 = (x_2510 & x_2528) ;
	assign x_2491 = (x_2472 & x_2490) ;
	assign x_2454 = (x_2435 & x_2453) ;
	assign x_4830 = (x_4792 & x_4829) ;
	assign x_4755 = (x_4717 & x_4754) ;
	assign x_4679 = (x_4641 & x_4678) ;
	assign x_4604 = (x_4566 & x_4603) ;
	assign x_4528 = (x_4490 & x_4527) ;
	assign x_4453 = (x_4415 & x_4452) ;
	assign x_4378 = (x_4340 & x_4377) ;
	assign x_4303 = (x_4265 & x_4302) ;
	assign x_4226 = (x_4188 & x_4225) ;
	assign x_4151 = (x_4113 & x_4150) ;
	assign x_4076 = (x_4038 & x_4075) ;
	assign x_4001 = (x_3963 & x_4000) ;
	assign x_3925 = (x_3887 & x_3924) ;
	assign x_3850 = (x_3812 & x_3849) ;
	assign x_3775 = (x_3737 & x_3774) ;
	assign x_3700 = (x_3662 & x_3699) ;
	assign x_3622 = (x_3584 & x_3621) ;
	assign x_3547 = (x_3509 & x_3546) ;
	assign x_3471 = (x_3433 & x_3470) ;
	assign x_3396 = (x_3358 & x_3395) ;
	assign x_3320 = (x_3282 & x_3319) ;
	assign x_3245 = (x_3207 & x_3244) ;
	assign x_3170 = (x_3132 & x_3169) ;
	assign x_3095 = (x_3057 & x_3094) ;
	assign x_3018 = (x_2980 & x_3017) ;
	assign x_2943 = (x_2905 & x_2942) ;
	assign x_2868 = (x_2830 & x_2867) ;
	assign x_2793 = (x_2755 & x_2792) ;
	assign x_2717 = (x_2679 & x_2716) ;
	assign x_2642 = (x_2604 & x_2641) ;
	assign x_2567 = (x_2529 & x_2566) ;
	assign x_2492 = (x_2454 & x_2491) ;
	assign x_4831 = (x_4755 & x_4830) ;
	assign x_4680 = (x_4604 & x_4679) ;
	assign x_4529 = (x_4453 & x_4528) ;
	assign x_4379 = (x_4303 & x_4378) ;
	assign x_4227 = (x_4151 & x_4226) ;
	assign x_4077 = (x_4001 & x_4076) ;
	assign x_3926 = (x_3850 & x_3925) ;
	assign x_3776 = (x_3700 & x_3775) ;
	assign x_3623 = (x_3547 & x_3622) ;
	assign x_3472 = (x_3396 & x_3471) ;
	assign x_3321 = (x_3245 & x_3320) ;
	assign x_3171 = (x_3095 & x_3170) ;
	assign x_3019 = (x_2943 & x_3018) ;
	assign x_2869 = (x_2793 & x_2868) ;
	assign x_2718 = (x_2642 & x_2717) ;
	assign x_2568 = (x_2492 & x_2567) ;
	assign x_4832 = (x_4680 & x_4831) ;
	assign x_4530 = (x_4379 & x_4529) ;
	assign x_4228 = (x_4077 & x_4227) ;
	assign x_3927 = (x_3776 & x_3926) ;
	assign x_3624 = (x_3472 & x_3623) ;
	assign x_3322 = (x_3171 & x_3321) ;
	assign x_3020 = (x_2869 & x_3019) ;
	assign x_2719 = (x_2568 & x_2718) ;
	assign x_4833 = (x_4530 & x_4832) ;
	assign x_4229 = (x_3927 & x_4228) ;
	assign x_3625 = (x_3322 & x_3624) ;
	assign x_3021 = (x_2719 & x_3020) ;
	assign x_4834 = (x_4229 & x_4833) ;
	assign x_3626 = (x_3021 & x_3625) ;
	assign x_4835 = (x_3626 & x_4834) ;
	assign v_1034 = 0 ;
	assign v_1033 = 0 ;
	assign v_994 = 0 ;
	assign v_985 = 0 ;
	assign v_976 = 0 ;
	assign v_967 = 0 ;
	assign v_958 = 0 ;
	assign v_949 = 0 ;
	assign v_908 = 0 ;
	assign v_865 = 0 ;
	assign v_856 = 0 ;
	assign v_847 = 0 ;
	assign v_838 = 0 ;
	assign v_829 = 0 ;
	assign v_806 = 0 ;
	assign v_783 = 0 ;
	assign v_694 = 0 ;
	assign o_1 = x_4835 ;
endmodule
