// Benchmark "SKOLEMFORMULA" written by ABC on Fri May 27 20:54:56 2022

module SKOLEMFORMULA ( 
    i0, i1,
    i2, i3  );
  input  i0, i1;
  output i2, i3;
  assign i2 = 1'b1;
  assign i3 = i1;
endmodule


