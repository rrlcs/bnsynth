// Verilog file written by procedure writeCombinationalCircuitInVerilog
//Skolem functions to be generated for i_ variables
module formula ( x_0,i_1,i_2,i_3,x_4,x_5,x_6,i_7,i_8,i_9,i_10,i_11,i_12,out);
input x_0;
input i_1;
input i_2;
input i_3;
input x_4;
input x_5;
input x_6;
input i_7;
input i_8;
input i_9;
input i_10;
input i_11;
input i_12;
output out;
wire c1;
assign c1 = x_0 ^ x_5;
wire carry1;
assign carry1 = (x_0 & x_5);
wire c2;
assign c2 = ((carry1 ^ x_4) ^ x_6);
wire carry2;
assign carry2 = (x_4 & x_6) | (carry1 & (x_4 ^ x_6));
wire a1;
assign a1 = ~(c1 ^ i_7);
wire a2;
assign a2 = ~(c2 ^ i_8);
wire a3;
assign a3 = ~(carry2 ^ i_3);
wire c3;
assign c3 = ~i_9;
wire a4;
assign a4 = ~(c3 ^ i_1);
wire c4;
assign c4 = x_0 | i_12 ;
wire a5;
assign a5 = ~(i_10 ^ c4);
wire c5;
assign c5 = x_4 & i_10 ;
wire a6;
assign a6 = ~(i_11 ^ c5);
wire c6;
assign c6 = x_5 | i_11 ;
wire a7;
assign a7 = ~(i_12 ^ c6);
assign out = ((((((a1 & a2) & a3) &a4) & a5) & a6) & a7);
endmodule
