// Benchmark "SKOLEMFORMULA" written by ABC on Fri May 20 19:55:17 2022

module SKOLEMFORMULA ( 
    i0, i1,
    i2  );
  input  i0, i1;
  output i2;
  assign i2 = i0 & i1;
endmodule


