module formula(v_1,v_2,v_3,v_4,v_5,v_6,v_7,v_8,v_9,v_10,v_11,v_12,v_13,v_14,v_15,v_16,v_17,v_18,v_19,v_20,v_21,v_22,v_23,v_24,v_25,v_26,v_27,v_28,v_29,v_30,v_31,v_32,v_33,v_34,v_35,v_36,v_37,v_38,v_39,v_40,v_41,v_42,v_43,v_44,v_45,v_46,v_47,v_48,v_49,v_50,v_51,v_52,v_53,v_54,v_55,v_56,v_57,v_58,v_59,v_60,v_61,v_62,v_63,v_64,v_65,v_66,v_67,v_68,v_69,v_70,v_71,v_72,v_73,v_74,v_75,v_76,v_77,v_78,v_79,v_80,v_81,v_82,v_83,v_84,v_85,v_86,v_87,v_88,v_89,v_90,v_91,v_92,v_93,v_94,v_95,v_96,v_97,v_98,v_99,v_100,v_101,v_102,v_103,v_104,v_105,v_106,v_107,v_108,v_109,v_110,v_111,v_112,v_113,v_114,v_115,v_116,v_117,v_118,v_119,v_120,v_121,v_122,v_123,v_124,v_125,v_126,v_127,v_128,v_129,v_130,v_131,v_132,v_133,v_134,v_135,v_136,v_137,v_138,v_139,v_140,v_141,v_142,v_143,v_144,v_145,v_146,v_147,v_148,v_149,v_150,v_151,v_152,v_153,v_154,v_155,v_156,v_157,v_158,v_159,v_160,v_161,v_162,v_163,v_164,v_165,v_166,v_167,v_168,v_169,v_170,v_171,v_172,v_173,v_174,v_175,v_176,v_177,v_178,v_179,v_180,o_1);
	input v_1;
	input v_2;
	input v_3;
	input v_4;
	input v_5;
	input v_6;
	input v_7;
	input v_8;
	input v_9;
	input v_10;
	input v_11;
	input v_12;
	input v_13;
	input v_14;
	input v_15;
	input v_16;
	input v_17;
	input v_18;
	input v_19;
	input v_20;
	input v_21;
	input v_22;
	input v_23;
	input v_24;
	input v_25;
	input v_26;
	input v_27;
	input v_28;
	input v_29;
	input v_30;
	input v_31;
	input v_32;
	input v_33;
	input v_34;
	input v_35;
	input v_36;
	input v_37;
	input v_38;
	input v_39;
	input v_40;
	input v_41;
	input v_42;
	input v_43;
	input v_44;
	input v_45;
	input v_46;
	input v_47;
	input v_48;
	input v_49;
	input v_50;
	input v_51;
	input v_52;
	input v_53;
	input v_54;
	input v_55;
	input v_56;
	input v_57;
	input v_58;
	input v_59;
	input v_60;
	input v_61;
	input v_62;
	input v_63;
	input v_64;
	input v_65;
	input v_66;
	input v_67;
	input v_68;
	input v_69;
	input v_70;
	input v_71;
	input v_72;
	input v_73;
	input v_74;
	input v_75;
	input v_76;
	input v_77;
	input v_78;
	input v_79;
	input v_80;
	input v_81;
	input v_82;
	input v_83;
	input v_84;
	input v_85;
	input v_86;
	input v_87;
	input v_88;
	input v_89;
	input v_90;
	input v_91;
	input v_92;
	input v_93;
	input v_94;
	input v_95;
	input v_96;
	input v_97;
	input v_98;
	input v_99;
	input v_100;
	input v_101;
	input v_102;
	input v_103;
	input v_104;
	input v_105;
	input v_106;
	input v_107;
	input v_108;
	input v_109;
	input v_110;
	input v_111;
	input v_112;
	input v_113;
	input v_114;
	input v_115;
	input v_116;
	input v_117;
	input v_118;
	input v_119;
	input v_120;
	input v_121;
	input v_122;
	input v_123;
	input v_124;
	input v_125;
	input v_126;
	input v_127;
	input v_128;
	input v_129;
	input v_130;
	input v_131;
	input v_132;
	input v_133;
	input v_134;
	input v_135;
	input v_136;
	input v_137;
	input v_138;
	input v_139;
	input v_140;
	input v_141;
	input v_142;
	input v_143;
	input v_144;
	input v_145;
	input v_146;
	input v_147;
	input v_148;
	input v_149;
	input v_150;
	input v_151;
	input v_152;
	input v_153;
	input v_154;
	input v_155;
	input v_156;
	input v_157;
	input v_158;
	input v_159;
	input v_160;
	input v_161;
	input v_162;
	input v_163;
	input v_164;
	input v_165;
	input v_166;
	input v_167;
	input v_168;
	input v_169;
	input v_170;
	input v_171;
	input v_172;
	input v_173;
	input v_174;
	input v_175;
	input v_176;
	input v_177;
	input v_178;
	input v_179;
	input v_180;
	wire x_1;
	wire x_2;
	wire x_3;
	wire x_4;
	wire x_5;
	wire x_6;
	wire x_7;
	wire x_8;
	wire x_9;
	wire x_10;
	wire x_11;
	wire x_12;
	wire x_13;
	wire x_14;
	wire x_15;
	wire x_16;
	wire x_17;
	wire x_18;
	wire x_19;
	wire x_20;
	wire x_21;
	wire x_22;
	wire x_23;
	wire x_24;
	wire x_25;
	wire x_26;
	wire x_27;
	wire x_28;
	wire x_29;
	wire x_30;
	wire x_31;
	wire x_32;
	wire x_33;
	wire x_34;
	wire x_35;
	wire x_36;
	wire x_37;
	wire x_38;
	wire x_39;
	wire x_40;
	wire x_41;
	wire x_42;
	wire x_43;
	wire x_44;
	wire x_45;
	wire x_46;
	wire x_47;
	wire x_48;
	wire x_49;
	wire x_50;
	wire x_51;
	wire x_52;
	wire x_53;
	wire x_54;
	wire x_55;
	wire x_56;
	wire x_57;
	wire x_58;
	wire x_59;
	wire x_60;
	wire x_61;
	wire x_62;
	wire x_63;
	wire x_64;
	wire x_65;
	wire x_66;
	wire x_67;
	wire x_68;
	wire x_69;
	wire x_70;
	wire x_71;
	wire x_72;
	wire x_73;
	wire x_74;
	wire x_75;
	wire x_76;
	wire x_77;
	wire x_78;
	wire x_79;
	wire x_80;
	wire x_81;
	wire x_82;
	wire x_83;
	wire x_84;
	wire x_85;
	wire x_86;
	wire x_87;
	wire x_88;
	wire x_89;
	wire x_90;
	wire x_91;
	wire x_92;
	wire x_93;
	wire x_94;
	wire x_95;
	wire x_96;
	wire x_97;
	wire x_98;
	wire x_99;
	wire x_100;
	wire x_101;
	wire x_102;
	wire x_103;
	wire x_104;
	wire x_105;
	wire x_106;
	wire x_107;
	wire x_108;
	wire x_109;
	wire x_110;
	wire x_111;
	wire x_112;
	wire x_113;
	wire x_114;
	wire x_115;
	wire x_116;
	wire x_117;
	wire x_118;
	wire x_119;
	wire x_120;
	wire x_121;
	wire x_122;
	wire x_123;
	wire x_124;
	wire x_125;
	wire x_126;
	wire x_127;
	wire x_128;
	wire x_129;
	wire x_130;
	wire x_131;
	wire x_132;
	wire x_133;
	wire x_134;
	wire x_135;
	wire x_136;
	wire x_137;
	wire x_138;
	wire x_139;
	wire x_140;
	wire x_141;
	wire x_142;
	wire x_143;
	wire x_144;
	wire x_145;
	wire x_146;
	wire x_147;
	wire x_148;
	wire x_149;
	wire x_150;
	wire x_151;
	wire x_152;
	wire x_153;
	wire x_154;
	wire x_155;
	wire x_156;
	wire x_157;
	wire x_158;
	wire x_159;
	wire x_160;
	wire x_161;
	wire x_162;
	wire x_163;
	wire x_164;
	wire x_165;
	wire x_166;
	wire x_167;
	wire x_168;
	wire x_169;
	wire x_170;
	wire x_171;
	wire x_172;
	wire x_173;
	wire x_174;
	wire x_175;
	wire x_176;
	wire x_177;
	wire x_178;
	wire x_179;
	wire x_180;
	wire x_181;
	wire x_182;
	wire x_183;
	wire x_184;
	wire x_185;
	wire x_186;
	wire x_187;
	wire x_188;
	wire x_189;
	wire x_190;
	wire x_191;
	wire x_192;
	wire x_193;
	wire x_194;
	wire x_195;
	wire x_196;
	wire x_197;
	wire x_198;
	wire x_199;
	wire x_200;
	wire x_201;
	wire x_202;
	wire x_203;
	wire x_204;
	wire x_205;
	wire x_206;
	wire x_207;
	wire x_208;
	wire x_209;
	wire x_210;
	wire x_211;
	wire x_212;
	wire x_213;
	wire x_214;
	wire x_215;
	wire x_216;
	wire x_217;
	wire x_218;
	wire x_219;
	wire x_220;
	wire x_221;
	wire x_222;
	wire x_223;
	wire x_224;
	wire x_225;
	wire x_226;
	wire x_227;
	wire x_228;
	wire x_229;
	wire x_230;
	wire x_231;
	wire x_232;
	wire x_233;
	wire x_234;
	wire x_235;
	wire x_236;
	wire x_237;
	wire x_238;
	wire x_239;
	wire x_240;
	wire x_241;
	wire x_242;
	wire x_243;
	wire x_244;
	wire x_245;
	wire x_246;
	wire x_247;
	wire x_248;
	wire x_249;
	wire x_250;
	wire x_251;
	wire x_252;
	wire x_253;
	wire x_254;
	wire x_255;
	wire x_256;
	wire x_257;
	wire x_258;
	wire x_259;
	wire x_260;
	wire x_261;
	wire x_262;
	wire x_263;
	wire x_264;
	wire x_265;
	wire x_266;
	wire x_267;
	wire x_268;
	wire x_269;
	wire x_270;
	wire x_271;
	wire x_272;
	wire x_273;
	wire x_274;
	wire x_275;
	wire x_276;
	wire x_277;
	wire x_278;
	wire x_279;
	wire x_280;
	wire x_281;
	wire x_282;
	wire x_283;
	wire x_284;
	wire x_285;
	wire x_286;
	wire x_287;
	wire x_288;
	wire x_289;
	wire x_290;
	wire x_291;
	wire x_292;
	wire x_293;
	wire x_294;
	wire x_295;
	wire x_296;
	wire x_297;
	wire x_298;
	wire x_299;
	wire x_300;
	wire x_301;
	wire x_302;
	wire x_303;
	wire x_304;
	wire x_305;
	wire x_306;
	wire x_307;
	wire x_308;
	wire x_309;
	wire x_310;
	wire x_311;
	wire x_312;
	wire x_313;
	wire x_314;
	wire x_315;
	wire x_316;
	wire x_317;
	wire x_318;
	wire x_319;
	wire x_320;
	wire x_321;
	wire x_322;
	wire x_323;
	wire x_324;
	wire x_325;
	wire x_326;
	wire x_327;
	wire x_328;
	wire x_329;
	wire x_330;
	wire x_331;
	wire x_332;
	wire x_333;
	wire x_334;
	wire x_335;
	wire x_336;
	wire x_337;
	wire x_338;
	wire x_339;
	wire x_340;
	wire x_341;
	wire x_342;
	wire x_343;
	wire x_344;
	wire x_345;
	wire x_346;
	wire x_347;
	wire x_348;
	wire x_349;
	wire x_350;
	wire x_351;
	wire x_352;
	wire x_353;
	wire x_354;
	wire x_355;
	wire x_356;
	wire x_357;
	wire x_358;
	wire x_359;
	wire x_360;
	wire x_361;
	wire x_362;
	wire x_363;
	wire x_364;
	wire x_365;
	wire x_366;
	wire x_367;
	wire x_368;
	wire x_369;
	wire x_370;
	wire x_371;
	wire x_372;
	wire x_373;
	wire x_374;
	wire x_375;
	wire x_376;
	wire x_377;
	wire x_378;
	wire x_379;
	wire x_380;
	wire x_381;
	wire x_382;
	wire x_383;
	wire x_384;
	wire x_385;
	wire x_386;
	wire x_387;
	wire x_388;
	wire x_389;
	wire x_390;
	wire x_391;
	wire x_392;
	wire x_393;
	wire x_394;
	wire x_395;
	wire x_396;
	wire x_397;
	wire x_398;
	wire x_399;
	wire x_400;
	wire x_401;
	wire x_402;
	wire x_403;
	wire x_404;
	wire x_405;
	wire x_406;
	wire x_407;
	wire x_408;
	wire x_409;
	wire x_410;
	wire x_411;
	wire x_412;
	wire x_413;
	wire x_414;
	wire x_415;
	wire x_416;
	wire x_417;
	wire x_418;
	wire x_419;
	wire x_420;
	wire x_421;
	wire x_422;
	wire x_423;
	wire x_424;
	wire x_425;
	wire x_426;
	wire x_427;
	wire x_428;
	wire x_429;
	wire x_430;
	wire x_431;
	wire x_432;
	wire x_433;
	wire x_434;
	wire x_435;
	wire x_436;
	wire x_437;
	wire x_438;
	wire x_439;
	wire x_440;
	wire x_441;
	wire x_442;
	wire x_443;
	wire x_444;
	wire x_445;
	wire x_446;
	wire x_447;
	wire x_448;
	wire x_449;
	wire x_450;
	wire x_451;
	wire x_452;
	wire x_453;
	wire x_454;
	wire x_455;
	wire x_456;
	wire x_457;
	wire x_458;
	wire x_459;
	wire x_460;
	wire x_461;
	wire x_462;
	wire x_463;
	wire x_464;
	wire x_465;
	wire x_466;
	wire x_467;
	wire x_468;
	wire x_469;
	wire x_470;
	wire x_471;
	wire x_472;
	wire x_473;
	wire x_474;
	wire x_475;
	wire x_476;
	wire x_477;
	wire x_478;
	wire x_479;
	wire x_480;
	wire x_481;
	wire x_482;
	wire x_483;
	wire x_484;
	wire x_485;
	wire x_486;
	wire x_487;
	wire x_488;
	wire x_489;
	wire x_490;
	wire x_491;
	wire x_492;
	wire x_493;
	wire x_494;
	wire x_495;
	wire x_496;
	wire x_497;
	wire x_498;
	wire x_499;
	wire x_500;
	wire x_501;
	wire x_502;
	wire x_503;
	wire x_504;
	wire x_505;
	wire x_506;
	wire x_507;
	wire x_508;
	wire x_509;
	wire x_510;
	wire x_511;
	wire x_512;
	wire x_513;
	wire x_514;
	wire x_515;
	wire x_516;
	wire x_517;
	wire x_518;
	wire x_519;
	wire x_520;
	wire x_521;
	wire x_522;
	wire x_523;
	wire x_524;
	wire x_525;
	wire x_526;
	wire x_527;
	wire x_528;
	wire x_529;
	wire x_530;
	wire x_531;
	wire x_532;
	wire x_533;
	wire x_534;
	wire x_535;
	wire x_536;
	wire x_537;
	wire x_538;
	wire x_539;
	wire x_540;
	wire x_541;
	wire x_542;
	wire x_543;
	wire x_544;
	wire x_545;
	wire x_546;
	wire x_547;
	wire x_548;
	wire x_549;
	wire x_550;
	wire x_551;
	wire x_552;
	wire x_553;
	wire x_554;
	wire x_555;
	wire x_556;
	wire x_557;
	wire x_558;
	wire x_559;
	wire x_560;
	wire x_561;
	wire x_562;
	wire x_563;
	wire x_564;
	wire x_565;
	wire x_566;
	wire x_567;
	wire x_568;
	wire x_569;
	wire x_570;
	wire x_571;
	wire x_572;
	wire x_573;
	wire x_574;
	wire x_575;
	wire x_576;
	wire x_577;
	wire x_578;
	wire x_579;
	wire x_580;
	wire x_581;
	wire x_582;
	wire x_583;
	wire x_584;
	wire x_585;
	wire x_586;
	wire x_587;
	wire x_588;
	wire x_589;
	wire x_590;
	wire x_591;
	wire x_592;
	wire x_593;
	wire x_594;
	wire x_595;
	wire x_596;
	wire x_597;
	wire x_598;
	wire x_599;
	wire x_600;
	wire x_601;
	wire x_602;
	wire x_603;
	wire x_604;
	wire x_605;
	wire x_606;
	wire x_607;
	wire x_608;
	wire x_609;
	wire x_610;
	wire x_611;
	wire x_612;
	wire x_613;
	wire x_614;
	wire x_615;
	wire x_616;
	wire x_617;
	wire x_618;
	wire x_619;
	wire x_620;
	wire x_621;
	wire x_622;
	wire x_623;
	wire x_624;
	wire x_625;
	wire x_626;
	wire x_627;
	wire x_628;
	wire x_629;
	wire x_630;
	wire x_631;
	wire x_632;
	wire x_633;
	wire x_634;
	wire x_635;
	wire x_636;
	wire x_637;
	wire x_638;
	wire x_639;
	wire x_640;
	wire x_641;
	wire x_642;
	wire x_643;
	wire x_644;
	wire x_645;
	wire x_646;
	wire x_647;
	wire x_648;
	wire x_649;
	wire x_650;
	wire x_651;
	wire x_652;
	wire x_653;
	wire x_654;
	wire x_655;
	wire x_656;
	wire x_657;
	wire x_658;
	wire x_659;
	wire x_660;
	wire x_661;
	wire x_662;
	wire x_663;
	wire x_664;
	wire x_665;
	wire x_666;
	wire x_667;
	wire x_668;
	wire x_669;
	wire x_670;
	wire x_671;
	wire x_672;
	wire x_673;
	wire x_674;
	wire x_675;
	wire x_676;
	wire x_677;
	wire x_678;
	wire x_679;
	wire x_680;
	wire x_681;
	wire x_682;
	wire x_683;
	wire x_684;
	wire x_685;
	wire x_686;
	wire x_687;
	wire x_688;
	wire x_689;
	wire x_690;
	wire x_691;
	wire x_692;
	wire x_693;
	wire x_694;
	wire x_695;
	wire x_696;
	wire x_697;
	wire x_698;
	wire x_699;
	wire x_700;
	wire x_701;
	wire x_702;
	wire x_703;
	wire x_704;
	wire x_705;
	wire x_706;
	wire x_707;
	wire x_708;
	wire x_709;
	wire x_710;
	wire x_711;
	wire x_712;
	wire x_713;
	wire x_714;
	wire x_715;
	wire x_716;
	wire x_717;
	wire x_718;
	wire x_719;
	wire x_720;
	wire x_721;
	wire x_722;
	wire x_723;
	wire x_724;
	wire x_725;
	wire x_726;
	wire x_727;
	wire x_728;
	wire x_729;
	wire x_730;
	wire x_731;
	wire x_732;
	wire x_733;
	wire x_734;
	wire x_735;
	wire x_736;
	wire x_737;
	wire x_738;
	wire x_739;
	wire x_740;
	wire x_741;
	wire x_742;
	wire x_743;
	wire x_744;
	wire x_745;
	wire x_746;
	wire x_747;
	wire x_748;
	wire x_749;
	wire x_750;
	wire x_751;
	wire x_752;
	wire x_753;
	wire x_754;
	wire x_755;
	wire x_756;
	wire x_757;
	wire x_758;
	wire x_759;
	wire x_760;
	wire x_761;
	wire x_762;
	wire x_763;
	wire x_764;
	wire x_765;
	wire x_766;
	wire x_767;
	wire x_768;
	wire x_769;
	wire x_770;
	wire x_771;
	wire x_772;
	wire x_773;
	wire x_774;
	wire x_775;
	wire x_776;
	wire x_777;
	wire x_778;
	wire x_779;
	wire x_780;
	wire x_781;
	wire x_782;
	wire x_783;
	wire x_784;
	wire x_785;
	wire x_786;
	wire x_787;
	wire x_788;
	wire x_789;
	wire x_790;
	wire x_791;
	wire x_792;
	wire x_793;
	wire x_794;
	wire x_795;
	wire x_796;
	wire x_797;
	wire x_798;
	wire x_799;
	wire x_800;
	wire x_801;
	wire x_802;
	wire x_803;
	wire x_804;
	wire x_805;
	wire x_806;
	wire x_807;
	wire x_808;
	wire x_809;
	wire x_810;
	wire x_811;
	wire x_812;
	wire x_813;
	wire x_814;
	wire x_815;
	wire x_816;
	wire x_817;
	wire x_818;
	wire x_819;
	wire x_820;
	wire x_821;
	wire x_822;
	wire x_823;
	wire x_824;
	wire x_825;
	wire x_826;
	wire x_827;
	wire x_828;
	wire x_829;
	wire x_830;
	wire x_831;
	wire x_832;
	wire x_833;
	wire x_834;
	wire x_835;
	wire x_836;
	wire x_837;
	wire x_838;
	wire x_839;
	wire x_840;
	wire x_841;
	wire x_842;
	wire x_843;
	wire x_844;
	wire x_845;
	wire x_846;
	wire x_847;
	wire x_848;
	wire x_849;
	wire x_850;
	wire x_851;
	wire x_852;
	wire x_853;
	wire x_854;
	wire x_855;
	wire x_856;
	wire x_857;
	wire x_858;
	wire x_859;
	wire x_860;
	wire x_861;
	wire x_862;
	wire x_863;
	wire x_864;
	wire x_865;
	wire x_866;
	wire x_867;
	wire x_868;
	wire x_869;
	wire x_870;
	wire x_871;
	wire x_872;
	wire x_873;
	wire x_874;
	wire x_875;
	wire x_876;
	wire x_877;
	wire x_878;
	wire x_879;
	wire x_880;
	wire x_881;
	wire x_882;
	wire x_883;
	wire x_884;
	wire x_885;
	wire x_886;
	wire x_887;
	wire x_888;
	wire x_889;
	wire x_890;
	wire x_891;
	wire x_892;
	wire x_893;
	wire x_894;
	wire x_895;
	wire x_896;
	wire x_897;
	wire x_898;
	wire x_899;
	wire x_900;
	wire x_901;
	wire x_902;
	wire x_903;
	wire x_904;
	wire x_905;
	wire x_906;
	wire x_907;
	wire x_908;
	wire x_909;
	wire x_910;
	wire x_911;
	wire x_912;
	wire x_913;
	wire x_914;
	wire x_915;
	wire x_916;
	wire x_917;
	wire x_918;
	wire x_919;
	wire x_920;
	wire x_921;
	wire x_922;
	wire x_923;
	wire x_924;
	wire x_925;
	wire x_926;
	wire x_927;
	wire x_928;
	wire x_929;
	wire x_930;
	wire x_931;
	wire x_932;
	wire x_933;
	wire x_934;
	wire x_935;
	wire x_936;
	wire x_937;
	wire x_938;
	wire x_939;
	wire x_940;
	wire x_941;
	wire x_942;
	wire x_943;
	wire x_944;
	wire x_945;
	wire x_946;
	wire x_947;
	wire x_948;
	wire x_949;
	wire x_950;
	wire x_951;
	wire x_952;
	wire x_953;
	wire x_954;
	wire x_955;
	wire x_956;
	wire x_957;
	wire x_958;
	wire x_959;
	wire x_960;
	wire x_961;
	wire x_962;
	wire x_963;
	wire x_964;
	wire x_965;
	wire x_966;
	wire x_967;
	wire x_968;
	wire x_969;
	wire x_970;
	wire x_971;
	wire x_972;
	wire x_973;
	wire x_974;
	wire x_975;
	wire x_976;
	wire x_977;
	wire x_978;
	wire x_979;
	wire x_980;
	wire x_981;
	wire x_982;
	wire x_983;
	wire x_984;
	wire x_985;
	wire x_986;
	wire x_987;
	wire x_988;
	wire x_989;
	wire x_990;
	wire x_991;
	wire x_992;
	wire x_993;
	wire x_994;
	wire x_995;
	wire x_996;
	wire x_997;
	wire x_998;
	wire x_999;
	wire x_1000;
	wire x_1001;
	wire x_1002;
	wire x_1003;
	wire x_1004;
	wire x_1005;
	wire x_1006;
	wire x_1007;
	wire x_1008;
	wire x_1009;
	wire x_1010;
	wire x_1011;
	wire x_1012;
	wire x_1013;
	wire x_1014;
	wire x_1015;
	wire x_1016;
	wire x_1017;
	wire x_1018;
	wire x_1019;
	wire x_1020;
	wire x_1021;
	wire x_1022;
	wire x_1023;
	wire x_1024;
	wire x_1025;
	wire x_1026;
	wire x_1027;
	wire x_1028;
	wire x_1029;
	wire x_1030;
	wire x_1031;
	wire x_1032;
	wire x_1033;
	wire x_1034;
	wire x_1035;
	wire x_1036;
	wire x_1037;
	wire x_1038;
	wire x_1039;
	wire x_1040;
	wire x_1041;
	wire x_1042;
	wire x_1043;
	wire x_1044;
	wire x_1045;
	wire x_1046;
	wire x_1047;
	wire x_1048;
	wire x_1049;
	wire x_1050;
	wire x_1051;
	wire x_1052;
	wire x_1053;
	wire x_1054;
	wire x_1055;
	wire x_1056;
	wire x_1057;
	wire x_1058;
	wire x_1059;
	wire x_1060;
	wire x_1061;
	wire x_1062;
	wire x_1063;
	wire x_1064;
	wire x_1065;
	wire x_1066;
	wire x_1067;
	wire x_1068;
	wire x_1069;
	wire x_1070;
	wire x_1071;
	wire x_1072;
	wire x_1073;
	wire x_1074;
	wire x_1075;
	wire x_1076;
	wire x_1077;
	wire x_1078;
	wire x_1079;
	wire x_1080;
	wire x_1081;
	wire x_1082;
	wire x_1083;
	wire x_1084;
	wire x_1085;
	wire x_1086;
	wire x_1087;
	wire x_1088;
	wire x_1089;
	wire x_1090;
	wire x_1091;
	wire x_1092;
	wire x_1093;
	wire x_1094;
	wire x_1095;
	wire x_1096;
	wire x_1097;
	wire x_1098;
	wire x_1099;
	wire x_1100;
	wire x_1101;
	wire x_1102;
	wire x_1103;
	wire x_1104;
	wire x_1105;
	wire x_1106;
	wire x_1107;
	wire x_1108;
	wire x_1109;
	wire x_1110;
	wire x_1111;
	wire x_1112;
	wire x_1113;
	wire x_1114;
	wire x_1115;
	wire x_1116;
	wire x_1117;
	wire x_1118;
	wire x_1119;
	wire x_1120;
	wire x_1121;
	wire x_1122;
	wire x_1123;
	wire x_1124;
	wire x_1125;
	wire x_1126;
	wire x_1127;
	wire x_1128;
	wire x_1129;
	wire x_1130;
	wire x_1131;
	wire x_1132;
	wire x_1133;
	wire x_1134;
	wire x_1135;
	wire x_1136;
	wire x_1137;
	wire x_1138;
	wire x_1139;
	wire x_1140;
	wire x_1141;
	wire x_1142;
	wire x_1143;
	wire x_1144;
	wire x_1145;
	wire x_1146;
	wire x_1147;
	wire x_1148;
	wire x_1149;
	wire x_1150;
	wire x_1151;
	wire x_1152;
	wire x_1153;
	wire x_1154;
	wire x_1155;
	wire x_1156;
	wire x_1157;
	wire x_1158;
	wire x_1159;
	wire x_1160;
	wire x_1161;
	wire x_1162;
	wire x_1163;
	wire x_1164;
	wire x_1165;
	wire x_1166;
	wire x_1167;
	wire x_1168;
	wire x_1169;
	wire x_1170;
	wire x_1171;
	wire x_1172;
	wire x_1173;
	wire x_1174;
	wire x_1175;
	wire x_1176;
	wire x_1177;
	wire x_1178;
	wire x_1179;
	wire x_1180;
	wire x_1181;
	wire x_1182;
	wire x_1183;
	wire x_1184;
	wire x_1185;
	wire x_1186;
	wire x_1187;
	wire x_1188;
	wire x_1189;
	wire x_1190;
	wire x_1191;
	wire x_1192;
	wire x_1193;
	wire x_1194;
	wire x_1195;
	wire x_1196;
	wire x_1197;
	wire x_1198;
	wire x_1199;
	wire x_1200;
	wire x_1201;
	wire x_1202;
	wire x_1203;
	wire x_1204;
	wire x_1205;
	wire x_1206;
	wire x_1207;
	wire x_1208;
	wire x_1209;
	wire x_1210;
	wire x_1211;
	wire x_1212;
	wire x_1213;
	wire x_1214;
	wire x_1215;
	wire x_1216;
	wire x_1217;
	wire x_1218;
	wire x_1219;
	wire x_1220;
	wire x_1221;
	wire x_1222;
	wire x_1223;
	wire x_1224;
	wire x_1225;
	wire x_1226;
	wire x_1227;
	wire x_1228;
	wire x_1229;
	wire x_1230;
	wire x_1231;
	wire x_1232;
	wire x_1233;
	wire x_1234;
	wire x_1235;
	wire x_1236;
	wire x_1237;
	wire x_1238;
	wire x_1239;
	wire x_1240;
	wire x_1241;
	wire x_1242;
	wire x_1243;
	wire x_1244;
	wire x_1245;
	wire x_1246;
	wire x_1247;
	wire x_1248;
	wire x_1249;
	wire x_1250;
	wire x_1251;
	wire x_1252;
	wire x_1253;
	wire x_1254;
	wire x_1255;
	wire x_1256;
	wire x_1257;
	wire x_1258;
	wire x_1259;
	wire x_1260;
	wire x_1261;
	wire x_1262;
	wire x_1263;
	wire x_1264;
	wire x_1265;
	wire x_1266;
	wire x_1267;
	wire x_1268;
	wire x_1269;
	wire x_1270;
	wire x_1271;
	wire x_1272;
	wire x_1273;
	wire x_1274;
	wire x_1275;
	wire x_1276;
	wire x_1277;
	wire x_1278;
	wire x_1279;
	wire x_1280;
	wire x_1281;
	wire x_1282;
	wire x_1283;
	wire x_1284;
	wire x_1285;
	wire x_1286;
	wire x_1287;
	wire x_1288;
	wire x_1289;
	wire x_1290;
	wire x_1291;
	wire x_1292;
	wire x_1293;
	wire x_1294;
	wire x_1295;
	wire x_1296;
	wire x_1297;
	wire x_1298;
	wire x_1299;
	wire x_1300;
	wire x_1301;
	wire x_1302;
	wire x_1303;
	wire x_1304;
	wire x_1305;
	wire x_1306;
	wire x_1307;
	wire x_1308;
	wire x_1309;
	wire x_1310;
	wire x_1311;
	wire x_1312;
	wire x_1313;
	wire x_1314;
	wire x_1315;
	wire x_1316;
	wire x_1317;
	wire x_1318;
	wire x_1319;
	wire x_1320;
	wire x_1321;
	wire x_1322;
	wire x_1323;
	wire x_1324;
	wire x_1325;
	wire x_1326;
	wire x_1327;
	wire x_1328;
	wire x_1329;
	wire x_1330;
	wire x_1331;
	wire x_1332;
	wire x_1333;
	wire x_1334;
	wire x_1335;
	wire x_1336;
	wire x_1337;
	wire x_1338;
	wire x_1339;
	wire x_1340;
	wire x_1341;
	wire x_1342;
	wire x_1343;
	wire x_1344;
	wire x_1345;
	wire x_1346;
	wire x_1347;
	wire x_1348;
	wire x_1349;
	wire x_1350;
	wire x_1351;
	wire x_1352;
	wire x_1353;
	wire x_1354;
	wire x_1355;
	wire x_1356;
	wire x_1357;
	wire x_1358;
	wire x_1359;
	wire x_1360;
	wire x_1361;
	wire x_1362;
	wire x_1363;
	wire x_1364;
	wire x_1365;
	wire x_1366;
	wire x_1367;
	wire x_1368;
	wire x_1369;
	wire x_1370;
	wire x_1371;
	wire x_1372;
	wire x_1373;
	wire x_1374;
	wire x_1375;
	wire x_1376;
	wire x_1377;
	wire x_1378;
	wire x_1379;
	wire x_1380;
	wire x_1381;
	wire x_1382;
	wire x_1383;
	wire x_1384;
	wire x_1385;
	wire x_1386;
	wire x_1387;
	wire x_1388;
	wire x_1389;
	wire x_1390;
	wire x_1391;
	wire x_1392;
	wire x_1393;
	wire x_1394;
	wire x_1395;
	wire x_1396;
	wire x_1397;
	wire x_1398;
	wire x_1399;
	wire x_1400;
	wire x_1401;
	wire x_1402;
	wire x_1403;
	wire x_1404;
	wire x_1405;
	wire x_1406;
	wire x_1407;
	wire x_1408;
	wire x_1409;
	wire x_1410;
	wire x_1411;
	wire x_1412;
	wire x_1413;
	wire x_1414;
	wire x_1415;
	wire x_1416;
	wire x_1417;
	wire x_1418;
	wire x_1419;
	wire x_1420;
	wire x_1421;
	wire x_1422;
	wire x_1423;
	wire x_1424;
	wire x_1425;
	wire x_1426;
	wire x_1427;
	wire x_1428;
	wire x_1429;
	wire x_1430;
	wire x_1431;
	wire x_1432;
	wire x_1433;
	wire x_1434;
	wire x_1435;
	wire x_1436;
	wire x_1437;
	wire x_1438;
	wire x_1439;
	wire x_1440;
	wire x_1441;
	wire x_1442;
	wire x_1443;
	wire x_1444;
	wire x_1445;
	wire x_1446;
	wire x_1447;
	wire x_1448;
	wire x_1449;
	wire x_1450;
	wire x_1451;
	wire x_1452;
	wire x_1453;
	wire x_1454;
	wire x_1455;
	wire x_1456;
	wire x_1457;
	wire x_1458;
	wire x_1459;
	wire x_1460;
	wire x_1461;
	wire x_1462;
	wire x_1463;
	wire x_1464;
	wire x_1465;
	wire x_1466;
	wire x_1467;
	wire x_1468;
	wire x_1469;
	wire x_1470;
	wire x_1471;
	wire x_1472;
	wire x_1473;
	wire x_1474;
	wire x_1475;
	wire x_1476;
	wire x_1477;
	wire x_1478;
	wire x_1479;
	wire x_1480;
	wire x_1481;
	wire x_1482;
	wire x_1483;
	wire x_1484;
	wire x_1485;
	wire x_1486;
	wire x_1487;
	wire x_1488;
	wire x_1489;
	wire x_1490;
	wire x_1491;
	wire x_1492;
	wire x_1493;
	wire x_1494;
	wire x_1495;
	wire x_1496;
	wire x_1497;
	wire x_1498;
	wire x_1499;
	wire x_1500;
	wire x_1501;
	wire x_1502;
	wire x_1503;
	wire x_1504;
	wire x_1505;
	wire x_1506;
	wire x_1507;
	wire x_1508;
	wire x_1509;
	wire x_1510;
	wire x_1511;
	wire x_1512;
	wire x_1513;
	wire x_1514;
	wire x_1515;
	wire x_1516;
	wire x_1517;
	wire x_1518;
	wire x_1519;
	wire x_1520;
	wire x_1521;
	wire x_1522;
	wire x_1523;
	wire x_1524;
	wire x_1525;
	wire x_1526;
	wire x_1527;
	wire x_1528;
	wire x_1529;
	wire x_1530;
	wire x_1531;
	wire x_1532;
	wire x_1533;
	wire x_1534;
	wire x_1535;
	wire x_1536;
	wire x_1537;
	wire x_1538;
	wire x_1539;
	wire x_1540;
	wire x_1541;
	wire x_1542;
	wire x_1543;
	wire x_1544;
	wire x_1545;
	wire x_1546;
	wire x_1547;
	wire x_1548;
	wire x_1549;
	wire x_1550;
	wire x_1551;
	wire x_1552;
	wire x_1553;
	wire x_1554;
	wire x_1555;
	wire x_1556;
	wire x_1557;
	wire x_1558;
	wire x_1559;
	wire x_1560;
	wire x_1561;
	wire x_1562;
	wire x_1563;
	wire x_1564;
	wire x_1565;
	wire x_1566;
	wire x_1567;
	wire x_1568;
	wire x_1569;
	wire x_1570;
	wire x_1571;
	wire x_1572;
	wire x_1573;
	wire x_1574;
	wire x_1575;
	wire x_1576;
	wire x_1577;
	wire x_1578;
	wire x_1579;
	wire x_1580;
	wire x_1581;
	wire x_1582;
	wire x_1583;
	wire x_1584;
	wire x_1585;
	wire x_1586;
	wire x_1587;
	wire x_1588;
	wire x_1589;
	wire x_1590;
	wire x_1591;
	wire x_1592;
	wire x_1593;
	wire x_1594;
	wire x_1595;
	wire x_1596;
	wire x_1597;
	wire x_1598;
	wire x_1599;
	wire x_1600;
	wire x_1601;
	wire x_1602;
	wire x_1603;
	wire x_1604;
	wire x_1605;
	wire x_1606;
	wire x_1607;
	wire x_1608;
	wire x_1609;
	wire x_1610;
	wire x_1611;
	wire x_1612;
	wire x_1613;
	wire x_1614;
	wire x_1615;
	wire x_1616;
	wire x_1617;
	wire x_1618;
	wire x_1619;
	wire x_1620;
	wire x_1621;
	wire x_1622;
	wire x_1623;
	wire x_1624;
	wire x_1625;
	wire x_1626;
	wire x_1627;
	wire x_1628;
	wire x_1629;
	wire x_1630;
	wire x_1631;
	wire x_1632;
	wire x_1633;
	wire x_1634;
	wire x_1635;
	wire x_1636;
	wire x_1637;
	wire x_1638;
	wire x_1639;
	wire x_1640;
	wire x_1641;
	wire x_1642;
	wire x_1643;
	wire x_1644;
	wire x_1645;
	wire x_1646;
	wire x_1647;
	wire x_1648;
	wire x_1649;
	wire x_1650;
	wire x_1651;
	wire x_1652;
	wire x_1653;
	wire x_1654;
	wire x_1655;
	wire x_1656;
	wire x_1657;
	wire x_1658;
	wire x_1659;
	wire x_1660;
	wire x_1661;
	wire x_1662;
	wire x_1663;
	wire x_1664;
	wire x_1665;
	wire x_1666;
	wire x_1667;
	wire x_1668;
	wire x_1669;
	wire x_1670;
	wire x_1671;
	wire x_1672;
	wire x_1673;
	wire x_1674;
	wire x_1675;
	wire x_1676;
	wire x_1677;
	wire x_1678;
	wire x_1679;
	wire x_1680;
	wire x_1681;
	wire x_1682;
	wire x_1683;
	wire x_1684;
	wire x_1685;
	wire x_1686;
	wire x_1687;
	wire x_1688;
	wire x_1689;
	wire x_1690;
	wire x_1691;
	wire x_1692;
	wire x_1693;
	wire x_1694;
	wire x_1695;
	wire x_1696;
	wire x_1697;
	wire x_1698;
	wire x_1699;
	wire x_1700;
	wire x_1701;
	wire x_1702;
	wire x_1703;
	wire x_1704;
	wire x_1705;
	wire x_1706;
	wire x_1707;
	wire x_1708;
	wire x_1709;
	wire x_1710;
	wire x_1711;
	wire x_1712;
	wire x_1713;
	wire x_1714;
	wire x_1715;
	wire x_1716;
	wire x_1717;
	wire x_1718;
	wire x_1719;
	wire x_1720;
	wire x_1721;
	wire x_1722;
	wire x_1723;
	wire x_1724;
	wire x_1725;
	wire x_1726;
	wire x_1727;
	wire x_1728;
	wire x_1729;
	wire x_1730;
	wire x_1731;
	wire x_1732;
	wire x_1733;
	wire x_1734;
	wire x_1735;
	wire x_1736;
	wire x_1737;
	wire x_1738;
	wire x_1739;
	wire x_1740;
	wire x_1741;
	wire x_1742;
	wire x_1743;
	wire x_1744;
	wire x_1745;
	wire x_1746;
	wire x_1747;
	wire x_1748;
	wire x_1749;
	wire x_1750;
	wire x_1751;
	wire x_1752;
	wire x_1753;
	wire x_1754;
	wire x_1755;
	wire x_1756;
	wire x_1757;
	wire x_1758;
	wire x_1759;
	wire x_1760;
	wire x_1761;
	wire x_1762;
	wire x_1763;
	wire x_1764;
	wire x_1765;
	wire x_1766;
	wire x_1767;
	wire x_1768;
	wire x_1769;
	wire x_1770;
	wire x_1771;
	wire x_1772;
	wire x_1773;
	wire x_1774;
	wire x_1775;
	wire x_1776;
	wire x_1777;
	wire x_1778;
	wire x_1779;
	wire x_1780;
	wire x_1781;
	wire x_1782;
	wire x_1783;
	wire x_1784;
	wire x_1785;
	wire x_1786;
	wire x_1787;
	wire x_1788;
	wire x_1789;
	wire x_1790;
	wire x_1791;
	wire x_1792;
	wire x_1793;
	wire x_1794;
	wire x_1795;
	wire x_1796;
	wire x_1797;
	wire x_1798;
	wire x_1799;
	wire x_1800;
	wire x_1801;
	wire x_1802;
	wire x_1803;
	wire x_1804;
	wire x_1805;
	wire x_1806;
	wire x_1807;
	wire x_1808;
	wire x_1809;
	wire x_1810;
	wire x_1811;
	wire x_1812;
	wire x_1813;
	wire x_1814;
	wire x_1815;
	wire x_1816;
	wire x_1817;
	wire x_1818;
	wire x_1819;
	wire x_1820;
	wire x_1821;
	wire x_1822;
	wire x_1823;
	wire x_1824;
	wire x_1825;
	wire x_1826;
	wire x_1827;
	wire x_1828;
	wire x_1829;
	wire x_1830;
	wire x_1831;
	wire x_1832;
	wire x_1833;
	wire x_1834;
	wire x_1835;
	wire x_1836;
	wire x_1837;
	wire x_1838;
	wire x_1839;
	wire x_1840;
	wire x_1841;
	wire x_1842;
	wire x_1843;
	wire x_1844;
	wire x_1845;
	wire x_1846;
	wire x_1847;
	wire x_1848;
	wire x_1849;
	wire x_1850;
	wire x_1851;
	wire x_1852;
	wire x_1853;
	wire x_1854;
	wire x_1855;
	wire x_1856;
	wire x_1857;
	wire x_1858;
	wire x_1859;
	wire x_1860;
	wire x_1861;
	wire x_1862;
	wire x_1863;
	wire x_1864;
	wire x_1865;
	wire x_1866;
	wire x_1867;
	wire x_1868;
	wire x_1869;
	wire x_1870;
	wire x_1871;
	wire x_1872;
	wire x_1873;
	wire x_1874;
	wire x_1875;
	wire x_1876;
	wire x_1877;
	wire x_1878;
	wire x_1879;
	wire x_1880;
	wire x_1881;
	wire x_1882;
	wire x_1883;
	wire x_1884;
	wire x_1885;
	wire x_1886;
	wire x_1887;
	wire x_1888;
	wire x_1889;
	wire x_1890;
	wire x_1891;
	wire x_1892;
	wire x_1893;
	wire x_1894;
	wire x_1895;
	wire x_1896;
	wire x_1897;
	wire x_1898;
	wire x_1899;
	wire x_1900;
	wire x_1901;
	wire x_1902;
	wire x_1903;
	wire x_1904;
	wire x_1905;
	wire x_1906;
	wire x_1907;
	wire x_1908;
	wire x_1909;
	wire x_1910;
	wire x_1911;
	wire x_1912;
	wire x_1913;
	wire x_1914;
	wire x_1915;
	wire x_1916;
	wire x_1917;
	wire x_1918;
	wire x_1919;
	wire x_1920;
	wire x_1921;
	wire x_1922;
	wire x_1923;
	wire x_1924;
	wire x_1925;
	wire x_1926;
	wire x_1927;
	wire x_1928;
	wire x_1929;
	wire x_1930;
	wire x_1931;
	wire x_1932;
	wire x_1933;
	wire x_1934;
	wire x_1935;
	wire x_1936;
	wire x_1937;
	wire x_1938;
	wire x_1939;
	wire x_1940;
	wire x_1941;
	wire x_1942;
	wire x_1943;
	wire x_1944;
	wire x_1945;
	wire x_1946;
	wire x_1947;
	wire x_1948;
	wire x_1949;
	wire x_1950;
	wire x_1951;
	wire x_1952;
	wire x_1953;
	wire x_1954;
	wire x_1955;
	wire x_1956;
	wire x_1957;
	wire x_1958;
	wire x_1959;
	wire x_1960;
	wire x_1961;
	wire x_1962;
	wire x_1963;
	wire x_1964;
	wire x_1965;
	wire x_1966;
	wire x_1967;
	wire x_1968;
	wire x_1969;
	wire x_1970;
	wire x_1971;
	wire x_1972;
	wire x_1973;
	wire x_1974;
	wire x_1975;
	wire x_1976;
	wire x_1977;
	wire x_1978;
	wire x_1979;
	wire x_1980;
	wire x_1981;
	wire x_1982;
	wire x_1983;
	wire x_1984;
	wire x_1985;
	wire x_1986;
	wire x_1987;
	wire x_1988;
	wire x_1989;
	wire x_1990;
	wire x_1991;
	wire x_1992;
	wire x_1993;
	wire x_1994;
	wire x_1995;
	wire x_1996;
	wire x_1997;
	wire x_1998;
	wire x_1999;
	wire x_2000;
	wire x_2001;
	wire x_2002;
	wire x_2003;
	wire x_2004;
	wire x_2005;
	wire x_2006;
	wire x_2007;
	wire x_2008;
	wire x_2009;
	wire x_2010;
	wire x_2011;
	wire x_2012;
	wire x_2013;
	wire x_2014;
	wire x_2015;
	wire x_2016;
	wire x_2017;
	wire x_2018;
	wire x_2019;
	wire x_2020;
	wire x_2021;
	wire x_2022;
	wire x_2023;
	wire x_2024;
	wire x_2025;
	wire x_2026;
	wire x_2027;
	wire x_2028;
	wire x_2029;
	wire x_2030;
	wire x_2031;
	wire x_2032;
	wire x_2033;
	wire x_2034;
	wire x_2035;
	wire x_2036;
	wire x_2037;
	wire x_2038;
	wire x_2039;
	wire x_2040;
	wire x_2041;
	wire x_2042;
	wire x_2043;
	wire x_2044;
	wire x_2045;
	wire x_2046;
	wire x_2047;
	wire x_2048;
	wire x_2049;
	wire x_2050;
	wire x_2051;
	wire x_2052;
	wire x_2053;
	wire x_2054;
	wire x_2055;
	wire x_2056;
	wire x_2057;
	wire x_2058;
	wire x_2059;
	wire x_2060;
	wire x_2061;
	wire x_2062;
	wire x_2063;
	wire x_2064;
	wire x_2065;
	wire x_2066;
	wire x_2067;
	wire x_2068;
	wire x_2069;
	wire x_2070;
	wire x_2071;
	wire x_2072;
	wire x_2073;
	wire x_2074;
	wire x_2075;
	wire x_2076;
	wire x_2077;
	wire x_2078;
	wire x_2079;
	wire x_2080;
	wire x_2081;
	wire x_2082;
	wire x_2083;
	wire x_2084;
	wire x_2085;
	wire x_2086;
	wire x_2087;
	wire x_2088;
	wire x_2089;
	wire x_2090;
	wire x_2091;
	wire x_2092;
	wire x_2093;
	wire x_2094;
	wire x_2095;
	wire x_2096;
	wire x_2097;
	wire x_2098;
	wire x_2099;
	wire x_2100;
	wire x_2101;
	wire x_2102;
	wire x_2103;
	wire x_2104;
	wire x_2105;
	wire x_2106;
	wire x_2107;
	wire x_2108;
	wire x_2109;
	wire x_2110;
	wire x_2111;
	wire x_2112;
	wire x_2113;
	wire x_2114;
	wire x_2115;
	wire x_2116;
	wire x_2117;
	wire x_2118;
	wire x_2119;
	wire x_2120;
	wire x_2121;
	wire x_2122;
	wire x_2123;
	wire x_2124;
	wire x_2125;
	wire x_2126;
	wire x_2127;
	wire x_2128;
	wire x_2129;
	wire x_2130;
	wire x_2131;
	wire x_2132;
	wire x_2133;
	wire x_2134;
	wire x_2135;
	wire x_2136;
	wire x_2137;
	wire x_2138;
	wire x_2139;
	wire x_2140;
	wire x_2141;
	wire x_2142;
	wire x_2143;
	wire x_2144;
	wire x_2145;
	wire x_2146;
	wire x_2147;
	wire x_2148;
	wire x_2149;
	wire x_2150;
	wire x_2151;
	wire x_2152;
	wire x_2153;
	wire x_2154;
	wire x_2155;
	wire x_2156;
	wire x_2157;
	wire x_2158;
	wire x_2159;
	wire x_2160;
	wire x_2161;
	wire x_2162;
	wire x_2163;
	wire x_2164;
	wire x_2165;
	wire x_2166;
	wire x_2167;
	wire x_2168;
	wire x_2169;
	wire x_2170;
	wire x_2171;
	wire x_2172;
	wire x_2173;
	wire x_2174;
	wire x_2175;
	wire x_2176;
	wire x_2177;
	wire x_2178;
	wire x_2179;
	wire x_2180;
	wire x_2181;
	wire x_2182;
	wire x_2183;
	wire x_2184;
	wire x_2185;
	wire x_2186;
	wire x_2187;
	wire x_2188;
	wire x_2189;
	wire x_2190;
	wire x_2191;
	wire x_2192;
	wire x_2193;
	wire x_2194;
	wire x_2195;
	wire x_2196;
	wire x_2197;
	wire x_2198;
	wire x_2199;
	output o_1;
	assign x_1100 = ((((~v_38 | v_80) | ~v_152) | v_165) | ~v_114) ;
	assign x_1099 = ((((v_53 | v_30) | v_161) | v_170) | v_139) ;
	assign x_1091 = ((((v_36 | ~v_71) | v_136) | ~v_127) | ~v_118) ;
	assign x_1090 = ((((~v_18 | v_27) | v_101) | v_178) | ~v_156) ;
	assign x_1082 = ((((~v_60 | v_33) | v_162) | v_126) | v_155) ;
	assign x_1081 = ((((~v_6 | v_80) | v_173) | v_163) | v_132) ;
	assign x_1065 = ((((~v_52 | v_18) | v_131) | v_124) | ~v_160) ;
	assign x_1064 = ((((~v_10 | v_77) | v_93) | ~v_96) | v_92) ;
	assign x_1048 = ((((v_50 | ~v_47) | ~v_121) | ~v_158) | v_111) ;
	assign x_1047 = ((((~v_51 | v_73) | ~v_139) | v_122) | v_175) ;
	assign x_1031 = ((((v_61 | ~v_41) | ~v_136) | ~v_135) | ~v_137) ;
	assign x_1030 = ((((~v_9 | v_80) | ~v_160) | v_121) | v_120) ;
	assign x_1022 = ((((v_1 | ~v_73) | ~v_136) | ~v_157) | ~v_178) ;
	assign x_1021 = ((((~v_2 | ~v_25) | ~v_167) | ~v_82) | ~v_112) ;
	assign x_1013 = ((((v_42 | v_52) | ~v_148) | v_145) | v_169) ;
	assign x_1012 = ((((v_20 | v_50) | ~v_83) | v_166) | ~v_89) ;
	assign x_996 = ((((~v_76 | ~v_44) | ~v_157) | v_97) | v_121) ;
	assign x_995 = ((((~v_16 | v_73) | ~v_119) | v_109) | v_180) ;
	assign x_979 = ((((v_31 | ~v_78) | v_106) | v_81) | v_91) ;
	assign x_978 = ((((~v_2 | v_49) | ~v_89) | ~v_115) | v_140) ;
	assign x_962 = ((((v_56 | v_58) | ~v_169) | v_116) | ~v_126) ;
	assign x_961 = ((((v_34 | v_76) | v_122) | ~v_104) | ~v_125) ;
	assign x_953 = ((((~v_42 | ~v_75) | ~v_141) | v_125) | v_180) ;
	assign x_952 = ((((v_71 | v_79) | ~v_160) | v_93) | ~v_127) ;
	assign x_944 = ((((~v_29 | v_40) | ~v_89) | v_90) | ~v_178) ;
	assign x_943 = ((((~v_34 | ~v_80) | ~v_140) | v_146) | v_150) ;
	assign x_927 = ((((~v_47 | ~v_18) | v_109) | ~v_118) | ~v_85) ;
	assign x_926 = ((((~v_21 | ~v_71) | ~v_127) | v_176) | ~v_108) ;
	assign x_910 = ((((~v_20 | ~v_39) | ~v_167) | ~v_121) | ~v_123) ;
	assign x_909 = ((((v_19 | ~v_20) | ~v_86) | ~v_125) | ~v_108) ;
	assign x_893 = ((((~v_60 | v_26) | ~v_92) | ~v_127) | v_134) ;
	assign x_892 = ((((~v_60 | ~v_36) | v_88) | v_105) | ~v_94) ;
	assign x_876 = ((((~v_71 | v_23) | ~v_98) | v_111) | ~v_127) ;
	assign x_875 = ((((v_60 | v_15) | v_168) | v_102) | ~v_94) ;
	assign x_859 = ((((~v_63 | ~v_69) | v_145) | v_137) | v_95) ;
	assign x_858 = ((((v_64 | v_18) | ~v_81) | v_139) | ~v_133) ;
	assign x_842 = ((((v_25 | ~v_34) | v_136) | ~v_179) | v_141) ;
	assign x_841 = ((((v_26 | v_36) | ~v_93) | v_175) | ~v_125) ;
	assign x_825 = ((((~v_56 | ~v_59) | v_146) | ~v_84) | ~v_147) ;
	assign x_824 = ((((~v_59 | v_54) | ~v_84) | v_140) | v_82) ;
	assign x_816 = ((((~v_63 | v_8) | ~v_148) | v_179) | v_94) ;
	assign x_815 = ((((~v_33 | v_29) | ~v_170) | ~v_86) | ~v_136) ;
	assign x_807 = ((((~v_70 | v_10) | v_109) | v_153) | ~v_151) ;
	assign x_806 = ((((v_47 | v_61) | v_163) | ~v_149) | v_173) ;
	assign x_790 = ((((~v_12 | v_56) | ~v_97) | ~v_154) | v_139) ;
	assign x_789 = ((((~v_70 | ~v_65) | v_134) | ~v_137) | ~v_85) ;
	assign x_773 = ((((~v_44 | v_18) | v_87) | v_154) | ~v_156) ;
	assign x_772 = ((((v_53 | v_5) | v_105) | ~v_112) | v_147) ;
	assign x_756 = ((((~v_3 | ~v_48) | v_157) | v_173) | v_154) ;
	assign x_755 = ((((v_57 | v_9) | v_152) | ~v_140) | ~v_132) ;
	assign x_747 = ((((~v_54 | v_18) | v_156) | ~v_155) | ~v_146) ;
	assign x_746 = ((((~v_20 | v_8) | v_127) | ~v_170) | ~v_82) ;
	assign x_738 = ((((~v_15 | v_9) | v_161) | ~v_120) | ~v_168) ;
	assign x_737 = ((((v_61 | v_78) | v_97) | v_176) | v_147) ;
	assign x_721 = ((((~v_67 | ~v_56) | ~v_178) | v_130) | ~v_93) ;
	assign x_720 = ((((~v_28 | v_18) | ~v_113) | ~v_121) | v_132) ;
	assign x_704 = ((((~v_20 | v_13) | v_136) | v_147) | v_124) ;
	assign x_703 = ((((~v_61 | v_3) | ~v_100) | ~v_120) | v_145) ;
	assign x_687 = ((((v_75 | v_32) | v_136) | ~v_155) | ~v_142) ;
	assign x_686 = ((((~v_30 | v_16) | v_131) | ~v_142) | ~v_101) ;
	assign x_678 = ((((~v_68 | v_69) | ~v_112) | v_133) | v_114) ;
	assign x_677 = ((((~v_33 | v_51) | v_144) | ~v_103) | v_113) ;
	assign x_669 = ((((~v_5 | v_18) | v_118) | v_169) | ~v_153) ;
	assign x_668 = ((((~v_35 | ~v_24) | v_142) | v_171) | ~v_143) ;
	assign x_652 = ((((~v_44 | v_60) | ~v_162) | v_146) | v_159) ;
	assign x_651 = ((((~v_23 | v_38) | v_155) | ~v_97) | ~v_168) ;
	assign x_635 = ((((~v_13 | v_14) | ~v_121) | ~v_134) | ~v_168) ;
	assign x_634 = ((((~v_77 | v_50) | ~v_160) | ~v_144) | ~v_133) ;
	assign x_618 = ((((v_56 | v_69) | v_120) | ~v_143) | ~v_162) ;
	assign x_617 = ((((~v_75 | ~v_41) | ~v_114) | ~v_85) | ~v_105) ;
	assign x_601 = ((((~v_40 | ~v_5) | ~v_168) | ~v_145) | v_130) ;
	assign x_600 = ((((~v_25 | ~v_10) | ~v_164) | ~v_95) | ~v_129) ;
	assign x_584 = ((((v_48 | v_6) | ~v_83) | v_146) | ~v_131) ;
	assign x_583 = ((((~v_35 | ~v_32) | v_143) | ~v_105) | ~v_101) ;
	assign x_567 = ((((v_24 | v_7) | ~v_158) | ~v_105) | v_101) ;
	assign x_566 = ((((~v_64 | v_49) | ~v_164) | v_156) | ~v_179) ;
	assign x_550 = ((((~v_17 | ~v_44) | v_99) | v_101) | ~v_138) ;
	assign x_549 = ((((~v_21 | ~v_67) | v_175) | ~v_87) | ~v_85) ;
	assign x_541 = ((((v_14 | v_47) | ~v_128) | v_121) | v_98) ;
	assign x_540 = ((((~v_1 | v_49) | ~v_137) | ~v_120) | v_92) ;
	assign x_532 = ((((~v_48 | ~v_35) | ~v_87) | v_172) | v_178) ;
	assign x_531 = ((((v_52 | ~v_74) | ~v_173) | ~v_146) | v_169) ;
	assign x_515 = ((((v_40 | v_3) | ~v_155) | ~v_98) | v_93) ;
	assign x_514 = ((((v_52 | ~v_61) | ~v_115) | ~v_142) | v_82) ;
	assign x_498 = ((((~v_6 | ~v_57) | ~v_119) | ~v_84) | ~v_124) ;
	assign x_497 = ((((~v_37 | ~v_3) | v_144) | v_136) | v_92) ;
	assign x_481 = ((((v_15 | ~v_65) | v_159) | v_130) | v_168) ;
	assign x_480 = ((((v_55 | ~v_28) | ~v_113) | v_89) | v_167) ;
	assign x_472 = ((((~v_76 | ~v_38) | ~v_131) | ~v_153) | v_134) ;
	assign x_471 = ((((~v_70 | ~v_57) | ~v_165) | v_172) | ~v_134) ;
	assign x_463 = ((((~v_11 | ~v_42) | ~v_159) | v_136) | ~v_113) ;
	assign x_462 = ((((v_28 | v_56) | v_102) | v_167) | ~v_96) ;
	assign x_446 = ((((~v_43 | v_73) | ~v_170) | v_167) | v_83) ;
	assign x_445 = ((((v_5 | ~v_18) | v_94) | ~v_132) | ~v_162) ;
	assign x_429 = ((((v_33 | ~v_16) | v_164) | ~v_152) | v_158) ;
	assign x_428 = ((((v_4 | v_70) | ~v_101) | ~v_90) | ~v_123) ;
	assign x_412 = ((((~v_51 | v_34) | v_120) | v_95) | v_128) ;
	assign x_411 = ((((v_28 | ~v_21) | v_137) | ~v_108) | v_151) ;
	assign x_403 = ((((~v_60 | ~v_5) | v_84) | v_106) | ~v_146) ;
	assign x_402 = ((((~v_51 | v_18) | v_121) | v_170) | ~v_101) ;
	assign x_394 = ((((~v_80 | v_34) | v_139) | v_93) | ~v_148) ;
	assign x_393 = ((((~v_11 | v_77) | ~v_158) | v_132) | v_134) ;
	assign x_377 = ((((~v_15 | ~v_39) | v_105) | v_109) | ~v_118) ;
	assign x_376 = ((((v_68 | v_58) | v_175) | ~v_151) | ~v_155) ;
	assign x_360 = ((((v_77 | ~v_51) | v_111) | v_104) | v_178) ;
	assign x_359 = ((((~v_71 | ~v_5) | v_162) | v_85) | ~v_142) ;
	assign x_343 = ((((~v_78 | ~v_24) | v_128) | ~v_132) | v_129) ;
	assign x_342 = ((((~v_63 | v_56) | ~v_165) | v_176) | v_132) ;
	assign x_326 = ((((~v_49 | ~v_72) | v_176) | v_143) | v_125) ;
	assign x_325 = ((((v_19 | ~v_21) | ~v_139) | v_103) | ~v_124) ;
	assign x_309 = ((((v_55 | v_1) | ~v_118) | ~v_116) | ~v_130) ;
	assign x_308 = ((((v_11 | ~v_4) | ~v_131) | ~v_126) | ~v_102) ;
	assign x_292 = ((((~v_40 | v_43) | v_139) | v_88) | v_148) ;
	assign x_291 = ((((v_14 | v_39) | ~v_118) | v_87) | ~v_90) ;
	assign x_275 = ((((~v_38 | ~v_65) | ~v_118) | ~v_104) | v_114) ;
	assign x_274 = ((((~v_74 | v_27) | ~v_155) | v_105) | ~v_96) ;
	assign x_266 = ((((~v_10 | v_63) | v_169) | v_144) | ~v_138) ;
	assign x_265 = ((((~v_21 | v_27) | ~v_101) | ~v_178) | ~v_126) ;
	assign x_257 = ((((v_30 | ~v_79) | v_96) | v_115) | v_173) ;
	assign x_256 = ((((~v_77 | ~v_50) | ~v_81) | ~v_103) | v_151) ;
	assign x_240 = ((((v_14 | v_41) | ~v_99) | ~v_88) | v_83) ;
	assign x_239 = ((((~v_23 | ~v_30) | v_100) | v_105) | ~v_173) ;
	assign x_223 = ((((~v_58 | ~v_10) | ~v_89) | ~v_83) | ~v_81) ;
	assign x_222 = ((((~v_43 | ~v_78) | v_94) | ~v_146) | v_162) ;
	assign x_206 = ((((v_33 | v_25) | ~v_97) | v_104) | ~v_126) ;
	assign x_205 = ((((~v_56 | ~v_59) | ~v_95) | v_94) | v_108) ;
	assign x_197 = ((((~v_51 | ~v_35) | v_139) | v_143) | v_102) ;
	assign x_196 = ((((~v_41 | v_57) | ~v_170) | ~v_166) | v_143) ;
	assign x_188 = ((((v_59 | v_38) | v_162) | ~v_91) | ~v_89) ;
	assign x_187 = ((((~v_59 | v_6) | v_144) | v_173) | ~v_151) ;
	assign x_171 = ((((v_15 | v_4) | ~v_97) | ~v_138) | ~v_176) ;
	assign x_170 = ((((~v_6 | ~v_50) | ~v_176) | v_161) | v_166) ;
	assign x_154 = ((((~v_22 | v_36) | v_122) | ~v_84) | ~v_88) ;
	assign x_153 = ((((~v_45 | v_20) | v_91) | ~v_137) | ~v_157) ;
	assign x_137 = ((((~v_37 | ~v_27) | ~v_105) | ~v_102) | ~v_115) ;
	assign x_136 = ((((v_46 | ~v_65) | v_115) | v_153) | v_158) ;
	assign x_128 = ((((~v_11 | v_52) | v_124) | ~v_156) | v_104) ;
	assign x_127 = ((((v_71 | v_39) | ~v_160) | v_141) | v_151) ;
	assign x_119 = ((((v_2 | ~v_28) | v_83) | ~v_160) | v_153) ;
	assign x_118 = ((((v_53 | ~v_52) | ~v_131) | v_124) | ~v_83) ;
	assign x_102 = ((((v_3 | ~v_34) | ~v_154) | ~v_132) | v_134) ;
	assign x_101 = ((((v_31 | v_64) | v_134) | v_95) | ~v_117) ;
	assign x_85 = ((((~v_66 | ~v_2) | v_148) | ~v_103) | ~v_162) ;
	assign x_84 = ((((v_80 | v_47) | v_146) | ~v_99) | v_135) ;
	assign x_68 = ((((~v_12 | ~v_59) | ~v_143) | ~v_83) | ~v_177) ;
	assign x_67 = ((((~v_28 | v_17) | v_108) | v_90) | ~v_135) ;
	assign x_51 = ((((~v_70 | v_3) | ~v_91) | v_152) | v_148) ;
	assign x_50 = ((((v_75 | v_61) | v_150) | v_144) | v_114) ;
	assign x_34 = ((((v_52 | ~v_39) | ~v_107) | v_89) | v_103) ;
	assign x_33 = ((((~v_34 | v_5) | v_125) | ~v_159) | v_177) ;
	assign x_17 = ((((~v_54 | ~v_43) | ~v_165) | v_121) | v_143) ;
	assign x_16 = ((((v_20 | ~v_5) | v_142) | ~v_171) | v_156) ;
	assign x_2189 = (x_1099 & x_1100) ;
	assign x_1098 = ((((~v_10 | v_69) | v_91) | v_100) | v_101) ;
	assign x_1097 = ((((v_53 | ~v_2) | v_133) | ~v_125) | v_155) ;
	assign x_1096 = ((((~v_32 | v_11) | v_92) | v_109) | v_112) ;
	assign x_1095 = ((((~v_46 | v_37) | ~v_126) | v_135) | ~v_111) ;
	assign x_1094 = ((((~v_35 | ~v_36) | ~v_175) | v_133) | ~v_104) ;
	assign x_1093 = ((((v_19 | ~v_73) | ~v_161) | ~v_104) | v_155) ;
	assign x_1092 = ((((v_13 | v_52) | v_81) | ~v_104) | ~v_147) ;
	assign x_2181 = (x_1090 & x_1091) ;
	assign x_1089 = ((((v_43 | ~v_19) | v_179) | ~v_138) | ~v_160) ;
	assign x_1088 = ((((~v_12 | ~v_62) | v_127) | v_90) | ~v_166) ;
	assign x_1087 = ((((~v_35 | v_65) | ~v_121) | ~v_147) | ~v_150) ;
	assign x_1086 = ((((~v_11 | ~v_46) | ~v_166) | ~v_112) | ~v_160) ;
	assign x_1085 = ((((~v_9 | v_29) | ~v_134) | ~v_126) | v_141) ;
	assign x_1084 = ((((v_12 | v_21) | ~v_131) | v_125) | v_157) ;
	assign x_1083 = ((((~v_29 | ~v_4) | ~v_85) | v_98) | v_136) ;
	assign x_2172 = (x_1081 & x_1082) ;
	assign x_1080 = ((((~v_80 | v_56) | v_112) | v_138) | ~v_144) ;
	assign x_1079 = ((((~v_42 | v_61) | ~v_82) | ~v_94) | v_127) ;
	assign x_1078 = ((((v_75 | v_39) | ~v_89) | v_95) | v_166) ;
	assign x_1077 = ((((~v_29 | ~v_37) | v_137) | ~v_86) | ~v_114) ;
	assign x_1076 = ((((v_24 | v_11) | v_84) | v_146) | ~v_149) ;
	assign x_1075 = ((((v_55 | v_15) | ~v_106) | ~v_125) | ~v_132) ;
	assign x_1074 = ((((v_23 | v_3) | v_109) | v_149) | v_134) ;
	assign x_1073 = ((((v_33 | v_7) | ~v_149) | ~v_91) | v_142) ;
	assign x_1072 = ((((~v_27 | ~v_2) | v_130) | v_165) | ~v_172) ;
	assign x_1071 = ((((~v_41 | v_40) | v_145) | v_180) | ~v_157) ;
	assign x_1070 = ((((~v_39 | ~v_20) | ~v_166) | ~v_118) | ~v_110) ;
	assign x_1069 = ((((v_40 | ~v_43) | v_145) | ~v_97) | v_101) ;
	assign x_1068 = ((((~v_22 | ~v_54) | ~v_170) | ~v_88) | v_177) ;
	assign x_1067 = ((((v_23 | ~v_53) | v_104) | v_177) | ~v_110) ;
	assign x_1066 = ((((v_24 | v_29) | v_152) | ~v_107) | ~v_115) ;
	assign x_2155 = (x_1064 & x_1065) ;
	assign x_1063 = ((((~v_10 | v_60) | ~v_146) | ~v_86) | v_170) ;
	assign x_1062 = ((((~v_40 | ~v_21) | v_156) | v_144) | ~v_136) ;
	assign x_1061 = ((((v_70 | ~v_40) | ~v_154) | v_164) | ~v_146) ;
	assign x_1060 = ((((v_65 | v_50) | v_172) | v_155) | v_163) ;
	assign x_1059 = ((((v_60 | ~v_3) | ~v_132) | v_109) | ~v_148) ;
	assign x_1058 = ((((~v_9 | v_38) | ~v_146) | v_141) | ~v_165) ;
	assign x_1057 = ((((~v_30 | v_37) | v_84) | v_134) | ~v_110) ;
	assign x_1056 = ((((v_44 | v_21) | ~v_138) | v_94) | v_107) ;
	assign x_1055 = ((((v_75 | v_27) | ~v_150) | v_148) | ~v_122) ;
	assign x_1054 = ((((~v_9 | v_50) | ~v_153) | v_141) | ~v_126) ;
	assign x_1053 = ((((v_54 | v_21) | ~v_137) | v_109) | ~v_122) ;
	assign x_1052 = ((((~v_49 | v_43) | v_129) | v_120) | v_104) ;
	assign x_1051 = ((((~v_26 | v_56) | v_156) | ~v_92) | ~v_121) ;
	assign x_1050 = ((((~v_24 | v_23) | ~v_120) | ~v_102) | v_143) ;
	assign x_1049 = ((((v_55 | v_31) | v_110) | v_106) | v_176) ;
	assign x_2139 = (x_1047 & x_1048) ;
	assign x_1046 = ((((~v_52 | v_45) | v_103) | v_81) | v_87) ;
	assign x_1045 = ((((~v_16 | ~v_36) | ~v_83) | ~v_108) | v_128) ;
	assign x_1044 = ((((v_53 | v_26) | ~v_120) | ~v_170) | ~v_179) ;
	assign x_1043 = ((((v_2 | v_17) | ~v_84) | v_92) | v_137) ;
	assign x_1042 = ((((~v_70 | ~v_36) | ~v_120) | v_153) | v_94) ;
	assign x_1041 = ((((v_70 | ~v_40) | ~v_119) | v_108) | v_124) ;
	assign x_1040 = ((((~v_7 | ~v_2) | v_85) | ~v_108) | ~v_84) ;
	assign x_1039 = ((((v_66 | ~v_4) | ~v_90) | ~v_100) | ~v_174) ;
	assign x_1038 = ((((v_44 | v_36) | ~v_134) | v_152) | ~v_108) ;
	assign x_1037 = ((((~v_54 | v_26) | ~v_156) | v_93) | v_90) ;
	assign x_1036 = ((((v_41 | v_5) | v_111) | ~v_175) | ~v_109) ;
	assign x_1035 = ((((~v_58 | v_19) | v_171) | v_152) | ~v_112) ;
	assign x_1034 = ((((~v_29 | ~v_76) | v_167) | ~v_144) | ~v_88) ;
	assign x_1033 = ((((~v_47 | ~v_63) | v_153) | v_154) | v_106) ;
	assign x_1032 = ((((~v_21 | ~v_42) | ~v_154) | ~v_96) | ~v_112) ;
	assign x_2121 = (x_1030 & x_1031) ;
	assign x_1029 = ((((~v_45 | ~v_67) | ~v_84) | v_113) | ~v_178) ;
	assign x_1028 = ((((v_60 | v_67) | v_112) | ~v_137) | v_119) ;
	assign x_1027 = ((((~v_74 | ~v_59) | v_110) | v_143) | v_129) ;
	assign x_1026 = ((((v_75 | v_60) | ~v_84) | ~v_133) | v_115) ;
	assign x_1025 = ((((v_47 | ~v_57) | ~v_119) | v_101) | v_88) ;
	assign x_1024 = ((((v_8 | ~v_70) | v_85) | v_143) | ~v_152) ;
	assign x_1023 = ((((v_48 | v_64) | v_81) | ~v_103) | ~v_110) ;
	assign x_2113 = (x_1021 & x_1022) ;
	assign x_1020 = ((((~v_34 | v_6) | ~v_155) | v_154) | v_129) ;
	assign x_1019 = ((((~v_66 | ~v_14) | v_170) | ~v_168) | ~v_139) ;
	assign x_1018 = ((((v_25 | ~v_76) | ~v_175) | ~v_93) | v_113) ;
	assign x_1017 = ((((~v_18 | ~v_15) | ~v_146) | ~v_141) | ~v_93) ;
	assign x_1016 = ((((v_7 | v_43) | v_93) | v_103) | v_173) ;
	assign x_1015 = ((((~v_65 | ~v_21) | ~v_102) | ~v_88) | v_89) ;
	assign x_1014 = ((((v_5 | v_76) | v_121) | v_114) | ~v_135) ;
	assign x_2104 = (x_1012 & x_1013) ;
	assign x_1011 = ((((~v_25 | v_75) | v_141) | v_107) | ~v_127) ;
	assign x_1010 = ((((~v_13 | ~v_22) | v_169) | v_82) | v_136) ;
	assign x_1009 = ((((~v_27 | ~v_50) | ~v_123) | v_104) | ~v_128) ;
	assign x_1008 = ((((v_63 | v_9) | v_157) | v_103) | v_148) ;
	assign x_1007 = ((((v_35 | v_22) | v_125) | v_129) | ~v_127) ;
	assign x_1006 = ((((v_23 | ~v_10) | ~v_85) | v_158) | ~v_92) ;
	assign x_1005 = ((((~v_7 | v_54) | v_150) | ~v_153) | ~v_140) ;
	assign x_1004 = ((((v_7 | ~v_77) | v_144) | ~v_128) | ~v_115) ;
	assign x_1003 = ((((v_4 | ~v_34) | v_144) | v_129) | ~v_113) ;
	assign x_1002 = ((((~v_40 | v_54) | v_170) | ~v_150) | ~v_163) ;
	assign x_1001 = ((((v_43 | v_40) | v_95) | v_88) | ~v_121) ;
	assign x_1000 = ((((v_53 | v_25) | v_156) | v_132) | v_90) ;
	assign x_999 = ((((v_26 | ~v_25) | v_154) | v_143) | ~v_114) ;
	assign x_998 = ((((~v_50 | v_1) | v_156) | ~v_165) | v_133) ;
	assign x_997 = ((((v_64 | v_34) | v_113) | v_169) | ~v_174) ;
	assign x_2087 = (x_995 & x_996) ;
	assign x_994 = ((((~v_41 | v_22) | v_95) | v_118) | ~v_156) ;
	assign x_993 = ((((~v_8 | v_74) | v_95) | v_90) | v_161) ;
	assign x_992 = ((((v_69 | v_67) | v_128) | ~v_167) | v_82) ;
	assign x_991 = ((((~v_20 | ~v_2) | v_156) | ~v_165) | v_112) ;
	assign x_990 = ((((~v_9 | v_69) | v_88) | v_168) | ~v_96) ;
	assign x_989 = ((((~v_80 | ~v_1) | ~v_162) | v_120) | v_149) ;
	assign x_988 = ((((v_39 | v_35) | v_81) | v_180) | v_153) ;
	assign x_987 = ((((v_8 | v_71) | ~v_111) | ~v_115) | ~v_90) ;
	assign x_986 = ((((v_27 | ~v_53) | ~v_91) | ~v_121) | ~v_81) ;
	assign x_985 = ((((v_55 | v_41) | ~v_135) | v_95) | v_113) ;
	assign x_984 = ((((~v_75 | ~v_8) | ~v_122) | ~v_110) | v_117) ;
	assign x_983 = ((((v_45 | ~v_8) | ~v_107) | ~v_150) | v_141) ;
	assign x_982 = ((((~v_14 | ~v_24) | v_119) | ~v_106) | ~v_134) ;
	assign x_981 = ((((v_23 | ~v_68) | v_100) | v_146) | ~v_103) ;
	assign x_980 = ((((v_36 | ~v_22) | v_152) | v_145) | v_115) ;
	assign x_2071 = (x_978 & x_979) ;
	assign x_977 = ((((v_63 | v_30) | v_154) | v_148) | ~v_143) ;
	assign x_976 = ((((v_9 | ~v_24) | ~v_97) | ~v_139) | v_145) ;
	assign x_975 = ((((~v_70 | v_36) | ~v_106) | ~v_165) | ~v_113) ;
	assign x_974 = ((((v_50 | v_46) | ~v_162) | ~v_160) | v_93) ;
	assign x_973 = ((((~v_17 | ~v_23) | ~v_127) | v_105) | v_175) ;
	assign x_972 = ((((~v_51 | v_38) | v_98) | ~v_122) | v_111) ;
	assign x_971 = ((((v_46 | v_35) | ~v_117) | ~v_123) | ~v_105) ;
	assign x_970 = ((((v_14 | ~v_32) | ~v_87) | v_119) | v_129) ;
	assign x_969 = ((((v_17 | ~v_56) | v_98) | ~v_119) | ~v_151) ;
	assign x_968 = ((((v_16 | ~v_53) | v_175) | ~v_149) | v_90) ;
	assign x_967 = ((((v_37 | v_12) | v_124) | ~v_156) | ~v_155) ;
	assign x_966 = ((((v_52 | ~v_73) | v_128) | v_144) | ~v_87) ;
	assign x_965 = ((((v_58 | v_52) | v_165) | v_179) | v_91) ;
	assign x_964 = ((((v_76 | v_73) | v_157) | ~v_98) | v_120) ;
	assign x_963 = ((((v_58 | v_11) | v_150) | v_136) | ~v_108) ;
	assign x_2052 = (x_961 & x_962) ;
	assign x_960 = ((((v_77 | v_17) | ~v_106) | ~v_152) | v_105) ;
	assign x_959 = ((((v_10 | ~v_35) | ~v_147) | v_114) | ~v_156) ;
	assign x_958 = ((((~v_10 | v_8) | v_129) | ~v_122) | v_153) ;
	assign x_957 = ((((v_44 | v_38) | ~v_170) | v_125) | v_149) ;
	assign x_956 = ((((v_41 | ~v_47) | ~v_168) | v_110) | v_132) ;
	assign x_955 = ((((v_62 | v_12) | v_119) | v_114) | ~v_174) ;
	assign x_954 = ((((~v_38 | ~v_54) | v_152) | ~v_135) | ~v_162) ;
	assign x_2044 = (x_952 & x_953) ;
	assign x_951 = ((((v_15 | ~v_75) | ~v_161) | ~v_82) | ~v_175) ;
	assign x_950 = ((((v_30 | ~v_12) | ~v_96) | v_169) | ~v_174) ;
	assign x_949 = ((((v_15 | v_29) | v_101) | v_107) | ~v_159) ;
	assign x_948 = ((((~v_15 | ~v_32) | v_170) | ~v_173) | v_90) ;
	assign x_947 = ((((~v_17 | ~v_7) | ~v_154) | v_93) | ~v_152) ;
	assign x_946 = ((((v_4 | v_24) | ~v_87) | ~v_148) | ~v_101) ;
	assign x_945 = ((((v_42 | ~v_47) | v_118) | ~v_92) | ~v_141) ;
	assign x_2035 = (x_943 & x_944) ;
	assign x_942 = ((((v_30 | ~v_59) | ~v_142) | ~v_159) | ~v_102) ;
	assign x_941 = ((((v_33 | v_37) | v_163) | v_128) | ~v_141) ;
	assign x_940 = ((((~v_58 | ~v_49) | v_141) | ~v_178) | v_177) ;
	assign x_939 = ((((v_60 | ~v_18) | ~v_139) | ~v_87) | v_91) ;
	assign x_938 = ((((~v_25 | ~v_35) | ~v_110) | v_89) | v_145) ;
	assign x_937 = ((((v_39 | ~v_55) | ~v_109) | ~v_176) | v_115) ;
	assign x_936 = ((((v_54 | v_11) | v_158) | ~v_139) | ~v_130) ;
	assign x_935 = ((((~v_74 | ~v_69) | ~v_85) | ~v_84) | v_119) ;
	assign x_934 = ((((v_76 | v_44) | v_115) | ~v_108) | v_132) ;
	assign x_933 = ((((~v_78 | v_59) | v_148) | ~v_175) | v_150) ;
	assign x_932 = ((((~v_46 | ~v_71) | ~v_155) | ~v_104) | ~v_131) ;
	assign x_931 = ((((~v_39 | v_8) | ~v_116) | v_88) | ~v_133) ;
	assign x_930 = ((((~v_72 | ~v_37) | v_173) | ~v_112) | ~v_122) ;
	assign x_929 = ((((~v_33 | ~v_56) | v_167) | v_164) | v_159) ;
	assign x_928 = ((((v_13 | ~v_22) | ~v_88) | ~v_156) | ~v_102) ;
	assign x_2018 = (x_926 & x_927) ;
	assign x_925 = ((((~v_7 | v_5) | v_96) | v_93) | ~v_157) ;
	assign x_924 = ((((~v_55 | ~v_27) | v_146) | v_95) | v_134) ;
	assign x_923 = ((((v_64 | v_42) | v_110) | v_126) | ~v_139) ;
	assign x_922 = ((((v_64 | ~v_27) | v_137) | ~v_174) | ~v_138) ;
	assign x_921 = ((((v_60 | v_39) | v_160) | v_105) | v_99) ;
	assign x_920 = ((((v_62 | ~v_29) | ~v_90) | v_137) | v_118) ;
	assign x_919 = ((((v_36 | v_41) | v_158) | v_171) | ~v_96) ;
	assign x_918 = ((((v_22 | v_46) | v_168) | v_158) | ~v_144) ;
	assign x_917 = ((((~v_34 | ~v_48) | ~v_110) | ~v_139) | ~v_83) ;
	assign x_916 = ((((v_77 | v_15) | ~v_106) | ~v_177) | ~v_142) ;
	assign x_915 = ((((v_46 | v_5) | v_155) | ~v_169) | ~v_108) ;
	assign x_914 = ((((v_20 | v_40) | ~v_98) | ~v_138) | v_146) ;
	assign x_913 = ((((v_4 | v_58) | v_149) | v_158) | ~v_110) ;
	assign x_912 = ((((~v_39 | v_14) | ~v_169) | v_103) | ~v_115) ;
	assign x_911 = ((((~v_71 | ~v_62) | ~v_166) | ~v_141) | v_132) ;
	assign x_2002 = (x_909 & x_910) ;
	assign x_908 = ((((~v_56 | ~v_27) | ~v_92) | ~v_119) | v_116) ;
	assign x_907 = ((((~v_15 | v_66) | v_114) | ~v_153) | v_142) ;
	assign x_906 = ((((~v_34 | ~v_41) | v_152) | ~v_126) | v_109) ;
	assign x_905 = ((((~v_10 | ~v_18) | ~v_102) | v_170) | v_171) ;
	assign x_904 = ((((v_73 | v_12) | ~v_106) | v_122) | v_172) ;
	assign x_903 = ((((v_75 | v_36) | ~v_116) | ~v_174) | v_92) ;
	assign x_902 = ((((~v_13 | ~v_32) | ~v_114) | v_136) | ~v_84) ;
	assign x_901 = ((((v_77 | ~v_74) | ~v_139) | ~v_127) | v_153) ;
	assign x_900 = ((((~v_42 | v_67) | v_118) | ~v_145) | ~v_173) ;
	assign x_899 = ((((~v_20 | v_60) | v_165) | v_152) | ~v_154) ;
	assign x_898 = ((((v_76 | ~v_21) | ~v_167) | v_162) | ~v_153) ;
	assign x_897 = ((((v_57 | ~v_44) | v_141) | ~v_137) | v_143) ;
	assign x_896 = ((((~v_59 | v_22) | v_157) | v_93) | ~v_89) ;
	assign x_895 = ((((~v_15 | v_27) | ~v_94) | v_147) | ~v_83) ;
	assign x_894 = ((((~v_71 | v_44) | v_158) | ~v_98) | ~v_127) ;
	assign x_1984 = (x_892 & x_893) ;
	assign x_891 = ((((~v_58 | v_28) | v_102) | v_158) | ~v_157) ;
	assign x_890 = ((((~v_22 | v_44) | ~v_141) | v_124) | ~v_172) ;
	assign x_889 = ((((v_39 | ~v_59) | v_109) | ~v_179) | v_166) ;
	assign x_888 = ((((~v_79 | v_42) | ~v_116) | v_146) | ~v_180) ;
	assign x_887 = ((((v_56 | v_22) | v_127) | ~v_107) | ~v_171) ;
	assign x_886 = ((((~v_29 | ~v_40) | ~v_81) | v_92) | ~v_115) ;
	assign x_885 = ((((v_73 | ~v_8) | ~v_133) | v_103) | v_173) ;
	assign x_884 = ((((v_57 | v_19) | v_165) | v_160) | ~v_180) ;
	assign x_883 = ((((~v_37 | v_20) | v_178) | ~v_114) | ~v_162) ;
	assign x_882 = ((((v_59 | ~v_39) | v_135) | v_137) | ~v_86) ;
	assign x_881 = ((((v_24 | v_50) | ~v_145) | v_105) | ~v_106) ;
	assign x_880 = ((((v_71 | ~v_23) | ~v_152) | v_115) | v_87) ;
	assign x_879 = ((((v_21 | v_18) | ~v_161) | v_155) | ~v_101) ;
	assign x_878 = ((((v_43 | v_56) | v_139) | ~v_122) | v_116) ;
	assign x_877 = ((((v_57 | v_62) | ~v_104) | v_177) | ~v_94) ;
	assign x_1968 = (x_875 & x_876) ;
	assign x_874 = ((((v_53 | ~v_12) | v_154) | v_90) | ~v_178) ;
	assign x_873 = ((((v_8 | v_51) | v_99) | ~v_148) | ~v_161) ;
	assign x_872 = ((((~v_75 | v_14) | ~v_134) | ~v_96) | v_141) ;
	assign x_871 = ((((v_3 | ~v_67) | ~v_120) | ~v_87) | v_90) ;
	assign x_870 = ((((~v_80 | v_38) | ~v_111) | ~v_98) | ~v_151) ;
	assign x_869 = ((((~v_47 | ~v_76) | ~v_135) | v_86) | ~v_118) ;
	assign x_868 = ((((v_35 | v_71) | ~v_179) | v_176) | v_97) ;
	assign x_867 = ((((v_46 | ~v_72) | ~v_163) | ~v_157) | ~v_118) ;
	assign x_866 = ((((v_55 | ~v_74) | v_102) | v_117) | ~v_115) ;
	assign x_865 = ((((v_51 | v_74) | ~v_107) | ~v_88) | v_161) ;
	assign x_864 = ((((v_23 | ~v_71) | v_179) | ~v_149) | v_126) ;
	assign x_863 = ((((~v_67 | v_29) | ~v_173) | v_116) | ~v_172) ;
	assign x_862 = ((((v_36 | ~v_62) | ~v_136) | ~v_116) | ~v_123) ;
	assign x_861 = ((((v_50 | v_33) | ~v_143) | ~v_121) | v_173) ;
	assign x_860 = ((((~v_63 | v_23) | ~v_135) | ~v_81) | ~v_175) ;
	assign x_1951 = (x_858 & x_859) ;
	assign x_857 = ((((~v_12 | v_29) | v_100) | ~v_95) | ~v_175) ;
	assign x_856 = ((((v_66 | ~v_75) | v_81) | ~v_111) | ~v_171) ;
	assign x_855 = ((((v_23 | ~v_49) | ~v_116) | ~v_110) | ~v_151) ;
	assign x_854 = ((((~v_16 | ~v_55) | v_88) | v_177) | v_119) ;
	assign x_853 = ((((~v_52 | v_13) | v_105) | v_166) | ~v_158) ;
	assign x_852 = ((((v_46 | ~v_39) | v_146) | ~v_135) | ~v_150) ;
	assign x_851 = ((((~v_33 | v_80) | v_102) | v_104) | v_81) ;
	assign x_850 = ((((~v_10 | ~v_29) | ~v_161) | v_90) | ~v_151) ;
	assign x_849 = ((((~v_41 | v_54) | v_166) | ~v_93) | ~v_119) ;
	assign x_848 = ((((~v_80 | ~v_21) | ~v_109) | ~v_143) | v_138) ;
	assign x_847 = ((((v_27 | v_45) | v_101) | v_109) | ~v_125) ;
	assign x_846 = ((((v_74 | v_76) | ~v_169) | ~v_98) | ~v_162) ;
	assign x_845 = ((((~v_46 | v_26) | v_177) | ~v_90) | ~v_167) ;
	assign x_844 = ((((v_69 | v_47) | ~v_149) | ~v_120) | v_107) ;
	assign x_843 = ((((v_27 | ~v_51) | v_141) | v_82) | v_173) ;
	assign x_1935 = (x_841 & x_842) ;
	assign x_840 = ((((~v_46 | v_75) | v_136) | v_88) | ~v_122) ;
	assign x_839 = ((((v_63 | ~v_76) | v_131) | ~v_148) | ~v_93) ;
	assign x_838 = ((((v_7 | v_5) | v_133) | v_153) | ~v_118) ;
	assign x_837 = ((((~v_60 | v_12) | ~v_130) | v_149) | ~v_179) ;
	assign x_836 = ((((v_33 | v_47) | ~v_153) | v_126) | v_110) ;
	assign x_835 = ((((v_24 | v_20) | ~v_82) | v_131) | v_126) ;
	assign x_834 = ((((~v_21 | ~v_64) | v_172) | v_82) | v_162) ;
	assign x_833 = ((((v_42 | v_32) | v_111) | ~v_136) | ~v_112) ;
	assign x_832 = ((((~v_7 | v_47) | v_175) | v_163) | v_87) ;
	assign x_831 = ((((v_26 | ~v_68) | ~v_136) | v_91) | v_176) ;
	assign x_830 = ((((v_66 | v_61) | ~v_161) | v_135) | ~v_131) ;
	assign x_829 = ((((v_2 | v_17) | ~v_163) | v_94) | v_121) ;
	assign x_828 = ((((~v_32 | ~v_4) | ~v_144) | v_91) | v_89) ;
	assign x_827 = ((((v_34 | ~v_45) | v_175) | v_174) | ~v_96) ;
	assign x_826 = ((((v_57 | ~v_26) | ~v_106) | v_121) | ~v_105) ;
	assign x_1915 = (x_824 & x_825) ;
	assign x_823 = ((((v_51 | v_43) | ~v_169) | ~v_123) | v_101) ;
	assign x_822 = ((((v_43 | v_11) | ~v_154) | ~v_136) | v_152) ;
	assign x_821 = ((((~v_40 | v_73) | v_180) | v_133) | ~v_119) ;
	assign x_820 = ((((v_28 | ~v_44) | v_149) | ~v_85) | v_107) ;
	assign x_819 = ((((v_55 | v_67) | v_169) | v_135) | v_142) ;
	assign x_818 = ((((~v_44 | v_23) | v_133) | ~v_175) | ~v_104) ;
	assign x_817 = ((((~v_21 | v_17) | ~v_86) | v_152) | v_171) ;
	assign x_1907 = (x_815 & x_816) ;
	assign x_814 = ((((~v_6 | v_70) | ~v_179) | ~v_107) | v_121) ;
	assign x_813 = ((((v_56 | ~v_40) | v_165) | ~v_82) | v_98) ;
	assign x_812 = ((((~v_45 | v_27) | ~v_84) | v_118) | ~v_155) ;
	assign x_811 = ((((~v_58 | ~v_7) | ~v_166) | ~v_171) | v_131) ;
	assign x_810 = ((((~v_4 | v_31) | ~v_136) | v_107) | ~v_97) ;
	assign x_809 = ((((v_37 | v_68) | ~v_126) | ~v_175) | ~v_133) ;
	assign x_808 = ((((v_79 | ~v_76) | ~v_169) | v_163) | v_176) ;
	assign x_1898 = (x_806 & x_807) ;
	assign x_805 = ((((~v_67 | ~v_54) | ~v_108) | ~v_139) | v_90) ;
	assign x_804 = ((((~v_36 | ~v_68) | v_134) | v_124) | v_103) ;
	assign x_803 = ((((~v_80 | ~v_58) | ~v_162) | ~v_172) | v_124) ;
	assign x_802 = ((((~v_53 | ~v_22) | ~v_154) | ~v_82) | ~v_151) ;
	assign x_801 = ((((v_3 | ~v_68) | ~v_145) | ~v_165) | ~v_159) ;
	assign x_800 = ((((~v_35 | v_74) | v_176) | ~v_151) | v_141) ;
	assign x_799 = ((((v_35 | v_43) | ~v_121) | ~v_164) | v_93) ;
	assign x_798 = ((((~v_6 | ~v_11) | v_118) | ~v_91) | v_124) ;
	assign x_797 = ((((v_8 | ~v_21) | ~v_151) | ~v_101) | ~v_83) ;
	assign x_796 = ((((~v_37 | v_77) | v_108) | v_86) | v_137) ;
	assign x_795 = ((((v_53 | v_23) | ~v_122) | v_111) | ~v_113) ;
	assign x_794 = ((((~v_67 | v_60) | ~v_153) | ~v_89) | v_172) ;
	assign x_793 = ((((v_1 | ~v_63) | v_122) | v_140) | ~v_83) ;
	assign x_792 = ((((~v_9 | v_44) | v_150) | ~v_121) | v_157) ;
	assign x_791 = ((((v_68 | ~v_7) | ~v_90) | ~v_100) | v_93) ;
	assign x_1881 = (x_789 & x_790) ;
	assign x_788 = ((((~v_5 | v_62) | v_141) | ~v_161) | v_179) ;
	assign x_787 = ((((~v_61 | v_36) | v_147) | v_169) | ~v_107) ;
	assign x_786 = ((((v_11 | ~v_14) | ~v_85) | v_86) | ~v_89) ;
	assign x_785 = ((((~v_79 | v_66) | ~v_112) | ~v_158) | ~v_144) ;
	assign x_784 = ((((v_30 | ~v_76) | v_121) | ~v_125) | ~v_115) ;
	assign x_783 = ((((~v_40 | ~v_23) | v_122) | ~v_120) | v_147) ;
	assign x_782 = ((((~v_39 | v_15) | v_90) | v_147) | v_120) ;
	assign x_781 = ((((v_39 | ~v_38) | v_117) | ~v_178) | v_131) ;
	assign x_780 = ((((~v_65 | ~v_68) | ~v_167) | v_116) | v_118) ;
	assign x_779 = ((((v_65 | ~v_62) | v_160) | v_87) | ~v_84) ;
	assign x_778 = ((((~v_51 | v_22) | v_126) | ~v_165) | v_97) ;
	assign x_777 = ((((v_47 | v_48) | ~v_102) | v_154) | ~v_158) ;
	assign x_776 = ((((~v_14 | ~v_46) | ~v_153) | v_107) | ~v_174) ;
	assign x_775 = ((((v_16 | ~v_26) | v_132) | v_166) | ~v_116) ;
	assign x_774 = ((((~v_7 | ~v_21) | v_138) | ~v_153) | v_146) ;
	assign x_1865 = (x_772 & x_773) ;
	assign x_771 = ((((v_7 | ~v_9) | ~v_124) | ~v_99) | ~v_83) ;
	assign x_770 = ((((v_14 | ~v_13) | v_130) | v_97) | v_161) ;
	assign x_769 = ((((v_56 | ~v_27) | ~v_103) | ~v_156) | v_149) ;
	assign x_768 = ((((~v_43 | ~v_77) | v_163) | ~v_178) | ~v_149) ;
	assign x_767 = ((((~v_39 | v_49) | v_94) | v_116) | ~v_97) ;
	assign x_766 = ((((~v_33 | v_47) | v_147) | v_161) | ~v_125) ;
	assign x_765 = ((((~v_24 | ~v_63) | v_175) | v_130) | ~v_150) ;
	assign x_764 = ((((~v_5 | v_4) | v_122) | ~v_90) | ~v_133) ;
	assign x_763 = ((((~v_62 | v_5) | ~v_174) | v_151) | v_173) ;
	assign x_762 = ((((v_74 | ~v_69) | v_156) | ~v_127) | v_138) ;
	assign x_761 = ((((v_16 | ~v_11) | v_111) | ~v_171) | v_178) ;
	assign x_760 = ((((v_43 | ~v_60) | v_163) | v_152) | ~v_107) ;
	assign x_759 = ((((v_47 | ~v_69) | ~v_106) | ~v_126) | ~v_164) ;
	assign x_758 = ((((~v_71 | ~v_5) | v_124) | ~v_125) | v_105) ;
	assign x_757 = ((((v_67 | v_65) | ~v_143) | ~v_82) | v_85) ;
	assign x_1847 = (x_755 & x_756) ;
	assign x_754 = ((((v_28 | ~v_15) | v_153) | v_88) | ~v_87) ;
	assign x_753 = ((((~v_53 | ~v_46) | ~v_158) | v_85) | ~v_113) ;
	assign x_752 = ((((v_3 | v_14) | ~v_140) | ~v_171) | ~v_164) ;
	assign x_751 = ((((v_31 | v_2) | v_137) | ~v_83) | v_103) ;
	assign x_750 = ((((v_56 | ~v_7) | v_104) | v_107) | v_175) ;
	assign x_749 = ((((v_17 | ~v_74) | ~v_110) | ~v_114) | v_124) ;
	assign x_748 = ((((~v_69 | v_8) | v_147) | ~v_125) | v_89) ;
	assign x_1839 = (x_746 & x_747) ;
	assign x_745 = ((((v_29 | v_35) | v_133) | ~v_163) | v_120) ;
	assign x_744 = ((((v_26 | v_27) | ~v_152) | v_142) | v_103) ;
	assign x_743 = ((((v_70 | v_57) | v_132) | ~v_162) | ~v_167) ;
	assign x_742 = ((((~v_22 | v_67) | v_101) | ~v_159) | ~v_113) ;
	assign x_741 = ((((v_59 | ~v_65) | ~v_121) | ~v_155) | v_115) ;
	assign x_740 = ((((v_22 | ~v_2) | v_155) | v_161) | v_147) ;
	assign x_739 = ((((~v_10 | ~v_61) | v_165) | ~v_114) | v_163) ;
	assign x_1830 = (x_737 & x_738) ;
	assign x_736 = ((((~v_69 | ~v_4) | ~v_118) | ~v_171) | v_153) ;
	assign x_735 = ((((v_18 | v_39) | v_135) | ~v_147) | v_152) ;
	assign x_734 = ((((~v_21 | v_24) | ~v_162) | v_178) | ~v_160) ;
	assign x_733 = ((((v_34 | ~v_57) | ~v_146) | v_101) | ~v_103) ;
	assign x_732 = ((((~v_45 | ~v_43) | v_127) | v_173) | ~v_101) ;
	assign x_731 = ((((~v_40 | ~v_71) | v_117) | v_132) | ~v_105) ;
	assign x_730 = ((((~v_18 | ~v_32) | ~v_116) | ~v_156) | ~v_142) ;
	assign x_729 = ((((~v_17 | ~v_64) | ~v_175) | v_95) | ~v_97) ;
	assign x_728 = ((((v_19 | v_16) | v_122) | ~v_175) | v_151) ;
	assign x_727 = ((((~v_75 | ~v_59) | ~v_177) | v_150) | v_159) ;
	assign x_726 = ((((v_32 | v_27) | ~v_180) | ~v_150) | ~v_170) ;
	assign x_725 = ((((~v_65 | ~v_50) | ~v_130) | v_144) | ~v_97) ;
	assign x_724 = ((((v_74 | v_59) | ~v_160) | ~v_131) | ~v_156) ;
	assign x_723 = ((((v_12 | v_61) | ~v_110) | ~v_104) | ~v_120) ;
	assign x_722 = ((((v_52 | v_49) | ~v_133) | ~v_159) | ~v_129) ;
	assign x_1813 = (x_720 & x_721) ;
	assign x_719 = ((((~v_51 | ~v_27) | v_137) | v_150) | v_83) ;
	assign x_718 = ((((~v_41 | v_39) | ~v_150) | ~v_155) | v_93) ;
	assign x_717 = ((((v_67 | v_47) | v_96) | v_111) | v_144) ;
	assign x_716 = ((((~v_19 | v_73) | ~v_91) | v_156) | ~v_149) ;
	assign x_715 = ((((~v_38 | v_75) | ~v_134) | ~v_176) | v_81) ;
	assign x_714 = ((((v_50 | v_17) | v_126) | ~v_116) | v_145) ;
	assign x_713 = ((((~v_12 | ~v_72) | ~v_178) | v_138) | v_147) ;
	assign x_712 = ((((v_21 | ~v_73) | v_164) | ~v_169) | v_118) ;
	assign x_711 = ((((~v_57 | v_39) | v_145) | v_176) | v_103) ;
	assign x_710 = ((((v_32 | ~v_9) | ~v_154) | v_144) | ~v_146) ;
	assign x_709 = ((((~v_40 | ~v_56) | ~v_84) | ~v_81) | v_104) ;
	assign x_708 = ((((v_43 | v_60) | v_134) | ~v_132) | ~v_130) ;
	assign x_707 = ((((~v_11 | ~v_41) | ~v_173) | v_174) | ~v_131) ;
	assign x_706 = ((((~v_42 | v_51) | v_139) | v_131) | ~v_88) ;
	assign x_705 = ((((v_58 | ~v_31) | ~v_93) | ~v_108) | v_106) ;
	assign x_1797 = (x_703 & x_704) ;
	assign x_702 = ((((~v_79 | ~v_1) | ~v_180) | ~v_87) | v_163) ;
	assign x_701 = ((((v_33 | v_50) | ~v_105) | v_111) | v_143) ;
	assign x_700 = ((((v_44 | v_21) | v_169) | v_145) | ~v_118) ;
	assign x_699 = ((((~v_6 | ~v_50) | v_171) | ~v_157) | ~v_97) ;
	assign x_698 = ((((v_23 | ~v_45) | ~v_99) | ~v_112) | ~v_154) ;
	assign x_697 = ((((~v_2 | ~v_42) | v_171) | ~v_176) | v_84) ;
	assign x_696 = ((((~v_28 | v_26) | v_177) | ~v_129) | ~v_136) ;
	assign x_695 = ((((~v_66 | ~v_65) | v_160) | ~v_104) | ~v_145) ;
	assign x_694 = ((((~v_44 | ~v_51) | ~v_145) | v_111) | ~v_96) ;
	assign x_693 = ((((v_1 | v_46) | ~v_84) | v_95) | ~v_87) ;
	assign x_692 = ((((v_14 | v_23) | v_179) | ~v_85) | v_97) ;
	assign x_691 = ((((~v_50 | ~v_58) | ~v_131) | v_101) | ~v_139) ;
	assign x_690 = ((((v_41 | ~v_60) | ~v_121) | ~v_117) | v_165) ;
	assign x_689 = ((((v_42 | ~v_71) | v_152) | ~v_137) | ~v_116) ;
	assign x_688 = ((((~v_69 | ~v_13) | v_108) | ~v_133) | ~v_126) ;
	assign x_1778 = (x_686 & x_687) ;
	assign x_685 = ((((v_76 | ~v_80) | ~v_164) | ~v_178) | v_148) ;
	assign x_684 = ((((v_71 | ~v_47) | v_114) | v_160) | v_135) ;
	assign x_683 = ((((~v_5 | v_74) | ~v_138) | ~v_92) | ~v_96) ;
	assign x_682 = ((((v_36 | ~v_14) | ~v_126) | v_128) | ~v_99) ;
	assign x_681 = ((((v_41 | v_27) | v_134) | v_109) | ~v_91) ;
	assign x_680 = ((((~v_1 | v_9) | v_92) | v_105) | v_139) ;
	assign x_679 = ((((v_71 | ~v_69) | v_115) | ~v_167) | ~v_83) ;
	assign x_1770 = (x_677 & x_678) ;
	assign x_676 = ((((~v_54 | ~v_27) | ~v_104) | v_128) | ~v_140) ;
	assign x_675 = ((((~v_48 | v_41) | v_137) | v_171) | v_100) ;
	assign x_674 = ((((v_68 | v_11) | v_155) | ~v_174) | ~v_165) ;
	assign x_673 = ((((v_73 | ~v_57) | v_120) | v_94) | v_163) ;
	assign x_672 = ((((~v_69 | ~v_63) | v_179) | ~v_144) | v_125) ;
	assign x_671 = ((((v_10 | ~v_48) | v_82) | ~v_105) | ~v_135) ;
	assign x_670 = ((((v_51 | ~v_16) | v_133) | ~v_142) | v_177) ;
	assign x_1761 = (x_668 & x_669) ;
	assign x_667 = ((((v_7 | v_16) | ~v_107) | v_155) | v_126) ;
	assign x_666 = ((((v_28 | ~v_11) | v_112) | ~v_176) | v_119) ;
	assign x_665 = ((((v_41 | ~v_74) | v_165) | v_119) | ~v_127) ;
	assign x_664 = ((((~v_10 | v_29) | v_131) | ~v_155) | ~v_106) ;
	assign x_663 = ((((~v_46 | ~v_52) | ~v_124) | v_126) | v_91) ;
	assign x_662 = ((((v_50 | v_10) | v_169) | ~v_136) | ~v_127) ;
	assign x_661 = ((((v_35 | v_24) | v_153) | ~v_82) | v_138) ;
	assign x_660 = ((((~v_11 | v_17) | v_85) | ~v_136) | v_86) ;
	assign x_659 = ((((~v_20 | v_7) | v_178) | ~v_112) | ~v_171) ;
	assign x_658 = ((((v_19 | v_3) | ~v_136) | v_162) | ~v_84) ;
	assign x_657 = ((((v_50 | v_5) | ~v_158) | ~v_128) | ~v_119) ;
	assign x_656 = ((((~v_14 | ~v_30) | ~v_169) | v_143) | v_161) ;
	assign x_655 = ((((~v_52 | ~v_2) | v_139) | ~v_148) | v_122) ;
	assign x_654 = ((((~v_62 | v_38) | v_93) | ~v_116) | v_145) ;
	assign x_653 = ((((~v_38 | v_48) | v_150) | v_116) | v_164) ;
	assign x_1744 = (x_651 & x_652) ;
	assign x_650 = ((((v_15 | ~v_58) | v_106) | v_180) | ~v_108) ;
	assign x_649 = ((((~v_20 | ~v_80) | ~v_143) | v_83) | ~v_178) ;
	assign x_648 = ((((v_65 | ~v_31) | ~v_97) | v_154) | ~v_86) ;
	assign x_647 = ((((~v_11 | ~v_52) | ~v_96) | v_176) | ~v_177) ;
	assign x_646 = ((((~v_23 | v_64) | ~v_164) | ~v_178) | v_153) ;
	assign x_645 = ((((~v_58 | ~v_49) | v_164) | v_119) | ~v_137) ;
	assign x_644 = ((((~v_20 | ~v_55) | ~v_141) | v_155) | v_128) ;
	assign x_643 = ((((~v_34 | ~v_5) | ~v_92) | v_112) | v_83) ;
	assign x_642 = ((((~v_53 | v_33) | v_147) | ~v_149) | ~v_156) ;
	assign x_641 = ((((~v_71 | v_13) | ~v_156) | ~v_177) | ~v_99) ;
	assign x_640 = ((((~v_9 | v_62) | v_180) | v_128) | v_166) ;
	assign x_639 = ((((~v_29 | v_6) | ~v_156) | v_112) | ~v_127) ;
	assign x_638 = ((((~v_28 | ~v_45) | ~v_95) | v_140) | ~v_97) ;
	assign x_637 = ((((v_42 | v_9) | ~v_162) | ~v_137) | v_172) ;
	assign x_636 = ((((v_66 | v_68) | v_98) | v_167) | v_151) ;
	assign x_1728 = (x_634 & x_635) ;
	assign x_633 = ((((~v_17 | ~v_61) | v_148) | ~v_141) | ~v_84) ;
	assign x_632 = ((((v_8 | ~v_44) | ~v_90) | ~v_158) | ~v_112) ;
	assign x_631 = ((((v_64 | ~v_4) | ~v_113) | v_134) | ~v_137) ;
	assign x_630 = ((((v_44 | v_33) | v_168) | v_145) | ~v_90) ;
	assign x_629 = ((((~v_24 | ~v_72) | v_168) | v_93) | v_84) ;
	assign x_628 = ((((~v_31 | ~v_39) | v_84) | ~v_133) | v_155) ;
	assign x_627 = ((((~v_78 | v_11) | ~v_144) | v_108) | ~v_115) ;
	assign x_626 = ((((v_18 | v_7) | ~v_140) | v_105) | v_153) ;
	assign x_625 = ((((~v_50 | v_45) | ~v_179) | ~v_103) | v_142) ;
	assign x_624 = ((((~v_21 | ~v_58) | ~v_97) | v_177) | ~v_161) ;
	assign x_623 = ((((v_29 | v_73) | ~v_161) | ~v_130) | ~v_117) ;
	assign x_622 = ((((v_62 | v_16) | v_162) | v_138) | ~v_163) ;
	assign x_621 = ((((v_76 | ~v_8) | ~v_180) | ~v_179) | ~v_172) ;
	assign x_620 = ((((v_22 | v_54) | ~v_153) | ~v_165) | v_98) ;
	assign x_619 = ((((v_16 | ~v_74) | v_122) | v_96) | v_162) ;
	assign x_1710 = (x_617 & x_618) ;
	assign x_616 = ((((~v_70 | ~v_25) | ~v_146) | ~v_144) | ~v_123) ;
	assign x_615 = ((((v_46 | ~v_28) | ~v_123) | v_128) | ~v_91) ;
	assign x_614 = ((((v_27 | ~v_79) | ~v_127) | ~v_171) | v_117) ;
	assign x_613 = ((((v_44 | v_9) | ~v_111) | ~v_165) | ~v_126) ;
	assign x_612 = ((((~v_36 | v_14) | v_100) | v_163) | v_86) ;
	assign x_611 = ((((~v_72 | ~v_6) | v_114) | v_130) | v_142) ;
	assign x_610 = ((((v_5 | ~v_48) | ~v_135) | v_126) | ~v_170) ;
	assign x_609 = ((((~v_28 | v_8) | v_117) | v_133) | ~v_141) ;
	assign x_608 = ((((v_51 | v_49) | ~v_131) | v_137) | ~v_127) ;
	assign x_607 = ((((v_38 | v_21) | v_123) | ~v_112) | ~v_173) ;
	assign x_606 = ((((v_58 | v_16) | ~v_115) | v_126) | v_131) ;
	assign x_605 = ((((v_52 | ~v_27) | ~v_99) | v_173) | ~v_154) ;
	assign x_604 = ((((v_54 | ~v_39) | v_155) | v_122) | ~v_137) ;
	assign x_603 = ((((~v_30 | ~v_6) | ~v_101) | ~v_111) | v_109) ;
	assign x_602 = ((((~v_59 | ~v_63) | ~v_116) | ~v_140) | v_122) ;
	assign x_1694 = (x_600 & x_601) ;
	assign x_599 = ((((v_15 | v_76) | v_119) | v_115) | ~v_112) ;
	assign x_598 = ((((~v_23 | v_35) | v_111) | v_84) | v_158) ;
	assign x_597 = ((((v_57 | v_29) | v_127) | v_139) | v_99) ;
	assign x_596 = ((((~v_13 | ~v_6) | ~v_82) | ~v_92) | ~v_112) ;
	assign x_595 = ((((v_77 | v_60) | ~v_150) | ~v_90) | v_110) ;
	assign x_594 = ((((~v_34 | ~v_22) | ~v_178) | v_95) | v_149) ;
	assign x_593 = ((((~v_40 | ~v_11) | v_151) | ~v_91) | v_105) ;
	assign x_592 = ((((~v_45 | ~v_9) | ~v_152) | ~v_124) | ~v_87) ;
	assign x_591 = ((((~v_46 | v_75) | ~v_144) | ~v_95) | v_97) ;
	assign x_590 = ((((~v_77 | v_63) | v_88) | ~v_96) | ~v_179) ;
	assign x_589 = ((((~v_79 | ~v_9) | ~v_153) | ~v_137) | ~v_142) ;
	assign x_588 = ((((~v_13 | ~v_80) | ~v_97) | ~v_93) | v_155) ;
	assign x_587 = ((((v_66 | ~v_9) | ~v_151) | v_149) | v_130) ;
	assign x_586 = ((((~v_3 | v_32) | ~v_162) | ~v_171) | v_91) ;
	assign x_585 = ((((~v_63 | v_17) | ~v_83) | v_84) | ~v_162) ;
	assign x_1677 = (x_583 & x_584) ;
	assign x_582 = ((((v_63 | v_55) | ~v_93) | v_170) | ~v_103) ;
	assign x_581 = ((((v_56 | v_4) | ~v_123) | v_92) | v_173) ;
	assign x_580 = ((((~v_11 | ~v_50) | ~v_159) | v_143) | ~v_118) ;
	assign x_579 = ((((v_62 | v_65) | v_173) | v_132) | v_107) ;
	assign x_578 = ((((~v_39 | ~v_35) | ~v_141) | v_96) | v_116) ;
	assign x_577 = ((((~v_7 | v_63) | v_130) | ~v_164) | ~v_162) ;
	assign x_576 = ((((v_32 | v_42) | ~v_150) | ~v_122) | v_96) ;
	assign x_575 = ((((~v_29 | v_47) | v_174) | ~v_139) | ~v_172) ;
	assign x_574 = ((((~v_58 | v_40) | ~v_152) | v_154) | ~v_159) ;
	assign x_573 = ((((v_75 | v_54) | ~v_174) | v_151) | ~v_94) ;
	assign x_572 = ((((v_38 | ~v_21) | v_113) | ~v_139) | ~v_114) ;
	assign x_571 = ((((v_63 | ~v_52) | ~v_142) | v_125) | v_108) ;
	assign x_570 = ((((~v_27 | ~v_9) | ~v_131) | ~v_143) | v_108) ;
	assign x_569 = ((((~v_40 | v_38) | v_150) | ~v_124) | v_174) ;
	assign x_568 = ((((v_67 | ~v_49) | v_157) | ~v_125) | ~v_154) ;
	assign x_1661 = (x_566 & x_567) ;
	assign x_565 = ((((~v_70 | v_3) | ~v_118) | ~v_146) | ~v_127) ;
	assign x_564 = ((((v_31 | ~v_68) | v_134) | v_89) | v_139) ;
	assign x_563 = ((((v_35 | v_66) | ~v_92) | ~v_88) | v_169) ;
	assign x_562 = ((((~v_48 | ~v_54) | v_130) | v_167) | ~v_102) ;
	assign x_561 = ((((~v_5 | ~v_36) | ~v_116) | ~v_150) | v_164) ;
	assign x_560 = ((((v_16 | v_37) | v_140) | ~v_161) | ~v_172) ;
	assign x_559 = ((((v_54 | ~v_79) | v_94) | v_133) | v_173) ;
	assign x_558 = ((((v_75 | ~v_53) | ~v_157) | v_117) | ~v_116) ;
	assign x_557 = ((((v_59 | ~v_25) | ~v_138) | v_156) | v_179) ;
	assign x_556 = ((((~v_47 | v_41) | v_155) | ~v_157) | ~v_111) ;
	assign x_555 = ((((~v_51 | v_79) | v_120) | v_117) | v_170) ;
	assign x_554 = ((((~v_73 | ~v_34) | v_172) | ~v_129) | v_93) ;
	assign x_553 = ((((~v_33 | v_50) | ~v_137) | ~v_162) | ~v_156) ;
	assign x_552 = ((((~v_36 | ~v_19) | ~v_168) | v_148) | v_142) ;
	assign x_551 = ((((v_49 | ~v_73) | v_142) | v_103) | v_152) ;
	assign x_1640 = (x_549 & x_550) ;
	assign x_548 = ((((v_58 | ~v_67) | ~v_114) | ~v_107) | v_171) ;
	assign x_547 = ((((v_59 | v_9) | ~v_164) | v_141) | v_173) ;
	assign x_546 = ((((~v_31 | v_17) | v_92) | ~v_97) | ~v_107) ;
	assign x_545 = ((((~v_3 | ~v_13) | ~v_100) | v_141) | v_176) ;
	assign x_544 = ((((v_29 | ~v_39) | ~v_102) | ~v_148) | v_86) ;
	assign x_543 = ((((v_37 | v_48) | v_179) | ~v_136) | ~v_174) ;
	assign x_542 = ((((~v_8 | v_58) | ~v_143) | ~v_128) | v_173) ;
	assign x_1632 = (x_540 & x_541) ;
	assign x_539 = ((((v_66 | ~v_73) | v_175) | ~v_180) | v_128) ;
	assign x_538 = ((((~v_41 | v_75) | ~v_142) | ~v_101) | v_176) ;
	assign x_537 = ((((~v_34 | v_29) | ~v_167) | ~v_173) | ~v_115) ;
	assign x_536 = ((((~v_48 | v_43) | ~v_176) | ~v_87) | v_103) ;
	assign x_535 = ((((v_74 | v_28) | ~v_162) | v_93) | ~v_86) ;
	assign x_534 = ((((v_58 | ~v_2) | v_114) | ~v_122) | v_161) ;
	assign x_533 = ((((v_30 | ~v_11) | ~v_151) | v_147) | v_135) ;
	assign x_1623 = (x_531 & x_532) ;
	assign x_530 = ((((~v_3 | ~v_23) | ~v_128) | ~v_133) | v_137) ;
	assign x_529 = ((((v_16 | v_32) | v_95) | v_89) | v_152) ;
	assign x_528 = ((((~v_66 | v_37) | v_126) | v_101) | v_138) ;
	assign x_527 = ((((~v_39 | ~v_70) | v_96) | ~v_134) | ~v_153) ;
	assign x_526 = ((((v_45 | ~v_30) | ~v_135) | v_164) | v_176) ;
	assign x_525 = ((((~v_64 | ~v_33) | v_163) | v_120) | v_91) ;
	assign x_524 = ((((~v_60 | v_52) | v_162) | v_173) | ~v_117) ;
	assign x_523 = ((((v_79 | ~v_46) | v_128) | ~v_88) | v_175) ;
	assign x_522 = ((((~v_53 | v_50) | ~v_156) | ~v_104) | ~v_102) ;
	assign x_521 = ((((~v_27 | ~v_59) | v_147) | v_144) | ~v_130) ;
	assign x_520 = ((((v_7 | ~v_74) | v_112) | v_125) | v_158) ;
	assign x_519 = ((((~v_77 | ~v_1) | ~v_160) | v_169) | v_148) ;
	assign x_518 = ((((v_42 | ~v_8) | ~v_110) | v_97) | ~v_96) ;
	assign x_517 = ((((~v_56 | ~v_12) | ~v_114) | ~v_111) | v_89) ;
	assign x_516 = ((((v_59 | v_5) | ~v_146) | ~v_152) | v_164) ;
	assign x_1606 = (x_514 & x_515) ;
	assign x_513 = ((((v_47 | ~v_61) | ~v_169) | ~v_105) | v_152) ;
	assign x_512 = ((((~v_71 | ~v_6) | v_119) | ~v_136) | ~v_137) ;
	assign x_511 = ((((v_51 | ~v_7) | ~v_180) | v_142) | v_85) ;
	assign x_510 = ((((~v_44 | v_20) | v_96) | v_84) | ~v_112) ;
	assign x_509 = ((((~v_3 | ~v_9) | v_97) | v_138) | v_99) ;
	assign x_508 = ((((v_45 | v_63) | ~v_155) | v_124) | ~v_88) ;
	assign x_507 = ((((v_73 | v_3) | ~v_175) | ~v_86) | ~v_163) ;
	assign x_506 = ((((v_58 | ~v_24) | v_100) | v_114) | v_134) ;
	assign x_505 = ((((v_73 | ~v_50) | v_97) | v_139) | ~v_158) ;
	assign x_504 = ((((~v_67 | v_8) | v_85) | v_143) | v_116) ;
	assign x_503 = ((((v_56 | ~v_66) | ~v_104) | v_173) | v_111) ;
	assign x_502 = ((((v_1 | ~v_36) | v_93) | ~v_118) | v_146) ;
	assign x_501 = ((((~v_61 | v_8) | v_88) | v_154) | v_114) ;
	assign x_500 = ((((v_71 | v_29) | ~v_110) | v_96) | v_151) ;
	assign x_499 = ((((v_60 | v_31) | ~v_96) | ~v_107) | v_137) ;
	assign x_1590 = (x_497 & x_498) ;
	assign x_496 = ((((v_66 | v_24) | ~v_176) | v_158) | v_172) ;
	assign x_495 = ((((~v_27 | v_5) | v_135) | v_138) | v_110) ;
	assign x_494 = ((((~v_20 | ~v_80) | v_107) | ~v_180) | v_156) ;
	assign x_493 = ((((v_50 | ~v_70) | v_92) | ~v_180) | ~v_129) ;
	assign x_492 = ((((~v_9 | v_69) | ~v_143) | v_171) | ~v_113) ;
	assign x_491 = ((((v_47 | v_27) | ~v_157) | ~v_159) | ~v_87) ;
	assign x_490 = ((((~v_76 | ~v_48) | v_140) | v_171) | v_172) ;
	assign x_489 = ((((v_79 | v_24) | v_163) | v_99) | v_87) ;
	assign x_488 = ((((~v_47 | v_58) | ~v_89) | v_137) | ~v_171) ;
	assign x_487 = ((((~v_49 | ~v_10) | v_164) | v_112) | v_168) ;
	assign x_486 = ((((~v_41 | ~v_71) | v_119) | v_111) | v_158) ;
	assign x_485 = ((((~v_4 | ~v_69) | ~v_115) | ~v_81) | v_91) ;
	assign x_484 = ((((v_30 | v_79) | v_131) | ~v_151) | ~v_127) ;
	assign x_483 = ((((~v_43 | v_67) | ~v_170) | ~v_173) | v_162) ;
	assign x_482 = ((((~v_30 | ~v_21) | v_100) | ~v_147) | ~v_157) ;
	assign x_1572 = (x_480 & x_481) ;
	assign x_479 = ((((~v_56 | ~v_79) | v_156) | v_174) | v_175) ;
	assign x_478 = ((((v_36 | v_64) | v_158) | v_86) | ~v_123) ;
	assign x_477 = ((((v_73 | ~v_79) | ~v_98) | v_94) | ~v_111) ;
	assign x_476 = ((((v_37 | v_75) | ~v_83) | v_144) | v_146) ;
	assign x_475 = ((((v_1 | v_37) | ~v_127) | v_139) | v_110) ;
	assign x_474 = ((((~v_78 | v_33) | ~v_97) | ~v_167) | v_147) ;
	assign x_473 = ((((~v_7 | ~v_56) | v_100) | v_138) | v_103) ;
	assign x_1564 = (x_471 & x_472) ;
	assign x_470 = ((((v_32 | v_25) | v_113) | ~v_82) | v_150) ;
	assign x_469 = ((((~v_8 | ~v_43) | ~v_177) | v_114) | v_158) ;
	assign x_468 = ((((v_19 | ~v_8) | v_122) | ~v_117) | v_147) ;
	assign x_467 = ((((v_17 | v_40) | v_136) | ~v_168) | ~v_179) ;
	assign x_466 = ((((~v_22 | v_12) | ~v_86) | v_81) | v_161) ;
	assign x_465 = ((((v_58 | v_10) | v_135) | ~v_138) | v_130) ;
	assign x_464 = ((((~v_19 | v_62) | ~v_106) | v_154) | v_112) ;
	assign x_1555 = (x_462 & x_463) ;
	assign x_461 = ((((~v_31 | v_63) | v_117) | ~v_135) | v_153) ;
	assign x_460 = ((((~v_46 | v_22) | v_151) | v_173) | ~v_101) ;
	assign x_459 = ((((~v_15 | ~v_61) | v_147) | v_175) | v_114) ;
	assign x_458 = ((((~v_51 | v_41) | ~v_163) | v_164) | v_175) ;
	assign x_457 = ((((v_31 | v_16) | v_136) | v_173) | ~v_123) ;
	assign x_456 = ((((~v_37 | v_56) | ~v_127) | v_91) | ~v_87) ;
	assign x_455 = ((((~v_40 | v_34) | v_85) | ~v_126) | v_142) ;
	assign x_454 = ((((~v_56 | ~v_14) | ~v_167) | ~v_129) | v_138) ;
	assign x_453 = ((((v_28 | ~v_46) | v_167) | ~v_113) | ~v_121) ;
	assign x_452 = ((((v_19 | v_73) | ~v_173) | v_174) | ~v_136) ;
	assign x_451 = ((((v_2 | v_49) | ~v_100) | ~v_115) | v_137) ;
	assign x_450 = ((((v_73 | ~v_74) | v_93) | v_121) | v_174) ;
	assign x_449 = ((((~v_71 | v_5) | v_169) | v_133) | v_119) ;
	assign x_448 = ((((v_38 | v_58) | ~v_84) | v_92) | v_83) ;
	assign x_447 = ((((v_74 | ~v_27) | v_87) | ~v_137) | v_141) ;
	assign x_1538 = (x_445 & x_446) ;
	assign x_444 = ((((~v_19 | v_22) | v_172) | v_81) | v_151) ;
	assign x_443 = ((((~v_75 | ~v_29) | ~v_155) | v_93) | v_173) ;
	assign x_442 = ((((~v_5 | v_42) | ~v_165) | v_138) | v_133) ;
	assign x_441 = ((((v_58 | v_4) | ~v_111) | v_180) | ~v_100) ;
	assign x_440 = ((((~v_39 | v_25) | ~v_155) | v_92) | ~v_140) ;
	assign x_439 = ((((v_20 | v_75) | v_82) | ~v_111) | v_117) ;
	assign x_438 = ((((v_1 | v_69) | v_92) | ~v_116) | ~v_119) ;
	assign x_437 = ((((v_58 | ~v_40) | v_176) | v_168) | ~v_142) ;
	assign x_436 = ((((~v_53 | v_42) | ~v_111) | ~v_88) | ~v_149) ;
	assign x_435 = ((((v_10 | ~v_26) | ~v_93) | ~v_168) | ~v_160) ;
	assign x_434 = ((((~v_64 | v_26) | v_114) | v_119) | ~v_152) ;
	assign x_433 = ((((~v_40 | v_71) | ~v_97) | ~v_153) | v_129) ;
	assign x_432 = ((((v_80 | ~v_41) | ~v_153) | v_89) | ~v_122) ;
	assign x_431 = ((((v_25 | v_78) | ~v_116) | ~v_165) | v_153) ;
	assign x_430 = ((((v_80 | v_64) | v_119) | v_138) | v_133) ;
	assign x_1522 = (x_428 & x_429) ;
	assign x_427 = ((((~v_60 | ~v_33) | v_116) | v_115) | v_158) ;
	assign x_426 = ((((v_16 | v_76) | ~v_154) | ~v_103) | ~v_151) ;
	assign x_425 = ((((v_11 | v_46) | ~v_88) | ~v_111) | v_140) ;
	assign x_424 = ((((~v_49 | v_62) | ~v_115) | v_164) | ~v_156) ;
	assign x_423 = ((((v_65 | ~v_70) | v_173) | ~v_81) | v_112) ;
	assign x_422 = ((((~v_20 | ~v_61) | v_165) | ~v_159) | v_86) ;
	assign x_421 = ((((v_78 | v_24) | ~v_101) | v_129) | ~v_125) ;
	assign x_420 = ((((v_64 | v_29) | ~v_129) | v_125) | ~v_113) ;
	assign x_419 = ((((~v_43 | ~v_72) | ~v_120) | v_129) | v_126) ;
	assign x_418 = ((((v_66 | v_2) | v_142) | ~v_98) | v_95) ;
	assign x_417 = ((((~v_64 | ~v_4) | ~v_135) | v_81) | ~v_87) ;
	assign x_416 = ((((v_75 | v_40) | ~v_96) | v_138) | v_152) ;
	assign x_415 = ((((v_29 | ~v_51) | ~v_148) | v_141) | v_118) ;
	assign x_414 = ((((v_74 | v_7) | v_156) | ~v_95) | v_165) ;
	assign x_413 = ((((~v_2 | v_10) | v_164) | ~v_118) | ~v_121) ;
	assign x_1503 = (x_411 & x_412) ;
	assign x_410 = ((((~v_16 | ~v_29) | ~v_122) | v_172) | v_169) ;
	assign x_409 = ((((~v_62 | v_5) | v_104) | v_141) | ~v_129) ;
	assign x_408 = ((((v_8 | v_7) | v_174) | ~v_118) | v_164) ;
	assign x_407 = ((((~v_43 | ~v_41) | v_160) | v_106) | ~v_158) ;
	assign x_406 = ((((~v_46 | v_4) | v_125) | ~v_99) | ~v_180) ;
	assign x_405 = ((((v_58 | ~v_62) | ~v_154) | ~v_171) | ~v_143) ;
	assign x_404 = ((((~v_51 | v_60) | ~v_130) | ~v_88) | ~v_131) ;
	assign x_1495 = (x_402 & x_403) ;
	assign x_401 = ((((v_9 | ~v_21) | ~v_157) | ~v_121) | v_165) ;
	assign x_400 = ((((v_21 | v_29) | ~v_138) | v_122) | v_174) ;
	assign x_399 = ((((v_66 | v_42) | ~v_128) | v_163) | ~v_119) ;
	assign x_398 = ((((v_33 | v_55) | ~v_159) | v_176) | ~v_125) ;
	assign x_397 = ((((~v_26 | v_69) | ~v_125) | v_148) | v_99) ;
	assign x_396 = ((((~v_79 | ~v_46) | v_146) | ~v_93) | v_145) ;
	assign x_395 = ((((~v_39 | ~v_8) | ~v_148) | v_176) | ~v_119) ;
	assign x_1486 = (x_393 & x_394) ;
	assign x_392 = ((((v_11 | v_6) | v_171) | ~v_93) | ~v_144) ;
	assign x_391 = ((((~v_63 | v_33) | ~v_115) | v_113) | ~v_106) ;
	assign x_390 = ((((~v_46 | ~v_8) | v_121) | ~v_95) | ~v_147) ;
	assign x_389 = ((((v_54 | v_38) | v_121) | v_132) | ~v_122) ;
	assign x_388 = ((((~v_41 | ~v_21) | ~v_173) | ~v_156) | v_123) ;
	assign x_387 = ((((v_48 | ~v_8) | v_136) | v_175) | v_120) ;
	assign x_386 = ((((~v_23 | ~v_10) | ~v_88) | ~v_174) | v_121) ;
	assign x_385 = ((((v_45 | ~v_74) | ~v_86) | ~v_152) | v_117) ;
	assign x_384 = ((((~v_27 | v_41) | v_169) | v_132) | ~v_157) ;
	assign x_383 = ((((~v_1 | ~v_34) | ~v_95) | ~v_135) | v_144) ;
	assign x_382 = ((((v_52 | ~v_79) | v_164) | ~v_142) | ~v_141) ;
	assign x_381 = ((((v_43 | v_5) | v_150) | ~v_151) | v_116) ;
	assign x_380 = ((((~v_5 | ~v_13) | v_144) | v_153) | ~v_121) ;
	assign x_379 = ((((~v_71 | ~v_69) | v_143) | v_114) | ~v_174) ;
	assign x_378 = ((((v_63 | v_54) | ~v_145) | ~v_143) | ~v_138) ;
	assign x_1469 = (x_376 & x_377) ;
	assign x_375 = ((((~v_28 | v_72) | v_175) | v_91) | v_109) ;
	assign x_374 = ((((~v_9 | ~v_48) | ~v_177) | v_169) | ~v_122) ;
	assign x_373 = ((((v_80 | ~v_20) | ~v_137) | v_123) | v_114) ;
	assign x_372 = ((((~v_15 | v_34) | v_120) | ~v_179) | v_105) ;
	assign x_371 = ((((v_51 | v_30) | v_128) | v_112) | ~v_147) ;
	assign x_370 = ((((v_5 | v_37) | v_108) | ~v_144) | v_104) ;
	assign x_369 = ((((v_59 | ~v_63) | v_136) | v_130) | v_140) ;
	assign x_368 = ((((~v_39 | v_29) | ~v_112) | ~v_154) | v_92) ;
	assign x_367 = ((((~v_41 | v_11) | ~v_95) | v_132) | ~v_114) ;
	assign x_366 = ((((~v_10 | v_58) | v_88) | ~v_107) | ~v_109) ;
	assign x_365 = ((((v_12 | ~v_4) | ~v_153) | ~v_148) | ~v_93) ;
	assign x_364 = ((((v_55 | v_12) | ~v_157) | ~v_109) | ~v_144) ;
	assign x_363 = ((((v_26 | v_56) | ~v_154) | v_83) | ~v_109) ;
	assign x_362 = ((((v_24 | ~v_38) | v_164) | ~v_100) | v_145) ;
	assign x_361 = ((((~v_60 | ~v_9) | ~v_158) | ~v_115) | v_82) ;
	assign x_1453 = (x_359 & x_360) ;
	assign x_358 = ((((v_46 | ~v_47) | ~v_96) | v_143) | ~v_159) ;
	assign x_357 = ((((~v_52 | ~v_47) | ~v_110) | ~v_141) | v_168) ;
	assign x_356 = ((((v_75 | v_31) | ~v_88) | ~v_84) | v_110) ;
	assign x_355 = ((((v_28 | ~v_14) | v_180) | ~v_122) | v_142) ;
	assign x_354 = ((((~v_32 | ~v_66) | v_133) | v_115) | v_153) ;
	assign x_353 = ((((~v_22 | ~v_46) | v_102) | ~v_117) | v_158) ;
	assign x_352 = ((((v_16 | v_26) | v_106) | ~v_92) | v_122) ;
	assign x_351 = ((((v_39 | v_2) | v_133) | v_177) | v_173) ;
	assign x_350 = ((((v_51 | v_25) | v_132) | v_158) | v_116) ;
	assign x_349 = ((((v_46 | ~v_62) | v_177) | ~v_176) | ~v_134) ;
	assign x_348 = ((((~v_15 | ~v_35) | v_125) | ~v_135) | v_118) ;
	assign x_347 = ((((~v_15 | v_21) | v_109) | ~v_155) | v_159) ;
	assign x_346 = ((((v_78 | ~v_2) | v_83) | v_129) | ~v_118) ;
	assign x_345 = ((((v_43 | ~v_45) | ~v_93) | v_127) | ~v_161) ;
	assign x_344 = ((((~v_36 | v_18) | ~v_137) | ~v_150) | v_108) ;
	assign x_1435 = (x_342 & x_343) ;
	assign x_341 = ((((v_34 | ~v_40) | ~v_125) | ~v_89) | v_146) ;
	assign x_340 = ((((~v_8 | v_54) | ~v_143) | v_113) | ~v_144) ;
	assign x_339 = ((((~v_4 | ~v_52) | v_147) | ~v_113) | v_121) ;
	assign x_338 = ((((~v_23 | v_74) | v_115) | ~v_82) | ~v_141) ;
	assign x_337 = ((((v_9 | ~v_60) | ~v_117) | v_105) | ~v_126) ;
	assign x_336 = ((((~v_20 | v_61) | ~v_129) | ~v_170) | ~v_124) ;
	assign x_335 = ((((v_71 | v_6) | v_125) | ~v_104) | ~v_117) ;
	assign x_334 = ((((v_55 | v_70) | v_145) | ~v_130) | ~v_91) ;
	assign x_333 = ((((v_80 | v_38) | v_168) | ~v_98) | v_89) ;
	assign x_332 = ((((~v_2 | ~v_80) | ~v_128) | v_89) | v_110) ;
	assign x_331 = ((((~v_28 | ~v_70) | v_93) | v_170) | v_178) ;
	assign x_330 = ((((~v_61 | ~v_70) | ~v_109) | v_82) | v_162) ;
	assign x_329 = ((((v_76 | ~v_64) | ~v_88) | ~v_99) | ~v_142) ;
	assign x_328 = ((((v_15 | ~v_70) | v_113) | v_114) | v_151) ;
	assign x_327 = ((((v_66 | ~v_50) | ~v_108) | ~v_165) | v_138) ;
	assign x_1419 = (x_325 & x_326) ;
	assign x_324 = ((((v_1 | ~v_31) | ~v_104) | ~v_154) | v_107) ;
	assign x_323 = ((((~v_7 | v_10) | v_168) | ~v_99) | ~v_112) ;
	assign x_322 = ((((v_74 | v_10) | v_93) | ~v_162) | v_152) ;
	assign x_321 = ((((v_13 | v_28) | v_126) | ~v_113) | ~v_167) ;
	assign x_320 = ((((v_28 | ~v_63) | v_103) | ~v_85) | ~v_131) ;
	assign x_319 = ((((~v_68 | ~v_20) | ~v_110) | v_172) | v_152) ;
	assign x_318 = ((((v_53 | v_54) | ~v_139) | ~v_132) | v_140) ;
	assign x_317 = ((((~v_11 | v_16) | v_120) | v_155) | v_163) ;
	assign x_316 = ((((v_24 | ~v_50) | ~v_112) | v_92) | v_136) ;
	assign x_315 = ((((~v_3 | ~v_61) | ~v_108) | ~v_91) | v_92) ;
	assign x_314 = ((((~v_11 | ~v_72) | v_144) | v_145) | v_126) ;
	assign x_313 = ((((v_62 | ~v_28) | v_92) | ~v_143) | ~v_105) ;
	assign x_312 = ((((v_1 | ~v_40) | ~v_164) | ~v_114) | ~v_127) ;
	assign x_311 = ((((~v_27 | v_35) | v_178) | v_172) | v_168) ;
	assign x_310 = ((((v_18 | v_63) | v_98) | ~v_159) | v_157) ;
	assign x_1402 = (x_308 & x_309) ;
	assign x_307 = ((((~v_34 | ~v_80) | ~v_105) | v_170) | ~v_146) ;
	assign x_306 = ((((~v_24 | ~v_47) | v_176) | ~v_179) | ~v_151) ;
	assign x_305 = ((((~v_45 | v_12) | ~v_174) | ~v_140) | ~v_148) ;
	assign x_304 = ((((~v_6 | v_56) | v_93) | ~v_88) | ~v_165) ;
	assign x_303 = ((((~v_21 | ~v_43) | ~v_127) | ~v_171) | v_104) ;
	assign x_302 = ((((v_40 | v_31) | ~v_90) | v_123) | v_118) ;
	assign x_301 = ((((v_30 | v_63) | ~v_96) | ~v_163) | ~v_148) ;
	assign x_300 = ((((~v_29 | v_12) | v_100) | v_153) | v_132) ;
	assign x_299 = ((((v_65 | v_8) | v_109) | ~v_91) | v_104) ;
	assign x_298 = ((((~v_71 | ~v_66) | v_92) | v_134) | v_167) ;
	assign x_297 = ((((~v_6 | ~v_34) | v_93) | v_174) | ~v_162) ;
	assign x_296 = ((((v_66 | ~v_20) | ~v_162) | v_87) | ~v_128) ;
	assign x_295 = ((((~v_30 | ~v_71) | ~v_113) | v_138) | ~v_100) ;
	assign x_294 = ((((~v_37 | ~v_49) | v_145) | v_179) | ~v_134) ;
	assign x_293 = ((((~v_11 | v_17) | ~v_115) | v_81) | v_172) ;
	assign x_1386 = (x_291 & x_292) ;
	assign x_290 = ((((v_38 | ~v_32) | v_95) | v_147) | ~v_145) ;
	assign x_289 = ((((~v_50 | ~v_44) | v_151) | v_161) | v_116) ;
	assign x_288 = ((((v_33 | v_16) | ~v_172) | v_161) | v_178) ;
	assign x_287 = ((((~v_34 | ~v_40) | v_140) | ~v_143) | ~v_157) ;
	assign x_286 = ((((v_20 | v_8) | ~v_91) | ~v_85) | v_120) ;
	assign x_285 = ((((v_8 | ~v_5) | v_139) | v_141) | v_97) ;
	assign x_284 = ((((~v_64 | ~v_41) | ~v_142) | ~v_84) | v_114) ;
	assign x_283 = ((((v_33 | v_41) | ~v_102) | ~v_107) | ~v_87) ;
	assign x_282 = ((((v_77 | ~v_41) | ~v_134) | ~v_155) | v_143) ;
	assign x_281 = ((((v_25 | ~v_43) | ~v_150) | ~v_162) | v_149) ;
	assign x_280 = ((((~v_45 | ~v_2) | ~v_95) | ~v_146) | ~v_114) ;
	assign x_279 = ((((~v_45 | ~v_62) | v_105) | ~v_103) | ~v_151) ;
	assign x_278 = ((((v_77 | v_56) | ~v_176) | ~v_170) | ~v_122) ;
	assign x_277 = ((((v_30 | v_25) | ~v_110) | v_129) | v_175) ;
	assign x_276 = ((((v_70 | ~v_58) | v_175) | v_105) | ~v_136) ;
	assign x_1366 = (x_274 & x_275) ;
	assign x_273 = ((((v_23 | v_13) | v_133) | ~v_154) | ~v_81) ;
	assign x_272 = ((((~v_40 | v_28) | ~v_118) | ~v_167) | ~v_154) ;
	assign x_271 = ((((~v_9 | v_66) | ~v_83) | ~v_128) | ~v_177) ;
	assign x_270 = ((((v_36 | v_34) | v_177) | ~v_133) | v_155) ;
	assign x_269 = ((((~v_19 | ~v_29) | v_134) | ~v_157) | v_162) ;
	assign x_268 = ((((~v_76 | ~v_56) | ~v_116) | ~v_141) | ~v_148) ;
	assign x_267 = ((((~v_63 | ~v_16) | ~v_112) | ~v_174) | v_111) ;
	assign x_1358 = (x_265 & x_266) ;
	assign x_264 = ((((v_16 | ~v_78) | v_130) | v_124) | v_178) ;
	assign x_263 = ((((v_64 | ~v_13) | ~v_109) | v_116) | ~v_152) ;
	assign x_262 = ((((v_44 | ~v_64) | v_170) | v_157) | v_84) ;
	assign x_261 = ((((~v_72 | v_6) | ~v_106) | v_121) | ~v_119) ;
	assign x_260 = ((((~v_29 | v_18) | v_105) | v_158) | ~v_178) ;
	assign x_259 = ((((v_37 | v_23) | v_162) | v_135) | v_126) ;
	assign x_258 = ((((~v_24 | ~v_2) | v_107) | ~v_161) | v_132) ;
	assign x_1349 = (x_256 & x_257) ;
	assign x_255 = ((((v_3 | v_79) | ~v_110) | v_122) | ~v_128) ;
	assign x_254 = ((((~v_64 | ~v_80) | ~v_139) | ~v_150) | ~v_119) ;
	assign x_253 = ((((v_77 | v_39) | v_180) | ~v_150) | v_163) ;
	assign x_252 = ((((v_16 | v_56) | ~v_177) | v_178) | v_161) ;
	assign x_251 = ((((v_57 | v_36) | ~v_142) | v_156) | v_161) ;
	assign x_250 = ((((v_38 | ~v_73) | ~v_92) | ~v_87) | ~v_96) ;
	assign x_249 = ((((~v_61 | v_69) | v_150) | ~v_105) | v_159) ;
	assign x_248 = ((((v_70 | ~v_17) | ~v_176) | v_97) | ~v_148) ;
	assign x_247 = ((((~v_9 | v_2) | ~v_145) | ~v_83) | v_174) ;
	assign x_246 = ((((v_45 | v_44) | ~v_177) | v_157) | ~v_151) ;
	assign x_245 = ((((~v_37 | v_31) | ~v_158) | v_93) | v_151) ;
	assign x_244 = ((((v_8 | ~v_19) | ~v_120) | v_175) | v_119) ;
	assign x_243 = ((((~v_12 | v_32) | v_123) | ~v_138) | ~v_165) ;
	assign x_242 = ((((v_22 | ~v_59) | ~v_119) | v_165) | ~v_167) ;
	assign x_241 = ((((~v_15 | v_76) | v_178) | v_85) | v_155) ;
	assign x_1332 = (x_239 & x_240) ;
	assign x_238 = ((((v_41 | ~v_57) | v_95) | ~v_128) | v_113) ;
	assign x_237 = ((((v_4 | v_9) | v_144) | v_173) | ~v_128) ;
	assign x_236 = ((((~v_54 | v_10) | v_93) | v_157) | ~v_136) ;
	assign x_235 = ((((~v_54 | ~v_68) | v_138) | ~v_157) | v_177) ;
	assign x_234 = ((((~v_68 | v_16) | ~v_115) | ~v_110) | v_177) ;
	assign x_233 = ((((v_57 | ~v_66) | ~v_95) | ~v_85) | v_150) ;
	assign x_232 = ((((~v_8 | v_41) | ~v_112) | v_140) | v_123) ;
	assign x_231 = ((((~v_48 | v_3) | v_105) | v_164) | ~v_88) ;
	assign x_230 = ((((v_58 | ~v_41) | ~v_144) | ~v_173) | ~v_135) ;
	assign x_229 = ((((~v_10 | ~v_40) | ~v_117) | v_128) | ~v_142) ;
	assign x_228 = ((((v_31 | ~v_43) | v_136) | v_101) | v_102) ;
	assign x_227 = ((((~v_45 | ~v_6) | ~v_127) | v_107) | ~v_172) ;
	assign x_226 = ((((~v_42 | v_34) | ~v_114) | v_96) | v_122) ;
	assign x_225 = ((((~v_25 | ~v_5) | v_111) | ~v_132) | v_85) ;
	assign x_224 = ((((v_24 | v_39) | ~v_140) | v_130) | ~v_82) ;
	assign x_1316 = (x_222 & x_223) ;
	assign x_221 = ((((~v_23 | ~v_28) | v_95) | ~v_155) | ~v_117) ;
	assign x_220 = ((((v_55 | ~v_28) | v_161) | ~v_129) | ~v_128) ;
	assign x_219 = ((((~v_40 | v_35) | ~v_102) | ~v_110) | ~v_112) ;
	assign x_218 = ((((v_27 | ~v_75) | ~v_147) | ~v_160) | ~v_88) ;
	assign x_217 = ((((v_17 | ~v_30) | v_173) | v_139) | v_110) ;
	assign x_216 = ((((~v_24 | v_78) | ~v_124) | ~v_116) | ~v_174) ;
	assign x_215 = ((((~v_73 | ~v_46) | v_122) | ~v_141) | ~v_143) ;
	assign x_214 = ((((v_49 | v_65) | ~v_135) | ~v_104) | v_150) ;
	assign x_213 = ((((v_13 | v_78) | v_90) | ~v_92) | ~v_102) ;
	assign x_212 = ((((~v_32 | ~v_29) | ~v_178) | ~v_142) | v_128) ;
	assign x_211 = ((((v_41 | v_62) | ~v_137) | v_140) | ~v_149) ;
	assign x_210 = ((((~v_56 | v_40) | v_99) | ~v_132) | ~v_96) ;
	assign x_209 = ((((v_9 | v_41) | ~v_174) | ~v_168) | ~v_179) ;
	assign x_208 = ((((~v_4 | v_53) | ~v_117) | v_118) | v_175) ;
	assign x_207 = ((((~v_71 | ~v_77) | v_82) | v_159) | v_163) ;
	assign x_1298 = (x_205 & x_206) ;
	assign x_204 = ((((~v_7 | ~v_6) | v_103) | ~v_156) | v_112) ;
	assign x_203 = ((((v_38 | ~v_18) | v_90) | v_159) | v_88) ;
	assign x_202 = ((((v_16 | ~v_27) | ~v_87) | v_86) | v_127) ;
	assign x_201 = ((((v_63 | v_10) | v_131) | v_174) | ~v_117) ;
	assign x_200 = ((((v_68 | ~v_26) | v_96) | v_90) | v_107) ;
	assign x_199 = ((((v_48 | ~v_69) | v_112) | v_87) | ~v_109) ;
	assign x_198 = ((((~v_78 | v_37) | ~v_139) | ~v_84) | ~v_90) ;
	assign x_1290 = (x_196 & x_197) ;
	assign x_195 = ((((~v_16 | ~v_48) | v_175) | ~v_126) | ~v_92) ;
	assign x_194 = ((((~v_64 | ~v_66) | v_162) | v_107) | ~v_125) ;
	assign x_193 = ((((~v_16 | ~v_70) | ~v_149) | v_171) | ~v_83) ;
	assign x_192 = ((((v_35 | v_61) | v_99) | ~v_157) | v_152) ;
	assign x_191 = ((((~v_27 | v_5) | ~v_89) | v_140) | ~v_117) ;
	assign x_190 = ((((~v_12 | ~v_57) | ~v_134) | ~v_90) | ~v_82) ;
	assign x_189 = ((((~v_79 | ~v_27) | ~v_128) | ~v_97) | v_99) ;
	assign x_1281 = (x_187 & x_188) ;
	assign x_186 = ((((~v_12 | ~v_24) | v_90) | v_149) | v_171) ;
	assign x_185 = ((((~v_64 | v_25) | v_97) | ~v_122) | v_179) ;
	assign x_184 = ((((~v_36 | v_25) | ~v_122) | ~v_133) | ~v_129) ;
	assign x_183 = ((((v_38 | v_67) | v_83) | v_169) | v_175) ;
	assign x_182 = ((((v_37 | v_60) | ~v_136) | v_85) | ~v_110) ;
	assign x_181 = ((((v_15 | v_9) | v_142) | ~v_176) | ~v_149) ;
	assign x_180 = ((((v_57 | ~v_52) | ~v_142) | v_99) | ~v_179) ;
	assign x_179 = ((((~v_77 | v_31) | v_148) | v_83) | ~v_87) ;
	assign x_178 = ((((~v_74 | v_35) | ~v_136) | ~v_129) | ~v_89) ;
	assign x_177 = ((((v_3 | ~v_46) | ~v_113) | v_107) | v_91) ;
	assign x_176 = ((((v_13 | ~v_72) | v_142) | ~v_146) | v_130) ;
	assign x_175 = ((((v_10 | ~v_44) | v_151) | v_96) | ~v_118) ;
	assign x_174 = ((((v_50 | ~v_44) | ~v_115) | v_158) | ~v_113) ;
	assign x_173 = ((((v_25 | v_2) | v_94) | v_125) | v_134) ;
	assign x_172 = ((((~v_53 | ~v_63) | v_119) | ~v_92) | v_149) ;
	assign x_1264 = (x_170 & x_171) ;
	assign x_169 = ((((v_55 | ~v_59) | v_92) | ~v_154) | ~v_107) ;
	assign x_168 = ((((~v_10 | ~v_24) | v_93) | ~v_147) | v_97) ;
	assign x_167 = ((((v_15 | ~v_35) | v_109) | ~v_160) | ~v_177) ;
	assign x_166 = ((((v_68 | v_14) | v_160) | v_117) | ~v_168) ;
	assign x_165 = ((((~v_5 | ~v_3) | ~v_83) | ~v_133) | v_136) ;
	assign x_164 = ((((~v_61 | ~v_5) | v_128) | ~v_162) | v_170) ;
	assign x_163 = ((((~v_40 | v_3) | v_161) | v_166) | v_88) ;
	assign x_162 = ((((~v_53 | v_2) | v_81) | v_132) | ~v_115) ;
	assign x_161 = ((((~v_49 | ~v_37) | v_87) | ~v_140) | ~v_150) ;
	assign x_160 = ((((v_70 | v_38) | v_104) | ~v_109) | v_96) ;
	assign x_159 = ((((~v_42 | ~v_7) | v_174) | v_170) | ~v_117) ;
	assign x_158 = ((((v_77 | v_29) | v_134) | ~v_97) | v_91) ;
	assign x_157 = ((((v_66 | ~v_41) | ~v_165) | v_109) | ~v_134) ;
	assign x_156 = ((((~v_52 | v_32) | ~v_118) | v_103) | ~v_115) ;
	assign x_155 = ((((v_79 | ~v_31) | v_167) | v_168) | v_106) ;
	assign x_1248 = (x_153 & x_154) ;
	assign x_152 = ((((v_18 | v_24) | v_89) | ~v_123) | v_85) ;
	assign x_151 = ((((~v_28 | ~v_48) | v_87) | ~v_101) | v_94) ;
	assign x_150 = ((((~v_47 | v_7) | v_112) | v_179) | v_110) ;
	assign x_149 = ((((~v_56 | ~v_48) | v_132) | v_84) | ~v_180) ;
	assign x_148 = ((((~v_60 | ~v_46) | v_155) | ~v_162) | ~v_111) ;
	assign x_147 = ((((~v_37 | v_10) | ~v_148) | v_152) | v_113) ;
	assign x_146 = ((((v_4 | v_21) | ~v_145) | v_114) | ~v_139) ;
	assign x_145 = ((((~v_21 | ~v_23) | v_142) | v_141) | ~v_168) ;
	assign x_144 = ((((~v_64 | ~v_76) | v_100) | v_122) | ~v_172) ;
	assign x_143 = ((((v_49 | v_52) | v_138) | v_136) | ~v_92) ;
	assign x_142 = ((((~v_6 | v_55) | v_116) | v_104) | ~v_125) ;
	assign x_141 = ((((~v_49 | ~v_52) | ~v_174) | ~v_94) | v_90) ;
	assign x_140 = ((((v_35 | v_14) | v_90) | ~v_174) | ~v_169) ;
	assign x_139 = ((((~v_4 | ~v_70) | v_166) | v_145) | v_103) ;
	assign x_138 = ((((v_63 | v_65) | ~v_171) | ~v_176) | v_159) ;
	assign x_1229 = (x_136 & x_137) ;
	assign x_135 = ((((~v_17 | v_37) | ~v_161) | v_138) | v_157) ;
	assign x_134 = ((((~v_53 | v_4) | v_152) | v_104) | ~v_82) ;
	assign x_133 = ((((v_38 | v_65) | ~v_89) | ~v_81) | ~v_132) ;
	assign x_132 = ((((~v_18 | ~v_14) | ~v_94) | v_123) | v_168) ;
	assign x_131 = ((((~v_49 | v_35) | v_114) | ~v_127) | ~v_118) ;
	assign x_130 = ((((~v_64 | v_7) | ~v_175) | ~v_179) | ~v_128) ;
	assign x_129 = ((((v_13 | v_56) | v_101) | ~v_164) | ~v_173) ;
	assign x_1221 = (x_127 & x_128) ;
	assign x_126 = ((((~v_75 | ~v_67) | v_141) | v_112) | ~v_135) ;
	assign x_125 = ((((v_69 | v_52) | v_105) | v_145) | ~v_134) ;
	assign x_124 = ((((v_53 | ~v_25) | v_85) | v_154) | v_104) ;
	assign x_123 = ((((v_20 | ~v_41) | ~v_163) | ~v_112) | ~v_116) ;
	assign x_122 = ((((~v_72 | v_6) | ~v_131) | v_139) | ~v_145) ;
	assign x_121 = ((((~v_72 | v_65) | v_180) | v_148) | v_145) ;
	assign x_120 = ((((v_48 | ~v_49) | ~v_147) | ~v_94) | ~v_152) ;
	assign x_1212 = (x_118 & x_119) ;
	assign x_117 = ((((~v_52 | ~v_21) | ~v_147) | v_117) | v_93) ;
	assign x_116 = ((((~v_51 | v_20) | v_171) | v_175) | ~v_176) ;
	assign x_115 = ((((~v_22 | v_47) | v_173) | v_120) | ~v_123) ;
	assign x_114 = ((((v_17 | v_75) | v_115) | v_138) | ~v_81) ;
	assign x_113 = ((((~v_48 | ~v_69) | v_124) | v_154) | ~v_91) ;
	assign x_112 = ((((~v_45 | v_62) | ~v_112) | ~v_108) | v_150) ;
	assign x_111 = ((((v_34 | ~v_46) | ~v_113) | v_140) | ~v_139) ;
	assign x_110 = ((((~v_76 | ~v_11) | ~v_110) | v_155) | ~v_122) ;
	assign x_109 = ((((~v_66 | ~v_21) | v_101) | ~v_99) | ~v_164) ;
	assign x_108 = ((((v_78 | v_10) | v_108) | v_122) | v_138) ;
	assign x_107 = ((((v_46 | ~v_17) | v_145) | ~v_140) | v_94) ;
	assign x_106 = ((((v_27 | v_26) | v_81) | ~v_142) | ~v_179) ;
	assign x_105 = ((((~v_15 | ~v_57) | v_175) | ~v_178) | ~v_89) ;
	assign x_104 = ((((v_52 | v_40) | v_133) | ~v_124) | ~v_123) ;
	assign x_103 = ((((v_28 | v_2) | ~v_94) | ~v_86) | v_175) ;
	assign x_1195 = (x_101 & x_102) ;
	assign x_100 = ((((~v_51 | v_31) | v_112) | v_137) | ~v_86) ;
	assign x_99 = ((((~v_31 | ~v_61) | ~v_156) | ~v_177) | ~v_125) ;
	assign x_98 = ((((v_74 | ~v_15) | v_122) | ~v_137) | ~v_89) ;
	assign x_97 = ((((v_12 | ~v_17) | ~v_178) | ~v_162) | ~v_122) ;
	assign x_96 = ((((~v_26 | ~v_80) | v_88) | ~v_86) | ~v_95) ;
	assign x_95 = ((((v_57 | ~v_27) | v_176) | v_145) | ~v_123) ;
	assign x_94 = ((((~v_34 | v_58) | ~v_118) | v_101) | ~v_137) ;
	assign x_93 = ((((~v_76 | ~v_79) | ~v_114) | ~v_124) | ~v_104) ;
	assign x_92 = ((((v_22 | ~v_18) | ~v_95) | v_93) | ~v_100) ;
	assign x_91 = ((((~v_6 | v_34) | v_82) | ~v_155) | v_127) ;
	assign x_90 = ((((v_54 | v_38) | v_130) | ~v_136) | v_118) ;
	assign x_89 = ((((v_52 | v_61) | ~v_154) | v_153) | ~v_134) ;
	assign x_88 = ((((v_70 | ~v_8) | ~v_95) | v_169) | v_97) ;
	assign x_87 = ((((~v_65 | ~v_51) | ~v_96) | ~v_159) | ~v_148) ;
	assign x_86 = ((((v_37 | v_73) | v_173) | v_171) | v_180) ;
	assign x_1179 = (x_84 & x_85) ;
	assign x_83 = ((((~v_39 | ~v_71) | ~v_114) | v_124) | ~v_127) ;
	assign x_82 = ((((~v_20 | ~v_76) | ~v_85) | v_132) | ~v_144) ;
	assign x_81 = ((((v_77 | v_58) | ~v_144) | ~v_103) | ~v_109) ;
	assign x_80 = ((((~v_30 | v_53) | v_155) | v_104) | ~v_164) ;
	assign x_79 = ((((v_54 | v_24) | ~v_93) | v_111) | v_83) ;
	assign x_78 = ((((v_56 | v_3) | ~v_96) | ~v_119) | ~v_105) ;
	assign x_77 = ((((v_10 | v_30) | v_155) | ~v_104) | ~v_130) ;
	assign x_76 = ((((v_58 | v_34) | ~v_94) | ~v_106) | v_180) ;
	assign x_75 = ((((v_53 | v_67) | ~v_133) | v_173) | ~v_93) ;
	assign x_74 = ((((~v_26 | v_31) | ~v_161) | ~v_151) | v_165) ;
	assign x_73 = ((((~v_71 | v_56) | v_98) | ~v_143) | v_96) ;
	assign x_72 = ((((v_12 | ~v_68) | v_178) | v_144) | ~v_135) ;
	assign x_71 = ((((v_16 | ~v_34) | v_166) | v_157) | v_86) ;
	assign x_70 = ((((~v_1 | v_53) | ~v_155) | ~v_164) | ~v_176) ;
	assign x_69 = ((((v_74 | ~v_6) | ~v_96) | v_97) | v_137) ;
	assign x_1161 = (x_67 & x_68) ;
	assign x_66 = ((((~v_20 | ~v_17) | v_152) | v_95) | v_140) ;
	assign x_65 = ((((~v_31 | v_70) | v_119) | v_170) | ~v_84) ;
	assign x_64 = ((((~v_55 | ~v_15) | ~v_175) | v_119) | ~v_97) ;
	assign x_63 = ((((~v_28 | v_60) | ~v_169) | ~v_162) | ~v_96) ;
	assign x_62 = ((((~v_21 | v_72) | v_102) | v_157) | v_114) ;
	assign x_61 = ((((v_13 | v_80) | v_128) | ~v_133) | ~v_85) ;
	assign x_60 = ((((~v_8 | v_4) | v_179) | ~v_114) | v_118) ;
	assign x_59 = ((((~v_41 | ~v_14) | ~v_133) | ~v_134) | ~v_162) ;
	assign x_58 = ((((v_14 | ~v_48) | v_92) | v_128) | v_127) ;
	assign x_57 = ((((v_35 | ~v_42) | ~v_112) | v_154) | v_160) ;
	assign x_56 = ((((v_2 | ~v_19) | ~v_136) | ~v_82) | ~v_105) ;
	assign x_55 = ((((~v_1 | ~v_11) | v_120) | ~v_132) | ~v_143) ;
	assign x_54 = ((((~v_59 | ~v_35) | v_125) | v_126) | v_172) ;
	assign x_53 = ((((v_56 | ~v_37) | ~v_121) | ~v_127) | ~v_154) ;
	assign x_52 = ((((v_5 | v_64) | ~v_131) | v_109) | ~v_148) ;
	assign x_1145 = (x_50 & x_51) ;
	assign x_49 = ((((v_70 | v_68) | ~v_111) | v_153) | ~v_117) ;
	assign x_48 = ((((v_51 | ~v_61) | ~v_95) | v_123) | v_115) ;
	assign x_47 = ((((~v_79 | v_17) | v_137) | v_146) | ~v_171) ;
	assign x_46 = ((((~v_44 | ~v_26) | ~v_128) | ~v_143) | ~v_118) ;
	assign x_45 = ((((v_25 | v_41) | ~v_92) | v_102) | v_172) ;
	assign x_44 = ((((~v_78 | v_17) | ~v_98) | v_121) | ~v_143) ;
	assign x_43 = ((((v_25 | v_24) | v_90) | ~v_161) | v_115) ;
	assign x_42 = ((((v_68 | ~v_1) | ~v_106) | ~v_93) | ~v_85) ;
	assign x_41 = ((((~v_45 | v_80) | v_97) | ~v_106) | v_133) ;
	assign x_40 = ((((v_14 | v_58) | ~v_170) | ~v_132) | v_157) ;
	assign x_39 = ((((~v_52 | ~v_21) | v_162) | ~v_177) | ~v_110) ;
	assign x_38 = ((((v_10 | v_72) | ~v_172) | ~v_87) | v_122) ;
	assign x_37 = ((((~v_70 | v_72) | ~v_137) | v_112) | v_102) ;
	assign x_36 = ((((v_62 | v_56) | v_159) | ~v_173) | v_155) ;
	assign x_35 = ((((~v_73 | v_75) | ~v_155) | v_138) | v_162) ;
	assign x_1128 = (x_33 & x_34) ;
	assign x_32 = ((((~v_25 | v_39) | ~v_132) | ~v_152) | ~v_112) ;
	assign x_31 = ((((v_20 | ~v_44) | v_127) | v_158) | ~v_166) ;
	assign x_30 = ((((~v_45 | ~v_75) | ~v_155) | v_121) | v_113) ;
	assign x_29 = ((((v_33 | v_5) | ~v_158) | v_169) | ~v_122) ;
	assign x_28 = ((((v_56 | v_62) | ~v_144) | ~v_167) | v_113) ;
	assign x_27 = ((((~v_63 | v_37) | v_155) | ~v_161) | ~v_123) ;
	assign x_26 = ((((v_50 | ~v_27) | ~v_94) | v_108) | ~v_128) ;
	assign x_25 = ((((~v_65 | v_64) | v_94) | ~v_105) | ~v_175) ;
	assign x_24 = ((((v_2 | v_3) | v_123) | v_122) | v_126) ;
	assign x_23 = ((((~v_52 | v_55) | ~v_172) | v_107) | v_92) ;
	assign x_22 = ((((v_32 | v_43) | v_124) | ~v_100) | ~v_85) ;
	assign x_21 = ((((~v_49 | ~v_67) | v_151) | v_109) | v_98) ;
	assign x_20 = ((((~v_44 | v_41) | v_138) | v_107) | ~v_143) ;
	assign x_19 = ((((~v_63 | ~v_8) | v_172) | v_89) | v_135) ;
	assign x_18 = ((((v_32 | v_77) | v_83) | ~v_115) | ~v_163) ;
	assign x_1112 = (x_16 & x_17) ;
	assign x_15 = ((((v_23 | ~v_68) | v_94) | v_134) | v_106) ;
	assign x_14 = ((((~v_42 | ~v_66) | ~v_156) | v_161) | v_152) ;
	assign x_13 = ((((v_56 | ~v_79) | ~v_180) | ~v_125) | ~v_147) ;
	assign x_12 = ((((~v_20 | v_73) | v_149) | v_154) | ~v_176) ;
	assign x_11 = ((((v_2 | ~v_66) | v_129) | v_170) | ~v_120) ;
	assign x_10 = ((((~v_10 | v_70) | v_140) | v_148) | ~v_162) ;
	assign x_9 = ((((~v_78 | ~v_22) | ~v_136) | ~v_155) | ~v_129) ;
	assign x_8 = ((((~v_53 | ~v_14) | v_137) | v_140) | v_121) ;
	assign x_7 = ((((~v_70 | v_2) | v_151) | v_90) | ~v_145) ;
	assign x_6 = ((((v_23 | ~v_22) | ~v_152) | ~v_174) | v_138) ;
	assign x_5 = ((((v_36 | v_61) | v_126) | ~v_170) | v_134) ;
	assign x_4 = ((((~v_16 | ~v_43) | ~v_111) | ~v_149) | v_174) ;
	assign x_3 = ((((~v_22 | ~v_3) | v_141) | v_94) | v_85) ;
	assign x_2 = ((((v_74 | v_52) | ~v_128) | ~v_125) | ~v_141) ;
	assign x_1 = ((((v_24 | ~v_56) | ~v_85) | v_126) | v_147) ;
	assign x_2190 = (x_1098 & x_2189) ;
	assign x_2188 = (x_1096 & x_1097) ;
	assign x_2186 = (x_1094 & x_1095) ;
	assign x_2185 = (x_1092 & x_1093) ;
	assign x_2182 = (x_1089 & x_2181) ;
	assign x_2180 = (x_1087 & x_1088) ;
	assign x_2178 = (x_1085 & x_1086) ;
	assign x_2177 = (x_1083 & x_1084) ;
	assign x_2173 = (x_1080 & x_2172) ;
	assign x_2171 = (x_1078 & x_1079) ;
	assign x_2169 = (x_1076 & x_1077) ;
	assign x_2168 = (x_1074 & x_1075) ;
	assign x_2165 = (x_1072 & x_1073) ;
	assign x_2164 = (x_1070 & x_1071) ;
	assign x_2162 = (x_1068 & x_1069) ;
	assign x_2161 = (x_1066 & x_1067) ;
	assign x_2156 = (x_1063 & x_2155) ;
	assign x_2154 = (x_1061 & x_1062) ;
	assign x_2152 = (x_1059 & x_1060) ;
	assign x_2151 = (x_1057 & x_1058) ;
	assign x_2148 = (x_1055 & x_1056) ;
	assign x_2147 = (x_1053 & x_1054) ;
	assign x_2145 = (x_1051 & x_1052) ;
	assign x_2144 = (x_1049 & x_1050) ;
	assign x_2140 = (x_1046 & x_2139) ;
	assign x_2138 = (x_1044 & x_1045) ;
	assign x_2136 = (x_1042 & x_1043) ;
	assign x_2135 = (x_1040 & x_1041) ;
	assign x_2132 = (x_1038 & x_1039) ;
	assign x_2131 = (x_1036 & x_1037) ;
	assign x_2129 = (x_1034 & x_1035) ;
	assign x_2128 = (x_1032 & x_1033) ;
	assign x_2122 = (x_1029 & x_2121) ;
	assign x_2120 = (x_1027 & x_1028) ;
	assign x_2118 = (x_1025 & x_1026) ;
	assign x_2117 = (x_1023 & x_1024) ;
	assign x_2114 = (x_1020 & x_2113) ;
	assign x_2112 = (x_1018 & x_1019) ;
	assign x_2110 = (x_1016 & x_1017) ;
	assign x_2109 = (x_1014 & x_1015) ;
	assign x_2105 = (x_1011 & x_2104) ;
	assign x_2103 = (x_1009 & x_1010) ;
	assign x_2101 = (x_1007 & x_1008) ;
	assign x_2100 = (x_1005 & x_1006) ;
	assign x_2097 = (x_1003 & x_1004) ;
	assign x_2096 = (x_1001 & x_1002) ;
	assign x_2094 = (x_999 & x_1000) ;
	assign x_2093 = (x_997 & x_998) ;
	assign x_2088 = (x_994 & x_2087) ;
	assign x_2086 = (x_992 & x_993) ;
	assign x_2084 = (x_990 & x_991) ;
	assign x_2083 = (x_988 & x_989) ;
	assign x_2080 = (x_986 & x_987) ;
	assign x_2079 = (x_984 & x_985) ;
	assign x_2077 = (x_982 & x_983) ;
	assign x_2076 = (x_980 & x_981) ;
	assign x_2072 = (x_977 & x_2071) ;
	assign x_2070 = (x_975 & x_976) ;
	assign x_2068 = (x_973 & x_974) ;
	assign x_2067 = (x_971 & x_972) ;
	assign x_2064 = (x_969 & x_970) ;
	assign x_2063 = (x_967 & x_968) ;
	assign x_2061 = (x_965 & x_966) ;
	assign x_2060 = (x_963 & x_964) ;
	assign x_2053 = (x_960 & x_2052) ;
	assign x_2051 = (x_958 & x_959) ;
	assign x_2049 = (x_956 & x_957) ;
	assign x_2048 = (x_954 & x_955) ;
	assign x_2045 = (x_951 & x_2044) ;
	assign x_2043 = (x_949 & x_950) ;
	assign x_2041 = (x_947 & x_948) ;
	assign x_2040 = (x_945 & x_946) ;
	assign x_2036 = (x_942 & x_2035) ;
	assign x_2034 = (x_940 & x_941) ;
	assign x_2032 = (x_938 & x_939) ;
	assign x_2031 = (x_936 & x_937) ;
	assign x_2028 = (x_934 & x_935) ;
	assign x_2027 = (x_932 & x_933) ;
	assign x_2025 = (x_930 & x_931) ;
	assign x_2024 = (x_928 & x_929) ;
	assign x_2019 = (x_925 & x_2018) ;
	assign x_2017 = (x_923 & x_924) ;
	assign x_2015 = (x_921 & x_922) ;
	assign x_2014 = (x_919 & x_920) ;
	assign x_2011 = (x_917 & x_918) ;
	assign x_2010 = (x_915 & x_916) ;
	assign x_2008 = (x_913 & x_914) ;
	assign x_2007 = (x_911 & x_912) ;
	assign x_2003 = (x_908 & x_2002) ;
	assign x_2001 = (x_906 & x_907) ;
	assign x_1999 = (x_904 & x_905) ;
	assign x_1998 = (x_902 & x_903) ;
	assign x_1995 = (x_900 & x_901) ;
	assign x_1994 = (x_898 & x_899) ;
	assign x_1992 = (x_896 & x_897) ;
	assign x_1991 = (x_894 & x_895) ;
	assign x_1985 = (x_891 & x_1984) ;
	assign x_1983 = (x_889 & x_890) ;
	assign x_1981 = (x_887 & x_888) ;
	assign x_1980 = (x_885 & x_886) ;
	assign x_1977 = (x_883 & x_884) ;
	assign x_1976 = (x_881 & x_882) ;
	assign x_1974 = (x_879 & x_880) ;
	assign x_1973 = (x_877 & x_878) ;
	assign x_1969 = (x_874 & x_1968) ;
	assign x_1967 = (x_872 & x_873) ;
	assign x_1965 = (x_870 & x_871) ;
	assign x_1964 = (x_868 & x_869) ;
	assign x_1961 = (x_866 & x_867) ;
	assign x_1960 = (x_864 & x_865) ;
	assign x_1958 = (x_862 & x_863) ;
	assign x_1957 = (x_860 & x_861) ;
	assign x_1952 = (x_857 & x_1951) ;
	assign x_1950 = (x_855 & x_856) ;
	assign x_1948 = (x_853 & x_854) ;
	assign x_1947 = (x_851 & x_852) ;
	assign x_1944 = (x_849 & x_850) ;
	assign x_1943 = (x_847 & x_848) ;
	assign x_1941 = (x_845 & x_846) ;
	assign x_1940 = (x_843 & x_844) ;
	assign x_1936 = (x_840 & x_1935) ;
	assign x_1934 = (x_838 & x_839) ;
	assign x_1932 = (x_836 & x_837) ;
	assign x_1931 = (x_834 & x_835) ;
	assign x_1928 = (x_832 & x_833) ;
	assign x_1927 = (x_830 & x_831) ;
	assign x_1925 = (x_828 & x_829) ;
	assign x_1924 = (x_826 & x_827) ;
	assign x_1916 = (x_823 & x_1915) ;
	assign x_1914 = (x_821 & x_822) ;
	assign x_1912 = (x_819 & x_820) ;
	assign x_1911 = (x_817 & x_818) ;
	assign x_1908 = (x_814 & x_1907) ;
	assign x_1906 = (x_812 & x_813) ;
	assign x_1904 = (x_810 & x_811) ;
	assign x_1903 = (x_808 & x_809) ;
	assign x_1899 = (x_805 & x_1898) ;
	assign x_1897 = (x_803 & x_804) ;
	assign x_1895 = (x_801 & x_802) ;
	assign x_1894 = (x_799 & x_800) ;
	assign x_1891 = (x_797 & x_798) ;
	assign x_1890 = (x_795 & x_796) ;
	assign x_1888 = (x_793 & x_794) ;
	assign x_1887 = (x_791 & x_792) ;
	assign x_1882 = (x_788 & x_1881) ;
	assign x_1880 = (x_786 & x_787) ;
	assign x_1878 = (x_784 & x_785) ;
	assign x_1877 = (x_782 & x_783) ;
	assign x_1874 = (x_780 & x_781) ;
	assign x_1873 = (x_778 & x_779) ;
	assign x_1871 = (x_776 & x_777) ;
	assign x_1870 = (x_774 & x_775) ;
	assign x_1866 = (x_771 & x_1865) ;
	assign x_1864 = (x_769 & x_770) ;
	assign x_1862 = (x_767 & x_768) ;
	assign x_1861 = (x_765 & x_766) ;
	assign x_1858 = (x_763 & x_764) ;
	assign x_1857 = (x_761 & x_762) ;
	assign x_1855 = (x_759 & x_760) ;
	assign x_1854 = (x_757 & x_758) ;
	assign x_1848 = (x_754 & x_1847) ;
	assign x_1846 = (x_752 & x_753) ;
	assign x_1844 = (x_750 & x_751) ;
	assign x_1843 = (x_748 & x_749) ;
	assign x_1840 = (x_745 & x_1839) ;
	assign x_1838 = (x_743 & x_744) ;
	assign x_1836 = (x_741 & x_742) ;
	assign x_1835 = (x_739 & x_740) ;
	assign x_1831 = (x_736 & x_1830) ;
	assign x_1829 = (x_734 & x_735) ;
	assign x_1827 = (x_732 & x_733) ;
	assign x_1826 = (x_730 & x_731) ;
	assign x_1823 = (x_728 & x_729) ;
	assign x_1822 = (x_726 & x_727) ;
	assign x_1820 = (x_724 & x_725) ;
	assign x_1819 = (x_722 & x_723) ;
	assign x_1814 = (x_719 & x_1813) ;
	assign x_1812 = (x_717 & x_718) ;
	assign x_1810 = (x_715 & x_716) ;
	assign x_1809 = (x_713 & x_714) ;
	assign x_1806 = (x_711 & x_712) ;
	assign x_1805 = (x_709 & x_710) ;
	assign x_1803 = (x_707 & x_708) ;
	assign x_1802 = (x_705 & x_706) ;
	assign x_1798 = (x_702 & x_1797) ;
	assign x_1796 = (x_700 & x_701) ;
	assign x_1794 = (x_698 & x_699) ;
	assign x_1793 = (x_696 & x_697) ;
	assign x_1790 = (x_694 & x_695) ;
	assign x_1789 = (x_692 & x_693) ;
	assign x_1787 = (x_690 & x_691) ;
	assign x_1786 = (x_688 & x_689) ;
	assign x_1779 = (x_685 & x_1778) ;
	assign x_1777 = (x_683 & x_684) ;
	assign x_1775 = (x_681 & x_682) ;
	assign x_1774 = (x_679 & x_680) ;
	assign x_1771 = (x_676 & x_1770) ;
	assign x_1769 = (x_674 & x_675) ;
	assign x_1767 = (x_672 & x_673) ;
	assign x_1766 = (x_670 & x_671) ;
	assign x_1762 = (x_667 & x_1761) ;
	assign x_1760 = (x_665 & x_666) ;
	assign x_1758 = (x_663 & x_664) ;
	assign x_1757 = (x_661 & x_662) ;
	assign x_1754 = (x_659 & x_660) ;
	assign x_1753 = (x_657 & x_658) ;
	assign x_1751 = (x_655 & x_656) ;
	assign x_1750 = (x_653 & x_654) ;
	assign x_1745 = (x_650 & x_1744) ;
	assign x_1743 = (x_648 & x_649) ;
	assign x_1741 = (x_646 & x_647) ;
	assign x_1740 = (x_644 & x_645) ;
	assign x_1737 = (x_642 & x_643) ;
	assign x_1736 = (x_640 & x_641) ;
	assign x_1734 = (x_638 & x_639) ;
	assign x_1733 = (x_636 & x_637) ;
	assign x_1729 = (x_633 & x_1728) ;
	assign x_1727 = (x_631 & x_632) ;
	assign x_1725 = (x_629 & x_630) ;
	assign x_1724 = (x_627 & x_628) ;
	assign x_1721 = (x_625 & x_626) ;
	assign x_1720 = (x_623 & x_624) ;
	assign x_1718 = (x_621 & x_622) ;
	assign x_1717 = (x_619 & x_620) ;
	assign x_1711 = (x_616 & x_1710) ;
	assign x_1709 = (x_614 & x_615) ;
	assign x_1707 = (x_612 & x_613) ;
	assign x_1706 = (x_610 & x_611) ;
	assign x_1703 = (x_608 & x_609) ;
	assign x_1702 = (x_606 & x_607) ;
	assign x_1700 = (x_604 & x_605) ;
	assign x_1699 = (x_602 & x_603) ;
	assign x_1695 = (x_599 & x_1694) ;
	assign x_1693 = (x_597 & x_598) ;
	assign x_1691 = (x_595 & x_596) ;
	assign x_1690 = (x_593 & x_594) ;
	assign x_1687 = (x_591 & x_592) ;
	assign x_1686 = (x_589 & x_590) ;
	assign x_1684 = (x_587 & x_588) ;
	assign x_1683 = (x_585 & x_586) ;
	assign x_1678 = (x_582 & x_1677) ;
	assign x_1676 = (x_580 & x_581) ;
	assign x_1674 = (x_578 & x_579) ;
	assign x_1673 = (x_576 & x_577) ;
	assign x_1670 = (x_574 & x_575) ;
	assign x_1669 = (x_572 & x_573) ;
	assign x_1667 = (x_570 & x_571) ;
	assign x_1666 = (x_568 & x_569) ;
	assign x_1662 = (x_565 & x_1661) ;
	assign x_1660 = (x_563 & x_564) ;
	assign x_1658 = (x_561 & x_562) ;
	assign x_1657 = (x_559 & x_560) ;
	assign x_1654 = (x_557 & x_558) ;
	assign x_1653 = (x_555 & x_556) ;
	assign x_1651 = (x_553 & x_554) ;
	assign x_1650 = (x_551 & x_552) ;
	assign x_1641 = (x_548 & x_1640) ;
	assign x_1639 = (x_546 & x_547) ;
	assign x_1637 = (x_544 & x_545) ;
	assign x_1636 = (x_542 & x_543) ;
	assign x_1633 = (x_539 & x_1632) ;
	assign x_1631 = (x_537 & x_538) ;
	assign x_1629 = (x_535 & x_536) ;
	assign x_1628 = (x_533 & x_534) ;
	assign x_1624 = (x_530 & x_1623) ;
	assign x_1622 = (x_528 & x_529) ;
	assign x_1620 = (x_526 & x_527) ;
	assign x_1619 = (x_524 & x_525) ;
	assign x_1616 = (x_522 & x_523) ;
	assign x_1615 = (x_520 & x_521) ;
	assign x_1613 = (x_518 & x_519) ;
	assign x_1612 = (x_516 & x_517) ;
	assign x_1607 = (x_513 & x_1606) ;
	assign x_1605 = (x_511 & x_512) ;
	assign x_1603 = (x_509 & x_510) ;
	assign x_1602 = (x_507 & x_508) ;
	assign x_1599 = (x_505 & x_506) ;
	assign x_1598 = (x_503 & x_504) ;
	assign x_1596 = (x_501 & x_502) ;
	assign x_1595 = (x_499 & x_500) ;
	assign x_1591 = (x_496 & x_1590) ;
	assign x_1589 = (x_494 & x_495) ;
	assign x_1587 = (x_492 & x_493) ;
	assign x_1586 = (x_490 & x_491) ;
	assign x_1583 = (x_488 & x_489) ;
	assign x_1582 = (x_486 & x_487) ;
	assign x_1580 = (x_484 & x_485) ;
	assign x_1579 = (x_482 & x_483) ;
	assign x_1573 = (x_479 & x_1572) ;
	assign x_1571 = (x_477 & x_478) ;
	assign x_1569 = (x_475 & x_476) ;
	assign x_1568 = (x_473 & x_474) ;
	assign x_1565 = (x_470 & x_1564) ;
	assign x_1563 = (x_468 & x_469) ;
	assign x_1561 = (x_466 & x_467) ;
	assign x_1560 = (x_464 & x_465) ;
	assign x_1556 = (x_461 & x_1555) ;
	assign x_1554 = (x_459 & x_460) ;
	assign x_1552 = (x_457 & x_458) ;
	assign x_1551 = (x_455 & x_456) ;
	assign x_1548 = (x_453 & x_454) ;
	assign x_1547 = (x_451 & x_452) ;
	assign x_1545 = (x_449 & x_450) ;
	assign x_1544 = (x_447 & x_448) ;
	assign x_1539 = (x_444 & x_1538) ;
	assign x_1537 = (x_442 & x_443) ;
	assign x_1535 = (x_440 & x_441) ;
	assign x_1534 = (x_438 & x_439) ;
	assign x_1531 = (x_436 & x_437) ;
	assign x_1530 = (x_434 & x_435) ;
	assign x_1528 = (x_432 & x_433) ;
	assign x_1527 = (x_430 & x_431) ;
	assign x_1523 = (x_427 & x_1522) ;
	assign x_1521 = (x_425 & x_426) ;
	assign x_1519 = (x_423 & x_424) ;
	assign x_1518 = (x_421 & x_422) ;
	assign x_1515 = (x_419 & x_420) ;
	assign x_1514 = (x_417 & x_418) ;
	assign x_1512 = (x_415 & x_416) ;
	assign x_1511 = (x_413 & x_414) ;
	assign x_1504 = (x_410 & x_1503) ;
	assign x_1502 = (x_408 & x_409) ;
	assign x_1500 = (x_406 & x_407) ;
	assign x_1499 = (x_404 & x_405) ;
	assign x_1496 = (x_401 & x_1495) ;
	assign x_1494 = (x_399 & x_400) ;
	assign x_1492 = (x_397 & x_398) ;
	assign x_1491 = (x_395 & x_396) ;
	assign x_1487 = (x_392 & x_1486) ;
	assign x_1485 = (x_390 & x_391) ;
	assign x_1483 = (x_388 & x_389) ;
	assign x_1482 = (x_386 & x_387) ;
	assign x_1479 = (x_384 & x_385) ;
	assign x_1478 = (x_382 & x_383) ;
	assign x_1476 = (x_380 & x_381) ;
	assign x_1475 = (x_378 & x_379) ;
	assign x_1470 = (x_375 & x_1469) ;
	assign x_1468 = (x_373 & x_374) ;
	assign x_1466 = (x_371 & x_372) ;
	assign x_1465 = (x_369 & x_370) ;
	assign x_1462 = (x_367 & x_368) ;
	assign x_1461 = (x_365 & x_366) ;
	assign x_1459 = (x_363 & x_364) ;
	assign x_1458 = (x_361 & x_362) ;
	assign x_1454 = (x_358 & x_1453) ;
	assign x_1452 = (x_356 & x_357) ;
	assign x_1450 = (x_354 & x_355) ;
	assign x_1449 = (x_352 & x_353) ;
	assign x_1446 = (x_350 & x_351) ;
	assign x_1445 = (x_348 & x_349) ;
	assign x_1443 = (x_346 & x_347) ;
	assign x_1442 = (x_344 & x_345) ;
	assign x_1436 = (x_341 & x_1435) ;
	assign x_1434 = (x_339 & x_340) ;
	assign x_1432 = (x_337 & x_338) ;
	assign x_1431 = (x_335 & x_336) ;
	assign x_1428 = (x_333 & x_334) ;
	assign x_1427 = (x_331 & x_332) ;
	assign x_1425 = (x_329 & x_330) ;
	assign x_1424 = (x_327 & x_328) ;
	assign x_1420 = (x_324 & x_1419) ;
	assign x_1418 = (x_322 & x_323) ;
	assign x_1416 = (x_320 & x_321) ;
	assign x_1415 = (x_318 & x_319) ;
	assign x_1412 = (x_316 & x_317) ;
	assign x_1411 = (x_314 & x_315) ;
	assign x_1409 = (x_312 & x_313) ;
	assign x_1408 = (x_310 & x_311) ;
	assign x_1403 = (x_307 & x_1402) ;
	assign x_1401 = (x_305 & x_306) ;
	assign x_1399 = (x_303 & x_304) ;
	assign x_1398 = (x_301 & x_302) ;
	assign x_1395 = (x_299 & x_300) ;
	assign x_1394 = (x_297 & x_298) ;
	assign x_1392 = (x_295 & x_296) ;
	assign x_1391 = (x_293 & x_294) ;
	assign x_1387 = (x_290 & x_1386) ;
	assign x_1385 = (x_288 & x_289) ;
	assign x_1383 = (x_286 & x_287) ;
	assign x_1382 = (x_284 & x_285) ;
	assign x_1379 = (x_282 & x_283) ;
	assign x_1378 = (x_280 & x_281) ;
	assign x_1376 = (x_278 & x_279) ;
	assign x_1375 = (x_276 & x_277) ;
	assign x_1367 = (x_273 & x_1366) ;
	assign x_1365 = (x_271 & x_272) ;
	assign x_1363 = (x_269 & x_270) ;
	assign x_1362 = (x_267 & x_268) ;
	assign x_1359 = (x_264 & x_1358) ;
	assign x_1357 = (x_262 & x_263) ;
	assign x_1355 = (x_260 & x_261) ;
	assign x_1354 = (x_258 & x_259) ;
	assign x_1350 = (x_255 & x_1349) ;
	assign x_1348 = (x_253 & x_254) ;
	assign x_1346 = (x_251 & x_252) ;
	assign x_1345 = (x_249 & x_250) ;
	assign x_1342 = (x_247 & x_248) ;
	assign x_1341 = (x_245 & x_246) ;
	assign x_1339 = (x_243 & x_244) ;
	assign x_1338 = (x_241 & x_242) ;
	assign x_1333 = (x_238 & x_1332) ;
	assign x_1331 = (x_236 & x_237) ;
	assign x_1329 = (x_234 & x_235) ;
	assign x_1328 = (x_232 & x_233) ;
	assign x_1325 = (x_230 & x_231) ;
	assign x_1324 = (x_228 & x_229) ;
	assign x_1322 = (x_226 & x_227) ;
	assign x_1321 = (x_224 & x_225) ;
	assign x_1317 = (x_221 & x_1316) ;
	assign x_1315 = (x_219 & x_220) ;
	assign x_1313 = (x_217 & x_218) ;
	assign x_1312 = (x_215 & x_216) ;
	assign x_1309 = (x_213 & x_214) ;
	assign x_1308 = (x_211 & x_212) ;
	assign x_1306 = (x_209 & x_210) ;
	assign x_1305 = (x_207 & x_208) ;
	assign x_1299 = (x_204 & x_1298) ;
	assign x_1297 = (x_202 & x_203) ;
	assign x_1295 = (x_200 & x_201) ;
	assign x_1294 = (x_198 & x_199) ;
	assign x_1291 = (x_195 & x_1290) ;
	assign x_1289 = (x_193 & x_194) ;
	assign x_1287 = (x_191 & x_192) ;
	assign x_1286 = (x_189 & x_190) ;
	assign x_1282 = (x_186 & x_1281) ;
	assign x_1280 = (x_184 & x_185) ;
	assign x_1278 = (x_182 & x_183) ;
	assign x_1277 = (x_180 & x_181) ;
	assign x_1274 = (x_178 & x_179) ;
	assign x_1273 = (x_176 & x_177) ;
	assign x_1271 = (x_174 & x_175) ;
	assign x_1270 = (x_172 & x_173) ;
	assign x_1265 = (x_169 & x_1264) ;
	assign x_1263 = (x_167 & x_168) ;
	assign x_1261 = (x_165 & x_166) ;
	assign x_1260 = (x_163 & x_164) ;
	assign x_1257 = (x_161 & x_162) ;
	assign x_1256 = (x_159 & x_160) ;
	assign x_1254 = (x_157 & x_158) ;
	assign x_1253 = (x_155 & x_156) ;
	assign x_1249 = (x_152 & x_1248) ;
	assign x_1247 = (x_150 & x_151) ;
	assign x_1245 = (x_148 & x_149) ;
	assign x_1244 = (x_146 & x_147) ;
	assign x_1241 = (x_144 & x_145) ;
	assign x_1240 = (x_142 & x_143) ;
	assign x_1238 = (x_140 & x_141) ;
	assign x_1237 = (x_138 & x_139) ;
	assign x_1230 = (x_135 & x_1229) ;
	assign x_1228 = (x_133 & x_134) ;
	assign x_1226 = (x_131 & x_132) ;
	assign x_1225 = (x_129 & x_130) ;
	assign x_1222 = (x_126 & x_1221) ;
	assign x_1220 = (x_124 & x_125) ;
	assign x_1218 = (x_122 & x_123) ;
	assign x_1217 = (x_120 & x_121) ;
	assign x_1213 = (x_117 & x_1212) ;
	assign x_1211 = (x_115 & x_116) ;
	assign x_1209 = (x_113 & x_114) ;
	assign x_1208 = (x_111 & x_112) ;
	assign x_1205 = (x_109 & x_110) ;
	assign x_1204 = (x_107 & x_108) ;
	assign x_1202 = (x_105 & x_106) ;
	assign x_1201 = (x_103 & x_104) ;
	assign x_1196 = (x_100 & x_1195) ;
	assign x_1194 = (x_98 & x_99) ;
	assign x_1192 = (x_96 & x_97) ;
	assign x_1191 = (x_94 & x_95) ;
	assign x_1188 = (x_92 & x_93) ;
	assign x_1187 = (x_90 & x_91) ;
	assign x_1185 = (x_88 & x_89) ;
	assign x_1184 = (x_86 & x_87) ;
	assign x_1180 = (x_83 & x_1179) ;
	assign x_1178 = (x_81 & x_82) ;
	assign x_1176 = (x_79 & x_80) ;
	assign x_1175 = (x_77 & x_78) ;
	assign x_1172 = (x_75 & x_76) ;
	assign x_1171 = (x_73 & x_74) ;
	assign x_1169 = (x_71 & x_72) ;
	assign x_1168 = (x_69 & x_70) ;
	assign x_1162 = (x_66 & x_1161) ;
	assign x_1160 = (x_64 & x_65) ;
	assign x_1158 = (x_62 & x_63) ;
	assign x_1157 = (x_60 & x_61) ;
	assign x_1154 = (x_58 & x_59) ;
	assign x_1153 = (x_56 & x_57) ;
	assign x_1151 = (x_54 & x_55) ;
	assign x_1150 = (x_52 & x_53) ;
	assign x_1146 = (x_49 & x_1145) ;
	assign x_1144 = (x_47 & x_48) ;
	assign x_1142 = (x_45 & x_46) ;
	assign x_1141 = (x_43 & x_44) ;
	assign x_1138 = (x_41 & x_42) ;
	assign x_1137 = (x_39 & x_40) ;
	assign x_1135 = (x_37 & x_38) ;
	assign x_1134 = (x_35 & x_36) ;
	assign x_1129 = (x_32 & x_1128) ;
	assign x_1127 = (x_30 & x_31) ;
	assign x_1125 = (x_28 & x_29) ;
	assign x_1124 = (x_26 & x_27) ;
	assign x_1121 = (x_24 & x_25) ;
	assign x_1120 = (x_22 & x_23) ;
	assign x_1118 = (x_20 & x_21) ;
	assign x_1117 = (x_18 & x_19) ;
	assign x_1113 = (x_15 & x_1112) ;
	assign x_1111 = (x_13 & x_14) ;
	assign x_1109 = (x_11 & x_12) ;
	assign x_1108 = (x_9 & x_10) ;
	assign x_1105 = (x_7 & x_8) ;
	assign x_1104 = (x_5 & x_6) ;
	assign x_1102 = (x_3 & x_4) ;
	assign x_1101 = (x_1 & x_2) ;
	assign x_2191 = (x_2188 & x_2190) ;
	assign x_2187 = (x_2185 & x_2186) ;
	assign x_2183 = (x_2180 & x_2182) ;
	assign x_2179 = (x_2177 & x_2178) ;
	assign x_2174 = (x_2171 & x_2173) ;
	assign x_2170 = (x_2168 & x_2169) ;
	assign x_2166 = (x_2164 & x_2165) ;
	assign x_2163 = (x_2161 & x_2162) ;
	assign x_2157 = (x_2154 & x_2156) ;
	assign x_2153 = (x_2151 & x_2152) ;
	assign x_2149 = (x_2147 & x_2148) ;
	assign x_2146 = (x_2144 & x_2145) ;
	assign x_2141 = (x_2138 & x_2140) ;
	assign x_2137 = (x_2135 & x_2136) ;
	assign x_2133 = (x_2131 & x_2132) ;
	assign x_2130 = (x_2128 & x_2129) ;
	assign x_2123 = (x_2120 & x_2122) ;
	assign x_2119 = (x_2117 & x_2118) ;
	assign x_2115 = (x_2112 & x_2114) ;
	assign x_2111 = (x_2109 & x_2110) ;
	assign x_2106 = (x_2103 & x_2105) ;
	assign x_2102 = (x_2100 & x_2101) ;
	assign x_2098 = (x_2096 & x_2097) ;
	assign x_2095 = (x_2093 & x_2094) ;
	assign x_2089 = (x_2086 & x_2088) ;
	assign x_2085 = (x_2083 & x_2084) ;
	assign x_2081 = (x_2079 & x_2080) ;
	assign x_2078 = (x_2076 & x_2077) ;
	assign x_2073 = (x_2070 & x_2072) ;
	assign x_2069 = (x_2067 & x_2068) ;
	assign x_2065 = (x_2063 & x_2064) ;
	assign x_2062 = (x_2060 & x_2061) ;
	assign x_2054 = (x_2051 & x_2053) ;
	assign x_2050 = (x_2048 & x_2049) ;
	assign x_2046 = (x_2043 & x_2045) ;
	assign x_2042 = (x_2040 & x_2041) ;
	assign x_2037 = (x_2034 & x_2036) ;
	assign x_2033 = (x_2031 & x_2032) ;
	assign x_2029 = (x_2027 & x_2028) ;
	assign x_2026 = (x_2024 & x_2025) ;
	assign x_2020 = (x_2017 & x_2019) ;
	assign x_2016 = (x_2014 & x_2015) ;
	assign x_2012 = (x_2010 & x_2011) ;
	assign x_2009 = (x_2007 & x_2008) ;
	assign x_2004 = (x_2001 & x_2003) ;
	assign x_2000 = (x_1998 & x_1999) ;
	assign x_1996 = (x_1994 & x_1995) ;
	assign x_1993 = (x_1991 & x_1992) ;
	assign x_1986 = (x_1983 & x_1985) ;
	assign x_1982 = (x_1980 & x_1981) ;
	assign x_1978 = (x_1976 & x_1977) ;
	assign x_1975 = (x_1973 & x_1974) ;
	assign x_1970 = (x_1967 & x_1969) ;
	assign x_1966 = (x_1964 & x_1965) ;
	assign x_1962 = (x_1960 & x_1961) ;
	assign x_1959 = (x_1957 & x_1958) ;
	assign x_1953 = (x_1950 & x_1952) ;
	assign x_1949 = (x_1947 & x_1948) ;
	assign x_1945 = (x_1943 & x_1944) ;
	assign x_1942 = (x_1940 & x_1941) ;
	assign x_1937 = (x_1934 & x_1936) ;
	assign x_1933 = (x_1931 & x_1932) ;
	assign x_1929 = (x_1927 & x_1928) ;
	assign x_1926 = (x_1924 & x_1925) ;
	assign x_1917 = (x_1914 & x_1916) ;
	assign x_1913 = (x_1911 & x_1912) ;
	assign x_1909 = (x_1906 & x_1908) ;
	assign x_1905 = (x_1903 & x_1904) ;
	assign x_1900 = (x_1897 & x_1899) ;
	assign x_1896 = (x_1894 & x_1895) ;
	assign x_1892 = (x_1890 & x_1891) ;
	assign x_1889 = (x_1887 & x_1888) ;
	assign x_1883 = (x_1880 & x_1882) ;
	assign x_1879 = (x_1877 & x_1878) ;
	assign x_1875 = (x_1873 & x_1874) ;
	assign x_1872 = (x_1870 & x_1871) ;
	assign x_1867 = (x_1864 & x_1866) ;
	assign x_1863 = (x_1861 & x_1862) ;
	assign x_1859 = (x_1857 & x_1858) ;
	assign x_1856 = (x_1854 & x_1855) ;
	assign x_1849 = (x_1846 & x_1848) ;
	assign x_1845 = (x_1843 & x_1844) ;
	assign x_1841 = (x_1838 & x_1840) ;
	assign x_1837 = (x_1835 & x_1836) ;
	assign x_1832 = (x_1829 & x_1831) ;
	assign x_1828 = (x_1826 & x_1827) ;
	assign x_1824 = (x_1822 & x_1823) ;
	assign x_1821 = (x_1819 & x_1820) ;
	assign x_1815 = (x_1812 & x_1814) ;
	assign x_1811 = (x_1809 & x_1810) ;
	assign x_1807 = (x_1805 & x_1806) ;
	assign x_1804 = (x_1802 & x_1803) ;
	assign x_1799 = (x_1796 & x_1798) ;
	assign x_1795 = (x_1793 & x_1794) ;
	assign x_1791 = (x_1789 & x_1790) ;
	assign x_1788 = (x_1786 & x_1787) ;
	assign x_1780 = (x_1777 & x_1779) ;
	assign x_1776 = (x_1774 & x_1775) ;
	assign x_1772 = (x_1769 & x_1771) ;
	assign x_1768 = (x_1766 & x_1767) ;
	assign x_1763 = (x_1760 & x_1762) ;
	assign x_1759 = (x_1757 & x_1758) ;
	assign x_1755 = (x_1753 & x_1754) ;
	assign x_1752 = (x_1750 & x_1751) ;
	assign x_1746 = (x_1743 & x_1745) ;
	assign x_1742 = (x_1740 & x_1741) ;
	assign x_1738 = (x_1736 & x_1737) ;
	assign x_1735 = (x_1733 & x_1734) ;
	assign x_1730 = (x_1727 & x_1729) ;
	assign x_1726 = (x_1724 & x_1725) ;
	assign x_1722 = (x_1720 & x_1721) ;
	assign x_1719 = (x_1717 & x_1718) ;
	assign x_1712 = (x_1709 & x_1711) ;
	assign x_1708 = (x_1706 & x_1707) ;
	assign x_1704 = (x_1702 & x_1703) ;
	assign x_1701 = (x_1699 & x_1700) ;
	assign x_1696 = (x_1693 & x_1695) ;
	assign x_1692 = (x_1690 & x_1691) ;
	assign x_1688 = (x_1686 & x_1687) ;
	assign x_1685 = (x_1683 & x_1684) ;
	assign x_1679 = (x_1676 & x_1678) ;
	assign x_1675 = (x_1673 & x_1674) ;
	assign x_1671 = (x_1669 & x_1670) ;
	assign x_1668 = (x_1666 & x_1667) ;
	assign x_1663 = (x_1660 & x_1662) ;
	assign x_1659 = (x_1657 & x_1658) ;
	assign x_1655 = (x_1653 & x_1654) ;
	assign x_1652 = (x_1650 & x_1651) ;
	assign x_1642 = (x_1639 & x_1641) ;
	assign x_1638 = (x_1636 & x_1637) ;
	assign x_1634 = (x_1631 & x_1633) ;
	assign x_1630 = (x_1628 & x_1629) ;
	assign x_1625 = (x_1622 & x_1624) ;
	assign x_1621 = (x_1619 & x_1620) ;
	assign x_1617 = (x_1615 & x_1616) ;
	assign x_1614 = (x_1612 & x_1613) ;
	assign x_1608 = (x_1605 & x_1607) ;
	assign x_1604 = (x_1602 & x_1603) ;
	assign x_1600 = (x_1598 & x_1599) ;
	assign x_1597 = (x_1595 & x_1596) ;
	assign x_1592 = (x_1589 & x_1591) ;
	assign x_1588 = (x_1586 & x_1587) ;
	assign x_1584 = (x_1582 & x_1583) ;
	assign x_1581 = (x_1579 & x_1580) ;
	assign x_1574 = (x_1571 & x_1573) ;
	assign x_1570 = (x_1568 & x_1569) ;
	assign x_1566 = (x_1563 & x_1565) ;
	assign x_1562 = (x_1560 & x_1561) ;
	assign x_1557 = (x_1554 & x_1556) ;
	assign x_1553 = (x_1551 & x_1552) ;
	assign x_1549 = (x_1547 & x_1548) ;
	assign x_1546 = (x_1544 & x_1545) ;
	assign x_1540 = (x_1537 & x_1539) ;
	assign x_1536 = (x_1534 & x_1535) ;
	assign x_1532 = (x_1530 & x_1531) ;
	assign x_1529 = (x_1527 & x_1528) ;
	assign x_1524 = (x_1521 & x_1523) ;
	assign x_1520 = (x_1518 & x_1519) ;
	assign x_1516 = (x_1514 & x_1515) ;
	assign x_1513 = (x_1511 & x_1512) ;
	assign x_1505 = (x_1502 & x_1504) ;
	assign x_1501 = (x_1499 & x_1500) ;
	assign x_1497 = (x_1494 & x_1496) ;
	assign x_1493 = (x_1491 & x_1492) ;
	assign x_1488 = (x_1485 & x_1487) ;
	assign x_1484 = (x_1482 & x_1483) ;
	assign x_1480 = (x_1478 & x_1479) ;
	assign x_1477 = (x_1475 & x_1476) ;
	assign x_1471 = (x_1468 & x_1470) ;
	assign x_1467 = (x_1465 & x_1466) ;
	assign x_1463 = (x_1461 & x_1462) ;
	assign x_1460 = (x_1458 & x_1459) ;
	assign x_1455 = (x_1452 & x_1454) ;
	assign x_1451 = (x_1449 & x_1450) ;
	assign x_1447 = (x_1445 & x_1446) ;
	assign x_1444 = (x_1442 & x_1443) ;
	assign x_1437 = (x_1434 & x_1436) ;
	assign x_1433 = (x_1431 & x_1432) ;
	assign x_1429 = (x_1427 & x_1428) ;
	assign x_1426 = (x_1424 & x_1425) ;
	assign x_1421 = (x_1418 & x_1420) ;
	assign x_1417 = (x_1415 & x_1416) ;
	assign x_1413 = (x_1411 & x_1412) ;
	assign x_1410 = (x_1408 & x_1409) ;
	assign x_1404 = (x_1401 & x_1403) ;
	assign x_1400 = (x_1398 & x_1399) ;
	assign x_1396 = (x_1394 & x_1395) ;
	assign x_1393 = (x_1391 & x_1392) ;
	assign x_1388 = (x_1385 & x_1387) ;
	assign x_1384 = (x_1382 & x_1383) ;
	assign x_1380 = (x_1378 & x_1379) ;
	assign x_1377 = (x_1375 & x_1376) ;
	assign x_1368 = (x_1365 & x_1367) ;
	assign x_1364 = (x_1362 & x_1363) ;
	assign x_1360 = (x_1357 & x_1359) ;
	assign x_1356 = (x_1354 & x_1355) ;
	assign x_1351 = (x_1348 & x_1350) ;
	assign x_1347 = (x_1345 & x_1346) ;
	assign x_1343 = (x_1341 & x_1342) ;
	assign x_1340 = (x_1338 & x_1339) ;
	assign x_1334 = (x_1331 & x_1333) ;
	assign x_1330 = (x_1328 & x_1329) ;
	assign x_1326 = (x_1324 & x_1325) ;
	assign x_1323 = (x_1321 & x_1322) ;
	assign x_1318 = (x_1315 & x_1317) ;
	assign x_1314 = (x_1312 & x_1313) ;
	assign x_1310 = (x_1308 & x_1309) ;
	assign x_1307 = (x_1305 & x_1306) ;
	assign x_1300 = (x_1297 & x_1299) ;
	assign x_1296 = (x_1294 & x_1295) ;
	assign x_1292 = (x_1289 & x_1291) ;
	assign x_1288 = (x_1286 & x_1287) ;
	assign x_1283 = (x_1280 & x_1282) ;
	assign x_1279 = (x_1277 & x_1278) ;
	assign x_1275 = (x_1273 & x_1274) ;
	assign x_1272 = (x_1270 & x_1271) ;
	assign x_1266 = (x_1263 & x_1265) ;
	assign x_1262 = (x_1260 & x_1261) ;
	assign x_1258 = (x_1256 & x_1257) ;
	assign x_1255 = (x_1253 & x_1254) ;
	assign x_1250 = (x_1247 & x_1249) ;
	assign x_1246 = (x_1244 & x_1245) ;
	assign x_1242 = (x_1240 & x_1241) ;
	assign x_1239 = (x_1237 & x_1238) ;
	assign x_1231 = (x_1228 & x_1230) ;
	assign x_1227 = (x_1225 & x_1226) ;
	assign x_1223 = (x_1220 & x_1222) ;
	assign x_1219 = (x_1217 & x_1218) ;
	assign x_1214 = (x_1211 & x_1213) ;
	assign x_1210 = (x_1208 & x_1209) ;
	assign x_1206 = (x_1204 & x_1205) ;
	assign x_1203 = (x_1201 & x_1202) ;
	assign x_1197 = (x_1194 & x_1196) ;
	assign x_1193 = (x_1191 & x_1192) ;
	assign x_1189 = (x_1187 & x_1188) ;
	assign x_1186 = (x_1184 & x_1185) ;
	assign x_1181 = (x_1178 & x_1180) ;
	assign x_1177 = (x_1175 & x_1176) ;
	assign x_1173 = (x_1171 & x_1172) ;
	assign x_1170 = (x_1168 & x_1169) ;
	assign x_1163 = (x_1160 & x_1162) ;
	assign x_1159 = (x_1157 & x_1158) ;
	assign x_1155 = (x_1153 & x_1154) ;
	assign x_1152 = (x_1150 & x_1151) ;
	assign x_1147 = (x_1144 & x_1146) ;
	assign x_1143 = (x_1141 & x_1142) ;
	assign x_1139 = (x_1137 & x_1138) ;
	assign x_1136 = (x_1134 & x_1135) ;
	assign x_1130 = (x_1127 & x_1129) ;
	assign x_1126 = (x_1124 & x_1125) ;
	assign x_1122 = (x_1120 & x_1121) ;
	assign x_1119 = (x_1117 & x_1118) ;
	assign x_1114 = (x_1111 & x_1113) ;
	assign x_1110 = (x_1108 & x_1109) ;
	assign x_1106 = (x_1104 & x_1105) ;
	assign x_1103 = (x_1101 & x_1102) ;
	assign x_2192 = (x_2187 & x_2191) ;
	assign x_2184 = (x_2179 & x_2183) ;
	assign x_2175 = (x_2170 & x_2174) ;
	assign x_2167 = (x_2163 & x_2166) ;
	assign x_2158 = (x_2153 & x_2157) ;
	assign x_2150 = (x_2146 & x_2149) ;
	assign x_2142 = (x_2137 & x_2141) ;
	assign x_2134 = (x_2130 & x_2133) ;
	assign x_2124 = (x_2119 & x_2123) ;
	assign x_2116 = (x_2111 & x_2115) ;
	assign x_2107 = (x_2102 & x_2106) ;
	assign x_2099 = (x_2095 & x_2098) ;
	assign x_2090 = (x_2085 & x_2089) ;
	assign x_2082 = (x_2078 & x_2081) ;
	assign x_2074 = (x_2069 & x_2073) ;
	assign x_2066 = (x_2062 & x_2065) ;
	assign x_2055 = (x_2050 & x_2054) ;
	assign x_2047 = (x_2042 & x_2046) ;
	assign x_2038 = (x_2033 & x_2037) ;
	assign x_2030 = (x_2026 & x_2029) ;
	assign x_2021 = (x_2016 & x_2020) ;
	assign x_2013 = (x_2009 & x_2012) ;
	assign x_2005 = (x_2000 & x_2004) ;
	assign x_1997 = (x_1993 & x_1996) ;
	assign x_1987 = (x_1982 & x_1986) ;
	assign x_1979 = (x_1975 & x_1978) ;
	assign x_1971 = (x_1966 & x_1970) ;
	assign x_1963 = (x_1959 & x_1962) ;
	assign x_1954 = (x_1949 & x_1953) ;
	assign x_1946 = (x_1942 & x_1945) ;
	assign x_1938 = (x_1933 & x_1937) ;
	assign x_1930 = (x_1926 & x_1929) ;
	assign x_1918 = (x_1913 & x_1917) ;
	assign x_1910 = (x_1905 & x_1909) ;
	assign x_1901 = (x_1896 & x_1900) ;
	assign x_1893 = (x_1889 & x_1892) ;
	assign x_1884 = (x_1879 & x_1883) ;
	assign x_1876 = (x_1872 & x_1875) ;
	assign x_1868 = (x_1863 & x_1867) ;
	assign x_1860 = (x_1856 & x_1859) ;
	assign x_1850 = (x_1845 & x_1849) ;
	assign x_1842 = (x_1837 & x_1841) ;
	assign x_1833 = (x_1828 & x_1832) ;
	assign x_1825 = (x_1821 & x_1824) ;
	assign x_1816 = (x_1811 & x_1815) ;
	assign x_1808 = (x_1804 & x_1807) ;
	assign x_1800 = (x_1795 & x_1799) ;
	assign x_1792 = (x_1788 & x_1791) ;
	assign x_1781 = (x_1776 & x_1780) ;
	assign x_1773 = (x_1768 & x_1772) ;
	assign x_1764 = (x_1759 & x_1763) ;
	assign x_1756 = (x_1752 & x_1755) ;
	assign x_1747 = (x_1742 & x_1746) ;
	assign x_1739 = (x_1735 & x_1738) ;
	assign x_1731 = (x_1726 & x_1730) ;
	assign x_1723 = (x_1719 & x_1722) ;
	assign x_1713 = (x_1708 & x_1712) ;
	assign x_1705 = (x_1701 & x_1704) ;
	assign x_1697 = (x_1692 & x_1696) ;
	assign x_1689 = (x_1685 & x_1688) ;
	assign x_1680 = (x_1675 & x_1679) ;
	assign x_1672 = (x_1668 & x_1671) ;
	assign x_1664 = (x_1659 & x_1663) ;
	assign x_1656 = (x_1652 & x_1655) ;
	assign x_1643 = (x_1638 & x_1642) ;
	assign x_1635 = (x_1630 & x_1634) ;
	assign x_1626 = (x_1621 & x_1625) ;
	assign x_1618 = (x_1614 & x_1617) ;
	assign x_1609 = (x_1604 & x_1608) ;
	assign x_1601 = (x_1597 & x_1600) ;
	assign x_1593 = (x_1588 & x_1592) ;
	assign x_1585 = (x_1581 & x_1584) ;
	assign x_1575 = (x_1570 & x_1574) ;
	assign x_1567 = (x_1562 & x_1566) ;
	assign x_1558 = (x_1553 & x_1557) ;
	assign x_1550 = (x_1546 & x_1549) ;
	assign x_1541 = (x_1536 & x_1540) ;
	assign x_1533 = (x_1529 & x_1532) ;
	assign x_1525 = (x_1520 & x_1524) ;
	assign x_1517 = (x_1513 & x_1516) ;
	assign x_1506 = (x_1501 & x_1505) ;
	assign x_1498 = (x_1493 & x_1497) ;
	assign x_1489 = (x_1484 & x_1488) ;
	assign x_1481 = (x_1477 & x_1480) ;
	assign x_1472 = (x_1467 & x_1471) ;
	assign x_1464 = (x_1460 & x_1463) ;
	assign x_1456 = (x_1451 & x_1455) ;
	assign x_1448 = (x_1444 & x_1447) ;
	assign x_1438 = (x_1433 & x_1437) ;
	assign x_1430 = (x_1426 & x_1429) ;
	assign x_1422 = (x_1417 & x_1421) ;
	assign x_1414 = (x_1410 & x_1413) ;
	assign x_1405 = (x_1400 & x_1404) ;
	assign x_1397 = (x_1393 & x_1396) ;
	assign x_1389 = (x_1384 & x_1388) ;
	assign x_1381 = (x_1377 & x_1380) ;
	assign x_1369 = (x_1364 & x_1368) ;
	assign x_1361 = (x_1356 & x_1360) ;
	assign x_1352 = (x_1347 & x_1351) ;
	assign x_1344 = (x_1340 & x_1343) ;
	assign x_1335 = (x_1330 & x_1334) ;
	assign x_1327 = (x_1323 & x_1326) ;
	assign x_1319 = (x_1314 & x_1318) ;
	assign x_1311 = (x_1307 & x_1310) ;
	assign x_1301 = (x_1296 & x_1300) ;
	assign x_1293 = (x_1288 & x_1292) ;
	assign x_1284 = (x_1279 & x_1283) ;
	assign x_1276 = (x_1272 & x_1275) ;
	assign x_1267 = (x_1262 & x_1266) ;
	assign x_1259 = (x_1255 & x_1258) ;
	assign x_1251 = (x_1246 & x_1250) ;
	assign x_1243 = (x_1239 & x_1242) ;
	assign x_1232 = (x_1227 & x_1231) ;
	assign x_1224 = (x_1219 & x_1223) ;
	assign x_1215 = (x_1210 & x_1214) ;
	assign x_1207 = (x_1203 & x_1206) ;
	assign x_1198 = (x_1193 & x_1197) ;
	assign x_1190 = (x_1186 & x_1189) ;
	assign x_1182 = (x_1177 & x_1181) ;
	assign x_1174 = (x_1170 & x_1173) ;
	assign x_1164 = (x_1159 & x_1163) ;
	assign x_1156 = (x_1152 & x_1155) ;
	assign x_1148 = (x_1143 & x_1147) ;
	assign x_1140 = (x_1136 & x_1139) ;
	assign x_1131 = (x_1126 & x_1130) ;
	assign x_1123 = (x_1119 & x_1122) ;
	assign x_1115 = (x_1110 & x_1114) ;
	assign x_1107 = (x_1103 & x_1106) ;
	assign x_2193 = (x_2184 & x_2192) ;
	assign x_2176 = (x_2167 & x_2175) ;
	assign x_2159 = (x_2150 & x_2158) ;
	assign x_2143 = (x_2134 & x_2142) ;
	assign x_2125 = (x_2116 & x_2124) ;
	assign x_2108 = (x_2099 & x_2107) ;
	assign x_2091 = (x_2082 & x_2090) ;
	assign x_2075 = (x_2066 & x_2074) ;
	assign x_2056 = (x_2047 & x_2055) ;
	assign x_2039 = (x_2030 & x_2038) ;
	assign x_2022 = (x_2013 & x_2021) ;
	assign x_2006 = (x_1997 & x_2005) ;
	assign x_1988 = (x_1979 & x_1987) ;
	assign x_1972 = (x_1963 & x_1971) ;
	assign x_1955 = (x_1946 & x_1954) ;
	assign x_1939 = (x_1930 & x_1938) ;
	assign x_1919 = (x_1910 & x_1918) ;
	assign x_1902 = (x_1893 & x_1901) ;
	assign x_1885 = (x_1876 & x_1884) ;
	assign x_1869 = (x_1860 & x_1868) ;
	assign x_1851 = (x_1842 & x_1850) ;
	assign x_1834 = (x_1825 & x_1833) ;
	assign x_1817 = (x_1808 & x_1816) ;
	assign x_1801 = (x_1792 & x_1800) ;
	assign x_1782 = (x_1773 & x_1781) ;
	assign x_1765 = (x_1756 & x_1764) ;
	assign x_1748 = (x_1739 & x_1747) ;
	assign x_1732 = (x_1723 & x_1731) ;
	assign x_1714 = (x_1705 & x_1713) ;
	assign x_1698 = (x_1689 & x_1697) ;
	assign x_1681 = (x_1672 & x_1680) ;
	assign x_1665 = (x_1656 & x_1664) ;
	assign x_1644 = (x_1635 & x_1643) ;
	assign x_1627 = (x_1618 & x_1626) ;
	assign x_1610 = (x_1601 & x_1609) ;
	assign x_1594 = (x_1585 & x_1593) ;
	assign x_1576 = (x_1567 & x_1575) ;
	assign x_1559 = (x_1550 & x_1558) ;
	assign x_1542 = (x_1533 & x_1541) ;
	assign x_1526 = (x_1517 & x_1525) ;
	assign x_1507 = (x_1498 & x_1506) ;
	assign x_1490 = (x_1481 & x_1489) ;
	assign x_1473 = (x_1464 & x_1472) ;
	assign x_1457 = (x_1448 & x_1456) ;
	assign x_1439 = (x_1430 & x_1438) ;
	assign x_1423 = (x_1414 & x_1422) ;
	assign x_1406 = (x_1397 & x_1405) ;
	assign x_1390 = (x_1381 & x_1389) ;
	assign x_1370 = (x_1361 & x_1369) ;
	assign x_1353 = (x_1344 & x_1352) ;
	assign x_1336 = (x_1327 & x_1335) ;
	assign x_1320 = (x_1311 & x_1319) ;
	assign x_1302 = (x_1293 & x_1301) ;
	assign x_1285 = (x_1276 & x_1284) ;
	assign x_1268 = (x_1259 & x_1267) ;
	assign x_1252 = (x_1243 & x_1251) ;
	assign x_1233 = (x_1224 & x_1232) ;
	assign x_1216 = (x_1207 & x_1215) ;
	assign x_1199 = (x_1190 & x_1198) ;
	assign x_1183 = (x_1174 & x_1182) ;
	assign x_1165 = (x_1156 & x_1164) ;
	assign x_1149 = (x_1140 & x_1148) ;
	assign x_1132 = (x_1123 & x_1131) ;
	assign x_1116 = (x_1107 & x_1115) ;
	assign x_2194 = (x_2176 & x_2193) ;
	assign x_2160 = (x_2143 & x_2159) ;
	assign x_2126 = (x_2108 & x_2125) ;
	assign x_2092 = (x_2075 & x_2091) ;
	assign x_2057 = (x_2039 & x_2056) ;
	assign x_2023 = (x_2006 & x_2022) ;
	assign x_1989 = (x_1972 & x_1988) ;
	assign x_1956 = (x_1939 & x_1955) ;
	assign x_1920 = (x_1902 & x_1919) ;
	assign x_1886 = (x_1869 & x_1885) ;
	assign x_1852 = (x_1834 & x_1851) ;
	assign x_1818 = (x_1801 & x_1817) ;
	assign x_1783 = (x_1765 & x_1782) ;
	assign x_1749 = (x_1732 & x_1748) ;
	assign x_1715 = (x_1698 & x_1714) ;
	assign x_1682 = (x_1665 & x_1681) ;
	assign x_1645 = (x_1627 & x_1644) ;
	assign x_1611 = (x_1594 & x_1610) ;
	assign x_1577 = (x_1559 & x_1576) ;
	assign x_1543 = (x_1526 & x_1542) ;
	assign x_1508 = (x_1490 & x_1507) ;
	assign x_1474 = (x_1457 & x_1473) ;
	assign x_1440 = (x_1423 & x_1439) ;
	assign x_1407 = (x_1390 & x_1406) ;
	assign x_1371 = (x_1353 & x_1370) ;
	assign x_1337 = (x_1320 & x_1336) ;
	assign x_1303 = (x_1285 & x_1302) ;
	assign x_1269 = (x_1252 & x_1268) ;
	assign x_1234 = (x_1216 & x_1233) ;
	assign x_1200 = (x_1183 & x_1199) ;
	assign x_1166 = (x_1149 & x_1165) ;
	assign x_1133 = (x_1116 & x_1132) ;
	assign x_2195 = (x_2160 & x_2194) ;
	assign x_2127 = (x_2092 & x_2126) ;
	assign x_2058 = (x_2023 & x_2057) ;
	assign x_1990 = (x_1956 & x_1989) ;
	assign x_1921 = (x_1886 & x_1920) ;
	assign x_1853 = (x_1818 & x_1852) ;
	assign x_1784 = (x_1749 & x_1783) ;
	assign x_1716 = (x_1682 & x_1715) ;
	assign x_1646 = (x_1611 & x_1645) ;
	assign x_1578 = (x_1543 & x_1577) ;
	assign x_1509 = (x_1474 & x_1508) ;
	assign x_1441 = (x_1407 & x_1440) ;
	assign x_1372 = (x_1337 & x_1371) ;
	assign x_1304 = (x_1269 & x_1303) ;
	assign x_1235 = (x_1200 & x_1234) ;
	assign x_1167 = (x_1133 & x_1166) ;
	assign x_2196 = (x_2127 & x_2195) ;
	assign x_2059 = (x_1990 & x_2058) ;
	assign x_1922 = (x_1853 & x_1921) ;
	assign x_1785 = (x_1716 & x_1784) ;
	assign x_1647 = (x_1578 & x_1646) ;
	assign x_1510 = (x_1441 & x_1509) ;
	assign x_1373 = (x_1304 & x_1372) ;
	assign x_1236 = (x_1167 & x_1235) ;
	assign x_2197 = (x_2059 & x_2196) ;
	assign x_1923 = (x_1785 & x_1922) ;
	assign x_1648 = (x_1510 & x_1647) ;
	assign x_1374 = (x_1236 & x_1373) ;
	assign x_2198 = (x_1923 & x_2197) ;
	assign x_1649 = (x_1374 & x_1648) ;
	assign x_2199 = (x_1649 & x_2198) ;
	assign o_1 = x_2199 ;
endmodule
