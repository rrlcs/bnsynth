// skolem function for order file variables
// Generated using findDep.cpp 
module formula (v_2, v_3, v_8, v_9, v_10, v_11, v_12, v_73, v_74, v_75, v_76, v_77, v_138, v_139, v_140, v_141, v_142, v_203, v_204, v_209, v_210, v_215, v_216, v_221, v_222, v_227, v_228, v_233, v_234, v_239, v_240, v_245, v_246, v_251, v_252, v_257, v_258, v_263, v_264, v_269, v_270, v_271, v_272, v_273, v_334, v_335, v_336, v_337, v_338, v_399, v_400, v_405, v_406, v_411, v_412, v_417, v_418, v_423, v_424, v_429, v_430, v_435, v_436, v_441, v_442, v_447, v_448, v_453, v_454, v_459, v_460, v_461, v_462, v_463, v_464, v_466, v_467, v_468, v_469, v_470, v_471, v_472, v_473, v_474, v_475, v_476, v_477, v_478, v_479, v_480, v_481, v_482, v_483, v_484, v_485, v_516, v_523, v_525, v_526, v_527, v_528, v_529, v_530, v_531, v_532, v_549, v_564, v_566, v_611, v_612, v_620, v_649, v_657, v_696, v_702, v_730, v_731, v_739, v_760, v_768, v_798, v_799, v_807, v_828, v_836, v_866, v_867, v_875, v_896, v_904, v_912, v_913, v_915, v_919, v_922, v_923, v_925, v_929, v_930, v_931, v_960, v_962, v_968, v_971, v_972, v_992, v_994, v_1007, v_1009, v_1032, v_1039, v_1042, v_1043, v_1044, v_1047, v_1048, v_1049, v_1050, v_1067, v_1069, v_1083, v_1085, v_1087, v_1101, v_1103, v_1105, v_1107, v_1119, v_1122, v_1125, v_1153, v_1154, v_1162, v_1183, v_1191, v_1221, v_1222, v_1230, v_1251, v_1259, v_1289, v_1290, v_1298, v_1319, v_1327, v_1357, v_1358, v_1366, v_1387, v_1395, v_1403, v_1404, v_1407, v_1408, v_1409, v_1411, v_1418, v_1421, v_1422, v_1424, v_1428, v_1429, v_1430, v_1432, v_1437, v_1438, v_1439, v_1440, v_1513, v_1526, v_1529, v_1530, v_1532, v_1536, v_1537, v_1538, v_1603, v_1605, v_1617, v_1620, v_1621, v_1677, v_1679, v_1726, v_1728, v_1745, v_1746, v_1747, v_1749, v_1750, v_1751, v_1752, v_1770, v_1772, v_1786, v_1788, v_1790, v_1804, v_1806, v_1808, v_1810, v_1848, v_1849, v_1857, v_1878, v_1886, v_1916, v_1917, v_1925, v_1946, v_1954, v_1984, v_1985, v_1993, v_2014, v_2022, v_2052, v_2053, v_2061, v_2082, v_2090, v_2098, v_2099, v_2102, v_2103, v_2104, v_2106, v_2110, v_2113, v_2114, v_2116, v_2120, v_2121, v_2122, v_2124, v_2129, v_2130, v_2131, v_2132, v_2169, v_2171, v_2177, v_2180, v_2181, v_2183, v_2187, v_2188, v_2189, v_2217, v_2219, v_2225, v_2228, v_2229, v_2248, v_2250, v_2263, v_2265, v_2280, v_2334, v_2336, v_2362, v_2364, v_2366, v_2392, v_2394, v_2396, v_2398, v_2452, v_2453, v_2462, v_2493, v_2502, v_2530, v_2531, v_2532, v_2533, v_2543, v_2564, v_2574, v_2604, v_2605, v_2606, v_2607, v_2617, v_2638, v_2648, v_2678, v_2679, v_2680, v_2681, v_2691, v_2712, v_2722, v_2752, v_2753, v_2754, v_2755, v_2765, v_2786, v_2796, v_2804, v_2805, v_2808, v_2809, v_2810, v_2812, v_2816, v_2819, v_2820, v_2822, v_2826, v_2827, v_2828, v_2830, v_2835, v_2836, v_2837, v_2838, v_2875, v_2877, v_2882, v_2885, v_2886, v_2888, v_2892, v_2893, v_2894, v_2922, v_2924, v_2929, v_2932, v_2933, v_2952, v_2954, v_2967, v_2969, v_2988, v_3013, v_3028, v_3030, v_3044, v_3047, v_3050, v_3052, v_3080, v_3088, v_3109, v_3117, v_3147, v_3155, v_3176, v_3184, v_3214, v_3222, v_3243, v_3251, v_3259, v_3260, o_1);
input v_2;
input v_3;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_73;
input v_74;
input v_75;
input v_76;
input v_77;
input v_138;
input v_139;
input v_140;
input v_141;
input v_142;
input v_203;
input v_204;
input v_209;
input v_210;
input v_215;
input v_216;
input v_221;
input v_222;
input v_227;
input v_228;
input v_233;
input v_234;
input v_239;
input v_240;
input v_245;
input v_246;
input v_251;
input v_252;
input v_257;
input v_258;
input v_263;
input v_264;
input v_269;
input v_270;
input v_271;
input v_272;
input v_273;
input v_334;
input v_335;
input v_336;
input v_337;
input v_338;
input v_399;
input v_400;
input v_405;
input v_406;
input v_411;
input v_412;
input v_417;
input v_418;
input v_423;
input v_424;
input v_429;
input v_430;
input v_435;
input v_436;
input v_441;
input v_442;
input v_447;
input v_448;
input v_453;
input v_454;
input v_459;
input v_460;
input v_461;
input v_462;
input v_463;
input v_464;
input v_466;
input v_467;
input v_468;
input v_469;
input v_470;
input v_471;
input v_472;
input v_473;
input v_474;
input v_475;
input v_476;
input v_477;
input v_478;
input v_479;
input v_480;
input v_481;
input v_482;
input v_483;
input v_484;
input v_485;
input v_516;
input v_523;
input v_525;
input v_526;
input v_527;
input v_528;
input v_529;
input v_530;
input v_531;
input v_532;
input v_549;
input v_564;
input v_566;
input v_611;
input v_612;
input v_620;
input v_649;
input v_657;
input v_696;
input v_702;
input v_730;
input v_731;
input v_739;
input v_760;
input v_768;
input v_798;
input v_799;
input v_807;
input v_828;
input v_836;
input v_866;
input v_867;
input v_875;
input v_896;
input v_904;
input v_912;
input v_913;
input v_915;
input v_919;
input v_922;
input v_923;
input v_925;
input v_929;
input v_930;
input v_931;
input v_960;
input v_962;
input v_968;
input v_971;
input v_972;
input v_992;
input v_994;
input v_1007;
input v_1009;
input v_1032;
input v_1039;
input v_1042;
input v_1043;
input v_1044;
input v_1047;
input v_1048;
input v_1049;
input v_1050;
input v_1067;
input v_1069;
input v_1083;
input v_1085;
input v_1087;
input v_1101;
input v_1103;
input v_1105;
input v_1107;
input v_1119;
input v_1122;
input v_1125;
input v_1153;
input v_1154;
input v_1162;
input v_1183;
input v_1191;
input v_1221;
input v_1222;
input v_1230;
input v_1251;
input v_1259;
input v_1289;
input v_1290;
input v_1298;
input v_1319;
input v_1327;
input v_1357;
input v_1358;
input v_1366;
input v_1387;
input v_1395;
input v_1403;
input v_1404;
input v_1407;
input v_1408;
input v_1409;
input v_1411;
input v_1418;
input v_1421;
input v_1422;
input v_1424;
input v_1428;
input v_1429;
input v_1430;
input v_1432;
input v_1437;
input v_1438;
input v_1439;
input v_1440;
input v_1513;
input v_1526;
input v_1529;
input v_1530;
input v_1532;
input v_1536;
input v_1537;
input v_1538;
input v_1603;
input v_1605;
input v_1617;
input v_1620;
input v_1621;
input v_1677;
input v_1679;
input v_1726;
input v_1728;
input v_1745;
input v_1746;
input v_1747;
input v_1749;
input v_1750;
input v_1751;
input v_1752;
input v_1770;
input v_1772;
input v_1786;
input v_1788;
input v_1790;
input v_1804;
input v_1806;
input v_1808;
input v_1810;
input v_1848;
input v_1849;
input v_1857;
input v_1878;
input v_1886;
input v_1916;
input v_1917;
input v_1925;
input v_1946;
input v_1954;
input v_1984;
input v_1985;
input v_1993;
input v_2014;
input v_2022;
input v_2052;
input v_2053;
input v_2061;
input v_2082;
input v_2090;
input v_2098;
input v_2099;
input v_2102;
input v_2103;
input v_2104;
input v_2106;
input v_2110;
input v_2113;
input v_2114;
input v_2116;
input v_2120;
input v_2121;
input v_2122;
input v_2124;
input v_2129;
input v_2130;
input v_2131;
input v_2132;
input v_2169;
input v_2171;
input v_2177;
input v_2180;
input v_2181;
input v_2183;
input v_2187;
input v_2188;
input v_2189;
input v_2217;
input v_2219;
input v_2225;
input v_2228;
input v_2229;
input v_2248;
input v_2250;
input v_2263;
input v_2265;
input v_2280;
input v_2334;
input v_2336;
input v_2362;
input v_2364;
input v_2366;
input v_2392;
input v_2394;
input v_2396;
input v_2398;
input v_2452;
input v_2453;
input v_2462;
input v_2493;
input v_2502;
input v_2530;
input v_2531;
input v_2532;
input v_2533;
input v_2543;
input v_2564;
input v_2574;
input v_2604;
input v_2605;
input v_2606;
input v_2607;
input v_2617;
input v_2638;
input v_2648;
input v_2678;
input v_2679;
input v_2680;
input v_2681;
input v_2691;
input v_2712;
input v_2722;
input v_2752;
input v_2753;
input v_2754;
input v_2755;
input v_2765;
input v_2786;
input v_2796;
input v_2804;
input v_2805;
input v_2808;
input v_2809;
input v_2810;
input v_2812;
input v_2816;
input v_2819;
input v_2820;
input v_2822;
input v_2826;
input v_2827;
input v_2828;
input v_2830;
input v_2835;
input v_2836;
input v_2837;
input v_2838;
input v_2875;
input v_2877;
input v_2882;
input v_2885;
input v_2886;
input v_2888;
input v_2892;
input v_2893;
input v_2894;
input v_2922;
input v_2924;
input v_2929;
input v_2932;
input v_2933;
input v_2952;
input v_2954;
input v_2967;
input v_2969;
input v_2988;
input v_3013;
input v_3028;
input v_3030;
input v_3044;
input v_3047;
input v_3050;
input v_3052;
input v_3080;
input v_3088;
input v_3109;
input v_3117;
input v_3147;
input v_3155;
input v_3176;
input v_3184;
input v_3214;
input v_3222;
input v_3243;
input v_3251;
input v_3259;
input v_3260;
output o_1;
wire v_4;
wire v_5;
wire v_6;
wire v_7;
wire v_13;
wire v_14;
wire v_15;
wire v_16;
wire v_17;
wire v_18;
wire v_19;
wire v_20;
wire v_21;
wire v_22;
wire v_23;
wire v_24;
wire v_25;
wire v_26;
wire v_27;
wire v_28;
wire v_29;
wire v_30;
wire v_31;
wire v_32;
wire v_33;
wire v_34;
wire v_35;
wire v_36;
wire v_37;
wire v_38;
wire v_39;
wire v_40;
wire v_41;
wire v_42;
wire v_43;
wire v_44;
wire v_45;
wire v_46;
wire v_47;
wire v_48;
wire v_49;
wire v_50;
wire v_51;
wire v_52;
wire v_53;
wire v_54;
wire v_55;
wire v_56;
wire v_57;
wire v_58;
wire v_59;
wire v_60;
wire v_61;
wire v_62;
wire v_63;
wire v_64;
wire v_65;
wire v_66;
wire v_67;
wire v_68;
wire v_69;
wire v_70;
wire v_71;
wire v_72;
wire v_78;
wire v_79;
wire v_80;
wire v_81;
wire v_82;
wire v_83;
wire v_84;
wire v_85;
wire v_86;
wire v_87;
wire v_88;
wire v_89;
wire v_90;
wire v_91;
wire v_92;
wire v_93;
wire v_94;
wire v_95;
wire v_96;
wire v_97;
wire v_98;
wire v_99;
wire v_100;
wire v_101;
wire v_102;
wire v_103;
wire v_104;
wire v_105;
wire v_106;
wire v_107;
wire v_108;
wire v_109;
wire v_110;
wire v_111;
wire v_112;
wire v_113;
wire v_114;
wire v_115;
wire v_116;
wire v_117;
wire v_118;
wire v_119;
wire v_120;
wire v_121;
wire v_122;
wire v_123;
wire v_124;
wire v_125;
wire v_126;
wire v_127;
wire v_128;
wire v_129;
wire v_130;
wire v_131;
wire v_132;
wire v_133;
wire v_134;
wire v_135;
wire v_136;
wire v_137;
wire v_143;
wire v_144;
wire v_145;
wire v_146;
wire v_147;
wire v_148;
wire v_149;
wire v_150;
wire v_151;
wire v_152;
wire v_153;
wire v_154;
wire v_155;
wire v_156;
wire v_157;
wire v_158;
wire v_159;
wire v_160;
wire v_161;
wire v_162;
wire v_163;
wire v_164;
wire v_165;
wire v_166;
wire v_167;
wire v_168;
wire v_169;
wire v_170;
wire v_171;
wire v_172;
wire v_173;
wire v_174;
wire v_175;
wire v_176;
wire v_177;
wire v_178;
wire v_179;
wire v_180;
wire v_181;
wire v_182;
wire v_183;
wire v_184;
wire v_185;
wire v_186;
wire v_187;
wire v_188;
wire v_189;
wire v_190;
wire v_191;
wire v_192;
wire v_193;
wire v_194;
wire v_195;
wire v_196;
wire v_197;
wire v_198;
wire v_199;
wire v_200;
wire v_201;
wire v_202;
wire v_205;
wire v_206;
wire v_207;
wire v_208;
wire v_211;
wire v_212;
wire v_213;
wire v_214;
wire v_217;
wire v_218;
wire v_219;
wire v_220;
wire v_223;
wire v_224;
wire v_225;
wire v_226;
wire v_229;
wire v_230;
wire v_231;
wire v_232;
wire v_235;
wire v_236;
wire v_237;
wire v_238;
wire v_241;
wire v_242;
wire v_243;
wire v_244;
wire v_247;
wire v_248;
wire v_249;
wire v_250;
wire v_253;
wire v_254;
wire v_255;
wire v_256;
wire v_259;
wire v_260;
wire v_261;
wire v_262;
wire v_265;
wire v_266;
wire v_267;
wire v_268;
wire v_274;
wire v_275;
wire v_276;
wire v_277;
wire v_278;
wire v_279;
wire v_280;
wire v_281;
wire v_282;
wire v_283;
wire v_284;
wire v_285;
wire v_286;
wire v_287;
wire v_288;
wire v_289;
wire v_290;
wire v_291;
wire v_292;
wire v_293;
wire v_294;
wire v_295;
wire v_296;
wire v_297;
wire v_298;
wire v_299;
wire v_300;
wire v_301;
wire v_302;
wire v_303;
wire v_304;
wire v_305;
wire v_306;
wire v_307;
wire v_308;
wire v_309;
wire v_310;
wire v_311;
wire v_312;
wire v_313;
wire v_314;
wire v_315;
wire v_316;
wire v_317;
wire v_318;
wire v_319;
wire v_320;
wire v_321;
wire v_322;
wire v_323;
wire v_324;
wire v_325;
wire v_326;
wire v_327;
wire v_328;
wire v_329;
wire v_330;
wire v_331;
wire v_332;
wire v_333;
wire v_339;
wire v_340;
wire v_341;
wire v_342;
wire v_343;
wire v_344;
wire v_345;
wire v_346;
wire v_347;
wire v_348;
wire v_349;
wire v_350;
wire v_351;
wire v_352;
wire v_353;
wire v_354;
wire v_355;
wire v_356;
wire v_357;
wire v_358;
wire v_359;
wire v_360;
wire v_361;
wire v_362;
wire v_363;
wire v_364;
wire v_365;
wire v_366;
wire v_367;
wire v_368;
wire v_369;
wire v_370;
wire v_371;
wire v_372;
wire v_373;
wire v_374;
wire v_375;
wire v_376;
wire v_377;
wire v_378;
wire v_379;
wire v_380;
wire v_381;
wire v_382;
wire v_383;
wire v_384;
wire v_385;
wire v_386;
wire v_387;
wire v_388;
wire v_389;
wire v_390;
wire v_391;
wire v_392;
wire v_393;
wire v_394;
wire v_395;
wire v_396;
wire v_397;
wire v_398;
wire v_401;
wire v_402;
wire v_403;
wire v_404;
wire v_407;
wire v_408;
wire v_409;
wire v_410;
wire v_413;
wire v_414;
wire v_415;
wire v_416;
wire v_419;
wire v_420;
wire v_421;
wire v_422;
wire v_425;
wire v_426;
wire v_427;
wire v_428;
wire v_431;
wire v_432;
wire v_433;
wire v_434;
wire v_437;
wire v_438;
wire v_439;
wire v_440;
wire v_443;
wire v_444;
wire v_445;
wire v_446;
wire v_449;
wire v_450;
wire v_451;
wire v_452;
wire v_455;
wire v_456;
wire v_457;
wire v_458;
wire v_486;
wire v_487;
wire v_488;
wire v_489;
wire v_490;
wire v_491;
wire v_492;
wire v_493;
wire v_494;
wire v_495;
wire v_496;
wire v_497;
wire v_498;
wire v_499;
wire v_500;
wire v_501;
wire v_502;
wire v_503;
wire v_504;
wire v_505;
wire v_506;
wire v_507;
wire v_508;
wire v_509;
wire v_510;
wire v_511;
wire v_512;
wire v_513;
wire v_514;
wire v_515;
wire v_517;
wire v_518;
wire v_519;
wire v_520;
wire v_521;
wire v_522;
wire v_524;
wire v_533;
wire v_534;
wire v_535;
wire v_536;
wire v_537;
wire v_538;
wire v_539;
wire v_540;
wire v_541;
wire v_542;
wire v_543;
wire v_544;
wire v_545;
wire v_546;
wire v_547;
wire v_548;
wire v_550;
wire v_551;
wire v_552;
wire v_553;
wire v_554;
wire v_555;
wire v_556;
wire v_557;
wire v_558;
wire v_559;
wire v_560;
wire v_561;
wire v_562;
wire v_563;
wire v_565;
wire v_567;
wire v_568;
wire v_569;
wire v_570;
wire v_571;
wire v_572;
wire v_573;
wire v_574;
wire v_575;
wire v_576;
wire v_577;
wire v_578;
wire v_579;
wire v_580;
wire v_581;
wire v_582;
wire v_583;
wire v_584;
wire v_585;
wire v_586;
wire v_587;
wire v_588;
wire v_589;
wire v_590;
wire v_591;
wire v_592;
wire v_593;
wire v_594;
wire v_595;
wire v_596;
wire v_597;
wire v_598;
wire v_599;
wire v_600;
wire v_601;
wire v_602;
wire v_603;
wire v_604;
wire v_605;
wire v_606;
wire v_607;
wire v_608;
wire v_609;
wire v_610;
wire v_613;
wire v_614;
wire v_615;
wire v_616;
wire v_617;
wire v_618;
wire v_619;
wire v_621;
wire v_622;
wire v_623;
wire v_624;
wire v_625;
wire v_626;
wire v_627;
wire v_628;
wire v_629;
wire v_630;
wire v_631;
wire v_632;
wire v_633;
wire v_634;
wire v_635;
wire v_636;
wire v_637;
wire v_638;
wire v_639;
wire v_640;
wire v_641;
wire v_642;
wire v_643;
wire v_644;
wire v_645;
wire v_646;
wire v_647;
wire v_648;
wire v_650;
wire v_651;
wire v_652;
wire v_653;
wire v_654;
wire v_655;
wire v_656;
wire v_658;
wire v_659;
wire v_660;
wire v_661;
wire v_662;
wire v_663;
wire v_664;
wire v_665;
wire v_666;
wire v_667;
wire v_668;
wire v_669;
wire v_670;
wire v_671;
wire v_672;
wire v_673;
wire v_674;
wire v_675;
wire v_676;
wire v_677;
wire v_678;
wire v_679;
wire v_680;
wire v_681;
wire v_682;
wire v_683;
wire v_684;
wire v_685;
wire v_686;
wire v_687;
wire v_688;
wire v_689;
wire v_690;
wire v_691;
wire v_692;
wire v_693;
wire v_694;
wire v_695;
wire v_697;
wire v_698;
wire v_699;
wire v_700;
wire v_701;
wire v_703;
wire v_704;
wire v_705;
wire v_706;
wire v_707;
wire v_708;
wire v_709;
wire v_710;
wire v_711;
wire v_712;
wire v_713;
wire v_714;
wire v_715;
wire v_716;
wire v_717;
wire v_718;
wire v_719;
wire v_720;
wire v_721;
wire v_722;
wire v_723;
wire v_724;
wire v_725;
wire v_726;
wire v_727;
wire v_728;
wire v_729;
wire v_732;
wire v_733;
wire v_734;
wire v_735;
wire v_736;
wire v_737;
wire v_738;
wire v_740;
wire v_741;
wire v_742;
wire v_743;
wire v_744;
wire v_745;
wire v_746;
wire v_747;
wire v_748;
wire v_749;
wire v_750;
wire v_751;
wire v_752;
wire v_753;
wire v_754;
wire v_755;
wire v_756;
wire v_757;
wire v_758;
wire v_759;
wire v_761;
wire v_762;
wire v_763;
wire v_764;
wire v_765;
wire v_766;
wire v_767;
wire v_769;
wire v_770;
wire v_771;
wire v_772;
wire v_773;
wire v_774;
wire v_775;
wire v_776;
wire v_777;
wire v_778;
wire v_779;
wire v_780;
wire v_781;
wire v_782;
wire v_783;
wire v_784;
wire v_785;
wire v_786;
wire v_787;
wire v_788;
wire v_789;
wire v_790;
wire v_791;
wire v_792;
wire v_793;
wire v_794;
wire v_795;
wire v_796;
wire v_797;
wire v_800;
wire v_801;
wire v_802;
wire v_803;
wire v_804;
wire v_805;
wire v_806;
wire v_808;
wire v_809;
wire v_810;
wire v_811;
wire v_812;
wire v_813;
wire v_814;
wire v_815;
wire v_816;
wire v_817;
wire v_818;
wire v_819;
wire v_820;
wire v_821;
wire v_822;
wire v_823;
wire v_824;
wire v_825;
wire v_826;
wire v_827;
wire v_829;
wire v_830;
wire v_831;
wire v_832;
wire v_833;
wire v_834;
wire v_835;
wire v_837;
wire v_838;
wire v_839;
wire v_840;
wire v_841;
wire v_842;
wire v_843;
wire v_844;
wire v_845;
wire v_846;
wire v_847;
wire v_848;
wire v_849;
wire v_850;
wire v_851;
wire v_852;
wire v_853;
wire v_854;
wire v_855;
wire v_856;
wire v_857;
wire v_858;
wire v_859;
wire v_860;
wire v_861;
wire v_862;
wire v_863;
wire v_864;
wire v_865;
wire v_868;
wire v_869;
wire v_870;
wire v_871;
wire v_872;
wire v_873;
wire v_874;
wire v_876;
wire v_877;
wire v_878;
wire v_879;
wire v_880;
wire v_881;
wire v_882;
wire v_883;
wire v_884;
wire v_885;
wire v_886;
wire v_887;
wire v_888;
wire v_889;
wire v_890;
wire v_891;
wire v_892;
wire v_893;
wire v_894;
wire v_895;
wire v_897;
wire v_898;
wire v_899;
wire v_900;
wire v_901;
wire v_902;
wire v_903;
wire v_905;
wire v_906;
wire v_907;
wire v_908;
wire v_909;
wire v_910;
wire v_911;
wire v_914;
wire v_916;
wire v_917;
wire v_918;
wire v_920;
wire v_921;
wire v_924;
wire v_926;
wire v_927;
wire v_928;
wire v_932;
wire v_933;
wire v_934;
wire v_935;
wire v_936;
wire v_937;
wire v_938;
wire v_939;
wire v_940;
wire v_941;
wire v_942;
wire v_943;
wire v_944;
wire v_945;
wire v_946;
wire v_947;
wire v_948;
wire v_949;
wire v_950;
wire v_951;
wire v_952;
wire v_953;
wire v_954;
wire v_955;
wire v_956;
wire v_957;
wire v_958;
wire v_959;
wire v_961;
wire v_963;
wire v_964;
wire v_965;
wire v_966;
wire v_967;
wire v_969;
wire v_970;
wire v_973;
wire v_974;
wire v_975;
wire v_976;
wire v_977;
wire v_978;
wire v_979;
wire v_980;
wire v_981;
wire v_982;
wire v_983;
wire v_984;
wire v_985;
wire v_986;
wire v_987;
wire v_988;
wire v_989;
wire v_990;
wire v_991;
wire v_993;
wire v_995;
wire v_996;
wire v_997;
wire v_998;
wire v_999;
wire v_1000;
wire v_1001;
wire v_1002;
wire v_1003;
wire v_1004;
wire v_1005;
wire v_1006;
wire v_1008;
wire v_1010;
wire v_1011;
wire v_1012;
wire v_1013;
wire v_1014;
wire v_1015;
wire v_1016;
wire v_1017;
wire v_1018;
wire v_1019;
wire v_1020;
wire v_1021;
wire v_1022;
wire v_1023;
wire v_1024;
wire v_1025;
wire v_1026;
wire v_1027;
wire v_1028;
wire v_1029;
wire v_1030;
wire v_1031;
wire v_1033;
wire v_1034;
wire v_1035;
wire v_1036;
wire v_1037;
wire v_1038;
wire v_1040;
wire v_1041;
wire v_1045;
wire v_1046;
wire v_1051;
wire v_1052;
wire v_1053;
wire v_1054;
wire v_1055;
wire v_1056;
wire v_1057;
wire v_1058;
wire v_1059;
wire v_1060;
wire v_1061;
wire v_1062;
wire v_1063;
wire v_1064;
wire v_1065;
wire v_1066;
wire v_1068;
wire v_1070;
wire v_1071;
wire v_1072;
wire v_1073;
wire v_1074;
wire v_1075;
wire v_1076;
wire v_1077;
wire v_1078;
wire v_1079;
wire v_1080;
wire v_1081;
wire v_1082;
wire v_1084;
wire v_1086;
wire v_1088;
wire v_1089;
wire v_1090;
wire v_1091;
wire v_1092;
wire v_1093;
wire v_1094;
wire v_1095;
wire v_1096;
wire v_1097;
wire v_1098;
wire v_1099;
wire v_1100;
wire v_1102;
wire v_1104;
wire v_1106;
wire v_1108;
wire v_1109;
wire v_1110;
wire v_1111;
wire v_1112;
wire v_1113;
wire v_1114;
wire v_1115;
wire v_1116;
wire v_1117;
wire v_1118;
wire v_1120;
wire v_1121;
wire v_1123;
wire v_1124;
wire v_1126;
wire v_1127;
wire v_1128;
wire v_1129;
wire v_1130;
wire v_1131;
wire v_1132;
wire v_1133;
wire v_1134;
wire v_1135;
wire v_1136;
wire v_1137;
wire v_1138;
wire v_1139;
wire v_1140;
wire v_1141;
wire v_1142;
wire v_1143;
wire v_1144;
wire v_1145;
wire v_1146;
wire v_1147;
wire v_1148;
wire v_1149;
wire v_1150;
wire v_1151;
wire v_1152;
wire v_1155;
wire v_1156;
wire v_1157;
wire v_1158;
wire v_1159;
wire v_1160;
wire v_1161;
wire v_1163;
wire v_1164;
wire v_1165;
wire v_1166;
wire v_1167;
wire v_1168;
wire v_1169;
wire v_1170;
wire v_1171;
wire v_1172;
wire v_1173;
wire v_1174;
wire v_1175;
wire v_1176;
wire v_1177;
wire v_1178;
wire v_1179;
wire v_1180;
wire v_1181;
wire v_1182;
wire v_1184;
wire v_1185;
wire v_1186;
wire v_1187;
wire v_1188;
wire v_1189;
wire v_1190;
wire v_1192;
wire v_1193;
wire v_1194;
wire v_1195;
wire v_1196;
wire v_1197;
wire v_1198;
wire v_1199;
wire v_1200;
wire v_1201;
wire v_1202;
wire v_1203;
wire v_1204;
wire v_1205;
wire v_1206;
wire v_1207;
wire v_1208;
wire v_1209;
wire v_1210;
wire v_1211;
wire v_1212;
wire v_1213;
wire v_1214;
wire v_1215;
wire v_1216;
wire v_1217;
wire v_1218;
wire v_1219;
wire v_1220;
wire v_1223;
wire v_1224;
wire v_1225;
wire v_1226;
wire v_1227;
wire v_1228;
wire v_1229;
wire v_1231;
wire v_1232;
wire v_1233;
wire v_1234;
wire v_1235;
wire v_1236;
wire v_1237;
wire v_1238;
wire v_1239;
wire v_1240;
wire v_1241;
wire v_1242;
wire v_1243;
wire v_1244;
wire v_1245;
wire v_1246;
wire v_1247;
wire v_1248;
wire v_1249;
wire v_1250;
wire v_1252;
wire v_1253;
wire v_1254;
wire v_1255;
wire v_1256;
wire v_1257;
wire v_1258;
wire v_1260;
wire v_1261;
wire v_1262;
wire v_1263;
wire v_1264;
wire v_1265;
wire v_1266;
wire v_1267;
wire v_1268;
wire v_1269;
wire v_1270;
wire v_1271;
wire v_1272;
wire v_1273;
wire v_1274;
wire v_1275;
wire v_1276;
wire v_1277;
wire v_1278;
wire v_1279;
wire v_1280;
wire v_1281;
wire v_1282;
wire v_1283;
wire v_1284;
wire v_1285;
wire v_1286;
wire v_1287;
wire v_1288;
wire v_1291;
wire v_1292;
wire v_1293;
wire v_1294;
wire v_1295;
wire v_1296;
wire v_1297;
wire v_1299;
wire v_1300;
wire v_1301;
wire v_1302;
wire v_1303;
wire v_1304;
wire v_1305;
wire v_1306;
wire v_1307;
wire v_1308;
wire v_1309;
wire v_1310;
wire v_1311;
wire v_1312;
wire v_1313;
wire v_1314;
wire v_1315;
wire v_1316;
wire v_1317;
wire v_1318;
wire v_1320;
wire v_1321;
wire v_1322;
wire v_1323;
wire v_1324;
wire v_1325;
wire v_1326;
wire v_1328;
wire v_1329;
wire v_1330;
wire v_1331;
wire v_1332;
wire v_1333;
wire v_1334;
wire v_1335;
wire v_1336;
wire v_1337;
wire v_1338;
wire v_1339;
wire v_1340;
wire v_1341;
wire v_1342;
wire v_1343;
wire v_1344;
wire v_1345;
wire v_1346;
wire v_1347;
wire v_1348;
wire v_1349;
wire v_1350;
wire v_1351;
wire v_1352;
wire v_1353;
wire v_1354;
wire v_1355;
wire v_1356;
wire v_1359;
wire v_1360;
wire v_1361;
wire v_1362;
wire v_1363;
wire v_1364;
wire v_1365;
wire v_1367;
wire v_1368;
wire v_1369;
wire v_1370;
wire v_1371;
wire v_1372;
wire v_1373;
wire v_1374;
wire v_1375;
wire v_1376;
wire v_1377;
wire v_1378;
wire v_1379;
wire v_1380;
wire v_1381;
wire v_1382;
wire v_1383;
wire v_1384;
wire v_1385;
wire v_1386;
wire v_1388;
wire v_1389;
wire v_1390;
wire v_1391;
wire v_1392;
wire v_1393;
wire v_1394;
wire v_1396;
wire v_1397;
wire v_1398;
wire v_1399;
wire v_1400;
wire v_1401;
wire v_1402;
wire v_1405;
wire v_1406;
wire v_1410;
wire v_1412;
wire v_1413;
wire v_1414;
wire v_1415;
wire v_1416;
wire v_1417;
wire v_1419;
wire v_1420;
wire v_1423;
wire v_1425;
wire v_1426;
wire v_1427;
wire v_1431;
wire v_1433;
wire v_1434;
wire v_1435;
wire v_1436;
wire v_1441;
wire v_1442;
wire v_1443;
wire v_1444;
wire v_1445;
wire v_1446;
wire v_1447;
wire v_1448;
wire v_1449;
wire v_1450;
wire v_1451;
wire v_1452;
wire v_1453;
wire v_1454;
wire v_1455;
wire v_1456;
wire v_1457;
wire v_1458;
wire v_1459;
wire v_1460;
wire v_1461;
wire v_1462;
wire v_1463;
wire v_1464;
wire v_1465;
wire v_1466;
wire v_1467;
wire v_1468;
wire v_1469;
wire v_1470;
wire v_1471;
wire v_1472;
wire v_1473;
wire v_1474;
wire v_1475;
wire v_1476;
wire v_1477;
wire v_1478;
wire v_1479;
wire v_1480;
wire v_1481;
wire v_1482;
wire v_1483;
wire v_1484;
wire v_1485;
wire v_1486;
wire v_1487;
wire v_1488;
wire v_1489;
wire v_1490;
wire v_1491;
wire v_1492;
wire v_1493;
wire v_1494;
wire v_1495;
wire v_1496;
wire v_1497;
wire v_1498;
wire v_1499;
wire v_1500;
wire v_1501;
wire v_1502;
wire v_1503;
wire v_1504;
wire v_1505;
wire v_1506;
wire v_1507;
wire v_1508;
wire v_1509;
wire v_1510;
wire v_1511;
wire v_1512;
wire v_1514;
wire v_1515;
wire v_1516;
wire v_1517;
wire v_1518;
wire v_1519;
wire v_1520;
wire v_1521;
wire v_1522;
wire v_1523;
wire v_1524;
wire v_1525;
wire v_1527;
wire v_1528;
wire v_1531;
wire v_1533;
wire v_1534;
wire v_1535;
wire v_1539;
wire v_1540;
wire v_1541;
wire v_1542;
wire v_1543;
wire v_1544;
wire v_1545;
wire v_1546;
wire v_1547;
wire v_1548;
wire v_1549;
wire v_1550;
wire v_1551;
wire v_1552;
wire v_1553;
wire v_1554;
wire v_1555;
wire v_1556;
wire v_1557;
wire v_1558;
wire v_1559;
wire v_1560;
wire v_1561;
wire v_1562;
wire v_1563;
wire v_1564;
wire v_1565;
wire v_1566;
wire v_1567;
wire v_1568;
wire v_1569;
wire v_1570;
wire v_1571;
wire v_1572;
wire v_1573;
wire v_1574;
wire v_1575;
wire v_1576;
wire v_1577;
wire v_1578;
wire v_1579;
wire v_1580;
wire v_1581;
wire v_1582;
wire v_1583;
wire v_1584;
wire v_1585;
wire v_1586;
wire v_1587;
wire v_1588;
wire v_1589;
wire v_1590;
wire v_1591;
wire v_1592;
wire v_1593;
wire v_1594;
wire v_1595;
wire v_1596;
wire v_1597;
wire v_1598;
wire v_1599;
wire v_1600;
wire v_1601;
wire v_1602;
wire v_1604;
wire v_1606;
wire v_1607;
wire v_1608;
wire v_1609;
wire v_1610;
wire v_1611;
wire v_1612;
wire v_1613;
wire v_1614;
wire v_1615;
wire v_1616;
wire v_1618;
wire v_1619;
wire v_1622;
wire v_1623;
wire v_1624;
wire v_1625;
wire v_1626;
wire v_1627;
wire v_1628;
wire v_1629;
wire v_1630;
wire v_1631;
wire v_1632;
wire v_1633;
wire v_1634;
wire v_1635;
wire v_1636;
wire v_1637;
wire v_1638;
wire v_1639;
wire v_1640;
wire v_1641;
wire v_1642;
wire v_1643;
wire v_1644;
wire v_1645;
wire v_1646;
wire v_1647;
wire v_1648;
wire v_1649;
wire v_1650;
wire v_1651;
wire v_1652;
wire v_1653;
wire v_1654;
wire v_1655;
wire v_1656;
wire v_1657;
wire v_1658;
wire v_1659;
wire v_1660;
wire v_1661;
wire v_1662;
wire v_1663;
wire v_1664;
wire v_1665;
wire v_1666;
wire v_1667;
wire v_1668;
wire v_1669;
wire v_1670;
wire v_1671;
wire v_1672;
wire v_1673;
wire v_1674;
wire v_1675;
wire v_1676;
wire v_1678;
wire v_1680;
wire v_1681;
wire v_1682;
wire v_1683;
wire v_1684;
wire v_1685;
wire v_1686;
wire v_1687;
wire v_1688;
wire v_1689;
wire v_1690;
wire v_1691;
wire v_1692;
wire v_1693;
wire v_1694;
wire v_1695;
wire v_1696;
wire v_1697;
wire v_1698;
wire v_1699;
wire v_1700;
wire v_1701;
wire v_1702;
wire v_1703;
wire v_1704;
wire v_1705;
wire v_1706;
wire v_1707;
wire v_1708;
wire v_1709;
wire v_1710;
wire v_1711;
wire v_1712;
wire v_1713;
wire v_1714;
wire v_1715;
wire v_1716;
wire v_1717;
wire v_1718;
wire v_1719;
wire v_1720;
wire v_1721;
wire v_1722;
wire v_1723;
wire v_1724;
wire v_1725;
wire v_1727;
wire v_1729;
wire v_1730;
wire v_1731;
wire v_1732;
wire v_1733;
wire v_1734;
wire v_1735;
wire v_1736;
wire v_1737;
wire v_1738;
wire v_1739;
wire v_1740;
wire v_1741;
wire v_1742;
wire v_1743;
wire v_1744;
wire v_1748;
wire v_1753;
wire v_1754;
wire v_1755;
wire v_1756;
wire v_1757;
wire v_1758;
wire v_1759;
wire v_1760;
wire v_1761;
wire v_1762;
wire v_1763;
wire v_1764;
wire v_1765;
wire v_1766;
wire v_1767;
wire v_1768;
wire v_1769;
wire v_1771;
wire v_1773;
wire v_1774;
wire v_1775;
wire v_1776;
wire v_1777;
wire v_1778;
wire v_1779;
wire v_1780;
wire v_1781;
wire v_1782;
wire v_1783;
wire v_1784;
wire v_1785;
wire v_1787;
wire v_1789;
wire v_1791;
wire v_1792;
wire v_1793;
wire v_1794;
wire v_1795;
wire v_1796;
wire v_1797;
wire v_1798;
wire v_1799;
wire v_1800;
wire v_1801;
wire v_1802;
wire v_1803;
wire v_1805;
wire v_1807;
wire v_1809;
wire v_1811;
wire v_1812;
wire v_1813;
wire v_1814;
wire v_1815;
wire v_1816;
wire v_1817;
wire v_1818;
wire v_1819;
wire v_1820;
wire v_1821;
wire v_1822;
wire v_1823;
wire v_1824;
wire v_1825;
wire v_1826;
wire v_1827;
wire v_1828;
wire v_1829;
wire v_1830;
wire v_1831;
wire v_1832;
wire v_1833;
wire v_1834;
wire v_1835;
wire v_1836;
wire v_1837;
wire v_1838;
wire v_1839;
wire v_1840;
wire v_1841;
wire v_1842;
wire v_1843;
wire v_1844;
wire v_1845;
wire v_1846;
wire v_1847;
wire v_1850;
wire v_1851;
wire v_1852;
wire v_1853;
wire v_1854;
wire v_1855;
wire v_1856;
wire v_1858;
wire v_1859;
wire v_1860;
wire v_1861;
wire v_1862;
wire v_1863;
wire v_1864;
wire v_1865;
wire v_1866;
wire v_1867;
wire v_1868;
wire v_1869;
wire v_1870;
wire v_1871;
wire v_1872;
wire v_1873;
wire v_1874;
wire v_1875;
wire v_1876;
wire v_1877;
wire v_1879;
wire v_1880;
wire v_1881;
wire v_1882;
wire v_1883;
wire v_1884;
wire v_1885;
wire v_1887;
wire v_1888;
wire v_1889;
wire v_1890;
wire v_1891;
wire v_1892;
wire v_1893;
wire v_1894;
wire v_1895;
wire v_1896;
wire v_1897;
wire v_1898;
wire v_1899;
wire v_1900;
wire v_1901;
wire v_1902;
wire v_1903;
wire v_1904;
wire v_1905;
wire v_1906;
wire v_1907;
wire v_1908;
wire v_1909;
wire v_1910;
wire v_1911;
wire v_1912;
wire v_1913;
wire v_1914;
wire v_1915;
wire v_1918;
wire v_1919;
wire v_1920;
wire v_1921;
wire v_1922;
wire v_1923;
wire v_1924;
wire v_1926;
wire v_1927;
wire v_1928;
wire v_1929;
wire v_1930;
wire v_1931;
wire v_1932;
wire v_1933;
wire v_1934;
wire v_1935;
wire v_1936;
wire v_1937;
wire v_1938;
wire v_1939;
wire v_1940;
wire v_1941;
wire v_1942;
wire v_1943;
wire v_1944;
wire v_1945;
wire v_1947;
wire v_1948;
wire v_1949;
wire v_1950;
wire v_1951;
wire v_1952;
wire v_1953;
wire v_1955;
wire v_1956;
wire v_1957;
wire v_1958;
wire v_1959;
wire v_1960;
wire v_1961;
wire v_1962;
wire v_1963;
wire v_1964;
wire v_1965;
wire v_1966;
wire v_1967;
wire v_1968;
wire v_1969;
wire v_1970;
wire v_1971;
wire v_1972;
wire v_1973;
wire v_1974;
wire v_1975;
wire v_1976;
wire v_1977;
wire v_1978;
wire v_1979;
wire v_1980;
wire v_1981;
wire v_1982;
wire v_1983;
wire v_1986;
wire v_1987;
wire v_1988;
wire v_1989;
wire v_1990;
wire v_1991;
wire v_1992;
wire v_1994;
wire v_1995;
wire v_1996;
wire v_1997;
wire v_1998;
wire v_1999;
wire v_2000;
wire v_2001;
wire v_2002;
wire v_2003;
wire v_2004;
wire v_2005;
wire v_2006;
wire v_2007;
wire v_2008;
wire v_2009;
wire v_2010;
wire v_2011;
wire v_2012;
wire v_2013;
wire v_2015;
wire v_2016;
wire v_2017;
wire v_2018;
wire v_2019;
wire v_2020;
wire v_2021;
wire v_2023;
wire v_2024;
wire v_2025;
wire v_2026;
wire v_2027;
wire v_2028;
wire v_2029;
wire v_2030;
wire v_2031;
wire v_2032;
wire v_2033;
wire v_2034;
wire v_2035;
wire v_2036;
wire v_2037;
wire v_2038;
wire v_2039;
wire v_2040;
wire v_2041;
wire v_2042;
wire v_2043;
wire v_2044;
wire v_2045;
wire v_2046;
wire v_2047;
wire v_2048;
wire v_2049;
wire v_2050;
wire v_2051;
wire v_2054;
wire v_2055;
wire v_2056;
wire v_2057;
wire v_2058;
wire v_2059;
wire v_2060;
wire v_2062;
wire v_2063;
wire v_2064;
wire v_2065;
wire v_2066;
wire v_2067;
wire v_2068;
wire v_2069;
wire v_2070;
wire v_2071;
wire v_2072;
wire v_2073;
wire v_2074;
wire v_2075;
wire v_2076;
wire v_2077;
wire v_2078;
wire v_2079;
wire v_2080;
wire v_2081;
wire v_2083;
wire v_2084;
wire v_2085;
wire v_2086;
wire v_2087;
wire v_2088;
wire v_2089;
wire v_2091;
wire v_2092;
wire v_2093;
wire v_2094;
wire v_2095;
wire v_2096;
wire v_2097;
wire v_2100;
wire v_2101;
wire v_2105;
wire v_2107;
wire v_2108;
wire v_2109;
wire v_2111;
wire v_2112;
wire v_2115;
wire v_2117;
wire v_2118;
wire v_2119;
wire v_2123;
wire v_2125;
wire v_2126;
wire v_2127;
wire v_2128;
wire v_2133;
wire v_2134;
wire v_2135;
wire v_2136;
wire v_2137;
wire v_2138;
wire v_2139;
wire v_2140;
wire v_2141;
wire v_2142;
wire v_2143;
wire v_2144;
wire v_2145;
wire v_2146;
wire v_2147;
wire v_2148;
wire v_2149;
wire v_2150;
wire v_2151;
wire v_2152;
wire v_2153;
wire v_2154;
wire v_2155;
wire v_2156;
wire v_2157;
wire v_2158;
wire v_2159;
wire v_2160;
wire v_2161;
wire v_2162;
wire v_2163;
wire v_2164;
wire v_2165;
wire v_2166;
wire v_2167;
wire v_2168;
wire v_2170;
wire v_2172;
wire v_2173;
wire v_2174;
wire v_2175;
wire v_2176;
wire v_2178;
wire v_2179;
wire v_2182;
wire v_2184;
wire v_2185;
wire v_2186;
wire v_2190;
wire v_2191;
wire v_2192;
wire v_2193;
wire v_2194;
wire v_2195;
wire v_2196;
wire v_2197;
wire v_2198;
wire v_2199;
wire v_2200;
wire v_2201;
wire v_2202;
wire v_2203;
wire v_2204;
wire v_2205;
wire v_2206;
wire v_2207;
wire v_2208;
wire v_2209;
wire v_2210;
wire v_2211;
wire v_2212;
wire v_2213;
wire v_2214;
wire v_2215;
wire v_2216;
wire v_2218;
wire v_2220;
wire v_2221;
wire v_2222;
wire v_2223;
wire v_2224;
wire v_2226;
wire v_2227;
wire v_2230;
wire v_2231;
wire v_2232;
wire v_2233;
wire v_2234;
wire v_2235;
wire v_2236;
wire v_2237;
wire v_2238;
wire v_2239;
wire v_2240;
wire v_2241;
wire v_2242;
wire v_2243;
wire v_2244;
wire v_2245;
wire v_2246;
wire v_2247;
wire v_2249;
wire v_2251;
wire v_2252;
wire v_2253;
wire v_2254;
wire v_2255;
wire v_2256;
wire v_2257;
wire v_2258;
wire v_2259;
wire v_2260;
wire v_2261;
wire v_2262;
wire v_2264;
wire v_2266;
wire v_2267;
wire v_2268;
wire v_2269;
wire v_2270;
wire v_2271;
wire v_2272;
wire v_2273;
wire v_2274;
wire v_2275;
wire v_2276;
wire v_2277;
wire v_2278;
wire v_2279;
wire v_2281;
wire v_2282;
wire v_2283;
wire v_2284;
wire v_2285;
wire v_2286;
wire v_2287;
wire v_2288;
wire v_2289;
wire v_2290;
wire v_2291;
wire v_2292;
wire v_2293;
wire v_2294;
wire v_2295;
wire v_2296;
wire v_2297;
wire v_2298;
wire v_2299;
wire v_2300;
wire v_2301;
wire v_2302;
wire v_2303;
wire v_2304;
wire v_2305;
wire v_2306;
wire v_2307;
wire v_2308;
wire v_2309;
wire v_2310;
wire v_2311;
wire v_2312;
wire v_2313;
wire v_2314;
wire v_2315;
wire v_2316;
wire v_2317;
wire v_2318;
wire v_2319;
wire v_2320;
wire v_2321;
wire v_2322;
wire v_2323;
wire v_2324;
wire v_2325;
wire v_2326;
wire v_2327;
wire v_2328;
wire v_2329;
wire v_2330;
wire v_2331;
wire v_2332;
wire v_2333;
wire v_2335;
wire v_2337;
wire v_2338;
wire v_2339;
wire v_2340;
wire v_2341;
wire v_2342;
wire v_2343;
wire v_2344;
wire v_2345;
wire v_2346;
wire v_2347;
wire v_2348;
wire v_2349;
wire v_2350;
wire v_2351;
wire v_2352;
wire v_2353;
wire v_2354;
wire v_2355;
wire v_2356;
wire v_2357;
wire v_2358;
wire v_2359;
wire v_2360;
wire v_2361;
wire v_2363;
wire v_2365;
wire v_2367;
wire v_2368;
wire v_2369;
wire v_2370;
wire v_2371;
wire v_2372;
wire v_2373;
wire v_2374;
wire v_2375;
wire v_2376;
wire v_2377;
wire v_2378;
wire v_2379;
wire v_2380;
wire v_2381;
wire v_2382;
wire v_2383;
wire v_2384;
wire v_2385;
wire v_2386;
wire v_2387;
wire v_2388;
wire v_2389;
wire v_2390;
wire v_2391;
wire v_2393;
wire v_2395;
wire v_2397;
wire v_2399;
wire v_2400;
wire v_2401;
wire v_2402;
wire v_2403;
wire v_2404;
wire v_2405;
wire v_2406;
wire v_2407;
wire v_2408;
wire v_2409;
wire v_2410;
wire v_2411;
wire v_2412;
wire v_2413;
wire v_2414;
wire v_2415;
wire v_2416;
wire v_2417;
wire v_2418;
wire v_2419;
wire v_2420;
wire v_2421;
wire v_2422;
wire v_2423;
wire v_2424;
wire v_2425;
wire v_2426;
wire v_2427;
wire v_2428;
wire v_2429;
wire v_2430;
wire v_2431;
wire v_2432;
wire v_2433;
wire v_2434;
wire v_2435;
wire v_2436;
wire v_2437;
wire v_2438;
wire v_2439;
wire v_2440;
wire v_2441;
wire v_2442;
wire v_2443;
wire v_2444;
wire v_2445;
wire v_2446;
wire v_2447;
wire v_2448;
wire v_2449;
wire v_2450;
wire v_2451;
wire v_2454;
wire v_2455;
wire v_2456;
wire v_2457;
wire v_2458;
wire v_2459;
wire v_2460;
wire v_2461;
wire v_2463;
wire v_2464;
wire v_2465;
wire v_2466;
wire v_2467;
wire v_2468;
wire v_2469;
wire v_2470;
wire v_2471;
wire v_2472;
wire v_2473;
wire v_2474;
wire v_2475;
wire v_2476;
wire v_2477;
wire v_2478;
wire v_2479;
wire v_2480;
wire v_2481;
wire v_2482;
wire v_2483;
wire v_2484;
wire v_2485;
wire v_2486;
wire v_2487;
wire v_2488;
wire v_2489;
wire v_2490;
wire v_2491;
wire v_2492;
wire v_2494;
wire v_2495;
wire v_2496;
wire v_2497;
wire v_2498;
wire v_2499;
wire v_2500;
wire v_2501;
wire v_2503;
wire v_2504;
wire v_2505;
wire v_2506;
wire v_2507;
wire v_2508;
wire v_2509;
wire v_2510;
wire v_2511;
wire v_2512;
wire v_2513;
wire v_2514;
wire v_2515;
wire v_2516;
wire v_2517;
wire v_2518;
wire v_2519;
wire v_2520;
wire v_2521;
wire v_2522;
wire v_2523;
wire v_2524;
wire v_2525;
wire v_2526;
wire v_2527;
wire v_2528;
wire v_2529;
wire v_2534;
wire v_2535;
wire v_2536;
wire v_2537;
wire v_2538;
wire v_2539;
wire v_2540;
wire v_2541;
wire v_2542;
wire v_2544;
wire v_2545;
wire v_2546;
wire v_2547;
wire v_2548;
wire v_2549;
wire v_2550;
wire v_2551;
wire v_2552;
wire v_2553;
wire v_2554;
wire v_2555;
wire v_2556;
wire v_2557;
wire v_2558;
wire v_2559;
wire v_2560;
wire v_2561;
wire v_2562;
wire v_2563;
wire v_2565;
wire v_2566;
wire v_2567;
wire v_2568;
wire v_2569;
wire v_2570;
wire v_2571;
wire v_2572;
wire v_2573;
wire v_2575;
wire v_2576;
wire v_2577;
wire v_2578;
wire v_2579;
wire v_2580;
wire v_2581;
wire v_2582;
wire v_2583;
wire v_2584;
wire v_2585;
wire v_2586;
wire v_2587;
wire v_2588;
wire v_2589;
wire v_2590;
wire v_2591;
wire v_2592;
wire v_2593;
wire v_2594;
wire v_2595;
wire v_2596;
wire v_2597;
wire v_2598;
wire v_2599;
wire v_2600;
wire v_2601;
wire v_2602;
wire v_2603;
wire v_2608;
wire v_2609;
wire v_2610;
wire v_2611;
wire v_2612;
wire v_2613;
wire v_2614;
wire v_2615;
wire v_2616;
wire v_2618;
wire v_2619;
wire v_2620;
wire v_2621;
wire v_2622;
wire v_2623;
wire v_2624;
wire v_2625;
wire v_2626;
wire v_2627;
wire v_2628;
wire v_2629;
wire v_2630;
wire v_2631;
wire v_2632;
wire v_2633;
wire v_2634;
wire v_2635;
wire v_2636;
wire v_2637;
wire v_2639;
wire v_2640;
wire v_2641;
wire v_2642;
wire v_2643;
wire v_2644;
wire v_2645;
wire v_2646;
wire v_2647;
wire v_2649;
wire v_2650;
wire v_2651;
wire v_2652;
wire v_2653;
wire v_2654;
wire v_2655;
wire v_2656;
wire v_2657;
wire v_2658;
wire v_2659;
wire v_2660;
wire v_2661;
wire v_2662;
wire v_2663;
wire v_2664;
wire v_2665;
wire v_2666;
wire v_2667;
wire v_2668;
wire v_2669;
wire v_2670;
wire v_2671;
wire v_2672;
wire v_2673;
wire v_2674;
wire v_2675;
wire v_2676;
wire v_2677;
wire v_2682;
wire v_2683;
wire v_2684;
wire v_2685;
wire v_2686;
wire v_2687;
wire v_2688;
wire v_2689;
wire v_2690;
wire v_2692;
wire v_2693;
wire v_2694;
wire v_2695;
wire v_2696;
wire v_2697;
wire v_2698;
wire v_2699;
wire v_2700;
wire v_2701;
wire v_2702;
wire v_2703;
wire v_2704;
wire v_2705;
wire v_2706;
wire v_2707;
wire v_2708;
wire v_2709;
wire v_2710;
wire v_2711;
wire v_2713;
wire v_2714;
wire v_2715;
wire v_2716;
wire v_2717;
wire v_2718;
wire v_2719;
wire v_2720;
wire v_2721;
wire v_2723;
wire v_2724;
wire v_2725;
wire v_2726;
wire v_2727;
wire v_2728;
wire v_2729;
wire v_2730;
wire v_2731;
wire v_2732;
wire v_2733;
wire v_2734;
wire v_2735;
wire v_2736;
wire v_2737;
wire v_2738;
wire v_2739;
wire v_2740;
wire v_2741;
wire v_2742;
wire v_2743;
wire v_2744;
wire v_2745;
wire v_2746;
wire v_2747;
wire v_2748;
wire v_2749;
wire v_2750;
wire v_2751;
wire v_2756;
wire v_2757;
wire v_2758;
wire v_2759;
wire v_2760;
wire v_2761;
wire v_2762;
wire v_2763;
wire v_2764;
wire v_2766;
wire v_2767;
wire v_2768;
wire v_2769;
wire v_2770;
wire v_2771;
wire v_2772;
wire v_2773;
wire v_2774;
wire v_2775;
wire v_2776;
wire v_2777;
wire v_2778;
wire v_2779;
wire v_2780;
wire v_2781;
wire v_2782;
wire v_2783;
wire v_2784;
wire v_2785;
wire v_2787;
wire v_2788;
wire v_2789;
wire v_2790;
wire v_2791;
wire v_2792;
wire v_2793;
wire v_2794;
wire v_2795;
wire v_2797;
wire v_2798;
wire v_2799;
wire v_2800;
wire v_2801;
wire v_2802;
wire v_2803;
wire v_2806;
wire v_2807;
wire v_2811;
wire v_2813;
wire v_2814;
wire v_2815;
wire v_2817;
wire v_2818;
wire v_2821;
wire v_2823;
wire v_2824;
wire v_2825;
wire v_2829;
wire v_2831;
wire v_2832;
wire v_2833;
wire v_2834;
wire v_2839;
wire v_2840;
wire v_2841;
wire v_2842;
wire v_2843;
wire v_2844;
wire v_2845;
wire v_2846;
wire v_2847;
wire v_2848;
wire v_2849;
wire v_2850;
wire v_2851;
wire v_2852;
wire v_2853;
wire v_2854;
wire v_2855;
wire v_2856;
wire v_2857;
wire v_2858;
wire v_2859;
wire v_2860;
wire v_2861;
wire v_2862;
wire v_2863;
wire v_2864;
wire v_2865;
wire v_2866;
wire v_2867;
wire v_2868;
wire v_2869;
wire v_2870;
wire v_2871;
wire v_2872;
wire v_2873;
wire v_2874;
wire v_2876;
wire v_2878;
wire v_2879;
wire v_2880;
wire v_2881;
wire v_2883;
wire v_2884;
wire v_2887;
wire v_2889;
wire v_2890;
wire v_2891;
wire v_2895;
wire v_2896;
wire v_2897;
wire v_2898;
wire v_2899;
wire v_2900;
wire v_2901;
wire v_2902;
wire v_2903;
wire v_2904;
wire v_2905;
wire v_2906;
wire v_2907;
wire v_2908;
wire v_2909;
wire v_2910;
wire v_2911;
wire v_2912;
wire v_2913;
wire v_2914;
wire v_2915;
wire v_2916;
wire v_2917;
wire v_2918;
wire v_2919;
wire v_2920;
wire v_2921;
wire v_2923;
wire v_2925;
wire v_2926;
wire v_2927;
wire v_2928;
wire v_2930;
wire v_2931;
wire v_2934;
wire v_2935;
wire v_2936;
wire v_2937;
wire v_2938;
wire v_2939;
wire v_2940;
wire v_2941;
wire v_2942;
wire v_2943;
wire v_2944;
wire v_2945;
wire v_2946;
wire v_2947;
wire v_2948;
wire v_2949;
wire v_2950;
wire v_2951;
wire v_2953;
wire v_2955;
wire v_2956;
wire v_2957;
wire v_2958;
wire v_2959;
wire v_2960;
wire v_2961;
wire v_2962;
wire v_2963;
wire v_2964;
wire v_2965;
wire v_2966;
wire v_2968;
wire v_2970;
wire v_2971;
wire v_2972;
wire v_2973;
wire v_2974;
wire v_2975;
wire v_2976;
wire v_2977;
wire v_2978;
wire v_2979;
wire v_2980;
wire v_2981;
wire v_2982;
wire v_2983;
wire v_2984;
wire v_2985;
wire v_2986;
wire v_2987;
wire v_2989;
wire v_2990;
wire v_2991;
wire v_2992;
wire v_2993;
wire v_2994;
wire v_2995;
wire v_2996;
wire v_2997;
wire v_2998;
wire v_2999;
wire v_3000;
wire v_3001;
wire v_3002;
wire v_3003;
wire v_3004;
wire v_3005;
wire v_3006;
wire v_3007;
wire v_3008;
wire v_3009;
wire v_3010;
wire v_3011;
wire v_3012;
wire v_3014;
wire v_3015;
wire v_3016;
wire v_3017;
wire v_3018;
wire v_3019;
wire v_3020;
wire v_3021;
wire v_3022;
wire v_3023;
wire v_3024;
wire v_3025;
wire v_3026;
wire v_3027;
wire v_3029;
wire v_3031;
wire v_3032;
wire v_3033;
wire v_3034;
wire v_3035;
wire v_3036;
wire v_3037;
wire v_3038;
wire v_3039;
wire v_3040;
wire v_3041;
wire v_3042;
wire v_3043;
wire v_3045;
wire v_3046;
wire v_3048;
wire v_3049;
wire v_3051;
wire v_3053;
wire v_3054;
wire v_3055;
wire v_3056;
wire v_3057;
wire v_3058;
wire v_3059;
wire v_3060;
wire v_3061;
wire v_3062;
wire v_3063;
wire v_3064;
wire v_3065;
wire v_3066;
wire v_3067;
wire v_3068;
wire v_3069;
wire v_3070;
wire v_3071;
wire v_3072;
wire v_3073;
wire v_3074;
wire v_3075;
wire v_3076;
wire v_3077;
wire v_3078;
wire v_3079;
wire v_3081;
wire v_3082;
wire v_3083;
wire v_3084;
wire v_3085;
wire v_3086;
wire v_3087;
wire v_3089;
wire v_3090;
wire v_3091;
wire v_3092;
wire v_3093;
wire v_3094;
wire v_3095;
wire v_3096;
wire v_3097;
wire v_3098;
wire v_3099;
wire v_3100;
wire v_3101;
wire v_3102;
wire v_3103;
wire v_3104;
wire v_3105;
wire v_3106;
wire v_3107;
wire v_3108;
wire v_3110;
wire v_3111;
wire v_3112;
wire v_3113;
wire v_3114;
wire v_3115;
wire v_3116;
wire v_3118;
wire v_3119;
wire v_3120;
wire v_3121;
wire v_3122;
wire v_3123;
wire v_3124;
wire v_3125;
wire v_3126;
wire v_3127;
wire v_3128;
wire v_3129;
wire v_3130;
wire v_3131;
wire v_3132;
wire v_3133;
wire v_3134;
wire v_3135;
wire v_3136;
wire v_3137;
wire v_3138;
wire v_3139;
wire v_3140;
wire v_3141;
wire v_3142;
wire v_3143;
wire v_3144;
wire v_3145;
wire v_3146;
wire v_3148;
wire v_3149;
wire v_3150;
wire v_3151;
wire v_3152;
wire v_3153;
wire v_3154;
wire v_3156;
wire v_3157;
wire v_3158;
wire v_3159;
wire v_3160;
wire v_3161;
wire v_3162;
wire v_3163;
wire v_3164;
wire v_3165;
wire v_3166;
wire v_3167;
wire v_3168;
wire v_3169;
wire v_3170;
wire v_3171;
wire v_3172;
wire v_3173;
wire v_3174;
wire v_3175;
wire v_3177;
wire v_3178;
wire v_3179;
wire v_3180;
wire v_3181;
wire v_3182;
wire v_3183;
wire v_3185;
wire v_3186;
wire v_3187;
wire v_3188;
wire v_3189;
wire v_3190;
wire v_3191;
wire v_3192;
wire v_3193;
wire v_3194;
wire v_3195;
wire v_3196;
wire v_3197;
wire v_3198;
wire v_3199;
wire v_3200;
wire v_3201;
wire v_3202;
wire v_3203;
wire v_3204;
wire v_3205;
wire v_3206;
wire v_3207;
wire v_3208;
wire v_3209;
wire v_3210;
wire v_3211;
wire v_3212;
wire v_3213;
wire v_3215;
wire v_3216;
wire v_3217;
wire v_3218;
wire v_3219;
wire v_3220;
wire v_3221;
wire v_3223;
wire v_3224;
wire v_3225;
wire v_3226;
wire v_3227;
wire v_3228;
wire v_3229;
wire v_3230;
wire v_3231;
wire v_3232;
wire v_3233;
wire v_3234;
wire v_3235;
wire v_3236;
wire v_3237;
wire v_3238;
wire v_3239;
wire v_3240;
wire v_3241;
wire v_3242;
wire v_3244;
wire v_3245;
wire v_3246;
wire v_3247;
wire v_3248;
wire v_3249;
wire v_3250;
wire v_3252;
wire v_3253;
wire v_3254;
wire v_3255;
wire v_3256;
wire v_3257;
wire v_3258;
wire v_3261;
wire v_3262;
wire v_3263;
wire v_3264;
wire v_3265;
wire v_3266;
wire v_3267;
wire v_3268;
wire v_3269;
wire v_3270;
wire v_3271;
wire v_3272;
wire v_3273;
wire v_3274;
wire v_3275;
wire v_3276;
wire v_3277;
wire v_3278;
wire v_3279;
wire v_3280;
wire v_3281;
wire v_3282;
wire v_3283;
wire v_3284;
wire v_3285;
wire v_3286;
wire v_3287;
wire v_3288;
wire v_3289;
wire v_3290;
wire v_3291;
wire v_3292;
wire v_3293;
wire v_3294;
wire v_3295;
wire v_3296;
wire v_3297;
wire v_3298;
wire v_3299;
wire v_3300;
wire v_3301;
wire v_3302;
wire v_3303;
wire v_3304;
wire v_3305;
wire v_3306;
wire v_3307;
wire v_3308;
wire v_3309;
wire v_3310;
wire v_3311;
wire v_3312;
wire v_3313;
wire v_3314;
wire v_3315;
wire v_3316;
wire v_3317;
wire v_3318;
wire v_3319;
wire v_3320;
wire v_3321;
wire v_3322;
wire v_3323;
wire v_3324;
wire v_3325;
wire v_3326;
wire v_3327;
wire v_3328;
wire v_3329;
wire v_3330;
wire v_3331;
wire v_3332;
wire v_3333;
wire v_3334;
wire v_3335;
wire v_3336;
wire v_3337;
wire v_3338;
wire v_3339;
wire v_3340;
wire v_3341;
wire v_3342;
wire v_3343;
wire v_3344;
wire v_3345;
wire v_3346;
wire v_3347;
wire v_3348;
wire v_3349;
wire v_3350;
wire v_3351;
wire v_3352;
wire v_3353;
wire v_3354;
wire v_3355;
wire v_3356;
wire v_3357;
wire v_3358;
wire v_3359;
wire v_3360;
wire v_3361;
wire v_3362;
wire v_3363;
wire x_1;
wire x_2;
wire x_3;
wire x_4;
wire x_5;
wire x_6;
wire x_7;
wire x_8;
wire x_9;
wire x_10;
wire x_11;
wire x_12;
wire x_13;
wire x_14;
wire x_15;
wire x_16;
wire x_17;
wire x_18;
wire x_19;
wire x_20;
wire x_21;
wire x_22;
wire x_23;
wire x_24;
wire x_25;
wire x_26;
wire x_27;
wire x_28;
wire x_29;
wire x_30;
wire x_31;
wire x_32;
wire x_33;
wire x_34;
wire x_35;
wire x_36;
wire x_37;
wire x_38;
wire x_39;
wire x_40;
wire x_41;
wire x_42;
wire x_43;
wire x_44;
wire x_45;
wire x_46;
wire x_47;
wire x_48;
wire x_49;
wire x_50;
wire x_51;
wire x_52;
wire x_53;
wire x_54;
wire x_55;
wire x_56;
wire x_57;
wire x_58;
wire x_59;
wire x_60;
wire x_61;
wire x_62;
wire x_63;
wire x_64;
wire x_65;
wire x_66;
wire x_67;
wire x_68;
wire x_69;
wire x_70;
wire x_71;
wire x_72;
wire x_73;
wire x_74;
wire x_75;
wire x_76;
wire x_77;
wire x_78;
wire x_79;
wire x_80;
wire x_81;
wire x_82;
wire x_83;
wire x_84;
wire x_85;
wire x_86;
wire x_87;
wire x_88;
wire x_89;
wire x_90;
wire x_91;
wire x_92;
wire x_93;
wire x_94;
wire x_95;
wire x_96;
wire x_97;
wire x_98;
wire x_99;
wire x_100;
wire x_101;
wire x_102;
wire x_103;
wire x_104;
wire x_105;
wire x_106;
wire x_107;
wire x_108;
wire x_109;
wire x_110;
wire x_111;
wire x_112;
wire x_113;
wire x_114;
wire x_115;
wire x_116;
wire x_117;
wire x_118;
wire x_119;
wire x_120;
wire x_121;
wire x_122;
wire x_123;
wire x_124;
wire x_125;
wire x_126;
wire x_127;
wire x_128;
wire x_129;
wire x_130;
wire x_131;
wire x_132;
wire x_133;
wire x_134;
wire x_135;
wire x_136;
wire x_137;
wire x_138;
wire x_139;
wire x_140;
wire x_141;
wire x_142;
wire x_143;
wire x_144;
wire x_145;
wire x_146;
wire x_147;
wire x_148;
wire x_149;
wire x_150;
wire x_151;
wire x_152;
wire x_153;
wire x_154;
wire x_155;
wire x_156;
wire x_157;
wire x_158;
wire x_159;
wire x_160;
wire x_161;
wire x_162;
wire x_163;
wire x_164;
wire x_165;
wire x_166;
wire x_167;
wire x_168;
wire x_169;
wire x_170;
wire x_171;
wire x_172;
wire x_173;
wire x_174;
wire x_175;
wire x_176;
wire x_177;
wire x_178;
wire x_179;
wire x_180;
wire x_181;
wire x_182;
wire x_183;
wire x_184;
wire x_185;
wire x_186;
wire x_187;
wire x_188;
wire x_189;
wire x_190;
wire x_191;
wire x_192;
wire x_193;
wire x_194;
wire x_195;
wire x_196;
wire x_197;
wire x_198;
wire x_199;
wire x_200;
wire x_201;
wire x_202;
wire x_203;
wire x_204;
wire x_205;
wire x_206;
wire x_207;
wire x_208;
wire x_209;
wire x_210;
wire x_211;
wire x_212;
wire x_213;
wire x_214;
wire x_215;
wire x_216;
wire x_217;
wire x_218;
wire x_219;
wire x_220;
wire x_221;
wire x_222;
wire x_223;
wire x_224;
wire x_225;
wire x_226;
wire x_227;
wire x_228;
wire x_229;
wire x_230;
wire x_231;
wire x_232;
wire x_233;
wire x_234;
wire x_235;
wire x_236;
wire x_237;
wire x_238;
wire x_239;
wire x_240;
wire x_241;
wire x_242;
wire x_243;
wire x_244;
wire x_245;
wire x_246;
wire x_247;
wire x_248;
wire x_249;
wire x_250;
wire x_251;
wire x_252;
wire x_253;
wire x_254;
wire x_255;
wire x_256;
wire x_257;
wire x_258;
wire x_259;
wire x_260;
wire x_261;
wire x_262;
wire x_263;
wire x_264;
wire x_265;
wire x_266;
wire x_267;
wire x_268;
wire x_269;
wire x_270;
wire x_271;
wire x_272;
wire x_273;
wire x_274;
wire x_275;
wire x_276;
wire x_277;
wire x_278;
wire x_279;
wire x_280;
wire x_281;
wire x_282;
wire x_283;
wire x_284;
wire x_285;
wire x_286;
wire x_287;
wire x_288;
wire x_289;
wire x_290;
wire x_291;
wire x_292;
wire x_293;
wire x_294;
wire x_295;
wire x_296;
wire x_297;
wire x_298;
wire x_299;
wire x_300;
wire x_301;
wire x_302;
wire x_303;
wire x_304;
wire x_305;
wire x_306;
wire x_307;
wire x_308;
wire x_309;
wire x_310;
wire x_311;
wire x_312;
wire x_313;
wire x_314;
wire x_315;
wire x_316;
wire x_317;
wire x_318;
wire x_319;
wire x_320;
wire x_321;
wire x_322;
wire x_323;
wire x_324;
wire x_325;
wire x_326;
wire x_327;
wire x_328;
wire x_329;
wire x_330;
wire x_331;
wire x_332;
wire x_333;
wire x_334;
wire x_335;
wire x_336;
wire x_337;
wire x_338;
wire x_339;
wire x_340;
wire x_341;
wire x_342;
wire x_343;
wire x_344;
wire x_345;
wire x_346;
wire x_347;
wire x_348;
wire x_349;
wire x_350;
wire x_351;
wire x_352;
wire x_353;
wire x_354;
wire x_355;
wire x_356;
wire x_357;
wire x_358;
wire x_359;
wire x_360;
wire x_361;
wire x_362;
wire x_363;
wire x_364;
wire x_365;
wire x_366;
wire x_367;
wire x_368;
wire x_369;
wire x_370;
wire x_371;
wire x_372;
wire x_373;
wire x_374;
wire x_375;
wire x_376;
wire x_377;
wire x_378;
wire x_379;
wire x_380;
wire x_381;
wire x_382;
wire x_383;
wire x_384;
wire x_385;
wire x_386;
wire x_387;
wire x_388;
wire x_389;
wire x_390;
wire x_391;
wire x_392;
wire x_393;
wire x_394;
wire x_395;
wire x_396;
wire x_397;
wire x_398;
wire x_399;
wire x_400;
wire x_401;
wire x_402;
wire x_403;
wire x_404;
wire x_405;
wire x_406;
wire x_407;
wire x_408;
wire x_409;
wire x_410;
wire x_411;
wire x_412;
wire x_413;
wire x_414;
wire x_415;
wire x_416;
wire x_417;
wire x_418;
wire x_419;
wire x_420;
wire x_421;
wire x_422;
wire x_423;
wire x_424;
wire x_425;
wire x_426;
wire x_427;
wire x_428;
wire x_429;
wire x_430;
wire x_431;
wire x_432;
wire x_433;
wire x_434;
wire x_435;
wire x_436;
wire x_437;
wire x_438;
wire x_439;
wire x_440;
wire x_441;
wire x_442;
wire x_443;
wire x_444;
wire x_445;
wire x_446;
wire x_447;
wire x_448;
wire x_449;
wire x_450;
wire x_451;
wire x_452;
wire x_453;
wire x_454;
wire x_455;
wire x_456;
wire x_457;
wire x_458;
wire x_459;
wire x_460;
wire x_461;
wire x_462;
wire x_463;
wire x_464;
wire x_465;
wire x_466;
wire x_467;
wire x_468;
wire x_469;
wire x_470;
wire x_471;
wire x_472;
wire x_473;
wire x_474;
wire x_475;
wire x_476;
wire x_477;
wire x_478;
wire x_479;
wire x_480;
wire x_481;
wire x_482;
wire x_483;
wire x_484;
wire x_485;
wire x_486;
wire x_487;
wire x_488;
wire x_489;
wire x_490;
wire x_491;
wire x_492;
wire x_493;
wire x_494;
wire x_495;
wire x_496;
wire x_497;
wire x_498;
wire x_499;
wire x_500;
wire x_501;
wire x_502;
wire x_503;
wire x_504;
wire x_505;
wire x_506;
wire x_507;
wire x_508;
wire x_509;
wire x_510;
wire x_511;
wire x_512;
wire x_513;
wire x_514;
wire x_515;
wire x_516;
wire x_517;
wire x_518;
wire x_519;
wire x_520;
wire x_521;
wire x_522;
wire x_523;
wire x_524;
wire x_525;
wire x_526;
wire x_527;
wire x_528;
wire x_529;
wire x_530;
wire x_531;
wire x_532;
wire x_533;
wire x_534;
wire x_535;
wire x_536;
wire x_537;
wire x_538;
wire x_539;
wire x_540;
wire x_541;
wire x_542;
wire x_543;
wire x_544;
wire x_545;
wire x_546;
wire x_547;
wire x_548;
wire x_549;
wire x_550;
wire x_551;
wire x_552;
wire x_553;
wire x_554;
wire x_555;
wire x_556;
wire x_557;
wire x_558;
wire x_559;
wire x_560;
wire x_561;
wire x_562;
wire x_563;
wire x_564;
wire x_565;
wire x_566;
wire x_567;
wire x_568;
wire x_569;
wire x_570;
wire x_571;
wire x_572;
wire x_573;
wire x_574;
wire x_575;
wire x_576;
wire x_577;
wire x_578;
wire x_579;
wire x_580;
wire x_581;
wire x_582;
wire x_583;
wire x_584;
wire x_585;
wire x_586;
wire x_587;
wire x_588;
wire x_589;
wire x_590;
wire x_591;
wire x_592;
wire x_593;
wire x_594;
wire x_595;
wire x_596;
wire x_597;
wire x_598;
wire x_599;
wire x_600;
wire x_601;
wire x_602;
wire x_603;
wire x_604;
wire x_605;
wire x_606;
wire x_607;
wire x_608;
wire x_609;
wire x_610;
wire x_611;
wire x_612;
wire x_613;
wire x_614;
wire x_615;
wire x_616;
wire x_617;
wire x_618;
wire x_619;
wire x_620;
wire x_621;
wire x_622;
wire x_623;
wire x_624;
wire x_625;
wire x_626;
wire x_627;
wire x_628;
wire x_629;
wire x_630;
wire x_631;
wire x_632;
wire x_633;
wire x_634;
wire x_635;
wire x_636;
wire x_637;
wire x_638;
wire x_639;
wire x_640;
wire x_641;
wire x_642;
wire x_643;
wire x_644;
wire x_645;
wire x_646;
wire x_647;
wire x_648;
wire x_649;
wire x_650;
wire x_651;
wire x_652;
wire x_653;
wire x_654;
wire x_655;
wire x_656;
wire x_657;
wire x_658;
wire x_659;
wire x_660;
wire x_661;
wire x_662;
wire x_663;
wire x_664;
wire x_665;
wire x_666;
wire x_667;
wire x_668;
wire x_669;
wire x_670;
wire x_671;
wire x_672;
wire x_673;
wire x_674;
wire x_675;
wire x_676;
wire x_677;
wire x_678;
wire x_679;
wire x_680;
wire x_681;
wire x_682;
wire x_683;
wire x_684;
wire x_685;
wire x_686;
wire x_687;
wire x_688;
wire x_689;
wire x_690;
wire x_691;
wire x_692;
wire x_693;
wire x_694;
wire x_695;
wire x_696;
wire x_697;
wire x_698;
wire x_699;
wire x_700;
wire x_701;
wire x_702;
wire x_703;
wire x_704;
wire x_705;
wire x_706;
wire x_707;
wire x_708;
wire x_709;
wire x_710;
wire x_711;
wire x_712;
wire x_713;
wire x_714;
wire x_715;
wire x_716;
wire x_717;
wire x_718;
wire x_719;
wire x_720;
wire x_721;
wire x_722;
wire x_723;
wire x_724;
wire x_725;
wire x_726;
wire x_727;
wire x_728;
wire x_729;
wire x_730;
wire x_731;
wire x_732;
wire x_733;
wire x_734;
wire x_735;
wire x_736;
wire x_737;
wire x_738;
wire x_739;
wire x_740;
wire x_741;
wire x_742;
wire x_743;
wire x_744;
wire x_745;
wire x_746;
wire x_747;
wire x_748;
wire x_749;
wire x_750;
wire x_751;
wire x_752;
wire x_753;
wire x_754;
wire x_755;
wire x_756;
wire x_757;
wire x_758;
wire x_759;
wire x_760;
wire x_761;
wire x_762;
wire x_763;
wire x_764;
wire x_765;
wire x_766;
wire x_767;
wire x_768;
wire x_769;
wire x_770;
wire x_771;
wire x_772;
wire x_773;
wire x_774;
wire x_775;
wire x_776;
wire x_777;
wire x_778;
wire x_779;
wire x_780;
wire x_781;
wire x_782;
wire x_783;
wire x_784;
wire x_785;
wire x_786;
wire x_787;
wire x_788;
wire x_789;
wire x_790;
wire x_791;
wire x_792;
wire x_793;
wire x_794;
wire x_795;
wire x_796;
wire x_797;
wire x_798;
wire x_799;
wire x_800;
wire x_801;
wire x_802;
wire x_803;
wire x_804;
wire x_805;
wire x_806;
wire x_807;
wire x_808;
wire x_809;
wire x_810;
wire x_811;
wire x_812;
wire x_813;
wire x_814;
wire x_815;
wire x_816;
wire x_817;
wire x_818;
wire x_819;
wire x_820;
wire x_821;
wire x_822;
wire x_823;
wire x_824;
wire x_825;
wire x_826;
wire x_827;
wire x_828;
wire x_829;
wire x_830;
wire x_831;
wire x_832;
wire x_833;
wire x_834;
wire x_835;
wire x_836;
wire x_837;
wire x_838;
wire x_839;
wire x_840;
wire x_841;
wire x_842;
wire x_843;
wire x_844;
wire x_845;
wire x_846;
wire x_847;
wire x_848;
wire x_849;
wire x_850;
wire x_851;
wire x_852;
wire x_853;
wire x_854;
wire x_855;
wire x_856;
wire x_857;
wire x_858;
wire x_859;
wire x_860;
wire x_861;
wire x_862;
wire x_863;
wire x_864;
wire x_865;
wire x_866;
wire x_867;
wire x_868;
wire x_869;
wire x_870;
wire x_871;
wire x_872;
wire x_873;
wire x_874;
wire x_875;
wire x_876;
wire x_877;
wire x_878;
wire x_879;
wire x_880;
wire x_881;
wire x_882;
wire x_883;
wire x_884;
wire x_885;
wire x_886;
wire x_887;
wire x_888;
wire x_889;
wire x_890;
wire x_891;
wire x_892;
wire x_893;
wire x_894;
wire x_895;
wire x_896;
wire x_897;
wire x_898;
wire x_899;
wire x_900;
wire x_901;
wire x_902;
wire x_903;
wire x_904;
wire x_905;
wire x_906;
wire x_907;
wire x_908;
wire x_909;
wire x_910;
wire x_911;
wire x_912;
wire x_913;
wire x_914;
wire x_915;
wire x_916;
wire x_917;
wire x_918;
wire x_919;
wire x_920;
wire x_921;
wire x_922;
wire x_923;
wire x_924;
wire x_925;
wire x_926;
wire x_927;
wire x_928;
wire x_929;
wire x_930;
wire x_931;
wire x_932;
wire x_933;
wire x_934;
wire x_935;
wire x_936;
wire x_937;
wire x_938;
wire x_939;
wire x_940;
wire x_941;
wire x_942;
wire x_943;
wire x_944;
wire x_945;
wire x_946;
wire x_947;
wire x_948;
wire x_949;
wire x_950;
wire x_951;
wire x_952;
wire x_953;
wire x_954;
wire x_955;
wire x_956;
wire x_957;
wire x_958;
wire x_959;
wire x_960;
wire x_961;
wire x_962;
wire x_963;
wire x_964;
wire x_965;
wire x_966;
wire x_967;
wire x_968;
wire x_969;
wire x_970;
wire x_971;
wire x_972;
wire x_973;
wire x_974;
wire x_975;
wire x_976;
wire x_977;
wire x_978;
wire x_979;
wire x_980;
wire x_981;
wire x_982;
wire x_983;
wire x_984;
wire x_985;
wire x_986;
wire x_987;
wire x_988;
wire x_989;
wire x_990;
wire x_991;
wire x_992;
wire x_993;
wire x_994;
wire x_995;
wire x_996;
wire x_997;
wire x_998;
wire x_999;
wire x_1000;
wire x_1001;
wire x_1002;
wire x_1003;
wire x_1004;
wire x_1005;
wire x_1006;
wire x_1007;
wire x_1008;
wire x_1009;
wire x_1010;
wire x_1011;
wire x_1012;
wire x_1013;
wire x_1014;
wire x_1015;
wire x_1016;
wire x_1017;
wire x_1018;
wire x_1019;
wire x_1020;
wire x_1021;
wire x_1022;
wire x_1023;
wire x_1024;
wire x_1025;
wire x_1026;
wire x_1027;
wire x_1028;
wire x_1029;
wire x_1030;
wire x_1031;
wire x_1032;
wire x_1033;
wire x_1034;
wire x_1035;
wire x_1036;
wire x_1037;
wire x_1038;
wire x_1039;
wire x_1040;
wire x_1041;
wire x_1042;
wire x_1043;
wire x_1044;
wire x_1045;
wire x_1046;
wire x_1047;
wire x_1048;
wire x_1049;
wire x_1050;
wire x_1051;
wire x_1052;
wire x_1053;
wire x_1054;
wire x_1055;
wire x_1056;
wire x_1057;
wire x_1058;
wire x_1059;
wire x_1060;
wire x_1061;
wire x_1062;
wire x_1063;
wire x_1064;
wire x_1065;
wire x_1066;
wire x_1067;
wire x_1068;
wire x_1069;
wire x_1070;
wire x_1071;
wire x_1072;
wire x_1073;
wire x_1074;
wire x_1075;
wire x_1076;
wire x_1077;
wire x_1078;
wire x_1079;
wire x_1080;
wire x_1081;
wire x_1082;
wire x_1083;
wire x_1084;
wire x_1085;
wire x_1086;
wire x_1087;
wire x_1088;
wire x_1089;
wire x_1090;
wire x_1091;
wire x_1092;
wire x_1093;
wire x_1094;
wire x_1095;
wire x_1096;
wire x_1097;
wire x_1098;
wire x_1099;
wire x_1100;
wire x_1101;
wire x_1102;
wire x_1103;
wire x_1104;
wire x_1105;
wire x_1106;
wire x_1107;
wire x_1108;
wire x_1109;
wire x_1110;
wire x_1111;
wire x_1112;
wire x_1113;
wire x_1114;
wire x_1115;
wire x_1116;
wire x_1117;
wire x_1118;
wire x_1119;
wire x_1120;
wire x_1121;
wire x_1122;
wire x_1123;
wire x_1124;
wire x_1125;
wire x_1126;
wire x_1127;
wire x_1128;
wire x_1129;
wire x_1130;
wire x_1131;
wire x_1132;
wire x_1133;
wire x_1134;
wire x_1135;
wire x_1136;
wire x_1137;
wire x_1138;
wire x_1139;
wire x_1140;
wire x_1141;
wire x_1142;
wire x_1143;
wire x_1144;
wire x_1145;
wire x_1146;
wire x_1147;
wire x_1148;
wire x_1149;
wire x_1150;
wire x_1151;
wire x_1152;
wire x_1153;
wire x_1154;
wire x_1155;
wire x_1156;
wire x_1157;
wire x_1158;
wire x_1159;
wire x_1160;
wire x_1161;
wire x_1162;
wire x_1163;
wire x_1164;
wire x_1165;
wire x_1166;
wire x_1167;
wire x_1168;
wire x_1169;
wire x_1170;
wire x_1171;
wire x_1172;
wire x_1173;
wire x_1174;
wire x_1175;
wire x_1176;
wire x_1177;
wire x_1178;
wire x_1179;
wire x_1180;
wire x_1181;
wire x_1182;
wire x_1183;
wire x_1184;
wire x_1185;
wire x_1186;
wire x_1187;
wire x_1188;
wire x_1189;
wire x_1190;
wire x_1191;
wire x_1192;
wire x_1193;
wire x_1194;
wire x_1195;
wire x_1196;
wire x_1197;
wire x_1198;
wire x_1199;
wire x_1200;
wire x_1201;
wire x_1202;
wire x_1203;
wire x_1204;
wire x_1205;
wire x_1206;
wire x_1207;
wire x_1208;
wire x_1209;
wire x_1210;
wire x_1211;
wire x_1212;
wire x_1213;
wire x_1214;
wire x_1215;
wire x_1216;
wire x_1217;
wire x_1218;
wire x_1219;
wire x_1220;
wire x_1221;
wire x_1222;
wire x_1223;
wire x_1224;
wire x_1225;
wire x_1226;
wire x_1227;
wire x_1228;
wire x_1229;
wire x_1230;
wire x_1231;
wire x_1232;
wire x_1233;
wire x_1234;
wire x_1235;
wire x_1236;
wire x_1237;
wire x_1238;
wire x_1239;
wire x_1240;
wire x_1241;
wire x_1242;
wire x_1243;
wire x_1244;
wire x_1245;
wire x_1246;
wire x_1247;
wire x_1248;
wire x_1249;
wire x_1250;
wire x_1251;
wire x_1252;
wire x_1253;
wire x_1254;
wire x_1255;
wire x_1256;
wire x_1257;
wire x_1258;
wire x_1259;
wire x_1260;
wire x_1261;
wire x_1262;
wire x_1263;
wire x_1264;
wire x_1265;
wire x_1266;
wire x_1267;
wire x_1268;
wire x_1269;
wire x_1270;
wire x_1271;
wire x_1272;
wire x_1273;
wire x_1274;
wire x_1275;
wire x_1276;
wire x_1277;
wire x_1278;
wire x_1279;
wire x_1280;
wire x_1281;
wire x_1282;
wire x_1283;
wire x_1284;
wire x_1285;
wire x_1286;
wire x_1287;
wire x_1288;
wire x_1289;
wire x_1290;
wire x_1291;
wire x_1292;
wire x_1293;
wire x_1294;
wire x_1295;
wire x_1296;
wire x_1297;
wire x_1298;
wire x_1299;
wire x_1300;
wire x_1301;
wire x_1302;
wire x_1303;
wire x_1304;
wire x_1305;
wire x_1306;
wire x_1307;
wire x_1308;
wire x_1309;
wire x_1310;
wire x_1311;
wire x_1312;
wire x_1313;
wire x_1314;
wire x_1315;
wire x_1316;
wire x_1317;
wire x_1318;
wire x_1319;
wire x_1320;
wire x_1321;
wire x_1322;
wire x_1323;
wire x_1324;
wire x_1325;
wire x_1326;
wire x_1327;
wire x_1328;
wire x_1329;
wire x_1330;
wire x_1331;
wire x_1332;
wire x_1333;
wire x_1334;
wire x_1335;
wire x_1336;
wire x_1337;
wire x_1338;
wire x_1339;
wire x_1340;
wire x_1341;
wire x_1342;
wire x_1343;
wire x_1344;
wire x_1345;
wire x_1346;
wire x_1347;
wire x_1348;
wire x_1349;
wire x_1350;
wire x_1351;
wire x_1352;
wire x_1353;
wire x_1354;
wire x_1355;
wire x_1356;
wire x_1357;
wire x_1358;
wire x_1359;
wire x_1360;
wire x_1361;
wire x_1362;
wire x_1363;
wire x_1364;
wire x_1365;
wire x_1366;
wire x_1367;
wire x_1368;
wire x_1369;
wire x_1370;
wire x_1371;
wire x_1372;
wire x_1373;
wire x_1374;
wire x_1375;
wire x_1376;
wire x_1377;
wire x_1378;
wire x_1379;
wire x_1380;
wire x_1381;
wire x_1382;
wire x_1383;
wire x_1384;
wire x_1385;
wire x_1386;
wire x_1387;
wire x_1388;
wire x_1389;
wire x_1390;
wire x_1391;
wire x_1392;
wire x_1393;
wire x_1394;
wire x_1395;
wire x_1396;
wire x_1397;
wire x_1398;
wire x_1399;
wire x_1400;
wire x_1401;
wire x_1402;
wire x_1403;
wire x_1404;
wire x_1405;
wire x_1406;
wire x_1407;
wire x_1408;
wire x_1409;
wire x_1410;
wire x_1411;
wire x_1412;
wire x_1413;
wire x_1414;
wire x_1415;
wire x_1416;
wire x_1417;
wire x_1418;
wire x_1419;
wire x_1420;
wire x_1421;
wire x_1422;
wire x_1423;
wire x_1424;
wire x_1425;
wire x_1426;
wire x_1427;
wire x_1428;
wire x_1429;
wire x_1430;
wire x_1431;
wire x_1432;
wire x_1433;
wire x_1434;
wire x_1435;
wire x_1436;
wire x_1437;
wire x_1438;
wire x_1439;
wire x_1440;
wire x_1441;
wire x_1442;
wire x_1443;
wire x_1444;
wire x_1445;
wire x_1446;
wire x_1447;
wire x_1448;
wire x_1449;
wire x_1450;
wire x_1451;
wire x_1452;
wire x_1453;
wire x_1454;
wire x_1455;
wire x_1456;
wire x_1457;
wire x_1458;
wire x_1459;
wire x_1460;
wire x_1461;
wire x_1462;
wire x_1463;
wire x_1464;
wire x_1465;
wire x_1466;
wire x_1467;
wire x_1468;
wire x_1469;
wire x_1470;
wire x_1471;
wire x_1472;
wire x_1473;
wire x_1474;
wire x_1475;
wire x_1476;
wire x_1477;
wire x_1478;
wire x_1479;
wire x_1480;
wire x_1481;
wire x_1482;
wire x_1483;
wire x_1484;
wire x_1485;
wire x_1486;
wire x_1487;
wire x_1488;
wire x_1489;
wire x_1490;
wire x_1491;
wire x_1492;
wire x_1493;
wire x_1494;
wire x_1495;
wire x_1496;
wire x_1497;
wire x_1498;
wire x_1499;
wire x_1500;
wire x_1501;
wire x_1502;
wire x_1503;
wire x_1504;
wire x_1505;
wire x_1506;
wire x_1507;
wire x_1508;
wire x_1509;
wire x_1510;
wire x_1511;
wire x_1512;
wire x_1513;
wire x_1514;
wire x_1515;
wire x_1516;
wire x_1517;
wire x_1518;
wire x_1519;
wire x_1520;
wire x_1521;
wire x_1522;
wire x_1523;
wire x_1524;
wire x_1525;
wire x_1526;
wire x_1527;
wire x_1528;
wire x_1529;
wire x_1530;
wire x_1531;
wire x_1532;
wire x_1533;
wire x_1534;
wire x_1535;
wire x_1536;
wire x_1537;
wire x_1538;
wire x_1539;
wire x_1540;
wire x_1541;
wire x_1542;
wire x_1543;
wire x_1544;
wire x_1545;
wire x_1546;
wire x_1547;
wire x_1548;
wire x_1549;
wire x_1550;
wire x_1551;
wire x_1552;
wire x_1553;
wire x_1554;
wire x_1555;
wire x_1556;
wire x_1557;
wire x_1558;
wire x_1559;
wire x_1560;
wire x_1561;
wire x_1562;
wire x_1563;
wire x_1564;
wire x_1565;
wire x_1566;
wire x_1567;
wire x_1568;
wire x_1569;
wire x_1570;
wire x_1571;
wire x_1572;
wire x_1573;
wire x_1574;
wire x_1575;
wire x_1576;
wire x_1577;
wire x_1578;
wire x_1579;
wire x_1580;
wire x_1581;
wire x_1582;
wire x_1583;
wire x_1584;
wire x_1585;
wire x_1586;
wire x_1587;
wire x_1588;
wire x_1589;
wire x_1590;
wire x_1591;
wire x_1592;
wire x_1593;
wire x_1594;
wire x_1595;
wire x_1596;
wire x_1597;
wire x_1598;
wire x_1599;
wire x_1600;
wire x_1601;
wire x_1602;
wire x_1603;
wire x_1604;
wire x_1605;
wire x_1606;
wire x_1607;
wire x_1608;
wire x_1609;
wire x_1610;
wire x_1611;
wire x_1612;
wire x_1613;
wire x_1614;
wire x_1615;
wire x_1616;
wire x_1617;
wire x_1618;
wire x_1619;
wire x_1620;
wire x_1621;
wire x_1622;
wire x_1623;
wire x_1624;
wire x_1625;
wire x_1626;
wire x_1627;
wire x_1628;
wire x_1629;
wire x_1630;
wire x_1631;
wire x_1632;
wire x_1633;
wire x_1634;
wire x_1635;
wire x_1636;
wire x_1637;
wire x_1638;
wire x_1639;
wire x_1640;
wire x_1641;
wire x_1642;
wire x_1643;
wire x_1644;
wire x_1645;
wire x_1646;
wire x_1647;
wire x_1648;
wire x_1649;
wire x_1650;
wire x_1651;
wire x_1652;
wire x_1653;
wire x_1654;
wire x_1655;
wire x_1656;
wire x_1657;
wire x_1658;
wire x_1659;
wire x_1660;
wire x_1661;
wire x_1662;
wire x_1663;
wire x_1664;
wire x_1665;
wire x_1666;
wire x_1667;
wire x_1668;
wire x_1669;
wire x_1670;
wire x_1671;
wire x_1672;
wire x_1673;
wire x_1674;
wire x_1675;
wire x_1676;
wire x_1677;
wire x_1678;
wire x_1679;
wire x_1680;
wire x_1681;
wire x_1682;
wire x_1683;
wire x_1684;
wire x_1685;
wire x_1686;
wire x_1687;
wire x_1688;
wire x_1689;
wire x_1690;
wire x_1691;
wire x_1692;
wire x_1693;
wire x_1694;
wire x_1695;
wire x_1696;
wire x_1697;
wire x_1698;
wire x_1699;
wire x_1700;
wire x_1701;
wire x_1702;
wire x_1703;
wire x_1704;
wire x_1705;
wire x_1706;
wire x_1707;
wire x_1708;
wire x_1709;
wire x_1710;
wire x_1711;
wire x_1712;
wire x_1713;
wire x_1714;
wire x_1715;
wire x_1716;
wire x_1717;
wire x_1718;
wire x_1719;
wire x_1720;
wire x_1721;
wire x_1722;
wire x_1723;
wire x_1724;
wire x_1725;
wire x_1726;
wire x_1727;
wire x_1728;
wire x_1729;
wire x_1730;
wire x_1731;
wire x_1732;
wire x_1733;
wire x_1734;
wire x_1735;
wire x_1736;
wire x_1737;
wire x_1738;
wire x_1739;
wire x_1740;
wire x_1741;
wire x_1742;
wire x_1743;
wire x_1744;
wire x_1745;
wire x_1746;
wire x_1747;
wire x_1748;
wire x_1749;
wire x_1750;
wire x_1751;
wire x_1752;
wire x_1753;
wire x_1754;
wire x_1755;
wire x_1756;
wire x_1757;
wire x_1758;
wire x_1759;
wire x_1760;
wire x_1761;
wire x_1762;
wire x_1763;
wire x_1764;
wire x_1765;
wire x_1766;
wire x_1767;
wire x_1768;
wire x_1769;
wire x_1770;
wire x_1771;
wire x_1772;
wire x_1773;
wire x_1774;
wire x_1775;
wire x_1776;
wire x_1777;
wire x_1778;
wire x_1779;
wire x_1780;
wire x_1781;
wire x_1782;
wire x_1783;
wire x_1784;
wire x_1785;
wire x_1786;
wire x_1787;
wire x_1788;
wire x_1789;
wire x_1790;
wire x_1791;
wire x_1792;
wire x_1793;
wire x_1794;
wire x_1795;
wire x_1796;
wire x_1797;
wire x_1798;
wire x_1799;
wire x_1800;
wire x_1801;
wire x_1802;
wire x_1803;
wire x_1804;
wire x_1805;
wire x_1806;
wire x_1807;
wire x_1808;
wire x_1809;
wire x_1810;
wire x_1811;
wire x_1812;
wire x_1813;
wire x_1814;
wire x_1815;
wire x_1816;
wire x_1817;
wire x_1818;
wire x_1819;
wire x_1820;
wire x_1821;
wire x_1822;
wire x_1823;
wire x_1824;
wire x_1825;
wire x_1826;
wire x_1827;
wire x_1828;
wire x_1829;
wire x_1830;
wire x_1831;
wire x_1832;
wire x_1833;
wire x_1834;
wire x_1835;
wire x_1836;
wire x_1837;
wire x_1838;
wire x_1839;
wire x_1840;
wire x_1841;
wire x_1842;
wire x_1843;
wire x_1844;
wire x_1845;
wire x_1846;
wire x_1847;
wire x_1848;
wire x_1849;
wire x_1850;
wire x_1851;
wire x_1852;
wire x_1853;
wire x_1854;
wire x_1855;
wire x_1856;
wire x_1857;
wire x_1858;
wire x_1859;
wire x_1860;
wire x_1861;
wire x_1862;
wire x_1863;
wire x_1864;
wire x_1865;
wire x_1866;
wire x_1867;
wire x_1868;
wire x_1869;
wire x_1870;
wire x_1871;
wire x_1872;
wire x_1873;
wire x_1874;
wire x_1875;
wire x_1876;
wire x_1877;
wire x_1878;
wire x_1879;
wire x_1880;
wire x_1881;
wire x_1882;
wire x_1883;
wire x_1884;
wire x_1885;
wire x_1886;
wire x_1887;
wire x_1888;
wire x_1889;
wire x_1890;
wire x_1891;
wire x_1892;
wire x_1893;
wire x_1894;
wire x_1895;
wire x_1896;
wire x_1897;
wire x_1898;
wire x_1899;
wire x_1900;
wire x_1901;
wire x_1902;
wire x_1903;
wire x_1904;
wire x_1905;
wire x_1906;
wire x_1907;
wire x_1908;
wire x_1909;
wire x_1910;
wire x_1911;
wire x_1912;
wire x_1913;
wire x_1914;
wire x_1915;
wire x_1916;
wire x_1917;
wire x_1918;
wire x_1919;
wire x_1920;
wire x_1921;
wire x_1922;
wire x_1923;
wire x_1924;
wire x_1925;
wire x_1926;
wire x_1927;
wire x_1928;
wire x_1929;
wire x_1930;
wire x_1931;
wire x_1932;
wire x_1933;
wire x_1934;
wire x_1935;
wire x_1936;
wire x_1937;
wire x_1938;
wire x_1939;
wire x_1940;
wire x_1941;
wire x_1942;
wire x_1943;
wire x_1944;
wire x_1945;
wire x_1946;
wire x_1947;
wire x_1948;
wire x_1949;
wire x_1950;
wire x_1951;
wire x_1952;
wire x_1953;
wire x_1954;
wire x_1955;
wire x_1956;
wire x_1957;
wire x_1958;
wire x_1959;
wire x_1960;
wire x_1961;
wire x_1962;
wire x_1963;
wire x_1964;
wire x_1965;
wire x_1966;
wire x_1967;
wire x_1968;
wire x_1969;
wire x_1970;
wire x_1971;
wire x_1972;
wire x_1973;
wire x_1974;
wire x_1975;
wire x_1976;
wire x_1977;
wire x_1978;
wire x_1979;
wire x_1980;
wire x_1981;
wire x_1982;
wire x_1983;
wire x_1984;
wire x_1985;
wire x_1986;
wire x_1987;
wire x_1988;
wire x_1989;
wire x_1990;
wire x_1991;
wire x_1992;
wire x_1993;
wire x_1994;
wire x_1995;
wire x_1996;
wire x_1997;
wire x_1998;
wire x_1999;
wire x_2000;
wire x_2001;
wire x_2002;
wire x_2003;
wire x_2004;
wire x_2005;
wire x_2006;
wire x_2007;
wire x_2008;
wire x_2009;
wire x_2010;
wire x_2011;
wire x_2012;
wire x_2013;
wire x_2014;
wire x_2015;
wire x_2016;
wire x_2017;
wire x_2018;
wire x_2019;
wire x_2020;
wire x_2021;
wire x_2022;
wire x_2023;
wire x_2024;
wire x_2025;
wire x_2026;
wire x_2027;
wire x_2028;
wire x_2029;
wire x_2030;
wire x_2031;
wire x_2032;
wire x_2033;
wire x_2034;
wire x_2035;
wire x_2036;
wire x_2037;
wire x_2038;
wire x_2039;
wire x_2040;
wire x_2041;
wire x_2042;
wire x_2043;
wire x_2044;
wire x_2045;
wire x_2046;
wire x_2047;
wire x_2048;
wire x_2049;
wire x_2050;
wire x_2051;
wire x_2052;
wire x_2053;
wire x_2054;
wire x_2055;
wire x_2056;
wire x_2057;
wire x_2058;
wire x_2059;
wire x_2060;
wire x_2061;
wire x_2062;
wire x_2063;
wire x_2064;
wire x_2065;
wire x_2066;
wire x_2067;
wire x_2068;
wire x_2069;
wire x_2070;
wire x_2071;
wire x_2072;
wire x_2073;
wire x_2074;
wire x_2075;
wire x_2076;
wire x_2077;
wire x_2078;
wire x_2079;
wire x_2080;
wire x_2081;
wire x_2082;
wire x_2083;
wire x_2084;
wire x_2085;
wire x_2086;
wire x_2087;
wire x_2088;
wire x_2089;
wire x_2090;
wire x_2091;
wire x_2092;
wire x_2093;
wire x_2094;
wire x_2095;
wire x_2096;
wire x_2097;
wire x_2098;
wire x_2099;
wire x_2100;
wire x_2101;
wire x_2102;
wire x_2103;
wire x_2104;
wire x_2105;
wire x_2106;
wire x_2107;
wire x_2108;
wire x_2109;
wire x_2110;
wire x_2111;
wire x_2112;
wire x_2113;
wire x_2114;
wire x_2115;
wire x_2116;
wire x_2117;
wire x_2118;
wire x_2119;
wire x_2120;
wire x_2121;
wire x_2122;
wire x_2123;
wire x_2124;
wire x_2125;
wire x_2126;
wire x_2127;
wire x_2128;
wire x_2129;
wire x_2130;
wire x_2131;
wire x_2132;
wire x_2133;
wire x_2134;
wire x_2135;
wire x_2136;
wire x_2137;
wire x_2138;
wire x_2139;
wire x_2140;
wire x_2141;
wire x_2142;
wire x_2143;
wire x_2144;
wire x_2145;
wire x_2146;
wire x_2147;
wire x_2148;
wire x_2149;
wire x_2150;
wire x_2151;
wire x_2152;
wire x_2153;
wire x_2154;
wire x_2155;
wire x_2156;
wire x_2157;
wire x_2158;
wire x_2159;
wire x_2160;
wire x_2161;
wire x_2162;
wire x_2163;
wire x_2164;
wire x_2165;
wire x_2166;
wire x_2167;
wire x_2168;
wire x_2169;
wire x_2170;
wire x_2171;
wire x_2172;
wire x_2173;
wire x_2174;
wire x_2175;
wire x_2176;
wire x_2177;
wire x_2178;
wire x_2179;
wire x_2180;
wire x_2181;
wire x_2182;
wire x_2183;
wire x_2184;
wire x_2185;
wire x_2186;
wire x_2187;
wire x_2188;
wire x_2189;
wire x_2190;
wire x_2191;
wire x_2192;
wire x_2193;
wire x_2194;
wire x_2195;
wire x_2196;
wire x_2197;
wire x_2198;
wire x_2199;
wire x_2200;
wire x_2201;
wire x_2202;
wire x_2203;
wire x_2204;
wire x_2205;
wire x_2206;
wire x_2207;
wire x_2208;
wire x_2209;
wire x_2210;
wire x_2211;
wire x_2212;
wire x_2213;
wire x_2214;
wire x_2215;
wire x_2216;
wire x_2217;
wire x_2218;
wire x_2219;
wire x_2220;
wire x_2221;
wire x_2222;
wire x_2223;
wire x_2224;
wire x_2225;
wire x_2226;
wire x_2227;
wire x_2228;
wire x_2229;
wire x_2230;
wire x_2231;
wire x_2232;
wire x_2233;
wire x_2234;
wire x_2235;
wire x_2236;
wire x_2237;
wire x_2238;
wire x_2239;
wire x_2240;
wire x_2241;
wire x_2242;
wire x_2243;
wire x_2244;
wire x_2245;
wire x_2246;
wire x_2247;
wire x_2248;
wire x_2249;
wire x_2250;
wire x_2251;
wire x_2252;
wire x_2253;
wire x_2254;
wire x_2255;
wire x_2256;
wire x_2257;
wire x_2258;
wire x_2259;
wire x_2260;
wire x_2261;
wire x_2262;
wire x_2263;
wire x_2264;
wire x_2265;
wire x_2266;
wire x_2267;
wire x_2268;
wire x_2269;
wire x_2270;
wire x_2271;
wire x_2272;
wire x_2273;
wire x_2274;
wire x_2275;
wire x_2276;
wire x_2277;
wire x_2278;
wire x_2279;
wire x_2280;
wire x_2281;
wire x_2282;
wire x_2283;
wire x_2284;
wire x_2285;
wire x_2286;
wire x_2287;
wire x_2288;
wire x_2289;
wire x_2290;
wire x_2291;
wire x_2292;
wire x_2293;
wire x_2294;
wire x_2295;
wire x_2296;
wire x_2297;
wire x_2298;
wire x_2299;
wire x_2300;
wire x_2301;
wire x_2302;
wire x_2303;
wire x_2304;
wire x_2305;
wire x_2306;
wire x_2307;
wire x_2308;
wire x_2309;
wire x_2310;
wire x_2311;
wire x_2312;
wire x_2313;
wire x_2314;
wire x_2315;
wire x_2316;
wire x_2317;
wire x_2318;
wire x_2319;
wire x_2320;
wire x_2321;
wire x_2322;
wire x_2323;
wire x_2324;
wire x_2325;
wire x_2326;
wire x_2327;
wire x_2328;
wire x_2329;
wire x_2330;
wire x_2331;
wire x_2332;
wire x_2333;
wire x_2334;
wire x_2335;
wire x_2336;
wire x_2337;
wire x_2338;
wire x_2339;
wire x_2340;
wire x_2341;
wire x_2342;
wire x_2343;
wire x_2344;
wire x_2345;
wire x_2346;
wire x_2347;
wire x_2348;
wire x_2349;
wire x_2350;
wire x_2351;
wire x_2352;
wire x_2353;
wire x_2354;
wire x_2355;
wire x_2356;
wire x_2357;
wire x_2358;
wire x_2359;
wire x_2360;
wire x_2361;
wire x_2362;
wire x_2363;
wire x_2364;
wire x_2365;
wire x_2366;
wire x_2367;
wire x_2368;
wire x_2369;
wire x_2370;
wire x_2371;
wire x_2372;
wire x_2373;
wire x_2374;
wire x_2375;
wire x_2376;
wire x_2377;
wire x_2378;
wire x_2379;
wire x_2380;
wire x_2381;
wire x_2382;
wire x_2383;
wire x_2384;
wire x_2385;
wire x_2386;
wire x_2387;
wire x_2388;
wire x_2389;
wire x_2390;
wire x_2391;
wire x_2392;
wire x_2393;
wire x_2394;
wire x_2395;
wire x_2396;
wire x_2397;
wire x_2398;
wire x_2399;
wire x_2400;
wire x_2401;
wire x_2402;
wire x_2403;
wire x_2404;
wire x_2405;
wire x_2406;
wire x_2407;
wire x_2408;
wire x_2409;
wire x_2410;
wire x_2411;
wire x_2412;
wire x_2413;
wire x_2414;
wire x_2415;
wire x_2416;
wire x_2417;
wire x_2418;
wire x_2419;
wire x_2420;
wire x_2421;
wire x_2422;
wire x_2423;
wire x_2424;
wire x_2425;
wire x_2426;
wire x_2427;
wire x_2428;
wire x_2429;
wire x_2430;
wire x_2431;
wire x_2432;
wire x_2433;
wire x_2434;
wire x_2435;
wire x_2436;
wire x_2437;
wire x_2438;
wire x_2439;
wire x_2440;
wire x_2441;
wire x_2442;
wire x_2443;
wire x_2444;
wire x_2445;
wire x_2446;
wire x_2447;
wire x_2448;
wire x_2449;
wire x_2450;
wire x_2451;
wire x_2452;
wire x_2453;
wire x_2454;
wire x_2455;
wire x_2456;
wire x_2457;
wire x_2458;
wire x_2459;
wire x_2460;
wire x_2461;
wire x_2462;
wire x_2463;
wire x_2464;
wire x_2465;
wire x_2466;
wire x_2467;
wire x_2468;
wire x_2469;
wire x_2470;
wire x_2471;
wire x_2472;
wire x_2473;
wire x_2474;
wire x_2475;
wire x_2476;
wire x_2477;
wire x_2478;
wire x_2479;
wire x_2480;
wire x_2481;
wire x_2482;
wire x_2483;
wire x_2484;
wire x_2485;
wire x_2486;
wire x_2487;
wire x_2488;
wire x_2489;
wire x_2490;
wire x_2491;
wire x_2492;
wire x_2493;
wire x_2494;
wire x_2495;
wire x_2496;
wire x_2497;
wire x_2498;
wire x_2499;
wire x_2500;
wire x_2501;
wire x_2502;
wire x_2503;
wire x_2504;
wire x_2505;
wire x_2506;
wire x_2507;
wire x_2508;
wire x_2509;
wire x_2510;
wire x_2511;
wire x_2512;
wire x_2513;
wire x_2514;
wire x_2515;
wire x_2516;
wire x_2517;
wire x_2518;
wire x_2519;
wire x_2520;
wire x_2521;
wire x_2522;
wire x_2523;
wire x_2524;
wire x_2525;
wire x_2526;
wire x_2527;
wire x_2528;
wire x_2529;
wire x_2530;
wire x_2531;
wire x_2532;
wire x_2533;
wire x_2534;
wire x_2535;
wire x_2536;
wire x_2537;
wire x_2538;
wire x_2539;
wire x_2540;
wire x_2541;
wire x_2542;
wire x_2543;
wire x_2544;
wire x_2545;
wire x_2546;
wire x_2547;
wire x_2548;
wire x_2549;
wire x_2550;
wire x_2551;
wire x_2552;
wire x_2553;
wire x_2554;
wire x_2555;
wire x_2556;
wire x_2557;
wire x_2558;
wire x_2559;
wire x_2560;
wire x_2561;
wire x_2562;
wire x_2563;
wire x_2564;
wire x_2565;
wire x_2566;
wire x_2567;
wire x_2568;
wire x_2569;
wire x_2570;
wire x_2571;
wire x_2572;
wire x_2573;
wire x_2574;
wire x_2575;
wire x_2576;
wire x_2577;
wire x_2578;
wire x_2579;
wire x_2580;
wire x_2581;
wire x_2582;
wire x_2583;
wire x_2584;
wire x_2585;
wire x_2586;
wire x_2587;
wire x_2588;
wire x_2589;
wire x_2590;
wire x_2591;
wire x_2592;
wire x_2593;
wire x_2594;
wire x_2595;
wire x_2596;
wire x_2597;
wire x_2598;
wire x_2599;
wire x_2600;
wire x_2601;
wire x_2602;
wire x_2603;
wire x_2604;
wire x_2605;
wire x_2606;
wire x_2607;
wire x_2608;
wire x_2609;
wire x_2610;
wire x_2611;
wire x_2612;
wire x_2613;
wire x_2614;
wire x_2615;
wire x_2616;
wire x_2617;
wire x_2618;
wire x_2619;
wire x_2620;
wire x_2621;
wire x_2622;
wire x_2623;
wire x_2624;
wire x_2625;
wire x_2626;
wire x_2627;
wire x_2628;
wire x_2629;
wire x_2630;
wire x_2631;
wire x_2632;
wire x_2633;
wire x_2634;
wire x_2635;
wire x_2636;
wire x_2637;
wire x_2638;
wire x_2639;
wire x_2640;
wire x_2641;
wire x_2642;
wire x_2643;
wire x_2644;
wire x_2645;
wire x_2646;
wire x_2647;
wire x_2648;
wire x_2649;
wire x_2650;
wire x_2651;
wire x_2652;
wire x_2653;
wire x_2654;
wire x_2655;
wire x_2656;
wire x_2657;
wire x_2658;
wire x_2659;
wire x_2660;
wire x_2661;
wire x_2662;
wire x_2663;
wire x_2664;
wire x_2665;
wire x_2666;
wire x_2667;
wire x_2668;
wire x_2669;
wire x_2670;
wire x_2671;
wire x_2672;
wire x_2673;
wire x_2674;
wire x_2675;
wire x_2676;
wire x_2677;
wire x_2678;
wire x_2679;
wire x_2680;
wire x_2681;
wire x_2682;
wire x_2683;
wire x_2684;
wire x_2685;
wire x_2686;
wire x_2687;
wire x_2688;
wire x_2689;
wire x_2690;
wire x_2691;
wire x_2692;
wire x_2693;
wire x_2694;
wire x_2695;
wire x_2696;
wire x_2697;
wire x_2698;
wire x_2699;
wire x_2700;
wire x_2701;
wire x_2702;
wire x_2703;
wire x_2704;
wire x_2705;
wire x_2706;
wire x_2707;
wire x_2708;
wire x_2709;
wire x_2710;
wire x_2711;
wire x_2712;
wire x_2713;
wire x_2714;
wire x_2715;
wire x_2716;
wire x_2717;
wire x_2718;
wire x_2719;
wire x_2720;
wire x_2721;
wire x_2722;
wire x_2723;
wire x_2724;
wire x_2725;
wire x_2726;
wire x_2727;
wire x_2728;
wire x_2729;
wire x_2730;
wire x_2731;
wire x_2732;
wire x_2733;
wire x_2734;
wire x_2735;
wire x_2736;
wire x_2737;
wire x_2738;
wire x_2739;
wire x_2740;
wire x_2741;
wire x_2742;
wire x_2743;
wire x_2744;
wire x_2745;
wire x_2746;
wire x_2747;
wire x_2748;
wire x_2749;
wire x_2750;
wire x_2751;
wire x_2752;
wire x_2753;
wire x_2754;
wire x_2755;
wire x_2756;
wire x_2757;
wire x_2758;
wire x_2759;
wire x_2760;
wire x_2761;
wire x_2762;
wire x_2763;
wire x_2764;
wire x_2765;
wire x_2766;
wire x_2767;
wire x_2768;
wire x_2769;
wire x_2770;
wire x_2771;
wire x_2772;
wire x_2773;
wire x_2774;
wire x_2775;
wire x_2776;
wire x_2777;
wire x_2778;
wire x_2779;
wire x_2780;
wire x_2781;
wire x_2782;
wire x_2783;
wire x_2784;
wire x_2785;
wire x_2786;
wire x_2787;
wire x_2788;
wire x_2789;
wire x_2790;
wire x_2791;
wire x_2792;
wire x_2793;
wire x_2794;
wire x_2795;
wire x_2796;
wire x_2797;
wire x_2798;
wire x_2799;
wire x_2800;
wire x_2801;
wire x_2802;
wire x_2803;
wire x_2804;
wire x_2805;
wire x_2806;
wire x_2807;
wire x_2808;
wire x_2809;
wire x_2810;
wire x_2811;
wire x_2812;
wire x_2813;
wire x_2814;
wire x_2815;
wire x_2816;
wire x_2817;
wire x_2818;
wire x_2819;
wire x_2820;
wire x_2821;
wire x_2822;
wire x_2823;
wire x_2824;
wire x_2825;
wire x_2826;
wire x_2827;
wire x_2828;
wire x_2829;
wire x_2830;
wire x_2831;
wire x_2832;
wire x_2833;
wire x_2834;
wire x_2835;
wire x_2836;
wire x_2837;
wire x_2838;
wire x_2839;
wire x_2840;
wire x_2841;
wire x_2842;
wire x_2843;
wire x_2844;
wire x_2845;
wire x_2846;
wire x_2847;
wire x_2848;
wire x_2849;
wire x_2850;
wire x_2851;
wire x_2852;
wire x_2853;
wire x_2854;
wire x_2855;
wire x_2856;
wire x_2857;
wire x_2858;
wire x_2859;
wire x_2860;
wire x_2861;
wire x_2862;
wire x_2863;
wire x_2864;
wire x_2865;
wire x_2866;
wire x_2867;
wire x_2868;
wire x_2869;
wire x_2870;
wire x_2871;
wire x_2872;
wire x_2873;
wire x_2874;
wire x_2875;
wire x_2876;
wire x_2877;
wire x_2878;
wire x_2879;
wire x_2880;
wire x_2881;
wire x_2882;
wire x_2883;
wire x_2884;
wire x_2885;
wire x_2886;
wire x_2887;
wire x_2888;
wire x_2889;
wire x_2890;
wire x_2891;
wire x_2892;
wire x_2893;
wire x_2894;
wire x_2895;
wire x_2896;
wire x_2897;
wire x_2898;
wire x_2899;
wire x_2900;
wire x_2901;
wire x_2902;
wire x_2903;
wire x_2904;
wire x_2905;
wire x_2906;
wire x_2907;
wire x_2908;
wire x_2909;
wire x_2910;
wire x_2911;
wire x_2912;
wire x_2913;
wire x_2914;
wire x_2915;
wire x_2916;
wire x_2917;
wire x_2918;
wire x_2919;
wire x_2920;
wire x_2921;
wire x_2922;
wire x_2923;
wire x_2924;
wire x_2925;
wire x_2926;
wire x_2927;
wire x_2928;
wire x_2929;
wire x_2930;
wire x_2931;
wire x_2932;
wire x_2933;
wire x_2934;
wire x_2935;
wire x_2936;
wire x_2937;
wire x_2938;
wire x_2939;
wire x_2940;
wire x_2941;
wire x_2942;
wire x_2943;
wire x_2944;
wire x_2945;
wire x_2946;
wire x_2947;
wire x_2948;
wire x_2949;
wire x_2950;
wire x_2951;
wire x_2952;
wire x_2953;
wire x_2954;
wire x_2955;
wire x_2956;
wire x_2957;
wire x_2958;
wire x_2959;
wire x_2960;
wire x_2961;
wire x_2962;
wire x_2963;
wire x_2964;
wire x_2965;
wire x_2966;
wire x_2967;
wire x_2968;
wire x_2969;
wire x_2970;
wire x_2971;
wire x_2972;
wire x_2973;
wire x_2974;
wire x_2975;
wire x_2976;
wire x_2977;
wire x_2978;
wire x_2979;
wire x_2980;
wire x_2981;
wire x_2982;
wire x_2983;
wire x_2984;
wire x_2985;
wire x_2986;
wire x_2987;
wire x_2988;
wire x_2989;
wire x_2990;
wire x_2991;
wire x_2992;
wire x_2993;
wire x_2994;
wire x_2995;
wire x_2996;
wire x_2997;
wire x_2998;
wire x_2999;
wire x_3000;
wire x_3001;
wire x_3002;
wire x_3003;
wire x_3004;
wire x_3005;
wire x_3006;
wire x_3007;
wire x_3008;
wire x_3009;
wire x_3010;
wire x_3011;
wire x_3012;
wire x_3013;
wire x_3014;
wire x_3015;
wire x_3016;
wire x_3017;
wire x_3018;
wire x_3019;
wire x_3020;
wire x_3021;
wire x_3022;
wire x_3023;
wire x_3024;
wire x_3025;
wire x_3026;
wire x_3027;
wire x_3028;
wire x_3029;
wire x_3030;
wire x_3031;
wire x_3032;
wire x_3033;
wire x_3034;
wire x_3035;
wire x_3036;
wire x_3037;
wire x_3038;
wire x_3039;
wire x_3040;
wire x_3041;
wire x_3042;
wire x_3043;
wire x_3044;
wire x_3045;
wire x_3046;
wire x_3047;
wire x_3048;
wire x_3049;
wire x_3050;
wire x_3051;
wire x_3052;
wire x_3053;
wire x_3054;
wire x_3055;
wire x_3056;
wire x_3057;
wire x_3058;
wire x_3059;
wire x_3060;
wire x_3061;
wire x_3062;
wire x_3063;
wire x_3064;
wire x_3065;
wire x_3066;
wire x_3067;
wire x_3068;
wire x_3069;
wire x_3070;
wire x_3071;
wire x_3072;
wire x_3073;
wire x_3074;
wire x_3075;
wire x_3076;
wire x_3077;
wire x_3078;
wire x_3079;
wire x_3080;
wire x_3081;
wire x_3082;
wire x_3083;
wire x_3084;
wire x_3085;
wire x_3086;
wire x_3087;
wire x_3088;
wire x_3089;
wire x_3090;
wire x_3091;
wire x_3092;
wire x_3093;
wire x_3094;
wire x_3095;
wire x_3096;
wire x_3097;
wire x_3098;
wire x_3099;
wire x_3100;
wire x_3101;
wire x_3102;
wire x_3103;
wire x_3104;
wire x_3105;
wire x_3106;
wire x_3107;
wire x_3108;
wire x_3109;
wire x_3110;
wire x_3111;
wire x_3112;
wire x_3113;
wire x_3114;
wire x_3115;
wire x_3116;
wire x_3117;
wire x_3118;
wire x_3119;
wire x_3120;
wire x_3121;
wire x_3122;
wire x_3123;
wire x_3124;
wire x_3125;
wire x_3126;
wire x_3127;
wire x_3128;
wire x_3129;
wire x_3130;
wire x_3131;
wire x_3132;
wire x_3133;
wire x_3134;
wire x_3135;
wire x_3136;
wire x_3137;
wire x_3138;
wire x_3139;
wire x_3140;
wire x_3141;
wire x_3142;
wire x_3143;
wire x_3144;
wire x_3145;
wire x_3146;
wire x_3147;
wire x_3148;
wire x_3149;
wire x_3150;
wire x_3151;
wire x_3152;
wire x_3153;
wire x_3154;
wire x_3155;
wire x_3156;
wire x_3157;
wire x_3158;
wire x_3159;
wire x_3160;
wire x_3161;
wire x_3162;
wire x_3163;
wire x_3164;
wire x_3165;
wire x_3166;
wire x_3167;
wire x_3168;
wire x_3169;
wire x_3170;
wire x_3171;
wire x_3172;
wire x_3173;
wire x_3174;
wire x_3175;
wire x_3176;
wire x_3177;
wire x_3178;
wire x_3179;
wire x_3180;
wire x_3181;
wire x_3182;
wire x_3183;
wire x_3184;
wire x_3185;
wire x_3186;
wire x_3187;
wire x_3188;
wire x_3189;
wire x_3190;
wire x_3191;
wire x_3192;
wire x_3193;
wire x_3194;
wire x_3195;
wire x_3196;
wire x_3197;
wire x_3198;
wire x_3199;
wire x_3200;
wire x_3201;
wire x_3202;
wire x_3203;
wire x_3204;
wire x_3205;
wire x_3206;
wire x_3207;
wire x_3208;
wire x_3209;
wire x_3210;
wire x_3211;
wire x_3212;
wire x_3213;
wire x_3214;
wire x_3215;
wire x_3216;
wire x_3217;
wire x_3218;
wire x_3219;
wire x_3220;
wire x_3221;
wire x_3222;
wire x_3223;
wire x_3224;
wire x_3225;
wire x_3226;
wire x_3227;
wire x_3228;
wire x_3229;
wire x_3230;
wire x_3231;
wire x_3232;
wire x_3233;
wire x_3234;
wire x_3235;
wire x_3236;
wire x_3237;
wire x_3238;
wire x_3239;
wire x_3240;
wire x_3241;
wire x_3242;
wire x_3243;
wire x_3244;
wire x_3245;
wire x_3246;
wire x_3247;
wire x_3248;
wire x_3249;
wire x_3250;
wire x_3251;
wire x_3252;
wire x_3253;
wire x_3254;
wire x_3255;
wire x_3256;
wire x_3257;
wire x_3258;
wire x_3259;
wire x_3260;
wire x_3261;
wire x_3262;
wire x_3263;
wire x_3264;
wire x_3265;
wire x_3266;
wire x_3267;
wire x_3268;
wire x_3269;
wire x_3270;
wire x_3271;
wire x_3272;
wire x_3273;
wire x_3274;
wire x_3275;
wire x_3276;
wire x_3277;
wire x_3278;
wire x_3279;
wire x_3280;
wire x_3281;
wire x_3282;
wire x_3283;
wire x_3284;
wire x_3285;
wire x_3286;
wire x_3287;
wire x_3288;
wire x_3289;
wire x_3290;
wire x_3291;
wire x_3292;
wire x_3293;
wire x_3294;
wire x_3295;
wire x_3296;
wire x_3297;
wire x_3298;
wire x_3299;
wire x_3300;
wire x_3301;
wire x_3302;
wire x_3303;
wire x_3304;
wire x_3305;
wire x_3306;
wire x_3307;
wire x_3308;
wire x_3309;
wire x_3310;
wire x_3311;
wire x_3312;
wire x_3313;
wire x_3314;
wire x_3315;
wire x_3316;
wire x_3317;
wire x_3318;
wire x_3319;
wire x_3320;
wire x_3321;
wire x_3322;
wire x_3323;
wire x_3324;
wire x_3325;
wire x_3326;
wire x_3327;
wire x_3328;
wire x_3329;
wire x_3330;
wire x_3331;
wire x_3332;
wire x_3333;
wire x_3334;
wire x_3335;
wire x_3336;
wire x_3337;
wire x_3338;
wire x_3339;
wire x_3340;
wire x_3341;
wire x_3342;
wire x_3343;
wire x_3344;
wire x_3345;
wire x_3346;
wire x_3347;
wire x_3348;
wire x_3349;
wire x_3350;
wire x_3351;
wire x_3352;
wire x_3353;
wire x_3354;
wire x_3355;
wire x_3356;
wire x_3357;
wire x_3358;
wire x_3359;
wire x_3360;
wire x_3361;
wire x_3362;
wire x_3363;
wire x_3364;
wire x_3365;
wire x_3366;
wire x_3367;
wire x_3368;
wire x_3369;
wire x_3370;
wire x_3371;
wire x_3372;
wire x_3373;
wire x_3374;
wire x_3375;
wire x_3376;
wire x_3377;
wire x_3378;
wire x_3379;
wire x_3380;
wire x_3381;
wire x_3382;
wire x_3383;
wire x_3384;
wire x_3385;
wire x_3386;
wire x_3387;
wire x_3388;
wire x_3389;
wire x_3390;
wire x_3391;
wire x_3392;
wire x_3393;
wire x_3394;
wire x_3395;
wire x_3396;
wire x_3397;
wire x_3398;
wire x_3399;
wire x_3400;
wire x_3401;
wire x_3402;
wire x_3403;
wire x_3404;
wire x_3405;
wire x_3406;
wire x_3407;
wire x_3408;
wire x_3409;
wire x_3410;
wire x_3411;
wire x_3412;
wire x_3413;
wire x_3414;
wire x_3415;
wire x_3416;
wire x_3417;
wire x_3418;
wire x_3419;
wire x_3420;
wire x_3421;
wire x_3422;
wire x_3423;
wire x_3424;
wire x_3425;
wire x_3426;
wire x_3427;
wire x_3428;
wire x_3429;
wire x_3430;
wire x_3431;
wire x_3432;
wire x_3433;
wire x_3434;
wire x_3435;
wire x_3436;
wire x_3437;
wire x_3438;
wire x_3439;
wire x_3440;
wire x_3441;
wire x_3442;
wire x_3443;
wire x_3444;
wire x_3445;
wire x_3446;
wire x_3447;
wire x_3448;
wire x_3449;
wire x_3450;
wire x_3451;
wire x_3452;
wire x_3453;
wire x_3454;
wire x_3455;
wire x_3456;
wire x_3457;
wire x_3458;
wire x_3459;
wire x_3460;
wire x_3461;
wire x_3462;
wire x_3463;
wire x_3464;
wire x_3465;
wire x_3466;
wire x_3467;
wire x_3468;
wire x_3469;
wire x_3470;
wire x_3471;
wire x_3472;
wire x_3473;
wire x_3474;
wire x_3475;
wire x_3476;
wire x_3477;
wire x_3478;
wire x_3479;
wire x_3480;
wire x_3481;
wire x_3482;
wire x_3483;
wire x_3484;
wire x_3485;
wire x_3486;
wire x_3487;
wire x_3488;
wire x_3489;
wire x_3490;
wire x_3491;
wire x_3492;
wire x_3493;
wire x_3494;
wire x_3495;
wire x_3496;
wire x_3497;
wire x_3498;
wire x_3499;
wire x_3500;
wire x_3501;
wire x_3502;
wire x_3503;
wire x_3504;
wire x_3505;
wire x_3506;
wire x_3507;
wire x_3508;
wire x_3509;
wire x_3510;
wire x_3511;
wire x_3512;
wire x_3513;
wire x_3514;
wire x_3515;
wire x_3516;
wire x_3517;
wire x_3518;
wire x_3519;
wire x_3520;
wire x_3521;
wire x_3522;
wire x_3523;
wire x_3524;
wire x_3525;
wire x_3526;
wire x_3527;
wire x_3528;
wire x_3529;
wire x_3530;
wire x_3531;
wire x_3532;
wire x_3533;
wire x_3534;
wire x_3535;
wire x_3536;
wire x_3537;
wire x_3538;
wire x_3539;
wire x_3540;
wire x_3541;
wire x_3542;
wire x_3543;
wire x_3544;
wire x_3545;
wire x_3546;
wire x_3547;
wire x_3548;
wire x_3549;
wire x_3550;
wire x_3551;
wire x_3552;
wire x_3553;
wire x_3554;
wire x_3555;
wire x_3556;
wire x_3557;
wire x_3558;
wire x_3559;
wire x_3560;
wire x_3561;
wire x_3562;
wire x_3563;
wire x_3564;
wire x_3565;
wire x_3566;
wire x_3567;
wire x_3568;
wire x_3569;
wire x_3570;
wire x_3571;
wire x_3572;
wire x_3573;
wire x_3574;
wire x_3575;
wire x_3576;
wire x_3577;
wire x_3578;
wire x_3579;
wire x_3580;
wire x_3581;
wire x_3582;
wire x_3583;
wire x_3584;
wire x_3585;
wire x_3586;
wire x_3587;
wire x_3588;
wire x_3589;
wire x_3590;
wire x_3591;
wire x_3592;
wire x_3593;
wire x_3594;
wire x_3595;
wire x_3596;
wire x_3597;
wire x_3598;
wire x_3599;
wire x_3600;
wire x_3601;
wire x_3602;
wire x_3603;
wire x_3604;
wire x_3605;
wire x_3606;
wire x_3607;
wire x_3608;
wire x_3609;
wire x_3610;
wire x_3611;
wire x_3612;
wire x_3613;
wire x_3614;
wire x_3615;
wire x_3616;
wire x_3617;
wire x_3618;
wire x_3619;
wire x_3620;
wire x_3621;
wire x_3622;
wire x_3623;
wire x_3624;
wire x_3625;
wire x_3626;
wire x_3627;
wire x_3628;
wire x_3629;
wire x_3630;
wire x_3631;
wire x_3632;
wire x_3633;
wire x_3634;
wire x_3635;
wire x_3636;
wire x_3637;
wire x_3638;
wire x_3639;
wire x_3640;
wire x_3641;
wire x_3642;
wire x_3643;
wire x_3644;
wire x_3645;
wire x_3646;
wire x_3647;
wire x_3648;
wire x_3649;
wire x_3650;
wire x_3651;
wire x_3652;
wire x_3653;
wire x_3654;
wire x_3655;
wire x_3656;
wire x_3657;
wire x_3658;
wire x_3659;
wire x_3660;
wire x_3661;
wire x_3662;
wire x_3663;
wire x_3664;
wire x_3665;
wire x_3666;
wire x_3667;
wire x_3668;
wire x_3669;
wire x_3670;
wire x_3671;
wire x_3672;
wire x_3673;
wire x_3674;
wire x_3675;
wire x_3676;
wire x_3677;
wire x_3678;
wire x_3679;
wire x_3680;
wire x_3681;
wire x_3682;
wire x_3683;
wire x_3684;
wire x_3685;
wire x_3686;
wire x_3687;
wire x_3688;
wire x_3689;
wire x_3690;
wire x_3691;
wire x_3692;
wire x_3693;
wire x_3694;
wire x_3695;
wire x_3696;
wire x_3697;
wire x_3698;
wire x_3699;
wire x_3700;
wire x_3701;
wire x_3702;
wire x_3703;
wire x_3704;
wire x_3705;
wire x_3706;
wire x_3707;
wire x_3708;
wire x_3709;
wire x_3710;
wire x_3711;
wire x_3712;
wire x_3713;
wire x_3714;
wire x_3715;
wire x_3716;
wire x_3717;
wire x_3718;
wire x_3719;
wire x_3720;
wire x_3721;
wire x_3722;
wire x_3723;
wire x_3724;
wire x_3725;
wire x_3726;
wire x_3727;
wire x_3728;
wire x_3729;
wire x_3730;
wire x_3731;
wire x_3732;
wire x_3733;
wire x_3734;
wire x_3735;
wire x_3736;
wire x_3737;
wire x_3738;
wire x_3739;
wire x_3740;
wire x_3741;
wire x_3742;
wire x_3743;
wire x_3744;
wire x_3745;
wire x_3746;
wire x_3747;
wire x_3748;
wire x_3749;
wire x_3750;
wire x_3751;
wire x_3752;
wire x_3753;
wire x_3754;
wire x_3755;
wire x_3756;
wire x_3757;
wire x_3758;
wire x_3759;
wire x_3760;
wire x_3761;
wire x_3762;
wire x_3763;
wire x_3764;
wire x_3765;
wire x_3766;
wire x_3767;
wire x_3768;
wire x_3769;
wire x_3770;
wire x_3771;
wire x_3772;
wire x_3773;
wire x_3774;
wire x_3775;
wire x_3776;
wire x_3777;
wire x_3778;
wire x_3779;
wire x_3780;
wire x_3781;
wire x_3782;
wire x_3783;
wire x_3784;
wire x_3785;
wire x_3786;
wire x_3787;
wire x_3788;
wire x_3789;
wire x_3790;
wire x_3791;
wire x_3792;
wire x_3793;
wire x_3794;
wire x_3795;
wire x_3796;
wire x_3797;
wire x_3798;
wire x_3799;
wire x_3800;
wire x_3801;
wire x_3802;
wire x_3803;
wire x_3804;
wire x_3805;
wire x_3806;
wire x_3807;
wire x_3808;
wire x_3809;
wire x_3810;
wire x_3811;
wire x_3812;
wire x_3813;
wire x_3814;
wire x_3815;
wire x_3816;
wire x_3817;
wire x_3818;
wire x_3819;
wire x_3820;
wire x_3821;
wire x_3822;
wire x_3823;
wire x_3824;
wire x_3825;
wire x_3826;
wire x_3827;
wire x_3828;
wire x_3829;
wire x_3830;
wire x_3831;
wire x_3832;
wire x_3833;
wire x_3834;
wire x_3835;
wire x_3836;
wire x_3837;
wire x_3838;
wire x_3839;
wire x_3840;
wire x_3841;
wire x_3842;
wire x_3843;
wire x_3844;
wire x_3845;
wire x_3846;
wire x_3847;
wire x_3848;
wire x_3849;
wire x_3850;
wire x_3851;
wire x_3852;
wire x_3853;
wire x_3854;
wire x_3855;
wire x_3856;
wire x_3857;
wire x_3858;
wire x_3859;
wire x_3860;
wire x_3861;
wire x_3862;
wire x_3863;
wire x_3864;
wire x_3865;
wire x_3866;
wire x_3867;
wire x_3868;
wire x_3869;
wire x_3870;
wire x_3871;
wire x_3872;
wire x_3873;
wire x_3874;
wire x_3875;
wire x_3876;
wire x_3877;
wire x_3878;
wire x_3879;
wire x_3880;
wire x_3881;
wire x_3882;
wire x_3883;
wire x_3884;
wire x_3885;
wire x_3886;
wire x_3887;
wire x_3888;
wire x_3889;
wire x_3890;
wire x_3891;
wire x_3892;
wire x_3893;
wire x_3894;
wire x_3895;
wire x_3896;
wire x_3897;
wire x_3898;
wire x_3899;
wire x_3900;
wire x_3901;
wire x_3902;
wire x_3903;
wire x_3904;
wire x_3905;
wire x_3906;
wire x_3907;
wire x_3908;
wire x_3909;
wire x_3910;
wire x_3911;
wire x_3912;
wire x_3913;
wire x_3914;
wire x_3915;
wire x_3916;
wire x_3917;
wire x_3918;
wire x_3919;
wire x_3920;
wire x_3921;
wire x_3922;
wire x_3923;
wire x_3924;
wire x_3925;
wire x_3926;
wire x_3927;
wire x_3928;
wire x_3929;
wire x_3930;
wire x_3931;
wire x_3932;
wire x_3933;
wire x_3934;
wire x_3935;
wire x_3936;
wire x_3937;
wire x_3938;
wire x_3939;
wire x_3940;
wire x_3941;
wire x_3942;
wire x_3943;
wire x_3944;
wire x_3945;
wire x_3946;
wire x_3947;
wire x_3948;
wire x_3949;
wire x_3950;
wire x_3951;
wire x_3952;
wire x_3953;
wire x_3954;
wire x_3955;
wire x_3956;
wire x_3957;
wire x_3958;
wire x_3959;
wire x_3960;
wire x_3961;
wire x_3962;
wire x_3963;
wire x_3964;
wire x_3965;
wire x_3966;
wire x_3967;
wire x_3968;
wire x_3969;
wire x_3970;
wire x_3971;
wire x_3972;
wire x_3973;
wire x_3974;
wire x_3975;
wire x_3976;
wire x_3977;
wire x_3978;
wire x_3979;
wire x_3980;
wire x_3981;
wire x_3982;
wire x_3983;
wire x_3984;
wire x_3985;
wire x_3986;
wire x_3987;
wire x_3988;
wire x_3989;
wire x_3990;
wire x_3991;
wire x_3992;
wire x_3993;
wire x_3994;
wire x_3995;
wire x_3996;
wire x_3997;
wire x_3998;
wire x_3999;
wire x_4000;
wire x_4001;
wire x_4002;
wire x_4003;
wire x_4004;
wire x_4005;
wire x_4006;
wire x_4007;
wire x_4008;
wire x_4009;
wire x_4010;
wire x_4011;
wire x_4012;
wire x_4013;
wire x_4014;
wire x_4015;
wire x_4016;
wire x_4017;
wire x_4018;
wire x_4019;
wire x_4020;
wire x_4021;
wire x_4022;
wire x_4023;
wire x_4024;
wire x_4025;
wire x_4026;
wire x_4027;
wire x_4028;
wire x_4029;
wire x_4030;
wire x_4031;
wire x_4032;
wire x_4033;
wire x_4034;
wire x_4035;
wire x_4036;
wire x_4037;
wire x_4038;
wire x_4039;
wire x_4040;
wire x_4041;
wire x_4042;
wire x_4043;
wire x_4044;
wire x_4045;
wire x_4046;
wire x_4047;
wire x_4048;
wire x_4049;
wire x_4050;
wire x_4051;
wire x_4052;
wire x_4053;
wire x_4054;
wire x_4055;
wire x_4056;
wire x_4057;
wire x_4058;
wire x_4059;
wire x_4060;
wire x_4061;
wire x_4062;
wire x_4063;
wire x_4064;
wire x_4065;
wire x_4066;
wire x_4067;
wire x_4068;
wire x_4069;
wire x_4070;
wire x_4071;
wire x_4072;
wire x_4073;
wire x_4074;
wire x_4075;
wire x_4076;
wire x_4077;
wire x_4078;
wire x_4079;
wire x_4080;
wire x_4081;
wire x_4082;
wire x_4083;
wire x_4084;
wire x_4085;
wire x_4086;
wire x_4087;
wire x_4088;
wire x_4089;
wire x_4090;
wire x_4091;
wire x_4092;
wire x_4093;
wire x_4094;
wire x_4095;
wire x_4096;
wire x_4097;
wire x_4098;
wire x_4099;
wire x_4100;
wire x_4101;
wire x_4102;
wire x_4103;
wire x_4104;
wire x_4105;
wire x_4106;
wire x_4107;
wire x_4108;
wire x_4109;
wire x_4110;
wire x_4111;
wire x_4112;
wire x_4113;
wire x_4114;
wire x_4115;
wire x_4116;
wire x_4117;
wire x_4118;
wire x_4119;
wire x_4120;
wire x_4121;
wire x_4122;
wire x_4123;
wire x_4124;
wire x_4125;
wire x_4126;
wire x_4127;
wire x_4128;
wire x_4129;
wire x_4130;
wire x_4131;
wire x_4132;
wire x_4133;
wire x_4134;
wire x_4135;
wire x_4136;
wire x_4137;
wire x_4138;
wire x_4139;
wire x_4140;
wire x_4141;
wire x_4142;
wire x_4143;
wire x_4144;
wire x_4145;
wire x_4146;
wire x_4147;
wire x_4148;
wire x_4149;
wire x_4150;
wire x_4151;
wire x_4152;
wire x_4153;
wire x_4154;
wire x_4155;
wire x_4156;
wire x_4157;
wire x_4158;
wire x_4159;
wire x_4160;
wire x_4161;
wire x_4162;
wire x_4163;
wire x_4164;
wire x_4165;
wire x_4166;
wire x_4167;
wire x_4168;
wire x_4169;
wire x_4170;
wire x_4171;
wire x_4172;
wire x_4173;
wire x_4174;
wire x_4175;
wire x_4176;
wire x_4177;
wire x_4178;
wire x_4179;
wire x_4180;
wire x_4181;
wire x_4182;
wire x_4183;
wire x_4184;
wire x_4185;
wire x_4186;
wire x_4187;
wire x_4188;
wire x_4189;
wire x_4190;
wire x_4191;
wire x_4192;
wire x_4193;
wire x_4194;
wire x_4195;
wire x_4196;
wire x_4197;
wire x_4198;
wire x_4199;
wire x_4200;
wire x_4201;
wire x_4202;
wire x_4203;
wire x_4204;
wire x_4205;
wire x_4206;
wire x_4207;
wire x_4208;
wire x_4209;
wire x_4210;
wire x_4211;
wire x_4212;
wire x_4213;
wire x_4214;
wire x_4215;
wire x_4216;
wire x_4217;
wire x_4218;
wire x_4219;
wire x_4220;
wire x_4221;
wire x_4222;
wire x_4223;
wire x_4224;
wire x_4225;
wire x_4226;
wire x_4227;
wire x_4228;
wire x_4229;
wire x_4230;
wire x_4231;
wire x_4232;
wire x_4233;
wire x_4234;
wire x_4235;
wire x_4236;
wire x_4237;
wire x_4238;
wire x_4239;
wire x_4240;
wire x_4241;
wire x_4242;
wire x_4243;
wire x_4244;
wire x_4245;
wire x_4246;
wire x_4247;
wire x_4248;
wire x_4249;
wire x_4250;
wire x_4251;
wire x_4252;
wire x_4253;
wire x_4254;
wire x_4255;
wire x_4256;
wire x_4257;
wire x_4258;
wire x_4259;
wire x_4260;
wire x_4261;
wire x_4262;
wire x_4263;
wire x_4264;
wire x_4265;
wire x_4266;
wire x_4267;
wire x_4268;
wire x_4269;
wire x_4270;
wire x_4271;
wire x_4272;
wire x_4273;
wire x_4274;
wire x_4275;
wire x_4276;
wire x_4277;
wire x_4278;
wire x_4279;
wire x_4280;
wire x_4281;
wire x_4282;
wire x_4283;
wire x_4284;
wire x_4285;
wire x_4286;
wire x_4287;
wire x_4288;
wire x_4289;
wire x_4290;
wire x_4291;
wire x_4292;
wire x_4293;
wire x_4294;
wire x_4295;
wire x_4296;
wire x_4297;
wire x_4298;
wire x_4299;
wire x_4300;
wire x_4301;
wire x_4302;
wire x_4303;
wire x_4304;
wire x_4305;
wire x_4306;
wire x_4307;
wire x_4308;
wire x_4309;
wire x_4310;
wire x_4311;
wire x_4312;
wire x_4313;
wire x_4314;
wire x_4315;
wire x_4316;
wire x_4317;
wire x_4318;
wire x_4319;
wire x_4320;
wire x_4321;
wire x_4322;
wire x_4323;
wire x_4324;
wire x_4325;
wire x_4326;
wire x_4327;
wire x_4328;
wire x_4329;
wire x_4330;
wire x_4331;
wire x_4332;
wire x_4333;
wire x_4334;
wire x_4335;
wire x_4336;
wire x_4337;
wire x_4338;
wire x_4339;
wire x_4340;
wire x_4341;
wire x_4342;
wire x_4343;
wire x_4344;
wire x_4345;
wire x_4346;
wire x_4347;
wire x_4348;
wire x_4349;
wire x_4350;
wire x_4351;
wire x_4352;
wire x_4353;
wire x_4354;
wire x_4355;
wire x_4356;
wire x_4357;
wire x_4358;
wire x_4359;
wire x_4360;
wire x_4361;
wire x_4362;
wire x_4363;
wire x_4364;
wire x_4365;
wire x_4366;
wire x_4367;
wire x_4368;
wire x_4369;
wire x_4370;
wire x_4371;
wire x_4372;
wire x_4373;
wire x_4374;
wire x_4375;
wire x_4376;
wire x_4377;
wire x_4378;
wire x_4379;
wire x_4380;
wire x_4381;
wire x_4382;
wire x_4383;
wire x_4384;
wire x_4385;
wire x_4386;
wire x_4387;
wire x_4388;
wire x_4389;
wire x_4390;
wire x_4391;
wire x_4392;
wire x_4393;
wire x_4394;
wire x_4395;
wire x_4396;
wire x_4397;
wire x_4398;
wire x_4399;
wire x_4400;
wire x_4401;
wire x_4402;
wire x_4403;
wire x_4404;
wire x_4405;
wire x_4406;
wire x_4407;
wire x_4408;
wire x_4409;
wire x_4410;
wire x_4411;
wire x_4412;
wire x_4413;
wire x_4414;
wire x_4415;
wire x_4416;
wire x_4417;
wire x_4418;
wire x_4419;
wire x_4420;
wire x_4421;
wire x_4422;
wire x_4423;
wire x_4424;
wire x_4425;
wire x_4426;
wire x_4427;
wire x_4428;
wire x_4429;
wire x_4430;
wire x_4431;
wire x_4432;
wire x_4433;
wire x_4434;
wire x_4435;
wire x_4436;
wire x_4437;
wire x_4438;
wire x_4439;
wire x_4440;
wire x_4441;
wire x_4442;
wire x_4443;
wire x_4444;
wire x_4445;
wire x_4446;
wire x_4447;
wire x_4448;
wire x_4449;
wire x_4450;
wire x_4451;
wire x_4452;
wire x_4453;
wire x_4454;
wire x_4455;
wire x_4456;
wire x_4457;
wire x_4458;
wire x_4459;
wire x_4460;
wire x_4461;
wire x_4462;
wire x_4463;
wire x_4464;
wire x_4465;
wire x_4466;
wire x_4467;
wire x_4468;
wire x_4469;
wire x_4470;
wire x_4471;
wire x_4472;
wire x_4473;
wire x_4474;
wire x_4475;
wire x_4476;
wire x_4477;
wire x_4478;
wire x_4479;
wire x_4480;
wire x_4481;
wire x_4482;
wire x_4483;
wire x_4484;
wire x_4485;
wire x_4486;
wire x_4487;
wire x_4488;
wire x_4489;
wire x_4490;
wire x_4491;
wire x_4492;
wire x_4493;
wire x_4494;
wire x_4495;
wire x_4496;
wire x_4497;
wire x_4498;
wire x_4499;
wire x_4500;
wire x_4501;
wire x_4502;
wire x_4503;
wire x_4504;
wire x_4505;
wire x_4506;
wire x_4507;
wire x_4508;
wire x_4509;
wire x_4510;
wire x_4511;
wire x_4512;
wire x_4513;
wire x_4514;
wire x_4515;
wire x_4516;
wire x_4517;
wire x_4518;
wire x_4519;
wire x_4520;
wire x_4521;
wire x_4522;
wire x_4523;
wire x_4524;
wire x_4525;
wire x_4526;
wire x_4527;
wire x_4528;
wire x_4529;
wire x_4530;
wire x_4531;
wire x_4532;
wire x_4533;
wire x_4534;
wire x_4535;
wire x_4536;
wire x_4537;
wire x_4538;
wire x_4539;
wire x_4540;
wire x_4541;
wire x_4542;
wire x_4543;
wire x_4544;
wire x_4545;
wire x_4546;
wire x_4547;
wire x_4548;
wire x_4549;
wire x_4550;
wire x_4551;
wire x_4552;
wire x_4553;
wire x_4554;
wire x_4555;
wire x_4556;
wire x_4557;
wire x_4558;
wire x_4559;
wire x_4560;
wire x_4561;
wire x_4562;
wire x_4563;
wire x_4564;
wire x_4565;
wire x_4566;
wire x_4567;
wire x_4568;
wire x_4569;
wire x_4570;
wire x_4571;
wire x_4572;
wire x_4573;
wire x_4574;
wire x_4575;
wire x_4576;
wire x_4577;
wire x_4578;
wire x_4579;
wire x_4580;
wire x_4581;
wire x_4582;
wire x_4583;
wire x_4584;
wire x_4585;
wire x_4586;
wire x_4587;
wire x_4588;
wire x_4589;
wire x_4590;
wire x_4591;
wire x_4592;
wire x_4593;
wire x_4594;
wire x_4595;
wire x_4596;
wire x_4597;
wire x_4598;
wire x_4599;
wire x_4600;
wire x_4601;
wire x_4602;
wire x_4603;
wire x_4604;
wire x_4605;
wire x_4606;
wire x_4607;
wire x_4608;
wire x_4609;
wire x_4610;
wire x_4611;
wire x_4612;
wire x_4613;
wire x_4614;
wire x_4615;
wire x_4616;
wire x_4617;
wire x_4618;
wire x_4619;
wire x_4620;
wire x_4621;
wire x_4622;
wire x_4623;
wire x_4624;
wire x_4625;
wire x_4626;
wire x_4627;
wire x_4628;
wire x_4629;
wire x_4630;
wire x_4631;
wire x_4632;
wire x_4633;
wire x_4634;
wire x_4635;
wire x_4636;
wire x_4637;
wire x_4638;
wire x_4639;
wire x_4640;
wire x_4641;
wire x_4642;
wire x_4643;
wire x_4644;
wire x_4645;
wire x_4646;
wire x_4647;
wire x_4648;
wire x_4649;
wire x_4650;
wire x_4651;
wire x_4652;
wire x_4653;
wire x_4654;
wire x_4655;
wire x_4656;
wire x_4657;
wire x_4658;
wire x_4659;
wire x_4660;
wire x_4661;
wire x_4662;
wire x_4663;
wire x_4664;
wire x_4665;
wire x_4666;
wire x_4667;
wire x_4668;
wire x_4669;
wire x_4670;
wire x_4671;
wire x_4672;
wire x_4673;
wire x_4674;
wire x_4675;
wire x_4676;
wire x_4677;
wire x_4678;
wire x_4679;
wire x_4680;
wire x_4681;
wire x_4682;
wire x_4683;
wire x_4684;
wire x_4685;
wire x_4686;
wire x_4687;
wire x_4688;
wire x_4689;
wire x_4690;
wire x_4691;
wire x_4692;
wire x_4693;
wire x_4694;
wire x_4695;
wire x_4696;
wire x_4697;
wire x_4698;
wire x_4699;
wire x_4700;
wire x_4701;
wire x_4702;
wire x_4703;
wire x_4704;
wire x_4705;
wire x_4706;
wire x_4707;
wire x_4708;
wire x_4709;
wire x_4710;
wire x_4711;
wire x_4712;
wire x_4713;
wire x_4714;
wire x_4715;
wire x_4716;
wire x_4717;
wire x_4718;
wire x_4719;
wire x_4720;
wire x_4721;
wire x_4722;
wire x_4723;
wire x_4724;
wire x_4725;
wire x_4726;
wire x_4727;
wire x_4728;
wire x_4729;
wire x_4730;
wire x_4731;
wire x_4732;
wire x_4733;
wire x_4734;
wire x_4735;
wire x_4736;
wire x_4737;
wire x_4738;
wire x_4739;
wire x_4740;
wire x_4741;
wire x_4742;
wire x_4743;
wire x_4744;
wire x_4745;
wire x_4746;
wire x_4747;
wire x_4748;
wire x_4749;
wire x_4750;
wire x_4751;
wire x_4752;
wire x_4753;
wire x_4754;
wire x_4755;
wire x_4756;
wire x_4757;
wire x_4758;
wire x_4759;
wire x_4760;
wire x_4761;
wire x_4762;
wire x_4763;
wire x_4764;
wire x_4765;
wire x_4766;
wire x_4767;
wire x_4768;
wire x_4769;
wire x_4770;
wire x_4771;
wire x_4772;
wire x_4773;
wire x_4774;
wire x_4775;
wire x_4776;
wire x_4777;
wire x_4778;
wire x_4779;
wire x_4780;
wire x_4781;
wire x_4782;
wire x_4783;
wire x_4784;
wire x_4785;
wire x_4786;
wire x_4787;
wire x_4788;
wire x_4789;
wire x_4790;
wire x_4791;
wire x_4792;
wire x_4793;
wire x_4794;
wire x_4795;
wire x_4796;
wire x_4797;
wire x_4798;
wire x_4799;
wire x_4800;
wire x_4801;
wire x_4802;
wire x_4803;
wire x_4804;
wire x_4805;
wire x_4806;
wire x_4807;
wire x_4808;
wire x_4809;
wire x_4810;
wire x_4811;
wire x_4812;
wire x_4813;
wire x_4814;
wire x_4815;
wire x_4816;
wire x_4817;
wire x_4818;
wire x_4819;
wire x_4820;
wire x_4821;
wire x_4822;
wire x_4823;
wire x_4824;
wire x_4825;
wire x_4826;
wire x_4827;
wire x_4828;
wire x_4829;
wire x_4830;
wire x_4831;
wire x_4832;
wire x_4833;
wire x_4834;
wire x_4835;
wire x_4836;
wire x_4837;
wire x_4838;
wire x_4839;
wire x_4840;
wire x_4841;
wire x_4842;
wire x_4843;
wire x_4844;
wire x_4845;
wire x_4846;
wire x_4847;
wire x_4848;
wire x_4849;
wire x_4850;
wire x_4851;
wire x_4852;
wire x_4853;
wire x_4854;
wire x_4855;
wire x_4856;
wire x_4857;
wire x_4858;
wire x_4859;
wire x_4860;
wire x_4861;
wire x_4862;
wire x_4863;
wire x_4864;
wire x_4865;
wire x_4866;
wire x_4867;
wire x_4868;
wire x_4869;
wire x_4870;
wire x_4871;
wire x_4872;
wire x_4873;
wire x_4874;
wire x_4875;
wire x_4876;
wire x_4877;
wire x_4878;
wire x_4879;
wire x_4880;
wire x_4881;
wire x_4882;
wire x_4883;
wire x_4884;
wire x_4885;
wire x_4886;
wire x_4887;
wire x_4888;
wire x_4889;
wire x_4890;
wire x_4891;
wire x_4892;
wire x_4893;
wire x_4894;
wire x_4895;
wire x_4896;
wire x_4897;
wire x_4898;
wire x_4899;
wire x_4900;
wire x_4901;
wire x_4902;
wire x_4903;
wire x_4904;
wire x_4905;
wire x_4906;
wire x_4907;
wire x_4908;
wire x_4909;
wire x_4910;
wire x_4911;
wire x_4912;
wire x_4913;
wire x_4914;
wire x_4915;
wire x_4916;
wire x_4917;
wire x_4918;
wire x_4919;
wire x_4920;
wire x_4921;
wire x_4922;
wire x_4923;
wire x_4924;
wire x_4925;
wire x_4926;
wire x_4927;
wire x_4928;
wire x_4929;
wire x_4930;
wire x_4931;
wire x_4932;
wire x_4933;
wire x_4934;
wire x_4935;
wire x_4936;
wire x_4937;
wire x_4938;
wire x_4939;
wire x_4940;
wire x_4941;
wire x_4942;
wire x_4943;
wire x_4944;
wire x_4945;
wire x_4946;
wire x_4947;
wire x_4948;
wire x_4949;
wire x_4950;
wire x_4951;
wire x_4952;
wire x_4953;
wire x_4954;
wire x_4955;
wire x_4956;
wire x_4957;
wire x_4958;
wire x_4959;
wire x_4960;
wire x_4961;
wire x_4962;
wire x_4963;
wire x_4964;
wire x_4965;
wire x_4966;
wire x_4967;
wire x_4968;
wire x_4969;
wire x_4970;
wire x_4971;
wire x_4972;
wire x_4973;
wire x_4974;
wire x_4975;
wire x_4976;
wire x_4977;
wire x_4978;
wire x_4979;
wire x_4980;
wire x_4981;
wire x_4982;
wire x_4983;
wire x_4984;
wire x_4985;
wire x_4986;
wire x_4987;
wire x_4988;
wire x_4989;
wire x_4990;
wire x_4991;
wire x_4992;
wire x_4993;
wire x_4994;
wire x_4995;
wire x_4996;
wire x_4997;
wire x_4998;
wire x_4999;
wire x_5000;
wire x_5001;
wire x_5002;
wire x_5003;
wire x_5004;
wire x_5005;
wire x_5006;
wire x_5007;
wire x_5008;
wire x_5009;
wire x_5010;
wire x_5011;
wire x_5012;
wire x_5013;
wire x_5014;
wire x_5015;
wire x_5016;
wire x_5017;
wire x_5018;
wire x_5019;
wire x_5020;
wire x_5021;
wire x_5022;
wire x_5023;
wire x_5024;
wire x_5025;
wire x_5026;
wire x_5027;
wire x_5028;
wire x_5029;
wire x_5030;
wire x_5031;
wire x_5032;
wire x_5033;
wire x_5034;
wire x_5035;
wire x_5036;
wire x_5037;
wire x_5038;
wire x_5039;
wire x_5040;
wire x_5041;
wire x_5042;
wire x_5043;
wire x_5044;
wire x_5045;
wire x_5046;
wire x_5047;
wire x_5048;
wire x_5049;
wire x_5050;
wire x_5051;
wire x_5052;
wire x_5053;
wire x_5054;
wire x_5055;
wire x_5056;
wire x_5057;
wire x_5058;
wire x_5059;
wire x_5060;
wire x_5061;
wire x_5062;
wire x_5063;
wire x_5064;
wire x_5065;
wire x_5066;
wire x_5067;
wire x_5068;
wire x_5069;
wire x_5070;
wire x_5071;
wire x_5072;
wire x_5073;
wire x_5074;
wire x_5075;
wire x_5076;
wire x_5077;
wire x_5078;
wire x_5079;
wire x_5080;
wire x_5081;
wire x_5082;
wire x_5083;
wire x_5084;
wire x_5085;
wire x_5086;
wire x_5087;
wire x_5088;
wire x_5089;
wire x_5090;
wire x_5091;
wire x_5092;
wire x_5093;
wire x_5094;
wire x_5095;
wire x_5096;
wire x_5097;
wire x_5098;
wire x_5099;
wire x_5100;
wire x_5101;
wire x_5102;
wire x_5103;
wire x_5104;
wire x_5105;
wire x_5106;
wire x_5107;
wire x_5108;
wire x_5109;
wire x_5110;
wire x_5111;
wire x_5112;
wire x_5113;
wire x_5114;
wire x_5115;
wire x_5116;
wire x_5117;
wire x_5118;
wire x_5119;
wire x_5120;
wire x_5121;
wire x_5122;
wire x_5123;
wire x_5124;
wire x_5125;
wire x_5126;
wire x_5127;
wire x_5128;
wire x_5129;
wire x_5130;
wire x_5131;
wire x_5132;
wire x_5133;
wire x_5134;
wire x_5135;
wire x_5136;
wire x_5137;
wire x_5138;
wire x_5139;
wire x_5140;
wire x_5141;
wire x_5142;
wire x_5143;
wire x_5144;
wire x_5145;
wire x_5146;
wire x_5147;
wire x_5148;
wire x_5149;
wire x_5150;
wire x_5151;
wire x_5152;
wire x_5153;
wire x_5154;
wire x_5155;
wire x_5156;
wire x_5157;
wire x_5158;
wire x_5159;
wire x_5160;
wire x_5161;
wire x_5162;
wire x_5163;
wire x_5164;
wire x_5165;
wire x_5166;
wire x_5167;
wire x_5168;
wire x_5169;
wire x_5170;
wire x_5171;
wire x_5172;
wire x_5173;
wire x_5174;
wire x_5175;
wire x_5176;
wire x_5177;
wire x_5178;
wire x_5179;
wire x_5180;
wire x_5181;
wire x_5182;
wire x_5183;
wire x_5184;
wire x_5185;
wire x_5186;
wire x_5187;
wire x_5188;
wire x_5189;
wire x_5190;
wire x_5191;
wire x_5192;
wire x_5193;
wire x_5194;
wire x_5195;
wire x_5196;
wire x_5197;
wire x_5198;
wire x_5199;
wire x_5200;
wire x_5201;
wire x_5202;
wire x_5203;
wire x_5204;
wire x_5205;
wire x_5206;
wire x_5207;
wire x_5208;
wire x_5209;
wire x_5210;
wire x_5211;
wire x_5212;
wire x_5213;
wire x_5214;
wire x_5215;
wire x_5216;
wire x_5217;
wire x_5218;
wire x_5219;
wire x_5220;
wire x_5221;
wire x_5222;
wire x_5223;
wire x_5224;
wire x_5225;
wire x_5226;
wire x_5227;
wire x_5228;
wire x_5229;
wire x_5230;
wire x_5231;
wire x_5232;
wire x_5233;
wire x_5234;
wire x_5235;
wire x_5236;
wire x_5237;
wire x_5238;
wire x_5239;
wire x_5240;
wire x_5241;
wire x_5242;
wire x_5243;
wire x_5244;
wire x_5245;
wire x_5246;
wire x_5247;
wire x_5248;
wire x_5249;
wire x_5250;
wire x_5251;
wire x_5252;
wire x_5253;
wire x_5254;
wire x_5255;
assign v_486 = 1;
assign v_4 = ~v_2 & ~v_3;
assign v_5 = ~v_3 & v_2;
assign v_6 = ~v_2 & v_3;
assign v_7 = v_2 & v_3;
assign v_13 = ~v_11 & ~v_12;
assign v_14 = ~v_12 & v_11;
assign v_15 = ~v_11 & v_12;
assign v_16 = v_11 & v_12;
assign v_17 = ~v_10 & v_13;
assign v_18 = v_10 & v_13;
assign v_19 = ~v_10 & v_14;
assign v_20 = v_10 & v_14;
assign v_21 = ~v_10 & v_15;
assign v_22 = v_10 & v_15;
assign v_23 = ~v_10 & v_16;
assign v_24 = v_10 & v_16;
assign v_25 = ~v_9 & v_17;
assign v_26 = v_9 & v_17;
assign v_27 = ~v_9 & v_18;
assign v_28 = v_9 & v_18;
assign v_29 = ~v_9 & v_19;
assign v_30 = v_9 & v_19;
assign v_31 = ~v_9 & v_20;
assign v_32 = v_9 & v_20;
assign v_33 = ~v_9 & v_21;
assign v_34 = v_9 & v_21;
assign v_35 = ~v_9 & v_22;
assign v_36 = v_9 & v_22;
assign v_37 = ~v_9 & v_23;
assign v_38 = v_9 & v_23;
assign v_39 = ~v_9 & v_24;
assign v_40 = v_9 & v_24;
assign v_41 = ~v_8 & v_25;
assign v_42 = v_8 & v_25;
assign v_43 = ~v_8 & v_26;
assign v_44 = v_8 & v_26;
assign v_45 = ~v_8 & v_27;
assign v_46 = v_8 & v_27;
assign v_47 = ~v_8 & v_28;
assign v_48 = v_8 & v_28;
assign v_49 = ~v_8 & v_29;
assign v_50 = v_8 & v_29;
assign v_51 = ~v_8 & v_30;
assign v_52 = v_8 & v_30;
assign v_53 = ~v_8 & v_31;
assign v_54 = v_8 & v_31;
assign v_55 = ~v_8 & v_32;
assign v_56 = v_8 & v_32;
assign v_57 = ~v_8 & v_33;
assign v_58 = v_8 & v_33;
assign v_59 = ~v_8 & v_34;
assign v_60 = v_8 & v_34;
assign v_61 = ~v_8 & v_35;
assign v_62 = v_8 & v_35;
assign v_63 = ~v_8 & v_36;
assign v_64 = v_8 & v_36;
assign v_65 = ~v_8 & v_37;
assign v_66 = v_8 & v_37;
assign v_67 = ~v_8 & v_38;
assign v_68 = v_8 & v_38;
assign v_69 = ~v_8 & v_39;
assign v_70 = v_8 & v_39;
assign v_71 = ~v_8 & v_40;
assign v_72 = v_8 & v_40;
assign v_78 = ~v_76 & ~v_77;
assign v_79 = ~v_77 & v_76;
assign v_80 = ~v_76 & v_77;
assign v_81 = v_76 & v_77;
assign v_82 = ~v_75 & v_78;
assign v_83 = v_75 & v_78;
assign v_84 = ~v_75 & v_79;
assign v_85 = v_75 & v_79;
assign v_86 = ~v_75 & v_80;
assign v_87 = v_75 & v_80;
assign v_88 = ~v_75 & v_81;
assign v_89 = v_75 & v_81;
assign v_90 = ~v_74 & v_82;
assign v_91 = v_74 & v_82;
assign v_92 = ~v_74 & v_83;
assign v_93 = v_74 & v_83;
assign v_94 = ~v_74 & v_84;
assign v_95 = v_74 & v_84;
assign v_96 = ~v_74 & v_85;
assign v_97 = v_74 & v_85;
assign v_98 = ~v_74 & v_86;
assign v_99 = v_74 & v_86;
assign v_100 = ~v_74 & v_87;
assign v_101 = v_74 & v_87;
assign v_102 = ~v_74 & v_88;
assign v_103 = v_74 & v_88;
assign v_104 = ~v_74 & v_89;
assign v_105 = v_74 & v_89;
assign v_106 = ~v_73 & v_90;
assign v_107 = v_73 & v_90;
assign v_108 = ~v_73 & v_91;
assign v_109 = v_73 & v_91;
assign v_110 = ~v_73 & v_92;
assign v_111 = v_73 & v_92;
assign v_112 = ~v_73 & v_93;
assign v_113 = v_73 & v_93;
assign v_114 = ~v_73 & v_94;
assign v_115 = v_73 & v_94;
assign v_116 = ~v_73 & v_95;
assign v_117 = v_73 & v_95;
assign v_118 = ~v_73 & v_96;
assign v_119 = v_73 & v_96;
assign v_120 = ~v_73 & v_97;
assign v_121 = v_73 & v_97;
assign v_122 = ~v_73 & v_98;
assign v_123 = v_73 & v_98;
assign v_124 = ~v_73 & v_99;
assign v_125 = v_73 & v_99;
assign v_126 = ~v_73 & v_100;
assign v_127 = v_73 & v_100;
assign v_128 = ~v_73 & v_101;
assign v_129 = v_73 & v_101;
assign v_130 = ~v_73 & v_102;
assign v_131 = v_73 & v_102;
assign v_132 = ~v_73 & v_103;
assign v_133 = v_73 & v_103;
assign v_134 = ~v_73 & v_104;
assign v_135 = v_73 & v_104;
assign v_136 = ~v_73 & v_105;
assign v_137 = v_73 & v_105;
assign v_143 = ~v_141 & ~v_142;
assign v_144 = ~v_142 & v_141;
assign v_145 = ~v_141 & v_142;
assign v_146 = v_141 & v_142;
assign v_147 = ~v_140 & v_143;
assign v_148 = v_140 & v_143;
assign v_149 = ~v_140 & v_144;
assign v_150 = v_140 & v_144;
assign v_151 = ~v_140 & v_145;
assign v_152 = v_140 & v_145;
assign v_153 = ~v_140 & v_146;
assign v_154 = v_140 & v_146;
assign v_155 = ~v_139 & v_147;
assign v_156 = v_139 & v_147;
assign v_157 = ~v_139 & v_148;
assign v_158 = v_139 & v_148;
assign v_159 = ~v_139 & v_149;
assign v_160 = v_139 & v_149;
assign v_161 = ~v_139 & v_150;
assign v_162 = v_139 & v_150;
assign v_163 = ~v_139 & v_151;
assign v_164 = v_139 & v_151;
assign v_165 = ~v_139 & v_152;
assign v_166 = v_139 & v_152;
assign v_167 = ~v_139 & v_153;
assign v_168 = v_139 & v_153;
assign v_169 = ~v_139 & v_154;
assign v_170 = v_139 & v_154;
assign v_171 = ~v_138 & v_155;
assign v_172 = v_138 & v_155;
assign v_173 = ~v_138 & v_156;
assign v_174 = v_138 & v_156;
assign v_175 = ~v_138 & v_157;
assign v_176 = v_138 & v_157;
assign v_177 = ~v_138 & v_158;
assign v_178 = v_138 & v_158;
assign v_179 = ~v_138 & v_159;
assign v_180 = v_138 & v_159;
assign v_181 = ~v_138 & v_160;
assign v_182 = v_138 & v_160;
assign v_183 = ~v_138 & v_161;
assign v_184 = v_138 & v_161;
assign v_185 = ~v_138 & v_162;
assign v_186 = v_138 & v_162;
assign v_187 = ~v_138 & v_163;
assign v_188 = v_138 & v_163;
assign v_189 = ~v_138 & v_164;
assign v_190 = v_138 & v_164;
assign v_191 = ~v_138 & v_165;
assign v_192 = v_138 & v_165;
assign v_193 = ~v_138 & v_166;
assign v_194 = v_138 & v_166;
assign v_195 = ~v_138 & v_167;
assign v_196 = v_138 & v_167;
assign v_197 = ~v_138 & v_168;
assign v_198 = v_138 & v_168;
assign v_199 = ~v_138 & v_169;
assign v_200 = v_138 & v_169;
assign v_201 = ~v_138 & v_170;
assign v_202 = v_138 & v_170;
assign v_205 = ~v_203 & ~v_204;
assign v_206 = ~v_204 & v_203;
assign v_207 = ~v_203 & v_204;
assign v_208 = v_203 & v_204;
assign v_211 = ~v_209 & ~v_210;
assign v_212 = ~v_210 & v_209;
assign v_213 = ~v_209 & v_210;
assign v_214 = v_209 & v_210;
assign v_217 = ~v_215 & ~v_216;
assign v_218 = ~v_216 & v_215;
assign v_219 = ~v_215 & v_216;
assign v_220 = v_215 & v_216;
assign v_223 = ~v_221 & ~v_222;
assign v_224 = ~v_222 & v_221;
assign v_225 = ~v_221 & v_222;
assign v_226 = v_221 & v_222;
assign v_229 = ~v_227 & ~v_228;
assign v_230 = ~v_228 & v_227;
assign v_231 = ~v_227 & v_228;
assign v_232 = v_227 & v_228;
assign v_235 = ~v_233 & ~v_234;
assign v_236 = ~v_234 & v_233;
assign v_237 = ~v_233 & v_234;
assign v_238 = v_233 & v_234;
assign v_241 = ~v_239 & ~v_240;
assign v_242 = ~v_240 & v_239;
assign v_243 = ~v_239 & v_240;
assign v_244 = v_239 & v_240;
assign v_247 = ~v_245 & ~v_246;
assign v_248 = ~v_246 & v_245;
assign v_249 = ~v_245 & v_246;
assign v_250 = v_245 & v_246;
assign v_253 = ~v_251 & ~v_252;
assign v_254 = ~v_252 & v_251;
assign v_255 = ~v_251 & v_252;
assign v_256 = v_251 & v_252;
assign v_259 = ~v_257 & ~v_258;
assign v_260 = ~v_258 & v_257;
assign v_261 = ~v_257 & v_258;
assign v_262 = v_257 & v_258;
assign v_265 = ~v_263 & ~v_264;
assign v_266 = ~v_264 & v_263;
assign v_267 = ~v_263 & v_264;
assign v_268 = v_263 & v_264;
assign v_274 = ~v_272 & ~v_273;
assign v_275 = ~v_273 & v_272;
assign v_276 = ~v_272 & v_273;
assign v_277 = v_272 & v_273;
assign v_278 = ~v_271 & v_274;
assign v_279 = v_271 & v_274;
assign v_280 = ~v_271 & v_275;
assign v_281 = v_271 & v_275;
assign v_282 = ~v_271 & v_276;
assign v_283 = v_271 & v_276;
assign v_284 = ~v_271 & v_277;
assign v_285 = v_271 & v_277;
assign v_286 = ~v_270 & v_278;
assign v_287 = v_270 & v_278;
assign v_288 = ~v_270 & v_279;
assign v_289 = v_270 & v_279;
assign v_290 = ~v_270 & v_280;
assign v_291 = v_270 & v_280;
assign v_292 = ~v_270 & v_281;
assign v_293 = v_270 & v_281;
assign v_294 = ~v_270 & v_282;
assign v_295 = v_270 & v_282;
assign v_296 = ~v_270 & v_283;
assign v_297 = v_270 & v_283;
assign v_298 = ~v_270 & v_284;
assign v_299 = v_270 & v_284;
assign v_300 = ~v_270 & v_285;
assign v_301 = v_270 & v_285;
assign v_302 = ~v_269 & v_286;
assign v_303 = v_269 & v_286;
assign v_304 = ~v_269 & v_287;
assign v_305 = v_269 & v_287;
assign v_306 = ~v_269 & v_288;
assign v_307 = v_269 & v_288;
assign v_308 = ~v_269 & v_289;
assign v_309 = v_269 & v_289;
assign v_310 = ~v_269 & v_290;
assign v_311 = v_269 & v_290;
assign v_312 = ~v_269 & v_291;
assign v_313 = v_269 & v_291;
assign v_314 = ~v_269 & v_292;
assign v_315 = v_269 & v_292;
assign v_316 = ~v_269 & v_293;
assign v_317 = v_269 & v_293;
assign v_318 = ~v_269 & v_294;
assign v_319 = v_269 & v_294;
assign v_320 = ~v_269 & v_295;
assign v_321 = v_269 & v_295;
assign v_322 = ~v_269 & v_296;
assign v_323 = v_269 & v_296;
assign v_324 = ~v_269 & v_297;
assign v_325 = v_269 & v_297;
assign v_326 = ~v_269 & v_298;
assign v_327 = v_269 & v_298;
assign v_328 = ~v_269 & v_299;
assign v_329 = v_269 & v_299;
assign v_330 = ~v_269 & v_300;
assign v_331 = v_269 & v_300;
assign v_332 = ~v_269 & v_301;
assign v_333 = v_269 & v_301;
assign v_339 = ~v_337 & ~v_338;
assign v_340 = ~v_338 & v_337;
assign v_341 = ~v_337 & v_338;
assign v_342 = v_337 & v_338;
assign v_343 = ~v_336 & v_339;
assign v_344 = v_336 & v_339;
assign v_345 = ~v_336 & v_340;
assign v_346 = v_336 & v_340;
assign v_347 = ~v_336 & v_341;
assign v_348 = v_336 & v_341;
assign v_349 = ~v_336 & v_342;
assign v_350 = v_336 & v_342;
assign v_351 = ~v_335 & v_343;
assign v_352 = v_335 & v_343;
assign v_353 = ~v_335 & v_344;
assign v_354 = v_335 & v_344;
assign v_355 = ~v_335 & v_345;
assign v_356 = v_335 & v_345;
assign v_357 = ~v_335 & v_346;
assign v_358 = v_335 & v_346;
assign v_359 = ~v_335 & v_347;
assign v_360 = v_335 & v_347;
assign v_361 = ~v_335 & v_348;
assign v_362 = v_335 & v_348;
assign v_363 = ~v_335 & v_349;
assign v_364 = v_335 & v_349;
assign v_365 = ~v_335 & v_350;
assign v_366 = v_335 & v_350;
assign v_367 = ~v_334 & v_351;
assign v_368 = v_334 & v_351;
assign v_369 = ~v_334 & v_352;
assign v_370 = v_334 & v_352;
assign v_371 = ~v_334 & v_353;
assign v_372 = v_334 & v_353;
assign v_373 = ~v_334 & v_354;
assign v_374 = v_334 & v_354;
assign v_375 = ~v_334 & v_355;
assign v_376 = v_334 & v_355;
assign v_377 = ~v_334 & v_356;
assign v_378 = v_334 & v_356;
assign v_379 = ~v_334 & v_357;
assign v_380 = v_334 & v_357;
assign v_381 = ~v_334 & v_358;
assign v_382 = v_334 & v_358;
assign v_383 = ~v_334 & v_359;
assign v_384 = v_334 & v_359;
assign v_385 = ~v_334 & v_360;
assign v_386 = v_334 & v_360;
assign v_387 = ~v_334 & v_361;
assign v_388 = v_334 & v_361;
assign v_389 = ~v_334 & v_362;
assign v_390 = v_334 & v_362;
assign v_391 = ~v_334 & v_363;
assign v_392 = v_334 & v_363;
assign v_393 = ~v_334 & v_364;
assign v_394 = v_334 & v_364;
assign v_395 = ~v_334 & v_365;
assign v_396 = v_334 & v_365;
assign v_397 = ~v_334 & v_366;
assign v_398 = v_334 & v_366;
assign v_401 = ~v_399 & ~v_400;
assign v_402 = ~v_400 & v_399;
assign v_403 = ~v_399 & v_400;
assign v_404 = v_399 & v_400;
assign v_407 = ~v_405 & ~v_406;
assign v_408 = ~v_406 & v_405;
assign v_409 = ~v_405 & v_406;
assign v_410 = v_405 & v_406;
assign v_413 = ~v_411 & ~v_412;
assign v_414 = ~v_412 & v_411;
assign v_415 = ~v_411 & v_412;
assign v_416 = v_411 & v_412;
assign v_419 = ~v_417 & ~v_418;
assign v_420 = ~v_418 & v_417;
assign v_421 = ~v_417 & v_418;
assign v_422 = v_417 & v_418;
assign v_425 = ~v_423 & ~v_424;
assign v_426 = ~v_424 & v_423;
assign v_427 = ~v_423 & v_424;
assign v_428 = v_423 & v_424;
assign v_431 = ~v_429 & ~v_430;
assign v_432 = ~v_430 & v_429;
assign v_433 = ~v_429 & v_430;
assign v_434 = v_429 & v_430;
assign v_437 = ~v_435 & ~v_436;
assign v_438 = ~v_436 & v_435;
assign v_439 = ~v_435 & v_436;
assign v_440 = v_435 & v_436;
assign v_443 = ~v_441 & ~v_442;
assign v_444 = ~v_442 & v_441;
assign v_445 = ~v_441 & v_442;
assign v_446 = v_441 & v_442;
assign v_449 = ~v_447 & ~v_448;
assign v_450 = ~v_448 & v_447;
assign v_451 = ~v_447 & v_448;
assign v_452 = v_447 & v_448;
assign v_455 = ~v_453 & ~v_454;
assign v_456 = ~v_454 & v_453;
assign v_457 = ~v_453 & v_454;
assign v_458 = v_453 & v_454;
assign v_487 = ~v_461 & ~v_462;
assign v_488 = ~v_462 & v_461;
assign v_489 = ~v_461 & v_462;
assign v_490 = v_461 & v_462;
assign v_491 = ~v_459 & ~v_460;
assign v_492 = ~v_460 & v_459;
assign v_493 = ~v_459 & v_460;
assign v_494 = v_459 & v_460;
assign v_495 = ~v_463 & ~v_464;
assign v_496 = ~v_464 & v_463;
assign v_497 = ~v_463 & v_464;
assign v_498 = v_463 & v_464;
assign v_499 = ~v_487 & v_495;
assign v_500 = ~v_487 & ~v_488;
assign v_501 = v_496 & v_500;
assign v_502 = ~v_499 & ~v_501;
assign v_503 = v_490 & v_497;
assign v_504 = ~v_503 & v_502;
assign v_505 = ~v_41 & ~v_42;
assign v_506 = ~v_43 & v_505;
assign v_507 = ~v_44 & v_506;
assign v_508 = ~v_45 & v_507;
assign v_509 = ~v_46 & v_508;
assign v_510 = ~v_495 & v_487;
assign v_511 = ~v_495 & ~v_496;
assign v_512 = v_488 & v_511;
assign v_513 = ~v_510 & ~v_512;
assign v_514 = v_489 & v_498;
assign v_515 = ~v_514 & v_513;
assign v_517 = ~v_515 & v_42;
assign v_518 = v_43 & v_515;
assign v_519 = ~v_504 & v_44;
assign v_520 = v_45 & v_516;
assign v_521 = v_46 & v_504;
assign v_524 = ~v_504 & v_523;
assign v_533 = ~v_529 & v_524;
assign v_534 = ~v_529 & ~v_530;
assign v_535 = ~v_529 & v_533;
assign v_536 = ~v_106 & v_535;
assign v_537 = v_107 & v_536;
assign v_538 = v_529 & v_537;
assign v_539 = ~v_107 & v_536;
assign v_540 = v_529 & v_539;
assign v_541 = ~v_171 & v_535;
assign v_542 = v_172 & v_541;
assign v_543 = v_529 & v_542;
assign v_544 = ~v_172 & v_541;
assign v_545 = v_529 & v_544;
assign v_546 = v_524 & v_534;
assign v_547 = ~v_530 & v_534;
assign v_548 = ~v_529 & v_547;
assign v_550 = ~v_549 & v_546;
assign v_551 = ~v_106 & v_550;
assign v_552 = v_107 & v_551;
assign v_553 = v_549 & v_552;
assign v_554 = ~v_107 & v_551;
assign v_555 = v_549 & v_554;
assign v_556 = ~v_171 & v_550;
assign v_557 = v_172 & v_556;
assign v_558 = v_549 & v_557;
assign v_559 = ~v_172 & v_556;
assign v_560 = v_549 & v_559;
assign v_561 = v_524 & v_532;
assign v_562 = ~v_531 & v_532;
assign v_563 = ~v_530 & v_562;
assign v_565 = ~v_529 & ~v_564;
assign v_567 = ~v_566 & v_561;
assign v_568 = ~v_106 & v_567;
assign v_569 = v_107 & v_568;
assign v_570 = v_566 & v_569;
assign v_571 = ~v_107 & v_568;
assign v_572 = v_566 & v_571;
assign v_573 = ~v_171 & v_567;
assign v_574 = v_172 & v_573;
assign v_575 = v_566 & v_574;
assign v_576 = ~v_172 & v_573;
assign v_577 = v_566 & v_576;
assign v_578 = ~v_171 & ~v_172;
assign v_579 = ~v_173 & v_578;
assign v_580 = ~v_174 & v_579;
assign v_581 = ~v_175 & v_580;
assign v_582 = ~v_176 & v_581;
assign v_583 = ~v_177 & v_582;
assign v_584 = ~v_468 & ~v_469;
assign v_585 = ~v_469 & v_468;
assign v_586 = ~v_468 & v_469;
assign v_587 = v_468 & v_469;
assign v_588 = ~v_205 & v_584;
assign v_589 = ~v_205 & ~v_206;
assign v_590 = v_585 & v_589;
assign v_591 = ~v_588 & ~v_590;
assign v_592 = v_208 & v_586;
assign v_593 = ~v_592 & v_591;
assign v_594 = ~v_584 & v_211;
assign v_595 = ~v_584 & ~v_585;
assign v_596 = v_212 & v_595;
assign v_597 = ~v_594 & ~v_596;
assign v_598 = v_213 & v_587;
assign v_599 = ~v_598 & v_597;
assign v_600 = ~v_584 & v_217;
assign v_601 = v_218 & v_595;
assign v_602 = ~v_600 & ~v_601;
assign v_603 = v_219 & v_587;
assign v_604 = ~v_603 & v_602;
assign v_605 = ~v_223 & v_584;
assign v_606 = ~v_223 & ~v_224;
assign v_607 = v_585 & v_606;
assign v_608 = ~v_605 & ~v_607;
assign v_609 = v_226 & v_586;
assign v_610 = ~v_609 & v_608;
assign v_613 = ~v_599 & v_172;
assign v_614 = v_173 & v_604;
assign v_615 = ~v_610 & v_174;
assign v_616 = v_175 & v_611;
assign v_617 = v_176 & v_612;
assign v_618 = v_177 & v_593;
assign v_621 = ~v_106 & ~v_107;
assign v_622 = ~v_108 & v_621;
assign v_623 = ~v_109 & v_622;
assign v_624 = ~v_110 & v_623;
assign v_625 = ~v_111 & v_624;
assign v_626 = ~v_112 & v_625;
assign v_627 = ~v_235 & v_584;
assign v_628 = ~v_235 & ~v_236;
assign v_629 = v_585 & v_628;
assign v_630 = ~v_627 & ~v_629;
assign v_631 = v_238 & v_586;
assign v_632 = ~v_631 & v_630;
assign v_633 = ~v_584 & v_241;
assign v_634 = v_242 & v_595;
assign v_635 = ~v_633 & ~v_634;
assign v_636 = v_243 & v_587;
assign v_637 = ~v_636 & v_635;
assign v_638 = ~v_584 & v_247;
assign v_639 = v_248 & v_595;
assign v_640 = ~v_638 & ~v_639;
assign v_641 = v_249 & v_587;
assign v_642 = ~v_641 & v_640;
assign v_643 = ~v_253 & v_584;
assign v_644 = ~v_253 & ~v_254;
assign v_645 = v_585 & v_644;
assign v_646 = ~v_643 & ~v_645;
assign v_647 = v_256 & v_586;
assign v_648 = ~v_647 & v_646;
assign v_650 = ~v_637 & v_107;
assign v_651 = v_108 & v_642;
assign v_652 = ~v_648 & v_109;
assign v_653 = v_110 & v_649;
assign v_654 = v_111 & v_612;
assign v_655 = v_112 & v_632;
assign v_658 = v_620 & v_657;
assign v_659 = ~v_470 & ~v_471;
assign v_660 = ~v_471 & v_470;
assign v_661 = ~v_470 & v_471;
assign v_662 = v_470 & v_471;
assign v_663 = ~v_472 & ~v_473;
assign v_664 = ~v_473 & v_472;
assign v_665 = ~v_472 & v_473;
assign v_666 = v_472 & v_473;
assign v_667 = ~v_474 & ~v_475;
assign v_668 = ~v_475 & v_474;
assign v_669 = ~v_474 & v_475;
assign v_670 = v_474 & v_475;
assign v_671 = ~v_476 & ~v_477;
assign v_672 = ~v_477 & v_476;
assign v_673 = ~v_476 & v_477;
assign v_674 = v_476 & v_477;
assign v_675 = ~v_478 & ~v_479;
assign v_676 = ~v_479 & v_478;
assign v_677 = ~v_478 & v_479;
assign v_678 = v_478 & v_479;
assign v_679 = ~v_480 & ~v_481;
assign v_680 = ~v_481 & v_480;
assign v_681 = ~v_480 & v_481;
assign v_682 = v_480 & v_481;
assign v_683 = ~v_482 & ~v_483;
assign v_684 = ~v_483 & v_482;
assign v_685 = ~v_482 & v_483;
assign v_686 = v_482 & v_483;
assign v_687 = ~v_484 & ~v_485;
assign v_688 = ~v_485 & v_484;
assign v_689 = ~v_484 & v_485;
assign v_690 = v_484 & v_485;
assign v_691 = ~v_223 & v_174;
assign v_692 = v_175 & v_229;
assign v_693 = v_176 & v_495;
assign v_694 = v_177 & v_205;
assign v_697 = ~v_253 & v_109;
assign v_698 = v_110 & v_259;
assign v_699 = v_111 & v_495;
assign v_700 = v_112 & v_235;
assign v_703 = v_696 & v_702;
assign v_704 = ~v_566 & v_683;
assign v_705 = ~v_566 & ~v_704;
assign v_706 = ~v_566 & v_684;
assign v_707 = ~v_566 & v_685;
assign v_708 = ~v_566 & v_686;
assign v_709 = ~v_205 & ~v_705;
assign v_710 = v_589 & v_706;
assign v_711 = ~v_709 & ~v_710;
assign v_712 = v_208 & v_707;
assign v_713 = ~v_712 & v_711;
assign v_714 = v_211 & v_705;
assign v_715 = ~v_706 & v_705;
assign v_716 = v_212 & v_715;
assign v_717 = ~v_714 & ~v_716;
assign v_718 = v_213 & v_708;
assign v_719 = ~v_718 & v_717;
assign v_720 = v_217 & v_705;
assign v_721 = v_218 & v_715;
assign v_722 = ~v_720 & ~v_721;
assign v_723 = v_219 & v_708;
assign v_724 = ~v_723 & v_722;
assign v_725 = ~v_223 & ~v_705;
assign v_726 = v_606 & v_706;
assign v_727 = ~v_725 & ~v_726;
assign v_728 = v_226 & v_707;
assign v_729 = ~v_728 & v_727;
assign v_732 = ~v_719 & v_172;
assign v_733 = v_173 & v_724;
assign v_734 = ~v_729 & v_174;
assign v_735 = v_175 & v_730;
assign v_736 = v_176 & v_731;
assign v_737 = v_177 & v_713;
assign v_740 = ~v_235 & ~v_705;
assign v_741 = v_628 & v_706;
assign v_742 = ~v_740 & ~v_741;
assign v_743 = v_238 & v_707;
assign v_744 = ~v_743 & v_742;
assign v_745 = v_241 & v_705;
assign v_746 = v_242 & v_715;
assign v_747 = ~v_745 & ~v_746;
assign v_748 = v_243 & v_708;
assign v_749 = ~v_748 & v_747;
assign v_750 = v_247 & v_705;
assign v_751 = v_248 & v_715;
assign v_752 = ~v_750 & ~v_751;
assign v_753 = v_249 & v_708;
assign v_754 = ~v_753 & v_752;
assign v_755 = ~v_253 & ~v_705;
assign v_756 = v_644 & v_706;
assign v_757 = ~v_755 & ~v_756;
assign v_758 = v_256 & v_707;
assign v_759 = ~v_758 & v_757;
assign v_761 = ~v_749 & v_107;
assign v_762 = v_108 & v_754;
assign v_763 = ~v_759 & v_109;
assign v_764 = v_110 & v_760;
assign v_765 = v_111 & v_731;
assign v_766 = v_112 & v_744;
assign v_769 = v_739 & v_768;
assign v_770 = ~v_566 & v_769;
assign v_771 = v_532 & v_770;
assign v_772 = ~v_549 & v_679;
assign v_773 = ~v_549 & ~v_772;
assign v_774 = ~v_549 & v_680;
assign v_775 = ~v_549 & v_681;
assign v_776 = ~v_549 & v_682;
assign v_777 = ~v_205 & ~v_773;
assign v_778 = v_589 & v_774;
assign v_779 = ~v_777 & ~v_778;
assign v_780 = v_208 & v_775;
assign v_781 = ~v_780 & v_779;
assign v_782 = v_211 & v_773;
assign v_783 = ~v_774 & v_773;
assign v_784 = v_212 & v_783;
assign v_785 = ~v_782 & ~v_784;
assign v_786 = v_213 & v_776;
assign v_787 = ~v_786 & v_785;
assign v_788 = v_217 & v_773;
assign v_789 = v_218 & v_783;
assign v_790 = ~v_788 & ~v_789;
assign v_791 = v_219 & v_776;
assign v_792 = ~v_791 & v_790;
assign v_793 = ~v_223 & ~v_773;
assign v_794 = v_606 & v_774;
assign v_795 = ~v_793 & ~v_794;
assign v_796 = v_226 & v_775;
assign v_797 = ~v_796 & v_795;
assign v_800 = ~v_787 & v_172;
assign v_801 = v_173 & v_792;
assign v_802 = ~v_797 & v_174;
assign v_803 = v_175 & v_798;
assign v_804 = v_176 & v_799;
assign v_805 = v_177 & v_781;
assign v_808 = ~v_235 & ~v_773;
assign v_809 = v_628 & v_774;
assign v_810 = ~v_808 & ~v_809;
assign v_811 = v_238 & v_775;
assign v_812 = ~v_811 & v_810;
assign v_813 = v_241 & v_773;
assign v_814 = v_242 & v_783;
assign v_815 = ~v_813 & ~v_814;
assign v_816 = v_243 & v_776;
assign v_817 = ~v_816 & v_815;
assign v_818 = v_247 & v_773;
assign v_819 = v_248 & v_783;
assign v_820 = ~v_818 & ~v_819;
assign v_821 = v_249 & v_776;
assign v_822 = ~v_821 & v_820;
assign v_823 = ~v_253 & ~v_773;
assign v_824 = v_644 & v_774;
assign v_825 = ~v_823 & ~v_824;
assign v_826 = v_256 & v_775;
assign v_827 = ~v_826 & v_825;
assign v_829 = ~v_817 & v_107;
assign v_830 = v_108 & v_822;
assign v_831 = ~v_827 & v_109;
assign v_832 = v_110 & v_828;
assign v_833 = v_111 & v_799;
assign v_834 = v_112 & v_812;
assign v_837 = v_807 & v_836;
assign v_838 = ~v_549 & v_837;
assign v_839 = v_534 & v_838;
assign v_840 = ~v_529 & v_675;
assign v_841 = ~v_529 & ~v_840;
assign v_842 = ~v_529 & v_676;
assign v_843 = ~v_529 & v_677;
assign v_844 = ~v_529 & v_678;
assign v_845 = ~v_205 & ~v_841;
assign v_846 = v_589 & v_842;
assign v_847 = ~v_845 & ~v_846;
assign v_848 = v_208 & v_843;
assign v_849 = ~v_848 & v_847;
assign v_850 = v_211 & v_841;
assign v_851 = ~v_842 & v_841;
assign v_852 = v_212 & v_851;
assign v_853 = ~v_850 & ~v_852;
assign v_854 = v_213 & v_844;
assign v_855 = ~v_854 & v_853;
assign v_856 = v_217 & v_841;
assign v_857 = v_218 & v_851;
assign v_858 = ~v_856 & ~v_857;
assign v_859 = v_219 & v_844;
assign v_860 = ~v_859 & v_858;
assign v_861 = ~v_223 & ~v_841;
assign v_862 = v_606 & v_842;
assign v_863 = ~v_861 & ~v_862;
assign v_864 = v_226 & v_843;
assign v_865 = ~v_864 & v_863;
assign v_868 = ~v_855 & v_172;
assign v_869 = v_173 & v_860;
assign v_870 = ~v_865 & v_174;
assign v_871 = v_175 & v_866;
assign v_872 = v_176 & v_867;
assign v_873 = v_177 & v_849;
assign v_876 = ~v_235 & ~v_841;
assign v_877 = v_628 & v_842;
assign v_878 = ~v_876 & ~v_877;
assign v_879 = v_238 & v_843;
assign v_880 = ~v_879 & v_878;
assign v_881 = v_241 & v_841;
assign v_882 = v_242 & v_851;
assign v_883 = ~v_881 & ~v_882;
assign v_884 = v_243 & v_844;
assign v_885 = ~v_884 & v_883;
assign v_886 = v_247 & v_841;
assign v_887 = v_248 & v_851;
assign v_888 = ~v_886 & ~v_887;
assign v_889 = v_249 & v_844;
assign v_890 = ~v_889 & v_888;
assign v_891 = ~v_253 & ~v_841;
assign v_892 = v_644 & v_842;
assign v_893 = ~v_891 & ~v_892;
assign v_894 = v_256 & v_843;
assign v_895 = ~v_894 & v_893;
assign v_897 = ~v_885 & v_107;
assign v_898 = v_108 & v_890;
assign v_899 = ~v_895 & v_109;
assign v_900 = v_110 & v_896;
assign v_901 = v_111 & v_867;
assign v_902 = v_112 & v_880;
assign v_905 = v_875 & v_904;
assign v_906 = ~v_529 & v_905;
assign v_907 = ~v_529 & v_906;
assign v_908 = ~v_839 & ~v_907;
assign v_910 = v_839 & v_907;
assign v_911 = ~v_771 & v_908;
assign v_914 = v_771 & v_910;
assign v_916 = ~v_491 & v_915;
assign v_917 = v_524 & v_916;
assign v_918 = ~v_529 & v_907;
assign v_920 = v_907 & v_918;
assign v_921 = ~v_549 & ~v_907;
assign v_924 = v_839 & v_921;
assign v_926 = ~v_908 & v_923;
assign v_927 = ~v_908 & v_924;
assign v_928 = ~v_566 & v_908;
assign v_932 = v_771 & v_928;
assign v_933 = ~v_911 & ~v_929;
assign v_934 = ~v_911 & v_930;
assign v_935 = ~v_911 & v_931;
assign v_936 = ~v_911 & v_932;
assign v_937 = ~v_911 & v_929;
assign v_938 = v_917 & v_929;
assign v_939 = v_675 & v_930;
assign v_940 = ~v_929 & ~v_939;
assign v_941 = v_676 & v_930;
assign v_942 = v_677 & v_930;
assign v_943 = v_678 & v_930;
assign v_944 = v_679 & v_931;
assign v_945 = ~v_944 & v_940;
assign v_946 = v_680 & v_931;
assign v_947 = ~v_941 & ~v_946;
assign v_948 = v_681 & v_931;
assign v_949 = ~v_942 & ~v_948;
assign v_950 = v_682 & v_931;
assign v_951 = ~v_943 & ~v_950;
assign v_952 = v_683 & v_932;
assign v_953 = ~v_952 & v_945;
assign v_954 = v_684 & v_932;
assign v_955 = ~v_954 & v_947;
assign v_956 = v_685 & v_932;
assign v_957 = ~v_956 & v_949;
assign v_958 = v_686 & v_932;
assign v_959 = ~v_958 & v_951;
assign v_961 = v_915 & v_960;
assign v_963 = ~v_491 & ~v_492;
assign v_964 = ~v_962 & v_963;
assign v_965 = v_524 & v_964;
assign v_966 = ~v_549 & v_907;
assign v_967 = v_839 & v_966;
assign v_969 = ~v_909 & v_967;
assign v_970 = ~v_566 & v_909;
assign v_973 = v_771 & v_970;
assign v_974 = ~v_912 & ~v_971;
assign v_975 = ~v_912 & v_972;
assign v_976 = ~v_912 & v_973;
assign v_977 = ~v_912 & v_971;
assign v_978 = v_965 & v_971;
assign v_979 = v_679 & v_972;
assign v_980 = ~v_971 & ~v_979;
assign v_981 = v_680 & v_972;
assign v_982 = v_681 & v_972;
assign v_983 = v_682 & v_972;
assign v_984 = v_683 & v_973;
assign v_985 = ~v_984 & v_980;
assign v_986 = v_684 & v_973;
assign v_987 = ~v_981 & ~v_986;
assign v_988 = v_685 & v_973;
assign v_989 = ~v_982 & ~v_988;
assign v_990 = v_686 & v_973;
assign v_991 = ~v_983 & ~v_990;
assign v_993 = ~v_962 & v_992;
assign v_995 = ~v_994 & v_494;
assign v_996 = v_524 & v_995;
assign v_997 = ~v_566 & v_910;
assign v_998 = v_771 & v_997;
assign v_999 = ~v_913 & v_998;
assign v_1000 = ~v_913 & ~v_998;
assign v_1001 = ~v_998 & v_996;
assign v_1002 = v_683 & v_998;
assign v_1003 = ~v_1002 & v_998;
assign v_1004 = v_684 & v_998;
assign v_1005 = v_685 & v_998;
assign v_1006 = v_686 & v_998;
assign v_1008 = ~v_994 & v_1007;
assign v_1010 = ~v_1009 & v_671;
assign v_1011 = v_494 & v_524;
assign v_1012 = ~v_1007 & v_1011;
assign v_1013 = v_524 & v_963;
assign v_1014 = ~v_992 & v_1013;
assign v_1015 = ~v_1012 & ~v_1014;
assign v_1016 = ~v_491 & v_524;
assign v_1017 = ~v_960 & v_1016;
assign v_1018 = ~v_1017 & v_1015;
assign v_1019 = ~v_915 & v_524;
assign v_1020 = ~v_1019 & v_1018;
assign v_1021 = v_524 & v_1020;
assign v_1022 = ~v_504 & v_1021;
assign v_1023 = v_495 & v_500;
assign v_1024 = v_490 & v_496;
assign v_1025 = ~v_1023 & ~v_1024;
assign v_1026 = ~v_495 & v_488;
assign v_1027 = ~v_487 & ~v_1026;
assign v_1028 = v_489 & v_511;
assign v_1029 = ~v_1028 & v_1027;
assign v_1030 = v_490 & v_498;
assign v_1031 = ~v_1030 & v_1029;
assign v_1033 = ~v_1031 & v_42;
assign v_1034 = v_43 & v_1031;
assign v_1035 = ~v_1025 & v_44;
assign v_1036 = v_45 & v_1032;
assign v_1037 = v_46 & v_1025;
assign v_1040 = v_1022 & v_1039;
assign v_1041 = v_5 & v_487;
assign v_1045 = ~v_5 & v_498;
assign v_1046 = ~v_4 & v_1041;
assign v_1051 = ~v_1046 & v_1040;
assign v_1052 = ~v_1046 & ~v_1047;
assign v_1053 = ~v_1048 & v_1052;
assign v_1054 = ~v_1046 & v_1051;
assign v_1055 = ~v_106 & v_1054;
assign v_1056 = v_107 & v_1055;
assign v_1057 = v_1046 & v_1056;
assign v_1058 = ~v_107 & v_1055;
assign v_1059 = v_1046 & v_1058;
assign v_1060 = ~v_171 & v_1054;
assign v_1061 = v_172 & v_1060;
assign v_1062 = v_1046 & v_1061;
assign v_1063 = ~v_172 & v_1060;
assign v_1064 = v_1046 & v_1063;
assign v_1065 = v_1040 & v_1052;
assign v_1066 = ~v_1047 & v_1052;
assign v_1068 = ~v_1046 & ~v_1067;
assign v_1070 = ~v_1069 & v_1065;
assign v_1071 = ~v_106 & v_1070;
assign v_1072 = v_107 & v_1071;
assign v_1073 = v_1069 & v_1072;
assign v_1074 = ~v_107 & v_1071;
assign v_1075 = v_1069 & v_1074;
assign v_1076 = ~v_171 & v_1070;
assign v_1077 = v_172 & v_1076;
assign v_1078 = v_1069 & v_1077;
assign v_1079 = ~v_172 & v_1076;
assign v_1080 = v_1069 & v_1079;
assign v_1081 = v_1040 & v_1053;
assign v_1082 = ~v_1048 & v_1053;
assign v_1084 = ~v_1047 & ~v_1083;
assign v_1086 = ~v_1046 & ~v_1085;
assign v_1088 = ~v_1087 & v_1081;
assign v_1089 = ~v_106 & v_1088;
assign v_1090 = v_107 & v_1089;
assign v_1091 = v_1087 & v_1090;
assign v_1092 = ~v_107 & v_1089;
assign v_1093 = v_1087 & v_1092;
assign v_1094 = ~v_171 & v_1088;
assign v_1095 = v_172 & v_1094;
assign v_1096 = v_1087 & v_1095;
assign v_1097 = ~v_172 & v_1094;
assign v_1098 = v_1087 & v_1097;
assign v_1099 = v_1040 & v_1050;
assign v_1100 = ~v_1049 & v_1050;
assign v_1102 = ~v_1048 & ~v_1101;
assign v_1104 = ~v_1047 & ~v_1103;
assign v_1106 = ~v_1046 & ~v_1105;
assign v_1108 = ~v_1107 & v_1099;
assign v_1109 = ~v_106 & v_1108;
assign v_1110 = v_107 & v_1109;
assign v_1111 = v_1107 & v_1110;
assign v_1112 = ~v_107 & v_1109;
assign v_1113 = v_1107 & v_1112;
assign v_1114 = ~v_171 & v_1108;
assign v_1115 = v_172 & v_1114;
assign v_1116 = v_1107 & v_1115;
assign v_1117 = ~v_172 & v_1114;
assign v_1118 = v_1107 & v_1117;
assign v_1120 = v_176 & v_1119;
assign v_1123 = v_111 & v_1119;
assign v_1126 = v_1122 & v_1125;
assign v_1127 = ~v_1107 & v_687;
assign v_1128 = ~v_1107 & ~v_1127;
assign v_1129 = ~v_1107 & v_688;
assign v_1130 = ~v_1107 & v_689;
assign v_1131 = ~v_1107 & v_690;
assign v_1132 = ~v_205 & ~v_1128;
assign v_1133 = v_589 & v_1129;
assign v_1134 = ~v_1132 & ~v_1133;
assign v_1135 = v_208 & v_1130;
assign v_1136 = ~v_1135 & v_1134;
assign v_1137 = v_211 & v_1128;
assign v_1138 = ~v_1129 & v_1128;
assign v_1139 = v_212 & v_1138;
assign v_1140 = ~v_1137 & ~v_1139;
assign v_1141 = v_213 & v_1131;
assign v_1142 = ~v_1141 & v_1140;
assign v_1143 = v_217 & v_1128;
assign v_1144 = v_218 & v_1138;
assign v_1145 = ~v_1143 & ~v_1144;
assign v_1146 = v_219 & v_1131;
assign v_1147 = ~v_1146 & v_1145;
assign v_1148 = ~v_223 & ~v_1128;
assign v_1149 = v_606 & v_1129;
assign v_1150 = ~v_1148 & ~v_1149;
assign v_1151 = v_226 & v_1130;
assign v_1152 = ~v_1151 & v_1150;
assign v_1155 = ~v_1142 & v_172;
assign v_1156 = v_173 & v_1147;
assign v_1157 = ~v_1152 & v_174;
assign v_1158 = v_175 & v_1153;
assign v_1159 = v_176 & v_1154;
assign v_1160 = v_177 & v_1136;
assign v_1163 = ~v_235 & ~v_1128;
assign v_1164 = v_628 & v_1129;
assign v_1165 = ~v_1163 & ~v_1164;
assign v_1166 = v_238 & v_1130;
assign v_1167 = ~v_1166 & v_1165;
assign v_1168 = v_241 & v_1128;
assign v_1169 = v_242 & v_1138;
assign v_1170 = ~v_1168 & ~v_1169;
assign v_1171 = v_243 & v_1131;
assign v_1172 = ~v_1171 & v_1170;
assign v_1173 = v_247 & v_1128;
assign v_1174 = v_248 & v_1138;
assign v_1175 = ~v_1173 & ~v_1174;
assign v_1176 = v_249 & v_1131;
assign v_1177 = ~v_1176 & v_1175;
assign v_1178 = ~v_253 & ~v_1128;
assign v_1179 = v_644 & v_1129;
assign v_1180 = ~v_1178 & ~v_1179;
assign v_1181 = v_256 & v_1130;
assign v_1182 = ~v_1181 & v_1180;
assign v_1184 = ~v_1172 & v_107;
assign v_1185 = v_108 & v_1177;
assign v_1186 = ~v_1182 & v_109;
assign v_1187 = v_110 & v_1183;
assign v_1188 = v_111 & v_1154;
assign v_1189 = v_112 & v_1167;
assign v_1192 = v_1162 & v_1191;
assign v_1193 = ~v_1107 & v_1192;
assign v_1194 = v_1050 & v_1193;
assign v_1195 = ~v_1087 & v_683;
assign v_1196 = ~v_1087 & ~v_1195;
assign v_1197 = ~v_1087 & v_684;
assign v_1198 = ~v_1087 & v_685;
assign v_1199 = ~v_1087 & v_686;
assign v_1200 = ~v_205 & ~v_1196;
assign v_1201 = v_589 & v_1197;
assign v_1202 = ~v_1200 & ~v_1201;
assign v_1203 = v_208 & v_1198;
assign v_1204 = ~v_1203 & v_1202;
assign v_1205 = v_211 & v_1196;
assign v_1206 = ~v_1197 & v_1196;
assign v_1207 = v_212 & v_1206;
assign v_1208 = ~v_1205 & ~v_1207;
assign v_1209 = v_213 & v_1199;
assign v_1210 = ~v_1209 & v_1208;
assign v_1211 = v_217 & v_1196;
assign v_1212 = v_218 & v_1206;
assign v_1213 = ~v_1211 & ~v_1212;
assign v_1214 = v_219 & v_1199;
assign v_1215 = ~v_1214 & v_1213;
assign v_1216 = ~v_223 & ~v_1196;
assign v_1217 = v_606 & v_1197;
assign v_1218 = ~v_1216 & ~v_1217;
assign v_1219 = v_226 & v_1198;
assign v_1220 = ~v_1219 & v_1218;
assign v_1223 = ~v_1210 & v_172;
assign v_1224 = v_173 & v_1215;
assign v_1225 = ~v_1220 & v_174;
assign v_1226 = v_175 & v_1221;
assign v_1227 = v_176 & v_1222;
assign v_1228 = v_177 & v_1204;
assign v_1231 = ~v_235 & ~v_1196;
assign v_1232 = v_628 & v_1197;
assign v_1233 = ~v_1231 & ~v_1232;
assign v_1234 = v_238 & v_1198;
assign v_1235 = ~v_1234 & v_1233;
assign v_1236 = v_241 & v_1196;
assign v_1237 = v_242 & v_1206;
assign v_1238 = ~v_1236 & ~v_1237;
assign v_1239 = v_243 & v_1199;
assign v_1240 = ~v_1239 & v_1238;
assign v_1241 = v_247 & v_1196;
assign v_1242 = v_248 & v_1206;
assign v_1243 = ~v_1241 & ~v_1242;
assign v_1244 = v_249 & v_1199;
assign v_1245 = ~v_1244 & v_1243;
assign v_1246 = ~v_253 & ~v_1196;
assign v_1247 = v_644 & v_1197;
assign v_1248 = ~v_1246 & ~v_1247;
assign v_1249 = v_256 & v_1198;
assign v_1250 = ~v_1249 & v_1248;
assign v_1252 = ~v_1240 & v_107;
assign v_1253 = v_108 & v_1245;
assign v_1254 = ~v_1250 & v_109;
assign v_1255 = v_110 & v_1251;
assign v_1256 = v_111 & v_1222;
assign v_1257 = v_112 & v_1235;
assign v_1260 = v_1230 & v_1259;
assign v_1261 = ~v_1087 & v_1260;
assign v_1262 = v_1053 & v_1261;
assign v_1263 = ~v_1069 & v_679;
assign v_1264 = ~v_1069 & ~v_1263;
assign v_1265 = ~v_1069 & v_680;
assign v_1266 = ~v_1069 & v_681;
assign v_1267 = ~v_1069 & v_682;
assign v_1268 = ~v_205 & ~v_1264;
assign v_1269 = v_589 & v_1265;
assign v_1270 = ~v_1268 & ~v_1269;
assign v_1271 = v_208 & v_1266;
assign v_1272 = ~v_1271 & v_1270;
assign v_1273 = v_211 & v_1264;
assign v_1274 = ~v_1265 & v_1264;
assign v_1275 = v_212 & v_1274;
assign v_1276 = ~v_1273 & ~v_1275;
assign v_1277 = v_213 & v_1267;
assign v_1278 = ~v_1277 & v_1276;
assign v_1279 = v_217 & v_1264;
assign v_1280 = v_218 & v_1274;
assign v_1281 = ~v_1279 & ~v_1280;
assign v_1282 = v_219 & v_1267;
assign v_1283 = ~v_1282 & v_1281;
assign v_1284 = ~v_223 & ~v_1264;
assign v_1285 = v_606 & v_1265;
assign v_1286 = ~v_1284 & ~v_1285;
assign v_1287 = v_226 & v_1266;
assign v_1288 = ~v_1287 & v_1286;
assign v_1291 = ~v_1278 & v_172;
assign v_1292 = v_173 & v_1283;
assign v_1293 = ~v_1288 & v_174;
assign v_1294 = v_175 & v_1289;
assign v_1295 = v_176 & v_1290;
assign v_1296 = v_177 & v_1272;
assign v_1299 = ~v_235 & ~v_1264;
assign v_1300 = v_628 & v_1265;
assign v_1301 = ~v_1299 & ~v_1300;
assign v_1302 = v_238 & v_1266;
assign v_1303 = ~v_1302 & v_1301;
assign v_1304 = v_241 & v_1264;
assign v_1305 = v_242 & v_1274;
assign v_1306 = ~v_1304 & ~v_1305;
assign v_1307 = v_243 & v_1267;
assign v_1308 = ~v_1307 & v_1306;
assign v_1309 = v_247 & v_1264;
assign v_1310 = v_248 & v_1274;
assign v_1311 = ~v_1309 & ~v_1310;
assign v_1312 = v_249 & v_1267;
assign v_1313 = ~v_1312 & v_1311;
assign v_1314 = ~v_253 & ~v_1264;
assign v_1315 = v_644 & v_1265;
assign v_1316 = ~v_1314 & ~v_1315;
assign v_1317 = v_256 & v_1266;
assign v_1318 = ~v_1317 & v_1316;
assign v_1320 = ~v_1308 & v_107;
assign v_1321 = v_108 & v_1313;
assign v_1322 = ~v_1318 & v_109;
assign v_1323 = v_110 & v_1319;
assign v_1324 = v_111 & v_1290;
assign v_1325 = v_112 & v_1303;
assign v_1328 = v_1298 & v_1327;
assign v_1329 = ~v_1069 & v_1328;
assign v_1330 = v_1052 & v_1329;
assign v_1331 = ~v_1046 & v_675;
assign v_1332 = ~v_1046 & ~v_1331;
assign v_1333 = ~v_1046 & v_676;
assign v_1334 = ~v_1046 & v_677;
assign v_1335 = ~v_1046 & v_678;
assign v_1336 = ~v_205 & ~v_1332;
assign v_1337 = v_589 & v_1333;
assign v_1338 = ~v_1336 & ~v_1337;
assign v_1339 = v_208 & v_1334;
assign v_1340 = ~v_1339 & v_1338;
assign v_1341 = v_211 & v_1332;
assign v_1342 = ~v_1333 & v_1332;
assign v_1343 = v_212 & v_1342;
assign v_1344 = ~v_1341 & ~v_1343;
assign v_1345 = v_213 & v_1335;
assign v_1346 = ~v_1345 & v_1344;
assign v_1347 = v_217 & v_1332;
assign v_1348 = v_218 & v_1342;
assign v_1349 = ~v_1347 & ~v_1348;
assign v_1350 = v_219 & v_1335;
assign v_1351 = ~v_1350 & v_1349;
assign v_1352 = ~v_223 & ~v_1332;
assign v_1353 = v_606 & v_1333;
assign v_1354 = ~v_1352 & ~v_1353;
assign v_1355 = v_226 & v_1334;
assign v_1356 = ~v_1355 & v_1354;
assign v_1359 = ~v_1346 & v_172;
assign v_1360 = v_173 & v_1351;
assign v_1361 = ~v_1356 & v_174;
assign v_1362 = v_175 & v_1357;
assign v_1363 = v_176 & v_1358;
assign v_1364 = v_177 & v_1340;
assign v_1367 = ~v_235 & ~v_1332;
assign v_1368 = v_628 & v_1333;
assign v_1369 = ~v_1367 & ~v_1368;
assign v_1370 = v_238 & v_1334;
assign v_1371 = ~v_1370 & v_1369;
assign v_1372 = v_241 & v_1332;
assign v_1373 = v_242 & v_1342;
assign v_1374 = ~v_1372 & ~v_1373;
assign v_1375 = v_243 & v_1335;
assign v_1376 = ~v_1375 & v_1374;
assign v_1377 = v_247 & v_1332;
assign v_1378 = v_248 & v_1342;
assign v_1379 = ~v_1377 & ~v_1378;
assign v_1380 = v_249 & v_1335;
assign v_1381 = ~v_1380 & v_1379;
assign v_1382 = ~v_253 & ~v_1332;
assign v_1383 = v_644 & v_1333;
assign v_1384 = ~v_1382 & ~v_1383;
assign v_1385 = v_256 & v_1334;
assign v_1386 = ~v_1385 & v_1384;
assign v_1388 = ~v_1376 & v_107;
assign v_1389 = v_108 & v_1381;
assign v_1390 = ~v_1386 & v_109;
assign v_1391 = v_110 & v_1387;
assign v_1392 = v_111 & v_1358;
assign v_1393 = v_112 & v_1371;
assign v_1396 = v_1366 & v_1395;
assign v_1397 = ~v_1046 & v_1396;
assign v_1398 = ~v_1046 & v_1397;
assign v_1399 = ~v_1330 & ~v_1398;
assign v_1401 = v_1330 & v_1398;
assign v_1402 = ~v_1262 & v_1399;
assign v_1405 = v_1262 & v_1401;
assign v_1406 = ~v_1194 & v_1402;
assign v_1410 = v_1194 & v_1405;
assign v_1412 = v_1040 & v_1411;
assign v_1413 = v_491 & v_495;
assign v_1414 = v_491 & v_496;
assign v_1415 = v_491 & v_497;
assign v_1416 = v_491 & v_498;
assign v_1417 = ~v_1046 & v_1398;
assign v_1419 = v_1398 & v_1417;
assign v_1420 = ~v_1069 & ~v_1398;
assign v_1423 = v_1330 & v_1420;
assign v_1425 = ~v_1399 & v_1422;
assign v_1426 = ~v_1399 & v_1423;
assign v_1427 = ~v_1087 & v_1399;
assign v_1431 = v_1262 & v_1427;
assign v_1433 = ~v_1402 & v_1429;
assign v_1434 = ~v_1402 & v_1430;
assign v_1435 = ~v_1402 & v_1431;
assign v_1436 = ~v_1107 & v_1402;
assign v_1441 = v_1194 & v_1436;
assign v_1442 = ~v_1406 & v_1437;
assign v_1443 = ~v_1406 & v_1438;
assign v_1444 = ~v_1406 & v_1439;
assign v_1445 = ~v_1406 & v_1440;
assign v_1446 = ~v_1406 & v_1441;
assign v_1447 = v_1412 & v_1437;
assign v_1448 = v_675 & v_1438;
assign v_1449 = ~v_1437 & ~v_1448;
assign v_1450 = v_676 & v_1438;
assign v_1451 = v_677 & v_1438;
assign v_1452 = v_678 & v_1438;
assign v_1453 = v_679 & v_1439;
assign v_1454 = ~v_1453 & v_1449;
assign v_1455 = v_680 & v_1439;
assign v_1456 = ~v_1450 & ~v_1455;
assign v_1457 = v_681 & v_1439;
assign v_1458 = ~v_1451 & ~v_1457;
assign v_1459 = v_682 & v_1439;
assign v_1460 = ~v_1452 & ~v_1459;
assign v_1461 = v_683 & v_1440;
assign v_1462 = ~v_1461 & v_1454;
assign v_1463 = v_684 & v_1440;
assign v_1464 = ~v_1463 & v_1456;
assign v_1465 = v_685 & v_1440;
assign v_1466 = ~v_1465 & v_1458;
assign v_1467 = v_686 & v_1440;
assign v_1468 = ~v_1467 & v_1460;
assign v_1469 = v_687 & v_1441;
assign v_1470 = ~v_1469 & v_1462;
assign v_1471 = v_688 & v_1441;
assign v_1472 = ~v_1471 & v_1464;
assign v_1473 = v_689 & v_1441;
assign v_1474 = ~v_1473 & v_1466;
assign v_1475 = v_690 & v_1441;
assign v_1476 = ~v_1475 & v_1468;
assign v_1477 = ~v_491 & v_659;
assign v_1478 = ~v_491 & v_660;
assign v_1479 = ~v_491 & v_661;
assign v_1480 = ~v_491 & v_662;
assign v_1481 = v_675 & v_1413;
assign v_1482 = ~v_1477 & ~v_1481;
assign v_1483 = v_676 & v_1413;
assign v_1484 = ~v_1478 & ~v_1483;
assign v_1485 = v_677 & v_1413;
assign v_1486 = ~v_1479 & ~v_1485;
assign v_1487 = v_678 & v_1413;
assign v_1488 = ~v_1480 & ~v_1487;
assign v_1489 = v_679 & v_1414;
assign v_1490 = ~v_1489 & v_1482;
assign v_1491 = v_680 & v_1414;
assign v_1492 = ~v_1491 & v_1484;
assign v_1493 = v_681 & v_1414;
assign v_1494 = ~v_1493 & v_1486;
assign v_1495 = v_682 & v_1414;
assign v_1496 = ~v_1495 & v_1488;
assign v_1497 = v_683 & v_1415;
assign v_1498 = ~v_1497 & v_1490;
assign v_1499 = v_684 & v_1415;
assign v_1500 = ~v_1499 & v_1492;
assign v_1501 = v_685 & v_1415;
assign v_1502 = ~v_1501 & v_1494;
assign v_1503 = v_686 & v_1415;
assign v_1504 = ~v_1503 & v_1496;
assign v_1505 = v_687 & v_1416;
assign v_1506 = ~v_1505 & v_1498;
assign v_1507 = v_688 & v_1416;
assign v_1508 = ~v_1507 & v_1500;
assign v_1509 = v_689 & v_1416;
assign v_1510 = ~v_1509 & v_1502;
assign v_1511 = v_690 & v_1416;
assign v_1512 = ~v_1511 & v_1504;
assign v_1514 = v_1411 & v_1513;
assign v_1515 = ~v_491 & v_1514;
assign v_1516 = v_1040 & v_1515;
assign v_1517 = ~v_492 & ~v_963;
assign v_1518 = ~v_492 & v_963;
assign v_1519 = v_492 & v_495;
assign v_1520 = v_492 & v_496;
assign v_1521 = v_492 & v_497;
assign v_1522 = v_492 & v_498;
assign v_1523 = v_1516 & v_1517;
assign v_1524 = ~v_1069 & v_1398;
assign v_1525 = v_1330 & v_1524;
assign v_1527 = ~v_1400 & v_1525;
assign v_1528 = ~v_1087 & v_1400;
assign v_1531 = v_1262 & v_1528;
assign v_1533 = ~v_1403 & v_1530;
assign v_1534 = ~v_1403 & v_1531;
assign v_1535 = ~v_1107 & v_1403;
assign v_1539 = v_1194 & v_1535;
assign v_1540 = ~v_1407 & v_1536;
assign v_1541 = ~v_1407 & v_1537;
assign v_1542 = ~v_1407 & v_1538;
assign v_1543 = ~v_1407 & v_1539;
assign v_1544 = v_1516 & v_1536;
assign v_1545 = v_679 & v_1537;
assign v_1546 = ~v_1536 & ~v_1545;
assign v_1547 = v_680 & v_1537;
assign v_1548 = v_681 & v_1537;
assign v_1549 = v_682 & v_1537;
assign v_1550 = v_683 & v_1538;
assign v_1551 = ~v_1550 & v_1546;
assign v_1552 = v_684 & v_1538;
assign v_1553 = ~v_1547 & ~v_1552;
assign v_1554 = v_685 & v_1538;
assign v_1555 = ~v_1548 & ~v_1554;
assign v_1556 = v_686 & v_1538;
assign v_1557 = ~v_1549 & ~v_1556;
assign v_1558 = v_687 & v_1539;
assign v_1559 = ~v_1558 & v_1551;
assign v_1560 = v_688 & v_1539;
assign v_1561 = ~v_1560 & v_1553;
assign v_1562 = v_689 & v_1539;
assign v_1563 = ~v_1562 & v_1555;
assign v_1564 = v_690 & v_1539;
assign v_1565 = ~v_1564 & v_1557;
assign v_1566 = v_663 & v_1518;
assign v_1567 = ~v_1517 & ~v_1566;
assign v_1568 = v_664 & v_1518;
assign v_1569 = v_665 & v_1518;
assign v_1570 = v_666 & v_1518;
assign v_1571 = v_675 & v_1519;
assign v_1572 = ~v_1571 & v_1567;
assign v_1573 = v_676 & v_1519;
assign v_1574 = ~v_1568 & ~v_1573;
assign v_1575 = v_677 & v_1519;
assign v_1576 = ~v_1569 & ~v_1575;
assign v_1577 = v_678 & v_1519;
assign v_1578 = ~v_1570 & ~v_1577;
assign v_1579 = v_679 & v_1520;
assign v_1580 = ~v_1579 & v_1572;
assign v_1581 = v_680 & v_1520;
assign v_1582 = ~v_1581 & v_1574;
assign v_1583 = v_681 & v_1520;
assign v_1584 = ~v_1583 & v_1576;
assign v_1585 = v_682 & v_1520;
assign v_1586 = ~v_1585 & v_1578;
assign v_1587 = v_683 & v_1521;
assign v_1588 = ~v_1587 & v_1580;
assign v_1589 = v_684 & v_1521;
assign v_1590 = ~v_1589 & v_1582;
assign v_1591 = v_685 & v_1521;
assign v_1592 = ~v_1591 & v_1584;
assign v_1593 = v_686 & v_1521;
assign v_1594 = ~v_1593 & v_1586;
assign v_1595 = v_687 & v_1522;
assign v_1596 = ~v_1595 & v_1588;
assign v_1597 = v_688 & v_1522;
assign v_1598 = ~v_1597 & v_1590;
assign v_1599 = v_689 & v_1522;
assign v_1600 = ~v_1599 & v_1592;
assign v_1601 = v_690 & v_1522;
assign v_1602 = ~v_1601 & v_1594;
assign v_1604 = v_1514 & v_1603;
assign v_1606 = ~v_1605 & v_963;
assign v_1607 = v_1040 & v_1606;
assign v_1608 = ~v_493 & ~v_494;
assign v_1609 = ~v_493 & v_494;
assign v_1610 = v_493 & v_495;
assign v_1611 = v_493 & v_496;
assign v_1612 = v_493 & v_497;
assign v_1613 = v_493 & v_498;
assign v_1614 = v_1607 & v_1608;
assign v_1615 = ~v_1087 & v_1401;
assign v_1616 = v_1262 & v_1615;
assign v_1618 = ~v_1404 & v_1616;
assign v_1619 = ~v_1107 & v_1404;
assign v_1622 = v_1194 & v_1619;
assign v_1623 = ~v_1408 & v_1620;
assign v_1624 = ~v_1408 & v_1621;
assign v_1625 = ~v_1408 & v_1622;
assign v_1626 = v_1607 & v_1620;
assign v_1627 = v_683 & v_1621;
assign v_1628 = ~v_1620 & ~v_1627;
assign v_1629 = v_684 & v_1621;
assign v_1630 = v_685 & v_1621;
assign v_1631 = v_686 & v_1621;
assign v_1632 = v_687 & v_1622;
assign v_1633 = ~v_1632 & v_1628;
assign v_1634 = v_688 & v_1622;
assign v_1635 = ~v_1629 & ~v_1634;
assign v_1636 = v_689 & v_1622;
assign v_1637 = ~v_1630 & ~v_1636;
assign v_1638 = v_690 & v_1622;
assign v_1639 = ~v_1631 & ~v_1638;
assign v_1640 = v_667 & v_1609;
assign v_1641 = ~v_1608 & ~v_1640;
assign v_1642 = v_668 & v_1609;
assign v_1643 = v_669 & v_1609;
assign v_1644 = v_670 & v_1609;
assign v_1645 = v_675 & v_1610;
assign v_1646 = ~v_1645 & v_1641;
assign v_1647 = v_676 & v_1610;
assign v_1648 = ~v_1642 & ~v_1647;
assign v_1649 = v_677 & v_1610;
assign v_1650 = ~v_1643 & ~v_1649;
assign v_1651 = v_678 & v_1610;
assign v_1652 = ~v_1644 & ~v_1651;
assign v_1653 = v_679 & v_1611;
assign v_1654 = ~v_1653 & v_1646;
assign v_1655 = v_680 & v_1611;
assign v_1656 = ~v_1655 & v_1648;
assign v_1657 = v_681 & v_1611;
assign v_1658 = ~v_1657 & v_1650;
assign v_1659 = v_682 & v_1611;
assign v_1660 = ~v_1659 & v_1652;
assign v_1661 = v_683 & v_1612;
assign v_1662 = ~v_1661 & v_1654;
assign v_1663 = v_684 & v_1612;
assign v_1664 = ~v_1663 & v_1656;
assign v_1665 = v_685 & v_1612;
assign v_1666 = ~v_1665 & v_1658;
assign v_1667 = v_686 & v_1612;
assign v_1668 = ~v_1667 & v_1660;
assign v_1669 = v_687 & v_1613;
assign v_1670 = ~v_1669 & v_1662;
assign v_1671 = v_688 & v_1613;
assign v_1672 = ~v_1671 & v_1664;
assign v_1673 = v_689 & v_1613;
assign v_1674 = ~v_1673 & v_1666;
assign v_1675 = v_690 & v_1613;
assign v_1676 = ~v_1675 & v_1668;
assign v_1678 = ~v_1605 & v_1677;
assign v_1680 = ~v_1679 & v_494;
assign v_1681 = v_1040 & v_1680;
assign v_1682 = v_494 & v_495;
assign v_1683 = v_494 & v_496;
assign v_1684 = v_494 & v_497;
assign v_1685 = v_494 & v_498;
assign v_1686 = ~v_494 & v_1681;
assign v_1687 = ~v_1107 & v_1405;
assign v_1688 = v_1194 & v_1687;
assign v_1689 = ~v_1409 & ~v_1688;
assign v_1690 = ~v_1409 & v_1688;
assign v_1691 = ~v_1688 & v_1681;
assign v_1692 = v_687 & v_1688;
assign v_1693 = ~v_1692 & v_1688;
assign v_1694 = v_688 & v_1688;
assign v_1695 = v_689 & v_1688;
assign v_1696 = v_690 & v_1688;
assign v_1697 = v_675 & v_1682;
assign v_1698 = ~v_1697 & v_494;
assign v_1699 = v_676 & v_1682;
assign v_1700 = v_677 & v_1682;
assign v_1701 = v_678 & v_1682;
assign v_1702 = v_679 & v_1683;
assign v_1703 = ~v_1702 & v_1698;
assign v_1704 = v_680 & v_1683;
assign v_1705 = ~v_1699 & ~v_1704;
assign v_1706 = v_681 & v_1683;
assign v_1707 = ~v_1700 & ~v_1706;
assign v_1708 = v_682 & v_1683;
assign v_1709 = ~v_1701 & ~v_1708;
assign v_1710 = v_683 & v_1684;
assign v_1711 = ~v_1710 & v_1703;
assign v_1712 = v_684 & v_1684;
assign v_1713 = ~v_1712 & v_1705;
assign v_1714 = v_685 & v_1684;
assign v_1715 = ~v_1714 & v_1707;
assign v_1716 = v_686 & v_1684;
assign v_1717 = ~v_1716 & v_1709;
assign v_1718 = v_687 & v_1685;
assign v_1719 = ~v_1718 & v_1711;
assign v_1720 = v_688 & v_1685;
assign v_1721 = ~v_1720 & v_1713;
assign v_1722 = v_689 & v_1685;
assign v_1723 = ~v_1722 & v_1715;
assign v_1724 = v_690 & v_1685;
assign v_1725 = ~v_1724 & v_1717;
assign v_1727 = ~v_1679 & v_1726;
assign v_1729 = v_494 & v_1040;
assign v_1730 = ~v_1726 & v_1729;
assign v_1731 = v_963 & v_1040;
assign v_1732 = ~v_1677 & v_1731;
assign v_1733 = ~v_491 & v_1040;
assign v_1734 = ~v_1603 & v_1733;
assign v_1735 = ~v_1732 & ~v_1734;
assign v_1736 = ~v_1513 & v_1040;
assign v_1737 = ~v_1736 & v_1735;
assign v_1738 = ~v_1411 & v_1040;
assign v_1739 = ~v_1738 & v_1737;
assign v_1740 = ~v_1730 & v_1739;
assign v_1741 = v_1040 & v_1740;
assign v_1742 = ~v_1741 & v_1022;
assign v_1743 = v_504 & v_523;
assign v_1744 = ~v_1022 & v_491;
assign v_1748 = v_494 & v_1022;
assign v_1753 = v_4 & v_1748;
assign v_1754 = ~v_1749 & v_1743;
assign v_1755 = ~v_1749 & ~v_1750;
assign v_1756 = ~v_1751 & v_1755;
assign v_1757 = ~v_1749 & v_1754;
assign v_1758 = ~v_106 & v_1757;
assign v_1759 = v_107 & v_1758;
assign v_1760 = v_1749 & v_1759;
assign v_1761 = ~v_107 & v_1758;
assign v_1762 = v_1749 & v_1761;
assign v_1763 = ~v_171 & v_1757;
assign v_1764 = v_172 & v_1763;
assign v_1765 = v_1749 & v_1764;
assign v_1766 = ~v_172 & v_1763;
assign v_1767 = v_1749 & v_1766;
assign v_1768 = v_1743 & v_1755;
assign v_1769 = ~v_1750 & v_1755;
assign v_1771 = ~v_1749 & ~v_1770;
assign v_1773 = ~v_1772 & v_1768;
assign v_1774 = ~v_106 & v_1773;
assign v_1775 = v_107 & v_1774;
assign v_1776 = v_1772 & v_1775;
assign v_1777 = ~v_107 & v_1774;
assign v_1778 = v_1772 & v_1777;
assign v_1779 = ~v_171 & v_1773;
assign v_1780 = v_172 & v_1779;
assign v_1781 = v_1772 & v_1780;
assign v_1782 = ~v_172 & v_1779;
assign v_1783 = v_1772 & v_1782;
assign v_1784 = v_1743 & v_1756;
assign v_1785 = ~v_1751 & v_1756;
assign v_1787 = ~v_1750 & ~v_1786;
assign v_1789 = ~v_1749 & ~v_1788;
assign v_1791 = ~v_1790 & v_1784;
assign v_1792 = ~v_106 & v_1791;
assign v_1793 = v_107 & v_1792;
assign v_1794 = v_1790 & v_1793;
assign v_1795 = ~v_107 & v_1792;
assign v_1796 = v_1790 & v_1795;
assign v_1797 = ~v_171 & v_1791;
assign v_1798 = v_172 & v_1797;
assign v_1799 = v_1790 & v_1798;
assign v_1800 = ~v_172 & v_1797;
assign v_1801 = v_1790 & v_1800;
assign v_1802 = v_1743 & v_1753;
assign v_1803 = ~v_1752 & v_1753;
assign v_1805 = ~v_1751 & ~v_1804;
assign v_1807 = ~v_1750 & ~v_1806;
assign v_1809 = ~v_1749 & ~v_1808;
assign v_1811 = ~v_1810 & v_1802;
assign v_1812 = ~v_106 & v_1811;
assign v_1813 = v_107 & v_1812;
assign v_1814 = v_1810 & v_1813;
assign v_1815 = ~v_107 & v_1812;
assign v_1816 = v_1810 & v_1815;
assign v_1817 = ~v_171 & v_1811;
assign v_1818 = v_172 & v_1817;
assign v_1819 = v_1810 & v_1818;
assign v_1820 = ~v_172 & v_1817;
assign v_1821 = v_1810 & v_1820;
assign v_1822 = ~v_1810 & v_687;
assign v_1823 = ~v_1810 & ~v_1822;
assign v_1824 = ~v_1810 & v_688;
assign v_1825 = ~v_1810 & v_689;
assign v_1826 = ~v_1810 & v_690;
assign v_1827 = ~v_205 & ~v_1823;
assign v_1828 = v_589 & v_1824;
assign v_1829 = ~v_1827 & ~v_1828;
assign v_1830 = v_208 & v_1825;
assign v_1831 = ~v_1830 & v_1829;
assign v_1832 = v_211 & v_1823;
assign v_1833 = ~v_1824 & v_1823;
assign v_1834 = v_212 & v_1833;
assign v_1835 = ~v_1832 & ~v_1834;
assign v_1836 = v_213 & v_1826;
assign v_1837 = ~v_1836 & v_1835;
assign v_1838 = v_217 & v_1823;
assign v_1839 = v_218 & v_1833;
assign v_1840 = ~v_1838 & ~v_1839;
assign v_1841 = v_219 & v_1826;
assign v_1842 = ~v_1841 & v_1840;
assign v_1843 = ~v_223 & ~v_1823;
assign v_1844 = v_606 & v_1824;
assign v_1845 = ~v_1843 & ~v_1844;
assign v_1846 = v_226 & v_1825;
assign v_1847 = ~v_1846 & v_1845;
assign v_1850 = ~v_1837 & v_172;
assign v_1851 = v_173 & v_1842;
assign v_1852 = ~v_1847 & v_174;
assign v_1853 = v_175 & v_1848;
assign v_1854 = v_176 & v_1849;
assign v_1855 = v_177 & v_1831;
assign v_1858 = ~v_235 & ~v_1823;
assign v_1859 = v_628 & v_1824;
assign v_1860 = ~v_1858 & ~v_1859;
assign v_1861 = v_238 & v_1825;
assign v_1862 = ~v_1861 & v_1860;
assign v_1863 = v_241 & v_1823;
assign v_1864 = v_242 & v_1833;
assign v_1865 = ~v_1863 & ~v_1864;
assign v_1866 = v_243 & v_1826;
assign v_1867 = ~v_1866 & v_1865;
assign v_1868 = v_247 & v_1823;
assign v_1869 = v_248 & v_1833;
assign v_1870 = ~v_1868 & ~v_1869;
assign v_1871 = v_249 & v_1826;
assign v_1872 = ~v_1871 & v_1870;
assign v_1873 = ~v_253 & ~v_1823;
assign v_1874 = v_644 & v_1824;
assign v_1875 = ~v_1873 & ~v_1874;
assign v_1876 = v_256 & v_1825;
assign v_1877 = ~v_1876 & v_1875;
assign v_1879 = ~v_1867 & v_107;
assign v_1880 = v_108 & v_1872;
assign v_1881 = ~v_1877 & v_109;
assign v_1882 = v_110 & v_1878;
assign v_1883 = v_111 & v_1849;
assign v_1884 = v_112 & v_1862;
assign v_1887 = v_1857 & v_1886;
assign v_1888 = ~v_1810 & v_1887;
assign v_1889 = v_1753 & v_1888;
assign v_1890 = ~v_1790 & v_683;
assign v_1891 = ~v_1790 & ~v_1890;
assign v_1892 = ~v_1790 & v_684;
assign v_1893 = ~v_1790 & v_685;
assign v_1894 = ~v_1790 & v_686;
assign v_1895 = ~v_205 & ~v_1891;
assign v_1896 = v_589 & v_1892;
assign v_1897 = ~v_1895 & ~v_1896;
assign v_1898 = v_208 & v_1893;
assign v_1899 = ~v_1898 & v_1897;
assign v_1900 = v_211 & v_1891;
assign v_1901 = ~v_1892 & v_1891;
assign v_1902 = v_212 & v_1901;
assign v_1903 = ~v_1900 & ~v_1902;
assign v_1904 = v_213 & v_1894;
assign v_1905 = ~v_1904 & v_1903;
assign v_1906 = v_217 & v_1891;
assign v_1907 = v_218 & v_1901;
assign v_1908 = ~v_1906 & ~v_1907;
assign v_1909 = v_219 & v_1894;
assign v_1910 = ~v_1909 & v_1908;
assign v_1911 = ~v_223 & ~v_1891;
assign v_1912 = v_606 & v_1892;
assign v_1913 = ~v_1911 & ~v_1912;
assign v_1914 = v_226 & v_1893;
assign v_1915 = ~v_1914 & v_1913;
assign v_1918 = ~v_1905 & v_172;
assign v_1919 = v_173 & v_1910;
assign v_1920 = ~v_1915 & v_174;
assign v_1921 = v_175 & v_1916;
assign v_1922 = v_176 & v_1917;
assign v_1923 = v_177 & v_1899;
assign v_1926 = ~v_235 & ~v_1891;
assign v_1927 = v_628 & v_1892;
assign v_1928 = ~v_1926 & ~v_1927;
assign v_1929 = v_238 & v_1893;
assign v_1930 = ~v_1929 & v_1928;
assign v_1931 = v_241 & v_1891;
assign v_1932 = v_242 & v_1901;
assign v_1933 = ~v_1931 & ~v_1932;
assign v_1934 = v_243 & v_1894;
assign v_1935 = ~v_1934 & v_1933;
assign v_1936 = v_247 & v_1891;
assign v_1937 = v_248 & v_1901;
assign v_1938 = ~v_1936 & ~v_1937;
assign v_1939 = v_249 & v_1894;
assign v_1940 = ~v_1939 & v_1938;
assign v_1941 = ~v_253 & ~v_1891;
assign v_1942 = v_644 & v_1892;
assign v_1943 = ~v_1941 & ~v_1942;
assign v_1944 = v_256 & v_1893;
assign v_1945 = ~v_1944 & v_1943;
assign v_1947 = ~v_1935 & v_107;
assign v_1948 = v_108 & v_1940;
assign v_1949 = ~v_1945 & v_109;
assign v_1950 = v_110 & v_1946;
assign v_1951 = v_111 & v_1917;
assign v_1952 = v_112 & v_1930;
assign v_1955 = v_1925 & v_1954;
assign v_1956 = ~v_1790 & v_1955;
assign v_1957 = v_1756 & v_1956;
assign v_1958 = ~v_1772 & v_679;
assign v_1959 = ~v_1772 & ~v_1958;
assign v_1960 = ~v_1772 & v_680;
assign v_1961 = ~v_1772 & v_681;
assign v_1962 = ~v_1772 & v_682;
assign v_1963 = ~v_205 & ~v_1959;
assign v_1964 = v_589 & v_1960;
assign v_1965 = ~v_1963 & ~v_1964;
assign v_1966 = v_208 & v_1961;
assign v_1967 = ~v_1966 & v_1965;
assign v_1968 = v_211 & v_1959;
assign v_1969 = ~v_1960 & v_1959;
assign v_1970 = v_212 & v_1969;
assign v_1971 = ~v_1968 & ~v_1970;
assign v_1972 = v_213 & v_1962;
assign v_1973 = ~v_1972 & v_1971;
assign v_1974 = v_217 & v_1959;
assign v_1975 = v_218 & v_1969;
assign v_1976 = ~v_1974 & ~v_1975;
assign v_1977 = v_219 & v_1962;
assign v_1978 = ~v_1977 & v_1976;
assign v_1979 = ~v_223 & ~v_1959;
assign v_1980 = v_606 & v_1960;
assign v_1981 = ~v_1979 & ~v_1980;
assign v_1982 = v_226 & v_1961;
assign v_1983 = ~v_1982 & v_1981;
assign v_1986 = ~v_1973 & v_172;
assign v_1987 = v_173 & v_1978;
assign v_1988 = ~v_1983 & v_174;
assign v_1989 = v_175 & v_1984;
assign v_1990 = v_176 & v_1985;
assign v_1991 = v_177 & v_1967;
assign v_1994 = ~v_235 & ~v_1959;
assign v_1995 = v_628 & v_1960;
assign v_1996 = ~v_1994 & ~v_1995;
assign v_1997 = v_238 & v_1961;
assign v_1998 = ~v_1997 & v_1996;
assign v_1999 = v_241 & v_1959;
assign v_2000 = v_242 & v_1969;
assign v_2001 = ~v_1999 & ~v_2000;
assign v_2002 = v_243 & v_1962;
assign v_2003 = ~v_2002 & v_2001;
assign v_2004 = v_247 & v_1959;
assign v_2005 = v_248 & v_1969;
assign v_2006 = ~v_2004 & ~v_2005;
assign v_2007 = v_249 & v_1962;
assign v_2008 = ~v_2007 & v_2006;
assign v_2009 = ~v_253 & ~v_1959;
assign v_2010 = v_644 & v_1960;
assign v_2011 = ~v_2009 & ~v_2010;
assign v_2012 = v_256 & v_1961;
assign v_2013 = ~v_2012 & v_2011;
assign v_2015 = ~v_2003 & v_107;
assign v_2016 = v_108 & v_2008;
assign v_2017 = ~v_2013 & v_109;
assign v_2018 = v_110 & v_2014;
assign v_2019 = v_111 & v_1985;
assign v_2020 = v_112 & v_1998;
assign v_2023 = v_1993 & v_2022;
assign v_2024 = ~v_1772 & v_2023;
assign v_2025 = v_1755 & v_2024;
assign v_2026 = ~v_1749 & v_675;
assign v_2027 = ~v_1749 & ~v_2026;
assign v_2028 = ~v_1749 & v_676;
assign v_2029 = ~v_1749 & v_677;
assign v_2030 = ~v_1749 & v_678;
assign v_2031 = ~v_205 & ~v_2027;
assign v_2032 = v_589 & v_2028;
assign v_2033 = ~v_2031 & ~v_2032;
assign v_2034 = v_208 & v_2029;
assign v_2035 = ~v_2034 & v_2033;
assign v_2036 = v_211 & v_2027;
assign v_2037 = ~v_2028 & v_2027;
assign v_2038 = v_212 & v_2037;
assign v_2039 = ~v_2036 & ~v_2038;
assign v_2040 = v_213 & v_2030;
assign v_2041 = ~v_2040 & v_2039;
assign v_2042 = v_217 & v_2027;
assign v_2043 = v_218 & v_2037;
assign v_2044 = ~v_2042 & ~v_2043;
assign v_2045 = v_219 & v_2030;
assign v_2046 = ~v_2045 & v_2044;
assign v_2047 = ~v_223 & ~v_2027;
assign v_2048 = v_606 & v_2028;
assign v_2049 = ~v_2047 & ~v_2048;
assign v_2050 = v_226 & v_2029;
assign v_2051 = ~v_2050 & v_2049;
assign v_2054 = ~v_2041 & v_172;
assign v_2055 = v_173 & v_2046;
assign v_2056 = ~v_2051 & v_174;
assign v_2057 = v_175 & v_2052;
assign v_2058 = v_176 & v_2053;
assign v_2059 = v_177 & v_2035;
assign v_2062 = ~v_235 & ~v_2027;
assign v_2063 = v_628 & v_2028;
assign v_2064 = ~v_2062 & ~v_2063;
assign v_2065 = v_238 & v_2029;
assign v_2066 = ~v_2065 & v_2064;
assign v_2067 = v_241 & v_2027;
assign v_2068 = v_242 & v_2037;
assign v_2069 = ~v_2067 & ~v_2068;
assign v_2070 = v_243 & v_2030;
assign v_2071 = ~v_2070 & v_2069;
assign v_2072 = v_247 & v_2027;
assign v_2073 = v_248 & v_2037;
assign v_2074 = ~v_2072 & ~v_2073;
assign v_2075 = v_249 & v_2030;
assign v_2076 = ~v_2075 & v_2074;
assign v_2077 = ~v_253 & ~v_2027;
assign v_2078 = v_644 & v_2028;
assign v_2079 = ~v_2077 & ~v_2078;
assign v_2080 = v_256 & v_2029;
assign v_2081 = ~v_2080 & v_2079;
assign v_2083 = ~v_2071 & v_107;
assign v_2084 = v_108 & v_2076;
assign v_2085 = ~v_2081 & v_109;
assign v_2086 = v_110 & v_2082;
assign v_2087 = v_111 & v_2053;
assign v_2088 = v_112 & v_2066;
assign v_2091 = v_2061 & v_2090;
assign v_2092 = ~v_1749 & v_2091;
assign v_2093 = ~v_1749 & v_2092;
assign v_2094 = ~v_2025 & ~v_2093;
assign v_2096 = v_2025 & v_2093;
assign v_2097 = ~v_1957 & v_2094;
assign v_2100 = v_1957 & v_2096;
assign v_2101 = ~v_1889 & v_2097;
assign v_2105 = v_1889 & v_2100;
assign v_2107 = ~v_1744 & v_2106;
assign v_2108 = v_1743 & v_2107;
assign v_2109 = ~v_1749 & v_2093;
assign v_2111 = v_2093 & v_2109;
assign v_2112 = ~v_1772 & ~v_2093;
assign v_2115 = v_2025 & v_2112;
assign v_2117 = ~v_2094 & v_2114;
assign v_2118 = ~v_2094 & v_2115;
assign v_2119 = ~v_1790 & v_2094;
assign v_2123 = v_1957 & v_2119;
assign v_2125 = ~v_2097 & v_2121;
assign v_2126 = ~v_2097 & v_2122;
assign v_2127 = ~v_2097 & v_2123;
assign v_2128 = ~v_1810 & v_2097;
assign v_2133 = v_1889 & v_2128;
assign v_2134 = ~v_2101 & v_2129;
assign v_2135 = ~v_2101 & v_2130;
assign v_2136 = ~v_2101 & v_2131;
assign v_2137 = ~v_2101 & v_2132;
assign v_2138 = ~v_2101 & v_2133;
assign v_2139 = v_2108 & v_2129;
assign v_2140 = v_675 & v_2130;
assign v_2141 = ~v_2129 & ~v_2140;
assign v_2142 = v_676 & v_2130;
assign v_2143 = v_677 & v_2130;
assign v_2144 = v_678 & v_2130;
assign v_2145 = v_679 & v_2131;
assign v_2146 = ~v_2145 & v_2141;
assign v_2147 = v_680 & v_2131;
assign v_2148 = ~v_2142 & ~v_2147;
assign v_2149 = v_681 & v_2131;
assign v_2150 = ~v_2143 & ~v_2149;
assign v_2151 = v_682 & v_2131;
assign v_2152 = ~v_2144 & ~v_2151;
assign v_2153 = v_683 & v_2132;
assign v_2154 = ~v_2153 & v_2146;
assign v_2155 = v_684 & v_2132;
assign v_2156 = ~v_2155 & v_2148;
assign v_2157 = v_685 & v_2132;
assign v_2158 = ~v_2157 & v_2150;
assign v_2159 = v_686 & v_2132;
assign v_2160 = ~v_2159 & v_2152;
assign v_2161 = v_687 & v_2133;
assign v_2162 = ~v_2161 & v_2154;
assign v_2163 = v_688 & v_2133;
assign v_2164 = ~v_2163 & v_2156;
assign v_2165 = v_689 & v_2133;
assign v_2166 = ~v_2165 & v_2158;
assign v_2167 = v_690 & v_2133;
assign v_2168 = ~v_2167 & v_2160;
assign v_2170 = v_2106 & v_2169;
assign v_2172 = ~v_1744 & ~v_1745;
assign v_2173 = ~v_2171 & v_2172;
assign v_2174 = v_1743 & v_2173;
assign v_2175 = ~v_1772 & v_2093;
assign v_2176 = v_2025 & v_2175;
assign v_2178 = ~v_2095 & v_2176;
assign v_2179 = ~v_1790 & v_2095;
assign v_2182 = v_1957 & v_2179;
assign v_2184 = ~v_2098 & v_2181;
assign v_2185 = ~v_2098 & v_2182;
assign v_2186 = ~v_1810 & v_2098;
assign v_2190 = v_1889 & v_2186;
assign v_2191 = ~v_2102 & v_2187;
assign v_2192 = ~v_2102 & v_2188;
assign v_2193 = ~v_2102 & v_2189;
assign v_2194 = ~v_2102 & v_2190;
assign v_2195 = v_2174 & v_2187;
assign v_2196 = v_679 & v_2188;
assign v_2197 = ~v_2187 & ~v_2196;
assign v_2198 = v_680 & v_2188;
assign v_2199 = v_681 & v_2188;
assign v_2200 = v_682 & v_2188;
assign v_2201 = v_683 & v_2189;
assign v_2202 = ~v_2201 & v_2197;
assign v_2203 = v_684 & v_2189;
assign v_2204 = ~v_2198 & ~v_2203;
assign v_2205 = v_685 & v_2189;
assign v_2206 = ~v_2199 & ~v_2205;
assign v_2207 = v_686 & v_2189;
assign v_2208 = ~v_2200 & ~v_2207;
assign v_2209 = v_687 & v_2190;
assign v_2210 = ~v_2209 & v_2202;
assign v_2211 = v_688 & v_2190;
assign v_2212 = ~v_2211 & v_2204;
assign v_2213 = v_689 & v_2190;
assign v_2214 = ~v_2213 & v_2206;
assign v_2215 = v_690 & v_2190;
assign v_2216 = ~v_2215 & v_2208;
assign v_2218 = ~v_2171 & v_2217;
assign v_2220 = ~v_1746 & v_2172;
assign v_2221 = ~v_2219 & v_2220;
assign v_2222 = v_1743 & v_2221;
assign v_2223 = ~v_1790 & v_2096;
assign v_2224 = v_1957 & v_2223;
assign v_2226 = ~v_2099 & v_2224;
assign v_2227 = ~v_1810 & v_2099;
assign v_2230 = v_1889 & v_2227;
assign v_2231 = ~v_2103 & v_2228;
assign v_2232 = ~v_2103 & v_2229;
assign v_2233 = ~v_2103 & v_2230;
assign v_2234 = v_2222 & v_2228;
assign v_2235 = v_683 & v_2229;
assign v_2236 = ~v_2228 & ~v_2235;
assign v_2237 = v_684 & v_2229;
assign v_2238 = v_685 & v_2229;
assign v_2239 = v_686 & v_2229;
assign v_2240 = v_687 & v_2230;
assign v_2241 = ~v_2240 & v_2236;
assign v_2242 = v_688 & v_2230;
assign v_2243 = ~v_2237 & ~v_2242;
assign v_2244 = v_689 & v_2230;
assign v_2245 = ~v_2238 & ~v_2244;
assign v_2246 = v_690 & v_2230;
assign v_2247 = ~v_2239 & ~v_2246;
assign v_2249 = ~v_2219 & v_2248;
assign v_2251 = ~v_2250 & v_1748;
assign v_2252 = v_1743 & v_2251;
assign v_2253 = ~v_1810 & v_2100;
assign v_2254 = v_1889 & v_2253;
assign v_2255 = ~v_2104 & ~v_2254;
assign v_2256 = ~v_2104 & v_2254;
assign v_2257 = ~v_2254 & v_2252;
assign v_2258 = v_687 & v_2254;
assign v_2259 = ~v_2258 & v_2254;
assign v_2260 = v_688 & v_2254;
assign v_2261 = v_689 & v_2254;
assign v_2262 = v_690 & v_2254;
assign v_2264 = ~v_2250 & v_2263;
assign v_2266 = v_1743 & v_1748;
assign v_2267 = ~v_2263 & v_2266;
assign v_2268 = v_1743 & v_2220;
assign v_2269 = ~v_2248 & v_2268;
assign v_2270 = v_1743 & v_2172;
assign v_2271 = ~v_2217 & v_2270;
assign v_2272 = ~v_2269 & ~v_2271;
assign v_2273 = ~v_1744 & v_1743;
assign v_2274 = ~v_2169 & v_2273;
assign v_2275 = ~v_2274 & v_2272;
assign v_2276 = ~v_2106 & v_1743;
assign v_2277 = ~v_2276 & v_2275;
assign v_2278 = ~v_2267 & v_2277;
assign v_2279 = v_1743 & v_2278;
assign v_2281 = ~v_466 & ~v_467;
assign v_2282 = ~v_467 & v_466;
assign v_2283 = ~v_466 & v_467;
assign v_2284 = v_466 & v_467;
assign v_2285 = v_265 & v_1744;
assign v_2286 = v_265 & v_1745;
assign v_2287 = v_265 & v_1746;
assign v_2288 = v_265 & v_1747;
assign v_2289 = v_265 & v_1748;
assign v_2290 = v_266 & v_487;
assign v_2291 = v_266 & v_488;
assign v_2292 = v_266 & v_489;
assign v_2293 = v_266 & v_490;
assign v_2294 = v_267 & v_495;
assign v_2295 = v_267 & v_496;
assign v_2296 = v_267 & v_497;
assign v_2297 = v_267 & v_498;
assign v_2298 = v_268 & v_2281;
assign v_2299 = v_268 & v_2282;
assign v_2300 = v_268 & v_2283;
assign v_2301 = v_268 & v_2284;
assign v_2306 = ~v_2302 & v_2280;
assign v_2307 = ~v_2302 & ~v_2303;
assign v_2308 = ~v_2304 & v_2307;
assign v_2309 = ~v_2302 & v_2306;
assign v_2310 = ~v_302 & v_2309;
assign v_2311 = v_303 & v_2310;
assign v_2312 = v_2302 & v_2311;
assign v_2313 = ~v_303 & v_2310;
assign v_2314 = v_304 & v_2313;
assign v_2315 = v_2302 & v_2314;
assign v_2316 = ~v_304 & v_2313;
assign v_2317 = v_305 & v_2316;
assign v_2318 = v_2302 & v_2317;
assign v_2319 = ~v_305 & v_2316;
assign v_2320 = v_2302 & v_2319;
assign v_2321 = ~v_367 & v_2309;
assign v_2322 = v_368 & v_2321;
assign v_2323 = v_2302 & v_2322;
assign v_2324 = ~v_368 & v_2321;
assign v_2325 = v_369 & v_2324;
assign v_2326 = v_2302 & v_2325;
assign v_2327 = ~v_369 & v_2324;
assign v_2328 = v_370 & v_2327;
assign v_2329 = v_2302 & v_2328;
assign v_2330 = ~v_370 & v_2327;
assign v_2331 = v_2302 & v_2330;
assign v_2332 = v_2280 & v_2307;
assign v_2333 = ~v_2303 & v_2307;
assign v_2335 = ~v_2302 & ~v_2334;
assign v_2337 = ~v_2336 & v_2332;
assign v_2338 = ~v_302 & v_2337;
assign v_2339 = v_303 & v_2338;
assign v_2340 = v_2336 & v_2339;
assign v_2341 = ~v_303 & v_2338;
assign v_2342 = v_304 & v_2341;
assign v_2343 = v_2336 & v_2342;
assign v_2344 = ~v_304 & v_2341;
assign v_2345 = v_305 & v_2344;
assign v_2346 = v_2336 & v_2345;
assign v_2347 = ~v_305 & v_2344;
assign v_2348 = v_2336 & v_2347;
assign v_2349 = ~v_367 & v_2337;
assign v_2350 = v_368 & v_2349;
assign v_2351 = v_2336 & v_2350;
assign v_2352 = ~v_368 & v_2349;
assign v_2353 = v_369 & v_2352;
assign v_2354 = v_2336 & v_2353;
assign v_2355 = ~v_369 & v_2352;
assign v_2356 = v_370 & v_2355;
assign v_2357 = v_2336 & v_2356;
assign v_2358 = ~v_370 & v_2355;
assign v_2359 = v_2336 & v_2358;
assign v_2360 = v_2280 & v_2308;
assign v_2361 = ~v_2304 & v_2308;
assign v_2363 = ~v_2303 & ~v_2362;
assign v_2365 = ~v_2302 & ~v_2364;
assign v_2367 = ~v_2366 & v_2360;
assign v_2368 = ~v_302 & v_2367;
assign v_2369 = v_303 & v_2368;
assign v_2370 = v_2366 & v_2369;
assign v_2371 = ~v_303 & v_2368;
assign v_2372 = v_304 & v_2371;
assign v_2373 = v_2366 & v_2372;
assign v_2374 = ~v_304 & v_2371;
assign v_2375 = v_305 & v_2374;
assign v_2376 = v_2366 & v_2375;
assign v_2377 = ~v_305 & v_2374;
assign v_2378 = v_2366 & v_2377;
assign v_2379 = ~v_367 & v_2367;
assign v_2380 = v_368 & v_2379;
assign v_2381 = v_2366 & v_2380;
assign v_2382 = ~v_368 & v_2379;
assign v_2383 = v_369 & v_2382;
assign v_2384 = v_2366 & v_2383;
assign v_2385 = ~v_369 & v_2382;
assign v_2386 = v_370 & v_2385;
assign v_2387 = v_2366 & v_2386;
assign v_2388 = ~v_370 & v_2385;
assign v_2389 = v_2366 & v_2388;
assign v_2390 = v_2280 & v_2289;
assign v_2391 = ~v_2305 & v_2289;
assign v_2393 = ~v_2304 & ~v_2392;
assign v_2395 = ~v_2303 & ~v_2394;
assign v_2397 = ~v_2302 & ~v_2396;
assign v_2399 = ~v_2398 & v_2390;
assign v_2400 = ~v_302 & v_2399;
assign v_2401 = v_303 & v_2400;
assign v_2402 = v_2398 & v_2401;
assign v_2403 = ~v_303 & v_2400;
assign v_2404 = v_304 & v_2403;
assign v_2405 = v_2398 & v_2404;
assign v_2406 = ~v_304 & v_2403;
assign v_2407 = v_305 & v_2406;
assign v_2408 = v_2398 & v_2407;
assign v_2409 = ~v_305 & v_2406;
assign v_2410 = v_2398 & v_2409;
assign v_2411 = ~v_367 & v_2399;
assign v_2412 = v_368 & v_2411;
assign v_2413 = v_2398 & v_2412;
assign v_2414 = ~v_368 & v_2411;
assign v_2415 = v_369 & v_2414;
assign v_2416 = v_2398 & v_2415;
assign v_2417 = ~v_369 & v_2414;
assign v_2418 = v_370 & v_2417;
assign v_2419 = v_2398 & v_2418;
assign v_2420 = ~v_370 & v_2417;
assign v_2421 = v_2398 & v_2420;
assign v_2422 = ~v_367 & ~v_368;
assign v_2423 = ~v_369 & v_2422;
assign v_2424 = ~v_370 & v_2423;
assign v_2425 = ~v_371 & v_2424;
assign v_2426 = ~v_372 & v_2425;
assign v_2427 = ~v_373 & v_2426;
assign v_2428 = ~v_374 & v_2427;
assign v_2429 = ~v_375 & v_2428;
assign v_2430 = ~v_401 & v_584;
assign v_2431 = ~v_401 & ~v_402;
assign v_2432 = v_585 & v_2431;
assign v_2433 = ~v_2430 & ~v_2432;
assign v_2434 = v_404 & v_586;
assign v_2435 = ~v_2434 & v_2433;
assign v_2436 = ~v_584 & v_407;
assign v_2437 = v_408 & v_595;
assign v_2438 = ~v_2436 & ~v_2437;
assign v_2439 = v_409 & v_587;
assign v_2440 = ~v_2439 & v_2438;
assign v_2441 = ~v_584 & v_413;
assign v_2442 = v_414 & v_595;
assign v_2443 = ~v_2441 & ~v_2442;
assign v_2444 = v_415 & v_587;
assign v_2445 = ~v_2444 & v_2443;
assign v_2446 = ~v_419 & v_584;
assign v_2447 = ~v_419 & ~v_420;
assign v_2448 = v_585 & v_2447;
assign v_2449 = ~v_2446 & ~v_2448;
assign v_2450 = v_422 & v_586;
assign v_2451 = ~v_2450 & v_2449;
assign v_2454 = ~v_2440 & v_368;
assign v_2455 = v_369 & v_2445;
assign v_2456 = ~v_2451 & v_370;
assign v_2457 = v_371 & v_2452;
assign v_2458 = v_372 & v_612;
assign v_2459 = v_373 & v_2453;
assign v_2460 = v_375 & v_2435;
assign v_2463 = ~v_302 & ~v_303;
assign v_2464 = ~v_304 & v_2463;
assign v_2465 = ~v_305 & v_2464;
assign v_2466 = ~v_306 & v_2465;
assign v_2467 = ~v_307 & v_2466;
assign v_2468 = ~v_308 & v_2467;
assign v_2469 = ~v_309 & v_2468;
assign v_2470 = ~v_310 & v_2469;
assign v_2471 = ~v_431 & v_584;
assign v_2472 = ~v_431 & ~v_432;
assign v_2473 = v_585 & v_2472;
assign v_2474 = ~v_2471 & ~v_2473;
assign v_2475 = v_434 & v_586;
assign v_2476 = ~v_2475 & v_2474;
assign v_2477 = ~v_584 & v_437;
assign v_2478 = v_438 & v_595;
assign v_2479 = ~v_2477 & ~v_2478;
assign v_2480 = v_439 & v_587;
assign v_2481 = ~v_2480 & v_2479;
assign v_2482 = ~v_584 & v_443;
assign v_2483 = v_444 & v_595;
assign v_2484 = ~v_2482 & ~v_2483;
assign v_2485 = v_445 & v_587;
assign v_2486 = ~v_2485 & v_2484;
assign v_2487 = ~v_449 & v_584;
assign v_2488 = ~v_449 & ~v_450;
assign v_2489 = v_585 & v_2488;
assign v_2490 = ~v_2487 & ~v_2489;
assign v_2491 = v_452 & v_586;
assign v_2492 = ~v_2491 & v_2490;
assign v_2494 = ~v_2481 & v_303;
assign v_2495 = v_304 & v_2486;
assign v_2496 = ~v_2492 & v_305;
assign v_2497 = v_306 & v_2493;
assign v_2498 = v_307 & v_612;
assign v_2499 = v_308 & v_2453;
assign v_2500 = v_310 & v_2476;
assign v_2503 = v_2462 & v_2502;
assign v_2504 = ~v_2398 & v_687;
assign v_2505 = ~v_2398 & ~v_2504;
assign v_2506 = ~v_2398 & v_688;
assign v_2507 = ~v_2398 & v_689;
assign v_2508 = ~v_2398 & v_690;
assign v_2509 = ~v_401 & ~v_2505;
assign v_2510 = v_2431 & v_2506;
assign v_2511 = ~v_2509 & ~v_2510;
assign v_2512 = v_404 & v_2507;
assign v_2513 = ~v_2512 & v_2511;
assign v_2514 = v_407 & v_2505;
assign v_2515 = ~v_2506 & v_2505;
assign v_2516 = v_408 & v_2515;
assign v_2517 = ~v_2514 & ~v_2516;
assign v_2518 = v_409 & v_2508;
assign v_2519 = ~v_2518 & v_2517;
assign v_2520 = v_413 & v_2505;
assign v_2521 = v_414 & v_2515;
assign v_2522 = ~v_2520 & ~v_2521;
assign v_2523 = v_415 & v_2508;
assign v_2524 = ~v_2523 & v_2522;
assign v_2525 = ~v_419 & ~v_2505;
assign v_2526 = v_2447 & v_2506;
assign v_2527 = ~v_2525 & ~v_2526;
assign v_2528 = v_422 & v_2507;
assign v_2529 = ~v_2528 & v_2527;
assign v_2534 = ~v_2519 & v_368;
assign v_2535 = v_369 & v_2524;
assign v_2536 = ~v_2529 & v_370;
assign v_2537 = v_371 & v_2530;
assign v_2538 = v_372 & v_2531;
assign v_2539 = v_373 & v_2532;
assign v_2540 = v_374 & v_2533;
assign v_2541 = v_375 & v_2513;
assign v_2544 = ~v_431 & ~v_2505;
assign v_2545 = v_2472 & v_2506;
assign v_2546 = ~v_2544 & ~v_2545;
assign v_2547 = v_434 & v_2507;
assign v_2548 = ~v_2547 & v_2546;
assign v_2549 = v_437 & v_2505;
assign v_2550 = v_438 & v_2515;
assign v_2551 = ~v_2549 & ~v_2550;
assign v_2552 = v_439 & v_2508;
assign v_2553 = ~v_2552 & v_2551;
assign v_2554 = v_443 & v_2505;
assign v_2555 = v_444 & v_2515;
assign v_2556 = ~v_2554 & ~v_2555;
assign v_2557 = v_445 & v_2508;
assign v_2558 = ~v_2557 & v_2556;
assign v_2559 = ~v_449 & ~v_2505;
assign v_2560 = v_2488 & v_2506;
assign v_2561 = ~v_2559 & ~v_2560;
assign v_2562 = v_452 & v_2507;
assign v_2563 = ~v_2562 & v_2561;
assign v_2565 = ~v_2553 & v_303;
assign v_2566 = v_304 & v_2558;
assign v_2567 = ~v_2563 & v_305;
assign v_2568 = v_306 & v_2564;
assign v_2569 = v_307 & v_2531;
assign v_2570 = v_308 & v_2532;
assign v_2571 = v_309 & v_2533;
assign v_2572 = v_310 & v_2548;
assign v_2575 = v_2543 & v_2574;
assign v_2576 = ~v_2398 & v_2575;
assign v_2577 = v_2289 & v_2576;
assign v_2578 = ~v_2366 & v_683;
assign v_2579 = ~v_2366 & ~v_2578;
assign v_2580 = ~v_2366 & v_684;
assign v_2581 = ~v_2366 & v_685;
assign v_2582 = ~v_2366 & v_686;
assign v_2583 = ~v_401 & ~v_2579;
assign v_2584 = v_2431 & v_2580;
assign v_2585 = ~v_2583 & ~v_2584;
assign v_2586 = v_404 & v_2581;
assign v_2587 = ~v_2586 & v_2585;
assign v_2588 = v_407 & v_2579;
assign v_2589 = ~v_2580 & v_2579;
assign v_2590 = v_408 & v_2589;
assign v_2591 = ~v_2588 & ~v_2590;
assign v_2592 = v_409 & v_2582;
assign v_2593 = ~v_2592 & v_2591;
assign v_2594 = v_413 & v_2579;
assign v_2595 = v_414 & v_2589;
assign v_2596 = ~v_2594 & ~v_2595;
assign v_2597 = v_415 & v_2582;
assign v_2598 = ~v_2597 & v_2596;
assign v_2599 = ~v_419 & ~v_2579;
assign v_2600 = v_2447 & v_2580;
assign v_2601 = ~v_2599 & ~v_2600;
assign v_2602 = v_422 & v_2581;
assign v_2603 = ~v_2602 & v_2601;
assign v_2608 = ~v_2593 & v_368;
assign v_2609 = v_369 & v_2598;
assign v_2610 = ~v_2603 & v_370;
assign v_2611 = v_371 & v_2604;
assign v_2612 = v_372 & v_2605;
assign v_2613 = v_373 & v_2606;
assign v_2614 = v_374 & v_2607;
assign v_2615 = v_375 & v_2587;
assign v_2618 = ~v_431 & ~v_2579;
assign v_2619 = v_2472 & v_2580;
assign v_2620 = ~v_2618 & ~v_2619;
assign v_2621 = v_434 & v_2581;
assign v_2622 = ~v_2621 & v_2620;
assign v_2623 = v_437 & v_2579;
assign v_2624 = v_438 & v_2589;
assign v_2625 = ~v_2623 & ~v_2624;
assign v_2626 = v_439 & v_2582;
assign v_2627 = ~v_2626 & v_2625;
assign v_2628 = v_443 & v_2579;
assign v_2629 = v_444 & v_2589;
assign v_2630 = ~v_2628 & ~v_2629;
assign v_2631 = v_445 & v_2582;
assign v_2632 = ~v_2631 & v_2630;
assign v_2633 = ~v_449 & ~v_2579;
assign v_2634 = v_2488 & v_2580;
assign v_2635 = ~v_2633 & ~v_2634;
assign v_2636 = v_452 & v_2581;
assign v_2637 = ~v_2636 & v_2635;
assign v_2639 = ~v_2627 & v_303;
assign v_2640 = v_304 & v_2632;
assign v_2641 = ~v_2637 & v_305;
assign v_2642 = v_306 & v_2638;
assign v_2643 = v_307 & v_2605;
assign v_2644 = v_308 & v_2606;
assign v_2645 = v_309 & v_2607;
assign v_2646 = v_310 & v_2622;
assign v_2649 = v_2617 & v_2648;
assign v_2650 = ~v_2366 & v_2649;
assign v_2651 = v_2308 & v_2650;
assign v_2652 = ~v_2336 & v_679;
assign v_2653 = ~v_2336 & ~v_2652;
assign v_2654 = ~v_2336 & v_680;
assign v_2655 = ~v_2336 & v_681;
assign v_2656 = ~v_2336 & v_682;
assign v_2657 = ~v_401 & ~v_2653;
assign v_2658 = v_2431 & v_2654;
assign v_2659 = ~v_2657 & ~v_2658;
assign v_2660 = v_404 & v_2655;
assign v_2661 = ~v_2660 & v_2659;
assign v_2662 = v_407 & v_2653;
assign v_2663 = ~v_2654 & v_2653;
assign v_2664 = v_408 & v_2663;
assign v_2665 = ~v_2662 & ~v_2664;
assign v_2666 = v_409 & v_2656;
assign v_2667 = ~v_2666 & v_2665;
assign v_2668 = v_413 & v_2653;
assign v_2669 = v_414 & v_2663;
assign v_2670 = ~v_2668 & ~v_2669;
assign v_2671 = v_415 & v_2656;
assign v_2672 = ~v_2671 & v_2670;
assign v_2673 = ~v_419 & ~v_2653;
assign v_2674 = v_2447 & v_2654;
assign v_2675 = ~v_2673 & ~v_2674;
assign v_2676 = v_422 & v_2655;
assign v_2677 = ~v_2676 & v_2675;
assign v_2682 = ~v_2667 & v_368;
assign v_2683 = v_369 & v_2672;
assign v_2684 = ~v_2677 & v_370;
assign v_2685 = v_371 & v_2678;
assign v_2686 = v_372 & v_2679;
assign v_2687 = v_373 & v_2680;
assign v_2688 = v_374 & v_2681;
assign v_2689 = v_375 & v_2661;
assign v_2692 = ~v_431 & ~v_2653;
assign v_2693 = v_2472 & v_2654;
assign v_2694 = ~v_2692 & ~v_2693;
assign v_2695 = v_434 & v_2655;
assign v_2696 = ~v_2695 & v_2694;
assign v_2697 = v_437 & v_2653;
assign v_2698 = v_438 & v_2663;
assign v_2699 = ~v_2697 & ~v_2698;
assign v_2700 = v_439 & v_2656;
assign v_2701 = ~v_2700 & v_2699;
assign v_2702 = v_443 & v_2653;
assign v_2703 = v_444 & v_2663;
assign v_2704 = ~v_2702 & ~v_2703;
assign v_2705 = v_445 & v_2656;
assign v_2706 = ~v_2705 & v_2704;
assign v_2707 = ~v_449 & ~v_2653;
assign v_2708 = v_2488 & v_2654;
assign v_2709 = ~v_2707 & ~v_2708;
assign v_2710 = v_452 & v_2655;
assign v_2711 = ~v_2710 & v_2709;
assign v_2713 = ~v_2701 & v_303;
assign v_2714 = v_304 & v_2706;
assign v_2715 = ~v_2711 & v_305;
assign v_2716 = v_306 & v_2712;
assign v_2717 = v_307 & v_2679;
assign v_2718 = v_308 & v_2680;
assign v_2719 = v_309 & v_2681;
assign v_2720 = v_310 & v_2696;
assign v_2723 = v_2691 & v_2722;
assign v_2724 = ~v_2336 & v_2723;
assign v_2725 = v_2307 & v_2724;
assign v_2726 = ~v_2302 & v_675;
assign v_2727 = ~v_2302 & ~v_2726;
assign v_2728 = ~v_2302 & v_676;
assign v_2729 = ~v_2302 & v_677;
assign v_2730 = ~v_2302 & v_678;
assign v_2731 = ~v_401 & ~v_2727;
assign v_2732 = v_2431 & v_2728;
assign v_2733 = ~v_2731 & ~v_2732;
assign v_2734 = v_404 & v_2729;
assign v_2735 = ~v_2734 & v_2733;
assign v_2736 = v_407 & v_2727;
assign v_2737 = ~v_2728 & v_2727;
assign v_2738 = v_408 & v_2737;
assign v_2739 = ~v_2736 & ~v_2738;
assign v_2740 = v_409 & v_2730;
assign v_2741 = ~v_2740 & v_2739;
assign v_2742 = v_413 & v_2727;
assign v_2743 = v_414 & v_2737;
assign v_2744 = ~v_2742 & ~v_2743;
assign v_2745 = v_415 & v_2730;
assign v_2746 = ~v_2745 & v_2744;
assign v_2747 = ~v_419 & ~v_2727;
assign v_2748 = v_2447 & v_2728;
assign v_2749 = ~v_2747 & ~v_2748;
assign v_2750 = v_422 & v_2729;
assign v_2751 = ~v_2750 & v_2749;
assign v_2756 = ~v_2741 & v_368;
assign v_2757 = v_369 & v_2746;
assign v_2758 = ~v_2751 & v_370;
assign v_2759 = v_371 & v_2752;
assign v_2760 = v_372 & v_2753;
assign v_2761 = v_373 & v_2754;
assign v_2762 = v_374 & v_2755;
assign v_2763 = v_375 & v_2735;
assign v_2766 = ~v_431 & ~v_2727;
assign v_2767 = v_2472 & v_2728;
assign v_2768 = ~v_2766 & ~v_2767;
assign v_2769 = v_434 & v_2729;
assign v_2770 = ~v_2769 & v_2768;
assign v_2771 = v_437 & v_2727;
assign v_2772 = v_438 & v_2737;
assign v_2773 = ~v_2771 & ~v_2772;
assign v_2774 = v_439 & v_2730;
assign v_2775 = ~v_2774 & v_2773;
assign v_2776 = v_443 & v_2727;
assign v_2777 = v_444 & v_2737;
assign v_2778 = ~v_2776 & ~v_2777;
assign v_2779 = v_445 & v_2730;
assign v_2780 = ~v_2779 & v_2778;
assign v_2781 = ~v_449 & ~v_2727;
assign v_2782 = v_2488 & v_2728;
assign v_2783 = ~v_2781 & ~v_2782;
assign v_2784 = v_452 & v_2729;
assign v_2785 = ~v_2784 & v_2783;
assign v_2787 = ~v_2775 & v_303;
assign v_2788 = v_304 & v_2780;
assign v_2789 = ~v_2785 & v_305;
assign v_2790 = v_306 & v_2786;
assign v_2791 = v_307 & v_2753;
assign v_2792 = v_308 & v_2754;
assign v_2793 = v_309 & v_2755;
assign v_2794 = v_310 & v_2770;
assign v_2797 = v_2765 & v_2796;
assign v_2798 = ~v_2302 & v_2797;
assign v_2799 = ~v_2302 & v_2798;
assign v_2800 = ~v_2725 & ~v_2799;
assign v_2802 = v_2725 & v_2799;
assign v_2803 = ~v_2651 & v_2800;
assign v_2806 = v_2651 & v_2802;
assign v_2807 = ~v_2577 & v_2803;
assign v_2811 = v_2577 & v_2806;
assign v_2813 = ~v_1744 & v_2812;
assign v_2814 = v_2280 & v_2813;
assign v_2815 = ~v_2302 & v_2799;
assign v_2817 = v_2799 & v_2815;
assign v_2818 = ~v_2336 & ~v_2799;
assign v_2821 = v_2725 & v_2818;
assign v_2823 = ~v_2800 & v_2820;
assign v_2824 = ~v_2800 & v_2821;
assign v_2825 = ~v_2366 & v_2800;
assign v_2829 = v_2651 & v_2825;
assign v_2831 = ~v_2803 & v_2827;
assign v_2832 = ~v_2803 & v_2828;
assign v_2833 = ~v_2803 & v_2829;
assign v_2834 = ~v_2398 & v_2803;
assign v_2839 = v_2577 & v_2834;
assign v_2840 = ~v_2807 & v_2835;
assign v_2841 = ~v_2807 & v_2836;
assign v_2842 = ~v_2807 & v_2837;
assign v_2843 = ~v_2807 & v_2838;
assign v_2844 = ~v_2807 & v_2839;
assign v_2845 = v_2814 & v_2835;
assign v_2846 = v_675 & v_2836;
assign v_2847 = ~v_2835 & ~v_2846;
assign v_2848 = v_676 & v_2836;
assign v_2849 = v_677 & v_2836;
assign v_2850 = v_678 & v_2836;
assign v_2851 = v_679 & v_2837;
assign v_2852 = ~v_2851 & v_2847;
assign v_2853 = v_680 & v_2837;
assign v_2854 = ~v_2848 & ~v_2853;
assign v_2855 = v_681 & v_2837;
assign v_2856 = ~v_2849 & ~v_2855;
assign v_2857 = v_682 & v_2837;
assign v_2858 = ~v_2850 & ~v_2857;
assign v_2859 = v_683 & v_2838;
assign v_2860 = ~v_2859 & v_2852;
assign v_2861 = v_684 & v_2838;
assign v_2862 = ~v_2861 & v_2854;
assign v_2863 = v_685 & v_2838;
assign v_2864 = ~v_2863 & v_2856;
assign v_2865 = v_686 & v_2838;
assign v_2866 = ~v_2865 & v_2858;
assign v_2867 = v_687 & v_2839;
assign v_2868 = ~v_2867 & v_2860;
assign v_2869 = v_688 & v_2839;
assign v_2870 = ~v_2869 & v_2862;
assign v_2871 = v_689 & v_2839;
assign v_2872 = ~v_2871 & v_2864;
assign v_2873 = v_690 & v_2839;
assign v_2874 = ~v_2873 & v_2866;
assign v_2876 = v_2812 & v_2875;
assign v_2878 = ~v_2877 & v_2172;
assign v_2879 = v_2280 & v_2878;
assign v_2880 = ~v_2336 & v_2799;
assign v_2881 = v_2725 & v_2880;
assign v_2883 = ~v_2801 & v_2881;
assign v_2884 = ~v_2366 & v_2801;
assign v_2887 = v_2651 & v_2884;
assign v_2889 = ~v_2804 & v_2886;
assign v_2890 = ~v_2804 & v_2887;
assign v_2891 = ~v_2398 & v_2804;
assign v_2895 = v_2577 & v_2891;
assign v_2896 = ~v_2808 & v_2892;
assign v_2897 = ~v_2808 & v_2893;
assign v_2898 = ~v_2808 & v_2894;
assign v_2899 = ~v_2808 & v_2895;
assign v_2900 = v_2879 & v_2892;
assign v_2901 = v_679 & v_2893;
assign v_2902 = ~v_2892 & ~v_2901;
assign v_2903 = v_680 & v_2893;
assign v_2904 = v_681 & v_2893;
assign v_2905 = v_682 & v_2893;
assign v_2906 = v_683 & v_2894;
assign v_2907 = ~v_2906 & v_2902;
assign v_2908 = v_684 & v_2894;
assign v_2909 = ~v_2903 & ~v_2908;
assign v_2910 = v_685 & v_2894;
assign v_2911 = ~v_2904 & ~v_2910;
assign v_2912 = v_686 & v_2894;
assign v_2913 = ~v_2905 & ~v_2912;
assign v_2914 = v_687 & v_2895;
assign v_2915 = ~v_2914 & v_2907;
assign v_2916 = v_688 & v_2895;
assign v_2917 = ~v_2916 & v_2909;
assign v_2918 = v_689 & v_2895;
assign v_2919 = ~v_2918 & v_2911;
assign v_2920 = v_690 & v_2895;
assign v_2921 = ~v_2920 & v_2913;
assign v_2923 = ~v_2877 & v_2922;
assign v_2925 = ~v_2924 & v_2220;
assign v_2926 = v_2280 & v_2925;
assign v_2927 = ~v_2366 & v_2802;
assign v_2928 = v_2651 & v_2927;
assign v_2930 = ~v_2805 & v_2928;
assign v_2931 = ~v_2398 & v_2805;
assign v_2934 = v_2577 & v_2931;
assign v_2935 = ~v_2809 & v_2932;
assign v_2936 = ~v_2809 & v_2933;
assign v_2937 = ~v_2809 & v_2934;
assign v_2938 = v_2926 & v_2932;
assign v_2939 = v_683 & v_2933;
assign v_2940 = ~v_2932 & ~v_2939;
assign v_2941 = v_684 & v_2933;
assign v_2942 = v_685 & v_2933;
assign v_2943 = v_686 & v_2933;
assign v_2944 = v_687 & v_2934;
assign v_2945 = ~v_2944 & v_2940;
assign v_2946 = v_688 & v_2934;
assign v_2947 = ~v_2941 & ~v_2946;
assign v_2948 = v_689 & v_2934;
assign v_2949 = ~v_2942 & ~v_2948;
assign v_2950 = v_690 & v_2934;
assign v_2951 = ~v_2943 & ~v_2950;
assign v_2953 = ~v_2924 & v_2952;
assign v_2955 = ~v_2954 & v_1748;
assign v_2956 = v_2280 & v_2955;
assign v_2957 = ~v_2398 & v_2806;
assign v_2958 = v_2577 & v_2957;
assign v_2959 = ~v_2810 & ~v_2958;
assign v_2960 = ~v_2810 & v_2958;
assign v_2961 = ~v_2958 & v_2956;
assign v_2962 = v_687 & v_2958;
assign v_2963 = ~v_2962 & v_2958;
assign v_2964 = v_688 & v_2958;
assign v_2965 = v_689 & v_2958;
assign v_2966 = v_690 & v_2958;
assign v_2968 = ~v_2954 & v_2967;
assign v_2970 = v_1748 & v_2280;
assign v_2971 = ~v_2967 & v_2970;
assign v_2972 = v_2220 & v_2280;
assign v_2973 = ~v_2952 & v_2972;
assign v_2974 = v_2172 & v_2280;
assign v_2975 = ~v_2922 & v_2974;
assign v_2976 = ~v_2973 & ~v_2975;
assign v_2977 = ~v_1744 & v_2280;
assign v_2978 = ~v_2875 & v_2977;
assign v_2979 = ~v_2978 & v_2976;
assign v_2980 = ~v_2812 & v_2280;
assign v_2981 = ~v_2980 & v_2979;
assign v_2982 = ~v_2971 & v_2981;
assign v_2983 = ~v_2982 & v_2280;
assign v_2984 = ~v_487 & v_44;
assign v_2985 = v_45 & v_487;
assign v_2986 = v_46 & v_487;
assign v_2989 = ~v_487 & v_5;
assign v_2990 = v_5 & v_488;
assign v_2991 = v_5 & v_489;
assign v_2992 = v_5 & v_490;
assign v_2993 = ~v_4 & v_2989;
assign v_2994 = ~v_4 & v_2990;
assign v_2995 = ~v_4 & v_2991;
assign v_2996 = ~v_4 & v_2992;
assign v_2997 = v_2988 & v_2993;
assign v_2998 = ~v_2994 & v_2993;
assign v_2999 = v_2993 & v_2997;
assign v_3000 = ~v_106 & v_2999;
assign v_3001 = v_107 & v_3000;
assign v_3002 = ~v_2993 & v_3001;
assign v_3003 = ~v_107 & v_3000;
assign v_3004 = ~v_2993 & v_3003;
assign v_3005 = ~v_171 & v_2999;
assign v_3006 = v_172 & v_3005;
assign v_3007 = ~v_2993 & v_3006;
assign v_3008 = ~v_172 & v_3005;
assign v_3009 = ~v_2993 & v_3008;
assign v_3010 = v_2988 & v_2998;
assign v_3011 = ~v_2994 & v_2998;
assign v_3012 = v_2993 & v_3011;
assign v_3014 = ~v_3013 & v_3010;
assign v_3015 = ~v_106 & v_3014;
assign v_3016 = v_107 & v_3015;
assign v_3017 = v_3013 & v_3016;
assign v_3018 = ~v_107 & v_3015;
assign v_3019 = v_3013 & v_3018;
assign v_3020 = ~v_171 & v_3014;
assign v_3021 = v_172 & v_3020;
assign v_3022 = v_3013 & v_3021;
assign v_3023 = ~v_172 & v_3020;
assign v_3024 = v_3013 & v_3023;
assign v_3025 = v_2988 & v_2996;
assign v_3026 = ~v_2995 & v_2996;
assign v_3027 = ~v_2994 & v_3026;
assign v_3029 = ~v_3028 & v_2993;
assign v_3031 = ~v_3030 & v_3025;
assign v_3032 = ~v_106 & v_3031;
assign v_3033 = v_107 & v_3032;
assign v_3034 = v_3030 & v_3033;
assign v_3035 = ~v_107 & v_3032;
assign v_3036 = v_3030 & v_3035;
assign v_3037 = ~v_171 & v_3031;
assign v_3038 = v_172 & v_3037;
assign v_3039 = v_3030 & v_3038;
assign v_3040 = ~v_172 & v_3037;
assign v_3041 = v_3030 & v_3040;
assign v_3042 = v_176 & v_584;
assign v_3045 = v_111 & v_584;
assign v_3048 = v_3044 & v_3047;
assign v_3053 = v_3050 & v_3052;
assign v_3054 = ~v_3030 & v_683;
assign v_3055 = ~v_3030 & ~v_3054;
assign v_3056 = ~v_3030 & v_684;
assign v_3057 = ~v_3030 & v_685;
assign v_3058 = ~v_3030 & v_686;
assign v_3059 = ~v_205 & ~v_3055;
assign v_3060 = v_589 & v_3056;
assign v_3061 = ~v_3059 & ~v_3060;
assign v_3062 = v_208 & v_3057;
assign v_3063 = ~v_3062 & v_3061;
assign v_3064 = v_211 & v_3055;
assign v_3065 = ~v_3056 & v_3055;
assign v_3066 = v_212 & v_3065;
assign v_3067 = ~v_3064 & ~v_3066;
assign v_3068 = v_213 & v_3058;
assign v_3069 = ~v_3068 & v_3067;
assign v_3070 = v_217 & v_3055;
assign v_3071 = v_218 & v_3065;
assign v_3072 = ~v_3070 & ~v_3071;
assign v_3073 = v_219 & v_3058;
assign v_3074 = ~v_3073 & v_3072;
assign v_3075 = ~v_223 & ~v_3055;
assign v_3076 = v_606 & v_3056;
assign v_3077 = ~v_3075 & ~v_3076;
assign v_3078 = v_226 & v_3057;
assign v_3079 = ~v_3078 & v_3077;
assign v_3081 = ~v_3069 & v_172;
assign v_3082 = v_173 & v_3074;
assign v_3083 = ~v_3079 & v_174;
assign v_3084 = v_175 & v_3080;
assign v_3085 = ~v_3055 & v_176;
assign v_3086 = v_177 & v_3063;
assign v_3089 = ~v_235 & ~v_3055;
assign v_3090 = v_628 & v_3056;
assign v_3091 = ~v_3089 & ~v_3090;
assign v_3092 = v_238 & v_3057;
assign v_3093 = ~v_3092 & v_3091;
assign v_3094 = v_241 & v_3055;
assign v_3095 = v_242 & v_3065;
assign v_3096 = ~v_3094 & ~v_3095;
assign v_3097 = v_243 & v_3058;
assign v_3098 = ~v_3097 & v_3096;
assign v_3099 = v_247 & v_3055;
assign v_3100 = v_248 & v_3065;
assign v_3101 = ~v_3099 & ~v_3100;
assign v_3102 = v_249 & v_3058;
assign v_3103 = ~v_3102 & v_3101;
assign v_3104 = ~v_253 & ~v_3055;
assign v_3105 = v_644 & v_3056;
assign v_3106 = ~v_3104 & ~v_3105;
assign v_3107 = v_256 & v_3057;
assign v_3108 = ~v_3107 & v_3106;
assign v_3110 = ~v_3098 & v_107;
assign v_3111 = v_108 & v_3103;
assign v_3112 = ~v_3108 & v_109;
assign v_3113 = v_110 & v_3109;
assign v_3114 = ~v_3055 & v_111;
assign v_3115 = v_112 & v_3093;
assign v_3118 = v_3088 & v_3117;
assign v_3119 = ~v_3030 & v_3118;
assign v_3120 = v_2996 & v_3119;
assign v_3121 = ~v_3013 & v_679;
assign v_3122 = ~v_3013 & ~v_3121;
assign v_3123 = ~v_3013 & v_680;
assign v_3124 = ~v_3013 & v_681;
assign v_3125 = ~v_3013 & v_682;
assign v_3126 = ~v_205 & ~v_3122;
assign v_3127 = v_589 & v_3123;
assign v_3128 = ~v_3126 & ~v_3127;
assign v_3129 = v_208 & v_3124;
assign v_3130 = ~v_3129 & v_3128;
assign v_3131 = v_211 & v_3122;
assign v_3132 = ~v_3123 & v_3122;
assign v_3133 = v_212 & v_3132;
assign v_3134 = ~v_3131 & ~v_3133;
assign v_3135 = v_213 & v_3125;
assign v_3136 = ~v_3135 & v_3134;
assign v_3137 = v_217 & v_3122;
assign v_3138 = v_218 & v_3132;
assign v_3139 = ~v_3137 & ~v_3138;
assign v_3140 = v_219 & v_3125;
assign v_3141 = ~v_3140 & v_3139;
assign v_3142 = ~v_223 & ~v_3122;
assign v_3143 = v_606 & v_3123;
assign v_3144 = ~v_3142 & ~v_3143;
assign v_3145 = v_226 & v_3124;
assign v_3146 = ~v_3145 & v_3144;
assign v_3148 = ~v_3136 & v_172;
assign v_3149 = v_173 & v_3141;
assign v_3150 = ~v_3146 & v_174;
assign v_3151 = v_175 & v_3147;
assign v_3152 = ~v_3122 & v_176;
assign v_3153 = v_177 & v_3130;
assign v_3156 = ~v_235 & ~v_3122;
assign v_3157 = v_628 & v_3123;
assign v_3158 = ~v_3156 & ~v_3157;
assign v_3159 = v_238 & v_3124;
assign v_3160 = ~v_3159 & v_3158;
assign v_3161 = v_241 & v_3122;
assign v_3162 = v_242 & v_3132;
assign v_3163 = ~v_3161 & ~v_3162;
assign v_3164 = v_243 & v_3125;
assign v_3165 = ~v_3164 & v_3163;
assign v_3166 = v_247 & v_3122;
assign v_3167 = v_248 & v_3132;
assign v_3168 = ~v_3166 & ~v_3167;
assign v_3169 = v_249 & v_3125;
assign v_3170 = ~v_3169 & v_3168;
assign v_3171 = ~v_253 & ~v_3122;
assign v_3172 = v_644 & v_3123;
assign v_3173 = ~v_3171 & ~v_3172;
assign v_3174 = v_256 & v_3124;
assign v_3175 = ~v_3174 & v_3173;
assign v_3177 = ~v_3165 & v_107;
assign v_3178 = v_108 & v_3170;
assign v_3179 = ~v_3175 & v_109;
assign v_3180 = v_110 & v_3176;
assign v_3181 = ~v_3122 & v_111;
assign v_3182 = v_112 & v_3160;
assign v_3185 = v_3155 & v_3184;
assign v_3186 = ~v_3013 & v_3185;
assign v_3187 = v_2998 & v_3186;
assign v_3188 = v_675 & v_2993;
assign v_3189 = ~v_3188 & v_2993;
assign v_3190 = v_676 & v_2993;
assign v_3191 = v_677 & v_2993;
assign v_3192 = v_678 & v_2993;
assign v_3193 = ~v_205 & ~v_3189;
assign v_3194 = v_589 & v_3190;
assign v_3195 = ~v_3193 & ~v_3194;
assign v_3196 = v_208 & v_3191;
assign v_3197 = ~v_3196 & v_3195;
assign v_3198 = v_211 & v_3189;
assign v_3199 = ~v_3190 & v_3189;
assign v_3200 = v_212 & v_3199;
assign v_3201 = ~v_3198 & ~v_3200;
assign v_3202 = v_213 & v_3192;
assign v_3203 = ~v_3202 & v_3201;
assign v_3204 = v_217 & v_3189;
assign v_3205 = v_218 & v_3199;
assign v_3206 = ~v_3204 & ~v_3205;
assign v_3207 = v_219 & v_3192;
assign v_3208 = ~v_3207 & v_3206;
assign v_3209 = ~v_223 & ~v_3189;
assign v_3210 = v_606 & v_3190;
assign v_3211 = ~v_3209 & ~v_3210;
assign v_3212 = v_226 & v_3191;
assign v_3213 = ~v_3212 & v_3211;
assign v_3215 = ~v_3203 & v_172;
assign v_3216 = v_173 & v_3208;
assign v_3217 = ~v_3213 & v_174;
assign v_3218 = v_175 & v_3214;
assign v_3219 = ~v_3189 & v_176;
assign v_3220 = v_177 & v_3197;
assign v_3223 = ~v_235 & ~v_3189;
assign v_3224 = v_628 & v_3190;
assign v_3225 = ~v_3223 & ~v_3224;
assign v_3226 = v_238 & v_3191;
assign v_3227 = ~v_3226 & v_3225;
assign v_3228 = v_241 & v_3189;
assign v_3229 = v_242 & v_3199;
assign v_3230 = ~v_3228 & ~v_3229;
assign v_3231 = v_243 & v_3192;
assign v_3232 = ~v_3231 & v_3230;
assign v_3233 = v_247 & v_3189;
assign v_3234 = v_248 & v_3199;
assign v_3235 = ~v_3233 & ~v_3234;
assign v_3236 = v_249 & v_3192;
assign v_3237 = ~v_3236 & v_3235;
assign v_3238 = ~v_253 & ~v_3189;
assign v_3239 = v_644 & v_3190;
assign v_3240 = ~v_3238 & ~v_3239;
assign v_3241 = v_256 & v_3191;
assign v_3242 = ~v_3241 & v_3240;
assign v_3244 = ~v_3232 & v_107;
assign v_3245 = v_108 & v_3237;
assign v_3246 = ~v_3242 & v_109;
assign v_3247 = v_110 & v_3243;
assign v_3248 = ~v_3189 & v_111;
assign v_3249 = v_112 & v_3227;
assign v_3252 = v_3222 & v_3251;
assign v_3253 = v_2993 & v_3252;
assign v_3254 = v_2993 & v_3253;
assign v_3255 = ~v_3187 & ~v_3254;
assign v_3257 = v_3187 & v_3254;
assign v_3258 = ~v_3120 & v_3255;
assign v_3261 = v_3120 & v_3257;
assign v_3262 = ~v_3258 & v_2988;
assign v_3263 = ~v_3262 & v_2988;
assign v_522 = v_3264 | v_3265;
assign v_619 = v_3266 | v_3267;
assign v_656 = v_3268 | v_3269;
assign v_695 = v_3270 | v_3271;
assign v_701 = v_3272 | v_3273;
assign v_738 = v_3274 | v_3275;
assign v_767 = v_3276 | v_3277;
assign v_806 = v_3278 | v_3279;
assign v_835 = v_3280 | v_3281;
assign v_874 = v_3282 | v_3283;
assign v_903 = v_3284 | v_3285;
assign v_1038 = v_3286 | v_3287;
assign v_1121 = v_3288 | v_3289;
assign v_1124 = v_3290 | v_3291;
assign v_1161 = v_3292 | v_3293;
assign v_1190 = v_3294 | v_3295;
assign v_1229 = v_3296 | v_3297;
assign v_1258 = v_3298 | v_3299;
assign v_1297 = v_3300 | v_3301;
assign v_1326 = v_3302 | v_3303;
assign v_1365 = v_3304 | v_3305;
assign v_1394 = v_3306 | v_3307;
assign v_1856 = v_3308 | v_3309;
assign v_1885 = v_3310 | v_3311;
assign v_1924 = v_3312 | v_3313;
assign v_1953 = v_3314 | v_3315;
assign v_1992 = v_3316 | v_3317;
assign v_2021 = v_3318 | v_3319;
assign v_2060 = v_3320 | v_3321;
assign v_2089 = v_3322 | v_3323;
assign v_2302 = v_2285 | v_2290 | v_2294 | v_2298;
assign v_2303 = v_2286 | v_2291 | v_2295 | v_2299;
assign v_2304 = v_2287 | v_2292 | v_2296 | v_2300;
assign v_2305 = v_2288 | v_2293 | v_2297 | v_2301;
assign v_2461 = v_3324 | v_3325;
assign v_2501 = v_3326 | v_3327;
assign v_2542 = v_3328 | v_3329;
assign v_2573 = v_3330 | v_3331;
assign v_2616 = v_3332 | v_3333;
assign v_2647 = v_3334 | v_3335;
assign v_2690 = v_3336 | v_3337;
assign v_2721 = v_3338 | v_3339;
assign v_2764 = v_3340 | v_3341;
assign v_2795 = v_3342 | v_3343;
assign v_2987 = v_41 | v_43 | v_2984 | v_2985 | v_2986;
assign v_3043 = v_3344 | v_3345;
assign v_3046 = v_3346 | v_3347;
assign v_3049 = v_3348 | v_3349;
assign v_3051 = v_3350 | v_3351;
assign v_3087 = v_3352 | v_3353;
assign v_3116 = v_3354 | v_3355;
assign v_3154 = v_3356 | v_3357;
assign v_3183 = v_3358 | v_3359;
assign v_3221 = v_3360 | v_3361;
assign v_3250 = v_3362 | v_3363;
assign v_3264 = v_41 | v_517 | v_518 | v_519 | v_520;
assign v_3265 = v_521;
assign v_3266 = v_171 | v_613 | v_614 | v_615 | v_616;
assign v_3267 = v_617 | v_618;
assign v_3268 = v_106 | v_650 | v_651 | v_652 | v_653;
assign v_3269 = v_654 | v_655;
assign v_3270 = v_171 | v_173 | v_691 | v_692 | v_693;
assign v_3271 = v_694;
assign v_3272 = v_106 | v_108 | v_697 | v_698 | v_699;
assign v_3273 = v_700;
assign v_3274 = v_171 | v_732 | v_733 | v_734 | v_735;
assign v_3275 = v_736 | v_737;
assign v_3276 = v_106 | v_761 | v_762 | v_763 | v_764;
assign v_3277 = v_765 | v_766;
assign v_3278 = v_171 | v_800 | v_801 | v_802 | v_803;
assign v_3279 = v_804 | v_805;
assign v_3280 = v_106 | v_829 | v_830 | v_831 | v_832;
assign v_3281 = v_833 | v_834;
assign v_3282 = v_171 | v_868 | v_869 | v_870 | v_871;
assign v_3283 = v_872 | v_873;
assign v_3284 = v_106 | v_897 | v_898 | v_899 | v_900;
assign v_3285 = v_901 | v_902;
assign v_3286 = v_41 | v_1033 | v_1034 | v_1035 | v_1036;
assign v_3287 = v_1037;
assign v_3288 = v_171 | v_613 | v_614 | v_615 | v_616;
assign v_3289 = v_618 | v_1120;
assign v_3290 = v_106 | v_650 | v_651 | v_652 | v_653;
assign v_3291 = v_655 | v_1123;
assign v_3292 = v_171 | v_1155 | v_1156 | v_1157 | v_1158;
assign v_3293 = v_1159 | v_1160;
assign v_3294 = v_106 | v_1184 | v_1185 | v_1186 | v_1187;
assign v_3295 = v_1188 | v_1189;
assign v_3296 = v_171 | v_1223 | v_1224 | v_1225 | v_1226;
assign v_3297 = v_1227 | v_1228;
assign v_3298 = v_106 | v_1252 | v_1253 | v_1254 | v_1255;
assign v_3299 = v_1256 | v_1257;
assign v_3300 = v_171 | v_1291 | v_1292 | v_1293 | v_1294;
assign v_3301 = v_1295 | v_1296;
assign v_3302 = v_106 | v_1320 | v_1321 | v_1322 | v_1323;
assign v_3303 = v_1324 | v_1325;
assign v_3304 = v_171 | v_1359 | v_1360 | v_1361 | v_1362;
assign v_3305 = v_1363 | v_1364;
assign v_3306 = v_106 | v_1388 | v_1389 | v_1390 | v_1391;
assign v_3307 = v_1392 | v_1393;
assign v_3308 = v_171 | v_1850 | v_1851 | v_1852 | v_1853;
assign v_3309 = v_1854 | v_1855;
assign v_3310 = v_106 | v_1879 | v_1880 | v_1881 | v_1882;
assign v_3311 = v_1883 | v_1884;
assign v_3312 = v_171 | v_1918 | v_1919 | v_1920 | v_1921;
assign v_3313 = v_1922 | v_1923;
assign v_3314 = v_106 | v_1947 | v_1948 | v_1949 | v_1950;
assign v_3315 = v_1951 | v_1952;
assign v_3316 = v_171 | v_1986 | v_1987 | v_1988 | v_1989;
assign v_3317 = v_1990 | v_1991;
assign v_3318 = v_106 | v_2015 | v_2016 | v_2017 | v_2018;
assign v_3319 = v_2019 | v_2020;
assign v_3320 = v_171 | v_2054 | v_2055 | v_2056 | v_2057;
assign v_3321 = v_2058 | v_2059;
assign v_3322 = v_106 | v_2083 | v_2084 | v_2085 | v_2086;
assign v_3323 = v_2087 | v_2088;
assign v_3324 = v_367 | v_374 | v_2454 | v_2455 | v_2456;
assign v_3325 = v_2457 | v_2458 | v_2459 | v_2460;
assign v_3326 = v_302 | v_309 | v_2494 | v_2495 | v_2496;
assign v_3327 = v_2497 | v_2498 | v_2499 | v_2500;
assign v_3328 = v_367 | v_2534 | v_2535 | v_2536 | v_2537;
assign v_3329 = v_2538 | v_2539 | v_2540 | v_2541;
assign v_3330 = v_302 | v_2565 | v_2566 | v_2567 | v_2568;
assign v_3331 = v_2569 | v_2570 | v_2571 | v_2572;
assign v_3332 = v_367 | v_2608 | v_2609 | v_2610 | v_2611;
assign v_3333 = v_2612 | v_2613 | v_2614 | v_2615;
assign v_3334 = v_302 | v_2639 | v_2640 | v_2641 | v_2642;
assign v_3335 = v_2643 | v_2644 | v_2645 | v_2646;
assign v_3336 = v_367 | v_2682 | v_2683 | v_2684 | v_2685;
assign v_3337 = v_2686 | v_2687 | v_2688 | v_2689;
assign v_3338 = v_302 | v_2713 | v_2714 | v_2715 | v_2716;
assign v_3339 = v_2717 | v_2718 | v_2719 | v_2720;
assign v_3340 = v_367 | v_2756 | v_2757 | v_2758 | v_2759;
assign v_3341 = v_2760 | v_2761 | v_2762 | v_2763;
assign v_3342 = v_302 | v_2787 | v_2788 | v_2789 | v_2790;
assign v_3343 = v_2791 | v_2792 | v_2793 | v_2794;
assign v_3344 = v_171 | v_613 | v_614 | v_615 | v_616;
assign v_3345 = v_618 | v_3042;
assign v_3346 = v_106 | v_650 | v_651 | v_652 | v_653;
assign v_3347 = v_655 | v_3045;
assign v_3348 = v_171 | v_173 | v_176 | v_691 | v_692;
assign v_3349 = v_694;
assign v_3350 = v_106 | v_108 | v_111 | v_697 | v_698;
assign v_3351 = v_700;
assign v_3352 = v_171 | v_3081 | v_3082 | v_3083 | v_3084;
assign v_3353 = v_3085 | v_3086;
assign v_3354 = v_106 | v_3110 | v_3111 | v_3112 | v_3113;
assign v_3355 = v_3114 | v_3115;
assign v_3356 = v_171 | v_3148 | v_3149 | v_3150 | v_3151;
assign v_3357 = v_3152 | v_3153;
assign v_3358 = v_106 | v_3177 | v_3178 | v_3179 | v_3180;
assign v_3359 = v_3181 | v_3182;
assign v_3360 = v_171 | v_3215 | v_3216 | v_3217 | v_3218;
assign v_3361 = v_3219 | v_3220;
assign v_3362 = v_106 | v_3244 | v_3245 | v_3246 | v_3247;
assign v_3363 = v_3248 | v_3249;
assign v_909 = v_907 ^ v_839;
assign v_1400 = v_1398 ^ v_1330;
assign v_2095 = v_2093 ^ v_2025;
assign v_2801 = v_2799 ^ v_2725;
assign v_3256 = v_3254 ^ v_3187;
assign x_1 = v_516 | ~v_487 | ~v_495;
assign x_2 = v_495 | ~v_487 | ~v_516;
assign x_3 = v_487 | ~v_495 | ~v_516;
assign x_4 = v_516 | ~v_488 | ~v_496;
assign x_5 = v_496 | ~v_488 | ~v_516;
assign x_6 = v_488 | ~v_496 | ~v_516;
assign x_7 = v_516 | ~v_489 | ~v_497;
assign x_8 = v_497 | ~v_489 | ~v_516;
assign x_9 = v_489 | ~v_497 | ~v_516;
assign x_10 = v_516 | ~v_490 | ~v_498;
assign x_11 = v_498 | ~v_490 | ~v_516;
assign x_12 = v_490 | ~v_498 | ~v_516;
assign x_13 = v_487 | v_488 | v_489 | v_490 | ~v_516;
assign x_14 = v_495 | v_496 | v_497 | v_498 | ~v_516;
assign x_15 = v_509 | v_522 | ~v_523;
assign x_16 = v_504 | ~v_509 | ~v_523;
assign x_17 = v_504 | v_522 | ~v_523;
assign x_18 = v_523 | ~v_504 | ~v_522;
assign x_19 = v_523 | ~v_504 | ~v_509;
assign x_20 = v_509 | v_523 | ~v_522;
assign x_21 = v_487 | ~v_5 | ~v_525;
assign x_22 = v_5 | v_495 | ~v_525;
assign x_23 = v_487 | v_495 | ~v_525;
assign x_24 = v_525 | ~v_487 | ~v_495;
assign x_25 = v_5 | v_525 | ~v_495;
assign x_26 = v_525 | ~v_5 | ~v_487;
assign x_27 = v_488 | ~v_5 | ~v_526;
assign x_28 = v_5 | v_496 | ~v_526;
assign x_29 = v_488 | v_496 | ~v_526;
assign x_30 = v_526 | ~v_488 | ~v_496;
assign x_31 = v_5 | v_526 | ~v_496;
assign x_32 = v_526 | ~v_5 | ~v_488;
assign x_33 = v_489 | ~v_5 | ~v_527;
assign x_34 = v_5 | v_497 | ~v_527;
assign x_35 = v_489 | v_497 | ~v_527;
assign x_36 = v_527 | ~v_489 | ~v_497;
assign x_37 = v_5 | v_527 | ~v_497;
assign x_38 = v_527 | ~v_5 | ~v_489;
assign x_39 = v_490 | ~v_5 | ~v_528;
assign x_40 = v_5 | v_498 | ~v_528;
assign x_41 = v_490 | v_498 | ~v_528;
assign x_42 = v_528 | ~v_490 | ~v_498;
assign x_43 = v_5 | v_528 | ~v_498;
assign x_44 = v_528 | ~v_5 | ~v_490;
assign x_45 = v_491 | ~v_4 | ~v_529;
assign x_46 = v_4 | v_525 | ~v_529;
assign x_47 = v_491 | v_525 | ~v_529;
assign x_48 = v_529 | ~v_491 | ~v_525;
assign x_49 = v_4 | v_529 | ~v_525;
assign x_50 = v_529 | ~v_4 | ~v_491;
assign x_51 = v_492 | ~v_4 | ~v_530;
assign x_52 = v_4 | v_526 | ~v_530;
assign x_53 = v_492 | v_526 | ~v_530;
assign x_54 = v_530 | ~v_492 | ~v_526;
assign x_55 = v_4 | v_530 | ~v_526;
assign x_56 = v_530 | ~v_4 | ~v_492;
assign x_57 = v_493 | ~v_4 | ~v_531;
assign x_58 = v_4 | v_527 | ~v_531;
assign x_59 = v_493 | v_527 | ~v_531;
assign x_60 = v_531 | ~v_493 | ~v_527;
assign x_61 = v_4 | v_531 | ~v_527;
assign x_62 = v_531 | ~v_4 | ~v_493;
assign x_63 = v_494 | ~v_4 | ~v_532;
assign x_64 = v_4 | v_528 | ~v_532;
assign x_65 = v_494 | v_528 | ~v_532;
assign x_66 = v_532 | ~v_494 | ~v_528;
assign x_67 = v_4 | v_532 | ~v_528;
assign x_68 = v_532 | ~v_4 | ~v_494;
assign x_69 = ~v_529 | ~v_530;
assign x_70 = ~v_529 | ~v_531;
assign x_71 = ~v_529 | ~v_532;
assign x_72 = ~v_530 | ~v_531;
assign x_73 = ~v_530 | ~v_532;
assign x_74 = ~v_531 | ~v_532;
assign x_75 = v_532 | ~v_548 | ~v_549;
assign x_76 = ~v_532 | ~v_547 | ~v_549;
assign x_77 = ~v_547 | ~v_548 | ~v_549;
assign x_78 = v_547 | v_548 | v_549;
assign x_79 = v_547 | v_549 | ~v_532;
assign x_80 = v_532 | v_548 | v_549;
assign x_81 = v_532 | ~v_563 | ~v_564;
assign x_82 = ~v_532 | ~v_562 | ~v_564;
assign x_83 = ~v_562 | ~v_563 | ~v_564;
assign x_84 = v_562 | v_563 | v_564;
assign x_85 = v_562 | v_564 | ~v_532;
assign x_86 = v_532 | v_563 | v_564;
assign x_87 = v_534 | ~v_565 | ~v_566;
assign x_88 = v_564 | ~v_534 | ~v_566;
assign x_89 = v_564 | ~v_565 | ~v_566;
assign x_90 = v_565 | v_566 | ~v_564;
assign x_91 = v_566 | ~v_534 | ~v_564;
assign x_92 = v_534 | v_565 | v_566;
assign x_93 = v_611 | ~v_229 | ~v_584;
assign x_94 = v_584 | ~v_229 | ~v_611;
assign x_95 = v_229 | ~v_584 | ~v_611;
assign x_96 = v_611 | ~v_230 | ~v_585;
assign x_97 = v_585 | ~v_230 | ~v_611;
assign x_98 = v_230 | ~v_585 | ~v_611;
assign x_99 = v_611 | ~v_231 | ~v_586;
assign x_100 = v_586 | ~v_231 | ~v_611;
assign x_101 = v_231 | ~v_586 | ~v_611;
assign x_102 = v_611 | ~v_232 | ~v_587;
assign x_103 = v_587 | ~v_232 | ~v_611;
assign x_104 = v_232 | ~v_587 | ~v_611;
assign x_105 = v_229 | v_230 | v_231 | v_232 | ~v_611;
assign x_106 = v_584 | v_585 | v_586 | v_587 | ~v_611;
assign x_107 = v_612 | ~v_495 | ~v_584;
assign x_108 = v_584 | ~v_495 | ~v_612;
assign x_109 = v_495 | ~v_584 | ~v_612;
assign x_110 = v_612 | ~v_496 | ~v_585;
assign x_111 = v_585 | ~v_496 | ~v_612;
assign x_112 = v_496 | ~v_585 | ~v_612;
assign x_113 = v_612 | ~v_497 | ~v_586;
assign x_114 = v_586 | ~v_497 | ~v_612;
assign x_115 = v_497 | ~v_586 | ~v_612;
assign x_116 = v_612 | ~v_498 | ~v_587;
assign x_117 = v_587 | ~v_498 | ~v_612;
assign x_118 = v_498 | ~v_587 | ~v_612;
assign x_119 = v_495 | v_496 | v_497 | v_498 | ~v_612;
assign x_120 = v_584 | v_585 | v_586 | v_587 | ~v_612;
assign x_121 = v_583 | v_619 | ~v_620;
assign x_122 = v_593 | ~v_583 | ~v_620;
assign x_123 = v_593 | v_619 | ~v_620;
assign x_124 = v_620 | ~v_593 | ~v_619;
assign x_125 = v_620 | ~v_583 | ~v_593;
assign x_126 = v_583 | v_620 | ~v_619;
assign x_127 = v_649 | ~v_259 | ~v_584;
assign x_128 = v_584 | ~v_259 | ~v_649;
assign x_129 = v_259 | ~v_584 | ~v_649;
assign x_130 = v_649 | ~v_260 | ~v_585;
assign x_131 = v_585 | ~v_260 | ~v_649;
assign x_132 = v_260 | ~v_585 | ~v_649;
assign x_133 = v_649 | ~v_261 | ~v_586;
assign x_134 = v_586 | ~v_261 | ~v_649;
assign x_135 = v_261 | ~v_586 | ~v_649;
assign x_136 = v_649 | ~v_262 | ~v_587;
assign x_137 = v_587 | ~v_262 | ~v_649;
assign x_138 = v_262 | ~v_587 | ~v_649;
assign x_139 = v_259 | v_260 | v_261 | v_262 | ~v_649;
assign x_140 = v_584 | v_585 | v_586 | v_587 | ~v_649;
assign x_141 = v_626 | v_656 | ~v_657;
assign x_142 = v_632 | ~v_626 | ~v_657;
assign x_143 = v_632 | v_656 | ~v_657;
assign x_144 = v_657 | ~v_632 | ~v_656;
assign x_145 = v_657 | ~v_626 | ~v_632;
assign x_146 = v_626 | v_657 | ~v_656;
assign x_147 = v_583 | v_695 | ~v_696;
assign x_148 = v_205 | ~v_583 | ~v_696;
assign x_149 = v_205 | v_695 | ~v_696;
assign x_150 = v_696 | ~v_205 | ~v_695;
assign x_151 = v_696 | ~v_205 | ~v_583;
assign x_152 = v_583 | v_696 | ~v_695;
assign x_153 = v_626 | v_701 | ~v_702;
assign x_154 = v_235 | ~v_626 | ~v_702;
assign x_155 = v_235 | v_701 | ~v_702;
assign x_156 = v_702 | ~v_235 | ~v_701;
assign x_157 = v_702 | ~v_235 | ~v_626;
assign x_158 = v_626 | v_702 | ~v_701;
assign x_159 = v_705 | v_730 | ~v_229;
assign x_160 = v_229 | v_705 | ~v_730;
assign x_161 = ~v_229 | ~v_705 | ~v_730;
assign x_162 = v_730 | ~v_230 | ~v_706;
assign x_163 = v_706 | ~v_230 | ~v_730;
assign x_164 = v_230 | ~v_706 | ~v_730;
assign x_165 = v_730 | ~v_231 | ~v_707;
assign x_166 = v_707 | ~v_231 | ~v_730;
assign x_167 = v_231 | ~v_707 | ~v_730;
assign x_168 = v_730 | ~v_232 | ~v_708;
assign x_169 = v_708 | ~v_232 | ~v_730;
assign x_170 = v_232 | ~v_708 | ~v_730;
assign x_171 = v_230 | v_231 | v_232 | ~v_705 | ~v_730;
assign x_172 = v_229 | v_706 | v_707 | v_708 | ~v_730;
assign x_173 = v_705 | v_731 | ~v_495;
assign x_174 = v_495 | v_705 | ~v_731;
assign x_175 = ~v_495 | ~v_705 | ~v_731;
assign x_176 = v_731 | ~v_496 | ~v_706;
assign x_177 = v_706 | ~v_496 | ~v_731;
assign x_178 = v_496 | ~v_706 | ~v_731;
assign x_179 = v_731 | ~v_497 | ~v_707;
assign x_180 = v_707 | ~v_497 | ~v_731;
assign x_181 = v_497 | ~v_707 | ~v_731;
assign x_182 = v_731 | ~v_498 | ~v_708;
assign x_183 = v_708 | ~v_498 | ~v_731;
assign x_184 = v_498 | ~v_708 | ~v_731;
assign x_185 = v_496 | v_497 | v_498 | ~v_705 | ~v_731;
assign x_186 = v_495 | v_706 | v_707 | v_708 | ~v_731;
assign x_187 = v_583 | v_738 | ~v_739;
assign x_188 = v_713 | ~v_583 | ~v_739;
assign x_189 = v_713 | v_738 | ~v_739;
assign x_190 = v_739 | ~v_713 | ~v_738;
assign x_191 = v_739 | ~v_583 | ~v_713;
assign x_192 = v_583 | v_739 | ~v_738;
assign x_193 = v_705 | v_760 | ~v_259;
assign x_194 = v_259 | v_705 | ~v_760;
assign x_195 = ~v_259 | ~v_705 | ~v_760;
assign x_196 = v_760 | ~v_260 | ~v_706;
assign x_197 = v_706 | ~v_260 | ~v_760;
assign x_198 = v_260 | ~v_706 | ~v_760;
assign x_199 = v_760 | ~v_261 | ~v_707;
assign x_200 = v_707 | ~v_261 | ~v_760;
assign x_201 = v_261 | ~v_707 | ~v_760;
assign x_202 = v_760 | ~v_262 | ~v_708;
assign x_203 = v_708 | ~v_262 | ~v_760;
assign x_204 = v_262 | ~v_708 | ~v_760;
assign x_205 = v_260 | v_261 | v_262 | ~v_705 | ~v_760;
assign x_206 = v_259 | v_706 | v_707 | v_708 | ~v_760;
assign x_207 = v_626 | v_767 | ~v_768;
assign x_208 = v_744 | ~v_626 | ~v_768;
assign x_209 = v_744 | v_767 | ~v_768;
assign x_210 = v_768 | ~v_744 | ~v_767;
assign x_211 = v_768 | ~v_626 | ~v_744;
assign x_212 = v_626 | v_768 | ~v_767;
assign x_213 = v_773 | v_798 | ~v_229;
assign x_214 = v_229 | v_773 | ~v_798;
assign x_215 = ~v_229 | ~v_773 | ~v_798;
assign x_216 = v_798 | ~v_230 | ~v_774;
assign x_217 = v_774 | ~v_230 | ~v_798;
assign x_218 = v_230 | ~v_774 | ~v_798;
assign x_219 = v_798 | ~v_231 | ~v_775;
assign x_220 = v_775 | ~v_231 | ~v_798;
assign x_221 = v_231 | ~v_775 | ~v_798;
assign x_222 = v_798 | ~v_232 | ~v_776;
assign x_223 = v_776 | ~v_232 | ~v_798;
assign x_224 = v_232 | ~v_776 | ~v_798;
assign x_225 = v_230 | v_231 | v_232 | ~v_773 | ~v_798;
assign x_226 = v_229 | v_774 | v_775 | v_776 | ~v_798;
assign x_227 = v_773 | v_799 | ~v_495;
assign x_228 = v_495 | v_773 | ~v_799;
assign x_229 = ~v_495 | ~v_773 | ~v_799;
assign x_230 = v_799 | ~v_496 | ~v_774;
assign x_231 = v_774 | ~v_496 | ~v_799;
assign x_232 = v_496 | ~v_774 | ~v_799;
assign x_233 = v_799 | ~v_497 | ~v_775;
assign x_234 = v_775 | ~v_497 | ~v_799;
assign x_235 = v_497 | ~v_775 | ~v_799;
assign x_236 = v_799 | ~v_498 | ~v_776;
assign x_237 = v_776 | ~v_498 | ~v_799;
assign x_238 = v_498 | ~v_776 | ~v_799;
assign x_239 = v_496 | v_497 | v_498 | ~v_773 | ~v_799;
assign x_240 = v_495 | v_774 | v_775 | v_776 | ~v_799;
assign x_241 = v_583 | v_806 | ~v_807;
assign x_242 = v_781 | ~v_583 | ~v_807;
assign x_243 = v_781 | v_806 | ~v_807;
assign x_244 = v_807 | ~v_781 | ~v_806;
assign x_245 = v_807 | ~v_583 | ~v_781;
assign x_246 = v_583 | v_807 | ~v_806;
assign x_247 = v_773 | v_828 | ~v_259;
assign x_248 = v_259 | v_773 | ~v_828;
assign x_249 = ~v_259 | ~v_773 | ~v_828;
assign x_250 = v_828 | ~v_260 | ~v_774;
assign x_251 = v_774 | ~v_260 | ~v_828;
assign x_252 = v_260 | ~v_774 | ~v_828;
assign x_253 = v_828 | ~v_261 | ~v_775;
assign x_254 = v_775 | ~v_261 | ~v_828;
assign x_255 = v_261 | ~v_775 | ~v_828;
assign x_256 = v_828 | ~v_262 | ~v_776;
assign x_257 = v_776 | ~v_262 | ~v_828;
assign x_258 = v_262 | ~v_776 | ~v_828;
assign x_259 = v_260 | v_261 | v_262 | ~v_773 | ~v_828;
assign x_260 = v_259 | v_774 | v_775 | v_776 | ~v_828;
assign x_261 = v_626 | v_835 | ~v_836;
assign x_262 = v_812 | ~v_626 | ~v_836;
assign x_263 = v_812 | v_835 | ~v_836;
assign x_264 = v_836 | ~v_812 | ~v_835;
assign x_265 = v_836 | ~v_626 | ~v_812;
assign x_266 = v_626 | v_836 | ~v_835;
assign x_267 = v_841 | v_866 | ~v_229;
assign x_268 = v_229 | v_841 | ~v_866;
assign x_269 = ~v_229 | ~v_841 | ~v_866;
assign x_270 = v_866 | ~v_230 | ~v_842;
assign x_271 = v_842 | ~v_230 | ~v_866;
assign x_272 = v_230 | ~v_842 | ~v_866;
assign x_273 = v_866 | ~v_231 | ~v_843;
assign x_274 = v_843 | ~v_231 | ~v_866;
assign x_275 = v_231 | ~v_843 | ~v_866;
assign x_276 = v_866 | ~v_232 | ~v_844;
assign x_277 = v_844 | ~v_232 | ~v_866;
assign x_278 = v_232 | ~v_844 | ~v_866;
assign x_279 = v_230 | v_231 | v_232 | ~v_841 | ~v_866;
assign x_280 = v_229 | v_842 | v_843 | v_844 | ~v_866;
assign x_281 = v_841 | v_867 | ~v_495;
assign x_282 = v_495 | v_841 | ~v_867;
assign x_283 = ~v_495 | ~v_841 | ~v_867;
assign x_284 = v_867 | ~v_496 | ~v_842;
assign x_285 = v_842 | ~v_496 | ~v_867;
assign x_286 = v_496 | ~v_842 | ~v_867;
assign x_287 = v_867 | ~v_497 | ~v_843;
assign x_288 = v_843 | ~v_497 | ~v_867;
assign x_289 = v_497 | ~v_843 | ~v_867;
assign x_290 = v_867 | ~v_498 | ~v_844;
assign x_291 = v_844 | ~v_498 | ~v_867;
assign x_292 = v_498 | ~v_844 | ~v_867;
assign x_293 = v_496 | v_497 | v_498 | ~v_841 | ~v_867;
assign x_294 = v_495 | v_842 | v_843 | v_844 | ~v_867;
assign x_295 = v_583 | v_874 | ~v_875;
assign x_296 = v_849 | ~v_583 | ~v_875;
assign x_297 = v_849 | v_874 | ~v_875;
assign x_298 = v_875 | ~v_849 | ~v_874;
assign x_299 = v_875 | ~v_583 | ~v_849;
assign x_300 = v_583 | v_875 | ~v_874;
assign x_301 = v_841 | v_896 | ~v_259;
assign x_302 = v_259 | v_841 | ~v_896;
assign x_303 = ~v_259 | ~v_841 | ~v_896;
assign x_304 = v_896 | ~v_260 | ~v_842;
assign x_305 = v_842 | ~v_260 | ~v_896;
assign x_306 = v_260 | ~v_842 | ~v_896;
assign x_307 = v_896 | ~v_261 | ~v_843;
assign x_308 = v_843 | ~v_261 | ~v_896;
assign x_309 = v_261 | ~v_843 | ~v_896;
assign x_310 = v_896 | ~v_262 | ~v_844;
assign x_311 = v_844 | ~v_262 | ~v_896;
assign x_312 = v_262 | ~v_844 | ~v_896;
assign x_313 = v_260 | v_261 | v_262 | ~v_841 | ~v_896;
assign x_314 = v_259 | v_842 | v_843 | v_844 | ~v_896;
assign x_315 = v_626 | v_903 | ~v_904;
assign x_316 = v_880 | ~v_626 | ~v_904;
assign x_317 = v_880 | v_903 | ~v_904;
assign x_318 = v_904 | ~v_880 | ~v_903;
assign x_319 = v_904 | ~v_626 | ~v_880;
assign x_320 = v_626 | v_904 | ~v_903;
assign x_321 = ~v_908 | ~v_909;
assign x_322 = ~v_908 | ~v_910;
assign x_323 = ~v_909 | ~v_910;
assign x_324 = v_908 | ~v_771 | ~v_912;
assign x_325 = v_771 | v_909 | ~v_912;
assign x_326 = v_908 | v_909 | ~v_912;
assign x_327 = v_912 | ~v_908 | ~v_909;
assign x_328 = v_771 | v_912 | ~v_909;
assign x_329 = v_912 | ~v_771 | ~v_908;
assign x_330 = v_909 | ~v_771 | ~v_913;
assign x_331 = v_771 | v_910 | ~v_913;
assign x_332 = v_909 | v_910 | ~v_913;
assign x_333 = v_913 | ~v_909 | ~v_910;
assign x_334 = v_771 | v_913 | ~v_910;
assign x_335 = v_913 | ~v_771 | ~v_909;
assign x_336 = ~v_911 | ~v_912;
assign x_337 = ~v_911 | ~v_913;
assign x_338 = ~v_911 | ~v_914;
assign x_339 = ~v_912 | ~v_913;
assign x_340 = ~v_912 | ~v_914;
assign x_341 = ~v_913 | ~v_914;
assign x_342 = v_915 | ~v_491 | ~v_911;
assign x_343 = v_911 | ~v_491 | ~v_915;
assign x_344 = v_491 | ~v_911 | ~v_915;
assign x_345 = v_915 | ~v_492 | ~v_912;
assign x_346 = v_912 | ~v_492 | ~v_915;
assign x_347 = v_492 | ~v_912 | ~v_915;
assign x_348 = v_915 | ~v_493 | ~v_913;
assign x_349 = v_913 | ~v_493 | ~v_915;
assign x_350 = v_493 | ~v_913 | ~v_915;
assign x_351 = v_915 | ~v_494 | ~v_914;
assign x_352 = v_914 | ~v_494 | ~v_915;
assign x_353 = v_494 | ~v_914 | ~v_915;
assign x_354 = v_491 | v_492 | v_493 | v_494 | ~v_915;
assign x_355 = v_911 | v_912 | v_913 | v_914 | ~v_915;
assign x_356 = v_549 | v_907 | ~v_919;
assign x_357 = ~v_907 | ~v_918 | ~v_919;
assign x_358 = v_549 | ~v_918 | ~v_919;
assign x_359 = v_918 | v_919 | ~v_549;
assign x_360 = v_918 | v_919 | ~v_907;
assign x_361 = v_907 | v_919 | ~v_549;
assign x_362 = v_919 | ~v_839 | ~v_922;
assign x_363 = v_839 | ~v_918 | ~v_922;
assign x_364 = v_919 | ~v_918 | ~v_922;
assign x_365 = v_918 | v_922 | ~v_919;
assign x_366 = v_839 | v_918 | v_922;
assign x_367 = v_922 | ~v_839 | ~v_919;
assign x_368 = v_920 | ~v_839 | ~v_923;
assign x_369 = v_839 | v_918 | ~v_923;
assign x_370 = v_918 | v_920 | ~v_923;
assign x_371 = v_923 | ~v_918 | ~v_920;
assign x_372 = v_839 | v_923 | ~v_918;
assign x_373 = v_923 | ~v_839 | ~v_920;
assign x_374 = v_566 | ~v_908 | ~v_925;
assign x_375 = v_908 | v_922 | ~v_925;
assign x_376 = v_566 | v_922 | ~v_925;
assign x_377 = v_925 | ~v_566 | ~v_922;
assign x_378 = v_908 | v_925 | ~v_922;
assign x_379 = v_925 | ~v_566 | ~v_908;
assign x_380 = v_925 | ~v_771 | ~v_929;
assign x_381 = v_771 | v_922 | ~v_929;
assign x_382 = v_922 | v_925 | ~v_929;
assign x_383 = v_929 | ~v_922 | ~v_925;
assign x_384 = v_771 | v_929 | ~v_922;
assign x_385 = v_929 | ~v_771 | ~v_925;
assign x_386 = v_926 | ~v_771 | ~v_930;
assign x_387 = v_771 | v_923 | ~v_930;
assign x_388 = v_923 | v_926 | ~v_930;
assign x_389 = v_930 | ~v_923 | ~v_926;
assign x_390 = v_771 | v_930 | ~v_923;
assign x_391 = v_930 | ~v_771 | ~v_926;
assign x_392 = v_927 | ~v_771 | ~v_931;
assign x_393 = v_771 | v_924 | ~v_931;
assign x_394 = v_924 | v_927 | ~v_931;
assign x_395 = v_931 | ~v_924 | ~v_927;
assign x_396 = v_771 | v_931 | ~v_924;
assign x_397 = v_931 | ~v_771 | ~v_927;
assign x_398 = v_953 | v_960 | ~v_659;
assign x_399 = v_659 | v_953 | ~v_960;
assign x_400 = ~v_659 | ~v_953 | ~v_960;
assign x_401 = v_955 | v_960 | ~v_660;
assign x_402 = v_660 | v_955 | ~v_960;
assign x_403 = ~v_660 | ~v_955 | ~v_960;
assign x_404 = v_957 | v_960 | ~v_661;
assign x_405 = v_661 | v_957 | ~v_960;
assign x_406 = ~v_661 | ~v_957 | ~v_960;
assign x_407 = v_959 | v_960 | ~v_662;
assign x_408 = v_662 | v_959 | ~v_960;
assign x_409 = ~v_662 | ~v_959 | ~v_960;
assign x_410 = ~v_953 | ~v_955 | ~v_957 | ~v_959 | ~v_960;
assign x_411 = v_659 | v_660 | v_661 | v_662 | ~v_960;
assign x_412 = v_491 | ~v_961 | ~v_962;
assign x_413 = ~v_491 | ~v_915 | ~v_962;
assign x_414 = ~v_915 | ~v_961 | ~v_962;
assign x_415 = v_915 | v_961 | v_962;
assign x_416 = v_915 | v_962 | ~v_491;
assign x_417 = v_491 | v_961 | v_962;
assign x_418 = v_566 | ~v_909 | ~v_968;
assign x_419 = v_909 | ~v_967 | ~v_968;
assign x_420 = v_566 | ~v_967 | ~v_968;
assign x_421 = v_967 | v_968 | ~v_566;
assign x_422 = v_909 | v_967 | v_968;
assign x_423 = v_968 | ~v_566 | ~v_909;
assign x_424 = v_968 | ~v_771 | ~v_971;
assign x_425 = v_771 | ~v_967 | ~v_971;
assign x_426 = v_968 | ~v_967 | ~v_971;
assign x_427 = v_967 | v_971 | ~v_968;
assign x_428 = v_771 | v_967 | v_971;
assign x_429 = v_971 | ~v_771 | ~v_968;
assign x_430 = v_969 | ~v_771 | ~v_972;
assign x_431 = v_771 | v_967 | ~v_972;
assign x_432 = v_967 | v_969 | ~v_972;
assign x_433 = v_972 | ~v_967 | ~v_969;
assign x_434 = v_771 | v_972 | ~v_967;
assign x_435 = v_972 | ~v_771 | ~v_969;
assign x_436 = v_985 | v_992 | ~v_663;
assign x_437 = v_663 | v_985 | ~v_992;
assign x_438 = ~v_663 | ~v_985 | ~v_992;
assign x_439 = v_987 | v_992 | ~v_664;
assign x_440 = v_664 | v_987 | ~v_992;
assign x_441 = ~v_664 | ~v_987 | ~v_992;
assign x_442 = v_989 | v_992 | ~v_665;
assign x_443 = v_665 | v_989 | ~v_992;
assign x_444 = ~v_665 | ~v_989 | ~v_992;
assign x_445 = v_991 | v_992 | ~v_666;
assign x_446 = v_666 | v_991 | ~v_992;
assign x_447 = ~v_666 | ~v_991 | ~v_992;
assign x_448 = ~v_985 | ~v_987 | ~v_989 | ~v_991 | ~v_992;
assign x_449 = v_663 | v_664 | v_665 | v_666 | ~v_992;
assign x_450 = ~v_963 | ~v_993 | ~v_994;
assign x_451 = v_962 | v_963 | ~v_994;
assign x_452 = v_962 | ~v_993 | ~v_994;
assign x_453 = v_993 | v_994 | ~v_962;
assign x_454 = v_963 | v_994 | ~v_962;
assign x_455 = v_993 | v_994 | ~v_963;
assign x_456 = v_1003 | v_1007 | ~v_667;
assign x_457 = v_667 | v_1003 | ~v_1007;
assign x_458 = ~v_667 | ~v_1003 | ~v_1007;
assign x_459 = v_1007 | ~v_668 | ~v_1004;
assign x_460 = v_1004 | ~v_668 | ~v_1007;
assign x_461 = v_668 | ~v_1004 | ~v_1007;
assign x_462 = v_1007 | ~v_669 | ~v_1005;
assign x_463 = v_1005 | ~v_669 | ~v_1007;
assign x_464 = v_669 | ~v_1005 | ~v_1007;
assign x_465 = v_1007 | ~v_670 | ~v_1006;
assign x_466 = v_1006 | ~v_670 | ~v_1007;
assign x_467 = v_670 | ~v_1006 | ~v_1007;
assign x_468 = v_668 | v_669 | v_670 | ~v_1003 | ~v_1007;
assign x_469 = v_667 | v_1004 | v_1005 | v_1006 | ~v_1007;
assign x_470 = ~v_494 | ~v_1008 | ~v_1009;
assign x_471 = v_494 | v_994 | ~v_1009;
assign x_472 = v_994 | ~v_1008 | ~v_1009;
assign x_473 = v_1008 | v_1009 | ~v_994;
assign x_474 = v_494 | v_1009 | ~v_994;
assign x_475 = v_1008 | v_1009 | ~v_494;
assign x_476 = ~v_495 | ~v_496;
assign x_477 = ~v_495 | ~v_497;
assign x_478 = ~v_495 | ~v_498;
assign x_479 = ~v_496 | ~v_497;
assign x_480 = ~v_496 | ~v_498;
assign x_481 = ~v_497 | ~v_498;
assign x_482 = v_1032 | ~v_488 | ~v_495;
assign x_483 = v_495 | ~v_488 | ~v_1032;
assign x_484 = v_488 | ~v_495 | ~v_1032;
assign x_485 = v_1032 | ~v_489 | ~v_496;
assign x_486 = v_496 | ~v_489 | ~v_1032;
assign x_487 = v_489 | ~v_496 | ~v_1032;
assign x_488 = v_1032 | ~v_490 | ~v_497;
assign x_489 = v_497 | ~v_490 | ~v_1032;
assign x_490 = v_490 | ~v_497 | ~v_1032;
assign x_491 = v_488 | v_489 | v_490 | ~v_1032;
assign x_492 = v_495 | v_496 | v_497 | ~v_1032;
assign x_493 = v_509 | v_1038 | ~v_1039;
assign x_494 = v_1025 | ~v_509 | ~v_1039;
assign x_495 = v_1025 | v_1038 | ~v_1039;
assign x_496 = v_1039 | ~v_1025 | ~v_1038;
assign x_497 = v_1039 | ~v_509 | ~v_1025;
assign x_498 = v_509 | v_1039 | ~v_1038;
assign x_499 = v_488 | ~v_5 | ~v_1042;
assign x_500 = v_5 | v_495 | ~v_1042;
assign x_501 = v_488 | v_495 | ~v_1042;
assign x_502 = v_1042 | ~v_488 | ~v_495;
assign x_503 = v_5 | v_1042 | ~v_495;
assign x_504 = v_1042 | ~v_5 | ~v_488;
assign x_505 = v_489 | ~v_5 | ~v_1043;
assign x_506 = v_5 | v_496 | ~v_1043;
assign x_507 = v_489 | v_496 | ~v_1043;
assign x_508 = v_1043 | ~v_489 | ~v_496;
assign x_509 = v_5 | v_1043 | ~v_496;
assign x_510 = v_1043 | ~v_5 | ~v_489;
assign x_511 = v_490 | ~v_5 | ~v_1044;
assign x_512 = v_5 | v_497 | ~v_1044;
assign x_513 = v_490 | v_497 | ~v_1044;
assign x_514 = v_1044 | ~v_490 | ~v_497;
assign x_515 = v_5 | v_1044 | ~v_497;
assign x_516 = v_1044 | ~v_5 | ~v_490;
assign x_517 = ~v_491 | ~v_492;
assign x_518 = ~v_491 | ~v_493;
assign x_519 = ~v_491 | ~v_494;
assign x_520 = ~v_492 | ~v_493;
assign x_521 = ~v_492 | ~v_494;
assign x_522 = ~v_493 | ~v_494;
assign x_523 = v_491 | ~v_4 | ~v_1047;
assign x_524 = v_4 | v_1042 | ~v_1047;
assign x_525 = v_491 | v_1042 | ~v_1047;
assign x_526 = v_1047 | ~v_491 | ~v_1042;
assign x_527 = v_4 | v_1047 | ~v_1042;
assign x_528 = v_1047 | ~v_4 | ~v_491;
assign x_529 = v_492 | ~v_4 | ~v_1048;
assign x_530 = v_4 | v_1043 | ~v_1048;
assign x_531 = v_492 | v_1043 | ~v_1048;
assign x_532 = v_1048 | ~v_492 | ~v_1043;
assign x_533 = v_4 | v_1048 | ~v_1043;
assign x_534 = v_1048 | ~v_4 | ~v_492;
assign x_535 = v_493 | ~v_4 | ~v_1049;
assign x_536 = v_4 | v_1044 | ~v_1049;
assign x_537 = v_493 | v_1044 | ~v_1049;
assign x_538 = v_1049 | ~v_493 | ~v_1044;
assign x_539 = v_4 | v_1049 | ~v_1044;
assign x_540 = v_1049 | ~v_4 | ~v_493;
assign x_541 = v_494 | ~v_4 | ~v_1050;
assign x_542 = v_4 | v_1045 | ~v_1050;
assign x_543 = v_494 | v_1045 | ~v_1050;
assign x_544 = v_1050 | ~v_494 | ~v_1045;
assign x_545 = v_4 | v_1050 | ~v_1045;
assign x_546 = v_1050 | ~v_4 | ~v_494;
assign x_547 = ~v_1046 | ~v_1047;
assign x_548 = ~v_1046 | ~v_1048;
assign x_549 = ~v_1046 | ~v_1049;
assign x_550 = ~v_1046 | ~v_1050;
assign x_551 = ~v_1047 | ~v_1048;
assign x_552 = ~v_1047 | ~v_1049;
assign x_553 = ~v_1047 | ~v_1050;
assign x_554 = ~v_1048 | ~v_1049;
assign x_555 = ~v_1048 | ~v_1050;
assign x_556 = ~v_1049 | ~v_1050;
assign x_557 = v_1050 | ~v_1066 | ~v_1067;
assign x_558 = ~v_1050 | ~v_1052 | ~v_1067;
assign x_559 = ~v_1052 | ~v_1066 | ~v_1067;
assign x_560 = v_1052 | v_1066 | v_1067;
assign x_561 = v_1052 | v_1067 | ~v_1050;
assign x_562 = v_1050 | v_1066 | v_1067;
assign x_563 = v_1053 | ~v_1068 | ~v_1069;
assign x_564 = v_1067 | ~v_1053 | ~v_1069;
assign x_565 = v_1067 | ~v_1068 | ~v_1069;
assign x_566 = v_1068 | v_1069 | ~v_1067;
assign x_567 = v_1069 | ~v_1053 | ~v_1067;
assign x_568 = v_1053 | v_1068 | v_1069;
assign x_569 = v_1050 | ~v_1082 | ~v_1083;
assign x_570 = ~v_1050 | ~v_1053 | ~v_1083;
assign x_571 = ~v_1053 | ~v_1082 | ~v_1083;
assign x_572 = v_1053 | v_1082 | v_1083;
assign x_573 = v_1053 | v_1083 | ~v_1050;
assign x_574 = v_1050 | v_1082 | v_1083;
assign x_575 = v_1053 | ~v_1084 | ~v_1085;
assign x_576 = v_1083 | ~v_1053 | ~v_1085;
assign x_577 = v_1083 | ~v_1084 | ~v_1085;
assign x_578 = v_1084 | v_1085 | ~v_1083;
assign x_579 = v_1085 | ~v_1053 | ~v_1083;
assign x_580 = v_1053 | v_1084 | v_1085;
assign x_581 = v_1052 | ~v_1086 | ~v_1087;
assign x_582 = v_1085 | ~v_1052 | ~v_1087;
assign x_583 = v_1085 | ~v_1086 | ~v_1087;
assign x_584 = v_1086 | v_1087 | ~v_1085;
assign x_585 = v_1087 | ~v_1052 | ~v_1085;
assign x_586 = v_1052 | v_1086 | v_1087;
assign x_587 = v_1050 | ~v_1100 | ~v_1101;
assign x_588 = ~v_1050 | ~v_1101;
assign x_589 = ~v_1050 | ~v_1100 | ~v_1101;
assign x_590 = v_1050 | v_1100 | v_1101;
assign x_591 = v_1050 | v_1100 | v_1101;
assign x_592 = v_1053 | ~v_1102 | ~v_1103;
assign x_593 = v_1101 | ~v_1053 | ~v_1103;
assign x_594 = v_1101 | ~v_1102 | ~v_1103;
assign x_595 = v_1102 | v_1103 | ~v_1101;
assign x_596 = v_1103 | ~v_1053 | ~v_1101;
assign x_597 = v_1053 | v_1102 | v_1103;
assign x_598 = v_1052 | ~v_1104 | ~v_1105;
assign x_599 = v_1103 | ~v_1052 | ~v_1105;
assign x_600 = v_1103 | ~v_1104 | ~v_1105;
assign x_601 = v_1104 | v_1105 | ~v_1103;
assign x_602 = v_1105 | ~v_1052 | ~v_1103;
assign x_603 = v_1052 | v_1104 | v_1105;
assign x_604 = ~v_1046 | ~v_1106 | ~v_1107;
assign x_605 = v_1046 | v_1105 | ~v_1107;
assign x_606 = v_1105 | ~v_1106 | ~v_1107;
assign x_607 = v_1106 | v_1107 | ~v_1105;
assign x_608 = v_1046 | v_1107 | ~v_1105;
assign x_609 = v_1106 | v_1107 | ~v_1046;
assign x_610 = v_1119 | ~v_495 | ~v_585;
assign x_611 = v_585 | ~v_495 | ~v_1119;
assign x_612 = v_495 | ~v_585 | ~v_1119;
assign x_613 = v_1119 | ~v_496 | ~v_586;
assign x_614 = v_586 | ~v_496 | ~v_1119;
assign x_615 = v_496 | ~v_586 | ~v_1119;
assign x_616 = v_1119 | ~v_497 | ~v_587;
assign x_617 = v_587 | ~v_497 | ~v_1119;
assign x_618 = v_497 | ~v_587 | ~v_1119;
assign x_619 = v_495 | v_496 | v_497 | ~v_1119;
assign x_620 = v_585 | v_586 | v_587 | ~v_1119;
assign x_621 = v_583 | v_1121 | ~v_1122;
assign x_622 = v_593 | ~v_583 | ~v_1122;
assign x_623 = v_593 | v_1121 | ~v_1122;
assign x_624 = v_1122 | ~v_593 | ~v_1121;
assign x_625 = v_1122 | ~v_583 | ~v_593;
assign x_626 = v_583 | v_1122 | ~v_1121;
assign x_627 = v_626 | v_1124 | ~v_1125;
assign x_628 = v_632 | ~v_626 | ~v_1125;
assign x_629 = v_632 | v_1124 | ~v_1125;
assign x_630 = v_1125 | ~v_632 | ~v_1124;
assign x_631 = v_1125 | ~v_626 | ~v_632;
assign x_632 = v_626 | v_1125 | ~v_1124;
assign x_633 = v_1128 | v_1153 | ~v_229;
assign x_634 = v_229 | v_1128 | ~v_1153;
assign x_635 = ~v_229 | ~v_1128 | ~v_1153;
assign x_636 = v_1153 | ~v_230 | ~v_1129;
assign x_637 = v_1129 | ~v_230 | ~v_1153;
assign x_638 = v_230 | ~v_1129 | ~v_1153;
assign x_639 = v_1153 | ~v_231 | ~v_1130;
assign x_640 = v_1130 | ~v_231 | ~v_1153;
assign x_641 = v_231 | ~v_1130 | ~v_1153;
assign x_642 = v_1153 | ~v_232 | ~v_1131;
assign x_643 = v_1131 | ~v_232 | ~v_1153;
assign x_644 = v_232 | ~v_1131 | ~v_1153;
assign x_645 = v_230 | v_231 | v_232 | ~v_1128 | ~v_1153;
assign x_646 = v_229 | v_1129 | v_1130 | v_1131 | ~v_1153;
assign x_647 = v_1154 | ~v_495 | ~v_1129;
assign x_648 = v_1129 | ~v_495 | ~v_1154;
assign x_649 = v_495 | ~v_1129 | ~v_1154;
assign x_650 = v_1154 | ~v_496 | ~v_1130;
assign x_651 = v_1130 | ~v_496 | ~v_1154;
assign x_652 = v_496 | ~v_1130 | ~v_1154;
assign x_653 = v_1154 | ~v_497 | ~v_1131;
assign x_654 = v_1131 | ~v_497 | ~v_1154;
assign x_655 = v_497 | ~v_1131 | ~v_1154;
assign x_656 = v_495 | v_496 | v_497 | ~v_1154;
assign x_657 = v_1129 | v_1130 | v_1131 | ~v_1154;
assign x_658 = v_583 | v_1161 | ~v_1162;
assign x_659 = v_1136 | ~v_583 | ~v_1162;
assign x_660 = v_1136 | v_1161 | ~v_1162;
assign x_661 = v_1162 | ~v_1136 | ~v_1161;
assign x_662 = v_1162 | ~v_583 | ~v_1136;
assign x_663 = v_583 | v_1162 | ~v_1161;
assign x_664 = v_1128 | v_1183 | ~v_259;
assign x_665 = v_259 | v_1128 | ~v_1183;
assign x_666 = ~v_259 | ~v_1128 | ~v_1183;
assign x_667 = v_1183 | ~v_260 | ~v_1129;
assign x_668 = v_1129 | ~v_260 | ~v_1183;
assign x_669 = v_260 | ~v_1129 | ~v_1183;
assign x_670 = v_1183 | ~v_261 | ~v_1130;
assign x_671 = v_1130 | ~v_261 | ~v_1183;
assign x_672 = v_261 | ~v_1130 | ~v_1183;
assign x_673 = v_1183 | ~v_262 | ~v_1131;
assign x_674 = v_1131 | ~v_262 | ~v_1183;
assign x_675 = v_262 | ~v_1131 | ~v_1183;
assign x_676 = v_260 | v_261 | v_262 | ~v_1128 | ~v_1183;
assign x_677 = v_259 | v_1129 | v_1130 | v_1131 | ~v_1183;
assign x_678 = v_626 | v_1190 | ~v_1191;
assign x_679 = v_1167 | ~v_626 | ~v_1191;
assign x_680 = v_1167 | v_1190 | ~v_1191;
assign x_681 = v_1191 | ~v_1167 | ~v_1190;
assign x_682 = v_1191 | ~v_626 | ~v_1167;
assign x_683 = v_626 | v_1191 | ~v_1190;
assign x_684 = v_1196 | v_1221 | ~v_229;
assign x_685 = v_229 | v_1196 | ~v_1221;
assign x_686 = ~v_229 | ~v_1196 | ~v_1221;
assign x_687 = v_1221 | ~v_230 | ~v_1197;
assign x_688 = v_1197 | ~v_230 | ~v_1221;
assign x_689 = v_230 | ~v_1197 | ~v_1221;
assign x_690 = v_1221 | ~v_231 | ~v_1198;
assign x_691 = v_1198 | ~v_231 | ~v_1221;
assign x_692 = v_231 | ~v_1198 | ~v_1221;
assign x_693 = v_1221 | ~v_232 | ~v_1199;
assign x_694 = v_1199 | ~v_232 | ~v_1221;
assign x_695 = v_232 | ~v_1199 | ~v_1221;
assign x_696 = v_230 | v_231 | v_232 | ~v_1196 | ~v_1221;
assign x_697 = v_229 | v_1197 | v_1198 | v_1199 | ~v_1221;
assign x_698 = v_1222 | ~v_495 | ~v_1197;
assign x_699 = v_1197 | ~v_495 | ~v_1222;
assign x_700 = v_495 | ~v_1197 | ~v_1222;
assign x_701 = v_1222 | ~v_496 | ~v_1198;
assign x_702 = v_1198 | ~v_496 | ~v_1222;
assign x_703 = v_496 | ~v_1198 | ~v_1222;
assign x_704 = v_1222 | ~v_497 | ~v_1199;
assign x_705 = v_1199 | ~v_497 | ~v_1222;
assign x_706 = v_497 | ~v_1199 | ~v_1222;
assign x_707 = v_495 | v_496 | v_497 | ~v_1222;
assign x_708 = v_1197 | v_1198 | v_1199 | ~v_1222;
assign x_709 = v_583 | v_1229 | ~v_1230;
assign x_710 = v_1204 | ~v_583 | ~v_1230;
assign x_711 = v_1204 | v_1229 | ~v_1230;
assign x_712 = v_1230 | ~v_1204 | ~v_1229;
assign x_713 = v_1230 | ~v_583 | ~v_1204;
assign x_714 = v_583 | v_1230 | ~v_1229;
assign x_715 = v_1196 | v_1251 | ~v_259;
assign x_716 = v_259 | v_1196 | ~v_1251;
assign x_717 = ~v_259 | ~v_1196 | ~v_1251;
assign x_718 = v_1251 | ~v_260 | ~v_1197;
assign x_719 = v_1197 | ~v_260 | ~v_1251;
assign x_720 = v_260 | ~v_1197 | ~v_1251;
assign x_721 = v_1251 | ~v_261 | ~v_1198;
assign x_722 = v_1198 | ~v_261 | ~v_1251;
assign x_723 = v_261 | ~v_1198 | ~v_1251;
assign x_724 = v_1251 | ~v_262 | ~v_1199;
assign x_725 = v_1199 | ~v_262 | ~v_1251;
assign x_726 = v_262 | ~v_1199 | ~v_1251;
assign x_727 = v_260 | v_261 | v_262 | ~v_1196 | ~v_1251;
assign x_728 = v_259 | v_1197 | v_1198 | v_1199 | ~v_1251;
assign x_729 = v_626 | v_1258 | ~v_1259;
assign x_730 = v_1235 | ~v_626 | ~v_1259;
assign x_731 = v_1235 | v_1258 | ~v_1259;
assign x_732 = v_1259 | ~v_1235 | ~v_1258;
assign x_733 = v_1259 | ~v_626 | ~v_1235;
assign x_734 = v_626 | v_1259 | ~v_1258;
assign x_735 = v_1264 | v_1289 | ~v_229;
assign x_736 = v_229 | v_1264 | ~v_1289;
assign x_737 = ~v_229 | ~v_1264 | ~v_1289;
assign x_738 = v_1289 | ~v_230 | ~v_1265;
assign x_739 = v_1265 | ~v_230 | ~v_1289;
assign x_740 = v_230 | ~v_1265 | ~v_1289;
assign x_741 = v_1289 | ~v_231 | ~v_1266;
assign x_742 = v_1266 | ~v_231 | ~v_1289;
assign x_743 = v_231 | ~v_1266 | ~v_1289;
assign x_744 = v_1289 | ~v_232 | ~v_1267;
assign x_745 = v_1267 | ~v_232 | ~v_1289;
assign x_746 = v_232 | ~v_1267 | ~v_1289;
assign x_747 = v_230 | v_231 | v_232 | ~v_1264 | ~v_1289;
assign x_748 = v_229 | v_1265 | v_1266 | v_1267 | ~v_1289;
assign x_749 = v_1290 | ~v_495 | ~v_1265;
assign x_750 = v_1265 | ~v_495 | ~v_1290;
assign x_751 = v_495 | ~v_1265 | ~v_1290;
assign x_752 = v_1290 | ~v_496 | ~v_1266;
assign x_753 = v_1266 | ~v_496 | ~v_1290;
assign x_754 = v_496 | ~v_1266 | ~v_1290;
assign x_755 = v_1290 | ~v_497 | ~v_1267;
assign x_756 = v_1267 | ~v_497 | ~v_1290;
assign x_757 = v_497 | ~v_1267 | ~v_1290;
assign x_758 = v_495 | v_496 | v_497 | ~v_1290;
assign x_759 = v_1265 | v_1266 | v_1267 | ~v_1290;
assign x_760 = v_583 | v_1297 | ~v_1298;
assign x_761 = v_1272 | ~v_583 | ~v_1298;
assign x_762 = v_1272 | v_1297 | ~v_1298;
assign x_763 = v_1298 | ~v_1272 | ~v_1297;
assign x_764 = v_1298 | ~v_583 | ~v_1272;
assign x_765 = v_583 | v_1298 | ~v_1297;
assign x_766 = v_1264 | v_1319 | ~v_259;
assign x_767 = v_259 | v_1264 | ~v_1319;
assign x_768 = ~v_259 | ~v_1264 | ~v_1319;
assign x_769 = v_1319 | ~v_260 | ~v_1265;
assign x_770 = v_1265 | ~v_260 | ~v_1319;
assign x_771 = v_260 | ~v_1265 | ~v_1319;
assign x_772 = v_1319 | ~v_261 | ~v_1266;
assign x_773 = v_1266 | ~v_261 | ~v_1319;
assign x_774 = v_261 | ~v_1266 | ~v_1319;
assign x_775 = v_1319 | ~v_262 | ~v_1267;
assign x_776 = v_1267 | ~v_262 | ~v_1319;
assign x_777 = v_262 | ~v_1267 | ~v_1319;
assign x_778 = v_260 | v_261 | v_262 | ~v_1264 | ~v_1319;
assign x_779 = v_259 | v_1265 | v_1266 | v_1267 | ~v_1319;
assign x_780 = v_626 | v_1326 | ~v_1327;
assign x_781 = v_1303 | ~v_626 | ~v_1327;
assign x_782 = v_1303 | v_1326 | ~v_1327;
assign x_783 = v_1327 | ~v_1303 | ~v_1326;
assign x_784 = v_1327 | ~v_626 | ~v_1303;
assign x_785 = v_626 | v_1327 | ~v_1326;
assign x_786 = v_1332 | v_1357 | ~v_229;
assign x_787 = v_229 | v_1332 | ~v_1357;
assign x_788 = ~v_229 | ~v_1332 | ~v_1357;
assign x_789 = v_1357 | ~v_230 | ~v_1333;
assign x_790 = v_1333 | ~v_230 | ~v_1357;
assign x_791 = v_230 | ~v_1333 | ~v_1357;
assign x_792 = v_1357 | ~v_231 | ~v_1334;
assign x_793 = v_1334 | ~v_231 | ~v_1357;
assign x_794 = v_231 | ~v_1334 | ~v_1357;
assign x_795 = v_1357 | ~v_232 | ~v_1335;
assign x_796 = v_1335 | ~v_232 | ~v_1357;
assign x_797 = v_232 | ~v_1335 | ~v_1357;
assign x_798 = v_230 | v_231 | v_232 | ~v_1332 | ~v_1357;
assign x_799 = v_229 | v_1333 | v_1334 | v_1335 | ~v_1357;
assign x_800 = v_1358 | ~v_495 | ~v_1333;
assign x_801 = v_1333 | ~v_495 | ~v_1358;
assign x_802 = v_495 | ~v_1333 | ~v_1358;
assign x_803 = v_1358 | ~v_496 | ~v_1334;
assign x_804 = v_1334 | ~v_496 | ~v_1358;
assign x_805 = v_496 | ~v_1334 | ~v_1358;
assign x_806 = v_1358 | ~v_497 | ~v_1335;
assign x_807 = v_1335 | ~v_497 | ~v_1358;
assign x_808 = v_497 | ~v_1335 | ~v_1358;
assign x_809 = v_495 | v_496 | v_497 | ~v_1358;
assign x_810 = v_1333 | v_1334 | v_1335 | ~v_1358;
assign x_811 = v_583 | v_1365 | ~v_1366;
assign x_812 = v_1340 | ~v_583 | ~v_1366;
assign x_813 = v_1340 | v_1365 | ~v_1366;
assign x_814 = v_1366 | ~v_1340 | ~v_1365;
assign x_815 = v_1366 | ~v_583 | ~v_1340;
assign x_816 = v_583 | v_1366 | ~v_1365;
assign x_817 = v_1332 | v_1387 | ~v_259;
assign x_818 = v_259 | v_1332 | ~v_1387;
assign x_819 = ~v_259 | ~v_1332 | ~v_1387;
assign x_820 = v_1387 | ~v_260 | ~v_1333;
assign x_821 = v_1333 | ~v_260 | ~v_1387;
assign x_822 = v_260 | ~v_1333 | ~v_1387;
assign x_823 = v_1387 | ~v_261 | ~v_1334;
assign x_824 = v_1334 | ~v_261 | ~v_1387;
assign x_825 = v_261 | ~v_1334 | ~v_1387;
assign x_826 = v_1387 | ~v_262 | ~v_1335;
assign x_827 = v_1335 | ~v_262 | ~v_1387;
assign x_828 = v_262 | ~v_1335 | ~v_1387;
assign x_829 = v_260 | v_261 | v_262 | ~v_1332 | ~v_1387;
assign x_830 = v_259 | v_1333 | v_1334 | v_1335 | ~v_1387;
assign x_831 = v_626 | v_1394 | ~v_1395;
assign x_832 = v_1371 | ~v_626 | ~v_1395;
assign x_833 = v_1371 | v_1394 | ~v_1395;
assign x_834 = v_1395 | ~v_1371 | ~v_1394;
assign x_835 = v_1395 | ~v_626 | ~v_1371;
assign x_836 = v_626 | v_1395 | ~v_1394;
assign x_837 = ~v_1399 | ~v_1400;
assign x_838 = ~v_1399 | ~v_1401;
assign x_839 = ~v_1400 | ~v_1401;
assign x_840 = v_1399 | ~v_1262 | ~v_1403;
assign x_841 = v_1262 | v_1400 | ~v_1403;
assign x_842 = v_1399 | v_1400 | ~v_1403;
assign x_843 = v_1403 | ~v_1399 | ~v_1400;
assign x_844 = v_1262 | v_1403 | ~v_1400;
assign x_845 = v_1403 | ~v_1262 | ~v_1399;
assign x_846 = v_1400 | ~v_1262 | ~v_1404;
assign x_847 = v_1262 | v_1401 | ~v_1404;
assign x_848 = v_1400 | v_1401 | ~v_1404;
assign x_849 = v_1404 | ~v_1400 | ~v_1401;
assign x_850 = v_1262 | v_1404 | ~v_1401;
assign x_851 = v_1404 | ~v_1262 | ~v_1400;
assign x_852 = ~v_1402 | ~v_1403;
assign x_853 = ~v_1402 | ~v_1404;
assign x_854 = ~v_1402 | ~v_1405;
assign x_855 = ~v_1403 | ~v_1404;
assign x_856 = ~v_1403 | ~v_1405;
assign x_857 = ~v_1404 | ~v_1405;
assign x_858 = v_1402 | ~v_1194 | ~v_1407;
assign x_859 = v_1194 | v_1403 | ~v_1407;
assign x_860 = v_1402 | v_1403 | ~v_1407;
assign x_861 = v_1407 | ~v_1402 | ~v_1403;
assign x_862 = v_1194 | v_1407 | ~v_1403;
assign x_863 = v_1407 | ~v_1194 | ~v_1402;
assign x_864 = v_1403 | ~v_1194 | ~v_1408;
assign x_865 = v_1194 | v_1404 | ~v_1408;
assign x_866 = v_1403 | v_1404 | ~v_1408;
assign x_867 = v_1408 | ~v_1403 | ~v_1404;
assign x_868 = v_1194 | v_1408 | ~v_1404;
assign x_869 = v_1408 | ~v_1194 | ~v_1403;
assign x_870 = v_1404 | ~v_1194 | ~v_1409;
assign x_871 = v_1194 | v_1405 | ~v_1409;
assign x_872 = v_1404 | v_1405 | ~v_1409;
assign x_873 = v_1409 | ~v_1404 | ~v_1405;
assign x_874 = v_1194 | v_1409 | ~v_1405;
assign x_875 = v_1409 | ~v_1194 | ~v_1404;
assign x_876 = ~v_1406 | ~v_1407;
assign x_877 = ~v_1406 | ~v_1408;
assign x_878 = ~v_1406 | ~v_1409;
assign x_879 = ~v_1406 | ~v_1410;
assign x_880 = ~v_1407 | ~v_1408;
assign x_881 = ~v_1407 | ~v_1409;
assign x_882 = ~v_1407 | ~v_1410;
assign x_883 = ~v_1408 | ~v_1409;
assign x_884 = ~v_1408 | ~v_1410;
assign x_885 = ~v_1409 | ~v_1410;
assign x_886 = v_1411 | ~v_491 | ~v_1407;
assign x_887 = v_1407 | ~v_491 | ~v_1411;
assign x_888 = v_491 | ~v_1407 | ~v_1411;
assign x_889 = v_1411 | ~v_492 | ~v_1408;
assign x_890 = v_1408 | ~v_492 | ~v_1411;
assign x_891 = v_492 | ~v_1408 | ~v_1411;
assign x_892 = v_1411 | ~v_493 | ~v_1409;
assign x_893 = v_1409 | ~v_493 | ~v_1411;
assign x_894 = v_493 | ~v_1409 | ~v_1411;
assign x_895 = v_1411 | ~v_494 | ~v_1410;
assign x_896 = v_1410 | ~v_494 | ~v_1411;
assign x_897 = v_494 | ~v_1410 | ~v_1411;
assign x_898 = v_491 | v_492 | v_493 | v_494 | ~v_1411;
assign x_899 = v_1407 | v_1408 | v_1409 | v_1410 | ~v_1411;
assign x_900 = v_1069 | v_1398 | ~v_1418;
assign x_901 = ~v_1398 | ~v_1417 | ~v_1418;
assign x_902 = v_1069 | ~v_1417 | ~v_1418;
assign x_903 = v_1417 | v_1418 | ~v_1069;
assign x_904 = v_1417 | v_1418 | ~v_1398;
assign x_905 = v_1398 | v_1418 | ~v_1069;
assign x_906 = v_1418 | ~v_1330 | ~v_1421;
assign x_907 = v_1330 | ~v_1417 | ~v_1421;
assign x_908 = v_1418 | ~v_1417 | ~v_1421;
assign x_909 = v_1417 | v_1421 | ~v_1418;
assign x_910 = v_1330 | v_1417 | v_1421;
assign x_911 = v_1421 | ~v_1330 | ~v_1418;
assign x_912 = v_1419 | ~v_1330 | ~v_1422;
assign x_913 = v_1330 | v_1417 | ~v_1422;
assign x_914 = v_1417 | v_1419 | ~v_1422;
assign x_915 = v_1422 | ~v_1417 | ~v_1419;
assign x_916 = v_1330 | v_1422 | ~v_1417;
assign x_917 = v_1422 | ~v_1330 | ~v_1419;
assign x_918 = v_1087 | ~v_1399 | ~v_1424;
assign x_919 = v_1399 | v_1421 | ~v_1424;
assign x_920 = v_1087 | v_1421 | ~v_1424;
assign x_921 = v_1424 | ~v_1087 | ~v_1421;
assign x_922 = v_1399 | v_1424 | ~v_1421;
assign x_923 = v_1424 | ~v_1087 | ~v_1399;
assign x_924 = v_1424 | ~v_1262 | ~v_1428;
assign x_925 = v_1262 | v_1421 | ~v_1428;
assign x_926 = v_1421 | v_1424 | ~v_1428;
assign x_927 = v_1428 | ~v_1421 | ~v_1424;
assign x_928 = v_1262 | v_1428 | ~v_1421;
assign x_929 = v_1428 | ~v_1262 | ~v_1424;
assign x_930 = v_1425 | ~v_1262 | ~v_1429;
assign x_931 = v_1262 | v_1422 | ~v_1429;
assign x_932 = v_1422 | v_1425 | ~v_1429;
assign x_933 = v_1429 | ~v_1422 | ~v_1425;
assign x_934 = v_1262 | v_1429 | ~v_1422;
assign x_935 = v_1429 | ~v_1262 | ~v_1425;
assign x_936 = v_1426 | ~v_1262 | ~v_1430;
assign x_937 = v_1262 | v_1423 | ~v_1430;
assign x_938 = v_1423 | v_1426 | ~v_1430;
assign x_939 = v_1430 | ~v_1423 | ~v_1426;
assign x_940 = v_1262 | v_1430 | ~v_1423;
assign x_941 = v_1430 | ~v_1262 | ~v_1426;
assign x_942 = v_1107 | ~v_1402 | ~v_1432;
assign x_943 = v_1402 | v_1428 | ~v_1432;
assign x_944 = v_1107 | v_1428 | ~v_1432;
assign x_945 = v_1432 | ~v_1107 | ~v_1428;
assign x_946 = v_1402 | v_1432 | ~v_1428;
assign x_947 = v_1432 | ~v_1107 | ~v_1402;
assign x_948 = v_1432 | ~v_1194 | ~v_1437;
assign x_949 = v_1194 | v_1428 | ~v_1437;
assign x_950 = v_1428 | v_1432 | ~v_1437;
assign x_951 = v_1437 | ~v_1428 | ~v_1432;
assign x_952 = v_1194 | v_1437 | ~v_1428;
assign x_953 = v_1437 | ~v_1194 | ~v_1432;
assign x_954 = v_1433 | ~v_1194 | ~v_1438;
assign x_955 = v_1194 | v_1429 | ~v_1438;
assign x_956 = v_1429 | v_1433 | ~v_1438;
assign x_957 = v_1438 | ~v_1429 | ~v_1433;
assign x_958 = v_1194 | v_1438 | ~v_1429;
assign x_959 = v_1438 | ~v_1194 | ~v_1433;
assign x_960 = v_1434 | ~v_1194 | ~v_1439;
assign x_961 = v_1194 | v_1430 | ~v_1439;
assign x_962 = v_1430 | v_1434 | ~v_1439;
assign x_963 = v_1439 | ~v_1430 | ~v_1434;
assign x_964 = v_1194 | v_1439 | ~v_1430;
assign x_965 = v_1439 | ~v_1194 | ~v_1434;
assign x_966 = v_1435 | ~v_1194 | ~v_1440;
assign x_967 = v_1194 | v_1431 | ~v_1440;
assign x_968 = v_1431 | v_1435 | ~v_1440;
assign x_969 = v_1440 | ~v_1431 | ~v_1435;
assign x_970 = v_1194 | v_1440 | ~v_1431;
assign x_971 = v_1440 | ~v_1194 | ~v_1435;
assign x_972 = v_1470 | v_1506 | v_1513;
assign x_973 = v_1506 | ~v_1470 | ~v_1513;
assign x_974 = v_1470 | ~v_1506 | ~v_1513;
assign x_975 = v_1472 | v_1508 | v_1513;
assign x_976 = v_1508 | ~v_1472 | ~v_1513;
assign x_977 = v_1472 | ~v_1508 | ~v_1513;
assign x_978 = v_1474 | v_1510 | v_1513;
assign x_979 = v_1510 | ~v_1474 | ~v_1513;
assign x_980 = v_1474 | ~v_1510 | ~v_1513;
assign x_981 = v_1476 | v_1512 | v_1513;
assign x_982 = v_1512 | ~v_1476 | ~v_1513;
assign x_983 = v_1476 | ~v_1512 | ~v_1513;
assign x_984 = ~v_1506 | ~v_1508 | ~v_1510 | ~v_1512 | ~v_1513;
assign x_985 = ~v_1470 | ~v_1472 | ~v_1474 | ~v_1476 | ~v_1513;
assign x_986 = v_1087 | ~v_1400 | ~v_1526;
assign x_987 = v_1400 | ~v_1525 | ~v_1526;
assign x_988 = v_1087 | ~v_1525 | ~v_1526;
assign x_989 = v_1525 | v_1526 | ~v_1087;
assign x_990 = v_1400 | v_1525 | v_1526;
assign x_991 = v_1526 | ~v_1087 | ~v_1400;
assign x_992 = v_1526 | ~v_1262 | ~v_1529;
assign x_993 = v_1262 | ~v_1525 | ~v_1529;
assign x_994 = v_1526 | ~v_1525 | ~v_1529;
assign x_995 = v_1525 | v_1529 | ~v_1526;
assign x_996 = v_1262 | v_1525 | v_1529;
assign x_997 = v_1529 | ~v_1262 | ~v_1526;
assign x_998 = v_1527 | ~v_1262 | ~v_1530;
assign x_999 = v_1262 | v_1525 | ~v_1530;
assign x_1000 = v_1525 | v_1527 | ~v_1530;
assign x_1001 = v_1530 | ~v_1525 | ~v_1527;
assign x_1002 = v_1262 | v_1530 | ~v_1525;
assign x_1003 = v_1530 | ~v_1262 | ~v_1527;
assign x_1004 = v_1107 | ~v_1403 | ~v_1532;
assign x_1005 = v_1403 | v_1529 | ~v_1532;
assign x_1006 = v_1107 | v_1529 | ~v_1532;
assign x_1007 = v_1532 | ~v_1107 | ~v_1529;
assign x_1008 = v_1403 | v_1532 | ~v_1529;
assign x_1009 = v_1532 | ~v_1107 | ~v_1403;
assign x_1010 = v_1532 | ~v_1194 | ~v_1536;
assign x_1011 = v_1194 | v_1529 | ~v_1536;
assign x_1012 = v_1529 | v_1532 | ~v_1536;
assign x_1013 = v_1536 | ~v_1529 | ~v_1532;
assign x_1014 = v_1194 | v_1536 | ~v_1529;
assign x_1015 = v_1536 | ~v_1194 | ~v_1532;
assign x_1016 = v_1533 | ~v_1194 | ~v_1537;
assign x_1017 = v_1194 | v_1530 | ~v_1537;
assign x_1018 = v_1530 | v_1533 | ~v_1537;
assign x_1019 = v_1537 | ~v_1530 | ~v_1533;
assign x_1020 = v_1194 | v_1537 | ~v_1530;
assign x_1021 = v_1537 | ~v_1194 | ~v_1533;
assign x_1022 = v_1534 | ~v_1194 | ~v_1538;
assign x_1023 = v_1194 | v_1531 | ~v_1538;
assign x_1024 = v_1531 | v_1534 | ~v_1538;
assign x_1025 = v_1538 | ~v_1531 | ~v_1534;
assign x_1026 = v_1194 | v_1538 | ~v_1531;
assign x_1027 = v_1538 | ~v_1194 | ~v_1534;
assign x_1028 = v_1559 | v_1596 | v_1603;
assign x_1029 = v_1596 | ~v_1559 | ~v_1603;
assign x_1030 = v_1559 | ~v_1596 | ~v_1603;
assign x_1031 = v_1561 | v_1598 | v_1603;
assign x_1032 = v_1598 | ~v_1561 | ~v_1603;
assign x_1033 = v_1561 | ~v_1598 | ~v_1603;
assign x_1034 = v_1563 | v_1600 | v_1603;
assign x_1035 = v_1600 | ~v_1563 | ~v_1603;
assign x_1036 = v_1563 | ~v_1600 | ~v_1603;
assign x_1037 = v_1565 | v_1602 | v_1603;
assign x_1038 = v_1602 | ~v_1565 | ~v_1603;
assign x_1039 = v_1565 | ~v_1602 | ~v_1603;
assign x_1040 = ~v_1596 | ~v_1598 | ~v_1600 | ~v_1602 | ~v_1603;
assign x_1041 = ~v_1559 | ~v_1561 | ~v_1563 | ~v_1565 | ~v_1603;
assign x_1042 = v_491 | ~v_1604 | ~v_1605;
assign x_1043 = ~v_491 | ~v_1514 | ~v_1605;
assign x_1044 = ~v_1514 | ~v_1604 | ~v_1605;
assign x_1045 = v_1514 | v_1604 | v_1605;
assign x_1046 = v_1514 | v_1605 | ~v_491;
assign x_1047 = v_491 | v_1604 | v_1605;
assign x_1048 = v_1107 | ~v_1404 | ~v_1617;
assign x_1049 = v_1404 | ~v_1616 | ~v_1617;
assign x_1050 = v_1107 | ~v_1616 | ~v_1617;
assign x_1051 = v_1616 | v_1617 | ~v_1107;
assign x_1052 = v_1404 | v_1616 | v_1617;
assign x_1053 = v_1617 | ~v_1107 | ~v_1404;
assign x_1054 = v_1617 | ~v_1194 | ~v_1620;
assign x_1055 = v_1194 | ~v_1616 | ~v_1620;
assign x_1056 = v_1617 | ~v_1616 | ~v_1620;
assign x_1057 = v_1616 | v_1620 | ~v_1617;
assign x_1058 = v_1194 | v_1616 | v_1620;
assign x_1059 = v_1620 | ~v_1194 | ~v_1617;
assign x_1060 = v_1618 | ~v_1194 | ~v_1621;
assign x_1061 = v_1194 | v_1616 | ~v_1621;
assign x_1062 = v_1616 | v_1618 | ~v_1621;
assign x_1063 = v_1621 | ~v_1616 | ~v_1618;
assign x_1064 = v_1194 | v_1621 | ~v_1616;
assign x_1065 = v_1621 | ~v_1194 | ~v_1618;
assign x_1066 = v_1633 | v_1670 | v_1677;
assign x_1067 = v_1670 | ~v_1633 | ~v_1677;
assign x_1068 = v_1633 | ~v_1670 | ~v_1677;
assign x_1069 = v_1635 | v_1672 | v_1677;
assign x_1070 = v_1672 | ~v_1635 | ~v_1677;
assign x_1071 = v_1635 | ~v_1672 | ~v_1677;
assign x_1072 = v_1637 | v_1674 | v_1677;
assign x_1073 = v_1674 | ~v_1637 | ~v_1677;
assign x_1074 = v_1637 | ~v_1674 | ~v_1677;
assign x_1075 = v_1639 | v_1676 | v_1677;
assign x_1076 = v_1676 | ~v_1639 | ~v_1677;
assign x_1077 = v_1639 | ~v_1676 | ~v_1677;
assign x_1078 = ~v_1670 | ~v_1672 | ~v_1674 | ~v_1676 | ~v_1677;
assign x_1079 = ~v_1633 | ~v_1635 | ~v_1637 | ~v_1639 | ~v_1677;
assign x_1080 = ~v_963 | ~v_1678 | ~v_1679;
assign x_1081 = v_963 | v_1605 | ~v_1679;
assign x_1082 = v_1605 | ~v_1678 | ~v_1679;
assign x_1083 = v_1678 | v_1679 | ~v_1605;
assign x_1084 = v_963 | v_1679 | ~v_1605;
assign x_1085 = v_1678 | v_1679 | ~v_963;
assign x_1086 = v_1693 | v_1719 | v_1726;
assign x_1087 = v_1719 | ~v_1693 | ~v_1726;
assign x_1088 = v_1693 | ~v_1719 | ~v_1726;
assign x_1089 = v_1721 | v_1726 | ~v_1694;
assign x_1090 = v_1694 | v_1721 | ~v_1726;
assign x_1091 = ~v_1694 | ~v_1721 | ~v_1726;
assign x_1092 = v_1723 | v_1726 | ~v_1695;
assign x_1093 = v_1695 | v_1723 | ~v_1726;
assign x_1094 = ~v_1695 | ~v_1723 | ~v_1726;
assign x_1095 = v_1725 | v_1726 | ~v_1696;
assign x_1096 = v_1696 | v_1725 | ~v_1726;
assign x_1097 = ~v_1696 | ~v_1725 | ~v_1726;
assign x_1098 = ~v_1719 | ~v_1721 | ~v_1723 | ~v_1725 | ~v_1726;
assign x_1099 = v_1694 | v_1695 | v_1696 | ~v_1693 | ~v_1726;
assign x_1100 = ~v_494 | ~v_1727 | ~v_1728;
assign x_1101 = v_494 | v_1679 | ~v_1728;
assign x_1102 = v_1679 | ~v_1727 | ~v_1728;
assign x_1103 = v_1727 | v_1728 | ~v_1679;
assign x_1104 = v_494 | v_1728 | ~v_1679;
assign x_1105 = v_1727 | v_1728 | ~v_494;
assign x_1106 = v_491 | ~v_1022 | ~v_1745;
assign x_1107 = v_492 | v_1022 | ~v_1745;
assign x_1108 = v_491 | v_492 | ~v_1745;
assign x_1109 = v_1745 | ~v_491 | ~v_492;
assign x_1110 = v_1022 | v_1745 | ~v_492;
assign x_1111 = v_1745 | ~v_491 | ~v_1022;
assign x_1112 = v_492 | ~v_1022 | ~v_1746;
assign x_1113 = v_493 | v_1022 | ~v_1746;
assign x_1114 = v_492 | v_493 | ~v_1746;
assign x_1115 = v_1746 | ~v_492 | ~v_493;
assign x_1116 = v_1022 | v_1746 | ~v_493;
assign x_1117 = v_1746 | ~v_492 | ~v_1022;
assign x_1118 = v_493 | ~v_1022 | ~v_1747;
assign x_1119 = v_494 | v_1022 | ~v_1747;
assign x_1120 = v_493 | v_494 | ~v_1747;
assign x_1121 = v_1747 | ~v_493 | ~v_494;
assign x_1122 = v_1022 | v_1747 | ~v_494;
assign x_1123 = v_1747 | ~v_493 | ~v_1022;
assign x_1124 = v_1744 | ~v_4 | ~v_1749;
assign x_1125 = v_4 | v_525 | ~v_1749;
assign x_1126 = v_525 | v_1744 | ~v_1749;
assign x_1127 = v_1749 | ~v_525 | ~v_1744;
assign x_1128 = v_4 | v_1749 | ~v_525;
assign x_1129 = v_1749 | ~v_4 | ~v_1744;
assign x_1130 = v_1745 | ~v_4 | ~v_1750;
assign x_1131 = v_4 | v_526 | ~v_1750;
assign x_1132 = v_526 | v_1745 | ~v_1750;
assign x_1133 = v_1750 | ~v_526 | ~v_1745;
assign x_1134 = v_4 | v_1750 | ~v_526;
assign x_1135 = v_1750 | ~v_4 | ~v_1745;
assign x_1136 = v_1746 | ~v_4 | ~v_1751;
assign x_1137 = v_4 | v_527 | ~v_1751;
assign x_1138 = v_527 | v_1746 | ~v_1751;
assign x_1139 = v_1751 | ~v_527 | ~v_1746;
assign x_1140 = v_4 | v_1751 | ~v_527;
assign x_1141 = v_1751 | ~v_4 | ~v_1746;
assign x_1142 = v_1747 | ~v_4 | ~v_1752;
assign x_1143 = v_4 | v_528 | ~v_1752;
assign x_1144 = v_528 | v_1747 | ~v_1752;
assign x_1145 = v_1752 | ~v_528 | ~v_1747;
assign x_1146 = v_4 | v_1752 | ~v_528;
assign x_1147 = v_1752 | ~v_4 | ~v_1747;
assign x_1148 = ~v_1749 | ~v_1750;
assign x_1149 = ~v_1749 | ~v_1751;
assign x_1150 = ~v_1749 | ~v_1752;
assign x_1151 = ~v_1749 | ~v_1753;
assign x_1152 = ~v_1750 | ~v_1751;
assign x_1153 = ~v_1750 | ~v_1752;
assign x_1154 = ~v_1750 | ~v_1753;
assign x_1155 = ~v_1751 | ~v_1752;
assign x_1156 = ~v_1751 | ~v_1753;
assign x_1157 = ~v_1752 | ~v_1753;
assign x_1158 = v_1753 | ~v_1769 | ~v_1770;
assign x_1159 = ~v_1753 | ~v_1755 | ~v_1770;
assign x_1160 = ~v_1755 | ~v_1769 | ~v_1770;
assign x_1161 = v_1755 | v_1769 | v_1770;
assign x_1162 = v_1755 | v_1770 | ~v_1753;
assign x_1163 = v_1753 | v_1769 | v_1770;
assign x_1164 = v_1756 | ~v_1771 | ~v_1772;
assign x_1165 = v_1770 | ~v_1756 | ~v_1772;
assign x_1166 = v_1770 | ~v_1771 | ~v_1772;
assign x_1167 = v_1771 | v_1772 | ~v_1770;
assign x_1168 = v_1772 | ~v_1756 | ~v_1770;
assign x_1169 = v_1756 | v_1771 | v_1772;
assign x_1170 = v_1753 | ~v_1785 | ~v_1786;
assign x_1171 = ~v_1753 | ~v_1756 | ~v_1786;
assign x_1172 = ~v_1756 | ~v_1785 | ~v_1786;
assign x_1173 = v_1756 | v_1785 | v_1786;
assign x_1174 = v_1756 | v_1786 | ~v_1753;
assign x_1175 = v_1753 | v_1785 | v_1786;
assign x_1176 = v_1756 | ~v_1787 | ~v_1788;
assign x_1177 = v_1786 | ~v_1756 | ~v_1788;
assign x_1178 = v_1786 | ~v_1787 | ~v_1788;
assign x_1179 = v_1787 | v_1788 | ~v_1786;
assign x_1180 = v_1788 | ~v_1756 | ~v_1786;
assign x_1181 = v_1756 | v_1787 | v_1788;
assign x_1182 = v_1755 | ~v_1789 | ~v_1790;
assign x_1183 = v_1788 | ~v_1755 | ~v_1790;
assign x_1184 = v_1788 | ~v_1789 | ~v_1790;
assign x_1185 = v_1789 | v_1790 | ~v_1788;
assign x_1186 = v_1790 | ~v_1755 | ~v_1788;
assign x_1187 = v_1755 | v_1789 | v_1790;
assign x_1188 = v_1753 | ~v_1803 | ~v_1804;
assign x_1189 = ~v_1753 | ~v_1804;
assign x_1190 = ~v_1753 | ~v_1803 | ~v_1804;
assign x_1191 = v_1753 | v_1803 | v_1804;
assign x_1192 = v_1753 | v_1803 | v_1804;
assign x_1193 = v_1756 | ~v_1805 | ~v_1806;
assign x_1194 = v_1804 | ~v_1756 | ~v_1806;
assign x_1195 = v_1804 | ~v_1805 | ~v_1806;
assign x_1196 = v_1805 | v_1806 | ~v_1804;
assign x_1197 = v_1806 | ~v_1756 | ~v_1804;
assign x_1198 = v_1756 | v_1805 | v_1806;
assign x_1199 = v_1755 | ~v_1807 | ~v_1808;
assign x_1200 = v_1806 | ~v_1755 | ~v_1808;
assign x_1201 = v_1806 | ~v_1807 | ~v_1808;
assign x_1202 = v_1807 | v_1808 | ~v_1806;
assign x_1203 = v_1808 | ~v_1755 | ~v_1806;
assign x_1204 = v_1755 | v_1807 | v_1808;
assign x_1205 = ~v_1749 | ~v_1809 | ~v_1810;
assign x_1206 = v_1749 | v_1808 | ~v_1810;
assign x_1207 = v_1808 | ~v_1809 | ~v_1810;
assign x_1208 = v_1809 | v_1810 | ~v_1808;
assign x_1209 = v_1749 | v_1810 | ~v_1808;
assign x_1210 = v_1809 | v_1810 | ~v_1749;
assign x_1211 = v_1823 | v_1848 | ~v_229;
assign x_1212 = v_229 | v_1823 | ~v_1848;
assign x_1213 = ~v_229 | ~v_1823 | ~v_1848;
assign x_1214 = v_1848 | ~v_230 | ~v_1824;
assign x_1215 = v_1824 | ~v_230 | ~v_1848;
assign x_1216 = v_230 | ~v_1824 | ~v_1848;
assign x_1217 = v_1848 | ~v_231 | ~v_1825;
assign x_1218 = v_1825 | ~v_231 | ~v_1848;
assign x_1219 = v_231 | ~v_1825 | ~v_1848;
assign x_1220 = v_1848 | ~v_232 | ~v_1826;
assign x_1221 = v_1826 | ~v_232 | ~v_1848;
assign x_1222 = v_232 | ~v_1826 | ~v_1848;
assign x_1223 = v_230 | v_231 | v_232 | ~v_1823 | ~v_1848;
assign x_1224 = v_229 | v_1824 | v_1825 | v_1826 | ~v_1848;
assign x_1225 = v_1823 | v_1849 | ~v_495;
assign x_1226 = v_495 | v_1823 | ~v_1849;
assign x_1227 = ~v_495 | ~v_1823 | ~v_1849;
assign x_1228 = v_1849 | ~v_496 | ~v_1824;
assign x_1229 = v_1824 | ~v_496 | ~v_1849;
assign x_1230 = v_496 | ~v_1824 | ~v_1849;
assign x_1231 = v_1849 | ~v_497 | ~v_1825;
assign x_1232 = v_1825 | ~v_497 | ~v_1849;
assign x_1233 = v_497 | ~v_1825 | ~v_1849;
assign x_1234 = v_1849 | ~v_498 | ~v_1826;
assign x_1235 = v_1826 | ~v_498 | ~v_1849;
assign x_1236 = v_498 | ~v_1826 | ~v_1849;
assign x_1237 = v_496 | v_497 | v_498 | ~v_1823 | ~v_1849;
assign x_1238 = v_495 | v_1824 | v_1825 | v_1826 | ~v_1849;
assign x_1239 = v_583 | v_1856 | ~v_1857;
assign x_1240 = v_1831 | ~v_583 | ~v_1857;
assign x_1241 = v_1831 | v_1856 | ~v_1857;
assign x_1242 = v_1857 | ~v_1831 | ~v_1856;
assign x_1243 = v_1857 | ~v_583 | ~v_1831;
assign x_1244 = v_583 | v_1857 | ~v_1856;
assign x_1245 = v_1823 | v_1878 | ~v_259;
assign x_1246 = v_259 | v_1823 | ~v_1878;
assign x_1247 = ~v_259 | ~v_1823 | ~v_1878;
assign x_1248 = v_1878 | ~v_260 | ~v_1824;
assign x_1249 = v_1824 | ~v_260 | ~v_1878;
assign x_1250 = v_260 | ~v_1824 | ~v_1878;
assign x_1251 = v_1878 | ~v_261 | ~v_1825;
assign x_1252 = v_1825 | ~v_261 | ~v_1878;
assign x_1253 = v_261 | ~v_1825 | ~v_1878;
assign x_1254 = v_1878 | ~v_262 | ~v_1826;
assign x_1255 = v_1826 | ~v_262 | ~v_1878;
assign x_1256 = v_262 | ~v_1826 | ~v_1878;
assign x_1257 = v_260 | v_261 | v_262 | ~v_1823 | ~v_1878;
assign x_1258 = v_259 | v_1824 | v_1825 | v_1826 | ~v_1878;
assign x_1259 = v_626 | v_1885 | ~v_1886;
assign x_1260 = v_1862 | ~v_626 | ~v_1886;
assign x_1261 = v_1862 | v_1885 | ~v_1886;
assign x_1262 = v_1886 | ~v_1862 | ~v_1885;
assign x_1263 = v_1886 | ~v_626 | ~v_1862;
assign x_1264 = v_626 | v_1886 | ~v_1885;
assign x_1265 = v_1891 | v_1916 | ~v_229;
assign x_1266 = v_229 | v_1891 | ~v_1916;
assign x_1267 = ~v_229 | ~v_1891 | ~v_1916;
assign x_1268 = v_1916 | ~v_230 | ~v_1892;
assign x_1269 = v_1892 | ~v_230 | ~v_1916;
assign x_1270 = v_230 | ~v_1892 | ~v_1916;
assign x_1271 = v_1916 | ~v_231 | ~v_1893;
assign x_1272 = v_1893 | ~v_231 | ~v_1916;
assign x_1273 = v_231 | ~v_1893 | ~v_1916;
assign x_1274 = v_1916 | ~v_232 | ~v_1894;
assign x_1275 = v_1894 | ~v_232 | ~v_1916;
assign x_1276 = v_232 | ~v_1894 | ~v_1916;
assign x_1277 = v_230 | v_231 | v_232 | ~v_1891 | ~v_1916;
assign x_1278 = v_229 | v_1892 | v_1893 | v_1894 | ~v_1916;
assign x_1279 = v_1891 | v_1917 | ~v_495;
assign x_1280 = v_495 | v_1891 | ~v_1917;
assign x_1281 = ~v_495 | ~v_1891 | ~v_1917;
assign x_1282 = v_1917 | ~v_496 | ~v_1892;
assign x_1283 = v_1892 | ~v_496 | ~v_1917;
assign x_1284 = v_496 | ~v_1892 | ~v_1917;
assign x_1285 = v_1917 | ~v_497 | ~v_1893;
assign x_1286 = v_1893 | ~v_497 | ~v_1917;
assign x_1287 = v_497 | ~v_1893 | ~v_1917;
assign x_1288 = v_1917 | ~v_498 | ~v_1894;
assign x_1289 = v_1894 | ~v_498 | ~v_1917;
assign x_1290 = v_498 | ~v_1894 | ~v_1917;
assign x_1291 = v_496 | v_497 | v_498 | ~v_1891 | ~v_1917;
assign x_1292 = v_495 | v_1892 | v_1893 | v_1894 | ~v_1917;
assign x_1293 = v_583 | v_1924 | ~v_1925;
assign x_1294 = v_1899 | ~v_583 | ~v_1925;
assign x_1295 = v_1899 | v_1924 | ~v_1925;
assign x_1296 = v_1925 | ~v_1899 | ~v_1924;
assign x_1297 = v_1925 | ~v_583 | ~v_1899;
assign x_1298 = v_583 | v_1925 | ~v_1924;
assign x_1299 = v_1891 | v_1946 | ~v_259;
assign x_1300 = v_259 | v_1891 | ~v_1946;
assign x_1301 = ~v_259 | ~v_1891 | ~v_1946;
assign x_1302 = v_1946 | ~v_260 | ~v_1892;
assign x_1303 = v_1892 | ~v_260 | ~v_1946;
assign x_1304 = v_260 | ~v_1892 | ~v_1946;
assign x_1305 = v_1946 | ~v_261 | ~v_1893;
assign x_1306 = v_1893 | ~v_261 | ~v_1946;
assign x_1307 = v_261 | ~v_1893 | ~v_1946;
assign x_1308 = v_1946 | ~v_262 | ~v_1894;
assign x_1309 = v_1894 | ~v_262 | ~v_1946;
assign x_1310 = v_262 | ~v_1894 | ~v_1946;
assign x_1311 = v_260 | v_261 | v_262 | ~v_1891 | ~v_1946;
assign x_1312 = v_259 | v_1892 | v_1893 | v_1894 | ~v_1946;
assign x_1313 = v_626 | v_1953 | ~v_1954;
assign x_1314 = v_1930 | ~v_626 | ~v_1954;
assign x_1315 = v_1930 | v_1953 | ~v_1954;
assign x_1316 = v_1954 | ~v_1930 | ~v_1953;
assign x_1317 = v_1954 | ~v_626 | ~v_1930;
assign x_1318 = v_626 | v_1954 | ~v_1953;
assign x_1319 = v_1959 | v_1984 | ~v_229;
assign x_1320 = v_229 | v_1959 | ~v_1984;
assign x_1321 = ~v_229 | ~v_1959 | ~v_1984;
assign x_1322 = v_1984 | ~v_230 | ~v_1960;
assign x_1323 = v_1960 | ~v_230 | ~v_1984;
assign x_1324 = v_230 | ~v_1960 | ~v_1984;
assign x_1325 = v_1984 | ~v_231 | ~v_1961;
assign x_1326 = v_1961 | ~v_231 | ~v_1984;
assign x_1327 = v_231 | ~v_1961 | ~v_1984;
assign x_1328 = v_1984 | ~v_232 | ~v_1962;
assign x_1329 = v_1962 | ~v_232 | ~v_1984;
assign x_1330 = v_232 | ~v_1962 | ~v_1984;
assign x_1331 = v_230 | v_231 | v_232 | ~v_1959 | ~v_1984;
assign x_1332 = v_229 | v_1960 | v_1961 | v_1962 | ~v_1984;
assign x_1333 = v_1959 | v_1985 | ~v_495;
assign x_1334 = v_495 | v_1959 | ~v_1985;
assign x_1335 = ~v_495 | ~v_1959 | ~v_1985;
assign x_1336 = v_1985 | ~v_496 | ~v_1960;
assign x_1337 = v_1960 | ~v_496 | ~v_1985;
assign x_1338 = v_496 | ~v_1960 | ~v_1985;
assign x_1339 = v_1985 | ~v_497 | ~v_1961;
assign x_1340 = v_1961 | ~v_497 | ~v_1985;
assign x_1341 = v_497 | ~v_1961 | ~v_1985;
assign x_1342 = v_1985 | ~v_498 | ~v_1962;
assign x_1343 = v_1962 | ~v_498 | ~v_1985;
assign x_1344 = v_498 | ~v_1962 | ~v_1985;
assign x_1345 = v_496 | v_497 | v_498 | ~v_1959 | ~v_1985;
assign x_1346 = v_495 | v_1960 | v_1961 | v_1962 | ~v_1985;
assign x_1347 = v_583 | v_1992 | ~v_1993;
assign x_1348 = v_1967 | ~v_583 | ~v_1993;
assign x_1349 = v_1967 | v_1992 | ~v_1993;
assign x_1350 = v_1993 | ~v_1967 | ~v_1992;
assign x_1351 = v_1993 | ~v_583 | ~v_1967;
assign x_1352 = v_583 | v_1993 | ~v_1992;
assign x_1353 = v_1959 | v_2014 | ~v_259;
assign x_1354 = v_259 | v_1959 | ~v_2014;
assign x_1355 = ~v_259 | ~v_1959 | ~v_2014;
assign x_1356 = v_2014 | ~v_260 | ~v_1960;
assign x_1357 = v_1960 | ~v_260 | ~v_2014;
assign x_1358 = v_260 | ~v_1960 | ~v_2014;
assign x_1359 = v_2014 | ~v_261 | ~v_1961;
assign x_1360 = v_1961 | ~v_261 | ~v_2014;
assign x_1361 = v_261 | ~v_1961 | ~v_2014;
assign x_1362 = v_2014 | ~v_262 | ~v_1962;
assign x_1363 = v_1962 | ~v_262 | ~v_2014;
assign x_1364 = v_262 | ~v_1962 | ~v_2014;
assign x_1365 = v_260 | v_261 | v_262 | ~v_1959 | ~v_2014;
assign x_1366 = v_259 | v_1960 | v_1961 | v_1962 | ~v_2014;
assign x_1367 = v_626 | v_2021 | ~v_2022;
assign x_1368 = v_1998 | ~v_626 | ~v_2022;
assign x_1369 = v_1998 | v_2021 | ~v_2022;
assign x_1370 = v_2022 | ~v_1998 | ~v_2021;
assign x_1371 = v_2022 | ~v_626 | ~v_1998;
assign x_1372 = v_626 | v_2022 | ~v_2021;
assign x_1373 = v_2027 | v_2052 | ~v_229;
assign x_1374 = v_229 | v_2027 | ~v_2052;
assign x_1375 = ~v_229 | ~v_2027 | ~v_2052;
assign x_1376 = v_2052 | ~v_230 | ~v_2028;
assign x_1377 = v_2028 | ~v_230 | ~v_2052;
assign x_1378 = v_230 | ~v_2028 | ~v_2052;
assign x_1379 = v_2052 | ~v_231 | ~v_2029;
assign x_1380 = v_2029 | ~v_231 | ~v_2052;
assign x_1381 = v_231 | ~v_2029 | ~v_2052;
assign x_1382 = v_2052 | ~v_232 | ~v_2030;
assign x_1383 = v_2030 | ~v_232 | ~v_2052;
assign x_1384 = v_232 | ~v_2030 | ~v_2052;
assign x_1385 = v_230 | v_231 | v_232 | ~v_2027 | ~v_2052;
assign x_1386 = v_229 | v_2028 | v_2029 | v_2030 | ~v_2052;
assign x_1387 = v_2027 | v_2053 | ~v_495;
assign x_1388 = v_495 | v_2027 | ~v_2053;
assign x_1389 = ~v_495 | ~v_2027 | ~v_2053;
assign x_1390 = v_2053 | ~v_496 | ~v_2028;
assign x_1391 = v_2028 | ~v_496 | ~v_2053;
assign x_1392 = v_496 | ~v_2028 | ~v_2053;
assign x_1393 = v_2053 | ~v_497 | ~v_2029;
assign x_1394 = v_2029 | ~v_497 | ~v_2053;
assign x_1395 = v_497 | ~v_2029 | ~v_2053;
assign x_1396 = v_2053 | ~v_498 | ~v_2030;
assign x_1397 = v_2030 | ~v_498 | ~v_2053;
assign x_1398 = v_498 | ~v_2030 | ~v_2053;
assign x_1399 = v_496 | v_497 | v_498 | ~v_2027 | ~v_2053;
assign x_1400 = v_495 | v_2028 | v_2029 | v_2030 | ~v_2053;
assign x_1401 = v_583 | v_2060 | ~v_2061;
assign x_1402 = v_2035 | ~v_583 | ~v_2061;
assign x_1403 = v_2035 | v_2060 | ~v_2061;
assign x_1404 = v_2061 | ~v_2035 | ~v_2060;
assign x_1405 = v_2061 | ~v_583 | ~v_2035;
assign x_1406 = v_583 | v_2061 | ~v_2060;
assign x_1407 = v_2027 | v_2082 | ~v_259;
assign x_1408 = v_259 | v_2027 | ~v_2082;
assign x_1409 = ~v_259 | ~v_2027 | ~v_2082;
assign x_1410 = v_2082 | ~v_260 | ~v_2028;
assign x_1411 = v_2028 | ~v_260 | ~v_2082;
assign x_1412 = v_260 | ~v_2028 | ~v_2082;
assign x_1413 = v_2082 | ~v_261 | ~v_2029;
assign x_1414 = v_2029 | ~v_261 | ~v_2082;
assign x_1415 = v_261 | ~v_2029 | ~v_2082;
assign x_1416 = v_2082 | ~v_262 | ~v_2030;
assign x_1417 = v_2030 | ~v_262 | ~v_2082;
assign x_1418 = v_262 | ~v_2030 | ~v_2082;
assign x_1419 = v_260 | v_261 | v_262 | ~v_2027 | ~v_2082;
assign x_1420 = v_259 | v_2028 | v_2029 | v_2030 | ~v_2082;
assign x_1421 = v_626 | v_2089 | ~v_2090;
assign x_1422 = v_2066 | ~v_626 | ~v_2090;
assign x_1423 = v_2066 | v_2089 | ~v_2090;
assign x_1424 = v_2090 | ~v_2066 | ~v_2089;
assign x_1425 = v_2090 | ~v_626 | ~v_2066;
assign x_1426 = v_626 | v_2090 | ~v_2089;
assign x_1427 = ~v_2094 | ~v_2095;
assign x_1428 = ~v_2094 | ~v_2096;
assign x_1429 = ~v_2095 | ~v_2096;
assign x_1430 = v_2094 | ~v_1957 | ~v_2098;
assign x_1431 = v_1957 | v_2095 | ~v_2098;
assign x_1432 = v_2094 | v_2095 | ~v_2098;
assign x_1433 = v_2098 | ~v_2094 | ~v_2095;
assign x_1434 = v_1957 | v_2098 | ~v_2095;
assign x_1435 = v_2098 | ~v_1957 | ~v_2094;
assign x_1436 = v_2095 | ~v_1957 | ~v_2099;
assign x_1437 = v_1957 | v_2096 | ~v_2099;
assign x_1438 = v_2095 | v_2096 | ~v_2099;
assign x_1439 = v_2099 | ~v_2095 | ~v_2096;
assign x_1440 = v_1957 | v_2099 | ~v_2096;
assign x_1441 = v_2099 | ~v_1957 | ~v_2095;
assign x_1442 = ~v_2097 | ~v_2098;
assign x_1443 = ~v_2097 | ~v_2099;
assign x_1444 = ~v_2097 | ~v_2100;
assign x_1445 = ~v_2098 | ~v_2099;
assign x_1446 = ~v_2098 | ~v_2100;
assign x_1447 = ~v_2099 | ~v_2100;
assign x_1448 = v_2097 | ~v_1889 | ~v_2102;
assign x_1449 = v_1889 | v_2098 | ~v_2102;
assign x_1450 = v_2097 | v_2098 | ~v_2102;
assign x_1451 = v_2102 | ~v_2097 | ~v_2098;
assign x_1452 = v_1889 | v_2102 | ~v_2098;
assign x_1453 = v_2102 | ~v_1889 | ~v_2097;
assign x_1454 = v_2098 | ~v_1889 | ~v_2103;
assign x_1455 = v_1889 | v_2099 | ~v_2103;
assign x_1456 = v_2098 | v_2099 | ~v_2103;
assign x_1457 = v_2103 | ~v_2098 | ~v_2099;
assign x_1458 = v_1889 | v_2103 | ~v_2099;
assign x_1459 = v_2103 | ~v_1889 | ~v_2098;
assign x_1460 = v_2099 | ~v_1889 | ~v_2104;
assign x_1461 = v_1889 | v_2100 | ~v_2104;
assign x_1462 = v_2099 | v_2100 | ~v_2104;
assign x_1463 = v_2104 | ~v_2099 | ~v_2100;
assign x_1464 = v_1889 | v_2104 | ~v_2100;
assign x_1465 = v_2104 | ~v_1889 | ~v_2099;
assign x_1466 = ~v_2101 | ~v_2102;
assign x_1467 = ~v_2101 | ~v_2103;
assign x_1468 = ~v_2101 | ~v_2104;
assign x_1469 = ~v_2101 | ~v_2105;
assign x_1470 = ~v_2102 | ~v_2103;
assign x_1471 = ~v_2102 | ~v_2104;
assign x_1472 = ~v_2102 | ~v_2105;
assign x_1473 = ~v_2103 | ~v_2104;
assign x_1474 = ~v_2103 | ~v_2105;
assign x_1475 = ~v_2104 | ~v_2105;
assign x_1476 = v_2106 | ~v_1744 | ~v_2101;
assign x_1477 = v_2101 | ~v_1744 | ~v_2106;
assign x_1478 = v_1744 | ~v_2101 | ~v_2106;
assign x_1479 = v_2106 | ~v_1745 | ~v_2102;
assign x_1480 = v_2102 | ~v_1745 | ~v_2106;
assign x_1481 = v_1745 | ~v_2102 | ~v_2106;
assign x_1482 = v_2106 | ~v_1746 | ~v_2103;
assign x_1483 = v_2103 | ~v_1746 | ~v_2106;
assign x_1484 = v_1746 | ~v_2103 | ~v_2106;
assign x_1485 = v_2106 | ~v_1747 | ~v_2104;
assign x_1486 = v_2104 | ~v_1747 | ~v_2106;
assign x_1487 = v_1747 | ~v_2104 | ~v_2106;
assign x_1488 = v_2106 | ~v_1748 | ~v_2105;
assign x_1489 = v_2105 | ~v_1748 | ~v_2106;
assign x_1490 = v_1748 | ~v_2105 | ~v_2106;
assign x_1491 = v_1744 | v_1745 | v_1746 | v_1747 | v_1748 | ~v_2106;
assign x_1492 = v_2101 | v_2102 | v_2103 | v_2104 | v_2105 | ~v_2106;
assign x_1493 = v_1772 | v_2093 | ~v_2110;
assign x_1494 = ~v_2093 | ~v_2109 | ~v_2110;
assign x_1495 = v_1772 | ~v_2109 | ~v_2110;
assign x_1496 = v_2109 | v_2110 | ~v_1772;
assign x_1497 = v_2109 | v_2110 | ~v_2093;
assign x_1498 = v_2093 | v_2110 | ~v_1772;
assign x_1499 = v_2110 | ~v_2025 | ~v_2113;
assign x_1500 = v_2025 | ~v_2109 | ~v_2113;
assign x_1501 = v_2110 | ~v_2109 | ~v_2113;
assign x_1502 = v_2109 | v_2113 | ~v_2110;
assign x_1503 = v_2025 | v_2109 | v_2113;
assign x_1504 = v_2113 | ~v_2025 | ~v_2110;
assign x_1505 = v_2111 | ~v_2025 | ~v_2114;
assign x_1506 = v_2025 | v_2109 | ~v_2114;
assign x_1507 = v_2109 | v_2111 | ~v_2114;
assign x_1508 = v_2114 | ~v_2109 | ~v_2111;
assign x_1509 = v_2025 | v_2114 | ~v_2109;
assign x_1510 = v_2114 | ~v_2025 | ~v_2111;
assign x_1511 = v_1790 | ~v_2094 | ~v_2116;
assign x_1512 = v_2094 | v_2113 | ~v_2116;
assign x_1513 = v_1790 | v_2113 | ~v_2116;
assign x_1514 = v_2116 | ~v_1790 | ~v_2113;
assign x_1515 = v_2094 | v_2116 | ~v_2113;
assign x_1516 = v_2116 | ~v_1790 | ~v_2094;
assign x_1517 = v_2116 | ~v_1957 | ~v_2120;
assign x_1518 = v_1957 | v_2113 | ~v_2120;
assign x_1519 = v_2113 | v_2116 | ~v_2120;
assign x_1520 = v_2120 | ~v_2113 | ~v_2116;
assign x_1521 = v_1957 | v_2120 | ~v_2113;
assign x_1522 = v_2120 | ~v_1957 | ~v_2116;
assign x_1523 = v_2117 | ~v_1957 | ~v_2121;
assign x_1524 = v_1957 | v_2114 | ~v_2121;
assign x_1525 = v_2114 | v_2117 | ~v_2121;
assign x_1526 = v_2121 | ~v_2114 | ~v_2117;
assign x_1527 = v_1957 | v_2121 | ~v_2114;
assign x_1528 = v_2121 | ~v_1957 | ~v_2117;
assign x_1529 = v_2118 | ~v_1957 | ~v_2122;
assign x_1530 = v_1957 | v_2115 | ~v_2122;
assign x_1531 = v_2115 | v_2118 | ~v_2122;
assign x_1532 = v_2122 | ~v_2115 | ~v_2118;
assign x_1533 = v_1957 | v_2122 | ~v_2115;
assign x_1534 = v_2122 | ~v_1957 | ~v_2118;
assign x_1535 = v_1810 | ~v_2097 | ~v_2124;
assign x_1536 = v_2097 | v_2120 | ~v_2124;
assign x_1537 = v_1810 | v_2120 | ~v_2124;
assign x_1538 = v_2124 | ~v_1810 | ~v_2120;
assign x_1539 = v_2097 | v_2124 | ~v_2120;
assign x_1540 = v_2124 | ~v_1810 | ~v_2097;
assign x_1541 = v_2124 | ~v_1889 | ~v_2129;
assign x_1542 = v_1889 | v_2120 | ~v_2129;
assign x_1543 = v_2120 | v_2124 | ~v_2129;
assign x_1544 = v_2129 | ~v_2120 | ~v_2124;
assign x_1545 = v_1889 | v_2129 | ~v_2120;
assign x_1546 = v_2129 | ~v_1889 | ~v_2124;
assign x_1547 = v_2125 | ~v_1889 | ~v_2130;
assign x_1548 = v_1889 | v_2121 | ~v_2130;
assign x_1549 = v_2121 | v_2125 | ~v_2130;
assign x_1550 = v_2130 | ~v_2121 | ~v_2125;
assign x_1551 = v_1889 | v_2130 | ~v_2121;
assign x_1552 = v_2130 | ~v_1889 | ~v_2125;
assign x_1553 = v_2126 | ~v_1889 | ~v_2131;
assign x_1554 = v_1889 | v_2122 | ~v_2131;
assign x_1555 = v_2122 | v_2126 | ~v_2131;
assign x_1556 = v_2131 | ~v_2122 | ~v_2126;
assign x_1557 = v_1889 | v_2131 | ~v_2122;
assign x_1558 = v_2131 | ~v_1889 | ~v_2126;
assign x_1559 = v_2127 | ~v_1889 | ~v_2132;
assign x_1560 = v_1889 | v_2123 | ~v_2132;
assign x_1561 = v_2123 | v_2127 | ~v_2132;
assign x_1562 = v_2132 | ~v_2123 | ~v_2127;
assign x_1563 = v_1889 | v_2132 | ~v_2123;
assign x_1564 = v_2132 | ~v_1889 | ~v_2127;
assign x_1565 = v_2162 | v_2169 | ~v_659;
assign x_1566 = v_659 | v_2162 | ~v_2169;
assign x_1567 = ~v_659 | ~v_2162 | ~v_2169;
assign x_1568 = v_2164 | v_2169 | ~v_660;
assign x_1569 = v_660 | v_2164 | ~v_2169;
assign x_1570 = ~v_660 | ~v_2164 | ~v_2169;
assign x_1571 = v_2166 | v_2169 | ~v_661;
assign x_1572 = v_661 | v_2166 | ~v_2169;
assign x_1573 = ~v_661 | ~v_2166 | ~v_2169;
assign x_1574 = v_2168 | v_2169 | ~v_662;
assign x_1575 = v_662 | v_2168 | ~v_2169;
assign x_1576 = ~v_662 | ~v_2168 | ~v_2169;
assign x_1577 = ~v_2162 | ~v_2164 | ~v_2166 | ~v_2168 | ~v_2169;
assign x_1578 = v_659 | v_660 | v_661 | v_662 | ~v_2169;
assign x_1579 = v_1744 | ~v_2170 | ~v_2171;
assign x_1580 = ~v_1744 | ~v_2106 | ~v_2171;
assign x_1581 = ~v_2106 | ~v_2170 | ~v_2171;
assign x_1582 = v_2106 | v_2170 | v_2171;
assign x_1583 = v_2106 | v_2171 | ~v_1744;
assign x_1584 = v_1744 | v_2170 | v_2171;
assign x_1585 = v_1790 | ~v_2095 | ~v_2177;
assign x_1586 = v_2095 | ~v_2176 | ~v_2177;
assign x_1587 = v_1790 | ~v_2176 | ~v_2177;
assign x_1588 = v_2176 | v_2177 | ~v_1790;
assign x_1589 = v_2095 | v_2176 | v_2177;
assign x_1590 = v_2177 | ~v_1790 | ~v_2095;
assign x_1591 = v_2177 | ~v_1957 | ~v_2180;
assign x_1592 = v_1957 | ~v_2176 | ~v_2180;
assign x_1593 = v_2177 | ~v_2176 | ~v_2180;
assign x_1594 = v_2176 | v_2180 | ~v_2177;
assign x_1595 = v_1957 | v_2176 | v_2180;
assign x_1596 = v_2180 | ~v_1957 | ~v_2177;
assign x_1597 = v_2178 | ~v_1957 | ~v_2181;
assign x_1598 = v_1957 | v_2176 | ~v_2181;
assign x_1599 = v_2176 | v_2178 | ~v_2181;
assign x_1600 = v_2181 | ~v_2176 | ~v_2178;
assign x_1601 = v_1957 | v_2181 | ~v_2176;
assign x_1602 = v_2181 | ~v_1957 | ~v_2178;
assign x_1603 = v_1810 | ~v_2098 | ~v_2183;
assign x_1604 = v_2098 | v_2180 | ~v_2183;
assign x_1605 = v_1810 | v_2180 | ~v_2183;
assign x_1606 = v_2183 | ~v_1810 | ~v_2180;
assign x_1607 = v_2098 | v_2183 | ~v_2180;
assign x_1608 = v_2183 | ~v_1810 | ~v_2098;
assign x_1609 = v_2183 | ~v_1889 | ~v_2187;
assign x_1610 = v_1889 | v_2180 | ~v_2187;
assign x_1611 = v_2180 | v_2183 | ~v_2187;
assign x_1612 = v_2187 | ~v_2180 | ~v_2183;
assign x_1613 = v_1889 | v_2187 | ~v_2180;
assign x_1614 = v_2187 | ~v_1889 | ~v_2183;
assign x_1615 = v_2184 | ~v_1889 | ~v_2188;
assign x_1616 = v_1889 | v_2181 | ~v_2188;
assign x_1617 = v_2181 | v_2184 | ~v_2188;
assign x_1618 = v_2188 | ~v_2181 | ~v_2184;
assign x_1619 = v_1889 | v_2188 | ~v_2181;
assign x_1620 = v_2188 | ~v_1889 | ~v_2184;
assign x_1621 = v_2185 | ~v_1889 | ~v_2189;
assign x_1622 = v_1889 | v_2182 | ~v_2189;
assign x_1623 = v_2182 | v_2185 | ~v_2189;
assign x_1624 = v_2189 | ~v_2182 | ~v_2185;
assign x_1625 = v_1889 | v_2189 | ~v_2182;
assign x_1626 = v_2189 | ~v_1889 | ~v_2185;
assign x_1627 = v_2210 | v_2217 | ~v_663;
assign x_1628 = v_663 | v_2210 | ~v_2217;
assign x_1629 = ~v_663 | ~v_2210 | ~v_2217;
assign x_1630 = v_2212 | v_2217 | ~v_664;
assign x_1631 = v_664 | v_2212 | ~v_2217;
assign x_1632 = ~v_664 | ~v_2212 | ~v_2217;
assign x_1633 = v_2214 | v_2217 | ~v_665;
assign x_1634 = v_665 | v_2214 | ~v_2217;
assign x_1635 = ~v_665 | ~v_2214 | ~v_2217;
assign x_1636 = v_2216 | v_2217 | ~v_666;
assign x_1637 = v_666 | v_2216 | ~v_2217;
assign x_1638 = ~v_666 | ~v_2216 | ~v_2217;
assign x_1639 = ~v_2210 | ~v_2212 | ~v_2214 | ~v_2216 | ~v_2217;
assign x_1640 = v_663 | v_664 | v_665 | v_666 | ~v_2217;
assign x_1641 = ~v_2172 | ~v_2218 | ~v_2219;
assign x_1642 = v_2171 | v_2172 | ~v_2219;
assign x_1643 = v_2171 | ~v_2218 | ~v_2219;
assign x_1644 = v_2218 | v_2219 | ~v_2171;
assign x_1645 = v_2172 | v_2219 | ~v_2171;
assign x_1646 = v_2218 | v_2219 | ~v_2172;
assign x_1647 = v_1810 | ~v_2099 | ~v_2225;
assign x_1648 = v_2099 | ~v_2224 | ~v_2225;
assign x_1649 = v_1810 | ~v_2224 | ~v_2225;
assign x_1650 = v_2224 | v_2225 | ~v_1810;
assign x_1651 = v_2099 | v_2224 | v_2225;
assign x_1652 = v_2225 | ~v_1810 | ~v_2099;
assign x_1653 = v_2225 | ~v_1889 | ~v_2228;
assign x_1654 = v_1889 | ~v_2224 | ~v_2228;
assign x_1655 = v_2225 | ~v_2224 | ~v_2228;
assign x_1656 = v_2224 | v_2228 | ~v_2225;
assign x_1657 = v_1889 | v_2224 | v_2228;
assign x_1658 = v_2228 | ~v_1889 | ~v_2225;
assign x_1659 = v_2226 | ~v_1889 | ~v_2229;
assign x_1660 = v_1889 | v_2224 | ~v_2229;
assign x_1661 = v_2224 | v_2226 | ~v_2229;
assign x_1662 = v_2229 | ~v_2224 | ~v_2226;
assign x_1663 = v_1889 | v_2229 | ~v_2224;
assign x_1664 = v_2229 | ~v_1889 | ~v_2226;
assign x_1665 = v_2241 | v_2248 | ~v_667;
assign x_1666 = v_667 | v_2241 | ~v_2248;
assign x_1667 = ~v_667 | ~v_2241 | ~v_2248;
assign x_1668 = v_2243 | v_2248 | ~v_668;
assign x_1669 = v_668 | v_2243 | ~v_2248;
assign x_1670 = ~v_668 | ~v_2243 | ~v_2248;
assign x_1671 = v_2245 | v_2248 | ~v_669;
assign x_1672 = v_669 | v_2245 | ~v_2248;
assign x_1673 = ~v_669 | ~v_2245 | ~v_2248;
assign x_1674 = v_2247 | v_2248 | ~v_670;
assign x_1675 = v_670 | v_2247 | ~v_2248;
assign x_1676 = ~v_670 | ~v_2247 | ~v_2248;
assign x_1677 = ~v_2241 | ~v_2243 | ~v_2245 | ~v_2247 | ~v_2248;
assign x_1678 = v_667 | v_668 | v_669 | v_670 | ~v_2248;
assign x_1679 = ~v_2220 | ~v_2249 | ~v_2250;
assign x_1680 = v_2219 | v_2220 | ~v_2250;
assign x_1681 = v_2219 | ~v_2249 | ~v_2250;
assign x_1682 = v_2249 | v_2250 | ~v_2219;
assign x_1683 = v_2220 | v_2250 | ~v_2219;
assign x_1684 = v_2249 | v_2250 | ~v_2220;
assign x_1685 = v_2259 | v_2263 | ~v_671;
assign x_1686 = v_671 | v_2259 | ~v_2263;
assign x_1687 = ~v_671 | ~v_2259 | ~v_2263;
assign x_1688 = v_2263 | ~v_672 | ~v_2260;
assign x_1689 = v_2260 | ~v_672 | ~v_2263;
assign x_1690 = v_672 | ~v_2260 | ~v_2263;
assign x_1691 = v_2263 | ~v_673 | ~v_2261;
assign x_1692 = v_2261 | ~v_673 | ~v_2263;
assign x_1693 = v_673 | ~v_2261 | ~v_2263;
assign x_1694 = v_2263 | ~v_674 | ~v_2262;
assign x_1695 = v_2262 | ~v_674 | ~v_2263;
assign x_1696 = v_674 | ~v_2262 | ~v_2263;
assign x_1697 = v_672 | v_673 | v_674 | ~v_2259 | ~v_2263;
assign x_1698 = v_671 | v_2260 | v_2261 | v_2262 | ~v_2263;
assign x_1699 = ~v_1748 | ~v_2264 | ~v_2265;
assign x_1700 = v_1748 | v_2250 | ~v_2265;
assign x_1701 = v_2250 | ~v_2264 | ~v_2265;
assign x_1702 = v_2264 | v_2265 | ~v_2250;
assign x_1703 = v_1748 | v_2265 | ~v_2250;
assign x_1704 = v_2264 | v_2265 | ~v_1748;
assign x_1705 = v_504 | ~v_2280;
assign x_1706 = v_2279 | ~v_504 | ~v_2280;
assign x_1707 = v_504 | v_2279 | ~v_2280;
assign x_1708 = v_2280 | ~v_504 | ~v_2279;
assign x_1709 = v_2280 | ~v_504 | ~v_2279;
assign x_1710 = ~v_2289 | ~v_2302;
assign x_1711 = ~v_2289 | ~v_2303;
assign x_1712 = ~v_2289 | ~v_2304;
assign x_1713 = ~v_2289 | ~v_2305;
assign x_1714 = ~v_2302 | ~v_2303;
assign x_1715 = ~v_2302 | ~v_2304;
assign x_1716 = ~v_2302 | ~v_2305;
assign x_1717 = ~v_2303 | ~v_2304;
assign x_1718 = ~v_2303 | ~v_2305;
assign x_1719 = ~v_2304 | ~v_2305;
assign x_1720 = v_2289 | ~v_2333 | ~v_2334;
assign x_1721 = ~v_2289 | ~v_2307 | ~v_2334;
assign x_1722 = ~v_2307 | ~v_2333 | ~v_2334;
assign x_1723 = v_2307 | v_2333 | v_2334;
assign x_1724 = v_2307 | v_2334 | ~v_2289;
assign x_1725 = v_2289 | v_2333 | v_2334;
assign x_1726 = v_2308 | ~v_2335 | ~v_2336;
assign x_1727 = v_2334 | ~v_2308 | ~v_2336;
assign x_1728 = v_2334 | ~v_2335 | ~v_2336;
assign x_1729 = v_2335 | v_2336 | ~v_2334;
assign x_1730 = v_2336 | ~v_2308 | ~v_2334;
assign x_1731 = v_2308 | v_2335 | v_2336;
assign x_1732 = v_2289 | ~v_2361 | ~v_2362;
assign x_1733 = ~v_2289 | ~v_2308 | ~v_2362;
assign x_1734 = ~v_2308 | ~v_2361 | ~v_2362;
assign x_1735 = v_2308 | v_2361 | v_2362;
assign x_1736 = v_2308 | v_2362 | ~v_2289;
assign x_1737 = v_2289 | v_2361 | v_2362;
assign x_1738 = v_2308 | ~v_2363 | ~v_2364;
assign x_1739 = v_2362 | ~v_2308 | ~v_2364;
assign x_1740 = v_2362 | ~v_2363 | ~v_2364;
assign x_1741 = v_2363 | v_2364 | ~v_2362;
assign x_1742 = v_2364 | ~v_2308 | ~v_2362;
assign x_1743 = v_2308 | v_2363 | v_2364;
assign x_1744 = v_2307 | ~v_2365 | ~v_2366;
assign x_1745 = v_2364 | ~v_2307 | ~v_2366;
assign x_1746 = v_2364 | ~v_2365 | ~v_2366;
assign x_1747 = v_2365 | v_2366 | ~v_2364;
assign x_1748 = v_2366 | ~v_2307 | ~v_2364;
assign x_1749 = v_2307 | v_2365 | v_2366;
assign x_1750 = v_2289 | ~v_2391 | ~v_2392;
assign x_1751 = ~v_2289 | ~v_2392;
assign x_1752 = ~v_2289 | ~v_2391 | ~v_2392;
assign x_1753 = v_2289 | v_2391 | v_2392;
assign x_1754 = v_2289 | v_2391 | v_2392;
assign x_1755 = v_2308 | ~v_2393 | ~v_2394;
assign x_1756 = v_2392 | ~v_2308 | ~v_2394;
assign x_1757 = v_2392 | ~v_2393 | ~v_2394;
assign x_1758 = v_2393 | v_2394 | ~v_2392;
assign x_1759 = v_2394 | ~v_2308 | ~v_2392;
assign x_1760 = v_2308 | v_2393 | v_2394;
assign x_1761 = v_2307 | ~v_2395 | ~v_2396;
assign x_1762 = v_2394 | ~v_2307 | ~v_2396;
assign x_1763 = v_2394 | ~v_2395 | ~v_2396;
assign x_1764 = v_2395 | v_2396 | ~v_2394;
assign x_1765 = v_2396 | ~v_2307 | ~v_2394;
assign x_1766 = v_2307 | v_2395 | v_2396;
assign x_1767 = ~v_2302 | ~v_2397 | ~v_2398;
assign x_1768 = v_2302 | v_2396 | ~v_2398;
assign x_1769 = v_2396 | ~v_2397 | ~v_2398;
assign x_1770 = v_2397 | v_2398 | ~v_2396;
assign x_1771 = v_2302 | v_2398 | ~v_2396;
assign x_1772 = v_2397 | v_2398 | ~v_2302;
assign x_1773 = v_2452 | ~v_425 | ~v_584;
assign x_1774 = v_584 | ~v_425 | ~v_2452;
assign x_1775 = v_425 | ~v_584 | ~v_2452;
assign x_1776 = v_2452 | ~v_426 | ~v_585;
assign x_1777 = v_585 | ~v_426 | ~v_2452;
assign x_1778 = v_426 | ~v_585 | ~v_2452;
assign x_1779 = v_2452 | ~v_427 | ~v_586;
assign x_1780 = v_586 | ~v_427 | ~v_2452;
assign x_1781 = v_427 | ~v_586 | ~v_2452;
assign x_1782 = v_2452 | ~v_428 | ~v_587;
assign x_1783 = v_587 | ~v_428 | ~v_2452;
assign x_1784 = v_428 | ~v_587 | ~v_2452;
assign x_1785 = v_425 | v_426 | v_427 | v_428 | ~v_2452;
assign x_1786 = v_584 | v_585 | v_586 | v_587 | ~v_2452;
assign x_1787 = v_2453 | ~v_584 | ~v_2281;
assign x_1788 = v_2281 | ~v_584 | ~v_2453;
assign x_1789 = v_584 | ~v_2281 | ~v_2453;
assign x_1790 = v_2453 | ~v_585 | ~v_2282;
assign x_1791 = v_2282 | ~v_585 | ~v_2453;
assign x_1792 = v_585 | ~v_2282 | ~v_2453;
assign x_1793 = v_2453 | ~v_586 | ~v_2283;
assign x_1794 = v_2283 | ~v_586 | ~v_2453;
assign x_1795 = v_586 | ~v_2283 | ~v_2453;
assign x_1796 = v_2453 | ~v_587 | ~v_2284;
assign x_1797 = v_2284 | ~v_587 | ~v_2453;
assign x_1798 = v_587 | ~v_2284 | ~v_2453;
assign x_1799 = v_584 | v_585 | v_586 | v_587 | ~v_2453;
assign x_1800 = v_2281 | v_2282 | v_2283 | v_2284 | ~v_2453;
assign x_1801 = v_2429 | v_2461 | ~v_2462;
assign x_1802 = v_2435 | ~v_2429 | ~v_2462;
assign x_1803 = v_2435 | v_2461 | ~v_2462;
assign x_1804 = v_2462 | ~v_2435 | ~v_2461;
assign x_1805 = v_2462 | ~v_2429 | ~v_2435;
assign x_1806 = v_2429 | v_2462 | ~v_2461;
assign x_1807 = v_2493 | ~v_455 | ~v_584;
assign x_1808 = v_584 | ~v_455 | ~v_2493;
assign x_1809 = v_455 | ~v_584 | ~v_2493;
assign x_1810 = v_2493 | ~v_456 | ~v_585;
assign x_1811 = v_585 | ~v_456 | ~v_2493;
assign x_1812 = v_456 | ~v_585 | ~v_2493;
assign x_1813 = v_2493 | ~v_457 | ~v_586;
assign x_1814 = v_586 | ~v_457 | ~v_2493;
assign x_1815 = v_457 | ~v_586 | ~v_2493;
assign x_1816 = v_2493 | ~v_458 | ~v_587;
assign x_1817 = v_587 | ~v_458 | ~v_2493;
assign x_1818 = v_458 | ~v_587 | ~v_2493;
assign x_1819 = v_455 | v_456 | v_457 | v_458 | ~v_2493;
assign x_1820 = v_584 | v_585 | v_586 | v_587 | ~v_2493;
assign x_1821 = v_2470 | v_2501 | ~v_2502;
assign x_1822 = v_2476 | ~v_2470 | ~v_2502;
assign x_1823 = v_2476 | v_2501 | ~v_2502;
assign x_1824 = v_2502 | ~v_2476 | ~v_2501;
assign x_1825 = v_2502 | ~v_2470 | ~v_2476;
assign x_1826 = v_2470 | v_2502 | ~v_2501;
assign x_1827 = v_2505 | v_2530 | ~v_425;
assign x_1828 = v_425 | v_2505 | ~v_2530;
assign x_1829 = ~v_425 | ~v_2505 | ~v_2530;
assign x_1830 = v_2530 | ~v_426 | ~v_2506;
assign x_1831 = v_2506 | ~v_426 | ~v_2530;
assign x_1832 = v_426 | ~v_2506 | ~v_2530;
assign x_1833 = v_2530 | ~v_427 | ~v_2507;
assign x_1834 = v_2507 | ~v_427 | ~v_2530;
assign x_1835 = v_427 | ~v_2507 | ~v_2530;
assign x_1836 = v_2530 | ~v_428 | ~v_2508;
assign x_1837 = v_2508 | ~v_428 | ~v_2530;
assign x_1838 = v_428 | ~v_2508 | ~v_2530;
assign x_1839 = v_426 | v_427 | v_428 | ~v_2505 | ~v_2530;
assign x_1840 = v_425 | v_2506 | v_2507 | v_2508 | ~v_2530;
assign x_1841 = v_2505 | v_2531 | ~v_495;
assign x_1842 = v_495 | v_2505 | ~v_2531;
assign x_1843 = ~v_495 | ~v_2505 | ~v_2531;
assign x_1844 = v_2531 | ~v_496 | ~v_2506;
assign x_1845 = v_2506 | ~v_496 | ~v_2531;
assign x_1846 = v_496 | ~v_2506 | ~v_2531;
assign x_1847 = v_2531 | ~v_497 | ~v_2507;
assign x_1848 = v_2507 | ~v_497 | ~v_2531;
assign x_1849 = v_497 | ~v_2507 | ~v_2531;
assign x_1850 = v_2531 | ~v_498 | ~v_2508;
assign x_1851 = v_2508 | ~v_498 | ~v_2531;
assign x_1852 = v_498 | ~v_2508 | ~v_2531;
assign x_1853 = v_496 | v_497 | v_498 | ~v_2505 | ~v_2531;
assign x_1854 = v_495 | v_2506 | v_2507 | v_2508 | ~v_2531;
assign x_1855 = v_2505 | v_2532 | ~v_2281;
assign x_1856 = v_2281 | v_2505 | ~v_2532;
assign x_1857 = ~v_2281 | ~v_2505 | ~v_2532;
assign x_1858 = v_2532 | ~v_2282 | ~v_2506;
assign x_1859 = v_2506 | ~v_2282 | ~v_2532;
assign x_1860 = v_2282 | ~v_2506 | ~v_2532;
assign x_1861 = v_2532 | ~v_2283 | ~v_2507;
assign x_1862 = v_2507 | ~v_2283 | ~v_2532;
assign x_1863 = v_2283 | ~v_2507 | ~v_2532;
assign x_1864 = v_2532 | ~v_2284 | ~v_2508;
assign x_1865 = v_2508 | ~v_2284 | ~v_2532;
assign x_1866 = v_2284 | ~v_2508 | ~v_2532;
assign x_1867 = v_2282 | v_2283 | v_2284 | ~v_2505 | ~v_2532;
assign x_1868 = v_2281 | v_2506 | v_2507 | v_2508 | ~v_2532;
assign x_1869 = v_2505 | v_2533 | ~v_584;
assign x_1870 = v_584 | v_2505 | ~v_2533;
assign x_1871 = ~v_584 | ~v_2505 | ~v_2533;
assign x_1872 = v_2533 | ~v_585 | ~v_2506;
assign x_1873 = v_2506 | ~v_585 | ~v_2533;
assign x_1874 = v_585 | ~v_2506 | ~v_2533;
assign x_1875 = v_2533 | ~v_586 | ~v_2507;
assign x_1876 = v_2507 | ~v_586 | ~v_2533;
assign x_1877 = v_586 | ~v_2507 | ~v_2533;
assign x_1878 = v_2533 | ~v_587 | ~v_2508;
assign x_1879 = v_2508 | ~v_587 | ~v_2533;
assign x_1880 = v_587 | ~v_2508 | ~v_2533;
assign x_1881 = v_585 | v_586 | v_587 | ~v_2505 | ~v_2533;
assign x_1882 = v_584 | v_2506 | v_2507 | v_2508 | ~v_2533;
assign x_1883 = v_2429 | v_2542 | ~v_2543;
assign x_1884 = v_2513 | ~v_2429 | ~v_2543;
assign x_1885 = v_2513 | v_2542 | ~v_2543;
assign x_1886 = v_2543 | ~v_2513 | ~v_2542;
assign x_1887 = v_2543 | ~v_2429 | ~v_2513;
assign x_1888 = v_2429 | v_2543 | ~v_2542;
assign x_1889 = v_2505 | v_2564 | ~v_455;
assign x_1890 = v_455 | v_2505 | ~v_2564;
assign x_1891 = ~v_455 | ~v_2505 | ~v_2564;
assign x_1892 = v_2564 | ~v_456 | ~v_2506;
assign x_1893 = v_2506 | ~v_456 | ~v_2564;
assign x_1894 = v_456 | ~v_2506 | ~v_2564;
assign x_1895 = v_2564 | ~v_457 | ~v_2507;
assign x_1896 = v_2507 | ~v_457 | ~v_2564;
assign x_1897 = v_457 | ~v_2507 | ~v_2564;
assign x_1898 = v_2564 | ~v_458 | ~v_2508;
assign x_1899 = v_2508 | ~v_458 | ~v_2564;
assign x_1900 = v_458 | ~v_2508 | ~v_2564;
assign x_1901 = v_456 | v_457 | v_458 | ~v_2505 | ~v_2564;
assign x_1902 = v_455 | v_2506 | v_2507 | v_2508 | ~v_2564;
assign x_1903 = v_2470 | v_2573 | ~v_2574;
assign x_1904 = v_2548 | ~v_2470 | ~v_2574;
assign x_1905 = v_2548 | v_2573 | ~v_2574;
assign x_1906 = v_2574 | ~v_2548 | ~v_2573;
assign x_1907 = v_2574 | ~v_2470 | ~v_2548;
assign x_1908 = v_2470 | v_2574 | ~v_2573;
assign x_1909 = v_2579 | v_2604 | ~v_425;
assign x_1910 = v_425 | v_2579 | ~v_2604;
assign x_1911 = ~v_425 | ~v_2579 | ~v_2604;
assign x_1912 = v_2604 | ~v_426 | ~v_2580;
assign x_1913 = v_2580 | ~v_426 | ~v_2604;
assign x_1914 = v_426 | ~v_2580 | ~v_2604;
assign x_1915 = v_2604 | ~v_427 | ~v_2581;
assign x_1916 = v_2581 | ~v_427 | ~v_2604;
assign x_1917 = v_427 | ~v_2581 | ~v_2604;
assign x_1918 = v_2604 | ~v_428 | ~v_2582;
assign x_1919 = v_2582 | ~v_428 | ~v_2604;
assign x_1920 = v_428 | ~v_2582 | ~v_2604;
assign x_1921 = v_426 | v_427 | v_428 | ~v_2579 | ~v_2604;
assign x_1922 = v_425 | v_2580 | v_2581 | v_2582 | ~v_2604;
assign x_1923 = v_2579 | v_2605 | ~v_495;
assign x_1924 = v_495 | v_2579 | ~v_2605;
assign x_1925 = ~v_495 | ~v_2579 | ~v_2605;
assign x_1926 = v_2605 | ~v_496 | ~v_2580;
assign x_1927 = v_2580 | ~v_496 | ~v_2605;
assign x_1928 = v_496 | ~v_2580 | ~v_2605;
assign x_1929 = v_2605 | ~v_497 | ~v_2581;
assign x_1930 = v_2581 | ~v_497 | ~v_2605;
assign x_1931 = v_497 | ~v_2581 | ~v_2605;
assign x_1932 = v_2605 | ~v_498 | ~v_2582;
assign x_1933 = v_2582 | ~v_498 | ~v_2605;
assign x_1934 = v_498 | ~v_2582 | ~v_2605;
assign x_1935 = v_496 | v_497 | v_498 | ~v_2579 | ~v_2605;
assign x_1936 = v_495 | v_2580 | v_2581 | v_2582 | ~v_2605;
assign x_1937 = v_2579 | v_2606 | ~v_2281;
assign x_1938 = v_2281 | v_2579 | ~v_2606;
assign x_1939 = ~v_2281 | ~v_2579 | ~v_2606;
assign x_1940 = v_2606 | ~v_2282 | ~v_2580;
assign x_1941 = v_2580 | ~v_2282 | ~v_2606;
assign x_1942 = v_2282 | ~v_2580 | ~v_2606;
assign x_1943 = v_2606 | ~v_2283 | ~v_2581;
assign x_1944 = v_2581 | ~v_2283 | ~v_2606;
assign x_1945 = v_2283 | ~v_2581 | ~v_2606;
assign x_1946 = v_2606 | ~v_2284 | ~v_2582;
assign x_1947 = v_2582 | ~v_2284 | ~v_2606;
assign x_1948 = v_2284 | ~v_2582 | ~v_2606;
assign x_1949 = v_2282 | v_2283 | v_2284 | ~v_2579 | ~v_2606;
assign x_1950 = v_2281 | v_2580 | v_2581 | v_2582 | ~v_2606;
assign x_1951 = v_2579 | v_2607 | ~v_584;
assign x_1952 = v_584 | v_2579 | ~v_2607;
assign x_1953 = ~v_584 | ~v_2579 | ~v_2607;
assign x_1954 = v_2607 | ~v_585 | ~v_2580;
assign x_1955 = v_2580 | ~v_585 | ~v_2607;
assign x_1956 = v_585 | ~v_2580 | ~v_2607;
assign x_1957 = v_2607 | ~v_586 | ~v_2581;
assign x_1958 = v_2581 | ~v_586 | ~v_2607;
assign x_1959 = v_586 | ~v_2581 | ~v_2607;
assign x_1960 = v_2607 | ~v_587 | ~v_2582;
assign x_1961 = v_2582 | ~v_587 | ~v_2607;
assign x_1962 = v_587 | ~v_2582 | ~v_2607;
assign x_1963 = v_585 | v_586 | v_587 | ~v_2579 | ~v_2607;
assign x_1964 = v_584 | v_2580 | v_2581 | v_2582 | ~v_2607;
assign x_1965 = v_2429 | v_2616 | ~v_2617;
assign x_1966 = v_2587 | ~v_2429 | ~v_2617;
assign x_1967 = v_2587 | v_2616 | ~v_2617;
assign x_1968 = v_2617 | ~v_2587 | ~v_2616;
assign x_1969 = v_2617 | ~v_2429 | ~v_2587;
assign x_1970 = v_2429 | v_2617 | ~v_2616;
assign x_1971 = v_2579 | v_2638 | ~v_455;
assign x_1972 = v_455 | v_2579 | ~v_2638;
assign x_1973 = ~v_455 | ~v_2579 | ~v_2638;
assign x_1974 = v_2638 | ~v_456 | ~v_2580;
assign x_1975 = v_2580 | ~v_456 | ~v_2638;
assign x_1976 = v_456 | ~v_2580 | ~v_2638;
assign x_1977 = v_2638 | ~v_457 | ~v_2581;
assign x_1978 = v_2581 | ~v_457 | ~v_2638;
assign x_1979 = v_457 | ~v_2581 | ~v_2638;
assign x_1980 = v_2638 | ~v_458 | ~v_2582;
assign x_1981 = v_2582 | ~v_458 | ~v_2638;
assign x_1982 = v_458 | ~v_2582 | ~v_2638;
assign x_1983 = v_456 | v_457 | v_458 | ~v_2579 | ~v_2638;
assign x_1984 = v_455 | v_2580 | v_2581 | v_2582 | ~v_2638;
assign x_1985 = v_2470 | v_2647 | ~v_2648;
assign x_1986 = v_2622 | ~v_2470 | ~v_2648;
assign x_1987 = v_2622 | v_2647 | ~v_2648;
assign x_1988 = v_2648 | ~v_2622 | ~v_2647;
assign x_1989 = v_2648 | ~v_2470 | ~v_2622;
assign x_1990 = v_2470 | v_2648 | ~v_2647;
assign x_1991 = v_2653 | v_2678 | ~v_425;
assign x_1992 = v_425 | v_2653 | ~v_2678;
assign x_1993 = ~v_425 | ~v_2653 | ~v_2678;
assign x_1994 = v_2678 | ~v_426 | ~v_2654;
assign x_1995 = v_2654 | ~v_426 | ~v_2678;
assign x_1996 = v_426 | ~v_2654 | ~v_2678;
assign x_1997 = v_2678 | ~v_427 | ~v_2655;
assign x_1998 = v_2655 | ~v_427 | ~v_2678;
assign x_1999 = v_427 | ~v_2655 | ~v_2678;
assign x_2000 = v_2678 | ~v_428 | ~v_2656;
assign x_2001 = v_2656 | ~v_428 | ~v_2678;
assign x_2002 = v_428 | ~v_2656 | ~v_2678;
assign x_2003 = v_426 | v_427 | v_428 | ~v_2653 | ~v_2678;
assign x_2004 = v_425 | v_2654 | v_2655 | v_2656 | ~v_2678;
assign x_2005 = v_2653 | v_2679 | ~v_495;
assign x_2006 = v_495 | v_2653 | ~v_2679;
assign x_2007 = ~v_495 | ~v_2653 | ~v_2679;
assign x_2008 = v_2679 | ~v_496 | ~v_2654;
assign x_2009 = v_2654 | ~v_496 | ~v_2679;
assign x_2010 = v_496 | ~v_2654 | ~v_2679;
assign x_2011 = v_2679 | ~v_497 | ~v_2655;
assign x_2012 = v_2655 | ~v_497 | ~v_2679;
assign x_2013 = v_497 | ~v_2655 | ~v_2679;
assign x_2014 = v_2679 | ~v_498 | ~v_2656;
assign x_2015 = v_2656 | ~v_498 | ~v_2679;
assign x_2016 = v_498 | ~v_2656 | ~v_2679;
assign x_2017 = v_496 | v_497 | v_498 | ~v_2653 | ~v_2679;
assign x_2018 = v_495 | v_2654 | v_2655 | v_2656 | ~v_2679;
assign x_2019 = v_2653 | v_2680 | ~v_2281;
assign x_2020 = v_2281 | v_2653 | ~v_2680;
assign x_2021 = ~v_2281 | ~v_2653 | ~v_2680;
assign x_2022 = v_2680 | ~v_2282 | ~v_2654;
assign x_2023 = v_2654 | ~v_2282 | ~v_2680;
assign x_2024 = v_2282 | ~v_2654 | ~v_2680;
assign x_2025 = v_2680 | ~v_2283 | ~v_2655;
assign x_2026 = v_2655 | ~v_2283 | ~v_2680;
assign x_2027 = v_2283 | ~v_2655 | ~v_2680;
assign x_2028 = v_2680 | ~v_2284 | ~v_2656;
assign x_2029 = v_2656 | ~v_2284 | ~v_2680;
assign x_2030 = v_2284 | ~v_2656 | ~v_2680;
assign x_2031 = v_2282 | v_2283 | v_2284 | ~v_2653 | ~v_2680;
assign x_2032 = v_2281 | v_2654 | v_2655 | v_2656 | ~v_2680;
assign x_2033 = v_2653 | v_2681 | ~v_584;
assign x_2034 = v_584 | v_2653 | ~v_2681;
assign x_2035 = ~v_584 | ~v_2653 | ~v_2681;
assign x_2036 = v_2681 | ~v_585 | ~v_2654;
assign x_2037 = v_2654 | ~v_585 | ~v_2681;
assign x_2038 = v_585 | ~v_2654 | ~v_2681;
assign x_2039 = v_2681 | ~v_586 | ~v_2655;
assign x_2040 = v_2655 | ~v_586 | ~v_2681;
assign x_2041 = v_586 | ~v_2655 | ~v_2681;
assign x_2042 = v_2681 | ~v_587 | ~v_2656;
assign x_2043 = v_2656 | ~v_587 | ~v_2681;
assign x_2044 = v_587 | ~v_2656 | ~v_2681;
assign x_2045 = v_585 | v_586 | v_587 | ~v_2653 | ~v_2681;
assign x_2046 = v_584 | v_2654 | v_2655 | v_2656 | ~v_2681;
assign x_2047 = v_2429 | v_2690 | ~v_2691;
assign x_2048 = v_2661 | ~v_2429 | ~v_2691;
assign x_2049 = v_2661 | v_2690 | ~v_2691;
assign x_2050 = v_2691 | ~v_2661 | ~v_2690;
assign x_2051 = v_2691 | ~v_2429 | ~v_2661;
assign x_2052 = v_2429 | v_2691 | ~v_2690;
assign x_2053 = v_2653 | v_2712 | ~v_455;
assign x_2054 = v_455 | v_2653 | ~v_2712;
assign x_2055 = ~v_455 | ~v_2653 | ~v_2712;
assign x_2056 = v_2712 | ~v_456 | ~v_2654;
assign x_2057 = v_2654 | ~v_456 | ~v_2712;
assign x_2058 = v_456 | ~v_2654 | ~v_2712;
assign x_2059 = v_2712 | ~v_457 | ~v_2655;
assign x_2060 = v_2655 | ~v_457 | ~v_2712;
assign x_2061 = v_457 | ~v_2655 | ~v_2712;
assign x_2062 = v_2712 | ~v_458 | ~v_2656;
assign x_2063 = v_2656 | ~v_458 | ~v_2712;
assign x_2064 = v_458 | ~v_2656 | ~v_2712;
assign x_2065 = v_456 | v_457 | v_458 | ~v_2653 | ~v_2712;
assign x_2066 = v_455 | v_2654 | v_2655 | v_2656 | ~v_2712;
assign x_2067 = v_2470 | v_2721 | ~v_2722;
assign x_2068 = v_2696 | ~v_2470 | ~v_2722;
assign x_2069 = v_2696 | v_2721 | ~v_2722;
assign x_2070 = v_2722 | ~v_2696 | ~v_2721;
assign x_2071 = v_2722 | ~v_2470 | ~v_2696;
assign x_2072 = v_2470 | v_2722 | ~v_2721;
assign x_2073 = v_2727 | v_2752 | ~v_425;
assign x_2074 = v_425 | v_2727 | ~v_2752;
assign x_2075 = ~v_425 | ~v_2727 | ~v_2752;
assign x_2076 = v_2752 | ~v_426 | ~v_2728;
assign x_2077 = v_2728 | ~v_426 | ~v_2752;
assign x_2078 = v_426 | ~v_2728 | ~v_2752;
assign x_2079 = v_2752 | ~v_427 | ~v_2729;
assign x_2080 = v_2729 | ~v_427 | ~v_2752;
assign x_2081 = v_427 | ~v_2729 | ~v_2752;
assign x_2082 = v_2752 | ~v_428 | ~v_2730;
assign x_2083 = v_2730 | ~v_428 | ~v_2752;
assign x_2084 = v_428 | ~v_2730 | ~v_2752;
assign x_2085 = v_426 | v_427 | v_428 | ~v_2727 | ~v_2752;
assign x_2086 = v_425 | v_2728 | v_2729 | v_2730 | ~v_2752;
assign x_2087 = v_2727 | v_2753 | ~v_495;
assign x_2088 = v_495 | v_2727 | ~v_2753;
assign x_2089 = ~v_495 | ~v_2727 | ~v_2753;
assign x_2090 = v_2753 | ~v_496 | ~v_2728;
assign x_2091 = v_2728 | ~v_496 | ~v_2753;
assign x_2092 = v_496 | ~v_2728 | ~v_2753;
assign x_2093 = v_2753 | ~v_497 | ~v_2729;
assign x_2094 = v_2729 | ~v_497 | ~v_2753;
assign x_2095 = v_497 | ~v_2729 | ~v_2753;
assign x_2096 = v_2753 | ~v_498 | ~v_2730;
assign x_2097 = v_2730 | ~v_498 | ~v_2753;
assign x_2098 = v_498 | ~v_2730 | ~v_2753;
assign x_2099 = v_496 | v_497 | v_498 | ~v_2727 | ~v_2753;
assign x_2100 = v_495 | v_2728 | v_2729 | v_2730 | ~v_2753;
assign x_2101 = v_2727 | v_2754 | ~v_2281;
assign x_2102 = v_2281 | v_2727 | ~v_2754;
assign x_2103 = ~v_2281 | ~v_2727 | ~v_2754;
assign x_2104 = v_2754 | ~v_2282 | ~v_2728;
assign x_2105 = v_2728 | ~v_2282 | ~v_2754;
assign x_2106 = v_2282 | ~v_2728 | ~v_2754;
assign x_2107 = v_2754 | ~v_2283 | ~v_2729;
assign x_2108 = v_2729 | ~v_2283 | ~v_2754;
assign x_2109 = v_2283 | ~v_2729 | ~v_2754;
assign x_2110 = v_2754 | ~v_2284 | ~v_2730;
assign x_2111 = v_2730 | ~v_2284 | ~v_2754;
assign x_2112 = v_2284 | ~v_2730 | ~v_2754;
assign x_2113 = v_2282 | v_2283 | v_2284 | ~v_2727 | ~v_2754;
assign x_2114 = v_2281 | v_2728 | v_2729 | v_2730 | ~v_2754;
assign x_2115 = v_2727 | v_2755 | ~v_584;
assign x_2116 = v_584 | v_2727 | ~v_2755;
assign x_2117 = ~v_584 | ~v_2727 | ~v_2755;
assign x_2118 = v_2755 | ~v_585 | ~v_2728;
assign x_2119 = v_2728 | ~v_585 | ~v_2755;
assign x_2120 = v_585 | ~v_2728 | ~v_2755;
assign x_2121 = v_2755 | ~v_586 | ~v_2729;
assign x_2122 = v_2729 | ~v_586 | ~v_2755;
assign x_2123 = v_586 | ~v_2729 | ~v_2755;
assign x_2124 = v_2755 | ~v_587 | ~v_2730;
assign x_2125 = v_2730 | ~v_587 | ~v_2755;
assign x_2126 = v_587 | ~v_2730 | ~v_2755;
assign x_2127 = v_585 | v_586 | v_587 | ~v_2727 | ~v_2755;
assign x_2128 = v_584 | v_2728 | v_2729 | v_2730 | ~v_2755;
assign x_2129 = v_2429 | v_2764 | ~v_2765;
assign x_2130 = v_2735 | ~v_2429 | ~v_2765;
assign x_2131 = v_2735 | v_2764 | ~v_2765;
assign x_2132 = v_2765 | ~v_2735 | ~v_2764;
assign x_2133 = v_2765 | ~v_2429 | ~v_2735;
assign x_2134 = v_2429 | v_2765 | ~v_2764;
assign x_2135 = v_2727 | v_2786 | ~v_455;
assign x_2136 = v_455 | v_2727 | ~v_2786;
assign x_2137 = ~v_455 | ~v_2727 | ~v_2786;
assign x_2138 = v_2786 | ~v_456 | ~v_2728;
assign x_2139 = v_2728 | ~v_456 | ~v_2786;
assign x_2140 = v_456 | ~v_2728 | ~v_2786;
assign x_2141 = v_2786 | ~v_457 | ~v_2729;
assign x_2142 = v_2729 | ~v_457 | ~v_2786;
assign x_2143 = v_457 | ~v_2729 | ~v_2786;
assign x_2144 = v_2786 | ~v_458 | ~v_2730;
assign x_2145 = v_2730 | ~v_458 | ~v_2786;
assign x_2146 = v_458 | ~v_2730 | ~v_2786;
assign x_2147 = v_456 | v_457 | v_458 | ~v_2727 | ~v_2786;
assign x_2148 = v_455 | v_2728 | v_2729 | v_2730 | ~v_2786;
assign x_2149 = v_2470 | v_2795 | ~v_2796;
assign x_2150 = v_2770 | ~v_2470 | ~v_2796;
assign x_2151 = v_2770 | v_2795 | ~v_2796;
assign x_2152 = v_2796 | ~v_2770 | ~v_2795;
assign x_2153 = v_2796 | ~v_2470 | ~v_2770;
assign x_2154 = v_2470 | v_2796 | ~v_2795;
assign x_2155 = ~v_2800 | ~v_2801;
assign x_2156 = ~v_2800 | ~v_2802;
assign x_2157 = ~v_2801 | ~v_2802;
assign x_2158 = v_2800 | ~v_2651 | ~v_2804;
assign x_2159 = v_2651 | v_2801 | ~v_2804;
assign x_2160 = v_2800 | v_2801 | ~v_2804;
assign x_2161 = v_2804 | ~v_2800 | ~v_2801;
assign x_2162 = v_2651 | v_2804 | ~v_2801;
assign x_2163 = v_2804 | ~v_2651 | ~v_2800;
assign x_2164 = v_2801 | ~v_2651 | ~v_2805;
assign x_2165 = v_2651 | v_2802 | ~v_2805;
assign x_2166 = v_2801 | v_2802 | ~v_2805;
assign x_2167 = v_2805 | ~v_2801 | ~v_2802;
assign x_2168 = v_2651 | v_2805 | ~v_2802;
assign x_2169 = v_2805 | ~v_2651 | ~v_2801;
assign x_2170 = ~v_2803 | ~v_2804;
assign x_2171 = ~v_2803 | ~v_2805;
assign x_2172 = ~v_2803 | ~v_2806;
assign x_2173 = ~v_2804 | ~v_2805;
assign x_2174 = ~v_2804 | ~v_2806;
assign x_2175 = ~v_2805 | ~v_2806;
assign x_2176 = v_2803 | ~v_2577 | ~v_2808;
assign x_2177 = v_2577 | v_2804 | ~v_2808;
assign x_2178 = v_2803 | v_2804 | ~v_2808;
assign x_2179 = v_2808 | ~v_2803 | ~v_2804;
assign x_2180 = v_2577 | v_2808 | ~v_2804;
assign x_2181 = v_2808 | ~v_2577 | ~v_2803;
assign x_2182 = v_2804 | ~v_2577 | ~v_2809;
assign x_2183 = v_2577 | v_2805 | ~v_2809;
assign x_2184 = v_2804 | v_2805 | ~v_2809;
assign x_2185 = v_2809 | ~v_2804 | ~v_2805;
assign x_2186 = v_2577 | v_2809 | ~v_2805;
assign x_2187 = v_2809 | ~v_2577 | ~v_2804;
assign x_2188 = v_2805 | ~v_2577 | ~v_2810;
assign x_2189 = v_2577 | v_2806 | ~v_2810;
assign x_2190 = v_2805 | v_2806 | ~v_2810;
assign x_2191 = v_2810 | ~v_2805 | ~v_2806;
assign x_2192 = v_2577 | v_2810 | ~v_2806;
assign x_2193 = v_2810 | ~v_2577 | ~v_2805;
assign x_2194 = ~v_2807 | ~v_2808;
assign x_2195 = ~v_2807 | ~v_2809;
assign x_2196 = ~v_2807 | ~v_2810;
assign x_2197 = ~v_2807 | ~v_2811;
assign x_2198 = ~v_2808 | ~v_2809;
assign x_2199 = ~v_2808 | ~v_2810;
assign x_2200 = ~v_2808 | ~v_2811;
assign x_2201 = ~v_2809 | ~v_2810;
assign x_2202 = ~v_2809 | ~v_2811;
assign x_2203 = ~v_2810 | ~v_2811;
assign x_2204 = v_2812 | ~v_1744 | ~v_2807;
assign x_2205 = v_2807 | ~v_1744 | ~v_2812;
assign x_2206 = v_1744 | ~v_2807 | ~v_2812;
assign x_2207 = v_2812 | ~v_1745 | ~v_2808;
assign x_2208 = v_2808 | ~v_1745 | ~v_2812;
assign x_2209 = v_1745 | ~v_2808 | ~v_2812;
assign x_2210 = v_2812 | ~v_1746 | ~v_2809;
assign x_2211 = v_2809 | ~v_1746 | ~v_2812;
assign x_2212 = v_1746 | ~v_2809 | ~v_2812;
assign x_2213 = v_2812 | ~v_1747 | ~v_2810;
assign x_2214 = v_2810 | ~v_1747 | ~v_2812;
assign x_2215 = v_1747 | ~v_2810 | ~v_2812;
assign x_2216 = v_2812 | ~v_1748 | ~v_2811;
assign x_2217 = v_2811 | ~v_1748 | ~v_2812;
assign x_2218 = v_1748 | ~v_2811 | ~v_2812;
assign x_2219 = v_1744 | v_1745 | v_1746 | v_1747 | v_1748 | ~v_2812;
assign x_2220 = v_2807 | v_2808 | v_2809 | v_2810 | v_2811 | ~v_2812;
assign x_2221 = v_2336 | v_2799 | ~v_2816;
assign x_2222 = ~v_2799 | ~v_2815 | ~v_2816;
assign x_2223 = v_2336 | ~v_2815 | ~v_2816;
assign x_2224 = v_2815 | v_2816 | ~v_2336;
assign x_2225 = v_2815 | v_2816 | ~v_2799;
assign x_2226 = v_2799 | v_2816 | ~v_2336;
assign x_2227 = v_2816 | ~v_2725 | ~v_2819;
assign x_2228 = v_2725 | ~v_2815 | ~v_2819;
assign x_2229 = v_2816 | ~v_2815 | ~v_2819;
assign x_2230 = v_2815 | v_2819 | ~v_2816;
assign x_2231 = v_2725 | v_2815 | v_2819;
assign x_2232 = v_2819 | ~v_2725 | ~v_2816;
assign x_2233 = v_2817 | ~v_2725 | ~v_2820;
assign x_2234 = v_2725 | v_2815 | ~v_2820;
assign x_2235 = v_2815 | v_2817 | ~v_2820;
assign x_2236 = v_2820 | ~v_2815 | ~v_2817;
assign x_2237 = v_2725 | v_2820 | ~v_2815;
assign x_2238 = v_2820 | ~v_2725 | ~v_2817;
assign x_2239 = v_2366 | ~v_2800 | ~v_2822;
assign x_2240 = v_2800 | v_2819 | ~v_2822;
assign x_2241 = v_2366 | v_2819 | ~v_2822;
assign x_2242 = v_2822 | ~v_2366 | ~v_2819;
assign x_2243 = v_2800 | v_2822 | ~v_2819;
assign x_2244 = v_2822 | ~v_2366 | ~v_2800;
assign x_2245 = v_2822 | ~v_2651 | ~v_2826;
assign x_2246 = v_2651 | v_2819 | ~v_2826;
assign x_2247 = v_2819 | v_2822 | ~v_2826;
assign x_2248 = v_2826 | ~v_2819 | ~v_2822;
assign x_2249 = v_2651 | v_2826 | ~v_2819;
assign x_2250 = v_2826 | ~v_2651 | ~v_2822;
assign x_2251 = v_2823 | ~v_2651 | ~v_2827;
assign x_2252 = v_2651 | v_2820 | ~v_2827;
assign x_2253 = v_2820 | v_2823 | ~v_2827;
assign x_2254 = v_2827 | ~v_2820 | ~v_2823;
assign x_2255 = v_2651 | v_2827 | ~v_2820;
assign x_2256 = v_2827 | ~v_2651 | ~v_2823;
assign x_2257 = v_2824 | ~v_2651 | ~v_2828;
assign x_2258 = v_2651 | v_2821 | ~v_2828;
assign x_2259 = v_2821 | v_2824 | ~v_2828;
assign x_2260 = v_2828 | ~v_2821 | ~v_2824;
assign x_2261 = v_2651 | v_2828 | ~v_2821;
assign x_2262 = v_2828 | ~v_2651 | ~v_2824;
assign x_2263 = v_2398 | ~v_2803 | ~v_2830;
assign x_2264 = v_2803 | v_2826 | ~v_2830;
assign x_2265 = v_2398 | v_2826 | ~v_2830;
assign x_2266 = v_2830 | ~v_2398 | ~v_2826;
assign x_2267 = v_2803 | v_2830 | ~v_2826;
assign x_2268 = v_2830 | ~v_2398 | ~v_2803;
assign x_2269 = v_2830 | ~v_2577 | ~v_2835;
assign x_2270 = v_2577 | v_2826 | ~v_2835;
assign x_2271 = v_2826 | v_2830 | ~v_2835;
assign x_2272 = v_2835 | ~v_2826 | ~v_2830;
assign x_2273 = v_2577 | v_2835 | ~v_2826;
assign x_2274 = v_2835 | ~v_2577 | ~v_2830;
assign x_2275 = v_2831 | ~v_2577 | ~v_2836;
assign x_2276 = v_2577 | v_2827 | ~v_2836;
assign x_2277 = v_2827 | v_2831 | ~v_2836;
assign x_2278 = v_2836 | ~v_2827 | ~v_2831;
assign x_2279 = v_2577 | v_2836 | ~v_2827;
assign x_2280 = v_2836 | ~v_2577 | ~v_2831;
assign x_2281 = v_2832 | ~v_2577 | ~v_2837;
assign x_2282 = v_2577 | v_2828 | ~v_2837;
assign x_2283 = v_2828 | v_2832 | ~v_2837;
assign x_2284 = v_2837 | ~v_2828 | ~v_2832;
assign x_2285 = v_2577 | v_2837 | ~v_2828;
assign x_2286 = v_2837 | ~v_2577 | ~v_2832;
assign x_2287 = v_2833 | ~v_2577 | ~v_2838;
assign x_2288 = v_2577 | v_2829 | ~v_2838;
assign x_2289 = v_2829 | v_2833 | ~v_2838;
assign x_2290 = v_2838 | ~v_2829 | ~v_2833;
assign x_2291 = v_2577 | v_2838 | ~v_2829;
assign x_2292 = v_2838 | ~v_2577 | ~v_2833;
assign x_2293 = v_2868 | v_2875 | ~v_659;
assign x_2294 = v_659 | v_2868 | ~v_2875;
assign x_2295 = ~v_659 | ~v_2868 | ~v_2875;
assign x_2296 = v_2870 | v_2875 | ~v_660;
assign x_2297 = v_660 | v_2870 | ~v_2875;
assign x_2298 = ~v_660 | ~v_2870 | ~v_2875;
assign x_2299 = v_2872 | v_2875 | ~v_661;
assign x_2300 = v_661 | v_2872 | ~v_2875;
assign x_2301 = ~v_661 | ~v_2872 | ~v_2875;
assign x_2302 = v_2874 | v_2875 | ~v_662;
assign x_2303 = v_662 | v_2874 | ~v_2875;
assign x_2304 = ~v_662 | ~v_2874 | ~v_2875;
assign x_2305 = ~v_2868 | ~v_2870 | ~v_2872 | ~v_2874 | ~v_2875;
assign x_2306 = v_659 | v_660 | v_661 | v_662 | ~v_2875;
assign x_2307 = v_1744 | ~v_2876 | ~v_2877;
assign x_2308 = ~v_1744 | ~v_2812 | ~v_2877;
assign x_2309 = ~v_2812 | ~v_2876 | ~v_2877;
assign x_2310 = v_2812 | v_2876 | v_2877;
assign x_2311 = v_2812 | v_2877 | ~v_1744;
assign x_2312 = v_1744 | v_2876 | v_2877;
assign x_2313 = v_2366 | ~v_2801 | ~v_2882;
assign x_2314 = v_2801 | ~v_2881 | ~v_2882;
assign x_2315 = v_2366 | ~v_2881 | ~v_2882;
assign x_2316 = v_2881 | v_2882 | ~v_2366;
assign x_2317 = v_2801 | v_2881 | v_2882;
assign x_2318 = v_2882 | ~v_2366 | ~v_2801;
assign x_2319 = v_2882 | ~v_2651 | ~v_2885;
assign x_2320 = v_2651 | ~v_2881 | ~v_2885;
assign x_2321 = v_2882 | ~v_2881 | ~v_2885;
assign x_2322 = v_2881 | v_2885 | ~v_2882;
assign x_2323 = v_2651 | v_2881 | v_2885;
assign x_2324 = v_2885 | ~v_2651 | ~v_2882;
assign x_2325 = v_2883 | ~v_2651 | ~v_2886;
assign x_2326 = v_2651 | v_2881 | ~v_2886;
assign x_2327 = v_2881 | v_2883 | ~v_2886;
assign x_2328 = v_2886 | ~v_2881 | ~v_2883;
assign x_2329 = v_2651 | v_2886 | ~v_2881;
assign x_2330 = v_2886 | ~v_2651 | ~v_2883;
assign x_2331 = v_2398 | ~v_2804 | ~v_2888;
assign x_2332 = v_2804 | v_2885 | ~v_2888;
assign x_2333 = v_2398 | v_2885 | ~v_2888;
assign x_2334 = v_2888 | ~v_2398 | ~v_2885;
assign x_2335 = v_2804 | v_2888 | ~v_2885;
assign x_2336 = v_2888 | ~v_2398 | ~v_2804;
assign x_2337 = v_2888 | ~v_2577 | ~v_2892;
assign x_2338 = v_2577 | v_2885 | ~v_2892;
assign x_2339 = v_2885 | v_2888 | ~v_2892;
assign x_2340 = v_2892 | ~v_2885 | ~v_2888;
assign x_2341 = v_2577 | v_2892 | ~v_2885;
assign x_2342 = v_2892 | ~v_2577 | ~v_2888;
assign x_2343 = v_2889 | ~v_2577 | ~v_2893;
assign x_2344 = v_2577 | v_2886 | ~v_2893;
assign x_2345 = v_2886 | v_2889 | ~v_2893;
assign x_2346 = v_2893 | ~v_2886 | ~v_2889;
assign x_2347 = v_2577 | v_2893 | ~v_2886;
assign x_2348 = v_2893 | ~v_2577 | ~v_2889;
assign x_2349 = v_2890 | ~v_2577 | ~v_2894;
assign x_2350 = v_2577 | v_2887 | ~v_2894;
assign x_2351 = v_2887 | v_2890 | ~v_2894;
assign x_2352 = v_2894 | ~v_2887 | ~v_2890;
assign x_2353 = v_2577 | v_2894 | ~v_2887;
assign x_2354 = v_2894 | ~v_2577 | ~v_2890;
assign x_2355 = v_2915 | v_2922 | ~v_663;
assign x_2356 = v_663 | v_2915 | ~v_2922;
assign x_2357 = ~v_663 | ~v_2915 | ~v_2922;
assign x_2358 = v_2917 | v_2922 | ~v_664;
assign x_2359 = v_664 | v_2917 | ~v_2922;
assign x_2360 = ~v_664 | ~v_2917 | ~v_2922;
assign x_2361 = v_2919 | v_2922 | ~v_665;
assign x_2362 = v_665 | v_2919 | ~v_2922;
assign x_2363 = ~v_665 | ~v_2919 | ~v_2922;
assign x_2364 = v_2921 | v_2922 | ~v_666;
assign x_2365 = v_666 | v_2921 | ~v_2922;
assign x_2366 = ~v_666 | ~v_2921 | ~v_2922;
assign x_2367 = ~v_2915 | ~v_2917 | ~v_2919 | ~v_2921 | ~v_2922;
assign x_2368 = v_663 | v_664 | v_665 | v_666 | ~v_2922;
assign x_2369 = ~v_2172 | ~v_2923 | ~v_2924;
assign x_2370 = v_2172 | v_2877 | ~v_2924;
assign x_2371 = v_2877 | ~v_2923 | ~v_2924;
assign x_2372 = v_2923 | v_2924 | ~v_2877;
assign x_2373 = v_2172 | v_2924 | ~v_2877;
assign x_2374 = v_2923 | v_2924 | ~v_2172;
assign x_2375 = v_2398 | ~v_2805 | ~v_2929;
assign x_2376 = v_2805 | ~v_2928 | ~v_2929;
assign x_2377 = v_2398 | ~v_2928 | ~v_2929;
assign x_2378 = v_2928 | v_2929 | ~v_2398;
assign x_2379 = v_2805 | v_2928 | v_2929;
assign x_2380 = v_2929 | ~v_2398 | ~v_2805;
assign x_2381 = v_2929 | ~v_2577 | ~v_2932;
assign x_2382 = v_2577 | ~v_2928 | ~v_2932;
assign x_2383 = v_2929 | ~v_2928 | ~v_2932;
assign x_2384 = v_2928 | v_2932 | ~v_2929;
assign x_2385 = v_2577 | v_2928 | v_2932;
assign x_2386 = v_2932 | ~v_2577 | ~v_2929;
assign x_2387 = v_2930 | ~v_2577 | ~v_2933;
assign x_2388 = v_2577 | v_2928 | ~v_2933;
assign x_2389 = v_2928 | v_2930 | ~v_2933;
assign x_2390 = v_2933 | ~v_2928 | ~v_2930;
assign x_2391 = v_2577 | v_2933 | ~v_2928;
assign x_2392 = v_2933 | ~v_2577 | ~v_2930;
assign x_2393 = v_2945 | v_2952 | ~v_667;
assign x_2394 = v_667 | v_2945 | ~v_2952;
assign x_2395 = ~v_667 | ~v_2945 | ~v_2952;
assign x_2396 = v_2947 | v_2952 | ~v_668;
assign x_2397 = v_668 | v_2947 | ~v_2952;
assign x_2398 = ~v_668 | ~v_2947 | ~v_2952;
assign x_2399 = v_2949 | v_2952 | ~v_669;
assign x_2400 = v_669 | v_2949 | ~v_2952;
assign x_2401 = ~v_669 | ~v_2949 | ~v_2952;
assign x_2402 = v_2951 | v_2952 | ~v_670;
assign x_2403 = v_670 | v_2951 | ~v_2952;
assign x_2404 = ~v_670 | ~v_2951 | ~v_2952;
assign x_2405 = ~v_2945 | ~v_2947 | ~v_2949 | ~v_2951 | ~v_2952;
assign x_2406 = v_667 | v_668 | v_669 | v_670 | ~v_2952;
assign x_2407 = ~v_2220 | ~v_2953 | ~v_2954;
assign x_2408 = v_2220 | v_2924 | ~v_2954;
assign x_2409 = v_2924 | ~v_2953 | ~v_2954;
assign x_2410 = v_2953 | v_2954 | ~v_2924;
assign x_2411 = v_2220 | v_2954 | ~v_2924;
assign x_2412 = v_2953 | v_2954 | ~v_2220;
assign x_2413 = v_2963 | v_2967 | ~v_671;
assign x_2414 = v_671 | v_2963 | ~v_2967;
assign x_2415 = ~v_671 | ~v_2963 | ~v_2967;
assign x_2416 = v_2967 | ~v_672 | ~v_2964;
assign x_2417 = v_2964 | ~v_672 | ~v_2967;
assign x_2418 = v_672 | ~v_2964 | ~v_2967;
assign x_2419 = v_2967 | ~v_673 | ~v_2965;
assign x_2420 = v_2965 | ~v_673 | ~v_2967;
assign x_2421 = v_673 | ~v_2965 | ~v_2967;
assign x_2422 = v_2967 | ~v_674 | ~v_2966;
assign x_2423 = v_2966 | ~v_674 | ~v_2967;
assign x_2424 = v_674 | ~v_2966 | ~v_2967;
assign x_2425 = v_672 | v_673 | v_674 | ~v_2963 | ~v_2967;
assign x_2426 = v_671 | v_2964 | v_2965 | v_2966 | ~v_2967;
assign x_2427 = ~v_1748 | ~v_2968 | ~v_2969;
assign x_2428 = v_1748 | v_2954 | ~v_2969;
assign x_2429 = v_2954 | ~v_2968 | ~v_2969;
assign x_2430 = v_2968 | v_2969 | ~v_2954;
assign x_2431 = v_1748 | v_2969 | ~v_2954;
assign x_2432 = v_2968 | v_2969 | ~v_1748;
assign x_2433 = v_509 | v_2987 | ~v_2988;
assign x_2434 = v_487 | ~v_509 | ~v_2988;
assign x_2435 = v_487 | v_2987 | ~v_2988;
assign x_2436 = v_2988 | ~v_487 | ~v_2987;
assign x_2437 = v_2988 | ~v_487 | ~v_509;
assign x_2438 = v_509 | v_2988 | ~v_2987;
assign x_2439 = v_2993 | ~v_2994;
assign x_2440 = v_2993 | ~v_2995;
assign x_2441 = v_2993 | ~v_2996;
assign x_2442 = ~v_2994 | ~v_2995;
assign x_2443 = ~v_2994 | ~v_2996;
assign x_2444 = ~v_2995 | ~v_2996;
assign x_2445 = v_2996 | ~v_3012 | ~v_3013;
assign x_2446 = ~v_2996 | ~v_3011 | ~v_3013;
assign x_2447 = ~v_3011 | ~v_3012 | ~v_3013;
assign x_2448 = v_3011 | v_3012 | v_3013;
assign x_2449 = v_3011 | v_3013 | ~v_2996;
assign x_2450 = v_2996 | v_3012 | v_3013;
assign x_2451 = v_2996 | ~v_3027 | ~v_3028;
assign x_2452 = ~v_2996 | ~v_3026 | ~v_3028;
assign x_2453 = ~v_3026 | ~v_3027 | ~v_3028;
assign x_2454 = v_3026 | v_3027 | v_3028;
assign x_2455 = v_3026 | v_3028 | ~v_2996;
assign x_2456 = v_2996 | v_3027 | v_3028;
assign x_2457 = v_2998 | ~v_3029 | ~v_3030;
assign x_2458 = v_3028 | ~v_2998 | ~v_3030;
assign x_2459 = v_3028 | ~v_3029 | ~v_3030;
assign x_2460 = v_3029 | v_3030 | ~v_3028;
assign x_2461 = v_3030 | ~v_2998 | ~v_3028;
assign x_2462 = v_2998 | v_3029 | v_3030;
assign x_2463 = v_583 | v_3043 | ~v_3044;
assign x_2464 = v_593 | ~v_583 | ~v_3044;
assign x_2465 = v_593 | v_3043 | ~v_3044;
assign x_2466 = v_3044 | ~v_593 | ~v_3043;
assign x_2467 = v_3044 | ~v_583 | ~v_593;
assign x_2468 = v_583 | v_3044 | ~v_3043;
assign x_2469 = v_626 | v_3046 | ~v_3047;
assign x_2470 = v_632 | ~v_626 | ~v_3047;
assign x_2471 = v_632 | v_3046 | ~v_3047;
assign x_2472 = v_3047 | ~v_632 | ~v_3046;
assign x_2473 = v_3047 | ~v_626 | ~v_632;
assign x_2474 = v_626 | v_3047 | ~v_3046;
assign x_2475 = v_583 | v_3049 | ~v_3050;
assign x_2476 = v_205 | ~v_583 | ~v_3050;
assign x_2477 = v_205 | v_3049 | ~v_3050;
assign x_2478 = v_3050 | ~v_205 | ~v_3049;
assign x_2479 = v_3050 | ~v_205 | ~v_583;
assign x_2480 = v_583 | v_3050 | ~v_3049;
assign x_2481 = v_626 | v_3051 | ~v_3052;
assign x_2482 = v_235 | ~v_626 | ~v_3052;
assign x_2483 = v_235 | v_3051 | ~v_3052;
assign x_2484 = v_3052 | ~v_235 | ~v_3051;
assign x_2485 = v_3052 | ~v_235 | ~v_626;
assign x_2486 = v_626 | v_3052 | ~v_3051;
assign x_2487 = v_3055 | v_3080 | ~v_229;
assign x_2488 = v_229 | v_3055 | ~v_3080;
assign x_2489 = ~v_229 | ~v_3055 | ~v_3080;
assign x_2490 = v_3080 | ~v_230 | ~v_3056;
assign x_2491 = v_3056 | ~v_230 | ~v_3080;
assign x_2492 = v_230 | ~v_3056 | ~v_3080;
assign x_2493 = v_3080 | ~v_231 | ~v_3057;
assign x_2494 = v_3057 | ~v_231 | ~v_3080;
assign x_2495 = v_231 | ~v_3057 | ~v_3080;
assign x_2496 = v_3080 | ~v_232 | ~v_3058;
assign x_2497 = v_3058 | ~v_232 | ~v_3080;
assign x_2498 = v_232 | ~v_3058 | ~v_3080;
assign x_2499 = v_230 | v_231 | v_232 | ~v_3055 | ~v_3080;
assign x_2500 = v_229 | v_3056 | v_3057 | v_3058 | ~v_3080;
assign x_2501 = v_583 | v_3087 | ~v_3088;
assign x_2502 = v_3063 | ~v_583 | ~v_3088;
assign x_2503 = v_3063 | v_3087 | ~v_3088;
assign x_2504 = v_3088 | ~v_3063 | ~v_3087;
assign x_2505 = v_3088 | ~v_583 | ~v_3063;
assign x_2506 = v_583 | v_3088 | ~v_3087;
assign x_2507 = v_3055 | v_3109 | ~v_259;
assign x_2508 = v_259 | v_3055 | ~v_3109;
assign x_2509 = ~v_259 | ~v_3055 | ~v_3109;
assign x_2510 = v_3109 | ~v_260 | ~v_3056;
assign x_2511 = v_3056 | ~v_260 | ~v_3109;
assign x_2512 = v_260 | ~v_3056 | ~v_3109;
assign x_2513 = v_3109 | ~v_261 | ~v_3057;
assign x_2514 = v_3057 | ~v_261 | ~v_3109;
assign x_2515 = v_261 | ~v_3057 | ~v_3109;
assign x_2516 = v_3109 | ~v_262 | ~v_3058;
assign x_2517 = v_3058 | ~v_262 | ~v_3109;
assign x_2518 = v_262 | ~v_3058 | ~v_3109;
assign x_2519 = v_260 | v_261 | v_262 | ~v_3055 | ~v_3109;
assign x_2520 = v_259 | v_3056 | v_3057 | v_3058 | ~v_3109;
assign x_2521 = v_626 | v_3116 | ~v_3117;
assign x_2522 = v_3093 | ~v_626 | ~v_3117;
assign x_2523 = v_3093 | v_3116 | ~v_3117;
assign x_2524 = v_3117 | ~v_3093 | ~v_3116;
assign x_2525 = v_3117 | ~v_626 | ~v_3093;
assign x_2526 = v_626 | v_3117 | ~v_3116;
assign x_2527 = v_3122 | v_3147 | ~v_229;
assign x_2528 = v_229 | v_3122 | ~v_3147;
assign x_2529 = ~v_229 | ~v_3122 | ~v_3147;
assign x_2530 = v_3147 | ~v_230 | ~v_3123;
assign x_2531 = v_3123 | ~v_230 | ~v_3147;
assign x_2532 = v_230 | ~v_3123 | ~v_3147;
assign x_2533 = v_3147 | ~v_231 | ~v_3124;
assign x_2534 = v_3124 | ~v_231 | ~v_3147;
assign x_2535 = v_231 | ~v_3124 | ~v_3147;
assign x_2536 = v_3147 | ~v_232 | ~v_3125;
assign x_2537 = v_3125 | ~v_232 | ~v_3147;
assign x_2538 = v_232 | ~v_3125 | ~v_3147;
assign x_2539 = v_230 | v_231 | v_232 | ~v_3122 | ~v_3147;
assign x_2540 = v_229 | v_3123 | v_3124 | v_3125 | ~v_3147;
assign x_2541 = v_583 | v_3154 | ~v_3155;
assign x_2542 = v_3130 | ~v_583 | ~v_3155;
assign x_2543 = v_3130 | v_3154 | ~v_3155;
assign x_2544 = v_3155 | ~v_3130 | ~v_3154;
assign x_2545 = v_3155 | ~v_583 | ~v_3130;
assign x_2546 = v_583 | v_3155 | ~v_3154;
assign x_2547 = v_3122 | v_3176 | ~v_259;
assign x_2548 = v_259 | v_3122 | ~v_3176;
assign x_2549 = ~v_259 | ~v_3122 | ~v_3176;
assign x_2550 = v_3176 | ~v_260 | ~v_3123;
assign x_2551 = v_3123 | ~v_260 | ~v_3176;
assign x_2552 = v_260 | ~v_3123 | ~v_3176;
assign x_2553 = v_3176 | ~v_261 | ~v_3124;
assign x_2554 = v_3124 | ~v_261 | ~v_3176;
assign x_2555 = v_261 | ~v_3124 | ~v_3176;
assign x_2556 = v_3176 | ~v_262 | ~v_3125;
assign x_2557 = v_3125 | ~v_262 | ~v_3176;
assign x_2558 = v_262 | ~v_3125 | ~v_3176;
assign x_2559 = v_260 | v_261 | v_262 | ~v_3122 | ~v_3176;
assign x_2560 = v_259 | v_3123 | v_3124 | v_3125 | ~v_3176;
assign x_2561 = v_626 | v_3183 | ~v_3184;
assign x_2562 = v_3160 | ~v_626 | ~v_3184;
assign x_2563 = v_3160 | v_3183 | ~v_3184;
assign x_2564 = v_3184 | ~v_3160 | ~v_3183;
assign x_2565 = v_3184 | ~v_626 | ~v_3160;
assign x_2566 = v_626 | v_3184 | ~v_3183;
assign x_2567 = v_3189 | v_3214 | ~v_229;
assign x_2568 = v_229 | v_3189 | ~v_3214;
assign x_2569 = ~v_229 | ~v_3189 | ~v_3214;
assign x_2570 = v_3214 | ~v_230 | ~v_3190;
assign x_2571 = v_3190 | ~v_230 | ~v_3214;
assign x_2572 = v_230 | ~v_3190 | ~v_3214;
assign x_2573 = v_3214 | ~v_231 | ~v_3191;
assign x_2574 = v_3191 | ~v_231 | ~v_3214;
assign x_2575 = v_231 | ~v_3191 | ~v_3214;
assign x_2576 = v_3214 | ~v_232 | ~v_3192;
assign x_2577 = v_3192 | ~v_232 | ~v_3214;
assign x_2578 = v_232 | ~v_3192 | ~v_3214;
assign x_2579 = v_230 | v_231 | v_232 | ~v_3189 | ~v_3214;
assign x_2580 = v_229 | v_3190 | v_3191 | v_3192 | ~v_3214;
assign x_2581 = v_583 | v_3221 | ~v_3222;
assign x_2582 = v_3197 | ~v_583 | ~v_3222;
assign x_2583 = v_3197 | v_3221 | ~v_3222;
assign x_2584 = v_3222 | ~v_3197 | ~v_3221;
assign x_2585 = v_3222 | ~v_583 | ~v_3197;
assign x_2586 = v_583 | v_3222 | ~v_3221;
assign x_2587 = v_3189 | v_3243 | ~v_259;
assign x_2588 = v_259 | v_3189 | ~v_3243;
assign x_2589 = ~v_259 | ~v_3189 | ~v_3243;
assign x_2590 = v_3243 | ~v_260 | ~v_3190;
assign x_2591 = v_3190 | ~v_260 | ~v_3243;
assign x_2592 = v_260 | ~v_3190 | ~v_3243;
assign x_2593 = v_3243 | ~v_261 | ~v_3191;
assign x_2594 = v_3191 | ~v_261 | ~v_3243;
assign x_2595 = v_261 | ~v_3191 | ~v_3243;
assign x_2596 = v_3243 | ~v_262 | ~v_3192;
assign x_2597 = v_3192 | ~v_262 | ~v_3243;
assign x_2598 = v_262 | ~v_3192 | ~v_3243;
assign x_2599 = v_260 | v_261 | v_262 | ~v_3189 | ~v_3243;
assign x_2600 = v_259 | v_3190 | v_3191 | v_3192 | ~v_3243;
assign x_2601 = v_626 | v_3250 | ~v_3251;
assign x_2602 = v_3227 | ~v_626 | ~v_3251;
assign x_2603 = v_3227 | v_3250 | ~v_3251;
assign x_2604 = v_3251 | ~v_3227 | ~v_3250;
assign x_2605 = v_3251 | ~v_626 | ~v_3227;
assign x_2606 = v_626 | v_3251 | ~v_3250;
assign x_2607 = ~v_3255 | ~v_3256;
assign x_2608 = ~v_3255 | ~v_3257;
assign x_2609 = ~v_3256 | ~v_3257;
assign x_2610 = v_3255 | ~v_3120 | ~v_3259;
assign x_2611 = v_3120 | v_3256 | ~v_3259;
assign x_2612 = v_3255 | v_3256 | ~v_3259;
assign x_2613 = v_3259 | ~v_3255 | ~v_3256;
assign x_2614 = v_3120 | v_3259 | ~v_3256;
assign x_2615 = v_3259 | ~v_3120 | ~v_3255;
assign x_2616 = v_3256 | ~v_3120 | ~v_3260;
assign x_2617 = v_3120 | v_3257 | ~v_3260;
assign x_2618 = v_3256 | v_3257 | ~v_3260;
assign x_2619 = v_3260 | ~v_3256 | ~v_3257;
assign x_2620 = v_3120 | v_3260 | ~v_3257;
assign x_2621 = v_3260 | ~v_3120 | ~v_3256;
assign x_2622 = ~v_3258 | ~v_3259;
assign x_2623 = ~v_3258 | ~v_3260;
assign x_2624 = ~v_3258 | ~v_3261;
assign x_2625 = ~v_3259 | ~v_3260;
assign x_2626 = ~v_3259 | ~v_3261;
assign x_2627 = ~v_3260 | ~v_3261;
assign x_2628 = v_7 | v_538 | v_540 | v_543 | v_545 | v_553 | v_555 | v_558 | v_560 | v_570 | v_572 | v_575 | v_577 | v_938 | v_978 | v_1001 | v_1057 | v_1059 | v_1062 | v_1064 | v_1073 | v_1075 | v_1078 | v_1080 | v_1091 | v_1093 | v_1096 | v_1098 | v_1111 | v_1113 | v_1116 | v_1118 | v_1447 | v_1523 | v_1544 | v_1614 | v_1626 | v_1686 | v_1691 | v_1742 | v_1760 | v_1762 | v_1765 | v_1767 | v_1776 | v_1778 | v_1781 | v_1783 | v_1794 | v_1796 | v_1799 | v_1801 | v_1814 | v_1816 | v_1819 | v_1821 | v_2139 | v_2195 | v_2234 | v_2257 | v_2312 | v_2315 | v_2318 | v_2320 | v_2323 | v_2326 | v_2329 | v_2331 | v_2340 | v_2343 | v_2346 | v_2348 | v_2351 | v_2354 | v_2357 | v_2359 | v_2370 | v_2373 | v_2376 | v_2378 | v_2381 | v_2384 | v_2387 | v_2389 | v_2402 | v_2405 | v_2408 | v_2410 | v_2413 | v_2416 | v_2419 | v_2421 | v_2845 | v_2900 | v_2938 | v_2961 | v_2983 | v_3002 | v_3004 | v_3007 | v_3009 | v_3017 | v_3019 | v_3022 | v_3024 | v_3034 | v_3036 | v_3039 | v_3041 | ~v_3263;
assign x_2629 = x_1 & x_2;
assign x_2630 = x_4 & x_5;
assign x_2631 = x_3 & x_2630;
assign x_2632 = x_2629 & x_2631;
assign x_2633 = x_6 & x_7;
assign x_2634 = x_9 & x_10;
assign x_2635 = x_8 & x_2634;
assign x_2636 = x_2633 & x_2635;
assign x_2637 = x_2632 & x_2636;
assign x_2638 = x_11 & x_12;
assign x_2639 = x_14 & x_15;
assign x_2640 = x_13 & x_2639;
assign x_2641 = x_2638 & x_2640;
assign x_2642 = x_16 & x_17;
assign x_2643 = x_19 & x_20;
assign x_2644 = x_18 & x_2643;
assign x_2645 = x_2642 & x_2644;
assign x_2646 = x_2641 & x_2645;
assign x_2647 = x_2637 & x_2646;
assign x_2648 = x_21 & x_22;
assign x_2649 = x_24 & x_25;
assign x_2650 = x_23 & x_2649;
assign x_2651 = x_2648 & x_2650;
assign x_2652 = x_26 & x_27;
assign x_2653 = x_29 & x_30;
assign x_2654 = x_28 & x_2653;
assign x_2655 = x_2652 & x_2654;
assign x_2656 = x_2651 & x_2655;
assign x_2657 = x_31 & x_32;
assign x_2658 = x_34 & x_35;
assign x_2659 = x_33 & x_2658;
assign x_2660 = x_2657 & x_2659;
assign x_2661 = x_37 & x_38;
assign x_2662 = x_36 & x_2661;
assign x_2663 = x_40 & x_41;
assign x_2664 = x_39 & x_2663;
assign x_2665 = x_2662 & x_2664;
assign x_2666 = x_2660 & x_2665;
assign x_2667 = x_2656 & x_2666;
assign x_2668 = x_2647 & x_2667;
assign x_2669 = x_42 & x_43;
assign x_2670 = x_45 & x_46;
assign x_2671 = x_44 & x_2670;
assign x_2672 = x_2669 & x_2671;
assign x_2673 = x_47 & x_48;
assign x_2674 = x_50 & x_51;
assign x_2675 = x_49 & x_2674;
assign x_2676 = x_2673 & x_2675;
assign x_2677 = x_2672 & x_2676;
assign x_2678 = x_52 & x_53;
assign x_2679 = x_55 & x_56;
assign x_2680 = x_54 & x_2679;
assign x_2681 = x_2678 & x_2680;
assign x_2682 = x_57 & x_58;
assign x_2683 = x_60 & x_61;
assign x_2684 = x_59 & x_2683;
assign x_2685 = x_2682 & x_2684;
assign x_2686 = x_2681 & x_2685;
assign x_2687 = x_2677 & x_2686;
assign x_2688 = x_62 & x_63;
assign x_2689 = x_65 & x_66;
assign x_2690 = x_64 & x_2689;
assign x_2691 = x_2688 & x_2690;
assign x_2692 = x_67 & x_68;
assign x_2693 = x_70 & x_71;
assign x_2694 = x_69 & x_2693;
assign x_2695 = x_2692 & x_2694;
assign x_2696 = x_2691 & x_2695;
assign x_2697 = x_72 & x_73;
assign x_2698 = x_75 & x_76;
assign x_2699 = x_74 & x_2698;
assign x_2700 = x_2697 & x_2699;
assign x_2701 = x_78 & x_79;
assign x_2702 = x_77 & x_2701;
assign x_2703 = x_81 & x_82;
assign x_2704 = x_80 & x_2703;
assign x_2705 = x_2702 & x_2704;
assign x_2706 = x_2700 & x_2705;
assign x_2707 = x_2696 & x_2706;
assign x_2708 = x_2687 & x_2707;
assign x_2709 = x_2668 & x_2708;
assign x_2710 = x_83 & x_84;
assign x_2711 = x_86 & x_87;
assign x_2712 = x_85 & x_2711;
assign x_2713 = x_2710 & x_2712;
assign x_2714 = x_88 & x_89;
assign x_2715 = x_91 & x_92;
assign x_2716 = x_90 & x_2715;
assign x_2717 = x_2714 & x_2716;
assign x_2718 = x_2713 & x_2717;
assign x_2719 = x_93 & x_94;
assign x_2720 = x_96 & x_97;
assign x_2721 = x_95 & x_2720;
assign x_2722 = x_2719 & x_2721;
assign x_2723 = x_98 & x_99;
assign x_2724 = x_101 & x_102;
assign x_2725 = x_100 & x_2724;
assign x_2726 = x_2723 & x_2725;
assign x_2727 = x_2722 & x_2726;
assign x_2728 = x_2718 & x_2727;
assign x_2729 = x_103 & x_104;
assign x_2730 = x_106 & x_107;
assign x_2731 = x_105 & x_2730;
assign x_2732 = x_2729 & x_2731;
assign x_2733 = x_108 & x_109;
assign x_2734 = x_111 & x_112;
assign x_2735 = x_110 & x_2734;
assign x_2736 = x_2733 & x_2735;
assign x_2737 = x_2732 & x_2736;
assign x_2738 = x_113 & x_114;
assign x_2739 = x_116 & x_117;
assign x_2740 = x_115 & x_2739;
assign x_2741 = x_2738 & x_2740;
assign x_2742 = x_119 & x_120;
assign x_2743 = x_118 & x_2742;
assign x_2744 = x_122 & x_123;
assign x_2745 = x_121 & x_2744;
assign x_2746 = x_2743 & x_2745;
assign x_2747 = x_2741 & x_2746;
assign x_2748 = x_2737 & x_2747;
assign x_2749 = x_2728 & x_2748;
assign x_2750 = x_124 & x_125;
assign x_2751 = x_127 & x_128;
assign x_2752 = x_126 & x_2751;
assign x_2753 = x_2750 & x_2752;
assign x_2754 = x_129 & x_130;
assign x_2755 = x_132 & x_133;
assign x_2756 = x_131 & x_2755;
assign x_2757 = x_2754 & x_2756;
assign x_2758 = x_2753 & x_2757;
assign x_2759 = x_134 & x_135;
assign x_2760 = x_137 & x_138;
assign x_2761 = x_136 & x_2760;
assign x_2762 = x_2759 & x_2761;
assign x_2763 = x_139 & x_140;
assign x_2764 = x_142 & x_143;
assign x_2765 = x_141 & x_2764;
assign x_2766 = x_2763 & x_2765;
assign x_2767 = x_2762 & x_2766;
assign x_2768 = x_2758 & x_2767;
assign x_2769 = x_144 & x_145;
assign x_2770 = x_147 & x_148;
assign x_2771 = x_146 & x_2770;
assign x_2772 = x_2769 & x_2771;
assign x_2773 = x_149 & x_150;
assign x_2774 = x_152 & x_153;
assign x_2775 = x_151 & x_2774;
assign x_2776 = x_2773 & x_2775;
assign x_2777 = x_2772 & x_2776;
assign x_2778 = x_154 & x_155;
assign x_2779 = x_157 & x_158;
assign x_2780 = x_156 & x_2779;
assign x_2781 = x_2778 & x_2780;
assign x_2782 = x_160 & x_161;
assign x_2783 = x_159 & x_2782;
assign x_2784 = x_163 & x_164;
assign x_2785 = x_162 & x_2784;
assign x_2786 = x_2783 & x_2785;
assign x_2787 = x_2781 & x_2786;
assign x_2788 = x_2777 & x_2787;
assign x_2789 = x_2768 & x_2788;
assign x_2790 = x_2749 & x_2789;
assign x_2791 = x_2709 & x_2790;
assign x_2792 = x_165 & x_166;
assign x_2793 = x_168 & x_169;
assign x_2794 = x_167 & x_2793;
assign x_2795 = x_2792 & x_2794;
assign x_2796 = x_170 & x_171;
assign x_2797 = x_173 & x_174;
assign x_2798 = x_172 & x_2797;
assign x_2799 = x_2796 & x_2798;
assign x_2800 = x_2795 & x_2799;
assign x_2801 = x_175 & x_176;
assign x_2802 = x_178 & x_179;
assign x_2803 = x_177 & x_2802;
assign x_2804 = x_2801 & x_2803;
assign x_2805 = x_180 & x_181;
assign x_2806 = x_183 & x_184;
assign x_2807 = x_182 & x_2806;
assign x_2808 = x_2805 & x_2807;
assign x_2809 = x_2804 & x_2808;
assign x_2810 = x_2800 & x_2809;
assign x_2811 = x_185 & x_186;
assign x_2812 = x_188 & x_189;
assign x_2813 = x_187 & x_2812;
assign x_2814 = x_2811 & x_2813;
assign x_2815 = x_190 & x_191;
assign x_2816 = x_193 & x_194;
assign x_2817 = x_192 & x_2816;
assign x_2818 = x_2815 & x_2817;
assign x_2819 = x_2814 & x_2818;
assign x_2820 = x_195 & x_196;
assign x_2821 = x_198 & x_199;
assign x_2822 = x_197 & x_2821;
assign x_2823 = x_2820 & x_2822;
assign x_2824 = x_201 & x_202;
assign x_2825 = x_200 & x_2824;
assign x_2826 = x_204 & x_205;
assign x_2827 = x_203 & x_2826;
assign x_2828 = x_2825 & x_2827;
assign x_2829 = x_2823 & x_2828;
assign x_2830 = x_2819 & x_2829;
assign x_2831 = x_2810 & x_2830;
assign x_2832 = x_206 & x_207;
assign x_2833 = x_209 & x_210;
assign x_2834 = x_208 & x_2833;
assign x_2835 = x_2832 & x_2834;
assign x_2836 = x_211 & x_212;
assign x_2837 = x_214 & x_215;
assign x_2838 = x_213 & x_2837;
assign x_2839 = x_2836 & x_2838;
assign x_2840 = x_2835 & x_2839;
assign x_2841 = x_216 & x_217;
assign x_2842 = x_219 & x_220;
assign x_2843 = x_218 & x_2842;
assign x_2844 = x_2841 & x_2843;
assign x_2845 = x_221 & x_222;
assign x_2846 = x_224 & x_225;
assign x_2847 = x_223 & x_2846;
assign x_2848 = x_2845 & x_2847;
assign x_2849 = x_2844 & x_2848;
assign x_2850 = x_2840 & x_2849;
assign x_2851 = x_226 & x_227;
assign x_2852 = x_229 & x_230;
assign x_2853 = x_228 & x_2852;
assign x_2854 = x_2851 & x_2853;
assign x_2855 = x_231 & x_232;
assign x_2856 = x_234 & x_235;
assign x_2857 = x_233 & x_2856;
assign x_2858 = x_2855 & x_2857;
assign x_2859 = x_2854 & x_2858;
assign x_2860 = x_236 & x_237;
assign x_2861 = x_239 & x_240;
assign x_2862 = x_238 & x_2861;
assign x_2863 = x_2860 & x_2862;
assign x_2864 = x_242 & x_243;
assign x_2865 = x_241 & x_2864;
assign x_2866 = x_245 & x_246;
assign x_2867 = x_244 & x_2866;
assign x_2868 = x_2865 & x_2867;
assign x_2869 = x_2863 & x_2868;
assign x_2870 = x_2859 & x_2869;
assign x_2871 = x_2850 & x_2870;
assign x_2872 = x_2831 & x_2871;
assign x_2873 = x_247 & x_248;
assign x_2874 = x_250 & x_251;
assign x_2875 = x_249 & x_2874;
assign x_2876 = x_2873 & x_2875;
assign x_2877 = x_252 & x_253;
assign x_2878 = x_255 & x_256;
assign x_2879 = x_254 & x_2878;
assign x_2880 = x_2877 & x_2879;
assign x_2881 = x_2876 & x_2880;
assign x_2882 = x_257 & x_258;
assign x_2883 = x_260 & x_261;
assign x_2884 = x_259 & x_2883;
assign x_2885 = x_2882 & x_2884;
assign x_2886 = x_262 & x_263;
assign x_2887 = x_265 & x_266;
assign x_2888 = x_264 & x_2887;
assign x_2889 = x_2886 & x_2888;
assign x_2890 = x_2885 & x_2889;
assign x_2891 = x_2881 & x_2890;
assign x_2892 = x_267 & x_268;
assign x_2893 = x_270 & x_271;
assign x_2894 = x_269 & x_2893;
assign x_2895 = x_2892 & x_2894;
assign x_2896 = x_272 & x_273;
assign x_2897 = x_275 & x_276;
assign x_2898 = x_274 & x_2897;
assign x_2899 = x_2896 & x_2898;
assign x_2900 = x_2895 & x_2899;
assign x_2901 = x_277 & x_278;
assign x_2902 = x_280 & x_281;
assign x_2903 = x_279 & x_2902;
assign x_2904 = x_2901 & x_2903;
assign x_2905 = x_283 & x_284;
assign x_2906 = x_282 & x_2905;
assign x_2907 = x_286 & x_287;
assign x_2908 = x_285 & x_2907;
assign x_2909 = x_2906 & x_2908;
assign x_2910 = x_2904 & x_2909;
assign x_2911 = x_2900 & x_2910;
assign x_2912 = x_2891 & x_2911;
assign x_2913 = x_288 & x_289;
assign x_2914 = x_291 & x_292;
assign x_2915 = x_290 & x_2914;
assign x_2916 = x_2913 & x_2915;
assign x_2917 = x_293 & x_294;
assign x_2918 = x_296 & x_297;
assign x_2919 = x_295 & x_2918;
assign x_2920 = x_2917 & x_2919;
assign x_2921 = x_2916 & x_2920;
assign x_2922 = x_298 & x_299;
assign x_2923 = x_301 & x_302;
assign x_2924 = x_300 & x_2923;
assign x_2925 = x_2922 & x_2924;
assign x_2926 = x_303 & x_304;
assign x_2927 = x_306 & x_307;
assign x_2928 = x_305 & x_2927;
assign x_2929 = x_2926 & x_2928;
assign x_2930 = x_2925 & x_2929;
assign x_2931 = x_2921 & x_2930;
assign x_2932 = x_308 & x_309;
assign x_2933 = x_311 & x_312;
assign x_2934 = x_310 & x_2933;
assign x_2935 = x_2932 & x_2934;
assign x_2936 = x_313 & x_314;
assign x_2937 = x_316 & x_317;
assign x_2938 = x_315 & x_2937;
assign x_2939 = x_2936 & x_2938;
assign x_2940 = x_2935 & x_2939;
assign x_2941 = x_318 & x_319;
assign x_2942 = x_321 & x_322;
assign x_2943 = x_320 & x_2942;
assign x_2944 = x_2941 & x_2943;
assign x_2945 = x_324 & x_325;
assign x_2946 = x_323 & x_2945;
assign x_2947 = x_327 & x_328;
assign x_2948 = x_326 & x_2947;
assign x_2949 = x_2946 & x_2948;
assign x_2950 = x_2944 & x_2949;
assign x_2951 = x_2940 & x_2950;
assign x_2952 = x_2931 & x_2951;
assign x_2953 = x_2912 & x_2952;
assign x_2954 = x_2872 & x_2953;
assign x_2955 = x_2791 & x_2954;
assign x_2956 = x_329 & x_330;
assign x_2957 = x_332 & x_333;
assign x_2958 = x_331 & x_2957;
assign x_2959 = x_2956 & x_2958;
assign x_2960 = x_334 & x_335;
assign x_2961 = x_337 & x_338;
assign x_2962 = x_336 & x_2961;
assign x_2963 = x_2960 & x_2962;
assign x_2964 = x_2959 & x_2963;
assign x_2965 = x_339 & x_340;
assign x_2966 = x_342 & x_343;
assign x_2967 = x_341 & x_2966;
assign x_2968 = x_2965 & x_2967;
assign x_2969 = x_344 & x_345;
assign x_2970 = x_347 & x_348;
assign x_2971 = x_346 & x_2970;
assign x_2972 = x_2969 & x_2971;
assign x_2973 = x_2968 & x_2972;
assign x_2974 = x_2964 & x_2973;
assign x_2975 = x_349 & x_350;
assign x_2976 = x_352 & x_353;
assign x_2977 = x_351 & x_2976;
assign x_2978 = x_2975 & x_2977;
assign x_2979 = x_354 & x_355;
assign x_2980 = x_357 & x_358;
assign x_2981 = x_356 & x_2980;
assign x_2982 = x_2979 & x_2981;
assign x_2983 = x_2978 & x_2982;
assign x_2984 = x_359 & x_360;
assign x_2985 = x_362 & x_363;
assign x_2986 = x_361 & x_2985;
assign x_2987 = x_2984 & x_2986;
assign x_2988 = x_365 & x_366;
assign x_2989 = x_364 & x_2988;
assign x_2990 = x_368 & x_369;
assign x_2991 = x_367 & x_2990;
assign x_2992 = x_2989 & x_2991;
assign x_2993 = x_2987 & x_2992;
assign x_2994 = x_2983 & x_2993;
assign x_2995 = x_2974 & x_2994;
assign x_2996 = x_370 & x_371;
assign x_2997 = x_373 & x_374;
assign x_2998 = x_372 & x_2997;
assign x_2999 = x_2996 & x_2998;
assign x_3000 = x_375 & x_376;
assign x_3001 = x_378 & x_379;
assign x_3002 = x_377 & x_3001;
assign x_3003 = x_3000 & x_3002;
assign x_3004 = x_2999 & x_3003;
assign x_3005 = x_380 & x_381;
assign x_3006 = x_383 & x_384;
assign x_3007 = x_382 & x_3006;
assign x_3008 = x_3005 & x_3007;
assign x_3009 = x_385 & x_386;
assign x_3010 = x_388 & x_389;
assign x_3011 = x_387 & x_3010;
assign x_3012 = x_3009 & x_3011;
assign x_3013 = x_3008 & x_3012;
assign x_3014 = x_3004 & x_3013;
assign x_3015 = x_390 & x_391;
assign x_3016 = x_393 & x_394;
assign x_3017 = x_392 & x_3016;
assign x_3018 = x_3015 & x_3017;
assign x_3019 = x_395 & x_396;
assign x_3020 = x_398 & x_399;
assign x_3021 = x_397 & x_3020;
assign x_3022 = x_3019 & x_3021;
assign x_3023 = x_3018 & x_3022;
assign x_3024 = x_400 & x_401;
assign x_3025 = x_403 & x_404;
assign x_3026 = x_402 & x_3025;
assign x_3027 = x_3024 & x_3026;
assign x_3028 = x_406 & x_407;
assign x_3029 = x_405 & x_3028;
assign x_3030 = x_409 & x_410;
assign x_3031 = x_408 & x_3030;
assign x_3032 = x_3029 & x_3031;
assign x_3033 = x_3027 & x_3032;
assign x_3034 = x_3023 & x_3033;
assign x_3035 = x_3014 & x_3034;
assign x_3036 = x_2995 & x_3035;
assign x_3037 = x_411 & x_412;
assign x_3038 = x_414 & x_415;
assign x_3039 = x_413 & x_3038;
assign x_3040 = x_3037 & x_3039;
assign x_3041 = x_416 & x_417;
assign x_3042 = x_419 & x_420;
assign x_3043 = x_418 & x_3042;
assign x_3044 = x_3041 & x_3043;
assign x_3045 = x_3040 & x_3044;
assign x_3046 = x_421 & x_422;
assign x_3047 = x_424 & x_425;
assign x_3048 = x_423 & x_3047;
assign x_3049 = x_3046 & x_3048;
assign x_3050 = x_426 & x_427;
assign x_3051 = x_429 & x_430;
assign x_3052 = x_428 & x_3051;
assign x_3053 = x_3050 & x_3052;
assign x_3054 = x_3049 & x_3053;
assign x_3055 = x_3045 & x_3054;
assign x_3056 = x_431 & x_432;
assign x_3057 = x_434 & x_435;
assign x_3058 = x_433 & x_3057;
assign x_3059 = x_3056 & x_3058;
assign x_3060 = x_436 & x_437;
assign x_3061 = x_439 & x_440;
assign x_3062 = x_438 & x_3061;
assign x_3063 = x_3060 & x_3062;
assign x_3064 = x_3059 & x_3063;
assign x_3065 = x_441 & x_442;
assign x_3066 = x_444 & x_445;
assign x_3067 = x_443 & x_3066;
assign x_3068 = x_3065 & x_3067;
assign x_3069 = x_447 & x_448;
assign x_3070 = x_446 & x_3069;
assign x_3071 = x_450 & x_451;
assign x_3072 = x_449 & x_3071;
assign x_3073 = x_3070 & x_3072;
assign x_3074 = x_3068 & x_3073;
assign x_3075 = x_3064 & x_3074;
assign x_3076 = x_3055 & x_3075;
assign x_3077 = x_452 & x_453;
assign x_3078 = x_455 & x_456;
assign x_3079 = x_454 & x_3078;
assign x_3080 = x_3077 & x_3079;
assign x_3081 = x_457 & x_458;
assign x_3082 = x_460 & x_461;
assign x_3083 = x_459 & x_3082;
assign x_3084 = x_3081 & x_3083;
assign x_3085 = x_3080 & x_3084;
assign x_3086 = x_462 & x_463;
assign x_3087 = x_465 & x_466;
assign x_3088 = x_464 & x_3087;
assign x_3089 = x_3086 & x_3088;
assign x_3090 = x_467 & x_468;
assign x_3091 = x_470 & x_471;
assign x_3092 = x_469 & x_3091;
assign x_3093 = x_3090 & x_3092;
assign x_3094 = x_3089 & x_3093;
assign x_3095 = x_3085 & x_3094;
assign x_3096 = x_472 & x_473;
assign x_3097 = x_475 & x_476;
assign x_3098 = x_474 & x_3097;
assign x_3099 = x_3096 & x_3098;
assign x_3100 = x_477 & x_478;
assign x_3101 = x_480 & x_481;
assign x_3102 = x_479 & x_3101;
assign x_3103 = x_3100 & x_3102;
assign x_3104 = x_3099 & x_3103;
assign x_3105 = x_482 & x_483;
assign x_3106 = x_485 & x_486;
assign x_3107 = x_484 & x_3106;
assign x_3108 = x_3105 & x_3107;
assign x_3109 = x_488 & x_489;
assign x_3110 = x_487 & x_3109;
assign x_3111 = x_491 & x_492;
assign x_3112 = x_490 & x_3111;
assign x_3113 = x_3110 & x_3112;
assign x_3114 = x_3108 & x_3113;
assign x_3115 = x_3104 & x_3114;
assign x_3116 = x_3095 & x_3115;
assign x_3117 = x_3076 & x_3116;
assign x_3118 = x_3036 & x_3117;
assign x_3119 = x_493 & x_494;
assign x_3120 = x_496 & x_497;
assign x_3121 = x_495 & x_3120;
assign x_3122 = x_3119 & x_3121;
assign x_3123 = x_498 & x_499;
assign x_3124 = x_501 & x_502;
assign x_3125 = x_500 & x_3124;
assign x_3126 = x_3123 & x_3125;
assign x_3127 = x_3122 & x_3126;
assign x_3128 = x_503 & x_504;
assign x_3129 = x_506 & x_507;
assign x_3130 = x_505 & x_3129;
assign x_3131 = x_3128 & x_3130;
assign x_3132 = x_508 & x_509;
assign x_3133 = x_511 & x_512;
assign x_3134 = x_510 & x_3133;
assign x_3135 = x_3132 & x_3134;
assign x_3136 = x_3131 & x_3135;
assign x_3137 = x_3127 & x_3136;
assign x_3138 = x_513 & x_514;
assign x_3139 = x_516 & x_517;
assign x_3140 = x_515 & x_3139;
assign x_3141 = x_3138 & x_3140;
assign x_3142 = x_518 & x_519;
assign x_3143 = x_521 & x_522;
assign x_3144 = x_520 & x_3143;
assign x_3145 = x_3142 & x_3144;
assign x_3146 = x_3141 & x_3145;
assign x_3147 = x_523 & x_524;
assign x_3148 = x_526 & x_527;
assign x_3149 = x_525 & x_3148;
assign x_3150 = x_3147 & x_3149;
assign x_3151 = x_529 & x_530;
assign x_3152 = x_528 & x_3151;
assign x_3153 = x_532 & x_533;
assign x_3154 = x_531 & x_3153;
assign x_3155 = x_3152 & x_3154;
assign x_3156 = x_3150 & x_3155;
assign x_3157 = x_3146 & x_3156;
assign x_3158 = x_3137 & x_3157;
assign x_3159 = x_534 & x_535;
assign x_3160 = x_537 & x_538;
assign x_3161 = x_536 & x_3160;
assign x_3162 = x_3159 & x_3161;
assign x_3163 = x_539 & x_540;
assign x_3164 = x_542 & x_543;
assign x_3165 = x_541 & x_3164;
assign x_3166 = x_3163 & x_3165;
assign x_3167 = x_3162 & x_3166;
assign x_3168 = x_544 & x_545;
assign x_3169 = x_547 & x_548;
assign x_3170 = x_546 & x_3169;
assign x_3171 = x_3168 & x_3170;
assign x_3172 = x_549 & x_550;
assign x_3173 = x_552 & x_553;
assign x_3174 = x_551 & x_3173;
assign x_3175 = x_3172 & x_3174;
assign x_3176 = x_3171 & x_3175;
assign x_3177 = x_3167 & x_3176;
assign x_3178 = x_554 & x_555;
assign x_3179 = x_557 & x_558;
assign x_3180 = x_556 & x_3179;
assign x_3181 = x_3178 & x_3180;
assign x_3182 = x_559 & x_560;
assign x_3183 = x_562 & x_563;
assign x_3184 = x_561 & x_3183;
assign x_3185 = x_3182 & x_3184;
assign x_3186 = x_3181 & x_3185;
assign x_3187 = x_564 & x_565;
assign x_3188 = x_567 & x_568;
assign x_3189 = x_566 & x_3188;
assign x_3190 = x_3187 & x_3189;
assign x_3191 = x_570 & x_571;
assign x_3192 = x_569 & x_3191;
assign x_3193 = x_573 & x_574;
assign x_3194 = x_572 & x_3193;
assign x_3195 = x_3192 & x_3194;
assign x_3196 = x_3190 & x_3195;
assign x_3197 = x_3186 & x_3196;
assign x_3198 = x_3177 & x_3197;
assign x_3199 = x_3158 & x_3198;
assign x_3200 = x_575 & x_576;
assign x_3201 = x_578 & x_579;
assign x_3202 = x_577 & x_3201;
assign x_3203 = x_3200 & x_3202;
assign x_3204 = x_580 & x_581;
assign x_3205 = x_583 & x_584;
assign x_3206 = x_582 & x_3205;
assign x_3207 = x_3204 & x_3206;
assign x_3208 = x_3203 & x_3207;
assign x_3209 = x_585 & x_586;
assign x_3210 = x_588 & x_589;
assign x_3211 = x_587 & x_3210;
assign x_3212 = x_3209 & x_3211;
assign x_3213 = x_590 & x_591;
assign x_3214 = x_593 & x_594;
assign x_3215 = x_592 & x_3214;
assign x_3216 = x_3213 & x_3215;
assign x_3217 = x_3212 & x_3216;
assign x_3218 = x_3208 & x_3217;
assign x_3219 = x_595 & x_596;
assign x_3220 = x_598 & x_599;
assign x_3221 = x_597 & x_3220;
assign x_3222 = x_3219 & x_3221;
assign x_3223 = x_600 & x_601;
assign x_3224 = x_603 & x_604;
assign x_3225 = x_602 & x_3224;
assign x_3226 = x_3223 & x_3225;
assign x_3227 = x_3222 & x_3226;
assign x_3228 = x_605 & x_606;
assign x_3229 = x_608 & x_609;
assign x_3230 = x_607 & x_3229;
assign x_3231 = x_3228 & x_3230;
assign x_3232 = x_611 & x_612;
assign x_3233 = x_610 & x_3232;
assign x_3234 = x_614 & x_615;
assign x_3235 = x_613 & x_3234;
assign x_3236 = x_3233 & x_3235;
assign x_3237 = x_3231 & x_3236;
assign x_3238 = x_3227 & x_3237;
assign x_3239 = x_3218 & x_3238;
assign x_3240 = x_616 & x_617;
assign x_3241 = x_619 & x_620;
assign x_3242 = x_618 & x_3241;
assign x_3243 = x_3240 & x_3242;
assign x_3244 = x_621 & x_622;
assign x_3245 = x_624 & x_625;
assign x_3246 = x_623 & x_3245;
assign x_3247 = x_3244 & x_3246;
assign x_3248 = x_3243 & x_3247;
assign x_3249 = x_626 & x_627;
assign x_3250 = x_629 & x_630;
assign x_3251 = x_628 & x_3250;
assign x_3252 = x_3249 & x_3251;
assign x_3253 = x_632 & x_633;
assign x_3254 = x_631 & x_3253;
assign x_3255 = x_635 & x_636;
assign x_3256 = x_634 & x_3255;
assign x_3257 = x_3254 & x_3256;
assign x_3258 = x_3252 & x_3257;
assign x_3259 = x_3248 & x_3258;
assign x_3260 = x_637 & x_638;
assign x_3261 = x_640 & x_641;
assign x_3262 = x_639 & x_3261;
assign x_3263 = x_3260 & x_3262;
assign x_3264 = x_642 & x_643;
assign x_3265 = x_645 & x_646;
assign x_3266 = x_644 & x_3265;
assign x_3267 = x_3264 & x_3266;
assign x_3268 = x_3263 & x_3267;
assign x_3269 = x_647 & x_648;
assign x_3270 = x_650 & x_651;
assign x_3271 = x_649 & x_3270;
assign x_3272 = x_3269 & x_3271;
assign x_3273 = x_653 & x_654;
assign x_3274 = x_652 & x_3273;
assign x_3275 = x_656 & x_657;
assign x_3276 = x_655 & x_3275;
assign x_3277 = x_3274 & x_3276;
assign x_3278 = x_3272 & x_3277;
assign x_3279 = x_3268 & x_3278;
assign x_3280 = x_3259 & x_3279;
assign x_3281 = x_3239 & x_3280;
assign x_3282 = x_3199 & x_3281;
assign x_3283 = x_3118 & x_3282;
assign x_3284 = x_2955 & x_3283;
assign x_3285 = x_658 & x_659;
assign x_3286 = x_661 & x_662;
assign x_3287 = x_660 & x_3286;
assign x_3288 = x_3285 & x_3287;
assign x_3289 = x_663 & x_664;
assign x_3290 = x_666 & x_667;
assign x_3291 = x_665 & x_3290;
assign x_3292 = x_3289 & x_3291;
assign x_3293 = x_3288 & x_3292;
assign x_3294 = x_668 & x_669;
assign x_3295 = x_671 & x_672;
assign x_3296 = x_670 & x_3295;
assign x_3297 = x_3294 & x_3296;
assign x_3298 = x_673 & x_674;
assign x_3299 = x_676 & x_677;
assign x_3300 = x_675 & x_3299;
assign x_3301 = x_3298 & x_3300;
assign x_3302 = x_3297 & x_3301;
assign x_3303 = x_3293 & x_3302;
assign x_3304 = x_678 & x_679;
assign x_3305 = x_681 & x_682;
assign x_3306 = x_680 & x_3305;
assign x_3307 = x_3304 & x_3306;
assign x_3308 = x_683 & x_684;
assign x_3309 = x_686 & x_687;
assign x_3310 = x_685 & x_3309;
assign x_3311 = x_3308 & x_3310;
assign x_3312 = x_3307 & x_3311;
assign x_3313 = x_688 & x_689;
assign x_3314 = x_691 & x_692;
assign x_3315 = x_690 & x_3314;
assign x_3316 = x_3313 & x_3315;
assign x_3317 = x_694 & x_695;
assign x_3318 = x_693 & x_3317;
assign x_3319 = x_697 & x_698;
assign x_3320 = x_696 & x_3319;
assign x_3321 = x_3318 & x_3320;
assign x_3322 = x_3316 & x_3321;
assign x_3323 = x_3312 & x_3322;
assign x_3324 = x_3303 & x_3323;
assign x_3325 = x_699 & x_700;
assign x_3326 = x_702 & x_703;
assign x_3327 = x_701 & x_3326;
assign x_3328 = x_3325 & x_3327;
assign x_3329 = x_704 & x_705;
assign x_3330 = x_707 & x_708;
assign x_3331 = x_706 & x_3330;
assign x_3332 = x_3329 & x_3331;
assign x_3333 = x_3328 & x_3332;
assign x_3334 = x_709 & x_710;
assign x_3335 = x_712 & x_713;
assign x_3336 = x_711 & x_3335;
assign x_3337 = x_3334 & x_3336;
assign x_3338 = x_714 & x_715;
assign x_3339 = x_717 & x_718;
assign x_3340 = x_716 & x_3339;
assign x_3341 = x_3338 & x_3340;
assign x_3342 = x_3337 & x_3341;
assign x_3343 = x_3333 & x_3342;
assign x_3344 = x_719 & x_720;
assign x_3345 = x_722 & x_723;
assign x_3346 = x_721 & x_3345;
assign x_3347 = x_3344 & x_3346;
assign x_3348 = x_724 & x_725;
assign x_3349 = x_727 & x_728;
assign x_3350 = x_726 & x_3349;
assign x_3351 = x_3348 & x_3350;
assign x_3352 = x_3347 & x_3351;
assign x_3353 = x_729 & x_730;
assign x_3354 = x_732 & x_733;
assign x_3355 = x_731 & x_3354;
assign x_3356 = x_3353 & x_3355;
assign x_3357 = x_735 & x_736;
assign x_3358 = x_734 & x_3357;
assign x_3359 = x_738 & x_739;
assign x_3360 = x_737 & x_3359;
assign x_3361 = x_3358 & x_3360;
assign x_3362 = x_3356 & x_3361;
assign x_3363 = x_3352 & x_3362;
assign x_3364 = x_3343 & x_3363;
assign x_3365 = x_3324 & x_3364;
assign x_3366 = x_740 & x_741;
assign x_3367 = x_743 & x_744;
assign x_3368 = x_742 & x_3367;
assign x_3369 = x_3366 & x_3368;
assign x_3370 = x_745 & x_746;
assign x_3371 = x_748 & x_749;
assign x_3372 = x_747 & x_3371;
assign x_3373 = x_3370 & x_3372;
assign x_3374 = x_3369 & x_3373;
assign x_3375 = x_750 & x_751;
assign x_3376 = x_753 & x_754;
assign x_3377 = x_752 & x_3376;
assign x_3378 = x_3375 & x_3377;
assign x_3379 = x_755 & x_756;
assign x_3380 = x_758 & x_759;
assign x_3381 = x_757 & x_3380;
assign x_3382 = x_3379 & x_3381;
assign x_3383 = x_3378 & x_3382;
assign x_3384 = x_3374 & x_3383;
assign x_3385 = x_760 & x_761;
assign x_3386 = x_763 & x_764;
assign x_3387 = x_762 & x_3386;
assign x_3388 = x_3385 & x_3387;
assign x_3389 = x_765 & x_766;
assign x_3390 = x_768 & x_769;
assign x_3391 = x_767 & x_3390;
assign x_3392 = x_3389 & x_3391;
assign x_3393 = x_3388 & x_3392;
assign x_3394 = x_770 & x_771;
assign x_3395 = x_773 & x_774;
assign x_3396 = x_772 & x_3395;
assign x_3397 = x_3394 & x_3396;
assign x_3398 = x_776 & x_777;
assign x_3399 = x_775 & x_3398;
assign x_3400 = x_779 & x_780;
assign x_3401 = x_778 & x_3400;
assign x_3402 = x_3399 & x_3401;
assign x_3403 = x_3397 & x_3402;
assign x_3404 = x_3393 & x_3403;
assign x_3405 = x_3384 & x_3404;
assign x_3406 = x_781 & x_782;
assign x_3407 = x_784 & x_785;
assign x_3408 = x_783 & x_3407;
assign x_3409 = x_3406 & x_3408;
assign x_3410 = x_786 & x_787;
assign x_3411 = x_789 & x_790;
assign x_3412 = x_788 & x_3411;
assign x_3413 = x_3410 & x_3412;
assign x_3414 = x_3409 & x_3413;
assign x_3415 = x_791 & x_792;
assign x_3416 = x_794 & x_795;
assign x_3417 = x_793 & x_3416;
assign x_3418 = x_3415 & x_3417;
assign x_3419 = x_796 & x_797;
assign x_3420 = x_799 & x_800;
assign x_3421 = x_798 & x_3420;
assign x_3422 = x_3419 & x_3421;
assign x_3423 = x_3418 & x_3422;
assign x_3424 = x_3414 & x_3423;
assign x_3425 = x_801 & x_802;
assign x_3426 = x_804 & x_805;
assign x_3427 = x_803 & x_3426;
assign x_3428 = x_3425 & x_3427;
assign x_3429 = x_806 & x_807;
assign x_3430 = x_809 & x_810;
assign x_3431 = x_808 & x_3430;
assign x_3432 = x_3429 & x_3431;
assign x_3433 = x_3428 & x_3432;
assign x_3434 = x_811 & x_812;
assign x_3435 = x_814 & x_815;
assign x_3436 = x_813 & x_3435;
assign x_3437 = x_3434 & x_3436;
assign x_3438 = x_817 & x_818;
assign x_3439 = x_816 & x_3438;
assign x_3440 = x_820 & x_821;
assign x_3441 = x_819 & x_3440;
assign x_3442 = x_3439 & x_3441;
assign x_3443 = x_3437 & x_3442;
assign x_3444 = x_3433 & x_3443;
assign x_3445 = x_3424 & x_3444;
assign x_3446 = x_3405 & x_3445;
assign x_3447 = x_3365 & x_3446;
assign x_3448 = x_822 & x_823;
assign x_3449 = x_825 & x_826;
assign x_3450 = x_824 & x_3449;
assign x_3451 = x_3448 & x_3450;
assign x_3452 = x_827 & x_828;
assign x_3453 = x_830 & x_831;
assign x_3454 = x_829 & x_3453;
assign x_3455 = x_3452 & x_3454;
assign x_3456 = x_3451 & x_3455;
assign x_3457 = x_832 & x_833;
assign x_3458 = x_835 & x_836;
assign x_3459 = x_834 & x_3458;
assign x_3460 = x_3457 & x_3459;
assign x_3461 = x_837 & x_838;
assign x_3462 = x_840 & x_841;
assign x_3463 = x_839 & x_3462;
assign x_3464 = x_3461 & x_3463;
assign x_3465 = x_3460 & x_3464;
assign x_3466 = x_3456 & x_3465;
assign x_3467 = x_842 & x_843;
assign x_3468 = x_845 & x_846;
assign x_3469 = x_844 & x_3468;
assign x_3470 = x_3467 & x_3469;
assign x_3471 = x_847 & x_848;
assign x_3472 = x_850 & x_851;
assign x_3473 = x_849 & x_3472;
assign x_3474 = x_3471 & x_3473;
assign x_3475 = x_3470 & x_3474;
assign x_3476 = x_852 & x_853;
assign x_3477 = x_855 & x_856;
assign x_3478 = x_854 & x_3477;
assign x_3479 = x_3476 & x_3478;
assign x_3480 = x_858 & x_859;
assign x_3481 = x_857 & x_3480;
assign x_3482 = x_861 & x_862;
assign x_3483 = x_860 & x_3482;
assign x_3484 = x_3481 & x_3483;
assign x_3485 = x_3479 & x_3484;
assign x_3486 = x_3475 & x_3485;
assign x_3487 = x_3466 & x_3486;
assign x_3488 = x_863 & x_864;
assign x_3489 = x_866 & x_867;
assign x_3490 = x_865 & x_3489;
assign x_3491 = x_3488 & x_3490;
assign x_3492 = x_868 & x_869;
assign x_3493 = x_871 & x_872;
assign x_3494 = x_870 & x_3493;
assign x_3495 = x_3492 & x_3494;
assign x_3496 = x_3491 & x_3495;
assign x_3497 = x_873 & x_874;
assign x_3498 = x_876 & x_877;
assign x_3499 = x_875 & x_3498;
assign x_3500 = x_3497 & x_3499;
assign x_3501 = x_878 & x_879;
assign x_3502 = x_881 & x_882;
assign x_3503 = x_880 & x_3502;
assign x_3504 = x_3501 & x_3503;
assign x_3505 = x_3500 & x_3504;
assign x_3506 = x_3496 & x_3505;
assign x_3507 = x_883 & x_884;
assign x_3508 = x_886 & x_887;
assign x_3509 = x_885 & x_3508;
assign x_3510 = x_3507 & x_3509;
assign x_3511 = x_888 & x_889;
assign x_3512 = x_891 & x_892;
assign x_3513 = x_890 & x_3512;
assign x_3514 = x_3511 & x_3513;
assign x_3515 = x_3510 & x_3514;
assign x_3516 = x_893 & x_894;
assign x_3517 = x_896 & x_897;
assign x_3518 = x_895 & x_3517;
assign x_3519 = x_3516 & x_3518;
assign x_3520 = x_899 & x_900;
assign x_3521 = x_898 & x_3520;
assign x_3522 = x_902 & x_903;
assign x_3523 = x_901 & x_3522;
assign x_3524 = x_3521 & x_3523;
assign x_3525 = x_3519 & x_3524;
assign x_3526 = x_3515 & x_3525;
assign x_3527 = x_3506 & x_3526;
assign x_3528 = x_3487 & x_3527;
assign x_3529 = x_904 & x_905;
assign x_3530 = x_907 & x_908;
assign x_3531 = x_906 & x_3530;
assign x_3532 = x_3529 & x_3531;
assign x_3533 = x_909 & x_910;
assign x_3534 = x_912 & x_913;
assign x_3535 = x_911 & x_3534;
assign x_3536 = x_3533 & x_3535;
assign x_3537 = x_3532 & x_3536;
assign x_3538 = x_914 & x_915;
assign x_3539 = x_917 & x_918;
assign x_3540 = x_916 & x_3539;
assign x_3541 = x_3538 & x_3540;
assign x_3542 = x_919 & x_920;
assign x_3543 = x_922 & x_923;
assign x_3544 = x_921 & x_3543;
assign x_3545 = x_3542 & x_3544;
assign x_3546 = x_3541 & x_3545;
assign x_3547 = x_3537 & x_3546;
assign x_3548 = x_924 & x_925;
assign x_3549 = x_927 & x_928;
assign x_3550 = x_926 & x_3549;
assign x_3551 = x_3548 & x_3550;
assign x_3552 = x_929 & x_930;
assign x_3553 = x_932 & x_933;
assign x_3554 = x_931 & x_3553;
assign x_3555 = x_3552 & x_3554;
assign x_3556 = x_3551 & x_3555;
assign x_3557 = x_934 & x_935;
assign x_3558 = x_937 & x_938;
assign x_3559 = x_936 & x_3558;
assign x_3560 = x_3557 & x_3559;
assign x_3561 = x_940 & x_941;
assign x_3562 = x_939 & x_3561;
assign x_3563 = x_943 & x_944;
assign x_3564 = x_942 & x_3563;
assign x_3565 = x_3562 & x_3564;
assign x_3566 = x_3560 & x_3565;
assign x_3567 = x_3556 & x_3566;
assign x_3568 = x_3547 & x_3567;
assign x_3569 = x_945 & x_946;
assign x_3570 = x_948 & x_949;
assign x_3571 = x_947 & x_3570;
assign x_3572 = x_3569 & x_3571;
assign x_3573 = x_950 & x_951;
assign x_3574 = x_953 & x_954;
assign x_3575 = x_952 & x_3574;
assign x_3576 = x_3573 & x_3575;
assign x_3577 = x_3572 & x_3576;
assign x_3578 = x_955 & x_956;
assign x_3579 = x_958 & x_959;
assign x_3580 = x_957 & x_3579;
assign x_3581 = x_3578 & x_3580;
assign x_3582 = x_960 & x_961;
assign x_3583 = x_963 & x_964;
assign x_3584 = x_962 & x_3583;
assign x_3585 = x_3582 & x_3584;
assign x_3586 = x_3581 & x_3585;
assign x_3587 = x_3577 & x_3586;
assign x_3588 = x_965 & x_966;
assign x_3589 = x_968 & x_969;
assign x_3590 = x_967 & x_3589;
assign x_3591 = x_3588 & x_3590;
assign x_3592 = x_970 & x_971;
assign x_3593 = x_973 & x_974;
assign x_3594 = x_972 & x_3593;
assign x_3595 = x_3592 & x_3594;
assign x_3596 = x_3591 & x_3595;
assign x_3597 = x_975 & x_976;
assign x_3598 = x_978 & x_979;
assign x_3599 = x_977 & x_3598;
assign x_3600 = x_3597 & x_3599;
assign x_3601 = x_981 & x_982;
assign x_3602 = x_980 & x_3601;
assign x_3603 = x_984 & x_985;
assign x_3604 = x_983 & x_3603;
assign x_3605 = x_3602 & x_3604;
assign x_3606 = x_3600 & x_3605;
assign x_3607 = x_3596 & x_3606;
assign x_3608 = x_3587 & x_3607;
assign x_3609 = x_3568 & x_3608;
assign x_3610 = x_3528 & x_3609;
assign x_3611 = x_3447 & x_3610;
assign x_3612 = x_986 & x_987;
assign x_3613 = x_989 & x_990;
assign x_3614 = x_988 & x_3613;
assign x_3615 = x_3612 & x_3614;
assign x_3616 = x_991 & x_992;
assign x_3617 = x_994 & x_995;
assign x_3618 = x_993 & x_3617;
assign x_3619 = x_3616 & x_3618;
assign x_3620 = x_3615 & x_3619;
assign x_3621 = x_996 & x_997;
assign x_3622 = x_999 & x_1000;
assign x_3623 = x_998 & x_3622;
assign x_3624 = x_3621 & x_3623;
assign x_3625 = x_1001 & x_1002;
assign x_3626 = x_1004 & x_1005;
assign x_3627 = x_1003 & x_3626;
assign x_3628 = x_3625 & x_3627;
assign x_3629 = x_3624 & x_3628;
assign x_3630 = x_3620 & x_3629;
assign x_3631 = x_1006 & x_1007;
assign x_3632 = x_1009 & x_1010;
assign x_3633 = x_1008 & x_3632;
assign x_3634 = x_3631 & x_3633;
assign x_3635 = x_1011 & x_1012;
assign x_3636 = x_1014 & x_1015;
assign x_3637 = x_1013 & x_3636;
assign x_3638 = x_3635 & x_3637;
assign x_3639 = x_3634 & x_3638;
assign x_3640 = x_1016 & x_1017;
assign x_3641 = x_1019 & x_1020;
assign x_3642 = x_1018 & x_3641;
assign x_3643 = x_3640 & x_3642;
assign x_3644 = x_1022 & x_1023;
assign x_3645 = x_1021 & x_3644;
assign x_3646 = x_1025 & x_1026;
assign x_3647 = x_1024 & x_3646;
assign x_3648 = x_3645 & x_3647;
assign x_3649 = x_3643 & x_3648;
assign x_3650 = x_3639 & x_3649;
assign x_3651 = x_3630 & x_3650;
assign x_3652 = x_1027 & x_1028;
assign x_3653 = x_1030 & x_1031;
assign x_3654 = x_1029 & x_3653;
assign x_3655 = x_3652 & x_3654;
assign x_3656 = x_1032 & x_1033;
assign x_3657 = x_1035 & x_1036;
assign x_3658 = x_1034 & x_3657;
assign x_3659 = x_3656 & x_3658;
assign x_3660 = x_3655 & x_3659;
assign x_3661 = x_1037 & x_1038;
assign x_3662 = x_1040 & x_1041;
assign x_3663 = x_1039 & x_3662;
assign x_3664 = x_3661 & x_3663;
assign x_3665 = x_1042 & x_1043;
assign x_3666 = x_1045 & x_1046;
assign x_3667 = x_1044 & x_3666;
assign x_3668 = x_3665 & x_3667;
assign x_3669 = x_3664 & x_3668;
assign x_3670 = x_3660 & x_3669;
assign x_3671 = x_1047 & x_1048;
assign x_3672 = x_1050 & x_1051;
assign x_3673 = x_1049 & x_3672;
assign x_3674 = x_3671 & x_3673;
assign x_3675 = x_1052 & x_1053;
assign x_3676 = x_1055 & x_1056;
assign x_3677 = x_1054 & x_3676;
assign x_3678 = x_3675 & x_3677;
assign x_3679 = x_3674 & x_3678;
assign x_3680 = x_1057 & x_1058;
assign x_3681 = x_1060 & x_1061;
assign x_3682 = x_1059 & x_3681;
assign x_3683 = x_3680 & x_3682;
assign x_3684 = x_1063 & x_1064;
assign x_3685 = x_1062 & x_3684;
assign x_3686 = x_1066 & x_1067;
assign x_3687 = x_1065 & x_3686;
assign x_3688 = x_3685 & x_3687;
assign x_3689 = x_3683 & x_3688;
assign x_3690 = x_3679 & x_3689;
assign x_3691 = x_3670 & x_3690;
assign x_3692 = x_3651 & x_3691;
assign x_3693 = x_1068 & x_1069;
assign x_3694 = x_1071 & x_1072;
assign x_3695 = x_1070 & x_3694;
assign x_3696 = x_3693 & x_3695;
assign x_3697 = x_1073 & x_1074;
assign x_3698 = x_1076 & x_1077;
assign x_3699 = x_1075 & x_3698;
assign x_3700 = x_3697 & x_3699;
assign x_3701 = x_3696 & x_3700;
assign x_3702 = x_1078 & x_1079;
assign x_3703 = x_1081 & x_1082;
assign x_3704 = x_1080 & x_3703;
assign x_3705 = x_3702 & x_3704;
assign x_3706 = x_1083 & x_1084;
assign x_3707 = x_1086 & x_1087;
assign x_3708 = x_1085 & x_3707;
assign x_3709 = x_3706 & x_3708;
assign x_3710 = x_3705 & x_3709;
assign x_3711 = x_3701 & x_3710;
assign x_3712 = x_1088 & x_1089;
assign x_3713 = x_1091 & x_1092;
assign x_3714 = x_1090 & x_3713;
assign x_3715 = x_3712 & x_3714;
assign x_3716 = x_1093 & x_1094;
assign x_3717 = x_1096 & x_1097;
assign x_3718 = x_1095 & x_3717;
assign x_3719 = x_3716 & x_3718;
assign x_3720 = x_3715 & x_3719;
assign x_3721 = x_1098 & x_1099;
assign x_3722 = x_1101 & x_1102;
assign x_3723 = x_1100 & x_3722;
assign x_3724 = x_3721 & x_3723;
assign x_3725 = x_1104 & x_1105;
assign x_3726 = x_1103 & x_3725;
assign x_3727 = x_1107 & x_1108;
assign x_3728 = x_1106 & x_3727;
assign x_3729 = x_3726 & x_3728;
assign x_3730 = x_3724 & x_3729;
assign x_3731 = x_3720 & x_3730;
assign x_3732 = x_3711 & x_3731;
assign x_3733 = x_1109 & x_1110;
assign x_3734 = x_1112 & x_1113;
assign x_3735 = x_1111 & x_3734;
assign x_3736 = x_3733 & x_3735;
assign x_3737 = x_1114 & x_1115;
assign x_3738 = x_1117 & x_1118;
assign x_3739 = x_1116 & x_3738;
assign x_3740 = x_3737 & x_3739;
assign x_3741 = x_3736 & x_3740;
assign x_3742 = x_1119 & x_1120;
assign x_3743 = x_1122 & x_1123;
assign x_3744 = x_1121 & x_3743;
assign x_3745 = x_3742 & x_3744;
assign x_3746 = x_1124 & x_1125;
assign x_3747 = x_1127 & x_1128;
assign x_3748 = x_1126 & x_3747;
assign x_3749 = x_3746 & x_3748;
assign x_3750 = x_3745 & x_3749;
assign x_3751 = x_3741 & x_3750;
assign x_3752 = x_1129 & x_1130;
assign x_3753 = x_1132 & x_1133;
assign x_3754 = x_1131 & x_3753;
assign x_3755 = x_3752 & x_3754;
assign x_3756 = x_1134 & x_1135;
assign x_3757 = x_1137 & x_1138;
assign x_3758 = x_1136 & x_3757;
assign x_3759 = x_3756 & x_3758;
assign x_3760 = x_3755 & x_3759;
assign x_3761 = x_1139 & x_1140;
assign x_3762 = x_1142 & x_1143;
assign x_3763 = x_1141 & x_3762;
assign x_3764 = x_3761 & x_3763;
assign x_3765 = x_1145 & x_1146;
assign x_3766 = x_1144 & x_3765;
assign x_3767 = x_1148 & x_1149;
assign x_3768 = x_1147 & x_3767;
assign x_3769 = x_3766 & x_3768;
assign x_3770 = x_3764 & x_3769;
assign x_3771 = x_3760 & x_3770;
assign x_3772 = x_3751 & x_3771;
assign x_3773 = x_3732 & x_3772;
assign x_3774 = x_3692 & x_3773;
assign x_3775 = x_1150 & x_1151;
assign x_3776 = x_1153 & x_1154;
assign x_3777 = x_1152 & x_3776;
assign x_3778 = x_3775 & x_3777;
assign x_3779 = x_1155 & x_1156;
assign x_3780 = x_1158 & x_1159;
assign x_3781 = x_1157 & x_3780;
assign x_3782 = x_3779 & x_3781;
assign x_3783 = x_3778 & x_3782;
assign x_3784 = x_1160 & x_1161;
assign x_3785 = x_1163 & x_1164;
assign x_3786 = x_1162 & x_3785;
assign x_3787 = x_3784 & x_3786;
assign x_3788 = x_1165 & x_1166;
assign x_3789 = x_1168 & x_1169;
assign x_3790 = x_1167 & x_3789;
assign x_3791 = x_3788 & x_3790;
assign x_3792 = x_3787 & x_3791;
assign x_3793 = x_3783 & x_3792;
assign x_3794 = x_1170 & x_1171;
assign x_3795 = x_1173 & x_1174;
assign x_3796 = x_1172 & x_3795;
assign x_3797 = x_3794 & x_3796;
assign x_3798 = x_1175 & x_1176;
assign x_3799 = x_1178 & x_1179;
assign x_3800 = x_1177 & x_3799;
assign x_3801 = x_3798 & x_3800;
assign x_3802 = x_3797 & x_3801;
assign x_3803 = x_1180 & x_1181;
assign x_3804 = x_1183 & x_1184;
assign x_3805 = x_1182 & x_3804;
assign x_3806 = x_3803 & x_3805;
assign x_3807 = x_1186 & x_1187;
assign x_3808 = x_1185 & x_3807;
assign x_3809 = x_1189 & x_1190;
assign x_3810 = x_1188 & x_3809;
assign x_3811 = x_3808 & x_3810;
assign x_3812 = x_3806 & x_3811;
assign x_3813 = x_3802 & x_3812;
assign x_3814 = x_3793 & x_3813;
assign x_3815 = x_1191 & x_1192;
assign x_3816 = x_1194 & x_1195;
assign x_3817 = x_1193 & x_3816;
assign x_3818 = x_3815 & x_3817;
assign x_3819 = x_1196 & x_1197;
assign x_3820 = x_1199 & x_1200;
assign x_3821 = x_1198 & x_3820;
assign x_3822 = x_3819 & x_3821;
assign x_3823 = x_3818 & x_3822;
assign x_3824 = x_1201 & x_1202;
assign x_3825 = x_1204 & x_1205;
assign x_3826 = x_1203 & x_3825;
assign x_3827 = x_3824 & x_3826;
assign x_3828 = x_1206 & x_1207;
assign x_3829 = x_1209 & x_1210;
assign x_3830 = x_1208 & x_3829;
assign x_3831 = x_3828 & x_3830;
assign x_3832 = x_3827 & x_3831;
assign x_3833 = x_3823 & x_3832;
assign x_3834 = x_1211 & x_1212;
assign x_3835 = x_1214 & x_1215;
assign x_3836 = x_1213 & x_3835;
assign x_3837 = x_3834 & x_3836;
assign x_3838 = x_1216 & x_1217;
assign x_3839 = x_1219 & x_1220;
assign x_3840 = x_1218 & x_3839;
assign x_3841 = x_3838 & x_3840;
assign x_3842 = x_3837 & x_3841;
assign x_3843 = x_1221 & x_1222;
assign x_3844 = x_1224 & x_1225;
assign x_3845 = x_1223 & x_3844;
assign x_3846 = x_3843 & x_3845;
assign x_3847 = x_1227 & x_1228;
assign x_3848 = x_1226 & x_3847;
assign x_3849 = x_1230 & x_1231;
assign x_3850 = x_1229 & x_3849;
assign x_3851 = x_3848 & x_3850;
assign x_3852 = x_3846 & x_3851;
assign x_3853 = x_3842 & x_3852;
assign x_3854 = x_3833 & x_3853;
assign x_3855 = x_3814 & x_3854;
assign x_3856 = x_1232 & x_1233;
assign x_3857 = x_1235 & x_1236;
assign x_3858 = x_1234 & x_3857;
assign x_3859 = x_3856 & x_3858;
assign x_3860 = x_1237 & x_1238;
assign x_3861 = x_1240 & x_1241;
assign x_3862 = x_1239 & x_3861;
assign x_3863 = x_3860 & x_3862;
assign x_3864 = x_3859 & x_3863;
assign x_3865 = x_1242 & x_1243;
assign x_3866 = x_1245 & x_1246;
assign x_3867 = x_1244 & x_3866;
assign x_3868 = x_3865 & x_3867;
assign x_3869 = x_1247 & x_1248;
assign x_3870 = x_1250 & x_1251;
assign x_3871 = x_1249 & x_3870;
assign x_3872 = x_3869 & x_3871;
assign x_3873 = x_3868 & x_3872;
assign x_3874 = x_3864 & x_3873;
assign x_3875 = x_1252 & x_1253;
assign x_3876 = x_1255 & x_1256;
assign x_3877 = x_1254 & x_3876;
assign x_3878 = x_3875 & x_3877;
assign x_3879 = x_1257 & x_1258;
assign x_3880 = x_1260 & x_1261;
assign x_3881 = x_1259 & x_3880;
assign x_3882 = x_3879 & x_3881;
assign x_3883 = x_3878 & x_3882;
assign x_3884 = x_1262 & x_1263;
assign x_3885 = x_1265 & x_1266;
assign x_3886 = x_1264 & x_3885;
assign x_3887 = x_3884 & x_3886;
assign x_3888 = x_1268 & x_1269;
assign x_3889 = x_1267 & x_3888;
assign x_3890 = x_1271 & x_1272;
assign x_3891 = x_1270 & x_3890;
assign x_3892 = x_3889 & x_3891;
assign x_3893 = x_3887 & x_3892;
assign x_3894 = x_3883 & x_3893;
assign x_3895 = x_3874 & x_3894;
assign x_3896 = x_1273 & x_1274;
assign x_3897 = x_1276 & x_1277;
assign x_3898 = x_1275 & x_3897;
assign x_3899 = x_3896 & x_3898;
assign x_3900 = x_1278 & x_1279;
assign x_3901 = x_1281 & x_1282;
assign x_3902 = x_1280 & x_3901;
assign x_3903 = x_3900 & x_3902;
assign x_3904 = x_3899 & x_3903;
assign x_3905 = x_1283 & x_1284;
assign x_3906 = x_1286 & x_1287;
assign x_3907 = x_1285 & x_3906;
assign x_3908 = x_3905 & x_3907;
assign x_3909 = x_1289 & x_1290;
assign x_3910 = x_1288 & x_3909;
assign x_3911 = x_1292 & x_1293;
assign x_3912 = x_1291 & x_3911;
assign x_3913 = x_3910 & x_3912;
assign x_3914 = x_3908 & x_3913;
assign x_3915 = x_3904 & x_3914;
assign x_3916 = x_1294 & x_1295;
assign x_3917 = x_1297 & x_1298;
assign x_3918 = x_1296 & x_3917;
assign x_3919 = x_3916 & x_3918;
assign x_3920 = x_1299 & x_1300;
assign x_3921 = x_1302 & x_1303;
assign x_3922 = x_1301 & x_3921;
assign x_3923 = x_3920 & x_3922;
assign x_3924 = x_3919 & x_3923;
assign x_3925 = x_1304 & x_1305;
assign x_3926 = x_1307 & x_1308;
assign x_3927 = x_1306 & x_3926;
assign x_3928 = x_3925 & x_3927;
assign x_3929 = x_1310 & x_1311;
assign x_3930 = x_1309 & x_3929;
assign x_3931 = x_1313 & x_1314;
assign x_3932 = x_1312 & x_3931;
assign x_3933 = x_3930 & x_3932;
assign x_3934 = x_3928 & x_3933;
assign x_3935 = x_3924 & x_3934;
assign x_3936 = x_3915 & x_3935;
assign x_3937 = x_3895 & x_3936;
assign x_3938 = x_3855 & x_3937;
assign x_3939 = x_3774 & x_3938;
assign x_3940 = x_3611 & x_3939;
assign x_3941 = x_3284 & x_3940;
assign x_3942 = x_1315 & x_1316;
assign x_3943 = x_1318 & x_1319;
assign x_3944 = x_1317 & x_3943;
assign x_3945 = x_3942 & x_3944;
assign x_3946 = x_1320 & x_1321;
assign x_3947 = x_1323 & x_1324;
assign x_3948 = x_1322 & x_3947;
assign x_3949 = x_3946 & x_3948;
assign x_3950 = x_3945 & x_3949;
assign x_3951 = x_1325 & x_1326;
assign x_3952 = x_1328 & x_1329;
assign x_3953 = x_1327 & x_3952;
assign x_3954 = x_3951 & x_3953;
assign x_3955 = x_1330 & x_1331;
assign x_3956 = x_1333 & x_1334;
assign x_3957 = x_1332 & x_3956;
assign x_3958 = x_3955 & x_3957;
assign x_3959 = x_3954 & x_3958;
assign x_3960 = x_3950 & x_3959;
assign x_3961 = x_1335 & x_1336;
assign x_3962 = x_1338 & x_1339;
assign x_3963 = x_1337 & x_3962;
assign x_3964 = x_3961 & x_3963;
assign x_3965 = x_1340 & x_1341;
assign x_3966 = x_1343 & x_1344;
assign x_3967 = x_1342 & x_3966;
assign x_3968 = x_3965 & x_3967;
assign x_3969 = x_3964 & x_3968;
assign x_3970 = x_1345 & x_1346;
assign x_3971 = x_1348 & x_1349;
assign x_3972 = x_1347 & x_3971;
assign x_3973 = x_3970 & x_3972;
assign x_3974 = x_1351 & x_1352;
assign x_3975 = x_1350 & x_3974;
assign x_3976 = x_1354 & x_1355;
assign x_3977 = x_1353 & x_3976;
assign x_3978 = x_3975 & x_3977;
assign x_3979 = x_3973 & x_3978;
assign x_3980 = x_3969 & x_3979;
assign x_3981 = x_3960 & x_3980;
assign x_3982 = x_1356 & x_1357;
assign x_3983 = x_1359 & x_1360;
assign x_3984 = x_1358 & x_3983;
assign x_3985 = x_3982 & x_3984;
assign x_3986 = x_1361 & x_1362;
assign x_3987 = x_1364 & x_1365;
assign x_3988 = x_1363 & x_3987;
assign x_3989 = x_3986 & x_3988;
assign x_3990 = x_3985 & x_3989;
assign x_3991 = x_1366 & x_1367;
assign x_3992 = x_1369 & x_1370;
assign x_3993 = x_1368 & x_3992;
assign x_3994 = x_3991 & x_3993;
assign x_3995 = x_1371 & x_1372;
assign x_3996 = x_1374 & x_1375;
assign x_3997 = x_1373 & x_3996;
assign x_3998 = x_3995 & x_3997;
assign x_3999 = x_3994 & x_3998;
assign x_4000 = x_3990 & x_3999;
assign x_4001 = x_1376 & x_1377;
assign x_4002 = x_1379 & x_1380;
assign x_4003 = x_1378 & x_4002;
assign x_4004 = x_4001 & x_4003;
assign x_4005 = x_1381 & x_1382;
assign x_4006 = x_1384 & x_1385;
assign x_4007 = x_1383 & x_4006;
assign x_4008 = x_4005 & x_4007;
assign x_4009 = x_4004 & x_4008;
assign x_4010 = x_1386 & x_1387;
assign x_4011 = x_1389 & x_1390;
assign x_4012 = x_1388 & x_4011;
assign x_4013 = x_4010 & x_4012;
assign x_4014 = x_1392 & x_1393;
assign x_4015 = x_1391 & x_4014;
assign x_4016 = x_1395 & x_1396;
assign x_4017 = x_1394 & x_4016;
assign x_4018 = x_4015 & x_4017;
assign x_4019 = x_4013 & x_4018;
assign x_4020 = x_4009 & x_4019;
assign x_4021 = x_4000 & x_4020;
assign x_4022 = x_3981 & x_4021;
assign x_4023 = x_1397 & x_1398;
assign x_4024 = x_1400 & x_1401;
assign x_4025 = x_1399 & x_4024;
assign x_4026 = x_4023 & x_4025;
assign x_4027 = x_1402 & x_1403;
assign x_4028 = x_1405 & x_1406;
assign x_4029 = x_1404 & x_4028;
assign x_4030 = x_4027 & x_4029;
assign x_4031 = x_4026 & x_4030;
assign x_4032 = x_1407 & x_1408;
assign x_4033 = x_1410 & x_1411;
assign x_4034 = x_1409 & x_4033;
assign x_4035 = x_4032 & x_4034;
assign x_4036 = x_1412 & x_1413;
assign x_4037 = x_1415 & x_1416;
assign x_4038 = x_1414 & x_4037;
assign x_4039 = x_4036 & x_4038;
assign x_4040 = x_4035 & x_4039;
assign x_4041 = x_4031 & x_4040;
assign x_4042 = x_1417 & x_1418;
assign x_4043 = x_1420 & x_1421;
assign x_4044 = x_1419 & x_4043;
assign x_4045 = x_4042 & x_4044;
assign x_4046 = x_1422 & x_1423;
assign x_4047 = x_1425 & x_1426;
assign x_4048 = x_1424 & x_4047;
assign x_4049 = x_4046 & x_4048;
assign x_4050 = x_4045 & x_4049;
assign x_4051 = x_1427 & x_1428;
assign x_4052 = x_1430 & x_1431;
assign x_4053 = x_1429 & x_4052;
assign x_4054 = x_4051 & x_4053;
assign x_4055 = x_1433 & x_1434;
assign x_4056 = x_1432 & x_4055;
assign x_4057 = x_1436 & x_1437;
assign x_4058 = x_1435 & x_4057;
assign x_4059 = x_4056 & x_4058;
assign x_4060 = x_4054 & x_4059;
assign x_4061 = x_4050 & x_4060;
assign x_4062 = x_4041 & x_4061;
assign x_4063 = x_1438 & x_1439;
assign x_4064 = x_1441 & x_1442;
assign x_4065 = x_1440 & x_4064;
assign x_4066 = x_4063 & x_4065;
assign x_4067 = x_1443 & x_1444;
assign x_4068 = x_1446 & x_1447;
assign x_4069 = x_1445 & x_4068;
assign x_4070 = x_4067 & x_4069;
assign x_4071 = x_4066 & x_4070;
assign x_4072 = x_1448 & x_1449;
assign x_4073 = x_1451 & x_1452;
assign x_4074 = x_1450 & x_4073;
assign x_4075 = x_4072 & x_4074;
assign x_4076 = x_1453 & x_1454;
assign x_4077 = x_1456 & x_1457;
assign x_4078 = x_1455 & x_4077;
assign x_4079 = x_4076 & x_4078;
assign x_4080 = x_4075 & x_4079;
assign x_4081 = x_4071 & x_4080;
assign x_4082 = x_1458 & x_1459;
assign x_4083 = x_1461 & x_1462;
assign x_4084 = x_1460 & x_4083;
assign x_4085 = x_4082 & x_4084;
assign x_4086 = x_1463 & x_1464;
assign x_4087 = x_1466 & x_1467;
assign x_4088 = x_1465 & x_4087;
assign x_4089 = x_4086 & x_4088;
assign x_4090 = x_4085 & x_4089;
assign x_4091 = x_1468 & x_1469;
assign x_4092 = x_1471 & x_1472;
assign x_4093 = x_1470 & x_4092;
assign x_4094 = x_4091 & x_4093;
assign x_4095 = x_1474 & x_1475;
assign x_4096 = x_1473 & x_4095;
assign x_4097 = x_1477 & x_1478;
assign x_4098 = x_1476 & x_4097;
assign x_4099 = x_4096 & x_4098;
assign x_4100 = x_4094 & x_4099;
assign x_4101 = x_4090 & x_4100;
assign x_4102 = x_4081 & x_4101;
assign x_4103 = x_4062 & x_4102;
assign x_4104 = x_4022 & x_4103;
assign x_4105 = x_1479 & x_1480;
assign x_4106 = x_1482 & x_1483;
assign x_4107 = x_1481 & x_4106;
assign x_4108 = x_4105 & x_4107;
assign x_4109 = x_1484 & x_1485;
assign x_4110 = x_1487 & x_1488;
assign x_4111 = x_1486 & x_4110;
assign x_4112 = x_4109 & x_4111;
assign x_4113 = x_4108 & x_4112;
assign x_4114 = x_1489 & x_1490;
assign x_4115 = x_1492 & x_1493;
assign x_4116 = x_1491 & x_4115;
assign x_4117 = x_4114 & x_4116;
assign x_4118 = x_1494 & x_1495;
assign x_4119 = x_1497 & x_1498;
assign x_4120 = x_1496 & x_4119;
assign x_4121 = x_4118 & x_4120;
assign x_4122 = x_4117 & x_4121;
assign x_4123 = x_4113 & x_4122;
assign x_4124 = x_1499 & x_1500;
assign x_4125 = x_1502 & x_1503;
assign x_4126 = x_1501 & x_4125;
assign x_4127 = x_4124 & x_4126;
assign x_4128 = x_1504 & x_1505;
assign x_4129 = x_1507 & x_1508;
assign x_4130 = x_1506 & x_4129;
assign x_4131 = x_4128 & x_4130;
assign x_4132 = x_4127 & x_4131;
assign x_4133 = x_1509 & x_1510;
assign x_4134 = x_1512 & x_1513;
assign x_4135 = x_1511 & x_4134;
assign x_4136 = x_4133 & x_4135;
assign x_4137 = x_1515 & x_1516;
assign x_4138 = x_1514 & x_4137;
assign x_4139 = x_1518 & x_1519;
assign x_4140 = x_1517 & x_4139;
assign x_4141 = x_4138 & x_4140;
assign x_4142 = x_4136 & x_4141;
assign x_4143 = x_4132 & x_4142;
assign x_4144 = x_4123 & x_4143;
assign x_4145 = x_1520 & x_1521;
assign x_4146 = x_1523 & x_1524;
assign x_4147 = x_1522 & x_4146;
assign x_4148 = x_4145 & x_4147;
assign x_4149 = x_1525 & x_1526;
assign x_4150 = x_1528 & x_1529;
assign x_4151 = x_1527 & x_4150;
assign x_4152 = x_4149 & x_4151;
assign x_4153 = x_4148 & x_4152;
assign x_4154 = x_1530 & x_1531;
assign x_4155 = x_1533 & x_1534;
assign x_4156 = x_1532 & x_4155;
assign x_4157 = x_4154 & x_4156;
assign x_4158 = x_1535 & x_1536;
assign x_4159 = x_1538 & x_1539;
assign x_4160 = x_1537 & x_4159;
assign x_4161 = x_4158 & x_4160;
assign x_4162 = x_4157 & x_4161;
assign x_4163 = x_4153 & x_4162;
assign x_4164 = x_1540 & x_1541;
assign x_4165 = x_1543 & x_1544;
assign x_4166 = x_1542 & x_4165;
assign x_4167 = x_4164 & x_4166;
assign x_4168 = x_1545 & x_1546;
assign x_4169 = x_1548 & x_1549;
assign x_4170 = x_1547 & x_4169;
assign x_4171 = x_4168 & x_4170;
assign x_4172 = x_4167 & x_4171;
assign x_4173 = x_1550 & x_1551;
assign x_4174 = x_1553 & x_1554;
assign x_4175 = x_1552 & x_4174;
assign x_4176 = x_4173 & x_4175;
assign x_4177 = x_1556 & x_1557;
assign x_4178 = x_1555 & x_4177;
assign x_4179 = x_1559 & x_1560;
assign x_4180 = x_1558 & x_4179;
assign x_4181 = x_4178 & x_4180;
assign x_4182 = x_4176 & x_4181;
assign x_4183 = x_4172 & x_4182;
assign x_4184 = x_4163 & x_4183;
assign x_4185 = x_4144 & x_4184;
assign x_4186 = x_1561 & x_1562;
assign x_4187 = x_1564 & x_1565;
assign x_4188 = x_1563 & x_4187;
assign x_4189 = x_4186 & x_4188;
assign x_4190 = x_1566 & x_1567;
assign x_4191 = x_1569 & x_1570;
assign x_4192 = x_1568 & x_4191;
assign x_4193 = x_4190 & x_4192;
assign x_4194 = x_4189 & x_4193;
assign x_4195 = x_1571 & x_1572;
assign x_4196 = x_1574 & x_1575;
assign x_4197 = x_1573 & x_4196;
assign x_4198 = x_4195 & x_4197;
assign x_4199 = x_1576 & x_1577;
assign x_4200 = x_1579 & x_1580;
assign x_4201 = x_1578 & x_4200;
assign x_4202 = x_4199 & x_4201;
assign x_4203 = x_4198 & x_4202;
assign x_4204 = x_4194 & x_4203;
assign x_4205 = x_1581 & x_1582;
assign x_4206 = x_1584 & x_1585;
assign x_4207 = x_1583 & x_4206;
assign x_4208 = x_4205 & x_4207;
assign x_4209 = x_1586 & x_1587;
assign x_4210 = x_1589 & x_1590;
assign x_4211 = x_1588 & x_4210;
assign x_4212 = x_4209 & x_4211;
assign x_4213 = x_4208 & x_4212;
assign x_4214 = x_1591 & x_1592;
assign x_4215 = x_1594 & x_1595;
assign x_4216 = x_1593 & x_4215;
assign x_4217 = x_4214 & x_4216;
assign x_4218 = x_1597 & x_1598;
assign x_4219 = x_1596 & x_4218;
assign x_4220 = x_1600 & x_1601;
assign x_4221 = x_1599 & x_4220;
assign x_4222 = x_4219 & x_4221;
assign x_4223 = x_4217 & x_4222;
assign x_4224 = x_4213 & x_4223;
assign x_4225 = x_4204 & x_4224;
assign x_4226 = x_1602 & x_1603;
assign x_4227 = x_1605 & x_1606;
assign x_4228 = x_1604 & x_4227;
assign x_4229 = x_4226 & x_4228;
assign x_4230 = x_1607 & x_1608;
assign x_4231 = x_1610 & x_1611;
assign x_4232 = x_1609 & x_4231;
assign x_4233 = x_4230 & x_4232;
assign x_4234 = x_4229 & x_4233;
assign x_4235 = x_1612 & x_1613;
assign x_4236 = x_1615 & x_1616;
assign x_4237 = x_1614 & x_4236;
assign x_4238 = x_4235 & x_4237;
assign x_4239 = x_1617 & x_1618;
assign x_4240 = x_1620 & x_1621;
assign x_4241 = x_1619 & x_4240;
assign x_4242 = x_4239 & x_4241;
assign x_4243 = x_4238 & x_4242;
assign x_4244 = x_4234 & x_4243;
assign x_4245 = x_1622 & x_1623;
assign x_4246 = x_1625 & x_1626;
assign x_4247 = x_1624 & x_4246;
assign x_4248 = x_4245 & x_4247;
assign x_4249 = x_1627 & x_1628;
assign x_4250 = x_1630 & x_1631;
assign x_4251 = x_1629 & x_4250;
assign x_4252 = x_4249 & x_4251;
assign x_4253 = x_4248 & x_4252;
assign x_4254 = x_1632 & x_1633;
assign x_4255 = x_1635 & x_1636;
assign x_4256 = x_1634 & x_4255;
assign x_4257 = x_4254 & x_4256;
assign x_4258 = x_1638 & x_1639;
assign x_4259 = x_1637 & x_4258;
assign x_4260 = x_1641 & x_1642;
assign x_4261 = x_1640 & x_4260;
assign x_4262 = x_4259 & x_4261;
assign x_4263 = x_4257 & x_4262;
assign x_4264 = x_4253 & x_4263;
assign x_4265 = x_4244 & x_4264;
assign x_4266 = x_4225 & x_4265;
assign x_4267 = x_4185 & x_4266;
assign x_4268 = x_4104 & x_4267;
assign x_4269 = x_1643 & x_1644;
assign x_4270 = x_1646 & x_1647;
assign x_4271 = x_1645 & x_4270;
assign x_4272 = x_4269 & x_4271;
assign x_4273 = x_1648 & x_1649;
assign x_4274 = x_1651 & x_1652;
assign x_4275 = x_1650 & x_4274;
assign x_4276 = x_4273 & x_4275;
assign x_4277 = x_4272 & x_4276;
assign x_4278 = x_1653 & x_1654;
assign x_4279 = x_1656 & x_1657;
assign x_4280 = x_1655 & x_4279;
assign x_4281 = x_4278 & x_4280;
assign x_4282 = x_1658 & x_1659;
assign x_4283 = x_1661 & x_1662;
assign x_4284 = x_1660 & x_4283;
assign x_4285 = x_4282 & x_4284;
assign x_4286 = x_4281 & x_4285;
assign x_4287 = x_4277 & x_4286;
assign x_4288 = x_1663 & x_1664;
assign x_4289 = x_1666 & x_1667;
assign x_4290 = x_1665 & x_4289;
assign x_4291 = x_4288 & x_4290;
assign x_4292 = x_1668 & x_1669;
assign x_4293 = x_1671 & x_1672;
assign x_4294 = x_1670 & x_4293;
assign x_4295 = x_4292 & x_4294;
assign x_4296 = x_4291 & x_4295;
assign x_4297 = x_1673 & x_1674;
assign x_4298 = x_1676 & x_1677;
assign x_4299 = x_1675 & x_4298;
assign x_4300 = x_4297 & x_4299;
assign x_4301 = x_1679 & x_1680;
assign x_4302 = x_1678 & x_4301;
assign x_4303 = x_1682 & x_1683;
assign x_4304 = x_1681 & x_4303;
assign x_4305 = x_4302 & x_4304;
assign x_4306 = x_4300 & x_4305;
assign x_4307 = x_4296 & x_4306;
assign x_4308 = x_4287 & x_4307;
assign x_4309 = x_1684 & x_1685;
assign x_4310 = x_1687 & x_1688;
assign x_4311 = x_1686 & x_4310;
assign x_4312 = x_4309 & x_4311;
assign x_4313 = x_1689 & x_1690;
assign x_4314 = x_1692 & x_1693;
assign x_4315 = x_1691 & x_4314;
assign x_4316 = x_4313 & x_4315;
assign x_4317 = x_4312 & x_4316;
assign x_4318 = x_1694 & x_1695;
assign x_4319 = x_1697 & x_1698;
assign x_4320 = x_1696 & x_4319;
assign x_4321 = x_4318 & x_4320;
assign x_4322 = x_1699 & x_1700;
assign x_4323 = x_1702 & x_1703;
assign x_4324 = x_1701 & x_4323;
assign x_4325 = x_4322 & x_4324;
assign x_4326 = x_4321 & x_4325;
assign x_4327 = x_4317 & x_4326;
assign x_4328 = x_1704 & x_1705;
assign x_4329 = x_1707 & x_1708;
assign x_4330 = x_1706 & x_4329;
assign x_4331 = x_4328 & x_4330;
assign x_4332 = x_1709 & x_1710;
assign x_4333 = x_1712 & x_1713;
assign x_4334 = x_1711 & x_4333;
assign x_4335 = x_4332 & x_4334;
assign x_4336 = x_4331 & x_4335;
assign x_4337 = x_1714 & x_1715;
assign x_4338 = x_1717 & x_1718;
assign x_4339 = x_1716 & x_4338;
assign x_4340 = x_4337 & x_4339;
assign x_4341 = x_1720 & x_1721;
assign x_4342 = x_1719 & x_4341;
assign x_4343 = x_1723 & x_1724;
assign x_4344 = x_1722 & x_4343;
assign x_4345 = x_4342 & x_4344;
assign x_4346 = x_4340 & x_4345;
assign x_4347 = x_4336 & x_4346;
assign x_4348 = x_4327 & x_4347;
assign x_4349 = x_4308 & x_4348;
assign x_4350 = x_1725 & x_1726;
assign x_4351 = x_1728 & x_1729;
assign x_4352 = x_1727 & x_4351;
assign x_4353 = x_4350 & x_4352;
assign x_4354 = x_1730 & x_1731;
assign x_4355 = x_1733 & x_1734;
assign x_4356 = x_1732 & x_4355;
assign x_4357 = x_4354 & x_4356;
assign x_4358 = x_4353 & x_4357;
assign x_4359 = x_1735 & x_1736;
assign x_4360 = x_1738 & x_1739;
assign x_4361 = x_1737 & x_4360;
assign x_4362 = x_4359 & x_4361;
assign x_4363 = x_1740 & x_1741;
assign x_4364 = x_1743 & x_1744;
assign x_4365 = x_1742 & x_4364;
assign x_4366 = x_4363 & x_4365;
assign x_4367 = x_4362 & x_4366;
assign x_4368 = x_4358 & x_4367;
assign x_4369 = x_1745 & x_1746;
assign x_4370 = x_1748 & x_1749;
assign x_4371 = x_1747 & x_4370;
assign x_4372 = x_4369 & x_4371;
assign x_4373 = x_1750 & x_1751;
assign x_4374 = x_1753 & x_1754;
assign x_4375 = x_1752 & x_4374;
assign x_4376 = x_4373 & x_4375;
assign x_4377 = x_4372 & x_4376;
assign x_4378 = x_1755 & x_1756;
assign x_4379 = x_1758 & x_1759;
assign x_4380 = x_1757 & x_4379;
assign x_4381 = x_4378 & x_4380;
assign x_4382 = x_1761 & x_1762;
assign x_4383 = x_1760 & x_4382;
assign x_4384 = x_1764 & x_1765;
assign x_4385 = x_1763 & x_4384;
assign x_4386 = x_4383 & x_4385;
assign x_4387 = x_4381 & x_4386;
assign x_4388 = x_4377 & x_4387;
assign x_4389 = x_4368 & x_4388;
assign x_4390 = x_1766 & x_1767;
assign x_4391 = x_1769 & x_1770;
assign x_4392 = x_1768 & x_4391;
assign x_4393 = x_4390 & x_4392;
assign x_4394 = x_1771 & x_1772;
assign x_4395 = x_1774 & x_1775;
assign x_4396 = x_1773 & x_4395;
assign x_4397 = x_4394 & x_4396;
assign x_4398 = x_4393 & x_4397;
assign x_4399 = x_1776 & x_1777;
assign x_4400 = x_1779 & x_1780;
assign x_4401 = x_1778 & x_4400;
assign x_4402 = x_4399 & x_4401;
assign x_4403 = x_1781 & x_1782;
assign x_4404 = x_1784 & x_1785;
assign x_4405 = x_1783 & x_4404;
assign x_4406 = x_4403 & x_4405;
assign x_4407 = x_4402 & x_4406;
assign x_4408 = x_4398 & x_4407;
assign x_4409 = x_1786 & x_1787;
assign x_4410 = x_1789 & x_1790;
assign x_4411 = x_1788 & x_4410;
assign x_4412 = x_4409 & x_4411;
assign x_4413 = x_1791 & x_1792;
assign x_4414 = x_1794 & x_1795;
assign x_4415 = x_1793 & x_4414;
assign x_4416 = x_4413 & x_4415;
assign x_4417 = x_4412 & x_4416;
assign x_4418 = x_1796 & x_1797;
assign x_4419 = x_1799 & x_1800;
assign x_4420 = x_1798 & x_4419;
assign x_4421 = x_4418 & x_4420;
assign x_4422 = x_1802 & x_1803;
assign x_4423 = x_1801 & x_4422;
assign x_4424 = x_1805 & x_1806;
assign x_4425 = x_1804 & x_4424;
assign x_4426 = x_4423 & x_4425;
assign x_4427 = x_4421 & x_4426;
assign x_4428 = x_4417 & x_4427;
assign x_4429 = x_4408 & x_4428;
assign x_4430 = x_4389 & x_4429;
assign x_4431 = x_4349 & x_4430;
assign x_4432 = x_1807 & x_1808;
assign x_4433 = x_1810 & x_1811;
assign x_4434 = x_1809 & x_4433;
assign x_4435 = x_4432 & x_4434;
assign x_4436 = x_1812 & x_1813;
assign x_4437 = x_1815 & x_1816;
assign x_4438 = x_1814 & x_4437;
assign x_4439 = x_4436 & x_4438;
assign x_4440 = x_4435 & x_4439;
assign x_4441 = x_1817 & x_1818;
assign x_4442 = x_1820 & x_1821;
assign x_4443 = x_1819 & x_4442;
assign x_4444 = x_4441 & x_4443;
assign x_4445 = x_1822 & x_1823;
assign x_4446 = x_1825 & x_1826;
assign x_4447 = x_1824 & x_4446;
assign x_4448 = x_4445 & x_4447;
assign x_4449 = x_4444 & x_4448;
assign x_4450 = x_4440 & x_4449;
assign x_4451 = x_1827 & x_1828;
assign x_4452 = x_1830 & x_1831;
assign x_4453 = x_1829 & x_4452;
assign x_4454 = x_4451 & x_4453;
assign x_4455 = x_1832 & x_1833;
assign x_4456 = x_1835 & x_1836;
assign x_4457 = x_1834 & x_4456;
assign x_4458 = x_4455 & x_4457;
assign x_4459 = x_4454 & x_4458;
assign x_4460 = x_1837 & x_1838;
assign x_4461 = x_1840 & x_1841;
assign x_4462 = x_1839 & x_4461;
assign x_4463 = x_4460 & x_4462;
assign x_4464 = x_1843 & x_1844;
assign x_4465 = x_1842 & x_4464;
assign x_4466 = x_1846 & x_1847;
assign x_4467 = x_1845 & x_4466;
assign x_4468 = x_4465 & x_4467;
assign x_4469 = x_4463 & x_4468;
assign x_4470 = x_4459 & x_4469;
assign x_4471 = x_4450 & x_4470;
assign x_4472 = x_1848 & x_1849;
assign x_4473 = x_1851 & x_1852;
assign x_4474 = x_1850 & x_4473;
assign x_4475 = x_4472 & x_4474;
assign x_4476 = x_1853 & x_1854;
assign x_4477 = x_1856 & x_1857;
assign x_4478 = x_1855 & x_4477;
assign x_4479 = x_4476 & x_4478;
assign x_4480 = x_4475 & x_4479;
assign x_4481 = x_1858 & x_1859;
assign x_4482 = x_1861 & x_1862;
assign x_4483 = x_1860 & x_4482;
assign x_4484 = x_4481 & x_4483;
assign x_4485 = x_1863 & x_1864;
assign x_4486 = x_1866 & x_1867;
assign x_4487 = x_1865 & x_4486;
assign x_4488 = x_4485 & x_4487;
assign x_4489 = x_4484 & x_4488;
assign x_4490 = x_4480 & x_4489;
assign x_4491 = x_1868 & x_1869;
assign x_4492 = x_1871 & x_1872;
assign x_4493 = x_1870 & x_4492;
assign x_4494 = x_4491 & x_4493;
assign x_4495 = x_1873 & x_1874;
assign x_4496 = x_1876 & x_1877;
assign x_4497 = x_1875 & x_4496;
assign x_4498 = x_4495 & x_4497;
assign x_4499 = x_4494 & x_4498;
assign x_4500 = x_1878 & x_1879;
assign x_4501 = x_1881 & x_1882;
assign x_4502 = x_1880 & x_4501;
assign x_4503 = x_4500 & x_4502;
assign x_4504 = x_1884 & x_1885;
assign x_4505 = x_1883 & x_4504;
assign x_4506 = x_1887 & x_1888;
assign x_4507 = x_1886 & x_4506;
assign x_4508 = x_4505 & x_4507;
assign x_4509 = x_4503 & x_4508;
assign x_4510 = x_4499 & x_4509;
assign x_4511 = x_4490 & x_4510;
assign x_4512 = x_4471 & x_4511;
assign x_4513 = x_1889 & x_1890;
assign x_4514 = x_1892 & x_1893;
assign x_4515 = x_1891 & x_4514;
assign x_4516 = x_4513 & x_4515;
assign x_4517 = x_1894 & x_1895;
assign x_4518 = x_1897 & x_1898;
assign x_4519 = x_1896 & x_4518;
assign x_4520 = x_4517 & x_4519;
assign x_4521 = x_4516 & x_4520;
assign x_4522 = x_1899 & x_1900;
assign x_4523 = x_1902 & x_1903;
assign x_4524 = x_1901 & x_4523;
assign x_4525 = x_4522 & x_4524;
assign x_4526 = x_1904 & x_1905;
assign x_4527 = x_1907 & x_1908;
assign x_4528 = x_1906 & x_4527;
assign x_4529 = x_4526 & x_4528;
assign x_4530 = x_4525 & x_4529;
assign x_4531 = x_4521 & x_4530;
assign x_4532 = x_1909 & x_1910;
assign x_4533 = x_1912 & x_1913;
assign x_4534 = x_1911 & x_4533;
assign x_4535 = x_4532 & x_4534;
assign x_4536 = x_1914 & x_1915;
assign x_4537 = x_1917 & x_1918;
assign x_4538 = x_1916 & x_4537;
assign x_4539 = x_4536 & x_4538;
assign x_4540 = x_4535 & x_4539;
assign x_4541 = x_1919 & x_1920;
assign x_4542 = x_1922 & x_1923;
assign x_4543 = x_1921 & x_4542;
assign x_4544 = x_4541 & x_4543;
assign x_4545 = x_1925 & x_1926;
assign x_4546 = x_1924 & x_4545;
assign x_4547 = x_1928 & x_1929;
assign x_4548 = x_1927 & x_4547;
assign x_4549 = x_4546 & x_4548;
assign x_4550 = x_4544 & x_4549;
assign x_4551 = x_4540 & x_4550;
assign x_4552 = x_4531 & x_4551;
assign x_4553 = x_1930 & x_1931;
assign x_4554 = x_1933 & x_1934;
assign x_4555 = x_1932 & x_4554;
assign x_4556 = x_4553 & x_4555;
assign x_4557 = x_1935 & x_1936;
assign x_4558 = x_1938 & x_1939;
assign x_4559 = x_1937 & x_4558;
assign x_4560 = x_4557 & x_4559;
assign x_4561 = x_4556 & x_4560;
assign x_4562 = x_1940 & x_1941;
assign x_4563 = x_1943 & x_1944;
assign x_4564 = x_1942 & x_4563;
assign x_4565 = x_4562 & x_4564;
assign x_4566 = x_1946 & x_1947;
assign x_4567 = x_1945 & x_4566;
assign x_4568 = x_1949 & x_1950;
assign x_4569 = x_1948 & x_4568;
assign x_4570 = x_4567 & x_4569;
assign x_4571 = x_4565 & x_4570;
assign x_4572 = x_4561 & x_4571;
assign x_4573 = x_1951 & x_1952;
assign x_4574 = x_1954 & x_1955;
assign x_4575 = x_1953 & x_4574;
assign x_4576 = x_4573 & x_4575;
assign x_4577 = x_1956 & x_1957;
assign x_4578 = x_1959 & x_1960;
assign x_4579 = x_1958 & x_4578;
assign x_4580 = x_4577 & x_4579;
assign x_4581 = x_4576 & x_4580;
assign x_4582 = x_1961 & x_1962;
assign x_4583 = x_1964 & x_1965;
assign x_4584 = x_1963 & x_4583;
assign x_4585 = x_4582 & x_4584;
assign x_4586 = x_1967 & x_1968;
assign x_4587 = x_1966 & x_4586;
assign x_4588 = x_1970 & x_1971;
assign x_4589 = x_1969 & x_4588;
assign x_4590 = x_4587 & x_4589;
assign x_4591 = x_4585 & x_4590;
assign x_4592 = x_4581 & x_4591;
assign x_4593 = x_4572 & x_4592;
assign x_4594 = x_4552 & x_4593;
assign x_4595 = x_4512 & x_4594;
assign x_4596 = x_4431 & x_4595;
assign x_4597 = x_4268 & x_4596;
assign x_4598 = x_1972 & x_1973;
assign x_4599 = x_1975 & x_1976;
assign x_4600 = x_1974 & x_4599;
assign x_4601 = x_4598 & x_4600;
assign x_4602 = x_1977 & x_1978;
assign x_4603 = x_1980 & x_1981;
assign x_4604 = x_1979 & x_4603;
assign x_4605 = x_4602 & x_4604;
assign x_4606 = x_4601 & x_4605;
assign x_4607 = x_1982 & x_1983;
assign x_4608 = x_1985 & x_1986;
assign x_4609 = x_1984 & x_4608;
assign x_4610 = x_4607 & x_4609;
assign x_4611 = x_1987 & x_1988;
assign x_4612 = x_1990 & x_1991;
assign x_4613 = x_1989 & x_4612;
assign x_4614 = x_4611 & x_4613;
assign x_4615 = x_4610 & x_4614;
assign x_4616 = x_4606 & x_4615;
assign x_4617 = x_1992 & x_1993;
assign x_4618 = x_1995 & x_1996;
assign x_4619 = x_1994 & x_4618;
assign x_4620 = x_4617 & x_4619;
assign x_4621 = x_1997 & x_1998;
assign x_4622 = x_2000 & x_2001;
assign x_4623 = x_1999 & x_4622;
assign x_4624 = x_4621 & x_4623;
assign x_4625 = x_4620 & x_4624;
assign x_4626 = x_2002 & x_2003;
assign x_4627 = x_2005 & x_2006;
assign x_4628 = x_2004 & x_4627;
assign x_4629 = x_4626 & x_4628;
assign x_4630 = x_2008 & x_2009;
assign x_4631 = x_2007 & x_4630;
assign x_4632 = x_2011 & x_2012;
assign x_4633 = x_2010 & x_4632;
assign x_4634 = x_4631 & x_4633;
assign x_4635 = x_4629 & x_4634;
assign x_4636 = x_4625 & x_4635;
assign x_4637 = x_4616 & x_4636;
assign x_4638 = x_2013 & x_2014;
assign x_4639 = x_2016 & x_2017;
assign x_4640 = x_2015 & x_4639;
assign x_4641 = x_4638 & x_4640;
assign x_4642 = x_2018 & x_2019;
assign x_4643 = x_2021 & x_2022;
assign x_4644 = x_2020 & x_4643;
assign x_4645 = x_4642 & x_4644;
assign x_4646 = x_4641 & x_4645;
assign x_4647 = x_2023 & x_2024;
assign x_4648 = x_2026 & x_2027;
assign x_4649 = x_2025 & x_4648;
assign x_4650 = x_4647 & x_4649;
assign x_4651 = x_2028 & x_2029;
assign x_4652 = x_2031 & x_2032;
assign x_4653 = x_2030 & x_4652;
assign x_4654 = x_4651 & x_4653;
assign x_4655 = x_4650 & x_4654;
assign x_4656 = x_4646 & x_4655;
assign x_4657 = x_2033 & x_2034;
assign x_4658 = x_2036 & x_2037;
assign x_4659 = x_2035 & x_4658;
assign x_4660 = x_4657 & x_4659;
assign x_4661 = x_2038 & x_2039;
assign x_4662 = x_2041 & x_2042;
assign x_4663 = x_2040 & x_4662;
assign x_4664 = x_4661 & x_4663;
assign x_4665 = x_4660 & x_4664;
assign x_4666 = x_2043 & x_2044;
assign x_4667 = x_2046 & x_2047;
assign x_4668 = x_2045 & x_4667;
assign x_4669 = x_4666 & x_4668;
assign x_4670 = x_2049 & x_2050;
assign x_4671 = x_2048 & x_4670;
assign x_4672 = x_2052 & x_2053;
assign x_4673 = x_2051 & x_4672;
assign x_4674 = x_4671 & x_4673;
assign x_4675 = x_4669 & x_4674;
assign x_4676 = x_4665 & x_4675;
assign x_4677 = x_4656 & x_4676;
assign x_4678 = x_4637 & x_4677;
assign x_4679 = x_2054 & x_2055;
assign x_4680 = x_2057 & x_2058;
assign x_4681 = x_2056 & x_4680;
assign x_4682 = x_4679 & x_4681;
assign x_4683 = x_2059 & x_2060;
assign x_4684 = x_2062 & x_2063;
assign x_4685 = x_2061 & x_4684;
assign x_4686 = x_4683 & x_4685;
assign x_4687 = x_4682 & x_4686;
assign x_4688 = x_2064 & x_2065;
assign x_4689 = x_2067 & x_2068;
assign x_4690 = x_2066 & x_4689;
assign x_4691 = x_4688 & x_4690;
assign x_4692 = x_2069 & x_2070;
assign x_4693 = x_2072 & x_2073;
assign x_4694 = x_2071 & x_4693;
assign x_4695 = x_4692 & x_4694;
assign x_4696 = x_4691 & x_4695;
assign x_4697 = x_4687 & x_4696;
assign x_4698 = x_2074 & x_2075;
assign x_4699 = x_2077 & x_2078;
assign x_4700 = x_2076 & x_4699;
assign x_4701 = x_4698 & x_4700;
assign x_4702 = x_2079 & x_2080;
assign x_4703 = x_2082 & x_2083;
assign x_4704 = x_2081 & x_4703;
assign x_4705 = x_4702 & x_4704;
assign x_4706 = x_4701 & x_4705;
assign x_4707 = x_2084 & x_2085;
assign x_4708 = x_2087 & x_2088;
assign x_4709 = x_2086 & x_4708;
assign x_4710 = x_4707 & x_4709;
assign x_4711 = x_2090 & x_2091;
assign x_4712 = x_2089 & x_4711;
assign x_4713 = x_2093 & x_2094;
assign x_4714 = x_2092 & x_4713;
assign x_4715 = x_4712 & x_4714;
assign x_4716 = x_4710 & x_4715;
assign x_4717 = x_4706 & x_4716;
assign x_4718 = x_4697 & x_4717;
assign x_4719 = x_2095 & x_2096;
assign x_4720 = x_2098 & x_2099;
assign x_4721 = x_2097 & x_4720;
assign x_4722 = x_4719 & x_4721;
assign x_4723 = x_2100 & x_2101;
assign x_4724 = x_2103 & x_2104;
assign x_4725 = x_2102 & x_4724;
assign x_4726 = x_4723 & x_4725;
assign x_4727 = x_4722 & x_4726;
assign x_4728 = x_2105 & x_2106;
assign x_4729 = x_2108 & x_2109;
assign x_4730 = x_2107 & x_4729;
assign x_4731 = x_4728 & x_4730;
assign x_4732 = x_2110 & x_2111;
assign x_4733 = x_2113 & x_2114;
assign x_4734 = x_2112 & x_4733;
assign x_4735 = x_4732 & x_4734;
assign x_4736 = x_4731 & x_4735;
assign x_4737 = x_4727 & x_4736;
assign x_4738 = x_2115 & x_2116;
assign x_4739 = x_2118 & x_2119;
assign x_4740 = x_2117 & x_4739;
assign x_4741 = x_4738 & x_4740;
assign x_4742 = x_2120 & x_2121;
assign x_4743 = x_2123 & x_2124;
assign x_4744 = x_2122 & x_4743;
assign x_4745 = x_4742 & x_4744;
assign x_4746 = x_4741 & x_4745;
assign x_4747 = x_2125 & x_2126;
assign x_4748 = x_2128 & x_2129;
assign x_4749 = x_2127 & x_4748;
assign x_4750 = x_4747 & x_4749;
assign x_4751 = x_2131 & x_2132;
assign x_4752 = x_2130 & x_4751;
assign x_4753 = x_2134 & x_2135;
assign x_4754 = x_2133 & x_4753;
assign x_4755 = x_4752 & x_4754;
assign x_4756 = x_4750 & x_4755;
assign x_4757 = x_4746 & x_4756;
assign x_4758 = x_4737 & x_4757;
assign x_4759 = x_4718 & x_4758;
assign x_4760 = x_4678 & x_4759;
assign x_4761 = x_2136 & x_2137;
assign x_4762 = x_2139 & x_2140;
assign x_4763 = x_2138 & x_4762;
assign x_4764 = x_4761 & x_4763;
assign x_4765 = x_2141 & x_2142;
assign x_4766 = x_2144 & x_2145;
assign x_4767 = x_2143 & x_4766;
assign x_4768 = x_4765 & x_4767;
assign x_4769 = x_4764 & x_4768;
assign x_4770 = x_2146 & x_2147;
assign x_4771 = x_2149 & x_2150;
assign x_4772 = x_2148 & x_4771;
assign x_4773 = x_4770 & x_4772;
assign x_4774 = x_2151 & x_2152;
assign x_4775 = x_2154 & x_2155;
assign x_4776 = x_2153 & x_4775;
assign x_4777 = x_4774 & x_4776;
assign x_4778 = x_4773 & x_4777;
assign x_4779 = x_4769 & x_4778;
assign x_4780 = x_2156 & x_2157;
assign x_4781 = x_2159 & x_2160;
assign x_4782 = x_2158 & x_4781;
assign x_4783 = x_4780 & x_4782;
assign x_4784 = x_2161 & x_2162;
assign x_4785 = x_2164 & x_2165;
assign x_4786 = x_2163 & x_4785;
assign x_4787 = x_4784 & x_4786;
assign x_4788 = x_4783 & x_4787;
assign x_4789 = x_2166 & x_2167;
assign x_4790 = x_2169 & x_2170;
assign x_4791 = x_2168 & x_4790;
assign x_4792 = x_4789 & x_4791;
assign x_4793 = x_2172 & x_2173;
assign x_4794 = x_2171 & x_4793;
assign x_4795 = x_2175 & x_2176;
assign x_4796 = x_2174 & x_4795;
assign x_4797 = x_4794 & x_4796;
assign x_4798 = x_4792 & x_4797;
assign x_4799 = x_4788 & x_4798;
assign x_4800 = x_4779 & x_4799;
assign x_4801 = x_2177 & x_2178;
assign x_4802 = x_2180 & x_2181;
assign x_4803 = x_2179 & x_4802;
assign x_4804 = x_4801 & x_4803;
assign x_4805 = x_2182 & x_2183;
assign x_4806 = x_2185 & x_2186;
assign x_4807 = x_2184 & x_4806;
assign x_4808 = x_4805 & x_4807;
assign x_4809 = x_4804 & x_4808;
assign x_4810 = x_2187 & x_2188;
assign x_4811 = x_2190 & x_2191;
assign x_4812 = x_2189 & x_4811;
assign x_4813 = x_4810 & x_4812;
assign x_4814 = x_2192 & x_2193;
assign x_4815 = x_2195 & x_2196;
assign x_4816 = x_2194 & x_4815;
assign x_4817 = x_4814 & x_4816;
assign x_4818 = x_4813 & x_4817;
assign x_4819 = x_4809 & x_4818;
assign x_4820 = x_2197 & x_2198;
assign x_4821 = x_2200 & x_2201;
assign x_4822 = x_2199 & x_4821;
assign x_4823 = x_4820 & x_4822;
assign x_4824 = x_2202 & x_2203;
assign x_4825 = x_2205 & x_2206;
assign x_4826 = x_2204 & x_4825;
assign x_4827 = x_4824 & x_4826;
assign x_4828 = x_4823 & x_4827;
assign x_4829 = x_2207 & x_2208;
assign x_4830 = x_2210 & x_2211;
assign x_4831 = x_2209 & x_4830;
assign x_4832 = x_4829 & x_4831;
assign x_4833 = x_2213 & x_2214;
assign x_4834 = x_2212 & x_4833;
assign x_4835 = x_2216 & x_2217;
assign x_4836 = x_2215 & x_4835;
assign x_4837 = x_4834 & x_4836;
assign x_4838 = x_4832 & x_4837;
assign x_4839 = x_4828 & x_4838;
assign x_4840 = x_4819 & x_4839;
assign x_4841 = x_4800 & x_4840;
assign x_4842 = x_2218 & x_2219;
assign x_4843 = x_2221 & x_2222;
assign x_4844 = x_2220 & x_4843;
assign x_4845 = x_4842 & x_4844;
assign x_4846 = x_2223 & x_2224;
assign x_4847 = x_2226 & x_2227;
assign x_4848 = x_2225 & x_4847;
assign x_4849 = x_4846 & x_4848;
assign x_4850 = x_4845 & x_4849;
assign x_4851 = x_2228 & x_2229;
assign x_4852 = x_2231 & x_2232;
assign x_4853 = x_2230 & x_4852;
assign x_4854 = x_4851 & x_4853;
assign x_4855 = x_2233 & x_2234;
assign x_4856 = x_2236 & x_2237;
assign x_4857 = x_2235 & x_4856;
assign x_4858 = x_4855 & x_4857;
assign x_4859 = x_4854 & x_4858;
assign x_4860 = x_4850 & x_4859;
assign x_4861 = x_2238 & x_2239;
assign x_4862 = x_2241 & x_2242;
assign x_4863 = x_2240 & x_4862;
assign x_4864 = x_4861 & x_4863;
assign x_4865 = x_2243 & x_2244;
assign x_4866 = x_2246 & x_2247;
assign x_4867 = x_2245 & x_4866;
assign x_4868 = x_4865 & x_4867;
assign x_4869 = x_4864 & x_4868;
assign x_4870 = x_2248 & x_2249;
assign x_4871 = x_2251 & x_2252;
assign x_4872 = x_2250 & x_4871;
assign x_4873 = x_4870 & x_4872;
assign x_4874 = x_2254 & x_2255;
assign x_4875 = x_2253 & x_4874;
assign x_4876 = x_2257 & x_2258;
assign x_4877 = x_2256 & x_4876;
assign x_4878 = x_4875 & x_4877;
assign x_4879 = x_4873 & x_4878;
assign x_4880 = x_4869 & x_4879;
assign x_4881 = x_4860 & x_4880;
assign x_4882 = x_2259 & x_2260;
assign x_4883 = x_2262 & x_2263;
assign x_4884 = x_2261 & x_4883;
assign x_4885 = x_4882 & x_4884;
assign x_4886 = x_2264 & x_2265;
assign x_4887 = x_2267 & x_2268;
assign x_4888 = x_2266 & x_4887;
assign x_4889 = x_4886 & x_4888;
assign x_4890 = x_4885 & x_4889;
assign x_4891 = x_2269 & x_2270;
assign x_4892 = x_2272 & x_2273;
assign x_4893 = x_2271 & x_4892;
assign x_4894 = x_4891 & x_4893;
assign x_4895 = x_2274 & x_2275;
assign x_4896 = x_2277 & x_2278;
assign x_4897 = x_2276 & x_4896;
assign x_4898 = x_4895 & x_4897;
assign x_4899 = x_4894 & x_4898;
assign x_4900 = x_4890 & x_4899;
assign x_4901 = x_2279 & x_2280;
assign x_4902 = x_2282 & x_2283;
assign x_4903 = x_2281 & x_4902;
assign x_4904 = x_4901 & x_4903;
assign x_4905 = x_2284 & x_2285;
assign x_4906 = x_2287 & x_2288;
assign x_4907 = x_2286 & x_4906;
assign x_4908 = x_4905 & x_4907;
assign x_4909 = x_4904 & x_4908;
assign x_4910 = x_2289 & x_2290;
assign x_4911 = x_2292 & x_2293;
assign x_4912 = x_2291 & x_4911;
assign x_4913 = x_4910 & x_4912;
assign x_4914 = x_2295 & x_2296;
assign x_4915 = x_2294 & x_4914;
assign x_4916 = x_2298 & x_2299;
assign x_4917 = x_2297 & x_4916;
assign x_4918 = x_4915 & x_4917;
assign x_4919 = x_4913 & x_4918;
assign x_4920 = x_4909 & x_4919;
assign x_4921 = x_4900 & x_4920;
assign x_4922 = x_4881 & x_4921;
assign x_4923 = x_4841 & x_4922;
assign x_4924 = x_4760 & x_4923;
assign x_4925 = x_2300 & x_2301;
assign x_4926 = x_2303 & x_2304;
assign x_4927 = x_2302 & x_4926;
assign x_4928 = x_4925 & x_4927;
assign x_4929 = x_2305 & x_2306;
assign x_4930 = x_2308 & x_2309;
assign x_4931 = x_2307 & x_4930;
assign x_4932 = x_4929 & x_4931;
assign x_4933 = x_4928 & x_4932;
assign x_4934 = x_2310 & x_2311;
assign x_4935 = x_2313 & x_2314;
assign x_4936 = x_2312 & x_4935;
assign x_4937 = x_4934 & x_4936;
assign x_4938 = x_2315 & x_2316;
assign x_4939 = x_2318 & x_2319;
assign x_4940 = x_2317 & x_4939;
assign x_4941 = x_4938 & x_4940;
assign x_4942 = x_4937 & x_4941;
assign x_4943 = x_4933 & x_4942;
assign x_4944 = x_2320 & x_2321;
assign x_4945 = x_2323 & x_2324;
assign x_4946 = x_2322 & x_4945;
assign x_4947 = x_4944 & x_4946;
assign x_4948 = x_2325 & x_2326;
assign x_4949 = x_2328 & x_2329;
assign x_4950 = x_2327 & x_4949;
assign x_4951 = x_4948 & x_4950;
assign x_4952 = x_4947 & x_4951;
assign x_4953 = x_2330 & x_2331;
assign x_4954 = x_2333 & x_2334;
assign x_4955 = x_2332 & x_4954;
assign x_4956 = x_4953 & x_4955;
assign x_4957 = x_2336 & x_2337;
assign x_4958 = x_2335 & x_4957;
assign x_4959 = x_2339 & x_2340;
assign x_4960 = x_2338 & x_4959;
assign x_4961 = x_4958 & x_4960;
assign x_4962 = x_4956 & x_4961;
assign x_4963 = x_4952 & x_4962;
assign x_4964 = x_4943 & x_4963;
assign x_4965 = x_2341 & x_2342;
assign x_4966 = x_2344 & x_2345;
assign x_4967 = x_2343 & x_4966;
assign x_4968 = x_4965 & x_4967;
assign x_4969 = x_2346 & x_2347;
assign x_4970 = x_2349 & x_2350;
assign x_4971 = x_2348 & x_4970;
assign x_4972 = x_4969 & x_4971;
assign x_4973 = x_4968 & x_4972;
assign x_4974 = x_2351 & x_2352;
assign x_4975 = x_2354 & x_2355;
assign x_4976 = x_2353 & x_4975;
assign x_4977 = x_4974 & x_4976;
assign x_4978 = x_2356 & x_2357;
assign x_4979 = x_2359 & x_2360;
assign x_4980 = x_2358 & x_4979;
assign x_4981 = x_4978 & x_4980;
assign x_4982 = x_4977 & x_4981;
assign x_4983 = x_4973 & x_4982;
assign x_4984 = x_2361 & x_2362;
assign x_4985 = x_2364 & x_2365;
assign x_4986 = x_2363 & x_4985;
assign x_4987 = x_4984 & x_4986;
assign x_4988 = x_2366 & x_2367;
assign x_4989 = x_2369 & x_2370;
assign x_4990 = x_2368 & x_4989;
assign x_4991 = x_4988 & x_4990;
assign x_4992 = x_4987 & x_4991;
assign x_4993 = x_2371 & x_2372;
assign x_4994 = x_2374 & x_2375;
assign x_4995 = x_2373 & x_4994;
assign x_4996 = x_4993 & x_4995;
assign x_4997 = x_2377 & x_2378;
assign x_4998 = x_2376 & x_4997;
assign x_4999 = x_2380 & x_2381;
assign x_5000 = x_2379 & x_4999;
assign x_5001 = x_4998 & x_5000;
assign x_5002 = x_4996 & x_5001;
assign x_5003 = x_4992 & x_5002;
assign x_5004 = x_4983 & x_5003;
assign x_5005 = x_4964 & x_5004;
assign x_5006 = x_2382 & x_2383;
assign x_5007 = x_2385 & x_2386;
assign x_5008 = x_2384 & x_5007;
assign x_5009 = x_5006 & x_5008;
assign x_5010 = x_2387 & x_2388;
assign x_5011 = x_2390 & x_2391;
assign x_5012 = x_2389 & x_5011;
assign x_5013 = x_5010 & x_5012;
assign x_5014 = x_5009 & x_5013;
assign x_5015 = x_2392 & x_2393;
assign x_5016 = x_2395 & x_2396;
assign x_5017 = x_2394 & x_5016;
assign x_5018 = x_5015 & x_5017;
assign x_5019 = x_2397 & x_2398;
assign x_5020 = x_2400 & x_2401;
assign x_5021 = x_2399 & x_5020;
assign x_5022 = x_5019 & x_5021;
assign x_5023 = x_5018 & x_5022;
assign x_5024 = x_5014 & x_5023;
assign x_5025 = x_2402 & x_2403;
assign x_5026 = x_2405 & x_2406;
assign x_5027 = x_2404 & x_5026;
assign x_5028 = x_5025 & x_5027;
assign x_5029 = x_2407 & x_2408;
assign x_5030 = x_2410 & x_2411;
assign x_5031 = x_2409 & x_5030;
assign x_5032 = x_5029 & x_5031;
assign x_5033 = x_5028 & x_5032;
assign x_5034 = x_2412 & x_2413;
assign x_5035 = x_2415 & x_2416;
assign x_5036 = x_2414 & x_5035;
assign x_5037 = x_5034 & x_5036;
assign x_5038 = x_2418 & x_2419;
assign x_5039 = x_2417 & x_5038;
assign x_5040 = x_2421 & x_2422;
assign x_5041 = x_2420 & x_5040;
assign x_5042 = x_5039 & x_5041;
assign x_5043 = x_5037 & x_5042;
assign x_5044 = x_5033 & x_5043;
assign x_5045 = x_5024 & x_5044;
assign x_5046 = x_2423 & x_2424;
assign x_5047 = x_2426 & x_2427;
assign x_5048 = x_2425 & x_5047;
assign x_5049 = x_5046 & x_5048;
assign x_5050 = x_2428 & x_2429;
assign x_5051 = x_2431 & x_2432;
assign x_5052 = x_2430 & x_5051;
assign x_5053 = x_5050 & x_5052;
assign x_5054 = x_5049 & x_5053;
assign x_5055 = x_2433 & x_2434;
assign x_5056 = x_2436 & x_2437;
assign x_5057 = x_2435 & x_5056;
assign x_5058 = x_5055 & x_5057;
assign x_5059 = x_2438 & x_2439;
assign x_5060 = x_2441 & x_2442;
assign x_5061 = x_2440 & x_5060;
assign x_5062 = x_5059 & x_5061;
assign x_5063 = x_5058 & x_5062;
assign x_5064 = x_5054 & x_5063;
assign x_5065 = x_2443 & x_2444;
assign x_5066 = x_2446 & x_2447;
assign x_5067 = x_2445 & x_5066;
assign x_5068 = x_5065 & x_5067;
assign x_5069 = x_2448 & x_2449;
assign x_5070 = x_2451 & x_2452;
assign x_5071 = x_2450 & x_5070;
assign x_5072 = x_5069 & x_5071;
assign x_5073 = x_5068 & x_5072;
assign x_5074 = x_2453 & x_2454;
assign x_5075 = x_2456 & x_2457;
assign x_5076 = x_2455 & x_5075;
assign x_5077 = x_5074 & x_5076;
assign x_5078 = x_2459 & x_2460;
assign x_5079 = x_2458 & x_5078;
assign x_5080 = x_2462 & x_2463;
assign x_5081 = x_2461 & x_5080;
assign x_5082 = x_5079 & x_5081;
assign x_5083 = x_5077 & x_5082;
assign x_5084 = x_5073 & x_5083;
assign x_5085 = x_5064 & x_5084;
assign x_5086 = x_5045 & x_5085;
assign x_5087 = x_5005 & x_5086;
assign x_5088 = x_2464 & x_2465;
assign x_5089 = x_2467 & x_2468;
assign x_5090 = x_2466 & x_5089;
assign x_5091 = x_5088 & x_5090;
assign x_5092 = x_2469 & x_2470;
assign x_5093 = x_2472 & x_2473;
assign x_5094 = x_2471 & x_5093;
assign x_5095 = x_5092 & x_5094;
assign x_5096 = x_5091 & x_5095;
assign x_5097 = x_2474 & x_2475;
assign x_5098 = x_2477 & x_2478;
assign x_5099 = x_2476 & x_5098;
assign x_5100 = x_5097 & x_5099;
assign x_5101 = x_2479 & x_2480;
assign x_5102 = x_2482 & x_2483;
assign x_5103 = x_2481 & x_5102;
assign x_5104 = x_5101 & x_5103;
assign x_5105 = x_5100 & x_5104;
assign x_5106 = x_5096 & x_5105;
assign x_5107 = x_2484 & x_2485;
assign x_5108 = x_2487 & x_2488;
assign x_5109 = x_2486 & x_5108;
assign x_5110 = x_5107 & x_5109;
assign x_5111 = x_2489 & x_2490;
assign x_5112 = x_2492 & x_2493;
assign x_5113 = x_2491 & x_5112;
assign x_5114 = x_5111 & x_5113;
assign x_5115 = x_5110 & x_5114;
assign x_5116 = x_2494 & x_2495;
assign x_5117 = x_2497 & x_2498;
assign x_5118 = x_2496 & x_5117;
assign x_5119 = x_5116 & x_5118;
assign x_5120 = x_2500 & x_2501;
assign x_5121 = x_2499 & x_5120;
assign x_5122 = x_2503 & x_2504;
assign x_5123 = x_2502 & x_5122;
assign x_5124 = x_5121 & x_5123;
assign x_5125 = x_5119 & x_5124;
assign x_5126 = x_5115 & x_5125;
assign x_5127 = x_5106 & x_5126;
assign x_5128 = x_2505 & x_2506;
assign x_5129 = x_2508 & x_2509;
assign x_5130 = x_2507 & x_5129;
assign x_5131 = x_5128 & x_5130;
assign x_5132 = x_2510 & x_2511;
assign x_5133 = x_2513 & x_2514;
assign x_5134 = x_2512 & x_5133;
assign x_5135 = x_5132 & x_5134;
assign x_5136 = x_5131 & x_5135;
assign x_5137 = x_2515 & x_2516;
assign x_5138 = x_2518 & x_2519;
assign x_5139 = x_2517 & x_5138;
assign x_5140 = x_5137 & x_5139;
assign x_5141 = x_2520 & x_2521;
assign x_5142 = x_2523 & x_2524;
assign x_5143 = x_2522 & x_5142;
assign x_5144 = x_5141 & x_5143;
assign x_5145 = x_5140 & x_5144;
assign x_5146 = x_5136 & x_5145;
assign x_5147 = x_2525 & x_2526;
assign x_5148 = x_2528 & x_2529;
assign x_5149 = x_2527 & x_5148;
assign x_5150 = x_5147 & x_5149;
assign x_5151 = x_2530 & x_2531;
assign x_5152 = x_2533 & x_2534;
assign x_5153 = x_2532 & x_5152;
assign x_5154 = x_5151 & x_5153;
assign x_5155 = x_5150 & x_5154;
assign x_5156 = x_2535 & x_2536;
assign x_5157 = x_2538 & x_2539;
assign x_5158 = x_2537 & x_5157;
assign x_5159 = x_5156 & x_5158;
assign x_5160 = x_2541 & x_2542;
assign x_5161 = x_2540 & x_5160;
assign x_5162 = x_2544 & x_2545;
assign x_5163 = x_2543 & x_5162;
assign x_5164 = x_5161 & x_5163;
assign x_5165 = x_5159 & x_5164;
assign x_5166 = x_5155 & x_5165;
assign x_5167 = x_5146 & x_5166;
assign x_5168 = x_5127 & x_5167;
assign x_5169 = x_2546 & x_2547;
assign x_5170 = x_2549 & x_2550;
assign x_5171 = x_2548 & x_5170;
assign x_5172 = x_5169 & x_5171;
assign x_5173 = x_2551 & x_2552;
assign x_5174 = x_2554 & x_2555;
assign x_5175 = x_2553 & x_5174;
assign x_5176 = x_5173 & x_5175;
assign x_5177 = x_5172 & x_5176;
assign x_5178 = x_2556 & x_2557;
assign x_5179 = x_2559 & x_2560;
assign x_5180 = x_2558 & x_5179;
assign x_5181 = x_5178 & x_5180;
assign x_5182 = x_2561 & x_2562;
assign x_5183 = x_2564 & x_2565;
assign x_5184 = x_2563 & x_5183;
assign x_5185 = x_5182 & x_5184;
assign x_5186 = x_5181 & x_5185;
assign x_5187 = x_5177 & x_5186;
assign x_5188 = x_2566 & x_2567;
assign x_5189 = x_2569 & x_2570;
assign x_5190 = x_2568 & x_5189;
assign x_5191 = x_5188 & x_5190;
assign x_5192 = x_2571 & x_2572;
assign x_5193 = x_2574 & x_2575;
assign x_5194 = x_2573 & x_5193;
assign x_5195 = x_5192 & x_5194;
assign x_5196 = x_5191 & x_5195;
assign x_5197 = x_2576 & x_2577;
assign x_5198 = x_2579 & x_2580;
assign x_5199 = x_2578 & x_5198;
assign x_5200 = x_5197 & x_5199;
assign x_5201 = x_2582 & x_2583;
assign x_5202 = x_2581 & x_5201;
assign x_5203 = x_2585 & x_2586;
assign x_5204 = x_2584 & x_5203;
assign x_5205 = x_5202 & x_5204;
assign x_5206 = x_5200 & x_5205;
assign x_5207 = x_5196 & x_5206;
assign x_5208 = x_5187 & x_5207;
assign x_5209 = x_2587 & x_2588;
assign x_5210 = x_2590 & x_2591;
assign x_5211 = x_2589 & x_5210;
assign x_5212 = x_5209 & x_5211;
assign x_5213 = x_2592 & x_2593;
assign x_5214 = x_2595 & x_2596;
assign x_5215 = x_2594 & x_5214;
assign x_5216 = x_5213 & x_5215;
assign x_5217 = x_5212 & x_5216;
assign x_5218 = x_2597 & x_2598;
assign x_5219 = x_2600 & x_2601;
assign x_5220 = x_2599 & x_5219;
assign x_5221 = x_5218 & x_5220;
assign x_5222 = x_2603 & x_2604;
assign x_5223 = x_2602 & x_5222;
assign x_5224 = x_2606 & x_2607;
assign x_5225 = x_2605 & x_5224;
assign x_5226 = x_5223 & x_5225;
assign x_5227 = x_5221 & x_5226;
assign x_5228 = x_5217 & x_5227;
assign x_5229 = x_2608 & x_2609;
assign x_5230 = x_2611 & x_2612;
assign x_5231 = x_2610 & x_5230;
assign x_5232 = x_5229 & x_5231;
assign x_5233 = x_2613 & x_2614;
assign x_5234 = x_2616 & x_2617;
assign x_5235 = x_2615 & x_5234;
assign x_5236 = x_5233 & x_5235;
assign x_5237 = x_5232 & x_5236;
assign x_5238 = x_2618 & x_2619;
assign x_5239 = x_2621 & x_2622;
assign x_5240 = x_2620 & x_5239;
assign x_5241 = x_5238 & x_5240;
assign x_5242 = x_2624 & x_2625;
assign x_5243 = x_2623 & x_5242;
assign x_5244 = x_2627 & x_2628;
assign x_5245 = x_2626 & x_5244;
assign x_5246 = x_5243 & x_5245;
assign x_5247 = x_5241 & x_5246;
assign x_5248 = x_5237 & x_5247;
assign x_5249 = x_5228 & x_5248;
assign x_5250 = x_5208 & x_5249;
assign x_5251 = x_5168 & x_5250;
assign x_5252 = x_5087 & x_5251;
assign x_5253 = x_4924 & x_5252;
assign x_5254 = x_4597 & x_5253;
assign x_5255 = x_3941 & x_5254;
assign o_1 = x_5255;
endmodule
