// Benchmark "SKOLEMFORMULA" written by ABC on Thu Jul  1 18:41:40 2021

module SKOLEMFORMULA ( 
    i0, i1,
    i2  );
  input  i0, i1;
  output i2;
  assign i2 = i0 & i1;
endmodule
