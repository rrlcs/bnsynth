// skolem function for order file variables
// Generated using findDep.cpp 
module formula (v_169, v_182, v_1446, v_1456, v_1466, v_130, v_143, v_156, v_262, v_275, v_288, v_1336, v_1346, v_1356, v_487, v_500, v_513, v_876, v_1306, v_1316, v_1326, v_1056, v_223, v_236, v_249, v_806, v_819, v_832, v_4, v_3, v_97, v_110, v_123, v_140, v_153, v_166, v_179, v_12, v_15, v_220, v_233, v_246, v_259, v_272, v_285, v_6, v_8, v_2, v_400, v_419, v_432, v_445, v_458, v_471, v_484, v_497, v_510, v_523, v_544, v_559, v_631, v_703, v_580, v_601, v_616, v_688, v_686, v_639, v_633, v_646, v_803, v_816, v_829, v_1, v_10, v_44, v_33, v_886, v_880, v_899, v_893, v_906, v_953, v_944, v_963, v_658, v_13, v_17, v_20, v_23, v_653, v_655, v_667, v_1001, v_995, v_1008, v_955, v_946, v_965, v_930, v_924, v_937, v_529, v_547, v_562, v_586, v_604, v_619, v_25, v_65, v_64, v_67, v_87, v_100, v_113, v_1286, v_1296, v_684, v_76, v_315, v_409, v_422, v_435, v_448, v_461, v_474, v_694, v_303, v_70, v_69, v_72, v_74, v_309, v_61, v_62, v_96, v_109, v_122, v_139, v_152, v_165, v_178, v_191, v_208, v_219, v_232, v_245, v_258, v_271, v_284, v_297, v_373, v_388, v_399, v_418, v_431, v_444, v_457, v_470, v_483, v_496, v_509, v_522, v_543, v_558, v_573, v_576, v_579, v_600, v_615, v_630, v_760, v_775, v_784, v_793, v_802, v_815, v_828, v_841, v_1237, v_1260, v_1273, v_1284, v_1294, v_1304, v_1314, v_1324, v_1334, v_1344, v_1354, v_1364, v_1367, v_1374, v_1387, v_1400, v_1413, v_1426, v_1435, v_1444, v_1454, v_1464, v_1474, v_1487, v_1496, v_1505, v_1514, v_1523, v_1532, v_1541, v_1550, v_1559, v_1568, v_1577, v_1586, o_1);
input v_169;
input v_182;
input v_1446;
input v_1456;
input v_1466;
input v_130;
input v_143;
input v_156;
input v_262;
input v_275;
input v_288;
input v_1336;
input v_1346;
input v_1356;
input v_487;
input v_500;
input v_513;
input v_876;
input v_1306;
input v_1316;
input v_1326;
input v_1056;
input v_223;
input v_236;
input v_249;
input v_806;
input v_819;
input v_832;
input v_4;
input v_3;
input v_97;
input v_110;
input v_123;
input v_140;
input v_153;
input v_166;
input v_179;
input v_12;
input v_15;
input v_220;
input v_233;
input v_246;
input v_259;
input v_272;
input v_285;
input v_6;
input v_8;
input v_2;
input v_400;
input v_419;
input v_432;
input v_445;
input v_458;
input v_471;
input v_484;
input v_497;
input v_510;
input v_523;
input v_544;
input v_559;
input v_631;
input v_703;
input v_580;
input v_601;
input v_616;
input v_688;
input v_686;
input v_639;
input v_633;
input v_646;
input v_803;
input v_816;
input v_829;
input v_1;
input v_10;
input v_44;
input v_33;
input v_886;
input v_880;
input v_899;
input v_893;
input v_906;
input v_953;
input v_944;
input v_963;
input v_658;
input v_13;
input v_17;
input v_20;
input v_23;
input v_653;
input v_655;
input v_667;
input v_1001;
input v_995;
input v_1008;
input v_955;
input v_946;
input v_965;
input v_930;
input v_924;
input v_937;
input v_529;
input v_547;
input v_562;
input v_586;
input v_604;
input v_619;
input v_25;
input v_65;
input v_64;
input v_67;
input v_87;
input v_100;
input v_113;
input v_1286;
input v_1296;
input v_684;
input v_76;
input v_315;
input v_409;
input v_422;
input v_435;
input v_448;
input v_461;
input v_474;
input v_694;
input v_303;
input v_70;
input v_69;
input v_72;
input v_74;
input v_309;
input v_61;
input v_62;
input v_96;
input v_109;
input v_122;
input v_139;
input v_152;
input v_165;
input v_178;
input v_191;
input v_208;
input v_219;
input v_232;
input v_245;
input v_258;
input v_271;
input v_284;
input v_297;
input v_373;
input v_388;
input v_399;
input v_418;
input v_431;
input v_444;
input v_457;
input v_470;
input v_483;
input v_496;
input v_509;
input v_522;
input v_543;
input v_558;
input v_573;
input v_576;
input v_579;
input v_600;
input v_615;
input v_630;
input v_760;
input v_775;
input v_784;
input v_793;
input v_802;
input v_815;
input v_828;
input v_841;
input v_1237;
input v_1260;
input v_1273;
input v_1284;
input v_1294;
input v_1304;
input v_1314;
input v_1324;
input v_1334;
input v_1344;
input v_1354;
input v_1364;
input v_1367;
input v_1374;
input v_1387;
input v_1400;
input v_1413;
input v_1426;
input v_1435;
input v_1444;
input v_1454;
input v_1464;
input v_1474;
input v_1487;
input v_1496;
input v_1505;
input v_1514;
input v_1523;
input v_1532;
input v_1541;
input v_1550;
input v_1559;
input v_1568;
input v_1577;
input v_1586;
output o_1;
wire v_5;
wire v_7;
wire v_9;
wire v_11;
wire v_14;
wire v_16;
wire v_18;
wire v_19;
wire v_21;
wire v_22;
wire v_24;
wire v_26;
wire v_27;
wire v_28;
wire v_29;
wire v_30;
wire v_31;
wire v_32;
wire v_34;
wire v_35;
wire v_36;
wire v_37;
wire v_38;
wire v_39;
wire v_40;
wire v_41;
wire v_42;
wire v_43;
wire v_45;
wire v_46;
wire v_47;
wire v_48;
wire v_49;
wire v_50;
wire v_51;
wire v_52;
wire v_53;
wire v_54;
wire v_55;
wire v_56;
wire v_57;
wire v_58;
wire v_59;
wire v_60;
wire v_63;
wire v_66;
wire v_68;
wire v_71;
wire v_73;
wire v_75;
wire v_77;
wire v_78;
wire v_79;
wire v_80;
wire v_81;
wire v_82;
wire v_83;
wire v_84;
wire v_85;
wire v_86;
wire v_88;
wire v_89;
wire v_90;
wire v_91;
wire v_92;
wire v_93;
wire v_94;
wire v_95;
wire v_98;
wire v_99;
wire v_101;
wire v_102;
wire v_103;
wire v_104;
wire v_105;
wire v_106;
wire v_107;
wire v_108;
wire v_111;
wire v_112;
wire v_114;
wire v_115;
wire v_116;
wire v_117;
wire v_118;
wire v_119;
wire v_120;
wire v_121;
wire v_124;
wire v_125;
wire v_126;
wire v_127;
wire v_128;
wire v_129;
wire v_131;
wire v_132;
wire v_133;
wire v_134;
wire v_135;
wire v_136;
wire v_137;
wire v_138;
wire v_141;
wire v_142;
wire v_144;
wire v_145;
wire v_146;
wire v_147;
wire v_148;
wire v_149;
wire v_150;
wire v_151;
wire v_154;
wire v_155;
wire v_157;
wire v_158;
wire v_159;
wire v_160;
wire v_161;
wire v_162;
wire v_163;
wire v_164;
wire v_167;
wire v_168;
wire v_170;
wire v_171;
wire v_172;
wire v_173;
wire v_174;
wire v_175;
wire v_176;
wire v_177;
wire v_180;
wire v_181;
wire v_183;
wire v_184;
wire v_185;
wire v_186;
wire v_187;
wire v_188;
wire v_189;
wire v_190;
wire v_192;
wire v_193;
wire v_194;
wire v_195;
wire v_196;
wire v_197;
wire v_198;
wire v_199;
wire v_200;
wire v_201;
wire v_202;
wire v_203;
wire v_204;
wire v_205;
wire v_206;
wire v_207;
wire v_209;
wire v_210;
wire v_211;
wire v_212;
wire v_213;
wire v_214;
wire v_215;
wire v_216;
wire v_217;
wire v_218;
wire v_221;
wire v_222;
wire v_224;
wire v_225;
wire v_226;
wire v_227;
wire v_228;
wire v_229;
wire v_230;
wire v_231;
wire v_234;
wire v_235;
wire v_237;
wire v_238;
wire v_239;
wire v_240;
wire v_241;
wire v_242;
wire v_243;
wire v_244;
wire v_247;
wire v_248;
wire v_250;
wire v_251;
wire v_252;
wire v_253;
wire v_254;
wire v_255;
wire v_256;
wire v_257;
wire v_260;
wire v_261;
wire v_263;
wire v_264;
wire v_265;
wire v_266;
wire v_267;
wire v_268;
wire v_269;
wire v_270;
wire v_273;
wire v_274;
wire v_276;
wire v_277;
wire v_278;
wire v_279;
wire v_280;
wire v_281;
wire v_282;
wire v_283;
wire v_286;
wire v_287;
wire v_289;
wire v_290;
wire v_291;
wire v_292;
wire v_293;
wire v_294;
wire v_295;
wire v_296;
wire v_298;
wire v_299;
wire v_300;
wire v_301;
wire v_302;
wire v_304;
wire v_305;
wire v_306;
wire v_307;
wire v_308;
wire v_310;
wire v_311;
wire v_312;
wire v_313;
wire v_314;
wire v_316;
wire v_317;
wire v_318;
wire v_319;
wire v_320;
wire v_321;
wire v_322;
wire v_323;
wire v_324;
wire v_325;
wire v_326;
wire v_327;
wire v_328;
wire v_329;
wire v_330;
wire v_331;
wire v_332;
wire v_333;
wire v_334;
wire v_335;
wire v_336;
wire v_337;
wire v_338;
wire v_339;
wire v_340;
wire v_341;
wire v_342;
wire v_343;
wire v_344;
wire v_345;
wire v_346;
wire v_347;
wire v_348;
wire v_349;
wire v_350;
wire v_351;
wire v_352;
wire v_353;
wire v_354;
wire v_355;
wire v_356;
wire v_357;
wire v_358;
wire v_359;
wire v_360;
wire v_361;
wire v_362;
wire v_363;
wire v_364;
wire v_365;
wire v_366;
wire v_367;
wire v_368;
wire v_369;
wire v_370;
wire v_371;
wire v_372;
wire v_374;
wire v_375;
wire v_376;
wire v_377;
wire v_378;
wire v_379;
wire v_380;
wire v_381;
wire v_382;
wire v_383;
wire v_384;
wire v_385;
wire v_386;
wire v_387;
wire v_389;
wire v_390;
wire v_391;
wire v_392;
wire v_393;
wire v_394;
wire v_395;
wire v_396;
wire v_397;
wire v_398;
wire v_401;
wire v_402;
wire v_403;
wire v_404;
wire v_405;
wire v_406;
wire v_407;
wire v_408;
wire v_410;
wire v_411;
wire v_412;
wire v_413;
wire v_414;
wire v_415;
wire v_416;
wire v_417;
wire v_420;
wire v_421;
wire v_423;
wire v_424;
wire v_425;
wire v_426;
wire v_427;
wire v_428;
wire v_429;
wire v_430;
wire v_433;
wire v_434;
wire v_436;
wire v_437;
wire v_438;
wire v_439;
wire v_440;
wire v_441;
wire v_442;
wire v_443;
wire v_446;
wire v_447;
wire v_449;
wire v_450;
wire v_451;
wire v_452;
wire v_453;
wire v_454;
wire v_455;
wire v_456;
wire v_459;
wire v_460;
wire v_462;
wire v_463;
wire v_464;
wire v_465;
wire v_466;
wire v_467;
wire v_468;
wire v_469;
wire v_472;
wire v_473;
wire v_475;
wire v_476;
wire v_477;
wire v_478;
wire v_479;
wire v_480;
wire v_481;
wire v_482;
wire v_485;
wire v_486;
wire v_488;
wire v_489;
wire v_490;
wire v_491;
wire v_492;
wire v_493;
wire v_494;
wire v_495;
wire v_498;
wire v_499;
wire v_501;
wire v_502;
wire v_503;
wire v_504;
wire v_505;
wire v_506;
wire v_507;
wire v_508;
wire v_511;
wire v_512;
wire v_514;
wire v_515;
wire v_516;
wire v_517;
wire v_518;
wire v_519;
wire v_520;
wire v_521;
wire v_524;
wire v_525;
wire v_526;
wire v_527;
wire v_528;
wire v_530;
wire v_531;
wire v_532;
wire v_533;
wire v_534;
wire v_535;
wire v_536;
wire v_537;
wire v_538;
wire v_539;
wire v_540;
wire v_541;
wire v_542;
wire v_545;
wire v_546;
wire v_548;
wire v_549;
wire v_550;
wire v_551;
wire v_552;
wire v_553;
wire v_554;
wire v_555;
wire v_556;
wire v_557;
wire v_560;
wire v_561;
wire v_563;
wire v_564;
wire v_565;
wire v_566;
wire v_567;
wire v_568;
wire v_569;
wire v_570;
wire v_571;
wire v_572;
wire v_574;
wire v_575;
wire v_577;
wire v_578;
wire v_581;
wire v_582;
wire v_583;
wire v_584;
wire v_585;
wire v_587;
wire v_588;
wire v_589;
wire v_590;
wire v_591;
wire v_592;
wire v_593;
wire v_594;
wire v_595;
wire v_596;
wire v_597;
wire v_598;
wire v_599;
wire v_602;
wire v_603;
wire v_605;
wire v_606;
wire v_607;
wire v_608;
wire v_609;
wire v_610;
wire v_611;
wire v_612;
wire v_613;
wire v_614;
wire v_617;
wire v_618;
wire v_620;
wire v_621;
wire v_622;
wire v_623;
wire v_624;
wire v_625;
wire v_626;
wire v_627;
wire v_628;
wire v_629;
wire v_632;
wire v_634;
wire v_635;
wire v_636;
wire v_637;
wire v_638;
wire v_640;
wire v_641;
wire v_642;
wire v_643;
wire v_644;
wire v_645;
wire v_647;
wire v_648;
wire v_649;
wire v_650;
wire v_651;
wire v_652;
wire v_654;
wire v_656;
wire v_657;
wire v_659;
wire v_660;
wire v_661;
wire v_662;
wire v_663;
wire v_664;
wire v_665;
wire v_666;
wire v_668;
wire v_669;
wire v_670;
wire v_671;
wire v_672;
wire v_673;
wire v_674;
wire v_675;
wire v_676;
wire v_677;
wire v_678;
wire v_679;
wire v_680;
wire v_681;
wire v_682;
wire v_683;
wire v_685;
wire v_687;
wire v_689;
wire v_690;
wire v_691;
wire v_692;
wire v_693;
wire v_695;
wire v_696;
wire v_697;
wire v_698;
wire v_699;
wire v_700;
wire v_701;
wire v_702;
wire v_704;
wire v_705;
wire v_706;
wire v_707;
wire v_708;
wire v_709;
wire v_710;
wire v_711;
wire v_712;
wire v_713;
wire v_714;
wire v_715;
wire v_716;
wire v_717;
wire v_718;
wire v_719;
wire v_720;
wire v_721;
wire v_722;
wire v_723;
wire v_724;
wire v_725;
wire v_726;
wire v_727;
wire v_728;
wire v_729;
wire v_730;
wire v_731;
wire v_732;
wire v_733;
wire v_734;
wire v_735;
wire v_736;
wire v_737;
wire v_738;
wire v_739;
wire v_740;
wire v_741;
wire v_742;
wire v_743;
wire v_744;
wire v_745;
wire v_746;
wire v_747;
wire v_748;
wire v_749;
wire v_750;
wire v_751;
wire v_752;
wire v_753;
wire v_754;
wire v_755;
wire v_756;
wire v_757;
wire v_758;
wire v_759;
wire v_761;
wire v_762;
wire v_763;
wire v_764;
wire v_765;
wire v_766;
wire v_767;
wire v_768;
wire v_769;
wire v_770;
wire v_771;
wire v_772;
wire v_773;
wire v_774;
wire v_776;
wire v_777;
wire v_778;
wire v_779;
wire v_780;
wire v_781;
wire v_782;
wire v_783;
wire v_785;
wire v_786;
wire v_787;
wire v_788;
wire v_789;
wire v_790;
wire v_791;
wire v_792;
wire v_794;
wire v_795;
wire v_796;
wire v_797;
wire v_798;
wire v_799;
wire v_800;
wire v_801;
wire v_804;
wire v_805;
wire v_807;
wire v_808;
wire v_809;
wire v_810;
wire v_811;
wire v_812;
wire v_813;
wire v_814;
wire v_817;
wire v_818;
wire v_820;
wire v_821;
wire v_822;
wire v_823;
wire v_824;
wire v_825;
wire v_826;
wire v_827;
wire v_830;
wire v_831;
wire v_833;
wire v_834;
wire v_835;
wire v_836;
wire v_837;
wire v_838;
wire v_839;
wire v_840;
wire v_842;
wire v_843;
wire v_844;
wire v_845;
wire v_846;
wire v_847;
wire v_848;
wire v_849;
wire v_850;
wire v_851;
wire v_852;
wire v_853;
wire v_854;
wire v_855;
wire v_856;
wire v_857;
wire v_858;
wire v_859;
wire v_860;
wire v_861;
wire v_862;
wire v_863;
wire v_864;
wire v_865;
wire v_866;
wire v_867;
wire v_868;
wire v_869;
wire v_870;
wire v_871;
wire v_872;
wire v_873;
wire v_874;
wire v_875;
wire v_877;
wire v_878;
wire v_879;
wire v_881;
wire v_882;
wire v_883;
wire v_884;
wire v_885;
wire v_887;
wire v_888;
wire v_889;
wire v_890;
wire v_891;
wire v_892;
wire v_894;
wire v_895;
wire v_896;
wire v_897;
wire v_898;
wire v_900;
wire v_901;
wire v_902;
wire v_903;
wire v_904;
wire v_905;
wire v_907;
wire v_908;
wire v_909;
wire v_910;
wire v_911;
wire v_912;
wire v_913;
wire v_914;
wire v_915;
wire v_916;
wire v_917;
wire v_918;
wire v_919;
wire v_920;
wire v_921;
wire v_922;
wire v_923;
wire v_925;
wire v_926;
wire v_927;
wire v_928;
wire v_929;
wire v_931;
wire v_932;
wire v_933;
wire v_934;
wire v_935;
wire v_936;
wire v_938;
wire v_939;
wire v_940;
wire v_941;
wire v_942;
wire v_943;
wire v_945;
wire v_947;
wire v_948;
wire v_949;
wire v_950;
wire v_951;
wire v_952;
wire v_954;
wire v_956;
wire v_957;
wire v_958;
wire v_959;
wire v_960;
wire v_961;
wire v_962;
wire v_964;
wire v_966;
wire v_967;
wire v_968;
wire v_969;
wire v_970;
wire v_971;
wire v_972;
wire v_973;
wire v_974;
wire v_975;
wire v_976;
wire v_977;
wire v_978;
wire v_979;
wire v_980;
wire v_981;
wire v_982;
wire v_983;
wire v_984;
wire v_985;
wire v_986;
wire v_987;
wire v_988;
wire v_989;
wire v_990;
wire v_991;
wire v_992;
wire v_993;
wire v_994;
wire v_996;
wire v_997;
wire v_998;
wire v_999;
wire v_1000;
wire v_1002;
wire v_1003;
wire v_1004;
wire v_1005;
wire v_1006;
wire v_1007;
wire v_1009;
wire v_1010;
wire v_1011;
wire v_1012;
wire v_1013;
wire v_1014;
wire v_1015;
wire v_1016;
wire v_1017;
wire v_1018;
wire v_1019;
wire v_1020;
wire v_1021;
wire v_1022;
wire v_1023;
wire v_1024;
wire v_1025;
wire v_1026;
wire v_1027;
wire v_1028;
wire v_1029;
wire v_1030;
wire v_1031;
wire v_1032;
wire v_1033;
wire v_1034;
wire v_1035;
wire v_1036;
wire v_1037;
wire v_1038;
wire v_1039;
wire v_1040;
wire v_1041;
wire v_1042;
wire v_1043;
wire v_1044;
wire v_1045;
wire v_1046;
wire v_1047;
wire v_1048;
wire v_1049;
wire v_1050;
wire v_1051;
wire v_1052;
wire v_1053;
wire v_1054;
wire v_1055;
wire v_1057;
wire v_1058;
wire v_1059;
wire v_1060;
wire v_1061;
wire v_1062;
wire v_1063;
wire v_1064;
wire v_1065;
wire v_1066;
wire v_1067;
wire v_1068;
wire v_1069;
wire v_1070;
wire v_1071;
wire v_1072;
wire v_1073;
wire v_1074;
wire v_1075;
wire v_1076;
wire v_1077;
wire v_1078;
wire v_1079;
wire v_1080;
wire v_1081;
wire v_1082;
wire v_1083;
wire v_1084;
wire v_1085;
wire v_1086;
wire v_1087;
wire v_1088;
wire v_1089;
wire v_1090;
wire v_1091;
wire v_1092;
wire v_1093;
wire v_1094;
wire v_1095;
wire v_1096;
wire v_1097;
wire v_1098;
wire v_1099;
wire v_1100;
wire v_1101;
wire v_1102;
wire v_1103;
wire v_1104;
wire v_1105;
wire v_1106;
wire v_1107;
wire v_1108;
wire v_1109;
wire v_1110;
wire v_1111;
wire v_1112;
wire v_1113;
wire v_1114;
wire v_1115;
wire v_1116;
wire v_1117;
wire v_1118;
wire v_1119;
wire v_1120;
wire v_1121;
wire v_1122;
wire v_1123;
wire v_1124;
wire v_1125;
wire v_1126;
wire v_1127;
wire v_1128;
wire v_1129;
wire v_1130;
wire v_1131;
wire v_1132;
wire v_1133;
wire v_1134;
wire v_1135;
wire v_1136;
wire v_1137;
wire v_1138;
wire v_1139;
wire v_1140;
wire v_1141;
wire v_1142;
wire v_1143;
wire v_1144;
wire v_1145;
wire v_1146;
wire v_1147;
wire v_1148;
wire v_1149;
wire v_1150;
wire v_1151;
wire v_1152;
wire v_1153;
wire v_1154;
wire v_1155;
wire v_1156;
wire v_1157;
wire v_1158;
wire v_1159;
wire v_1160;
wire v_1161;
wire v_1162;
wire v_1163;
wire v_1164;
wire v_1165;
wire v_1166;
wire v_1167;
wire v_1168;
wire v_1169;
wire v_1170;
wire v_1171;
wire v_1172;
wire v_1173;
wire v_1174;
wire v_1175;
wire v_1176;
wire v_1177;
wire v_1178;
wire v_1179;
wire v_1180;
wire v_1181;
wire v_1182;
wire v_1183;
wire v_1184;
wire v_1185;
wire v_1186;
wire v_1187;
wire v_1188;
wire v_1189;
wire v_1190;
wire v_1191;
wire v_1192;
wire v_1193;
wire v_1194;
wire v_1195;
wire v_1196;
wire v_1197;
wire v_1198;
wire v_1199;
wire v_1200;
wire v_1201;
wire v_1202;
wire v_1203;
wire v_1204;
wire v_1205;
wire v_1206;
wire v_1207;
wire v_1208;
wire v_1209;
wire v_1210;
wire v_1211;
wire v_1212;
wire v_1213;
wire v_1214;
wire v_1215;
wire v_1216;
wire v_1217;
wire v_1218;
wire v_1219;
wire v_1220;
wire v_1221;
wire v_1222;
wire v_1223;
wire v_1224;
wire v_1225;
wire v_1226;
wire v_1227;
wire v_1228;
wire v_1229;
wire v_1230;
wire v_1231;
wire v_1232;
wire v_1233;
wire v_1234;
wire v_1235;
wire v_1236;
wire v_1238;
wire v_1239;
wire v_1240;
wire v_1241;
wire v_1242;
wire v_1243;
wire v_1244;
wire v_1245;
wire v_1246;
wire v_1247;
wire v_1248;
wire v_1249;
wire v_1250;
wire v_1251;
wire v_1252;
wire v_1253;
wire v_1254;
wire v_1255;
wire v_1256;
wire v_1257;
wire v_1258;
wire v_1259;
wire v_1261;
wire v_1262;
wire v_1263;
wire v_1264;
wire v_1265;
wire v_1266;
wire v_1267;
wire v_1268;
wire v_1269;
wire v_1270;
wire v_1271;
wire v_1272;
wire v_1274;
wire v_1275;
wire v_1276;
wire v_1277;
wire v_1278;
wire v_1279;
wire v_1280;
wire v_1281;
wire v_1282;
wire v_1283;
wire v_1285;
wire v_1287;
wire v_1288;
wire v_1289;
wire v_1290;
wire v_1291;
wire v_1292;
wire v_1293;
wire v_1295;
wire v_1297;
wire v_1298;
wire v_1299;
wire v_1300;
wire v_1301;
wire v_1302;
wire v_1303;
wire v_1305;
wire v_1307;
wire v_1308;
wire v_1309;
wire v_1310;
wire v_1311;
wire v_1312;
wire v_1313;
wire v_1315;
wire v_1317;
wire v_1318;
wire v_1319;
wire v_1320;
wire v_1321;
wire v_1322;
wire v_1323;
wire v_1325;
wire v_1327;
wire v_1328;
wire v_1329;
wire v_1330;
wire v_1331;
wire v_1332;
wire v_1333;
wire v_1335;
wire v_1337;
wire v_1338;
wire v_1339;
wire v_1340;
wire v_1341;
wire v_1342;
wire v_1343;
wire v_1345;
wire v_1347;
wire v_1348;
wire v_1349;
wire v_1350;
wire v_1351;
wire v_1352;
wire v_1353;
wire v_1355;
wire v_1357;
wire v_1358;
wire v_1359;
wire v_1360;
wire v_1361;
wire v_1362;
wire v_1363;
wire v_1365;
wire v_1366;
wire v_1368;
wire v_1369;
wire v_1370;
wire v_1371;
wire v_1372;
wire v_1373;
wire v_1375;
wire v_1376;
wire v_1377;
wire v_1378;
wire v_1379;
wire v_1380;
wire v_1381;
wire v_1382;
wire v_1383;
wire v_1384;
wire v_1385;
wire v_1386;
wire v_1388;
wire v_1389;
wire v_1390;
wire v_1391;
wire v_1392;
wire v_1393;
wire v_1394;
wire v_1395;
wire v_1396;
wire v_1397;
wire v_1398;
wire v_1399;
wire v_1401;
wire v_1402;
wire v_1403;
wire v_1404;
wire v_1405;
wire v_1406;
wire v_1407;
wire v_1408;
wire v_1409;
wire v_1410;
wire v_1411;
wire v_1412;
wire v_1414;
wire v_1415;
wire v_1416;
wire v_1417;
wire v_1418;
wire v_1419;
wire v_1420;
wire v_1421;
wire v_1422;
wire v_1423;
wire v_1424;
wire v_1425;
wire v_1427;
wire v_1428;
wire v_1429;
wire v_1430;
wire v_1431;
wire v_1432;
wire v_1433;
wire v_1434;
wire v_1436;
wire v_1437;
wire v_1438;
wire v_1439;
wire v_1440;
wire v_1441;
wire v_1442;
wire v_1443;
wire v_1445;
wire v_1447;
wire v_1448;
wire v_1449;
wire v_1450;
wire v_1451;
wire v_1452;
wire v_1453;
wire v_1455;
wire v_1457;
wire v_1458;
wire v_1459;
wire v_1460;
wire v_1461;
wire v_1462;
wire v_1463;
wire v_1465;
wire v_1467;
wire v_1468;
wire v_1469;
wire v_1470;
wire v_1471;
wire v_1472;
wire v_1473;
wire v_1475;
wire v_1476;
wire v_1477;
wire v_1478;
wire v_1479;
wire v_1480;
wire v_1481;
wire v_1482;
wire v_1483;
wire v_1484;
wire v_1485;
wire v_1486;
wire v_1488;
wire v_1489;
wire v_1490;
wire v_1491;
wire v_1492;
wire v_1493;
wire v_1494;
wire v_1495;
wire v_1497;
wire v_1498;
wire v_1499;
wire v_1500;
wire v_1501;
wire v_1502;
wire v_1503;
wire v_1504;
wire v_1506;
wire v_1507;
wire v_1508;
wire v_1509;
wire v_1510;
wire v_1511;
wire v_1512;
wire v_1513;
wire v_1515;
wire v_1516;
wire v_1517;
wire v_1518;
wire v_1519;
wire v_1520;
wire v_1521;
wire v_1522;
wire v_1524;
wire v_1525;
wire v_1526;
wire v_1527;
wire v_1528;
wire v_1529;
wire v_1530;
wire v_1531;
wire v_1533;
wire v_1534;
wire v_1535;
wire v_1536;
wire v_1537;
wire v_1538;
wire v_1539;
wire v_1540;
wire v_1542;
wire v_1543;
wire v_1544;
wire v_1545;
wire v_1546;
wire v_1547;
wire v_1548;
wire v_1549;
wire v_1551;
wire v_1552;
wire v_1553;
wire v_1554;
wire v_1555;
wire v_1556;
wire v_1557;
wire v_1558;
wire v_1560;
wire v_1561;
wire v_1562;
wire v_1563;
wire v_1564;
wire v_1565;
wire v_1566;
wire v_1567;
wire v_1569;
wire v_1570;
wire v_1571;
wire v_1572;
wire v_1573;
wire v_1574;
wire v_1575;
wire v_1576;
wire v_1578;
wire v_1579;
wire v_1580;
wire v_1581;
wire v_1582;
wire v_1583;
wire v_1584;
wire v_1585;
wire v_1587;
wire v_1588;
wire v_1589;
wire v_1590;
wire v_1591;
wire v_1592;
wire v_1593;
wire v_1594;
wire v_1595;
wire v_1596;
wire v_1597;
wire v_1598;
wire v_1599;
wire v_1600;
wire v_1601;
wire v_1602;
wire v_1603;
wire v_1604;
wire v_1605;
wire v_1606;
wire v_1607;
wire v_1608;
wire v_1609;
wire v_1610;
wire v_1611;
wire v_1612;
wire v_1613;
wire v_1614;
wire v_1615;
wire v_1616;
wire v_1617;
wire v_1618;
wire v_1619;
wire v_1620;
wire v_1621;
wire v_1622;
wire v_1623;
wire v_1624;
wire v_1625;
wire v_1626;
wire v_1627;
wire v_1628;
wire v_1629;
wire v_1630;
wire v_1631;
wire v_1632;
wire v_1633;
wire v_1634;
wire v_1635;
wire v_1636;
wire v_1637;
wire v_1638;
wire v_1639;
wire v_1640;
wire v_1641;
wire v_1642;
wire v_1643;
wire v_1644;
wire v_1645;
wire v_1646;
wire v_1647;
wire v_1648;
wire v_1649;
wire v_1650;
wire v_1651;
wire v_1652;
wire v_1653;
wire v_1654;
wire v_1655;
wire v_1656;
wire v_1657;
wire v_1658;
wire v_1659;
wire v_1660;
wire v_1661;
wire v_1662;
wire v_1663;
wire v_1664;
wire v_1665;
wire v_1666;
wire v_1667;
wire v_1668;
wire v_1669;
wire v_1670;
wire v_1671;
wire v_1672;
wire v_1673;
wire v_1674;
wire v_1675;
wire v_1676;
wire v_1677;
wire v_1678;
wire v_1679;
wire v_1680;
wire v_1681;
wire v_1682;
wire v_1683;
wire v_1684;
wire v_1685;
wire v_1686;
wire v_1687;
wire v_1688;
wire v_1689;
wire v_1690;
wire v_1691;
wire v_1692;
wire v_1693;
wire v_1694;
wire v_1695;
wire v_1696;
wire v_1697;
wire v_1698;
wire v_1699;
wire v_1700;
wire v_1701;
wire v_1702;
wire v_1703;
wire v_1704;
wire v_1705;
wire v_1706;
wire v_1707;
wire v_1708;
wire x_1;
assign v_1644 = 1;
assign v_5 = ~v_1 & ~v_2 & v_3 & v_4;
assign v_7 = ~v_1 & v_4 & v_6;
assign v_9 = ~v_1 & v_4 & v_8;
assign v_11 = v_2 & v_4 & ~v_10;
assign v_14 = ~v_1 & v_2 & v_4 & ~v_12 & ~v_13;
assign v_16 = ~v_1 & v_2 & v_4 & ~v_13 & ~v_15;
assign v_18 = ~v_1 & v_2 & v_4 & ~v_17;
assign v_19 = ~v_1 & v_4 & v_10 & ~v_17;
assign v_21 = ~v_1 & v_4 & v_10 & ~v_20;
assign v_22 = ~v_1 & v_4 & ~v_10 & v_17;
assign v_24 = ~v_1 & v_4 & v_23;
assign v_26 = v_25;
assign v_27 = v_4 & ~v_8 & ~v_10 & v_20;
assign v_28 = v_4 & v_8 & ~v_12 & v_13;
assign v_29 = v_4 & v_8 & v_13 & ~v_15;
assign v_30 = v_4 & v_6 & ~v_10;
assign v_31 = v_4 & v_6 & v_13;
assign v_32 = v_4 & v_6 & v_20;
assign v_34 = v_4 & v_33;
assign v_35 = v_4 & v_6 & v_17;
assign v_36 = v_4 & v_8 & v_17;
assign v_37 = v_4 & v_8 & v_13 & ~v_20;
assign v_38 = v_4 & v_8 & ~v_10 & ~v_20;
assign v_39 = v_4 & ~v_10 & v_23;
assign v_40 = ~v_2 & v_4 & ~v_8 & v_10 & v_13;
assign v_41 = v_3 & v_4 & ~v_10;
assign v_42 = ~v_2 & v_4 & v_12 & v_13 & v_17;
assign v_43 = ~v_2 & v_4 & v_13 & ~v_15 & v_17;
assign v_45 = v_4 & v_44;
assign v_46 = v_4 & v_17 & v_23;
assign v_47 = ~v_2 & v_3 & v_4 & v_17;
assign v_48 = ~v_2 & v_4 & ~v_8 & ~v_12 & v_20;
assign v_49 = v_1 & ~v_2 & v_4 & ~v_8 & v_20;
assign v_50 = ~v_1 & ~v_2 & v_4 & v_10 & ~v_15;
assign v_51 = v_1 & v_2 & v_4 & ~v_13 & v_17;
assign v_52 = v_1 & v_2 & v_4 & ~v_13 & v_20;
assign v_53 = v_2 & v_4 & v_13 & ~v_17;
assign v_54 = ~v_1 & v_3 & v_4 & ~v_13;
assign v_55 = v_3 & v_4 & v_8 & v_13;
assign v_56 = v_4 & v_13 & v_23;
assign v_57 = v_4 & v_8 & v_10 & ~v_13 & v_20;
assign v_58 = v_3 & v_4 & v_13 & ~v_20;
assign v_59 = v_2 & v_4 & v_13 & ~v_20;
assign v_63 = v_3 & v_4;
assign v_79 = v_63 & v_78;
assign v_80 = v_64 & ~v_65;
assign v_81 = ~v_67 & v_80;
assign v_82 = ~v_69 & ~v_70;
assign v_83 = ~v_72 & v_82;
assign v_84 = ~v_74 & v_83;
assign v_85 = v_76 & v_84;
assign v_86 = v_81 & v_85;
assign v_88 = v_86 & v_87;
assign v_94 = v_92 & v_93;
assign v_98 = v_4 & v_97;
assign v_99 = v_78 & v_98;
assign v_101 = v_86 & v_100;
assign v_107 = v_105 & v_106;
assign v_111 = v_4 & v_110;
assign v_112 = v_78 & v_111;
assign v_114 = v_86 & v_113;
assign v_120 = v_118 & v_119;
assign v_124 = v_4 & v_123;
assign v_127 = v_124 & v_126;
assign v_128 = v_72 & v_82;
assign v_129 = ~v_74 & v_128;
assign v_131 = v_129 & v_130;
assign v_137 = v_135 & v_136;
assign v_141 = v_4 & v_140;
assign v_142 = v_126 & v_141;
assign v_144 = v_129 & v_143;
assign v_150 = v_148 & v_149;
assign v_154 = v_4 & v_153;
assign v_155 = v_126 & v_154;
assign v_157 = v_129 & v_156;
assign v_163 = v_161 & v_162;
assign v_167 = v_4 & v_166;
assign v_168 = v_126 & v_167;
assign v_170 = v_129 & v_169;
assign v_176 = v_174 & v_175;
assign v_180 = v_4 & v_179;
assign v_181 = v_126 & v_180;
assign v_183 = v_129 & v_182;
assign v_189 = v_187 & v_188;
assign v_192 = v_4 & v_12;
assign v_196 = v_192 & v_195;
assign v_197 = ~v_64 & v_65;
assign v_198 = ~v_67 & v_197;
assign v_199 = v_85 & v_198;
assign v_200 = v_87 & v_199;
assign v_206 = v_204 & v_205;
assign v_209 = v_4 & v_15;
assign v_210 = v_195 & v_209;
assign v_211 = v_100 & v_199;
assign v_217 = v_215 & v_216;
assign v_221 = v_4 & v_220;
assign v_222 = v_126 & v_221;
assign v_224 = v_129 & v_223;
assign v_230 = v_228 & v_229;
assign v_234 = v_4 & v_233;
assign v_235 = v_126 & v_234;
assign v_237 = v_129 & v_236;
assign v_243 = v_241 & v_242;
assign v_247 = v_4 & v_246;
assign v_248 = v_126 & v_247;
assign v_250 = v_129 & v_249;
assign v_256 = v_254 & v_255;
assign v_260 = v_4 & v_259;
assign v_261 = v_126 & v_260;
assign v_263 = v_129 & v_262;
assign v_269 = v_267 & v_268;
assign v_273 = v_4 & v_272;
assign v_274 = v_126 & v_273;
assign v_276 = v_129 & v_275;
assign v_282 = v_280 & v_281;
assign v_286 = v_4 & v_285;
assign v_287 = v_126 & v_286;
assign v_289 = v_129 & v_288;
assign v_295 = v_293 & v_294;
assign v_298 = v_4 & v_8;
assign v_301 = v_2 & v_4;
assign v_306 = v_4 & v_6;
assign v_311 = v_304 & v_310;
assign v_317 = v_311 & v_316;
assign v_326 = v_306 & v_325;
assign v_327 = v_321 & v_326;
assign v_328 = v_63 & v_98;
assign v_329 = v_111 & v_328;
assign v_330 = v_192 & v_209;
assign v_331 = v_299 & v_305;
assign v_332 = v_313 & v_331;
assign v_333 = ~v_69 & v_70;
assign v_334 = ~v_72 & v_333;
assign v_335 = v_74 & v_334;
assign v_336 = v_332 & v_335;
assign v_337 = v_330 & v_336;
assign v_338 = v_329 & v_337;
assign v_340 = v_192 & v_214;
assign v_341 = v_336 & v_340;
assign v_344 = v_305 & v_306;
assign v_345 = v_313 & v_344;
assign v_346 = v_303 & v_345;
assign v_347 = v_298 & v_299;
assign v_348 = v_313 & v_347;
assign v_349 = v_309 & v_348;
assign v_351 = v_301 & v_331;
assign v_352 = v_315 & v_351;
assign v_354 = v_335 & v_353;
assign v_355 = v_315 & v_335;
assign v_356 = v_298 & v_306;
assign v_357 = v_313 & v_356;
assign v_358 = v_355 & v_357;
assign v_368 = v_360 & v_367;
assign v_371 = v_368 & v_370;
assign v_374 = v_203 & v_209;
assign v_375 = v_336 & v_374;
assign v_377 = v_298 & v_321;
assign v_378 = v_325 & v_377;
assign v_383 = v_367 & v_382;
assign v_386 = v_383 & v_385;
assign v_390 = v_301 & v_389;
assign v_392 = v_383 & v_391;
assign v_394 = v_331 & v_355;
assign v_396 = v_366 & v_395;
assign v_401 = v_4 & v_400;
assign v_405 = v_401 & v_404;
assign v_406 = v_69 & ~v_70;
assign v_407 = ~v_72 & v_406;
assign v_408 = ~v_74 & v_407;
assign v_410 = v_408 & v_409;
assign v_416 = v_414 & v_415;
assign v_420 = v_4 & v_419;
assign v_421 = v_404 & v_420;
assign v_423 = v_408 & v_422;
assign v_429 = v_427 & v_428;
assign v_433 = v_4 & v_432;
assign v_434 = v_404 & v_433;
assign v_436 = v_408 & v_435;
assign v_442 = v_440 & v_441;
assign v_446 = v_4 & v_445;
assign v_447 = v_404 & v_446;
assign v_449 = v_408 & v_448;
assign v_455 = v_453 & v_454;
assign v_459 = v_4 & v_458;
assign v_460 = v_404 & v_459;
assign v_462 = v_408 & v_461;
assign v_468 = v_466 & v_467;
assign v_472 = v_4 & v_471;
assign v_473 = v_404 & v_472;
assign v_475 = v_408 & v_474;
assign v_481 = v_479 & v_480;
assign v_485 = v_4 & v_484;
assign v_486 = v_126 & v_485;
assign v_488 = v_129 & v_487;
assign v_494 = v_492 & v_493;
assign v_498 = v_4 & v_497;
assign v_499 = v_126 & v_498;
assign v_501 = v_129 & v_500;
assign v_507 = v_505 & v_506;
assign v_511 = v_4 & v_510;
assign v_512 = v_126 & v_511;
assign v_514 = v_129 & v_513;
assign v_520 = v_518 & v_519;
assign v_524 = v_4 & v_523;
assign v_528 = v_524 & v_527;
assign v_530 = v_4 & v_529;
assign v_531 = v_64 & v_65;
assign v_532 = ~v_67 & v_531;
assign v_533 = v_85 & v_532;
assign v_534 = v_530 & v_533;
assign v_541 = v_538 & v_540;
assign v_545 = v_4 & v_544;
assign v_546 = v_527 & v_545;
assign v_548 = v_4 & v_547;
assign v_549 = v_533 & v_548;
assign v_556 = v_553 & v_555;
assign v_560 = v_4 & v_559;
assign v_561 = v_527 & v_560;
assign v_563 = v_4 & v_562;
assign v_564 = v_533 & v_563;
assign v_571 = v_568 & v_570;
assign v_581 = v_4 & v_580;
assign v_585 = v_581 & v_584;
assign v_587 = v_4 & v_586;
assign v_588 = ~v_64 & ~v_65;
assign v_589 = v_67 & v_588;
assign v_590 = v_85 & v_589;
assign v_591 = v_587 & v_590;
assign v_598 = v_595 & v_597;
assign v_602 = v_4 & v_601;
assign v_603 = v_584 & v_602;
assign v_605 = v_4 & v_604;
assign v_606 = v_590 & v_605;
assign v_613 = v_610 & v_612;
assign v_617 = v_4 & v_616;
assign v_618 = v_584 & v_617;
assign v_620 = v_4 & v_619;
assign v_621 = v_590 & v_620;
assign v_628 = v_625 & v_627;
assign v_632 = v_4 & v_631;
assign v_636 = v_4 & v_633;
assign v_638 = v_635 & v_637;
assign v_642 = v_4 & v_639;
assign v_644 = v_641 & v_643;
assign v_645 = v_638 & v_644;
assign v_649 = v_4 & v_646;
assign v_651 = v_648 & v_650;
assign v_652 = v_645 & v_651;
assign v_656 = v_4 & v_655;
assign v_657 = v_654 & v_656;
assign v_660 = v_657 & v_659;
assign v_661 = v_4 & v_658;
assign v_662 = v_4 & v_653;
assign v_664 = v_662 & v_663;
assign v_665 = v_661 & v_664;
assign v_669 = v_666 & v_668;
assign v_672 = v_670 & v_671;
assign v_675 = v_673 & v_674;
assign v_676 = v_672 & v_675;
assign v_679 = v_677 & v_678;
assign v_680 = v_676 & v_679;
assign v_681 = v_669 & v_680;
assign v_682 = v_652 & v_681;
assign v_683 = v_632 & v_682;
assign v_685 = v_683 & v_684;
assign v_687 = v_4 & v_686;
assign v_690 = v_687 & v_689;
assign v_691 = v_685 & v_690;
assign v_696 = v_4 & v_688;
assign v_697 = v_695 & v_696;
assign v_702 = v_698 & v_701;
assign v_704 = v_4 & v_703;
assign v_706 = v_696 & v_705;
assign v_707 = ~v_67 & v_588;
assign v_708 = ~v_76 & v_84;
assign v_709 = v_707 & v_708;
assign v_710 = v_706 & v_709;
assign v_714 = v_465 & v_636;
assign v_715 = v_459 & v_634;
assign v_717 = v_452 & v_642;
assign v_718 = v_446 & v_640;
assign v_721 = v_478 & v_649;
assign v_722 = v_472 & v_647;
assign v_729 = v_726 & v_728;
assign v_730 = v_4 & v_667;
assign v_732 = v_98 & v_426;
assign v_733 = v_104 & v_420;
assign v_735 = v_63 & v_413;
assign v_736 = v_91 & v_401;
assign v_739 = v_111 & v_439;
assign v_740 = v_117 & v_433;
assign v_749 = v_687 & v_696;
assign v_750 = v_694 & v_749;
assign v_752 = v_748 & v_751;
assign v_755 = v_87 & v_754;
assign v_758 = v_753 & v_757;
assign v_761 = v_695 & v_749;
assign v_763 = v_701 & v_762;
assign v_765 = v_709 & v_764;
assign v_769 = v_747 & v_768;
assign v_771 = v_692 & v_705;
assign v_773 = v_770 & v_772;
assign v_776 = v_78 & v_642;
assign v_777 = v_63 & v_86;
assign v_782 = v_780 & v_781;
assign v_785 = v_78 & v_636;
assign v_786 = v_86 & v_98;
assign v_791 = v_789 & v_790;
assign v_794 = v_78 & v_649;
assign v_795 = v_86 & v_111;
assign v_800 = v_798 & v_799;
assign v_804 = v_4 & v_803;
assign v_805 = v_126 & v_804;
assign v_807 = v_129 & v_806;
assign v_813 = v_811 & v_812;
assign v_817 = v_4 & v_816;
assign v_818 = v_126 & v_817;
assign v_820 = v_129 & v_819;
assign v_826 = v_824 & v_825;
assign v_830 = v_4 & v_829;
assign v_831 = v_126 & v_830;
assign v_833 = v_129 & v_832;
assign v_839 = v_837 & v_838;
assign v_842 = v_69 & v_70;
assign v_843 = v_72 & v_842;
assign v_844 = ~v_74 & v_843;
assign v_847 = v_845 & v_846;
assign v_849 = v_847 & v_848;
assign v_850 = v_4 & v_33;
assign v_851 = v_849 & v_850;
assign v_852 = v_844 & v_851;
assign v_853 = v_72 & v_406;
assign v_854 = ~v_74 & v_853;
assign v_855 = v_4 & v_10;
assign v_856 = v_1 & v_4;
assign v_857 = v_855 & v_856;
assign v_858 = v_4 & v_44;
assign v_859 = v_857 & v_858;
assign v_861 = v_859 & v_860;
assign v_862 = v_854 & v_861;
assign v_864 = v_72 & v_333;
assign v_865 = ~v_74 & v_864;
assign v_866 = v_846 & v_855;
assign v_867 = v_858 & v_866;
assign v_868 = v_860 & v_867;
assign v_869 = v_865 & v_868;
assign v_879 = v_871 & v_878;
assign v_881 = v_4 & v_880;
assign v_885 = v_882 & v_884;
assign v_887 = v_4 & v_886;
assign v_891 = v_888 & v_890;
assign v_892 = v_885 & v_891;
assign v_896 = v_4 & v_893;
assign v_898 = v_895 & v_897;
assign v_902 = v_4 & v_899;
assign v_904 = v_901 & v_903;
assign v_905 = v_898 & v_904;
assign v_909 = v_4 & v_906;
assign v_911 = v_908 & v_910;
assign v_912 = v_905 & v_911;
assign v_915 = v_913 & v_914;
assign v_918 = v_916 & v_917;
assign v_919 = v_915 & v_918;
assign v_922 = v_920 & v_921;
assign v_923 = v_919 & v_922;
assign v_925 = v_4 & v_924;
assign v_929 = v_926 & v_928;
assign v_931 = v_4 & v_930;
assign v_935 = v_932 & v_934;
assign v_936 = v_929 & v_935;
assign v_938 = v_4 & v_937;
assign v_942 = v_939 & v_941;
assign v_943 = v_936 & v_942;
assign v_947 = v_4 & v_946;
assign v_949 = v_4 & v_944;
assign v_952 = v_948 & v_951;
assign v_956 = v_4 & v_955;
assign v_958 = v_4 & v_953;
assign v_961 = v_957 & v_960;
assign v_962 = v_952 & v_961;
assign v_966 = v_4 & v_965;
assign v_968 = v_4 & v_963;
assign v_971 = v_967 & v_970;
assign v_972 = v_962 & v_971;
assign v_975 = v_973 & v_974;
assign v_978 = v_976 & v_977;
assign v_979 = v_975 & v_978;
assign v_982 = v_980 & v_981;
assign v_983 = v_979 & v_982;
assign v_986 = v_984 & v_985;
assign v_989 = v_987 & v_988;
assign v_990 = v_986 & v_989;
assign v_993 = v_991 & v_992;
assign v_994 = v_990 & v_993;
assign v_998 = v_4 & v_995;
assign v_1000 = v_997 & v_999;
assign v_1004 = v_4 & v_1001;
assign v_1006 = v_1003 & v_1005;
assign v_1007 = v_1000 & v_1006;
assign v_1011 = v_4 & v_1008;
assign v_1013 = v_1010 & v_1012;
assign v_1014 = v_1007 & v_1013;
assign v_1017 = v_1015 & v_1016;
assign v_1020 = v_1018 & v_1019;
assign v_1021 = v_1017 & v_1020;
assign v_1024 = v_1022 & v_1023;
assign v_1025 = v_1021 & v_1024;
assign v_1026 = v_1014 & v_1025;
assign v_1027 = v_994 & v_1026;
assign v_1028 = v_983 & v_1027;
assign v_1029 = v_972 & v_1028;
assign v_1030 = v_943 & v_1029;
assign v_1031 = v_923 & v_1030;
assign v_1032 = v_912 & v_1031;
assign v_1033 = v_892 & v_1032;
assign v_1034 = v_661 & v_1033;
assign v_1037 = v_879 & v_1036;
assign v_1038 = v_847 & v_858;
assign v_1039 = v_860 & v_1038;
assign v_1040 = v_750 & v_1039;
assign v_1041 = ~v_876 & v_1040;
assign v_1042 = v_335 & v_1041;
assign v_1044 = v_659 & v_1033;
assign v_1051 = v_1043 & v_1050;
assign v_1058 = v_1051 & v_1057;
assign v_1059 = v_848 & v_866;
assign v_1060 = v_860 & v_1059;
assign v_1061 = v_352 & v_1060;
assign v_1062 = v_335 & v_1061;
assign v_1068 = v_1063 & v_1067;
assign v_1069 = ~v_72 & v_842;
assign v_1070 = ~v_74 & v_1069;
assign v_1071 = v_849 & v_860;
assign v_1072 = v_1070 & v_1071;
assign v_1086 = v_1080 & v_1085;
assign v_1093 = v_1086 & v_1092;
assign v_1094 = v_846 & v_1093;
assign v_1095 = v_845 & v_856;
assign v_1096 = v_858 & v_1095;
assign v_1097 = v_860 & v_1096;
assign v_1098 = v_750 & v_1097;
assign v_1099 = v_876 & v_1098;
assign v_1100 = v_335 & v_1099;
assign v_1102 = v_180 & v_883;
assign v_1103 = v_186 & v_881;
assign v_1105 = v_167 & v_889;
assign v_1106 = v_173 & v_887;
assign v_1109 = v_634 & v_896;
assign v_1110 = v_636 & v_894;
assign v_1112 = v_640 & v_902;
assign v_1113 = v_642 & v_900;
assign v_1116 = v_647 & v_909;
assign v_1117 = v_649 & v_907;
assign v_1120 = v_104 & v_234;
assign v_1121 = v_98 & v_240;
assign v_1123 = v_91 & v_221;
assign v_1124 = v_63 & v_227;
assign v_1127 = v_117 & v_247;
assign v_1128 = v_111 & v_253;
assign v_1131 = v_498 & v_927;
assign v_1132 = v_504 & v_925;
assign v_1134 = v_485 & v_933;
assign v_1135 = v_491 & v_931;
assign v_1138 = v_511 & v_940;
assign v_1139 = v_517 & v_938;
assign v_1142 = v_949 & v_950;
assign v_1143 = v_945 & v_947;
assign v_1145 = v_958 & v_959;
assign v_1146 = v_954 & v_956;
assign v_1149 = v_968 & v_969;
assign v_1150 = v_964 & v_966;
assign v_1153 = v_141 & v_609;
assign v_1154 = v_147 & v_602;
assign v_1156 = v_124 & v_594;
assign v_1157 = v_134 & v_581;
assign v_1160 = v_154 & v_624;
assign v_1161 = v_160 & v_617;
assign v_1164 = v_611 & v_817;
assign v_1165 = v_605 & v_823;
assign v_1167 = v_596 & v_804;
assign v_1168 = v_587 & v_810;
assign v_1171 = v_626 & v_830;
assign v_1172 = v_620 & v_836;
assign v_1175 = v_552 & v_998;
assign v_1176 = v_545 & v_996;
assign v_1178 = v_537 & v_1004;
assign v_1179 = v_524 & v_1002;
assign v_1182 = v_567 & v_1011;
assign v_1183 = v_560 & v_1009;
assign v_1186 = v_273 & v_554;
assign v_1187 = v_279 & v_548;
assign v_1189 = v_260 & v_539;
assign v_1190 = v_266 & v_530;
assign v_1193 = v_286 & v_569;
assign v_1194 = v_292 & v_563;
assign v_1206 = v_1098 & v_1205;
assign v_1207 = v_335 & v_1206;
assign v_1211 = v_1208 & v_1210;
assign v_1213 = v_1040 & v_1212;
assign v_1214 = v_335 & v_1213;
assign v_1216 = v_848 & v_857;
assign v_1217 = v_860 & v_1216;
assign v_1218 = v_129 & v_1217;
assign v_1219 = ~v_1056 & v_1218;
assign v_1225 = v_1220 & v_1224;
assign v_1226 = v_848 & v_1095;
assign v_1227 = v_860 & v_1226;
assign v_1228 = v_349 & v_1227;
assign v_1229 = v_335 & v_1228;
assign v_1235 = v_1230 & v_1234;
assign v_1238 = v_335 & v_1040;
assign v_1239 = v_74 & v_83;
assign v_1240 = v_850 & v_1226;
assign v_1241 = v_1239 & v_1240;
assign v_1246 = v_1055 & v_1245;
assign v_1253 = v_845 & v_1252;
assign v_1254 = v_1093 & v_1253;
assign v_1255 = v_1036 & v_1254;
assign v_1256 = v_1249 & v_1255;
assign v_1258 = v_1067 & v_1257;
assign v_1262 = v_858 & v_1093;
assign v_1263 = v_1261 & v_1262;
assign v_1264 = v_1050 & v_1263;
assign v_1267 = v_335 & v_1098;
assign v_1271 = v_1055 & v_1270;
assign v_1274 = v_850 & v_1252;
assign v_1275 = v_1093 & v_1274;
assign v_1281 = v_1261 & v_1280;
assign v_1282 = v_1050 & v_1281;
assign v_1285 = v_404 & v_887;
assign v_1287 = v_408 & v_1286;
assign v_1292 = v_1290 & v_1291;
assign v_1295 = v_404 & v_881;
assign v_1297 = v_408 & v_1296;
assign v_1302 = v_1300 & v_1301;
assign v_1305 = v_126 & v_902;
assign v_1307 = v_129 & v_1306;
assign v_1312 = v_1310 & v_1311;
assign v_1315 = v_126 & v_896;
assign v_1317 = v_129 & v_1316;
assign v_1322 = v_1320 & v_1321;
assign v_1325 = v_126 & v_909;
assign v_1327 = v_129 & v_1326;
assign v_1332 = v_1330 & v_1331;
assign v_1335 = v_126 & v_958;
assign v_1337 = v_129 & v_1336;
assign v_1342 = v_1340 & v_1341;
assign v_1345 = v_126 & v_949;
assign v_1347 = v_129 & v_1346;
assign v_1352 = v_1350 & v_1351;
assign v_1355 = v_126 & v_968;
assign v_1357 = v_129 & v_1356;
assign v_1362 = v_1360 & v_1361;
assign v_1369 = v_1054 & v_1368;
assign v_1371 = v_4 & v_13;
assign v_1377 = v_4 & v_17;
assign v_1379 = v_1376 & v_1378;
assign v_1380 = v_1054 & v_1379;
assign v_1382 = v_1371 & v_1377;
assign v_1383 = v_1368 & v_1375;
assign v_1388 = v_4 & v_20;
assign v_1392 = v_1389 & v_1391;
assign v_1393 = v_1054 & v_1392;
assign v_1395 = v_1376 & v_1390;
assign v_1396 = v_1382 & v_1388;
assign v_1401 = v_4 & v_23;
assign v_1402 = v_1391 & v_1401;
assign v_1404 = v_1396 & v_1403;
assign v_1406 = v_1054 & v_1405;
assign v_1410 = v_1408 & v_1409;
assign v_1416 = v_662 & v_1415;
assign v_1417 = v_67 & v_531;
assign v_1418 = v_85 & v_1417;
assign v_1419 = v_87 & v_1418;
assign v_1424 = v_1422 & v_1423;
assign v_1427 = v_656 & v_1415;
assign v_1428 = v_100 & v_1418;
assign v_1433 = v_1431 & v_1432;
assign v_1436 = v_730 & v_1415;
assign v_1437 = v_113 & v_1418;
assign v_1442 = v_1440 & v_1441;
assign v_1445 = v_126 & v_1004;
assign v_1447 = v_129 & v_1446;
assign v_1452 = v_1450 & v_1451;
assign v_1455 = v_126 & v_998;
assign v_1457 = v_129 & v_1456;
assign v_1462 = v_1460 & v_1461;
assign v_1465 = v_126 & v_1011;
assign v_1467 = v_129 & v_1466;
assign v_1472 = v_1470 & v_1471;
assign v_1477 = v_956 & v_1476;
assign v_1478 = v_67 & v_197;
assign v_1479 = v_85 & v_1478;
assign v_1480 = v_87 & v_1479;
assign v_1485 = v_1483 & v_1484;
assign v_1488 = v_947 & v_1476;
assign v_1489 = v_100 & v_1479;
assign v_1494 = v_1492 & v_1493;
assign v_1497 = v_966 & v_1476;
assign v_1498 = v_113 & v_1479;
assign v_1503 = v_1501 & v_1502;
assign v_1506 = v_931 & v_1476;
assign v_1507 = v_956 & v_1479;
assign v_1512 = v_1510 & v_1511;
assign v_1515 = v_925 & v_1476;
assign v_1516 = v_947 & v_1479;
assign v_1521 = v_1519 & v_1520;
assign v_1524 = v_938 & v_1476;
assign v_1525 = v_966 & v_1479;
assign v_1530 = v_1528 & v_1529;
assign v_1533 = v_527 & v_530;
assign v_1534 = v_87 & v_533;
assign v_1539 = v_1537 & v_1538;
assign v_1542 = v_527 & v_548;
assign v_1543 = v_100 & v_533;
assign v_1548 = v_1546 & v_1547;
assign v_1551 = v_527 & v_563;
assign v_1552 = v_113 & v_533;
assign v_1557 = v_1555 & v_1556;
assign v_1560 = v_584 & v_587;
assign v_1561 = v_87 & v_590;
assign v_1566 = v_1564 & v_1565;
assign v_1569 = v_584 & v_605;
assign v_1570 = v_100 & v_590;
assign v_1575 = v_1573 & v_1574;
assign v_1578 = v_584 & v_620;
assign v_1579 = v_113 & v_590;
assign v_1584 = v_1582 & v_1583;
assign v_1588 = v_74 & v_1587;
assign v_1590 = v_1401 & v_1589;
assign v_1593 = ~v_69 & ~v_72;
assign v_1595 = v_1383 & v_1390;
assign v_1597 = v_1594 & v_1596;
assign v_1610 = ~v_1586;
assign v_1642 = v_1654 & v_1655;
assign v_1643 = v_1696 & v_1697;
assign v_1645 = v_1599 & v_1600 & v_1601 & v_1602 & v_1603;
assign v_1646 = v_1604 & v_1605 & v_1606 & v_1607 & v_1608;
assign v_1647 = v_1609 & v_1610 & v_1611 & v_1612 & v_1613;
assign v_1648 = v_1614 & v_1615 & v_1616 & v_1617 & v_1618;
assign v_1649 = v_1619 & v_1620 & v_1621 & v_1622 & v_1623;
assign v_1650 = v_1624 & v_1625 & v_1626 & v_1627 & v_1628;
assign v_1651 = v_1629 & v_1630 & v_1631 & v_1632 & v_1633;
assign v_1652 = v_1634 & v_1635 & v_1636 & v_1637 & v_1638;
assign v_1653 = v_1639 & v_1640 & v_1641;
assign v_1654 = v_1645 & v_1646 & v_1647 & v_1648 & v_1649;
assign v_1655 = v_1650 & v_1651 & v_1652 & v_1653;
assign v_1656 = v_61 & v_90 & v_95 & v_103 & v_108;
assign v_1657 = v_116 & v_121 & v_133 & v_138 & v_146;
assign v_1658 = v_151 & v_159 & v_164 & v_172 & v_177;
assign v_1659 = v_185 & v_190 & v_202 & v_207 & v_213;
assign v_1660 = v_218 & v_226 & v_231 & v_239 & v_244;
assign v_1661 = v_252 & v_257 & v_265 & v_270 & v_278;
assign v_1662 = v_283 & v_291 & v_296 & v_343 & v_372;
assign v_1663 = v_380 & v_387 & v_393 & v_398 & v_412;
assign v_1664 = v_417 & v_425 & v_430 & v_438 & v_443;
assign v_1665 = v_451 & v_456 & v_464 & v_469 & v_477;
assign v_1666 = v_482 & v_490 & v_495 & v_503 & v_508;
assign v_1667 = v_516 & v_521 & v_536 & v_542 & v_551;
assign v_1668 = v_557 & v_566 & v_572 & v_574 & v_575;
assign v_1669 = v_577 & v_578 & v_593 & v_599 & v_608;
assign v_1670 = v_614 & v_623 & v_629 & v_712 & v_759;
assign v_1671 = v_767 & v_774 & v_779 & v_783 & v_788;
assign v_1672 = v_792 & v_797 & v_801 & v_809 & v_814;
assign v_1673 = v_822 & v_827 & v_835 & v_840 & v_1074;
assign v_1674 = v_1236 & v_1248 & v_1259 & v_1266 & v_1272;
assign v_1675 = v_1278 & v_1283 & v_1289 & v_1293 & v_1299;
assign v_1676 = v_1303 & v_1309 & v_1313 & v_1319 & v_1323;
assign v_1677 = v_1329 & v_1333 & v_1339 & v_1343 & v_1349;
assign v_1678 = v_1353 & v_1359 & v_1363 & v_1365 & v_1366;
assign v_1679 = v_1370 & v_1373 & v_1381 & v_1386 & v_1394;
assign v_1680 = v_1399 & v_1407 & v_1412 & v_1421 & v_1425;
assign v_1681 = v_1430 & v_1434 & v_1439 & v_1443 & v_1449;
assign v_1682 = v_1453 & v_1459 & v_1463 & v_1469 & v_1473;
assign v_1683 = v_1482 & v_1486 & v_1491 & v_1495 & v_1500;
assign v_1684 = v_1504 & v_1509 & v_1513 & v_1518 & v_1522;
assign v_1685 = v_1527 & v_1531 & v_1536 & v_1540 & v_1545;
assign v_1686 = v_1549 & v_1554 & v_1558 & v_1563 & v_1567;
assign v_1687 = v_1572 & v_1576 & v_1581 & v_1585 & v_1592;
assign v_1688 = v_1598 & v_1642;
assign v_1689 = v_1656 & v_1657 & v_1658 & v_1659 & v_1660;
assign v_1690 = v_1661 & v_1662 & v_1663 & v_1664 & v_1665;
assign v_1691 = v_1666 & v_1667 & v_1668 & v_1669 & v_1670;
assign v_1692 = v_1671 & v_1672 & v_1673 & v_1674 & v_1675;
assign v_1693 = v_1676 & v_1677 & v_1678 & v_1679 & v_1680;
assign v_1694 = v_1681 & v_1682 & v_1683 & v_1684 & v_1685;
assign v_1695 = v_1686 & v_1687 & v_1688;
assign v_1696 = v_1689 & v_1690 & v_1691 & v_1692 & v_1693;
assign v_1697 = v_1694 & v_1695;
assign v_60 = v_1707 | v_1708;
assign v_66 = ~v_64 | v_65;
assign v_68 = v_66 | v_67;
assign v_71 = v_69 | v_70;
assign v_73 = v_71 | v_72;
assign v_75 = v_73 | v_74;
assign v_77 = v_75 | ~v_76;
assign v_78 = v_68 | v_77;
assign v_89 = v_79 | v_88;
assign v_90 = ~v_62 | v_89;
assign v_91 = ~v_3 | ~v_4;
assign v_92 = v_86 | v_91;
assign v_93 = v_78 | ~v_87;
assign v_95 = v_62 | v_94;
assign v_102 = v_99 | v_101;
assign v_103 = ~v_96 | v_102;
assign v_104 = ~v_4 | ~v_97;
assign v_105 = v_86 | v_104;
assign v_106 = v_78 | ~v_100;
assign v_108 = v_96 | v_107;
assign v_115 = v_112 | v_114;
assign v_116 = ~v_109 | v_115;
assign v_117 = ~v_4 | ~v_110;
assign v_118 = v_86 | v_117;
assign v_119 = v_78 | ~v_113;
assign v_121 = v_109 | v_120;
assign v_125 = v_71 | ~v_72;
assign v_126 = v_74 | v_125;
assign v_132 = v_127 | v_131;
assign v_133 = ~v_122 | v_132;
assign v_134 = ~v_4 | ~v_123;
assign v_135 = v_129 | v_134;
assign v_136 = v_126 | ~v_130;
assign v_138 = v_122 | v_137;
assign v_145 = v_142 | v_144;
assign v_146 = ~v_139 | v_145;
assign v_147 = ~v_4 | ~v_140;
assign v_148 = v_129 | v_147;
assign v_149 = v_126 | ~v_143;
assign v_151 = v_139 | v_150;
assign v_158 = v_155 | v_157;
assign v_159 = ~v_152 | v_158;
assign v_160 = ~v_4 | ~v_153;
assign v_161 = v_129 | v_160;
assign v_162 = v_126 | ~v_156;
assign v_164 = v_152 | v_163;
assign v_171 = v_168 | v_170;
assign v_172 = ~v_165 | v_171;
assign v_173 = ~v_4 | ~v_166;
assign v_174 = v_129 | v_173;
assign v_175 = v_126 | ~v_169;
assign v_177 = v_165 | v_176;
assign v_184 = v_181 | v_183;
assign v_185 = ~v_178 | v_184;
assign v_186 = ~v_4 | ~v_179;
assign v_187 = v_129 | v_186;
assign v_188 = v_126 | ~v_182;
assign v_190 = v_178 | v_189;
assign v_193 = v_64 | ~v_65;
assign v_194 = v_67 | v_193;
assign v_195 = v_77 | v_194;
assign v_201 = v_196 | v_200;
assign v_202 = ~v_191 | v_201;
assign v_203 = ~v_4 | ~v_12;
assign v_204 = v_199 | v_203;
assign v_205 = ~v_87 | v_195;
assign v_207 = v_191 | v_206;
assign v_212 = v_210 | v_211;
assign v_213 = ~v_208 | v_212;
assign v_214 = ~v_4 | ~v_15;
assign v_215 = v_199 | v_214;
assign v_216 = ~v_100 | v_195;
assign v_218 = v_208 | v_217;
assign v_225 = v_222 | v_224;
assign v_226 = ~v_219 | v_225;
assign v_227 = ~v_4 | ~v_220;
assign v_228 = v_129 | v_227;
assign v_229 = v_126 | ~v_223;
assign v_231 = v_219 | v_230;
assign v_238 = v_235 | v_237;
assign v_239 = ~v_232 | v_238;
assign v_240 = ~v_4 | ~v_233;
assign v_241 = v_129 | v_240;
assign v_242 = v_126 | ~v_236;
assign v_244 = v_232 | v_243;
assign v_251 = v_248 | v_250;
assign v_252 = ~v_245 | v_251;
assign v_253 = ~v_4 | ~v_246;
assign v_254 = v_129 | v_253;
assign v_255 = v_126 | ~v_249;
assign v_257 = v_245 | v_256;
assign v_264 = v_261 | v_263;
assign v_265 = ~v_258 | v_264;
assign v_266 = ~v_4 | ~v_259;
assign v_267 = v_129 | v_266;
assign v_268 = v_126 | ~v_262;
assign v_270 = v_258 | v_269;
assign v_277 = v_274 | v_276;
assign v_278 = ~v_271 | v_277;
assign v_279 = ~v_4 | ~v_272;
assign v_280 = v_129 | v_279;
assign v_281 = v_126 | ~v_275;
assign v_283 = v_271 | v_282;
assign v_290 = v_287 | v_289;
assign v_291 = ~v_284 | v_290;
assign v_292 = ~v_4 | ~v_285;
assign v_293 = v_129 | v_292;
assign v_294 = v_126 | ~v_288;
assign v_296 = v_284 | v_295;
assign v_299 = ~v_4 | ~v_6;
assign v_300 = v_298 | v_299;
assign v_302 = v_300 | v_301;
assign v_304 = v_302 | ~v_303;
assign v_305 = ~v_4 | ~v_8;
assign v_307 = v_305 | v_306;
assign v_308 = v_301 | v_307;
assign v_310 = v_308 | ~v_309;
assign v_312 = v_298 | v_306;
assign v_313 = ~v_2 | ~v_4;
assign v_314 = v_312 | v_313;
assign v_316 = v_314 | ~v_315;
assign v_318 = v_69 | ~v_70;
assign v_319 = v_72 | v_318;
assign v_320 = ~v_74 | v_319;
assign v_321 = v_317 | v_320;
assign v_322 = ~v_315 | v_320;
assign v_323 = v_299 | v_305;
assign v_324 = v_301 | v_323;
assign v_325 = v_322 | v_324;
assign v_339 = v_327 | v_338;
assign v_342 = v_339 | v_341;
assign v_343 = ~v_297 | v_342;
assign v_350 = v_346 | v_349;
assign v_353 = v_350 | v_352;
assign v_359 = v_299 | v_358;
assign v_360 = v_354 | v_359;
assign v_361 = v_91 | v_104;
assign v_362 = v_117 | v_361;
assign v_363 = v_203 | v_214;
assign v_364 = v_301 | v_312;
assign v_365 = v_320 | v_364;
assign v_366 = v_363 | v_365;
assign v_367 = v_362 | v_366;
assign v_369 = v_203 | v_209;
assign v_370 = v_365 | v_369;
assign v_372 = v_297 | v_371;
assign v_376 = v_338 | v_375;
assign v_379 = v_376 | v_378;
assign v_380 = ~v_373 | v_379;
assign v_381 = v_192 | v_214;
assign v_382 = v_365 | v_381;
assign v_384 = v_305 | v_354;
assign v_385 = v_358 | v_384;
assign v_387 = v_373 | v_386;
assign v_389 = v_312 | v_322;
assign v_391 = v_337 | v_390;
assign v_393 = ~v_388 | v_392;
assign v_395 = v_313 | v_394;
assign v_397 = v_376 | v_396;
assign v_398 = v_388 | v_397;
assign v_402 = ~v_69 | v_70;
assign v_403 = v_72 | v_402;
assign v_404 = v_74 | v_403;
assign v_411 = v_405 | v_410;
assign v_412 = ~v_399 | v_411;
assign v_413 = ~v_4 | ~v_400;
assign v_414 = v_408 | v_413;
assign v_415 = v_404 | ~v_409;
assign v_417 = v_399 | v_416;
assign v_424 = v_421 | v_423;
assign v_425 = ~v_418 | v_424;
assign v_426 = ~v_4 | ~v_419;
assign v_427 = v_408 | v_426;
assign v_428 = v_404 | ~v_422;
assign v_430 = v_418 | v_429;
assign v_437 = v_434 | v_436;
assign v_438 = ~v_431 | v_437;
assign v_439 = ~v_4 | ~v_432;
assign v_440 = v_408 | v_439;
assign v_441 = v_404 | ~v_435;
assign v_443 = v_431 | v_442;
assign v_450 = v_447 | v_449;
assign v_451 = ~v_444 | v_450;
assign v_452 = ~v_4 | ~v_445;
assign v_453 = v_408 | v_452;
assign v_454 = v_404 | ~v_448;
assign v_456 = v_444 | v_455;
assign v_463 = v_460 | v_462;
assign v_464 = ~v_457 | v_463;
assign v_465 = ~v_4 | ~v_458;
assign v_466 = v_408 | v_465;
assign v_467 = v_404 | ~v_461;
assign v_469 = v_457 | v_468;
assign v_476 = v_473 | v_475;
assign v_477 = ~v_470 | v_476;
assign v_478 = ~v_4 | ~v_471;
assign v_479 = v_408 | v_478;
assign v_480 = v_404 | ~v_474;
assign v_482 = v_470 | v_481;
assign v_489 = v_486 | v_488;
assign v_490 = ~v_483 | v_489;
assign v_491 = ~v_4 | ~v_484;
assign v_492 = v_129 | v_491;
assign v_493 = v_126 | ~v_487;
assign v_495 = v_483 | v_494;
assign v_502 = v_499 | v_501;
assign v_503 = ~v_496 | v_502;
assign v_504 = ~v_4 | ~v_497;
assign v_505 = v_129 | v_504;
assign v_506 = v_126 | ~v_500;
assign v_508 = v_496 | v_507;
assign v_515 = v_512 | v_514;
assign v_516 = ~v_509 | v_515;
assign v_517 = ~v_4 | ~v_510;
assign v_518 = v_129 | v_517;
assign v_519 = v_126 | ~v_513;
assign v_521 = v_509 | v_520;
assign v_525 = ~v_64 | ~v_65;
assign v_526 = v_67 | v_525;
assign v_527 = v_77 | v_526;
assign v_535 = v_528 | v_534;
assign v_536 = ~v_522 | v_535;
assign v_537 = ~v_4 | ~v_523;
assign v_538 = v_533 | v_537;
assign v_539 = ~v_4 | ~v_529;
assign v_540 = v_527 | v_539;
assign v_542 = v_522 | v_541;
assign v_550 = v_546 | v_549;
assign v_551 = ~v_543 | v_550;
assign v_552 = ~v_4 | ~v_544;
assign v_553 = v_533 | v_552;
assign v_554 = ~v_4 | ~v_547;
assign v_555 = v_527 | v_554;
assign v_557 = v_543 | v_556;
assign v_565 = v_561 | v_564;
assign v_566 = ~v_558 | v_565;
assign v_567 = ~v_4 | ~v_559;
assign v_568 = v_533 | v_567;
assign v_569 = ~v_4 | ~v_562;
assign v_570 = v_527 | v_569;
assign v_572 = v_558 | v_571;
assign v_574 = v_113 | ~v_573;
assign v_575 = ~v_113 | v_573;
assign v_577 = v_87 | ~v_576;
assign v_578 = ~v_87 | v_576;
assign v_582 = v_64 | v_65;
assign v_583 = ~v_67 | v_582;
assign v_584 = v_77 | v_583;
assign v_592 = v_585 | v_591;
assign v_593 = ~v_579 | v_592;
assign v_594 = ~v_4 | ~v_580;
assign v_595 = v_590 | v_594;
assign v_596 = ~v_4 | ~v_586;
assign v_597 = v_584 | v_596;
assign v_599 = v_579 | v_598;
assign v_607 = v_603 | v_606;
assign v_608 = ~v_600 | v_607;
assign v_609 = ~v_4 | ~v_601;
assign v_610 = v_590 | v_609;
assign v_611 = ~v_4 | ~v_604;
assign v_612 = v_584 | v_611;
assign v_614 = v_600 | v_613;
assign v_622 = v_618 | v_621;
assign v_623 = ~v_615 | v_622;
assign v_624 = ~v_4 | ~v_616;
assign v_625 = v_590 | v_624;
assign v_626 = ~v_4 | ~v_619;
assign v_627 = v_584 | v_626;
assign v_629 = v_615 | v_628;
assign v_634 = ~v_4 | ~v_633;
assign v_635 = v_459 | v_634;
assign v_637 = v_465 | v_636;
assign v_640 = ~v_4 | ~v_639;
assign v_641 = v_446 | v_640;
assign v_643 = v_452 | v_642;
assign v_647 = ~v_4 | ~v_646;
assign v_648 = v_472 | v_647;
assign v_650 = v_478 | v_649;
assign v_654 = ~v_4 | ~v_653;
assign v_659 = ~v_4 | ~v_658;
assign v_663 = ~v_4 | ~v_655;
assign v_666 = v_660 | v_665;
assign v_668 = ~v_4 | ~v_667;
assign v_670 = v_104 | v_420;
assign v_671 = v_98 | v_426;
assign v_673 = v_91 | v_401;
assign v_674 = v_63 | v_413;
assign v_677 = v_117 | v_433;
assign v_678 = v_111 | v_439;
assign v_689 = ~v_4 | ~v_688;
assign v_692 = ~v_4 | ~v_686;
assign v_693 = v_689 | v_692;
assign v_695 = v_693 | ~v_694;
assign v_698 = v_691 | v_697;
assign v_699 = v_67 | v_582;
assign v_700 = v_75 | v_76;
assign v_701 = v_699 | v_700;
assign v_705 = ~v_87 | v_704;
assign v_711 = v_702 | v_710;
assign v_712 = ~v_630 | v_711;
assign v_713 = ~v_4 | ~v_631;
assign v_716 = v_714 | v_715;
assign v_719 = v_717 | v_718;
assign v_720 = v_716 | v_719;
assign v_723 = v_721 | v_722;
assign v_724 = v_720 | v_723;
assign v_725 = v_662 | v_663;
assign v_726 = v_661 | v_725;
assign v_727 = v_654 | v_656;
assign v_728 = v_659 | v_727;
assign v_731 = v_729 | v_730;
assign v_734 = v_732 | v_733;
assign v_737 = v_735 | v_736;
assign v_738 = v_734 | v_737;
assign v_741 = v_739 | v_740;
assign v_742 = v_738 | v_741;
assign v_743 = v_731 | v_742;
assign v_744 = v_724 | v_743;
assign v_745 = v_713 | v_744;
assign v_746 = ~v_684 | v_745;
assign v_747 = v_692 | v_696;
assign v_748 = v_746 | v_747;
assign v_751 = v_689 | v_750;
assign v_753 = v_709 | v_752;
assign v_754 = ~v_4 | ~v_703;
assign v_756 = v_689 | v_755;
assign v_757 = v_701 | v_756;
assign v_759 = v_630 | v_758;
assign v_762 = v_690 | v_761;
assign v_764 = v_687 | v_755;
assign v_766 = v_763 | v_765;
assign v_767 = ~v_760 | v_766;
assign v_768 = v_693 | v_750;
assign v_770 = v_709 | v_769;
assign v_772 = v_701 | v_771;
assign v_774 = v_760 | v_773;
assign v_778 = v_776 | v_777;
assign v_779 = ~v_775 | v_778;
assign v_780 = v_86 | v_640;
assign v_781 = v_78 | v_91;
assign v_783 = v_775 | v_782;
assign v_787 = v_785 | v_786;
assign v_788 = ~v_784 | v_787;
assign v_789 = v_86 | v_634;
assign v_790 = v_78 | v_104;
assign v_792 = v_784 | v_791;
assign v_796 = v_794 | v_795;
assign v_797 = ~v_793 | v_796;
assign v_798 = v_86 | v_647;
assign v_799 = v_78 | v_117;
assign v_801 = v_793 | v_800;
assign v_808 = v_805 | v_807;
assign v_809 = ~v_802 | v_808;
assign v_810 = ~v_4 | ~v_803;
assign v_811 = v_129 | v_810;
assign v_812 = v_126 | ~v_806;
assign v_814 = v_802 | v_813;
assign v_821 = v_818 | v_820;
assign v_822 = ~v_815 | v_821;
assign v_823 = ~v_4 | ~v_816;
assign v_824 = v_129 | v_823;
assign v_825 = v_126 | ~v_819;
assign v_827 = v_815 | v_826;
assign v_834 = v_831 | v_833;
assign v_835 = ~v_828 | v_834;
assign v_836 = ~v_4 | ~v_829;
assign v_837 = v_129 | v_836;
assign v_838 = v_126 | ~v_832;
assign v_840 = v_828 | v_839;
assign v_845 = ~v_4 | ~v_10;
assign v_846 = ~v_1 | ~v_4;
assign v_848 = ~v_4 | ~v_44;
assign v_860 = ~v_4 | ~v_33;
assign v_863 = v_852 | v_862;
assign v_870 = v_863 | v_869;
assign v_871 = v_856 | v_870;
assign v_872 = v_846 | v_855;
assign v_873 = v_848 | v_872;
assign v_874 = v_850 | v_873;
assign v_875 = v_695 | v_874;
assign v_877 = v_875 | ~v_876;
assign v_878 = v_320 | v_877;
assign v_882 = v_186 | v_881;
assign v_883 = ~v_4 | ~v_880;
assign v_884 = v_180 | v_883;
assign v_888 = v_173 | v_887;
assign v_889 = ~v_4 | ~v_886;
assign v_890 = v_167 | v_889;
assign v_894 = ~v_4 | ~v_893;
assign v_895 = v_636 | v_894;
assign v_897 = v_634 | v_896;
assign v_900 = ~v_4 | ~v_899;
assign v_901 = v_642 | v_900;
assign v_903 = v_640 | v_902;
assign v_907 = ~v_4 | ~v_906;
assign v_908 = v_649 | v_907;
assign v_910 = v_647 | v_909;
assign v_913 = v_98 | v_240;
assign v_914 = v_104 | v_234;
assign v_916 = v_63 | v_227;
assign v_917 = v_91 | v_221;
assign v_920 = v_111 | v_253;
assign v_921 = v_117 | v_247;
assign v_926 = v_504 | v_925;
assign v_927 = ~v_4 | ~v_924;
assign v_928 = v_498 | v_927;
assign v_932 = v_491 | v_931;
assign v_933 = ~v_4 | ~v_930;
assign v_934 = v_485 | v_933;
assign v_939 = v_517 | v_938;
assign v_940 = ~v_4 | ~v_937;
assign v_941 = v_511 | v_940;
assign v_945 = ~v_4 | ~v_944;
assign v_948 = v_945 | v_947;
assign v_950 = ~v_4 | ~v_946;
assign v_951 = v_949 | v_950;
assign v_954 = ~v_4 | ~v_953;
assign v_957 = v_954 | v_956;
assign v_959 = ~v_4 | ~v_955;
assign v_960 = v_958 | v_959;
assign v_964 = ~v_4 | ~v_963;
assign v_967 = v_964 | v_966;
assign v_969 = ~v_4 | ~v_965;
assign v_970 = v_968 | v_969;
assign v_973 = v_147 | v_602;
assign v_974 = v_141 | v_609;
assign v_976 = v_134 | v_581;
assign v_977 = v_124 | v_594;
assign v_980 = v_160 | v_617;
assign v_981 = v_154 | v_624;
assign v_984 = v_605 | v_823;
assign v_985 = v_611 | v_817;
assign v_987 = v_587 | v_810;
assign v_988 = v_596 | v_804;
assign v_991 = v_620 | v_836;
assign v_992 = v_626 | v_830;
assign v_996 = ~v_4 | ~v_995;
assign v_997 = v_545 | v_996;
assign v_999 = v_552 | v_998;
assign v_1002 = ~v_4 | ~v_1001;
assign v_1003 = v_524 | v_1002;
assign v_1005 = v_537 | v_1004;
assign v_1009 = ~v_4 | ~v_1008;
assign v_1010 = v_560 | v_1009;
assign v_1012 = v_567 | v_1011;
assign v_1015 = v_279 | v_548;
assign v_1016 = v_273 | v_554;
assign v_1018 = v_266 | v_530;
assign v_1019 = v_260 | v_539;
assign v_1022 = v_292 | v_563;
assign v_1023 = v_286 | v_569;
assign v_1035 = v_875 | v_1034;
assign v_1036 = v_320 | v_1035;
assign v_1043 = v_1037 | v_1042;
assign v_1045 = v_855 | v_856;
assign v_1046 = v_848 | v_1045;
assign v_1047 = v_850 | v_1046;
assign v_1048 = v_695 | v_1047;
assign v_1049 = v_1044 | v_1048;
assign v_1050 = v_320 | v_1049;
assign v_1052 = v_845 | v_846;
assign v_1053 = v_858 | v_1052;
assign v_1054 = v_850 | v_1053;
assign v_1055 = v_126 | v_1054;
assign v_1057 = v_1055 | v_1056;
assign v_1063 = v_1058 | v_1062;
assign v_1064 = v_858 | v_872;
assign v_1065 = v_850 | v_1064;
assign v_1066 = v_310 | v_1065;
assign v_1067 = v_320 | v_1066;
assign v_1073 = v_1068 | v_1072;
assign v_1074 = ~v_841 | v_1073;
assign v_1075 = ~v_69 | ~v_70;
assign v_1076 = ~v_72 | v_1075;
assign v_1077 = v_74 | v_1076;
assign v_1078 = v_858 | v_1045;
assign v_1079 = v_860 | v_1078;
assign v_1080 = v_1077 | v_1079;
assign v_1081 = ~v_72 | v_402;
assign v_1082 = v_74 | v_1081;
assign v_1083 = v_848 | v_1052;
assign v_1084 = v_850 | v_1083;
assign v_1085 = v_1082 | v_1084;
assign v_1087 = ~v_72 | v_318;
assign v_1088 = v_74 | v_1087;
assign v_1089 = v_845 | v_856;
assign v_1090 = v_848 | v_1089;
assign v_1091 = v_850 | v_1090;
assign v_1092 = v_1088 | v_1091;
assign v_1101 = v_1094 | v_1100;
assign v_1104 = v_1102 | v_1103;
assign v_1107 = v_1105 | v_1106;
assign v_1108 = v_1104 | v_1107;
assign v_1111 = v_1109 | v_1110;
assign v_1114 = v_1112 | v_1113;
assign v_1115 = v_1111 | v_1114;
assign v_1118 = v_1116 | v_1117;
assign v_1119 = v_1115 | v_1118;
assign v_1122 = v_1120 | v_1121;
assign v_1125 = v_1123 | v_1124;
assign v_1126 = v_1122 | v_1125;
assign v_1129 = v_1127 | v_1128;
assign v_1130 = v_1126 | v_1129;
assign v_1133 = v_1131 | v_1132;
assign v_1136 = v_1134 | v_1135;
assign v_1137 = v_1133 | v_1136;
assign v_1140 = v_1138 | v_1139;
assign v_1141 = v_1137 | v_1140;
assign v_1144 = v_1142 | v_1143;
assign v_1147 = v_1145 | v_1146;
assign v_1148 = v_1144 | v_1147;
assign v_1151 = v_1149 | v_1150;
assign v_1152 = v_1148 | v_1151;
assign v_1155 = v_1153 | v_1154;
assign v_1158 = v_1156 | v_1157;
assign v_1159 = v_1155 | v_1158;
assign v_1162 = v_1160 | v_1161;
assign v_1163 = v_1159 | v_1162;
assign v_1166 = v_1164 | v_1165;
assign v_1169 = v_1167 | v_1168;
assign v_1170 = v_1166 | v_1169;
assign v_1173 = v_1171 | v_1172;
assign v_1174 = v_1170 | v_1173;
assign v_1177 = v_1175 | v_1176;
assign v_1180 = v_1178 | v_1179;
assign v_1181 = v_1177 | v_1180;
assign v_1184 = v_1182 | v_1183;
assign v_1185 = v_1181 | v_1184;
assign v_1188 = v_1186 | v_1187;
assign v_1191 = v_1189 | v_1190;
assign v_1192 = v_1188 | v_1191;
assign v_1195 = v_1193 | v_1194;
assign v_1196 = v_1192 | v_1195;
assign v_1197 = v_1185 | v_1196;
assign v_1198 = v_1174 | v_1197;
assign v_1199 = v_1163 | v_1198;
assign v_1200 = v_1152 | v_1199;
assign v_1201 = v_1141 | v_1200;
assign v_1202 = v_1130 | v_1201;
assign v_1203 = v_1119 | v_1202;
assign v_1204 = v_1108 | v_1203;
assign v_1205 = v_659 | v_1204;
assign v_1208 = v_1101 | v_1207;
assign v_1209 = v_876 | v_1048;
assign v_1210 = v_320 | v_1209;
assign v_1212 = v_661 | v_1204;
assign v_1215 = v_1211 | v_1214;
assign v_1220 = v_1215 | v_1219;
assign v_1221 = v_858 | v_1089;
assign v_1222 = v_850 | v_1221;
assign v_1223 = v_316 | v_1222;
assign v_1224 = v_320 | v_1223;
assign v_1230 = v_1225 | v_1229;
assign v_1231 = v_72 | v_1075;
assign v_1232 = v_74 | v_1231;
assign v_1233 = v_850 | v_1078;
assign v_1234 = v_1232 | v_1233;
assign v_1236 = v_841 | v_1235;
assign v_1242 = v_855 | v_1241;
assign v_1243 = v_870 | v_1242;
assign v_1244 = v_1207 | v_1243;
assign v_1245 = v_1238 | v_1244;
assign v_1247 = v_1229 | v_1246;
assign v_1248 = ~v_1237 | v_1247;
assign v_1249 = v_320 | v_1048;
assign v_1250 = v_73 | ~v_74;
assign v_1251 = v_860 | v_1064;
assign v_1252 = v_1250 | v_1251;
assign v_1257 = v_1218 | v_1256;
assign v_1259 = v_1237 | v_1258;
assign v_1261 = v_320 | v_875;
assign v_1265 = v_1218 | v_1264;
assign v_1266 = ~v_1260 | v_1265;
assign v_1268 = v_848 | v_870;
assign v_1269 = v_1267 | v_1268;
assign v_1270 = v_1214 | v_1269;
assign v_1272 = v_1260 | v_1271;
assign v_1276 = v_1267 | v_1275;
assign v_1277 = v_1214 | v_1276;
assign v_1278 = ~v_1273 | v_1277;
assign v_1279 = v_860 | v_1241;
assign v_1280 = v_870 | v_1279;
assign v_1283 = v_1273 | v_1282;
assign v_1288 = v_1285 | v_1287;
assign v_1289 = ~v_1284 | v_1288;
assign v_1290 = v_408 | v_889;
assign v_1291 = v_404 | ~v_1286;
assign v_1293 = v_1284 | v_1292;
assign v_1298 = v_1295 | v_1297;
assign v_1299 = ~v_1294 | v_1298;
assign v_1300 = v_408 | v_883;
assign v_1301 = v_404 | ~v_1296;
assign v_1303 = v_1294 | v_1302;
assign v_1308 = v_1305 | v_1307;
assign v_1309 = ~v_1304 | v_1308;
assign v_1310 = v_129 | v_900;
assign v_1311 = v_126 | ~v_1306;
assign v_1313 = v_1304 | v_1312;
assign v_1318 = v_1315 | v_1317;
assign v_1319 = ~v_1314 | v_1318;
assign v_1320 = v_129 | v_894;
assign v_1321 = v_126 | ~v_1316;
assign v_1323 = v_1314 | v_1322;
assign v_1328 = v_1325 | v_1327;
assign v_1329 = ~v_1324 | v_1328;
assign v_1330 = v_129 | v_907;
assign v_1331 = v_126 | ~v_1326;
assign v_1333 = v_1324 | v_1332;
assign v_1338 = v_1335 | v_1337;
assign v_1339 = ~v_1334 | v_1338;
assign v_1340 = v_129 | v_954;
assign v_1341 = v_126 | ~v_1336;
assign v_1343 = v_1334 | v_1342;
assign v_1348 = v_1345 | v_1347;
assign v_1349 = ~v_1344 | v_1348;
assign v_1350 = v_129 | v_945;
assign v_1351 = v_126 | ~v_1346;
assign v_1353 = v_1344 | v_1352;
assign v_1358 = v_1355 | v_1357;
assign v_1359 = ~v_1354 | v_1358;
assign v_1360 = v_129 | v_964;
assign v_1361 = v_126 | ~v_1356;
assign v_1363 = v_1354 | v_1362;
assign v_1365 = v_100 | ~v_1364;
assign v_1366 = ~v_100 | v_1364;
assign v_1368 = ~v_4 | ~v_13;
assign v_1370 = ~v_1367 | v_1369;
assign v_1372 = v_1217 | v_1371;
assign v_1373 = v_1367 | v_1372;
assign v_1375 = ~v_4 | ~v_17;
assign v_1376 = v_1368 | v_1375;
assign v_1378 = v_1371 | v_1377;
assign v_1381 = ~v_1374 | v_1380;
assign v_1384 = v_1382 | v_1383;
assign v_1385 = v_1217 | v_1384;
assign v_1386 = v_1374 | v_1385;
assign v_1389 = v_1382 | v_1388;
assign v_1390 = ~v_4 | ~v_20;
assign v_1391 = v_1376 | v_1390;
assign v_1394 = ~v_1387 | v_1393;
assign v_1397 = v_1395 | v_1396;
assign v_1398 = v_1217 | v_1397;
assign v_1399 = v_1387 | v_1398;
assign v_1403 = ~v_4 | ~v_23;
assign v_1405 = v_1402 | v_1404;
assign v_1407 = ~v_1400 | v_1406;
assign v_1408 = v_1396 | v_1403;
assign v_1409 = v_1391 | v_1401;
assign v_1411 = v_1217 | v_1410;
assign v_1412 = v_1400 | v_1411;
assign v_1414 = ~v_67 | v_525;
assign v_1415 = v_77 | v_1414;
assign v_1420 = v_1416 | v_1419;
assign v_1421 = ~v_1413 | v_1420;
assign v_1422 = v_654 | v_1418;
assign v_1423 = ~v_87 | v_1415;
assign v_1425 = v_1413 | v_1424;
assign v_1429 = v_1427 | v_1428;
assign v_1430 = ~v_1426 | v_1429;
assign v_1431 = v_663 | v_1418;
assign v_1432 = ~v_100 | v_1415;
assign v_1434 = v_1426 | v_1433;
assign v_1438 = v_1436 | v_1437;
assign v_1439 = ~v_1435 | v_1438;
assign v_1440 = v_668 | v_1418;
assign v_1441 = ~v_113 | v_1415;
assign v_1443 = v_1435 | v_1442;
assign v_1448 = v_1445 | v_1447;
assign v_1449 = ~v_1444 | v_1448;
assign v_1450 = v_129 | v_1002;
assign v_1451 = v_126 | ~v_1446;
assign v_1453 = v_1444 | v_1452;
assign v_1458 = v_1455 | v_1457;
assign v_1459 = ~v_1454 | v_1458;
assign v_1460 = v_129 | v_996;
assign v_1461 = v_126 | ~v_1456;
assign v_1463 = v_1454 | v_1462;
assign v_1468 = v_1465 | v_1467;
assign v_1469 = ~v_1464 | v_1468;
assign v_1470 = v_129 | v_1009;
assign v_1471 = v_126 | ~v_1466;
assign v_1473 = v_1464 | v_1472;
assign v_1475 = ~v_67 | v_193;
assign v_1476 = v_77 | v_1475;
assign v_1481 = v_1477 | v_1480;
assign v_1482 = ~v_1474 | v_1481;
assign v_1483 = v_959 | v_1479;
assign v_1484 = ~v_87 | v_1476;
assign v_1486 = v_1474 | v_1485;
assign v_1490 = v_1488 | v_1489;
assign v_1491 = ~v_1487 | v_1490;
assign v_1492 = v_950 | v_1479;
assign v_1493 = ~v_100 | v_1476;
assign v_1495 = v_1487 | v_1494;
assign v_1499 = v_1497 | v_1498;
assign v_1500 = ~v_1496 | v_1499;
assign v_1501 = v_969 | v_1479;
assign v_1502 = ~v_113 | v_1476;
assign v_1504 = v_1496 | v_1503;
assign v_1508 = v_1506 | v_1507;
assign v_1509 = ~v_1505 | v_1508;
assign v_1510 = v_933 | v_1479;
assign v_1511 = v_959 | v_1476;
assign v_1513 = v_1505 | v_1512;
assign v_1517 = v_1515 | v_1516;
assign v_1518 = ~v_1514 | v_1517;
assign v_1519 = v_927 | v_1479;
assign v_1520 = v_950 | v_1476;
assign v_1522 = v_1514 | v_1521;
assign v_1526 = v_1524 | v_1525;
assign v_1527 = ~v_1523 | v_1526;
assign v_1528 = v_940 | v_1479;
assign v_1529 = v_969 | v_1476;
assign v_1531 = v_1523 | v_1530;
assign v_1535 = v_1533 | v_1534;
assign v_1536 = ~v_1532 | v_1535;
assign v_1537 = v_533 | v_539;
assign v_1538 = ~v_87 | v_527;
assign v_1540 = v_1532 | v_1539;
assign v_1544 = v_1542 | v_1543;
assign v_1545 = ~v_1541 | v_1544;
assign v_1546 = v_533 | v_554;
assign v_1547 = ~v_100 | v_527;
assign v_1549 = v_1541 | v_1548;
assign v_1553 = v_1551 | v_1552;
assign v_1554 = ~v_1550 | v_1553;
assign v_1555 = v_533 | v_569;
assign v_1556 = ~v_113 | v_527;
assign v_1558 = v_1550 | v_1557;
assign v_1562 = v_1560 | v_1561;
assign v_1563 = ~v_1559 | v_1562;
assign v_1564 = v_590 | v_596;
assign v_1565 = ~v_87 | v_584;
assign v_1567 = v_1559 | v_1566;
assign v_1571 = v_1569 | v_1570;
assign v_1572 = ~v_1568 | v_1571;
assign v_1573 = v_590 | v_611;
assign v_1574 = ~v_100 | v_584;
assign v_1576 = v_1568 | v_1575;
assign v_1580 = v_1578 | v_1579;
assign v_1581 = ~v_1577 | v_1580;
assign v_1582 = v_590 | v_626;
assign v_1583 = ~v_113 | v_584;
assign v_1585 = v_1577 | v_1584;
assign v_1587 = v_69 | v_72;
assign v_1589 = v_1378 | v_1388;
assign v_1591 = v_1588 | v_1590;
assign v_1592 = ~v_1586 | v_1591;
assign v_1594 = ~v_74 | v_1593;
assign v_1596 = v_1403 | v_1595;
assign v_1598 = v_1586 | v_1597;
assign v_1599 = ~v_61 | ~v_62 | v_388 | v_841;
assign v_1600 = ~v_61 | ~v_297 | v_841;
assign v_1601 = ~v_61 | ~v_373 | v_841;
assign v_1602 = ~v_61 | ~v_388 | v_1237;
assign v_1603 = ~v_61 | v_191 | ~v_388 | v_841 | v_1367;
assign v_1604 = ~v_61 | v_208 | ~v_388 | v_841 | v_1367;
assign v_1605 = ~v_61 | ~v_388 | v_841 | v_1374;
assign v_1606 = ~v_61 | v_841 | ~v_1237 | v_1374;
assign v_1607 = ~v_61 | v_841 | ~v_1237 | v_1387;
assign v_1608 = ~v_61 | v_841 | v_1237 | ~v_1374;
assign v_1609 = ~v_61 | v_841 | ~v_1400;
assign v_1611 = ~v_61 | v_373 | v_1237 | ~v_1387;
assign v_1612 = ~v_61 | v_191 | ~v_373 | ~v_1367;
assign v_1613 = ~v_61 | v_208 | ~v_373 | ~v_1367;
assign v_1614 = ~v_61 | ~v_297 | v_1237;
assign v_1615 = ~v_61 | ~v_297 | ~v_1367;
assign v_1616 = ~v_61 | ~v_297 | ~v_1387;
assign v_1617 = ~v_61 | ~v_1273;
assign v_1618 = ~v_61 | ~v_297 | ~v_1374;
assign v_1619 = ~v_61 | ~v_373 | ~v_1374;
assign v_1620 = ~v_61 | ~v_373 | ~v_1367 | v_1387;
assign v_1621 = ~v_61 | ~v_373 | v_1237 | v_1387;
assign v_1622 = ~v_61 | v_1237 | ~v_1400;
assign v_1623 = ~v_61 | v_373 | v_388 | ~v_1237 | ~v_1367;
assign v_1624 = ~v_61 | ~v_62 | v_1237;
assign v_1625 = ~v_61 | ~v_191 | v_388 | ~v_1367 | ~v_1374;
assign v_1626 = ~v_61 | v_208 | v_388 | ~v_1367 | ~v_1374;
assign v_1627 = ~v_61 | ~v_1260;
assign v_1628 = ~v_61 | ~v_1374 | ~v_1400;
assign v_1629 = ~v_61 | ~v_62 | v_388 | ~v_1374;
assign v_1630 = ~v_61 | v_191 | v_373 | v_388 | ~v_1387;
assign v_1631 = ~v_61 | v_373 | v_388 | ~v_841 | ~v_1387;
assign v_1632 = ~v_61 | v_208 | v_388 | v_841 | ~v_1237;
assign v_1633 = ~v_61 | ~v_388 | ~v_841 | v_1367 | ~v_1374;
assign v_1634 = ~v_61 | ~v_388 | ~v_841 | v_1367 | ~v_1387;
assign v_1635 = ~v_61 | ~v_388 | ~v_1367 | v_1374;
assign v_1636 = ~v_61 | ~v_62 | v_841 | v_1367;
assign v_1637 = ~v_61 | ~v_62 | ~v_373 | ~v_1367;
assign v_1638 = ~v_61 | ~v_1367 | ~v_1400;
assign v_1639 = ~v_61 | ~v_373 | ~v_1237 | v_1367 | ~v_1387;
assign v_1640 = ~v_61 | ~v_62 | ~v_1367 | v_1387;
assign v_1641 = ~v_61 | ~v_388 | ~v_1367 | v_1387;
assign v_1698 = v_5 | v_7 | v_9 | v_11 | v_14;
assign v_1699 = v_16 | v_18 | v_19 | v_21 | v_22;
assign v_1700 = v_24 | v_26 | v_27 | v_28 | v_29;
assign v_1701 = v_30 | v_31 | v_32 | v_34 | v_35;
assign v_1702 = v_36 | v_37 | v_38 | v_39 | v_40;
assign v_1703 = v_41 | v_42 | v_43 | v_45 | v_46;
assign v_1704 = v_47 | v_48 | v_49 | v_50 | v_51;
assign v_1705 = v_52 | v_53 | v_54 | v_55 | v_56;
assign v_1706 = v_57 | v_58 | v_59;
assign v_1707 = v_1698 | v_1699 | v_1700 | v_1701 | v_1702;
assign v_1708 = v_1703 | v_1704 | v_1705 | v_1706;
assign x_1 = v_60 | v_1643;
assign o_1 = x_1;
endmodule
