// skolem function for order file variables
// Generated using findDep.cpp 
module formula (v_10415, v_98, v_721, v_731, v_741, v_751, v_761, v_771, v_793, v_804, v_838, v_850, v_862, v_874, v_886, v_898, v_922, v_940, v_984, v_996, v_1008, v_1020, v_1032, v_1044, v_1072, v_1085, v_1116, v_1128, v_1140, v_1152, v_1164, v_1176, v_1204, v_1221, v_1272, v_1284, v_1296, v_1308, v_1320, v_1332, v_1360, v_1373, v_1404, v_1416, v_1428, v_1440, v_1452, v_1464, v_1492, v_1511, v_1556, v_1568, v_1580, v_1592, v_1604, v_1616, v_1644, v_1657, v_1688, v_1700, v_1712, v_1724, v_1736, v_1748, v_1776, v_1793, v_1852, v_1864, v_1876, v_1888, v_1900, v_1912, v_1940, v_1953, v_1984, v_1996, v_2008, v_2020, v_2032, v_2044, v_2072, v_2090, v_2134, v_2146, v_2158, v_2170, v_2182, v_2194, v_2222, v_2235, v_2266, v_2278, v_2290, v_2302, v_2314, v_2326, v_2354, v_2371, v_2422, v_2434, v_2446, v_2458, v_2470, v_2482, v_2510, v_2523, v_2554, v_2566, v_2578, v_2590, v_2602, v_2614, v_2642, v_2662, v_2708, v_2720, v_2732, v_2744, v_2756, v_2768, v_2796, v_2809, v_2840, v_2852, v_2864, v_2876, v_2888, v_2900, v_2928, v_2945, v_3012, v_3024, v_3036, v_3048, v_3060, v_3072, v_3100, v_3113, v_3144, v_3156, v_3168, v_3180, v_3192, v_3204, v_3232, v_3250, v_3294, v_3306, v_3318, v_3330, v_3342, v_3354, v_3382, v_3395, v_3426, v_3438, v_3450, v_3462, v_3474, v_3486, v_3514, v_3531, v_3582, v_3594, v_3606, v_3618, v_3630, v_3642, v_3670, v_3683, v_3714, v_3726, v_3738, v_3750, v_3762, v_3774, v_3802, v_3821, v_3866, v_3878, v_3890, v_3902, v_3914, v_3926, v_3954, v_3967, v_3998, v_4010, v_4022, v_4034, v_4046, v_4058, v_4086, v_4103, v_4162, v_4174, v_4186, v_4198, v_4210, v_4222, v_4250, v_4263, v_4294, v_4306, v_4318, v_4330, v_4342, v_4354, v_4382, v_4400, v_4444, v_4456, v_4468, v_4480, v_4492, v_4504, v_4532, v_4545, v_4576, v_4588, v_4600, v_4612, v_4624, v_4636, v_4664, v_4681, v_4732, v_4744, v_4756, v_4768, v_4780, v_4792, v_4820, v_4833, v_4864, v_4876, v_4888, v_4900, v_4912, v_4924, v_4952, v_4973, v_5020, v_5032, v_5044, v_5056, v_5068, v_5080, v_5108, v_5121, v_5152, v_5164, v_5176, v_5188, v_5200, v_5212, v_5240, v_5257, v_5332, v_5344, v_5356, v_5368, v_5380, v_5392, v_5420, v_5433, v_5464, v_5476, v_5488, v_5500, v_5512, v_5524, v_5552, v_5570, v_5614, v_5626, v_5638, v_5650, v_5662, v_5674, v_5702, v_5715, v_5746, v_5758, v_5770, v_5782, v_5794, v_5806, v_5834, v_5851, v_5902, v_5914, v_5926, v_5938, v_5950, v_5962, v_5990, v_6003, v_6034, v_6046, v_6058, v_6070, v_6082, v_6094, v_6122, v_6141, v_6186, v_6198, v_6210, v_6222, v_6234, v_6246, v_6274, v_6287, v_6318, v_6330, v_6342, v_6354, v_6366, v_6378, v_6406, v_6423, v_6482, v_6494, v_6506, v_6518, v_6530, v_6542, v_6570, v_6583, v_6614, v_6626, v_6638, v_6650, v_6662, v_6674, v_6702, v_6720, v_6764, v_6776, v_6788, v_6800, v_6812, v_6824, v_6852, v_6865, v_6896, v_6908, v_6920, v_6932, v_6944, v_6956, v_6984, v_7001, v_7052, v_7064, v_7076, v_7088, v_7100, v_7112, v_7140, v_7153, v_7184, v_7196, v_7208, v_7220, v_7232, v_7244, v_7272, v_7292, v_7338, v_7350, v_7362, v_7374, v_7386, v_7398, v_7426, v_7439, v_7470, v_7482, v_7494, v_7506, v_7518, v_7530, v_7558, v_7575, v_7642, v_7654, v_7666, v_7678, v_7690, v_7702, v_7730, v_7743, v_7774, v_7786, v_7798, v_7810, v_7822, v_7834, v_7862, v_7880, v_7924, v_7936, v_7948, v_7960, v_7972, v_7984, v_8012, v_8025, v_8056, v_8068, v_8080, v_8092, v_8104, v_8116, v_8144, v_8161, v_8212, v_8224, v_8236, v_8248, v_8260, v_8272, v_8300, v_8313, v_8344, v_8356, v_8368, v_8380, v_8392, v_8404, v_8432, v_8451, v_8496, v_8508, v_8520, v_8532, v_8544, v_8556, v_8584, v_8597, v_8628, v_8640, v_8652, v_8664, v_8676, v_8688, v_8716, v_8733, v_8792, v_8804, v_8816, v_8828, v_8840, v_8852, v_8880, v_8893, v_8924, v_8936, v_8948, v_8960, v_8972, v_8984, v_9012, v_9030, v_9074, v_9086, v_9098, v_9110, v_9122, v_9134, v_9162, v_9175, v_9206, v_9218, v_9230, v_9242, v_9254, v_9266, v_9294, v_9311, v_9362, v_9374, v_9386, v_9398, v_9410, v_9422, v_9450, v_9463, v_9494, v_9506, v_9518, v_9530, v_9542, v_9554, v_9582, v_9604, v_9652, v_9664, v_9676, v_9688, v_9700, v_9712, v_9740, v_9753, v_9784, v_9796, v_9808, v_9820, v_9832, v_9844, v_9872, v_9, v_14, v_19, v_24, v_29, v_87, v_89, v_91, v_47, v_45, v_43, v_8, v_13, v_18, v_23, v_28, v_10414, v_10421, v_10427, v_10433, v_10439, v_10445, v_10451, v_4, v_10462, v_3, v_1, v_563, v_361, v_96, v_807, v_9903, v_9884, v_10200, v_10196, v_7, v_720, v_730, v_740, v_750, v_760, v_770, v_792, v_802, v_837, v_849, v_861, v_873, v_885, v_897, v_921, v_933, v_983, v_995, v_1007, v_1019, v_1031, v_1043, v_1071, v_1083, v_1115, v_1127, v_1139, v_1151, v_1163, v_1175, v_1203, v_1215, v_1271, v_1283, v_1295, v_1307, v_1319, v_1331, v_1359, v_1371, v_1403, v_1415, v_1427, v_1439, v_1451, v_1463, v_1491, v_1503, v_1555, v_1567, v_1579, v_1591, v_1603, v_1615, v_1643, v_1655, v_1687, v_1699, v_1711, v_1723, v_1735, v_1747, v_1775, v_1787, v_1851, v_1863, v_1875, v_1887, v_1899, v_1911, v_1939, v_1951, v_1983, v_1995, v_2007, v_2019, v_2031, v_2043, v_2071, v_2083, v_2133, v_2145, v_2157, v_2169, v_2181, v_2193, v_2221, v_2233, v_2265, v_2277, v_2289, v_2301, v_2313, v_2325, v_2353, v_2365, v_2421, v_2433, v_2445, v_2457, v_2469, v_2481, v_2509, v_2521, v_2553, v_2565, v_2577, v_2589, v_2601, v_2613, v_2641, v_2653, v_2707, v_2719, v_2731, v_2743, v_2755, v_2767, v_2795, v_2807, v_2839, v_2851, v_2863, v_2875, v_2887, v_2899, v_2927, v_2939, v_3011, v_3023, v_3035, v_3047, v_3059, v_3071, v_3099, v_3111, v_3143, v_3155, v_3167, v_3179, v_3191, v_3203, v_3231, v_3243, v_3293, v_3305, v_3317, v_3329, v_3341, v_3353, v_3381, v_3393, v_3425, v_3437, v_3449, v_3461, v_3473, v_3485, v_3513, v_3525, v_3581, v_3593, v_3605, v_3617, v_3629, v_3641, v_3669, v_3681, v_3713, v_3725, v_3737, v_3749, v_3761, v_3773, v_3801, v_3813, v_3865, v_3877, v_3889, v_3901, v_3913, v_3925, v_3953, v_3965, v_3997, v_4009, v_4021, v_4033, v_4045, v_4057, v_4085, v_4097, v_4161, v_4173, v_4185, v_4197, v_4209, v_4221, v_4249, v_4261, v_4293, v_4305, v_4317, v_4329, v_4341, v_4353, v_4381, v_4393, v_4443, v_4455, v_4467, v_4479, v_4491, v_4503, v_4531, v_4543, v_4575, v_4587, v_4599, v_4611, v_4623, v_4635, v_4663, v_4675, v_4731, v_4743, v_4755, v_4767, v_4779, v_4791, v_4819, v_4831, v_4863, v_4875, v_4887, v_4899, v_4911, v_4923, v_4951, v_4963, v_5019, v_5031, v_5043, v_5055, v_5067, v_5079, v_5107, v_5119, v_5151, v_5163, v_5175, v_5187, v_5199, v_5211, v_5239, v_5251, v_5331, v_5343, v_5355, v_5367, v_5379, v_5391, v_5419, v_5431, v_5463, v_5475, v_5487, v_5499, v_5511, v_5523, v_5551, v_5563, v_5613, v_5625, v_5637, v_5649, v_5661, v_5673, v_5701, v_5713, v_5745, v_5757, v_5769, v_5781, v_5793, v_5805, v_5833, v_5845, v_5901, v_5913, v_5925, v_5937, v_5949, v_5961, v_5989, v_6001, v_6033, v_6045, v_6057, v_6069, v_6081, v_6093, v_6121, v_6133, v_6185, v_6197, v_6209, v_6221, v_6233, v_6245, v_6273, v_6285, v_6317, v_6329, v_6341, v_6353, v_6365, v_6377, v_6405, v_6417, v_6481, v_6493, v_6505, v_6517, v_6529, v_6541, v_6569, v_6581, v_6613, v_6625, v_6637, v_6649, v_6661, v_6673, v_6701, v_6713, v_6763, v_6775, v_6787, v_6799, v_6811, v_6823, v_6851, v_6863, v_6895, v_6907, v_6919, v_6931, v_6943, v_6955, v_6983, v_6995, v_7051, v_7063, v_7075, v_7087, v_7099, v_7111, v_7139, v_7151, v_7183, v_7195, v_7207, v_7219, v_7231, v_7243, v_7271, v_7283, v_7337, v_7349, v_7361, v_7373, v_7385, v_7397, v_7425, v_7437, v_7469, v_7481, v_7493, v_7505, v_7517, v_7529, v_7557, v_7569, v_7641, v_7653, v_7665, v_7677, v_7689, v_7701, v_7729, v_7741, v_7773, v_7785, v_7797, v_7809, v_7821, v_7833, v_7861, v_7873, v_7923, v_7935, v_7947, v_7959, v_7971, v_7983, v_8011, v_8023, v_8055, v_8067, v_8079, v_8091, v_8103, v_8115, v_8143, v_8155, v_8211, v_8223, v_8235, v_8247, v_8259, v_8271, v_8299, v_8311, v_8343, v_8355, v_8367, v_8379, v_8391, v_8403, v_8431, v_8443, v_8495, v_8507, v_8519, v_8531, v_8543, v_8555, v_8583, v_8595, v_8627, v_8639, v_8651, v_8663, v_8675, v_8687, v_8715, v_8727, v_8791, v_8803, v_8815, v_8827, v_8839, v_8851, v_8879, v_8891, v_8923, v_8935, v_8947, v_8959, v_8971, v_8983, v_9011, v_9023, v_9073, v_9085, v_9097, v_9109, v_9121, v_9133, v_9161, v_9173, v_9205, v_9217, v_9229, v_9241, v_9253, v_9265, v_9293, v_9305, v_9361, v_9373, v_9385, v_9397, v_9409, v_9421, v_9449, v_9461, v_9493, v_9505, v_9517, v_9529, v_9541, v_9553, v_9581, v_9593, v_9651, v_9663, v_9675, v_9687, v_9699, v_9711, v_9739, v_9751, v_9783, v_9795, v_9807, v_9819, v_9831, v_9843, v_9871, v_9883, v_9948, v_9985, v_10022, v_10059, v_10096, v_10133, v_10168, v_10195, v_10224, v_10251, v_10278, v_10305, v_10332, v_10359, v_10386, v_10413, v_10420, v_10426, v_10432, v_10438, v_10444, v_10450, v_10456, v_10461, v_10465, v_34852, o_1);
input v_10415;
input v_98;
input v_721;
input v_731;
input v_741;
input v_751;
input v_761;
input v_771;
input v_793;
input v_804;
input v_838;
input v_850;
input v_862;
input v_874;
input v_886;
input v_898;
input v_922;
input v_940;
input v_984;
input v_996;
input v_1008;
input v_1020;
input v_1032;
input v_1044;
input v_1072;
input v_1085;
input v_1116;
input v_1128;
input v_1140;
input v_1152;
input v_1164;
input v_1176;
input v_1204;
input v_1221;
input v_1272;
input v_1284;
input v_1296;
input v_1308;
input v_1320;
input v_1332;
input v_1360;
input v_1373;
input v_1404;
input v_1416;
input v_1428;
input v_1440;
input v_1452;
input v_1464;
input v_1492;
input v_1511;
input v_1556;
input v_1568;
input v_1580;
input v_1592;
input v_1604;
input v_1616;
input v_1644;
input v_1657;
input v_1688;
input v_1700;
input v_1712;
input v_1724;
input v_1736;
input v_1748;
input v_1776;
input v_1793;
input v_1852;
input v_1864;
input v_1876;
input v_1888;
input v_1900;
input v_1912;
input v_1940;
input v_1953;
input v_1984;
input v_1996;
input v_2008;
input v_2020;
input v_2032;
input v_2044;
input v_2072;
input v_2090;
input v_2134;
input v_2146;
input v_2158;
input v_2170;
input v_2182;
input v_2194;
input v_2222;
input v_2235;
input v_2266;
input v_2278;
input v_2290;
input v_2302;
input v_2314;
input v_2326;
input v_2354;
input v_2371;
input v_2422;
input v_2434;
input v_2446;
input v_2458;
input v_2470;
input v_2482;
input v_2510;
input v_2523;
input v_2554;
input v_2566;
input v_2578;
input v_2590;
input v_2602;
input v_2614;
input v_2642;
input v_2662;
input v_2708;
input v_2720;
input v_2732;
input v_2744;
input v_2756;
input v_2768;
input v_2796;
input v_2809;
input v_2840;
input v_2852;
input v_2864;
input v_2876;
input v_2888;
input v_2900;
input v_2928;
input v_2945;
input v_3012;
input v_3024;
input v_3036;
input v_3048;
input v_3060;
input v_3072;
input v_3100;
input v_3113;
input v_3144;
input v_3156;
input v_3168;
input v_3180;
input v_3192;
input v_3204;
input v_3232;
input v_3250;
input v_3294;
input v_3306;
input v_3318;
input v_3330;
input v_3342;
input v_3354;
input v_3382;
input v_3395;
input v_3426;
input v_3438;
input v_3450;
input v_3462;
input v_3474;
input v_3486;
input v_3514;
input v_3531;
input v_3582;
input v_3594;
input v_3606;
input v_3618;
input v_3630;
input v_3642;
input v_3670;
input v_3683;
input v_3714;
input v_3726;
input v_3738;
input v_3750;
input v_3762;
input v_3774;
input v_3802;
input v_3821;
input v_3866;
input v_3878;
input v_3890;
input v_3902;
input v_3914;
input v_3926;
input v_3954;
input v_3967;
input v_3998;
input v_4010;
input v_4022;
input v_4034;
input v_4046;
input v_4058;
input v_4086;
input v_4103;
input v_4162;
input v_4174;
input v_4186;
input v_4198;
input v_4210;
input v_4222;
input v_4250;
input v_4263;
input v_4294;
input v_4306;
input v_4318;
input v_4330;
input v_4342;
input v_4354;
input v_4382;
input v_4400;
input v_4444;
input v_4456;
input v_4468;
input v_4480;
input v_4492;
input v_4504;
input v_4532;
input v_4545;
input v_4576;
input v_4588;
input v_4600;
input v_4612;
input v_4624;
input v_4636;
input v_4664;
input v_4681;
input v_4732;
input v_4744;
input v_4756;
input v_4768;
input v_4780;
input v_4792;
input v_4820;
input v_4833;
input v_4864;
input v_4876;
input v_4888;
input v_4900;
input v_4912;
input v_4924;
input v_4952;
input v_4973;
input v_5020;
input v_5032;
input v_5044;
input v_5056;
input v_5068;
input v_5080;
input v_5108;
input v_5121;
input v_5152;
input v_5164;
input v_5176;
input v_5188;
input v_5200;
input v_5212;
input v_5240;
input v_5257;
input v_5332;
input v_5344;
input v_5356;
input v_5368;
input v_5380;
input v_5392;
input v_5420;
input v_5433;
input v_5464;
input v_5476;
input v_5488;
input v_5500;
input v_5512;
input v_5524;
input v_5552;
input v_5570;
input v_5614;
input v_5626;
input v_5638;
input v_5650;
input v_5662;
input v_5674;
input v_5702;
input v_5715;
input v_5746;
input v_5758;
input v_5770;
input v_5782;
input v_5794;
input v_5806;
input v_5834;
input v_5851;
input v_5902;
input v_5914;
input v_5926;
input v_5938;
input v_5950;
input v_5962;
input v_5990;
input v_6003;
input v_6034;
input v_6046;
input v_6058;
input v_6070;
input v_6082;
input v_6094;
input v_6122;
input v_6141;
input v_6186;
input v_6198;
input v_6210;
input v_6222;
input v_6234;
input v_6246;
input v_6274;
input v_6287;
input v_6318;
input v_6330;
input v_6342;
input v_6354;
input v_6366;
input v_6378;
input v_6406;
input v_6423;
input v_6482;
input v_6494;
input v_6506;
input v_6518;
input v_6530;
input v_6542;
input v_6570;
input v_6583;
input v_6614;
input v_6626;
input v_6638;
input v_6650;
input v_6662;
input v_6674;
input v_6702;
input v_6720;
input v_6764;
input v_6776;
input v_6788;
input v_6800;
input v_6812;
input v_6824;
input v_6852;
input v_6865;
input v_6896;
input v_6908;
input v_6920;
input v_6932;
input v_6944;
input v_6956;
input v_6984;
input v_7001;
input v_7052;
input v_7064;
input v_7076;
input v_7088;
input v_7100;
input v_7112;
input v_7140;
input v_7153;
input v_7184;
input v_7196;
input v_7208;
input v_7220;
input v_7232;
input v_7244;
input v_7272;
input v_7292;
input v_7338;
input v_7350;
input v_7362;
input v_7374;
input v_7386;
input v_7398;
input v_7426;
input v_7439;
input v_7470;
input v_7482;
input v_7494;
input v_7506;
input v_7518;
input v_7530;
input v_7558;
input v_7575;
input v_7642;
input v_7654;
input v_7666;
input v_7678;
input v_7690;
input v_7702;
input v_7730;
input v_7743;
input v_7774;
input v_7786;
input v_7798;
input v_7810;
input v_7822;
input v_7834;
input v_7862;
input v_7880;
input v_7924;
input v_7936;
input v_7948;
input v_7960;
input v_7972;
input v_7984;
input v_8012;
input v_8025;
input v_8056;
input v_8068;
input v_8080;
input v_8092;
input v_8104;
input v_8116;
input v_8144;
input v_8161;
input v_8212;
input v_8224;
input v_8236;
input v_8248;
input v_8260;
input v_8272;
input v_8300;
input v_8313;
input v_8344;
input v_8356;
input v_8368;
input v_8380;
input v_8392;
input v_8404;
input v_8432;
input v_8451;
input v_8496;
input v_8508;
input v_8520;
input v_8532;
input v_8544;
input v_8556;
input v_8584;
input v_8597;
input v_8628;
input v_8640;
input v_8652;
input v_8664;
input v_8676;
input v_8688;
input v_8716;
input v_8733;
input v_8792;
input v_8804;
input v_8816;
input v_8828;
input v_8840;
input v_8852;
input v_8880;
input v_8893;
input v_8924;
input v_8936;
input v_8948;
input v_8960;
input v_8972;
input v_8984;
input v_9012;
input v_9030;
input v_9074;
input v_9086;
input v_9098;
input v_9110;
input v_9122;
input v_9134;
input v_9162;
input v_9175;
input v_9206;
input v_9218;
input v_9230;
input v_9242;
input v_9254;
input v_9266;
input v_9294;
input v_9311;
input v_9362;
input v_9374;
input v_9386;
input v_9398;
input v_9410;
input v_9422;
input v_9450;
input v_9463;
input v_9494;
input v_9506;
input v_9518;
input v_9530;
input v_9542;
input v_9554;
input v_9582;
input v_9604;
input v_9652;
input v_9664;
input v_9676;
input v_9688;
input v_9700;
input v_9712;
input v_9740;
input v_9753;
input v_9784;
input v_9796;
input v_9808;
input v_9820;
input v_9832;
input v_9844;
input v_9872;
input v_9;
input v_14;
input v_19;
input v_24;
input v_29;
input v_87;
input v_89;
input v_91;
input v_47;
input v_45;
input v_43;
input v_8;
input v_13;
input v_18;
input v_23;
input v_28;
input v_10414;
input v_10421;
input v_10427;
input v_10433;
input v_10439;
input v_10445;
input v_10451;
input v_4;
input v_10462;
input v_3;
input v_1;
input v_563;
input v_361;
input v_96;
input v_807;
input v_9903;
input v_9884;
input v_10200;
input v_10196;
input v_7;
input v_720;
input v_730;
input v_740;
input v_750;
input v_760;
input v_770;
input v_792;
input v_802;
input v_837;
input v_849;
input v_861;
input v_873;
input v_885;
input v_897;
input v_921;
input v_933;
input v_983;
input v_995;
input v_1007;
input v_1019;
input v_1031;
input v_1043;
input v_1071;
input v_1083;
input v_1115;
input v_1127;
input v_1139;
input v_1151;
input v_1163;
input v_1175;
input v_1203;
input v_1215;
input v_1271;
input v_1283;
input v_1295;
input v_1307;
input v_1319;
input v_1331;
input v_1359;
input v_1371;
input v_1403;
input v_1415;
input v_1427;
input v_1439;
input v_1451;
input v_1463;
input v_1491;
input v_1503;
input v_1555;
input v_1567;
input v_1579;
input v_1591;
input v_1603;
input v_1615;
input v_1643;
input v_1655;
input v_1687;
input v_1699;
input v_1711;
input v_1723;
input v_1735;
input v_1747;
input v_1775;
input v_1787;
input v_1851;
input v_1863;
input v_1875;
input v_1887;
input v_1899;
input v_1911;
input v_1939;
input v_1951;
input v_1983;
input v_1995;
input v_2007;
input v_2019;
input v_2031;
input v_2043;
input v_2071;
input v_2083;
input v_2133;
input v_2145;
input v_2157;
input v_2169;
input v_2181;
input v_2193;
input v_2221;
input v_2233;
input v_2265;
input v_2277;
input v_2289;
input v_2301;
input v_2313;
input v_2325;
input v_2353;
input v_2365;
input v_2421;
input v_2433;
input v_2445;
input v_2457;
input v_2469;
input v_2481;
input v_2509;
input v_2521;
input v_2553;
input v_2565;
input v_2577;
input v_2589;
input v_2601;
input v_2613;
input v_2641;
input v_2653;
input v_2707;
input v_2719;
input v_2731;
input v_2743;
input v_2755;
input v_2767;
input v_2795;
input v_2807;
input v_2839;
input v_2851;
input v_2863;
input v_2875;
input v_2887;
input v_2899;
input v_2927;
input v_2939;
input v_3011;
input v_3023;
input v_3035;
input v_3047;
input v_3059;
input v_3071;
input v_3099;
input v_3111;
input v_3143;
input v_3155;
input v_3167;
input v_3179;
input v_3191;
input v_3203;
input v_3231;
input v_3243;
input v_3293;
input v_3305;
input v_3317;
input v_3329;
input v_3341;
input v_3353;
input v_3381;
input v_3393;
input v_3425;
input v_3437;
input v_3449;
input v_3461;
input v_3473;
input v_3485;
input v_3513;
input v_3525;
input v_3581;
input v_3593;
input v_3605;
input v_3617;
input v_3629;
input v_3641;
input v_3669;
input v_3681;
input v_3713;
input v_3725;
input v_3737;
input v_3749;
input v_3761;
input v_3773;
input v_3801;
input v_3813;
input v_3865;
input v_3877;
input v_3889;
input v_3901;
input v_3913;
input v_3925;
input v_3953;
input v_3965;
input v_3997;
input v_4009;
input v_4021;
input v_4033;
input v_4045;
input v_4057;
input v_4085;
input v_4097;
input v_4161;
input v_4173;
input v_4185;
input v_4197;
input v_4209;
input v_4221;
input v_4249;
input v_4261;
input v_4293;
input v_4305;
input v_4317;
input v_4329;
input v_4341;
input v_4353;
input v_4381;
input v_4393;
input v_4443;
input v_4455;
input v_4467;
input v_4479;
input v_4491;
input v_4503;
input v_4531;
input v_4543;
input v_4575;
input v_4587;
input v_4599;
input v_4611;
input v_4623;
input v_4635;
input v_4663;
input v_4675;
input v_4731;
input v_4743;
input v_4755;
input v_4767;
input v_4779;
input v_4791;
input v_4819;
input v_4831;
input v_4863;
input v_4875;
input v_4887;
input v_4899;
input v_4911;
input v_4923;
input v_4951;
input v_4963;
input v_5019;
input v_5031;
input v_5043;
input v_5055;
input v_5067;
input v_5079;
input v_5107;
input v_5119;
input v_5151;
input v_5163;
input v_5175;
input v_5187;
input v_5199;
input v_5211;
input v_5239;
input v_5251;
input v_5331;
input v_5343;
input v_5355;
input v_5367;
input v_5379;
input v_5391;
input v_5419;
input v_5431;
input v_5463;
input v_5475;
input v_5487;
input v_5499;
input v_5511;
input v_5523;
input v_5551;
input v_5563;
input v_5613;
input v_5625;
input v_5637;
input v_5649;
input v_5661;
input v_5673;
input v_5701;
input v_5713;
input v_5745;
input v_5757;
input v_5769;
input v_5781;
input v_5793;
input v_5805;
input v_5833;
input v_5845;
input v_5901;
input v_5913;
input v_5925;
input v_5937;
input v_5949;
input v_5961;
input v_5989;
input v_6001;
input v_6033;
input v_6045;
input v_6057;
input v_6069;
input v_6081;
input v_6093;
input v_6121;
input v_6133;
input v_6185;
input v_6197;
input v_6209;
input v_6221;
input v_6233;
input v_6245;
input v_6273;
input v_6285;
input v_6317;
input v_6329;
input v_6341;
input v_6353;
input v_6365;
input v_6377;
input v_6405;
input v_6417;
input v_6481;
input v_6493;
input v_6505;
input v_6517;
input v_6529;
input v_6541;
input v_6569;
input v_6581;
input v_6613;
input v_6625;
input v_6637;
input v_6649;
input v_6661;
input v_6673;
input v_6701;
input v_6713;
input v_6763;
input v_6775;
input v_6787;
input v_6799;
input v_6811;
input v_6823;
input v_6851;
input v_6863;
input v_6895;
input v_6907;
input v_6919;
input v_6931;
input v_6943;
input v_6955;
input v_6983;
input v_6995;
input v_7051;
input v_7063;
input v_7075;
input v_7087;
input v_7099;
input v_7111;
input v_7139;
input v_7151;
input v_7183;
input v_7195;
input v_7207;
input v_7219;
input v_7231;
input v_7243;
input v_7271;
input v_7283;
input v_7337;
input v_7349;
input v_7361;
input v_7373;
input v_7385;
input v_7397;
input v_7425;
input v_7437;
input v_7469;
input v_7481;
input v_7493;
input v_7505;
input v_7517;
input v_7529;
input v_7557;
input v_7569;
input v_7641;
input v_7653;
input v_7665;
input v_7677;
input v_7689;
input v_7701;
input v_7729;
input v_7741;
input v_7773;
input v_7785;
input v_7797;
input v_7809;
input v_7821;
input v_7833;
input v_7861;
input v_7873;
input v_7923;
input v_7935;
input v_7947;
input v_7959;
input v_7971;
input v_7983;
input v_8011;
input v_8023;
input v_8055;
input v_8067;
input v_8079;
input v_8091;
input v_8103;
input v_8115;
input v_8143;
input v_8155;
input v_8211;
input v_8223;
input v_8235;
input v_8247;
input v_8259;
input v_8271;
input v_8299;
input v_8311;
input v_8343;
input v_8355;
input v_8367;
input v_8379;
input v_8391;
input v_8403;
input v_8431;
input v_8443;
input v_8495;
input v_8507;
input v_8519;
input v_8531;
input v_8543;
input v_8555;
input v_8583;
input v_8595;
input v_8627;
input v_8639;
input v_8651;
input v_8663;
input v_8675;
input v_8687;
input v_8715;
input v_8727;
input v_8791;
input v_8803;
input v_8815;
input v_8827;
input v_8839;
input v_8851;
input v_8879;
input v_8891;
input v_8923;
input v_8935;
input v_8947;
input v_8959;
input v_8971;
input v_8983;
input v_9011;
input v_9023;
input v_9073;
input v_9085;
input v_9097;
input v_9109;
input v_9121;
input v_9133;
input v_9161;
input v_9173;
input v_9205;
input v_9217;
input v_9229;
input v_9241;
input v_9253;
input v_9265;
input v_9293;
input v_9305;
input v_9361;
input v_9373;
input v_9385;
input v_9397;
input v_9409;
input v_9421;
input v_9449;
input v_9461;
input v_9493;
input v_9505;
input v_9517;
input v_9529;
input v_9541;
input v_9553;
input v_9581;
input v_9593;
input v_9651;
input v_9663;
input v_9675;
input v_9687;
input v_9699;
input v_9711;
input v_9739;
input v_9751;
input v_9783;
input v_9795;
input v_9807;
input v_9819;
input v_9831;
input v_9843;
input v_9871;
input v_9883;
input v_9948;
input v_9985;
input v_10022;
input v_10059;
input v_10096;
input v_10133;
input v_10168;
input v_10195;
input v_10224;
input v_10251;
input v_10278;
input v_10305;
input v_10332;
input v_10359;
input v_10386;
input v_10413;
input v_10420;
input v_10426;
input v_10432;
input v_10438;
input v_10444;
input v_10450;
input v_10456;
input v_10461;
input v_10465;
input v_34852;
output o_1;
wire v_2;
wire v_5;
wire v_6;
wire v_10;
wire v_11;
wire v_12;
wire v_15;
wire v_16;
wire v_17;
wire v_20;
wire v_21;
wire v_22;
wire v_25;
wire v_26;
wire v_27;
wire v_30;
wire v_31;
wire v_32;
wire v_33;
wire v_34;
wire v_35;
wire v_36;
wire v_37;
wire v_38;
wire v_39;
wire v_40;
wire v_41;
wire v_42;
wire v_44;
wire v_46;
wire v_48;
wire v_49;
wire v_50;
wire v_51;
wire v_52;
wire v_53;
wire v_54;
wire v_55;
wire v_56;
wire v_57;
wire v_58;
wire v_59;
wire v_60;
wire v_61;
wire v_62;
wire v_63;
wire v_64;
wire v_65;
wire v_66;
wire v_67;
wire v_68;
wire v_69;
wire v_70;
wire v_71;
wire v_72;
wire v_73;
wire v_74;
wire v_75;
wire v_76;
wire v_77;
wire v_78;
wire v_79;
wire v_80;
wire v_81;
wire v_82;
wire v_83;
wire v_84;
wire v_85;
wire v_86;
wire v_88;
wire v_90;
wire v_92;
wire v_93;
wire v_94;
wire v_95;
wire v_97;
wire v_99;
wire v_100;
wire v_101;
wire v_102;
wire v_103;
wire v_104;
wire v_105;
wire v_106;
wire v_107;
wire v_108;
wire v_109;
wire v_110;
wire v_111;
wire v_112;
wire v_113;
wire v_114;
wire v_115;
wire v_116;
wire v_117;
wire v_118;
wire v_119;
wire v_120;
wire v_121;
wire v_122;
wire v_123;
wire v_124;
wire v_125;
wire v_126;
wire v_127;
wire v_128;
wire v_129;
wire v_130;
wire v_131;
wire v_132;
wire v_133;
wire v_134;
wire v_135;
wire v_136;
wire v_137;
wire v_138;
wire v_139;
wire v_140;
wire v_141;
wire v_142;
wire v_143;
wire v_144;
wire v_145;
wire v_146;
wire v_147;
wire v_148;
wire v_149;
wire v_150;
wire v_151;
wire v_152;
wire v_153;
wire v_154;
wire v_155;
wire v_156;
wire v_157;
wire v_158;
wire v_159;
wire v_160;
wire v_161;
wire v_162;
wire v_163;
wire v_164;
wire v_165;
wire v_166;
wire v_167;
wire v_168;
wire v_169;
wire v_170;
wire v_171;
wire v_172;
wire v_173;
wire v_174;
wire v_175;
wire v_176;
wire v_177;
wire v_178;
wire v_179;
wire v_180;
wire v_181;
wire v_182;
wire v_183;
wire v_184;
wire v_185;
wire v_186;
wire v_187;
wire v_188;
wire v_189;
wire v_190;
wire v_191;
wire v_192;
wire v_193;
wire v_194;
wire v_195;
wire v_196;
wire v_197;
wire v_198;
wire v_199;
wire v_200;
wire v_201;
wire v_202;
wire v_203;
wire v_204;
wire v_205;
wire v_206;
wire v_207;
wire v_208;
wire v_209;
wire v_210;
wire v_211;
wire v_212;
wire v_213;
wire v_214;
wire v_215;
wire v_216;
wire v_217;
wire v_218;
wire v_219;
wire v_220;
wire v_221;
wire v_222;
wire v_223;
wire v_224;
wire v_225;
wire v_226;
wire v_227;
wire v_228;
wire v_229;
wire v_230;
wire v_231;
wire v_232;
wire v_233;
wire v_234;
wire v_235;
wire v_236;
wire v_237;
wire v_238;
wire v_239;
wire v_240;
wire v_241;
wire v_242;
wire v_243;
wire v_244;
wire v_245;
wire v_246;
wire v_247;
wire v_248;
wire v_249;
wire v_250;
wire v_251;
wire v_252;
wire v_253;
wire v_254;
wire v_255;
wire v_256;
wire v_257;
wire v_258;
wire v_259;
wire v_260;
wire v_261;
wire v_262;
wire v_263;
wire v_264;
wire v_265;
wire v_266;
wire v_267;
wire v_268;
wire v_269;
wire v_270;
wire v_271;
wire v_272;
wire v_273;
wire v_274;
wire v_275;
wire v_276;
wire v_277;
wire v_278;
wire v_279;
wire v_280;
wire v_281;
wire v_282;
wire v_283;
wire v_284;
wire v_285;
wire v_286;
wire v_287;
wire v_288;
wire v_289;
wire v_290;
wire v_291;
wire v_292;
wire v_293;
wire v_294;
wire v_295;
wire v_296;
wire v_297;
wire v_298;
wire v_299;
wire v_300;
wire v_301;
wire v_302;
wire v_303;
wire v_304;
wire v_305;
wire v_306;
wire v_307;
wire v_308;
wire v_309;
wire v_310;
wire v_311;
wire v_312;
wire v_313;
wire v_314;
wire v_315;
wire v_316;
wire v_317;
wire v_318;
wire v_319;
wire v_320;
wire v_321;
wire v_322;
wire v_323;
wire v_324;
wire v_325;
wire v_326;
wire v_327;
wire v_328;
wire v_329;
wire v_330;
wire v_331;
wire v_332;
wire v_333;
wire v_334;
wire v_335;
wire v_336;
wire v_337;
wire v_338;
wire v_339;
wire v_340;
wire v_341;
wire v_342;
wire v_343;
wire v_344;
wire v_345;
wire v_346;
wire v_347;
wire v_348;
wire v_349;
wire v_350;
wire v_351;
wire v_352;
wire v_353;
wire v_354;
wire v_355;
wire v_356;
wire v_357;
wire v_358;
wire v_359;
wire v_360;
wire v_362;
wire v_363;
wire v_364;
wire v_365;
wire v_366;
wire v_367;
wire v_368;
wire v_369;
wire v_370;
wire v_371;
wire v_372;
wire v_373;
wire v_374;
wire v_375;
wire v_376;
wire v_377;
wire v_378;
wire v_379;
wire v_380;
wire v_381;
wire v_382;
wire v_383;
wire v_384;
wire v_385;
wire v_386;
wire v_387;
wire v_388;
wire v_389;
wire v_390;
wire v_391;
wire v_392;
wire v_393;
wire v_394;
wire v_395;
wire v_396;
wire v_397;
wire v_398;
wire v_399;
wire v_400;
wire v_401;
wire v_402;
wire v_403;
wire v_404;
wire v_405;
wire v_406;
wire v_407;
wire v_408;
wire v_409;
wire v_410;
wire v_411;
wire v_412;
wire v_413;
wire v_414;
wire v_415;
wire v_416;
wire v_417;
wire v_418;
wire v_419;
wire v_420;
wire v_421;
wire v_422;
wire v_423;
wire v_424;
wire v_425;
wire v_426;
wire v_427;
wire v_428;
wire v_429;
wire v_430;
wire v_431;
wire v_432;
wire v_433;
wire v_434;
wire v_435;
wire v_436;
wire v_437;
wire v_438;
wire v_439;
wire v_440;
wire v_441;
wire v_442;
wire v_443;
wire v_444;
wire v_445;
wire v_446;
wire v_447;
wire v_448;
wire v_449;
wire v_450;
wire v_451;
wire v_452;
wire v_453;
wire v_454;
wire v_455;
wire v_456;
wire v_457;
wire v_458;
wire v_459;
wire v_460;
wire v_461;
wire v_462;
wire v_463;
wire v_464;
wire v_465;
wire v_466;
wire v_467;
wire v_468;
wire v_469;
wire v_470;
wire v_471;
wire v_472;
wire v_473;
wire v_474;
wire v_475;
wire v_476;
wire v_477;
wire v_478;
wire v_479;
wire v_480;
wire v_481;
wire v_482;
wire v_483;
wire v_484;
wire v_485;
wire v_486;
wire v_487;
wire v_488;
wire v_489;
wire v_490;
wire v_491;
wire v_492;
wire v_493;
wire v_494;
wire v_495;
wire v_496;
wire v_497;
wire v_498;
wire v_499;
wire v_500;
wire v_501;
wire v_502;
wire v_503;
wire v_504;
wire v_505;
wire v_506;
wire v_507;
wire v_508;
wire v_509;
wire v_510;
wire v_511;
wire v_512;
wire v_513;
wire v_514;
wire v_515;
wire v_516;
wire v_517;
wire v_518;
wire v_519;
wire v_520;
wire v_521;
wire v_522;
wire v_523;
wire v_524;
wire v_525;
wire v_526;
wire v_527;
wire v_528;
wire v_529;
wire v_530;
wire v_531;
wire v_532;
wire v_533;
wire v_534;
wire v_535;
wire v_536;
wire v_537;
wire v_538;
wire v_539;
wire v_540;
wire v_541;
wire v_542;
wire v_543;
wire v_544;
wire v_545;
wire v_546;
wire v_547;
wire v_548;
wire v_549;
wire v_550;
wire v_551;
wire v_552;
wire v_553;
wire v_554;
wire v_555;
wire v_556;
wire v_557;
wire v_558;
wire v_559;
wire v_560;
wire v_561;
wire v_562;
wire v_564;
wire v_565;
wire v_566;
wire v_567;
wire v_568;
wire v_569;
wire v_570;
wire v_571;
wire v_572;
wire v_573;
wire v_574;
wire v_575;
wire v_576;
wire v_577;
wire v_578;
wire v_579;
wire v_580;
wire v_581;
wire v_582;
wire v_583;
wire v_584;
wire v_585;
wire v_586;
wire v_587;
wire v_588;
wire v_589;
wire v_590;
wire v_591;
wire v_592;
wire v_593;
wire v_594;
wire v_595;
wire v_596;
wire v_597;
wire v_598;
wire v_599;
wire v_600;
wire v_601;
wire v_602;
wire v_603;
wire v_604;
wire v_605;
wire v_606;
wire v_607;
wire v_608;
wire v_609;
wire v_610;
wire v_611;
wire v_612;
wire v_613;
wire v_614;
wire v_615;
wire v_616;
wire v_617;
wire v_618;
wire v_619;
wire v_620;
wire v_621;
wire v_622;
wire v_623;
wire v_624;
wire v_625;
wire v_626;
wire v_627;
wire v_628;
wire v_629;
wire v_630;
wire v_631;
wire v_632;
wire v_633;
wire v_634;
wire v_635;
wire v_636;
wire v_637;
wire v_638;
wire v_639;
wire v_640;
wire v_641;
wire v_642;
wire v_643;
wire v_644;
wire v_645;
wire v_646;
wire v_647;
wire v_648;
wire v_649;
wire v_650;
wire v_651;
wire v_652;
wire v_653;
wire v_654;
wire v_655;
wire v_656;
wire v_657;
wire v_658;
wire v_659;
wire v_660;
wire v_661;
wire v_662;
wire v_663;
wire v_664;
wire v_665;
wire v_666;
wire v_667;
wire v_668;
wire v_669;
wire v_670;
wire v_671;
wire v_672;
wire v_673;
wire v_674;
wire v_675;
wire v_676;
wire v_677;
wire v_678;
wire v_679;
wire v_680;
wire v_681;
wire v_682;
wire v_683;
wire v_684;
wire v_685;
wire v_686;
wire v_687;
wire v_688;
wire v_689;
wire v_690;
wire v_691;
wire v_692;
wire v_693;
wire v_694;
wire v_695;
wire v_696;
wire v_697;
wire v_698;
wire v_699;
wire v_700;
wire v_701;
wire v_702;
wire v_703;
wire v_704;
wire v_705;
wire v_706;
wire v_707;
wire v_708;
wire v_709;
wire v_710;
wire v_711;
wire v_712;
wire v_713;
wire v_714;
wire v_715;
wire v_716;
wire v_717;
wire v_718;
wire v_719;
wire v_722;
wire v_723;
wire v_724;
wire v_725;
wire v_726;
wire v_727;
wire v_728;
wire v_729;
wire v_732;
wire v_733;
wire v_734;
wire v_735;
wire v_736;
wire v_737;
wire v_738;
wire v_739;
wire v_742;
wire v_743;
wire v_744;
wire v_745;
wire v_746;
wire v_747;
wire v_748;
wire v_749;
wire v_752;
wire v_753;
wire v_754;
wire v_755;
wire v_756;
wire v_757;
wire v_758;
wire v_759;
wire v_762;
wire v_763;
wire v_764;
wire v_765;
wire v_766;
wire v_767;
wire v_768;
wire v_769;
wire v_772;
wire v_773;
wire v_774;
wire v_775;
wire v_776;
wire v_777;
wire v_778;
wire v_779;
wire v_780;
wire v_781;
wire v_782;
wire v_783;
wire v_784;
wire v_785;
wire v_786;
wire v_787;
wire v_788;
wire v_789;
wire v_790;
wire v_791;
wire v_794;
wire v_795;
wire v_796;
wire v_797;
wire v_798;
wire v_799;
wire v_800;
wire v_801;
wire v_803;
wire v_805;
wire v_806;
wire v_808;
wire v_809;
wire v_810;
wire v_811;
wire v_812;
wire v_813;
wire v_814;
wire v_815;
wire v_816;
wire v_817;
wire v_818;
wire v_819;
wire v_820;
wire v_821;
wire v_822;
wire v_823;
wire v_824;
wire v_825;
wire v_826;
wire v_827;
wire v_828;
wire v_829;
wire v_830;
wire v_831;
wire v_832;
wire v_833;
wire v_834;
wire v_835;
wire v_836;
wire v_839;
wire v_840;
wire v_841;
wire v_842;
wire v_843;
wire v_844;
wire v_845;
wire v_846;
wire v_847;
wire v_848;
wire v_851;
wire v_852;
wire v_853;
wire v_854;
wire v_855;
wire v_856;
wire v_857;
wire v_858;
wire v_859;
wire v_860;
wire v_863;
wire v_864;
wire v_865;
wire v_866;
wire v_867;
wire v_868;
wire v_869;
wire v_870;
wire v_871;
wire v_872;
wire v_875;
wire v_876;
wire v_877;
wire v_878;
wire v_879;
wire v_880;
wire v_881;
wire v_882;
wire v_883;
wire v_884;
wire v_887;
wire v_888;
wire v_889;
wire v_890;
wire v_891;
wire v_892;
wire v_893;
wire v_894;
wire v_895;
wire v_896;
wire v_899;
wire v_900;
wire v_901;
wire v_902;
wire v_903;
wire v_904;
wire v_905;
wire v_906;
wire v_907;
wire v_908;
wire v_909;
wire v_910;
wire v_911;
wire v_912;
wire v_913;
wire v_914;
wire v_915;
wire v_916;
wire v_917;
wire v_918;
wire v_919;
wire v_920;
wire v_923;
wire v_924;
wire v_925;
wire v_926;
wire v_927;
wire v_928;
wire v_929;
wire v_930;
wire v_931;
wire v_932;
wire v_934;
wire v_935;
wire v_936;
wire v_937;
wire v_938;
wire v_939;
wire v_941;
wire v_942;
wire v_943;
wire v_944;
wire v_945;
wire v_946;
wire v_947;
wire v_948;
wire v_949;
wire v_950;
wire v_951;
wire v_952;
wire v_953;
wire v_954;
wire v_955;
wire v_956;
wire v_957;
wire v_958;
wire v_959;
wire v_960;
wire v_961;
wire v_962;
wire v_963;
wire v_964;
wire v_965;
wire v_966;
wire v_967;
wire v_968;
wire v_969;
wire v_970;
wire v_971;
wire v_972;
wire v_973;
wire v_974;
wire v_975;
wire v_976;
wire v_977;
wire v_978;
wire v_979;
wire v_980;
wire v_981;
wire v_982;
wire v_985;
wire v_986;
wire v_987;
wire v_988;
wire v_989;
wire v_990;
wire v_991;
wire v_992;
wire v_993;
wire v_994;
wire v_997;
wire v_998;
wire v_999;
wire v_1000;
wire v_1001;
wire v_1002;
wire v_1003;
wire v_1004;
wire v_1005;
wire v_1006;
wire v_1009;
wire v_1010;
wire v_1011;
wire v_1012;
wire v_1013;
wire v_1014;
wire v_1015;
wire v_1016;
wire v_1017;
wire v_1018;
wire v_1021;
wire v_1022;
wire v_1023;
wire v_1024;
wire v_1025;
wire v_1026;
wire v_1027;
wire v_1028;
wire v_1029;
wire v_1030;
wire v_1033;
wire v_1034;
wire v_1035;
wire v_1036;
wire v_1037;
wire v_1038;
wire v_1039;
wire v_1040;
wire v_1041;
wire v_1042;
wire v_1045;
wire v_1046;
wire v_1047;
wire v_1048;
wire v_1049;
wire v_1050;
wire v_1051;
wire v_1052;
wire v_1053;
wire v_1054;
wire v_1055;
wire v_1056;
wire v_1057;
wire v_1058;
wire v_1059;
wire v_1060;
wire v_1061;
wire v_1062;
wire v_1063;
wire v_1064;
wire v_1065;
wire v_1066;
wire v_1067;
wire v_1068;
wire v_1069;
wire v_1070;
wire v_1073;
wire v_1074;
wire v_1075;
wire v_1076;
wire v_1077;
wire v_1078;
wire v_1079;
wire v_1080;
wire v_1081;
wire v_1082;
wire v_1084;
wire v_1086;
wire v_1087;
wire v_1088;
wire v_1089;
wire v_1090;
wire v_1091;
wire v_1092;
wire v_1093;
wire v_1094;
wire v_1095;
wire v_1096;
wire v_1097;
wire v_1098;
wire v_1099;
wire v_1100;
wire v_1101;
wire v_1102;
wire v_1103;
wire v_1104;
wire v_1105;
wire v_1106;
wire v_1107;
wire v_1108;
wire v_1109;
wire v_1110;
wire v_1111;
wire v_1112;
wire v_1113;
wire v_1114;
wire v_1117;
wire v_1118;
wire v_1119;
wire v_1120;
wire v_1121;
wire v_1122;
wire v_1123;
wire v_1124;
wire v_1125;
wire v_1126;
wire v_1129;
wire v_1130;
wire v_1131;
wire v_1132;
wire v_1133;
wire v_1134;
wire v_1135;
wire v_1136;
wire v_1137;
wire v_1138;
wire v_1141;
wire v_1142;
wire v_1143;
wire v_1144;
wire v_1145;
wire v_1146;
wire v_1147;
wire v_1148;
wire v_1149;
wire v_1150;
wire v_1153;
wire v_1154;
wire v_1155;
wire v_1156;
wire v_1157;
wire v_1158;
wire v_1159;
wire v_1160;
wire v_1161;
wire v_1162;
wire v_1165;
wire v_1166;
wire v_1167;
wire v_1168;
wire v_1169;
wire v_1170;
wire v_1171;
wire v_1172;
wire v_1173;
wire v_1174;
wire v_1177;
wire v_1178;
wire v_1179;
wire v_1180;
wire v_1181;
wire v_1182;
wire v_1183;
wire v_1184;
wire v_1185;
wire v_1186;
wire v_1187;
wire v_1188;
wire v_1189;
wire v_1190;
wire v_1191;
wire v_1192;
wire v_1193;
wire v_1194;
wire v_1195;
wire v_1196;
wire v_1197;
wire v_1198;
wire v_1199;
wire v_1200;
wire v_1201;
wire v_1202;
wire v_1205;
wire v_1206;
wire v_1207;
wire v_1208;
wire v_1209;
wire v_1210;
wire v_1211;
wire v_1212;
wire v_1213;
wire v_1214;
wire v_1216;
wire v_1217;
wire v_1218;
wire v_1219;
wire v_1220;
wire v_1222;
wire v_1223;
wire v_1224;
wire v_1225;
wire v_1226;
wire v_1227;
wire v_1228;
wire v_1229;
wire v_1230;
wire v_1231;
wire v_1232;
wire v_1233;
wire v_1234;
wire v_1235;
wire v_1236;
wire v_1237;
wire v_1238;
wire v_1239;
wire v_1240;
wire v_1241;
wire v_1242;
wire v_1243;
wire v_1244;
wire v_1245;
wire v_1246;
wire v_1247;
wire v_1248;
wire v_1249;
wire v_1250;
wire v_1251;
wire v_1252;
wire v_1253;
wire v_1254;
wire v_1255;
wire v_1256;
wire v_1257;
wire v_1258;
wire v_1259;
wire v_1260;
wire v_1261;
wire v_1262;
wire v_1263;
wire v_1264;
wire v_1265;
wire v_1266;
wire v_1267;
wire v_1268;
wire v_1269;
wire v_1270;
wire v_1273;
wire v_1274;
wire v_1275;
wire v_1276;
wire v_1277;
wire v_1278;
wire v_1279;
wire v_1280;
wire v_1281;
wire v_1282;
wire v_1285;
wire v_1286;
wire v_1287;
wire v_1288;
wire v_1289;
wire v_1290;
wire v_1291;
wire v_1292;
wire v_1293;
wire v_1294;
wire v_1297;
wire v_1298;
wire v_1299;
wire v_1300;
wire v_1301;
wire v_1302;
wire v_1303;
wire v_1304;
wire v_1305;
wire v_1306;
wire v_1309;
wire v_1310;
wire v_1311;
wire v_1312;
wire v_1313;
wire v_1314;
wire v_1315;
wire v_1316;
wire v_1317;
wire v_1318;
wire v_1321;
wire v_1322;
wire v_1323;
wire v_1324;
wire v_1325;
wire v_1326;
wire v_1327;
wire v_1328;
wire v_1329;
wire v_1330;
wire v_1333;
wire v_1334;
wire v_1335;
wire v_1336;
wire v_1337;
wire v_1338;
wire v_1339;
wire v_1340;
wire v_1341;
wire v_1342;
wire v_1343;
wire v_1344;
wire v_1345;
wire v_1346;
wire v_1347;
wire v_1348;
wire v_1349;
wire v_1350;
wire v_1351;
wire v_1352;
wire v_1353;
wire v_1354;
wire v_1355;
wire v_1356;
wire v_1357;
wire v_1358;
wire v_1361;
wire v_1362;
wire v_1363;
wire v_1364;
wire v_1365;
wire v_1366;
wire v_1367;
wire v_1368;
wire v_1369;
wire v_1370;
wire v_1372;
wire v_1374;
wire v_1375;
wire v_1376;
wire v_1377;
wire v_1378;
wire v_1379;
wire v_1380;
wire v_1381;
wire v_1382;
wire v_1383;
wire v_1384;
wire v_1385;
wire v_1386;
wire v_1387;
wire v_1388;
wire v_1389;
wire v_1390;
wire v_1391;
wire v_1392;
wire v_1393;
wire v_1394;
wire v_1395;
wire v_1396;
wire v_1397;
wire v_1398;
wire v_1399;
wire v_1400;
wire v_1401;
wire v_1402;
wire v_1405;
wire v_1406;
wire v_1407;
wire v_1408;
wire v_1409;
wire v_1410;
wire v_1411;
wire v_1412;
wire v_1413;
wire v_1414;
wire v_1417;
wire v_1418;
wire v_1419;
wire v_1420;
wire v_1421;
wire v_1422;
wire v_1423;
wire v_1424;
wire v_1425;
wire v_1426;
wire v_1429;
wire v_1430;
wire v_1431;
wire v_1432;
wire v_1433;
wire v_1434;
wire v_1435;
wire v_1436;
wire v_1437;
wire v_1438;
wire v_1441;
wire v_1442;
wire v_1443;
wire v_1444;
wire v_1445;
wire v_1446;
wire v_1447;
wire v_1448;
wire v_1449;
wire v_1450;
wire v_1453;
wire v_1454;
wire v_1455;
wire v_1456;
wire v_1457;
wire v_1458;
wire v_1459;
wire v_1460;
wire v_1461;
wire v_1462;
wire v_1465;
wire v_1466;
wire v_1467;
wire v_1468;
wire v_1469;
wire v_1470;
wire v_1471;
wire v_1472;
wire v_1473;
wire v_1474;
wire v_1475;
wire v_1476;
wire v_1477;
wire v_1478;
wire v_1479;
wire v_1480;
wire v_1481;
wire v_1482;
wire v_1483;
wire v_1484;
wire v_1485;
wire v_1486;
wire v_1487;
wire v_1488;
wire v_1489;
wire v_1490;
wire v_1493;
wire v_1494;
wire v_1495;
wire v_1496;
wire v_1497;
wire v_1498;
wire v_1499;
wire v_1500;
wire v_1501;
wire v_1502;
wire v_1504;
wire v_1505;
wire v_1506;
wire v_1507;
wire v_1508;
wire v_1509;
wire v_1510;
wire v_1512;
wire v_1513;
wire v_1514;
wire v_1515;
wire v_1516;
wire v_1517;
wire v_1518;
wire v_1519;
wire v_1520;
wire v_1521;
wire v_1522;
wire v_1523;
wire v_1524;
wire v_1525;
wire v_1526;
wire v_1527;
wire v_1528;
wire v_1529;
wire v_1530;
wire v_1531;
wire v_1532;
wire v_1533;
wire v_1534;
wire v_1535;
wire v_1536;
wire v_1537;
wire v_1538;
wire v_1539;
wire v_1540;
wire v_1541;
wire v_1542;
wire v_1543;
wire v_1544;
wire v_1545;
wire v_1546;
wire v_1547;
wire v_1548;
wire v_1549;
wire v_1550;
wire v_1551;
wire v_1552;
wire v_1553;
wire v_1554;
wire v_1557;
wire v_1558;
wire v_1559;
wire v_1560;
wire v_1561;
wire v_1562;
wire v_1563;
wire v_1564;
wire v_1565;
wire v_1566;
wire v_1569;
wire v_1570;
wire v_1571;
wire v_1572;
wire v_1573;
wire v_1574;
wire v_1575;
wire v_1576;
wire v_1577;
wire v_1578;
wire v_1581;
wire v_1582;
wire v_1583;
wire v_1584;
wire v_1585;
wire v_1586;
wire v_1587;
wire v_1588;
wire v_1589;
wire v_1590;
wire v_1593;
wire v_1594;
wire v_1595;
wire v_1596;
wire v_1597;
wire v_1598;
wire v_1599;
wire v_1600;
wire v_1601;
wire v_1602;
wire v_1605;
wire v_1606;
wire v_1607;
wire v_1608;
wire v_1609;
wire v_1610;
wire v_1611;
wire v_1612;
wire v_1613;
wire v_1614;
wire v_1617;
wire v_1618;
wire v_1619;
wire v_1620;
wire v_1621;
wire v_1622;
wire v_1623;
wire v_1624;
wire v_1625;
wire v_1626;
wire v_1627;
wire v_1628;
wire v_1629;
wire v_1630;
wire v_1631;
wire v_1632;
wire v_1633;
wire v_1634;
wire v_1635;
wire v_1636;
wire v_1637;
wire v_1638;
wire v_1639;
wire v_1640;
wire v_1641;
wire v_1642;
wire v_1645;
wire v_1646;
wire v_1647;
wire v_1648;
wire v_1649;
wire v_1650;
wire v_1651;
wire v_1652;
wire v_1653;
wire v_1654;
wire v_1656;
wire v_1658;
wire v_1659;
wire v_1660;
wire v_1661;
wire v_1662;
wire v_1663;
wire v_1664;
wire v_1665;
wire v_1666;
wire v_1667;
wire v_1668;
wire v_1669;
wire v_1670;
wire v_1671;
wire v_1672;
wire v_1673;
wire v_1674;
wire v_1675;
wire v_1676;
wire v_1677;
wire v_1678;
wire v_1679;
wire v_1680;
wire v_1681;
wire v_1682;
wire v_1683;
wire v_1684;
wire v_1685;
wire v_1686;
wire v_1689;
wire v_1690;
wire v_1691;
wire v_1692;
wire v_1693;
wire v_1694;
wire v_1695;
wire v_1696;
wire v_1697;
wire v_1698;
wire v_1701;
wire v_1702;
wire v_1703;
wire v_1704;
wire v_1705;
wire v_1706;
wire v_1707;
wire v_1708;
wire v_1709;
wire v_1710;
wire v_1713;
wire v_1714;
wire v_1715;
wire v_1716;
wire v_1717;
wire v_1718;
wire v_1719;
wire v_1720;
wire v_1721;
wire v_1722;
wire v_1725;
wire v_1726;
wire v_1727;
wire v_1728;
wire v_1729;
wire v_1730;
wire v_1731;
wire v_1732;
wire v_1733;
wire v_1734;
wire v_1737;
wire v_1738;
wire v_1739;
wire v_1740;
wire v_1741;
wire v_1742;
wire v_1743;
wire v_1744;
wire v_1745;
wire v_1746;
wire v_1749;
wire v_1750;
wire v_1751;
wire v_1752;
wire v_1753;
wire v_1754;
wire v_1755;
wire v_1756;
wire v_1757;
wire v_1758;
wire v_1759;
wire v_1760;
wire v_1761;
wire v_1762;
wire v_1763;
wire v_1764;
wire v_1765;
wire v_1766;
wire v_1767;
wire v_1768;
wire v_1769;
wire v_1770;
wire v_1771;
wire v_1772;
wire v_1773;
wire v_1774;
wire v_1777;
wire v_1778;
wire v_1779;
wire v_1780;
wire v_1781;
wire v_1782;
wire v_1783;
wire v_1784;
wire v_1785;
wire v_1786;
wire v_1788;
wire v_1789;
wire v_1790;
wire v_1791;
wire v_1792;
wire v_1794;
wire v_1795;
wire v_1796;
wire v_1797;
wire v_1798;
wire v_1799;
wire v_1800;
wire v_1801;
wire v_1802;
wire v_1803;
wire v_1804;
wire v_1805;
wire v_1806;
wire v_1807;
wire v_1808;
wire v_1809;
wire v_1810;
wire v_1811;
wire v_1812;
wire v_1813;
wire v_1814;
wire v_1815;
wire v_1816;
wire v_1817;
wire v_1818;
wire v_1819;
wire v_1820;
wire v_1821;
wire v_1822;
wire v_1823;
wire v_1824;
wire v_1825;
wire v_1826;
wire v_1827;
wire v_1828;
wire v_1829;
wire v_1830;
wire v_1831;
wire v_1832;
wire v_1833;
wire v_1834;
wire v_1835;
wire v_1836;
wire v_1837;
wire v_1838;
wire v_1839;
wire v_1840;
wire v_1841;
wire v_1842;
wire v_1843;
wire v_1844;
wire v_1845;
wire v_1846;
wire v_1847;
wire v_1848;
wire v_1849;
wire v_1850;
wire v_1853;
wire v_1854;
wire v_1855;
wire v_1856;
wire v_1857;
wire v_1858;
wire v_1859;
wire v_1860;
wire v_1861;
wire v_1862;
wire v_1865;
wire v_1866;
wire v_1867;
wire v_1868;
wire v_1869;
wire v_1870;
wire v_1871;
wire v_1872;
wire v_1873;
wire v_1874;
wire v_1877;
wire v_1878;
wire v_1879;
wire v_1880;
wire v_1881;
wire v_1882;
wire v_1883;
wire v_1884;
wire v_1885;
wire v_1886;
wire v_1889;
wire v_1890;
wire v_1891;
wire v_1892;
wire v_1893;
wire v_1894;
wire v_1895;
wire v_1896;
wire v_1897;
wire v_1898;
wire v_1901;
wire v_1902;
wire v_1903;
wire v_1904;
wire v_1905;
wire v_1906;
wire v_1907;
wire v_1908;
wire v_1909;
wire v_1910;
wire v_1913;
wire v_1914;
wire v_1915;
wire v_1916;
wire v_1917;
wire v_1918;
wire v_1919;
wire v_1920;
wire v_1921;
wire v_1922;
wire v_1923;
wire v_1924;
wire v_1925;
wire v_1926;
wire v_1927;
wire v_1928;
wire v_1929;
wire v_1930;
wire v_1931;
wire v_1932;
wire v_1933;
wire v_1934;
wire v_1935;
wire v_1936;
wire v_1937;
wire v_1938;
wire v_1941;
wire v_1942;
wire v_1943;
wire v_1944;
wire v_1945;
wire v_1946;
wire v_1947;
wire v_1948;
wire v_1949;
wire v_1950;
wire v_1952;
wire v_1954;
wire v_1955;
wire v_1956;
wire v_1957;
wire v_1958;
wire v_1959;
wire v_1960;
wire v_1961;
wire v_1962;
wire v_1963;
wire v_1964;
wire v_1965;
wire v_1966;
wire v_1967;
wire v_1968;
wire v_1969;
wire v_1970;
wire v_1971;
wire v_1972;
wire v_1973;
wire v_1974;
wire v_1975;
wire v_1976;
wire v_1977;
wire v_1978;
wire v_1979;
wire v_1980;
wire v_1981;
wire v_1982;
wire v_1985;
wire v_1986;
wire v_1987;
wire v_1988;
wire v_1989;
wire v_1990;
wire v_1991;
wire v_1992;
wire v_1993;
wire v_1994;
wire v_1997;
wire v_1998;
wire v_1999;
wire v_2000;
wire v_2001;
wire v_2002;
wire v_2003;
wire v_2004;
wire v_2005;
wire v_2006;
wire v_2009;
wire v_2010;
wire v_2011;
wire v_2012;
wire v_2013;
wire v_2014;
wire v_2015;
wire v_2016;
wire v_2017;
wire v_2018;
wire v_2021;
wire v_2022;
wire v_2023;
wire v_2024;
wire v_2025;
wire v_2026;
wire v_2027;
wire v_2028;
wire v_2029;
wire v_2030;
wire v_2033;
wire v_2034;
wire v_2035;
wire v_2036;
wire v_2037;
wire v_2038;
wire v_2039;
wire v_2040;
wire v_2041;
wire v_2042;
wire v_2045;
wire v_2046;
wire v_2047;
wire v_2048;
wire v_2049;
wire v_2050;
wire v_2051;
wire v_2052;
wire v_2053;
wire v_2054;
wire v_2055;
wire v_2056;
wire v_2057;
wire v_2058;
wire v_2059;
wire v_2060;
wire v_2061;
wire v_2062;
wire v_2063;
wire v_2064;
wire v_2065;
wire v_2066;
wire v_2067;
wire v_2068;
wire v_2069;
wire v_2070;
wire v_2073;
wire v_2074;
wire v_2075;
wire v_2076;
wire v_2077;
wire v_2078;
wire v_2079;
wire v_2080;
wire v_2081;
wire v_2082;
wire v_2084;
wire v_2085;
wire v_2086;
wire v_2087;
wire v_2088;
wire v_2089;
wire v_2091;
wire v_2092;
wire v_2093;
wire v_2094;
wire v_2095;
wire v_2096;
wire v_2097;
wire v_2098;
wire v_2099;
wire v_2100;
wire v_2101;
wire v_2102;
wire v_2103;
wire v_2104;
wire v_2105;
wire v_2106;
wire v_2107;
wire v_2108;
wire v_2109;
wire v_2110;
wire v_2111;
wire v_2112;
wire v_2113;
wire v_2114;
wire v_2115;
wire v_2116;
wire v_2117;
wire v_2118;
wire v_2119;
wire v_2120;
wire v_2121;
wire v_2122;
wire v_2123;
wire v_2124;
wire v_2125;
wire v_2126;
wire v_2127;
wire v_2128;
wire v_2129;
wire v_2130;
wire v_2131;
wire v_2132;
wire v_2135;
wire v_2136;
wire v_2137;
wire v_2138;
wire v_2139;
wire v_2140;
wire v_2141;
wire v_2142;
wire v_2143;
wire v_2144;
wire v_2147;
wire v_2148;
wire v_2149;
wire v_2150;
wire v_2151;
wire v_2152;
wire v_2153;
wire v_2154;
wire v_2155;
wire v_2156;
wire v_2159;
wire v_2160;
wire v_2161;
wire v_2162;
wire v_2163;
wire v_2164;
wire v_2165;
wire v_2166;
wire v_2167;
wire v_2168;
wire v_2171;
wire v_2172;
wire v_2173;
wire v_2174;
wire v_2175;
wire v_2176;
wire v_2177;
wire v_2178;
wire v_2179;
wire v_2180;
wire v_2183;
wire v_2184;
wire v_2185;
wire v_2186;
wire v_2187;
wire v_2188;
wire v_2189;
wire v_2190;
wire v_2191;
wire v_2192;
wire v_2195;
wire v_2196;
wire v_2197;
wire v_2198;
wire v_2199;
wire v_2200;
wire v_2201;
wire v_2202;
wire v_2203;
wire v_2204;
wire v_2205;
wire v_2206;
wire v_2207;
wire v_2208;
wire v_2209;
wire v_2210;
wire v_2211;
wire v_2212;
wire v_2213;
wire v_2214;
wire v_2215;
wire v_2216;
wire v_2217;
wire v_2218;
wire v_2219;
wire v_2220;
wire v_2223;
wire v_2224;
wire v_2225;
wire v_2226;
wire v_2227;
wire v_2228;
wire v_2229;
wire v_2230;
wire v_2231;
wire v_2232;
wire v_2234;
wire v_2236;
wire v_2237;
wire v_2238;
wire v_2239;
wire v_2240;
wire v_2241;
wire v_2242;
wire v_2243;
wire v_2244;
wire v_2245;
wire v_2246;
wire v_2247;
wire v_2248;
wire v_2249;
wire v_2250;
wire v_2251;
wire v_2252;
wire v_2253;
wire v_2254;
wire v_2255;
wire v_2256;
wire v_2257;
wire v_2258;
wire v_2259;
wire v_2260;
wire v_2261;
wire v_2262;
wire v_2263;
wire v_2264;
wire v_2267;
wire v_2268;
wire v_2269;
wire v_2270;
wire v_2271;
wire v_2272;
wire v_2273;
wire v_2274;
wire v_2275;
wire v_2276;
wire v_2279;
wire v_2280;
wire v_2281;
wire v_2282;
wire v_2283;
wire v_2284;
wire v_2285;
wire v_2286;
wire v_2287;
wire v_2288;
wire v_2291;
wire v_2292;
wire v_2293;
wire v_2294;
wire v_2295;
wire v_2296;
wire v_2297;
wire v_2298;
wire v_2299;
wire v_2300;
wire v_2303;
wire v_2304;
wire v_2305;
wire v_2306;
wire v_2307;
wire v_2308;
wire v_2309;
wire v_2310;
wire v_2311;
wire v_2312;
wire v_2315;
wire v_2316;
wire v_2317;
wire v_2318;
wire v_2319;
wire v_2320;
wire v_2321;
wire v_2322;
wire v_2323;
wire v_2324;
wire v_2327;
wire v_2328;
wire v_2329;
wire v_2330;
wire v_2331;
wire v_2332;
wire v_2333;
wire v_2334;
wire v_2335;
wire v_2336;
wire v_2337;
wire v_2338;
wire v_2339;
wire v_2340;
wire v_2341;
wire v_2342;
wire v_2343;
wire v_2344;
wire v_2345;
wire v_2346;
wire v_2347;
wire v_2348;
wire v_2349;
wire v_2350;
wire v_2351;
wire v_2352;
wire v_2355;
wire v_2356;
wire v_2357;
wire v_2358;
wire v_2359;
wire v_2360;
wire v_2361;
wire v_2362;
wire v_2363;
wire v_2364;
wire v_2366;
wire v_2367;
wire v_2368;
wire v_2369;
wire v_2370;
wire v_2372;
wire v_2373;
wire v_2374;
wire v_2375;
wire v_2376;
wire v_2377;
wire v_2378;
wire v_2379;
wire v_2380;
wire v_2381;
wire v_2382;
wire v_2383;
wire v_2384;
wire v_2385;
wire v_2386;
wire v_2387;
wire v_2388;
wire v_2389;
wire v_2390;
wire v_2391;
wire v_2392;
wire v_2393;
wire v_2394;
wire v_2395;
wire v_2396;
wire v_2397;
wire v_2398;
wire v_2399;
wire v_2400;
wire v_2401;
wire v_2402;
wire v_2403;
wire v_2404;
wire v_2405;
wire v_2406;
wire v_2407;
wire v_2408;
wire v_2409;
wire v_2410;
wire v_2411;
wire v_2412;
wire v_2413;
wire v_2414;
wire v_2415;
wire v_2416;
wire v_2417;
wire v_2418;
wire v_2419;
wire v_2420;
wire v_2423;
wire v_2424;
wire v_2425;
wire v_2426;
wire v_2427;
wire v_2428;
wire v_2429;
wire v_2430;
wire v_2431;
wire v_2432;
wire v_2435;
wire v_2436;
wire v_2437;
wire v_2438;
wire v_2439;
wire v_2440;
wire v_2441;
wire v_2442;
wire v_2443;
wire v_2444;
wire v_2447;
wire v_2448;
wire v_2449;
wire v_2450;
wire v_2451;
wire v_2452;
wire v_2453;
wire v_2454;
wire v_2455;
wire v_2456;
wire v_2459;
wire v_2460;
wire v_2461;
wire v_2462;
wire v_2463;
wire v_2464;
wire v_2465;
wire v_2466;
wire v_2467;
wire v_2468;
wire v_2471;
wire v_2472;
wire v_2473;
wire v_2474;
wire v_2475;
wire v_2476;
wire v_2477;
wire v_2478;
wire v_2479;
wire v_2480;
wire v_2483;
wire v_2484;
wire v_2485;
wire v_2486;
wire v_2487;
wire v_2488;
wire v_2489;
wire v_2490;
wire v_2491;
wire v_2492;
wire v_2493;
wire v_2494;
wire v_2495;
wire v_2496;
wire v_2497;
wire v_2498;
wire v_2499;
wire v_2500;
wire v_2501;
wire v_2502;
wire v_2503;
wire v_2504;
wire v_2505;
wire v_2506;
wire v_2507;
wire v_2508;
wire v_2511;
wire v_2512;
wire v_2513;
wire v_2514;
wire v_2515;
wire v_2516;
wire v_2517;
wire v_2518;
wire v_2519;
wire v_2520;
wire v_2522;
wire v_2524;
wire v_2525;
wire v_2526;
wire v_2527;
wire v_2528;
wire v_2529;
wire v_2530;
wire v_2531;
wire v_2532;
wire v_2533;
wire v_2534;
wire v_2535;
wire v_2536;
wire v_2537;
wire v_2538;
wire v_2539;
wire v_2540;
wire v_2541;
wire v_2542;
wire v_2543;
wire v_2544;
wire v_2545;
wire v_2546;
wire v_2547;
wire v_2548;
wire v_2549;
wire v_2550;
wire v_2551;
wire v_2552;
wire v_2555;
wire v_2556;
wire v_2557;
wire v_2558;
wire v_2559;
wire v_2560;
wire v_2561;
wire v_2562;
wire v_2563;
wire v_2564;
wire v_2567;
wire v_2568;
wire v_2569;
wire v_2570;
wire v_2571;
wire v_2572;
wire v_2573;
wire v_2574;
wire v_2575;
wire v_2576;
wire v_2579;
wire v_2580;
wire v_2581;
wire v_2582;
wire v_2583;
wire v_2584;
wire v_2585;
wire v_2586;
wire v_2587;
wire v_2588;
wire v_2591;
wire v_2592;
wire v_2593;
wire v_2594;
wire v_2595;
wire v_2596;
wire v_2597;
wire v_2598;
wire v_2599;
wire v_2600;
wire v_2603;
wire v_2604;
wire v_2605;
wire v_2606;
wire v_2607;
wire v_2608;
wire v_2609;
wire v_2610;
wire v_2611;
wire v_2612;
wire v_2615;
wire v_2616;
wire v_2617;
wire v_2618;
wire v_2619;
wire v_2620;
wire v_2621;
wire v_2622;
wire v_2623;
wire v_2624;
wire v_2625;
wire v_2626;
wire v_2627;
wire v_2628;
wire v_2629;
wire v_2630;
wire v_2631;
wire v_2632;
wire v_2633;
wire v_2634;
wire v_2635;
wire v_2636;
wire v_2637;
wire v_2638;
wire v_2639;
wire v_2640;
wire v_2643;
wire v_2644;
wire v_2645;
wire v_2646;
wire v_2647;
wire v_2648;
wire v_2649;
wire v_2650;
wire v_2651;
wire v_2652;
wire v_2654;
wire v_2655;
wire v_2656;
wire v_2657;
wire v_2658;
wire v_2659;
wire v_2660;
wire v_2661;
wire v_2663;
wire v_2664;
wire v_2665;
wire v_2666;
wire v_2667;
wire v_2668;
wire v_2669;
wire v_2670;
wire v_2671;
wire v_2672;
wire v_2673;
wire v_2674;
wire v_2675;
wire v_2676;
wire v_2677;
wire v_2678;
wire v_2679;
wire v_2680;
wire v_2681;
wire v_2682;
wire v_2683;
wire v_2684;
wire v_2685;
wire v_2686;
wire v_2687;
wire v_2688;
wire v_2689;
wire v_2690;
wire v_2691;
wire v_2692;
wire v_2693;
wire v_2694;
wire v_2695;
wire v_2696;
wire v_2697;
wire v_2698;
wire v_2699;
wire v_2700;
wire v_2701;
wire v_2702;
wire v_2703;
wire v_2704;
wire v_2705;
wire v_2706;
wire v_2709;
wire v_2710;
wire v_2711;
wire v_2712;
wire v_2713;
wire v_2714;
wire v_2715;
wire v_2716;
wire v_2717;
wire v_2718;
wire v_2721;
wire v_2722;
wire v_2723;
wire v_2724;
wire v_2725;
wire v_2726;
wire v_2727;
wire v_2728;
wire v_2729;
wire v_2730;
wire v_2733;
wire v_2734;
wire v_2735;
wire v_2736;
wire v_2737;
wire v_2738;
wire v_2739;
wire v_2740;
wire v_2741;
wire v_2742;
wire v_2745;
wire v_2746;
wire v_2747;
wire v_2748;
wire v_2749;
wire v_2750;
wire v_2751;
wire v_2752;
wire v_2753;
wire v_2754;
wire v_2757;
wire v_2758;
wire v_2759;
wire v_2760;
wire v_2761;
wire v_2762;
wire v_2763;
wire v_2764;
wire v_2765;
wire v_2766;
wire v_2769;
wire v_2770;
wire v_2771;
wire v_2772;
wire v_2773;
wire v_2774;
wire v_2775;
wire v_2776;
wire v_2777;
wire v_2778;
wire v_2779;
wire v_2780;
wire v_2781;
wire v_2782;
wire v_2783;
wire v_2784;
wire v_2785;
wire v_2786;
wire v_2787;
wire v_2788;
wire v_2789;
wire v_2790;
wire v_2791;
wire v_2792;
wire v_2793;
wire v_2794;
wire v_2797;
wire v_2798;
wire v_2799;
wire v_2800;
wire v_2801;
wire v_2802;
wire v_2803;
wire v_2804;
wire v_2805;
wire v_2806;
wire v_2808;
wire v_2810;
wire v_2811;
wire v_2812;
wire v_2813;
wire v_2814;
wire v_2815;
wire v_2816;
wire v_2817;
wire v_2818;
wire v_2819;
wire v_2820;
wire v_2821;
wire v_2822;
wire v_2823;
wire v_2824;
wire v_2825;
wire v_2826;
wire v_2827;
wire v_2828;
wire v_2829;
wire v_2830;
wire v_2831;
wire v_2832;
wire v_2833;
wire v_2834;
wire v_2835;
wire v_2836;
wire v_2837;
wire v_2838;
wire v_2841;
wire v_2842;
wire v_2843;
wire v_2844;
wire v_2845;
wire v_2846;
wire v_2847;
wire v_2848;
wire v_2849;
wire v_2850;
wire v_2853;
wire v_2854;
wire v_2855;
wire v_2856;
wire v_2857;
wire v_2858;
wire v_2859;
wire v_2860;
wire v_2861;
wire v_2862;
wire v_2865;
wire v_2866;
wire v_2867;
wire v_2868;
wire v_2869;
wire v_2870;
wire v_2871;
wire v_2872;
wire v_2873;
wire v_2874;
wire v_2877;
wire v_2878;
wire v_2879;
wire v_2880;
wire v_2881;
wire v_2882;
wire v_2883;
wire v_2884;
wire v_2885;
wire v_2886;
wire v_2889;
wire v_2890;
wire v_2891;
wire v_2892;
wire v_2893;
wire v_2894;
wire v_2895;
wire v_2896;
wire v_2897;
wire v_2898;
wire v_2901;
wire v_2902;
wire v_2903;
wire v_2904;
wire v_2905;
wire v_2906;
wire v_2907;
wire v_2908;
wire v_2909;
wire v_2910;
wire v_2911;
wire v_2912;
wire v_2913;
wire v_2914;
wire v_2915;
wire v_2916;
wire v_2917;
wire v_2918;
wire v_2919;
wire v_2920;
wire v_2921;
wire v_2922;
wire v_2923;
wire v_2924;
wire v_2925;
wire v_2926;
wire v_2929;
wire v_2930;
wire v_2931;
wire v_2932;
wire v_2933;
wire v_2934;
wire v_2935;
wire v_2936;
wire v_2937;
wire v_2938;
wire v_2940;
wire v_2941;
wire v_2942;
wire v_2943;
wire v_2944;
wire v_2946;
wire v_2947;
wire v_2948;
wire v_2949;
wire v_2950;
wire v_2951;
wire v_2952;
wire v_2953;
wire v_2954;
wire v_2955;
wire v_2956;
wire v_2957;
wire v_2958;
wire v_2959;
wire v_2960;
wire v_2961;
wire v_2962;
wire v_2963;
wire v_2964;
wire v_2965;
wire v_2966;
wire v_2967;
wire v_2968;
wire v_2969;
wire v_2970;
wire v_2971;
wire v_2972;
wire v_2973;
wire v_2974;
wire v_2975;
wire v_2976;
wire v_2977;
wire v_2978;
wire v_2979;
wire v_2980;
wire v_2981;
wire v_2982;
wire v_2983;
wire v_2984;
wire v_2985;
wire v_2986;
wire v_2987;
wire v_2988;
wire v_2989;
wire v_2990;
wire v_2991;
wire v_2992;
wire v_2993;
wire v_2994;
wire v_2995;
wire v_2996;
wire v_2997;
wire v_2998;
wire v_2999;
wire v_3000;
wire v_3001;
wire v_3002;
wire v_3003;
wire v_3004;
wire v_3005;
wire v_3006;
wire v_3007;
wire v_3008;
wire v_3009;
wire v_3010;
wire v_3013;
wire v_3014;
wire v_3015;
wire v_3016;
wire v_3017;
wire v_3018;
wire v_3019;
wire v_3020;
wire v_3021;
wire v_3022;
wire v_3025;
wire v_3026;
wire v_3027;
wire v_3028;
wire v_3029;
wire v_3030;
wire v_3031;
wire v_3032;
wire v_3033;
wire v_3034;
wire v_3037;
wire v_3038;
wire v_3039;
wire v_3040;
wire v_3041;
wire v_3042;
wire v_3043;
wire v_3044;
wire v_3045;
wire v_3046;
wire v_3049;
wire v_3050;
wire v_3051;
wire v_3052;
wire v_3053;
wire v_3054;
wire v_3055;
wire v_3056;
wire v_3057;
wire v_3058;
wire v_3061;
wire v_3062;
wire v_3063;
wire v_3064;
wire v_3065;
wire v_3066;
wire v_3067;
wire v_3068;
wire v_3069;
wire v_3070;
wire v_3073;
wire v_3074;
wire v_3075;
wire v_3076;
wire v_3077;
wire v_3078;
wire v_3079;
wire v_3080;
wire v_3081;
wire v_3082;
wire v_3083;
wire v_3084;
wire v_3085;
wire v_3086;
wire v_3087;
wire v_3088;
wire v_3089;
wire v_3090;
wire v_3091;
wire v_3092;
wire v_3093;
wire v_3094;
wire v_3095;
wire v_3096;
wire v_3097;
wire v_3098;
wire v_3101;
wire v_3102;
wire v_3103;
wire v_3104;
wire v_3105;
wire v_3106;
wire v_3107;
wire v_3108;
wire v_3109;
wire v_3110;
wire v_3112;
wire v_3114;
wire v_3115;
wire v_3116;
wire v_3117;
wire v_3118;
wire v_3119;
wire v_3120;
wire v_3121;
wire v_3122;
wire v_3123;
wire v_3124;
wire v_3125;
wire v_3126;
wire v_3127;
wire v_3128;
wire v_3129;
wire v_3130;
wire v_3131;
wire v_3132;
wire v_3133;
wire v_3134;
wire v_3135;
wire v_3136;
wire v_3137;
wire v_3138;
wire v_3139;
wire v_3140;
wire v_3141;
wire v_3142;
wire v_3145;
wire v_3146;
wire v_3147;
wire v_3148;
wire v_3149;
wire v_3150;
wire v_3151;
wire v_3152;
wire v_3153;
wire v_3154;
wire v_3157;
wire v_3158;
wire v_3159;
wire v_3160;
wire v_3161;
wire v_3162;
wire v_3163;
wire v_3164;
wire v_3165;
wire v_3166;
wire v_3169;
wire v_3170;
wire v_3171;
wire v_3172;
wire v_3173;
wire v_3174;
wire v_3175;
wire v_3176;
wire v_3177;
wire v_3178;
wire v_3181;
wire v_3182;
wire v_3183;
wire v_3184;
wire v_3185;
wire v_3186;
wire v_3187;
wire v_3188;
wire v_3189;
wire v_3190;
wire v_3193;
wire v_3194;
wire v_3195;
wire v_3196;
wire v_3197;
wire v_3198;
wire v_3199;
wire v_3200;
wire v_3201;
wire v_3202;
wire v_3205;
wire v_3206;
wire v_3207;
wire v_3208;
wire v_3209;
wire v_3210;
wire v_3211;
wire v_3212;
wire v_3213;
wire v_3214;
wire v_3215;
wire v_3216;
wire v_3217;
wire v_3218;
wire v_3219;
wire v_3220;
wire v_3221;
wire v_3222;
wire v_3223;
wire v_3224;
wire v_3225;
wire v_3226;
wire v_3227;
wire v_3228;
wire v_3229;
wire v_3230;
wire v_3233;
wire v_3234;
wire v_3235;
wire v_3236;
wire v_3237;
wire v_3238;
wire v_3239;
wire v_3240;
wire v_3241;
wire v_3242;
wire v_3244;
wire v_3245;
wire v_3246;
wire v_3247;
wire v_3248;
wire v_3249;
wire v_3251;
wire v_3252;
wire v_3253;
wire v_3254;
wire v_3255;
wire v_3256;
wire v_3257;
wire v_3258;
wire v_3259;
wire v_3260;
wire v_3261;
wire v_3262;
wire v_3263;
wire v_3264;
wire v_3265;
wire v_3266;
wire v_3267;
wire v_3268;
wire v_3269;
wire v_3270;
wire v_3271;
wire v_3272;
wire v_3273;
wire v_3274;
wire v_3275;
wire v_3276;
wire v_3277;
wire v_3278;
wire v_3279;
wire v_3280;
wire v_3281;
wire v_3282;
wire v_3283;
wire v_3284;
wire v_3285;
wire v_3286;
wire v_3287;
wire v_3288;
wire v_3289;
wire v_3290;
wire v_3291;
wire v_3292;
wire v_3295;
wire v_3296;
wire v_3297;
wire v_3298;
wire v_3299;
wire v_3300;
wire v_3301;
wire v_3302;
wire v_3303;
wire v_3304;
wire v_3307;
wire v_3308;
wire v_3309;
wire v_3310;
wire v_3311;
wire v_3312;
wire v_3313;
wire v_3314;
wire v_3315;
wire v_3316;
wire v_3319;
wire v_3320;
wire v_3321;
wire v_3322;
wire v_3323;
wire v_3324;
wire v_3325;
wire v_3326;
wire v_3327;
wire v_3328;
wire v_3331;
wire v_3332;
wire v_3333;
wire v_3334;
wire v_3335;
wire v_3336;
wire v_3337;
wire v_3338;
wire v_3339;
wire v_3340;
wire v_3343;
wire v_3344;
wire v_3345;
wire v_3346;
wire v_3347;
wire v_3348;
wire v_3349;
wire v_3350;
wire v_3351;
wire v_3352;
wire v_3355;
wire v_3356;
wire v_3357;
wire v_3358;
wire v_3359;
wire v_3360;
wire v_3361;
wire v_3362;
wire v_3363;
wire v_3364;
wire v_3365;
wire v_3366;
wire v_3367;
wire v_3368;
wire v_3369;
wire v_3370;
wire v_3371;
wire v_3372;
wire v_3373;
wire v_3374;
wire v_3375;
wire v_3376;
wire v_3377;
wire v_3378;
wire v_3379;
wire v_3380;
wire v_3383;
wire v_3384;
wire v_3385;
wire v_3386;
wire v_3387;
wire v_3388;
wire v_3389;
wire v_3390;
wire v_3391;
wire v_3392;
wire v_3394;
wire v_3396;
wire v_3397;
wire v_3398;
wire v_3399;
wire v_3400;
wire v_3401;
wire v_3402;
wire v_3403;
wire v_3404;
wire v_3405;
wire v_3406;
wire v_3407;
wire v_3408;
wire v_3409;
wire v_3410;
wire v_3411;
wire v_3412;
wire v_3413;
wire v_3414;
wire v_3415;
wire v_3416;
wire v_3417;
wire v_3418;
wire v_3419;
wire v_3420;
wire v_3421;
wire v_3422;
wire v_3423;
wire v_3424;
wire v_3427;
wire v_3428;
wire v_3429;
wire v_3430;
wire v_3431;
wire v_3432;
wire v_3433;
wire v_3434;
wire v_3435;
wire v_3436;
wire v_3439;
wire v_3440;
wire v_3441;
wire v_3442;
wire v_3443;
wire v_3444;
wire v_3445;
wire v_3446;
wire v_3447;
wire v_3448;
wire v_3451;
wire v_3452;
wire v_3453;
wire v_3454;
wire v_3455;
wire v_3456;
wire v_3457;
wire v_3458;
wire v_3459;
wire v_3460;
wire v_3463;
wire v_3464;
wire v_3465;
wire v_3466;
wire v_3467;
wire v_3468;
wire v_3469;
wire v_3470;
wire v_3471;
wire v_3472;
wire v_3475;
wire v_3476;
wire v_3477;
wire v_3478;
wire v_3479;
wire v_3480;
wire v_3481;
wire v_3482;
wire v_3483;
wire v_3484;
wire v_3487;
wire v_3488;
wire v_3489;
wire v_3490;
wire v_3491;
wire v_3492;
wire v_3493;
wire v_3494;
wire v_3495;
wire v_3496;
wire v_3497;
wire v_3498;
wire v_3499;
wire v_3500;
wire v_3501;
wire v_3502;
wire v_3503;
wire v_3504;
wire v_3505;
wire v_3506;
wire v_3507;
wire v_3508;
wire v_3509;
wire v_3510;
wire v_3511;
wire v_3512;
wire v_3515;
wire v_3516;
wire v_3517;
wire v_3518;
wire v_3519;
wire v_3520;
wire v_3521;
wire v_3522;
wire v_3523;
wire v_3524;
wire v_3526;
wire v_3527;
wire v_3528;
wire v_3529;
wire v_3530;
wire v_3532;
wire v_3533;
wire v_3534;
wire v_3535;
wire v_3536;
wire v_3537;
wire v_3538;
wire v_3539;
wire v_3540;
wire v_3541;
wire v_3542;
wire v_3543;
wire v_3544;
wire v_3545;
wire v_3546;
wire v_3547;
wire v_3548;
wire v_3549;
wire v_3550;
wire v_3551;
wire v_3552;
wire v_3553;
wire v_3554;
wire v_3555;
wire v_3556;
wire v_3557;
wire v_3558;
wire v_3559;
wire v_3560;
wire v_3561;
wire v_3562;
wire v_3563;
wire v_3564;
wire v_3565;
wire v_3566;
wire v_3567;
wire v_3568;
wire v_3569;
wire v_3570;
wire v_3571;
wire v_3572;
wire v_3573;
wire v_3574;
wire v_3575;
wire v_3576;
wire v_3577;
wire v_3578;
wire v_3579;
wire v_3580;
wire v_3583;
wire v_3584;
wire v_3585;
wire v_3586;
wire v_3587;
wire v_3588;
wire v_3589;
wire v_3590;
wire v_3591;
wire v_3592;
wire v_3595;
wire v_3596;
wire v_3597;
wire v_3598;
wire v_3599;
wire v_3600;
wire v_3601;
wire v_3602;
wire v_3603;
wire v_3604;
wire v_3607;
wire v_3608;
wire v_3609;
wire v_3610;
wire v_3611;
wire v_3612;
wire v_3613;
wire v_3614;
wire v_3615;
wire v_3616;
wire v_3619;
wire v_3620;
wire v_3621;
wire v_3622;
wire v_3623;
wire v_3624;
wire v_3625;
wire v_3626;
wire v_3627;
wire v_3628;
wire v_3631;
wire v_3632;
wire v_3633;
wire v_3634;
wire v_3635;
wire v_3636;
wire v_3637;
wire v_3638;
wire v_3639;
wire v_3640;
wire v_3643;
wire v_3644;
wire v_3645;
wire v_3646;
wire v_3647;
wire v_3648;
wire v_3649;
wire v_3650;
wire v_3651;
wire v_3652;
wire v_3653;
wire v_3654;
wire v_3655;
wire v_3656;
wire v_3657;
wire v_3658;
wire v_3659;
wire v_3660;
wire v_3661;
wire v_3662;
wire v_3663;
wire v_3664;
wire v_3665;
wire v_3666;
wire v_3667;
wire v_3668;
wire v_3671;
wire v_3672;
wire v_3673;
wire v_3674;
wire v_3675;
wire v_3676;
wire v_3677;
wire v_3678;
wire v_3679;
wire v_3680;
wire v_3682;
wire v_3684;
wire v_3685;
wire v_3686;
wire v_3687;
wire v_3688;
wire v_3689;
wire v_3690;
wire v_3691;
wire v_3692;
wire v_3693;
wire v_3694;
wire v_3695;
wire v_3696;
wire v_3697;
wire v_3698;
wire v_3699;
wire v_3700;
wire v_3701;
wire v_3702;
wire v_3703;
wire v_3704;
wire v_3705;
wire v_3706;
wire v_3707;
wire v_3708;
wire v_3709;
wire v_3710;
wire v_3711;
wire v_3712;
wire v_3715;
wire v_3716;
wire v_3717;
wire v_3718;
wire v_3719;
wire v_3720;
wire v_3721;
wire v_3722;
wire v_3723;
wire v_3724;
wire v_3727;
wire v_3728;
wire v_3729;
wire v_3730;
wire v_3731;
wire v_3732;
wire v_3733;
wire v_3734;
wire v_3735;
wire v_3736;
wire v_3739;
wire v_3740;
wire v_3741;
wire v_3742;
wire v_3743;
wire v_3744;
wire v_3745;
wire v_3746;
wire v_3747;
wire v_3748;
wire v_3751;
wire v_3752;
wire v_3753;
wire v_3754;
wire v_3755;
wire v_3756;
wire v_3757;
wire v_3758;
wire v_3759;
wire v_3760;
wire v_3763;
wire v_3764;
wire v_3765;
wire v_3766;
wire v_3767;
wire v_3768;
wire v_3769;
wire v_3770;
wire v_3771;
wire v_3772;
wire v_3775;
wire v_3776;
wire v_3777;
wire v_3778;
wire v_3779;
wire v_3780;
wire v_3781;
wire v_3782;
wire v_3783;
wire v_3784;
wire v_3785;
wire v_3786;
wire v_3787;
wire v_3788;
wire v_3789;
wire v_3790;
wire v_3791;
wire v_3792;
wire v_3793;
wire v_3794;
wire v_3795;
wire v_3796;
wire v_3797;
wire v_3798;
wire v_3799;
wire v_3800;
wire v_3803;
wire v_3804;
wire v_3805;
wire v_3806;
wire v_3807;
wire v_3808;
wire v_3809;
wire v_3810;
wire v_3811;
wire v_3812;
wire v_3814;
wire v_3815;
wire v_3816;
wire v_3817;
wire v_3818;
wire v_3819;
wire v_3820;
wire v_3822;
wire v_3823;
wire v_3824;
wire v_3825;
wire v_3826;
wire v_3827;
wire v_3828;
wire v_3829;
wire v_3830;
wire v_3831;
wire v_3832;
wire v_3833;
wire v_3834;
wire v_3835;
wire v_3836;
wire v_3837;
wire v_3838;
wire v_3839;
wire v_3840;
wire v_3841;
wire v_3842;
wire v_3843;
wire v_3844;
wire v_3845;
wire v_3846;
wire v_3847;
wire v_3848;
wire v_3849;
wire v_3850;
wire v_3851;
wire v_3852;
wire v_3853;
wire v_3854;
wire v_3855;
wire v_3856;
wire v_3857;
wire v_3858;
wire v_3859;
wire v_3860;
wire v_3861;
wire v_3862;
wire v_3863;
wire v_3864;
wire v_3867;
wire v_3868;
wire v_3869;
wire v_3870;
wire v_3871;
wire v_3872;
wire v_3873;
wire v_3874;
wire v_3875;
wire v_3876;
wire v_3879;
wire v_3880;
wire v_3881;
wire v_3882;
wire v_3883;
wire v_3884;
wire v_3885;
wire v_3886;
wire v_3887;
wire v_3888;
wire v_3891;
wire v_3892;
wire v_3893;
wire v_3894;
wire v_3895;
wire v_3896;
wire v_3897;
wire v_3898;
wire v_3899;
wire v_3900;
wire v_3903;
wire v_3904;
wire v_3905;
wire v_3906;
wire v_3907;
wire v_3908;
wire v_3909;
wire v_3910;
wire v_3911;
wire v_3912;
wire v_3915;
wire v_3916;
wire v_3917;
wire v_3918;
wire v_3919;
wire v_3920;
wire v_3921;
wire v_3922;
wire v_3923;
wire v_3924;
wire v_3927;
wire v_3928;
wire v_3929;
wire v_3930;
wire v_3931;
wire v_3932;
wire v_3933;
wire v_3934;
wire v_3935;
wire v_3936;
wire v_3937;
wire v_3938;
wire v_3939;
wire v_3940;
wire v_3941;
wire v_3942;
wire v_3943;
wire v_3944;
wire v_3945;
wire v_3946;
wire v_3947;
wire v_3948;
wire v_3949;
wire v_3950;
wire v_3951;
wire v_3952;
wire v_3955;
wire v_3956;
wire v_3957;
wire v_3958;
wire v_3959;
wire v_3960;
wire v_3961;
wire v_3962;
wire v_3963;
wire v_3964;
wire v_3966;
wire v_3968;
wire v_3969;
wire v_3970;
wire v_3971;
wire v_3972;
wire v_3973;
wire v_3974;
wire v_3975;
wire v_3976;
wire v_3977;
wire v_3978;
wire v_3979;
wire v_3980;
wire v_3981;
wire v_3982;
wire v_3983;
wire v_3984;
wire v_3985;
wire v_3986;
wire v_3987;
wire v_3988;
wire v_3989;
wire v_3990;
wire v_3991;
wire v_3992;
wire v_3993;
wire v_3994;
wire v_3995;
wire v_3996;
wire v_3999;
wire v_4000;
wire v_4001;
wire v_4002;
wire v_4003;
wire v_4004;
wire v_4005;
wire v_4006;
wire v_4007;
wire v_4008;
wire v_4011;
wire v_4012;
wire v_4013;
wire v_4014;
wire v_4015;
wire v_4016;
wire v_4017;
wire v_4018;
wire v_4019;
wire v_4020;
wire v_4023;
wire v_4024;
wire v_4025;
wire v_4026;
wire v_4027;
wire v_4028;
wire v_4029;
wire v_4030;
wire v_4031;
wire v_4032;
wire v_4035;
wire v_4036;
wire v_4037;
wire v_4038;
wire v_4039;
wire v_4040;
wire v_4041;
wire v_4042;
wire v_4043;
wire v_4044;
wire v_4047;
wire v_4048;
wire v_4049;
wire v_4050;
wire v_4051;
wire v_4052;
wire v_4053;
wire v_4054;
wire v_4055;
wire v_4056;
wire v_4059;
wire v_4060;
wire v_4061;
wire v_4062;
wire v_4063;
wire v_4064;
wire v_4065;
wire v_4066;
wire v_4067;
wire v_4068;
wire v_4069;
wire v_4070;
wire v_4071;
wire v_4072;
wire v_4073;
wire v_4074;
wire v_4075;
wire v_4076;
wire v_4077;
wire v_4078;
wire v_4079;
wire v_4080;
wire v_4081;
wire v_4082;
wire v_4083;
wire v_4084;
wire v_4087;
wire v_4088;
wire v_4089;
wire v_4090;
wire v_4091;
wire v_4092;
wire v_4093;
wire v_4094;
wire v_4095;
wire v_4096;
wire v_4098;
wire v_4099;
wire v_4100;
wire v_4101;
wire v_4102;
wire v_4104;
wire v_4105;
wire v_4106;
wire v_4107;
wire v_4108;
wire v_4109;
wire v_4110;
wire v_4111;
wire v_4112;
wire v_4113;
wire v_4114;
wire v_4115;
wire v_4116;
wire v_4117;
wire v_4118;
wire v_4119;
wire v_4120;
wire v_4121;
wire v_4122;
wire v_4123;
wire v_4124;
wire v_4125;
wire v_4126;
wire v_4127;
wire v_4128;
wire v_4129;
wire v_4130;
wire v_4131;
wire v_4132;
wire v_4133;
wire v_4134;
wire v_4135;
wire v_4136;
wire v_4137;
wire v_4138;
wire v_4139;
wire v_4140;
wire v_4141;
wire v_4142;
wire v_4143;
wire v_4144;
wire v_4145;
wire v_4146;
wire v_4147;
wire v_4148;
wire v_4149;
wire v_4150;
wire v_4151;
wire v_4152;
wire v_4153;
wire v_4154;
wire v_4155;
wire v_4156;
wire v_4157;
wire v_4158;
wire v_4159;
wire v_4160;
wire v_4163;
wire v_4164;
wire v_4165;
wire v_4166;
wire v_4167;
wire v_4168;
wire v_4169;
wire v_4170;
wire v_4171;
wire v_4172;
wire v_4175;
wire v_4176;
wire v_4177;
wire v_4178;
wire v_4179;
wire v_4180;
wire v_4181;
wire v_4182;
wire v_4183;
wire v_4184;
wire v_4187;
wire v_4188;
wire v_4189;
wire v_4190;
wire v_4191;
wire v_4192;
wire v_4193;
wire v_4194;
wire v_4195;
wire v_4196;
wire v_4199;
wire v_4200;
wire v_4201;
wire v_4202;
wire v_4203;
wire v_4204;
wire v_4205;
wire v_4206;
wire v_4207;
wire v_4208;
wire v_4211;
wire v_4212;
wire v_4213;
wire v_4214;
wire v_4215;
wire v_4216;
wire v_4217;
wire v_4218;
wire v_4219;
wire v_4220;
wire v_4223;
wire v_4224;
wire v_4225;
wire v_4226;
wire v_4227;
wire v_4228;
wire v_4229;
wire v_4230;
wire v_4231;
wire v_4232;
wire v_4233;
wire v_4234;
wire v_4235;
wire v_4236;
wire v_4237;
wire v_4238;
wire v_4239;
wire v_4240;
wire v_4241;
wire v_4242;
wire v_4243;
wire v_4244;
wire v_4245;
wire v_4246;
wire v_4247;
wire v_4248;
wire v_4251;
wire v_4252;
wire v_4253;
wire v_4254;
wire v_4255;
wire v_4256;
wire v_4257;
wire v_4258;
wire v_4259;
wire v_4260;
wire v_4262;
wire v_4264;
wire v_4265;
wire v_4266;
wire v_4267;
wire v_4268;
wire v_4269;
wire v_4270;
wire v_4271;
wire v_4272;
wire v_4273;
wire v_4274;
wire v_4275;
wire v_4276;
wire v_4277;
wire v_4278;
wire v_4279;
wire v_4280;
wire v_4281;
wire v_4282;
wire v_4283;
wire v_4284;
wire v_4285;
wire v_4286;
wire v_4287;
wire v_4288;
wire v_4289;
wire v_4290;
wire v_4291;
wire v_4292;
wire v_4295;
wire v_4296;
wire v_4297;
wire v_4298;
wire v_4299;
wire v_4300;
wire v_4301;
wire v_4302;
wire v_4303;
wire v_4304;
wire v_4307;
wire v_4308;
wire v_4309;
wire v_4310;
wire v_4311;
wire v_4312;
wire v_4313;
wire v_4314;
wire v_4315;
wire v_4316;
wire v_4319;
wire v_4320;
wire v_4321;
wire v_4322;
wire v_4323;
wire v_4324;
wire v_4325;
wire v_4326;
wire v_4327;
wire v_4328;
wire v_4331;
wire v_4332;
wire v_4333;
wire v_4334;
wire v_4335;
wire v_4336;
wire v_4337;
wire v_4338;
wire v_4339;
wire v_4340;
wire v_4343;
wire v_4344;
wire v_4345;
wire v_4346;
wire v_4347;
wire v_4348;
wire v_4349;
wire v_4350;
wire v_4351;
wire v_4352;
wire v_4355;
wire v_4356;
wire v_4357;
wire v_4358;
wire v_4359;
wire v_4360;
wire v_4361;
wire v_4362;
wire v_4363;
wire v_4364;
wire v_4365;
wire v_4366;
wire v_4367;
wire v_4368;
wire v_4369;
wire v_4370;
wire v_4371;
wire v_4372;
wire v_4373;
wire v_4374;
wire v_4375;
wire v_4376;
wire v_4377;
wire v_4378;
wire v_4379;
wire v_4380;
wire v_4383;
wire v_4384;
wire v_4385;
wire v_4386;
wire v_4387;
wire v_4388;
wire v_4389;
wire v_4390;
wire v_4391;
wire v_4392;
wire v_4394;
wire v_4395;
wire v_4396;
wire v_4397;
wire v_4398;
wire v_4399;
wire v_4401;
wire v_4402;
wire v_4403;
wire v_4404;
wire v_4405;
wire v_4406;
wire v_4407;
wire v_4408;
wire v_4409;
wire v_4410;
wire v_4411;
wire v_4412;
wire v_4413;
wire v_4414;
wire v_4415;
wire v_4416;
wire v_4417;
wire v_4418;
wire v_4419;
wire v_4420;
wire v_4421;
wire v_4422;
wire v_4423;
wire v_4424;
wire v_4425;
wire v_4426;
wire v_4427;
wire v_4428;
wire v_4429;
wire v_4430;
wire v_4431;
wire v_4432;
wire v_4433;
wire v_4434;
wire v_4435;
wire v_4436;
wire v_4437;
wire v_4438;
wire v_4439;
wire v_4440;
wire v_4441;
wire v_4442;
wire v_4445;
wire v_4446;
wire v_4447;
wire v_4448;
wire v_4449;
wire v_4450;
wire v_4451;
wire v_4452;
wire v_4453;
wire v_4454;
wire v_4457;
wire v_4458;
wire v_4459;
wire v_4460;
wire v_4461;
wire v_4462;
wire v_4463;
wire v_4464;
wire v_4465;
wire v_4466;
wire v_4469;
wire v_4470;
wire v_4471;
wire v_4472;
wire v_4473;
wire v_4474;
wire v_4475;
wire v_4476;
wire v_4477;
wire v_4478;
wire v_4481;
wire v_4482;
wire v_4483;
wire v_4484;
wire v_4485;
wire v_4486;
wire v_4487;
wire v_4488;
wire v_4489;
wire v_4490;
wire v_4493;
wire v_4494;
wire v_4495;
wire v_4496;
wire v_4497;
wire v_4498;
wire v_4499;
wire v_4500;
wire v_4501;
wire v_4502;
wire v_4505;
wire v_4506;
wire v_4507;
wire v_4508;
wire v_4509;
wire v_4510;
wire v_4511;
wire v_4512;
wire v_4513;
wire v_4514;
wire v_4515;
wire v_4516;
wire v_4517;
wire v_4518;
wire v_4519;
wire v_4520;
wire v_4521;
wire v_4522;
wire v_4523;
wire v_4524;
wire v_4525;
wire v_4526;
wire v_4527;
wire v_4528;
wire v_4529;
wire v_4530;
wire v_4533;
wire v_4534;
wire v_4535;
wire v_4536;
wire v_4537;
wire v_4538;
wire v_4539;
wire v_4540;
wire v_4541;
wire v_4542;
wire v_4544;
wire v_4546;
wire v_4547;
wire v_4548;
wire v_4549;
wire v_4550;
wire v_4551;
wire v_4552;
wire v_4553;
wire v_4554;
wire v_4555;
wire v_4556;
wire v_4557;
wire v_4558;
wire v_4559;
wire v_4560;
wire v_4561;
wire v_4562;
wire v_4563;
wire v_4564;
wire v_4565;
wire v_4566;
wire v_4567;
wire v_4568;
wire v_4569;
wire v_4570;
wire v_4571;
wire v_4572;
wire v_4573;
wire v_4574;
wire v_4577;
wire v_4578;
wire v_4579;
wire v_4580;
wire v_4581;
wire v_4582;
wire v_4583;
wire v_4584;
wire v_4585;
wire v_4586;
wire v_4589;
wire v_4590;
wire v_4591;
wire v_4592;
wire v_4593;
wire v_4594;
wire v_4595;
wire v_4596;
wire v_4597;
wire v_4598;
wire v_4601;
wire v_4602;
wire v_4603;
wire v_4604;
wire v_4605;
wire v_4606;
wire v_4607;
wire v_4608;
wire v_4609;
wire v_4610;
wire v_4613;
wire v_4614;
wire v_4615;
wire v_4616;
wire v_4617;
wire v_4618;
wire v_4619;
wire v_4620;
wire v_4621;
wire v_4622;
wire v_4625;
wire v_4626;
wire v_4627;
wire v_4628;
wire v_4629;
wire v_4630;
wire v_4631;
wire v_4632;
wire v_4633;
wire v_4634;
wire v_4637;
wire v_4638;
wire v_4639;
wire v_4640;
wire v_4641;
wire v_4642;
wire v_4643;
wire v_4644;
wire v_4645;
wire v_4646;
wire v_4647;
wire v_4648;
wire v_4649;
wire v_4650;
wire v_4651;
wire v_4652;
wire v_4653;
wire v_4654;
wire v_4655;
wire v_4656;
wire v_4657;
wire v_4658;
wire v_4659;
wire v_4660;
wire v_4661;
wire v_4662;
wire v_4665;
wire v_4666;
wire v_4667;
wire v_4668;
wire v_4669;
wire v_4670;
wire v_4671;
wire v_4672;
wire v_4673;
wire v_4674;
wire v_4676;
wire v_4677;
wire v_4678;
wire v_4679;
wire v_4680;
wire v_4682;
wire v_4683;
wire v_4684;
wire v_4685;
wire v_4686;
wire v_4687;
wire v_4688;
wire v_4689;
wire v_4690;
wire v_4691;
wire v_4692;
wire v_4693;
wire v_4694;
wire v_4695;
wire v_4696;
wire v_4697;
wire v_4698;
wire v_4699;
wire v_4700;
wire v_4701;
wire v_4702;
wire v_4703;
wire v_4704;
wire v_4705;
wire v_4706;
wire v_4707;
wire v_4708;
wire v_4709;
wire v_4710;
wire v_4711;
wire v_4712;
wire v_4713;
wire v_4714;
wire v_4715;
wire v_4716;
wire v_4717;
wire v_4718;
wire v_4719;
wire v_4720;
wire v_4721;
wire v_4722;
wire v_4723;
wire v_4724;
wire v_4725;
wire v_4726;
wire v_4727;
wire v_4728;
wire v_4729;
wire v_4730;
wire v_4733;
wire v_4734;
wire v_4735;
wire v_4736;
wire v_4737;
wire v_4738;
wire v_4739;
wire v_4740;
wire v_4741;
wire v_4742;
wire v_4745;
wire v_4746;
wire v_4747;
wire v_4748;
wire v_4749;
wire v_4750;
wire v_4751;
wire v_4752;
wire v_4753;
wire v_4754;
wire v_4757;
wire v_4758;
wire v_4759;
wire v_4760;
wire v_4761;
wire v_4762;
wire v_4763;
wire v_4764;
wire v_4765;
wire v_4766;
wire v_4769;
wire v_4770;
wire v_4771;
wire v_4772;
wire v_4773;
wire v_4774;
wire v_4775;
wire v_4776;
wire v_4777;
wire v_4778;
wire v_4781;
wire v_4782;
wire v_4783;
wire v_4784;
wire v_4785;
wire v_4786;
wire v_4787;
wire v_4788;
wire v_4789;
wire v_4790;
wire v_4793;
wire v_4794;
wire v_4795;
wire v_4796;
wire v_4797;
wire v_4798;
wire v_4799;
wire v_4800;
wire v_4801;
wire v_4802;
wire v_4803;
wire v_4804;
wire v_4805;
wire v_4806;
wire v_4807;
wire v_4808;
wire v_4809;
wire v_4810;
wire v_4811;
wire v_4812;
wire v_4813;
wire v_4814;
wire v_4815;
wire v_4816;
wire v_4817;
wire v_4818;
wire v_4821;
wire v_4822;
wire v_4823;
wire v_4824;
wire v_4825;
wire v_4826;
wire v_4827;
wire v_4828;
wire v_4829;
wire v_4830;
wire v_4832;
wire v_4834;
wire v_4835;
wire v_4836;
wire v_4837;
wire v_4838;
wire v_4839;
wire v_4840;
wire v_4841;
wire v_4842;
wire v_4843;
wire v_4844;
wire v_4845;
wire v_4846;
wire v_4847;
wire v_4848;
wire v_4849;
wire v_4850;
wire v_4851;
wire v_4852;
wire v_4853;
wire v_4854;
wire v_4855;
wire v_4856;
wire v_4857;
wire v_4858;
wire v_4859;
wire v_4860;
wire v_4861;
wire v_4862;
wire v_4865;
wire v_4866;
wire v_4867;
wire v_4868;
wire v_4869;
wire v_4870;
wire v_4871;
wire v_4872;
wire v_4873;
wire v_4874;
wire v_4877;
wire v_4878;
wire v_4879;
wire v_4880;
wire v_4881;
wire v_4882;
wire v_4883;
wire v_4884;
wire v_4885;
wire v_4886;
wire v_4889;
wire v_4890;
wire v_4891;
wire v_4892;
wire v_4893;
wire v_4894;
wire v_4895;
wire v_4896;
wire v_4897;
wire v_4898;
wire v_4901;
wire v_4902;
wire v_4903;
wire v_4904;
wire v_4905;
wire v_4906;
wire v_4907;
wire v_4908;
wire v_4909;
wire v_4910;
wire v_4913;
wire v_4914;
wire v_4915;
wire v_4916;
wire v_4917;
wire v_4918;
wire v_4919;
wire v_4920;
wire v_4921;
wire v_4922;
wire v_4925;
wire v_4926;
wire v_4927;
wire v_4928;
wire v_4929;
wire v_4930;
wire v_4931;
wire v_4932;
wire v_4933;
wire v_4934;
wire v_4935;
wire v_4936;
wire v_4937;
wire v_4938;
wire v_4939;
wire v_4940;
wire v_4941;
wire v_4942;
wire v_4943;
wire v_4944;
wire v_4945;
wire v_4946;
wire v_4947;
wire v_4948;
wire v_4949;
wire v_4950;
wire v_4953;
wire v_4954;
wire v_4955;
wire v_4956;
wire v_4957;
wire v_4958;
wire v_4959;
wire v_4960;
wire v_4961;
wire v_4962;
wire v_4964;
wire v_4965;
wire v_4966;
wire v_4967;
wire v_4968;
wire v_4969;
wire v_4970;
wire v_4971;
wire v_4972;
wire v_4974;
wire v_4975;
wire v_4976;
wire v_4977;
wire v_4978;
wire v_4979;
wire v_4980;
wire v_4981;
wire v_4982;
wire v_4983;
wire v_4984;
wire v_4985;
wire v_4986;
wire v_4987;
wire v_4988;
wire v_4989;
wire v_4990;
wire v_4991;
wire v_4992;
wire v_4993;
wire v_4994;
wire v_4995;
wire v_4996;
wire v_4997;
wire v_4998;
wire v_4999;
wire v_5000;
wire v_5001;
wire v_5002;
wire v_5003;
wire v_5004;
wire v_5005;
wire v_5006;
wire v_5007;
wire v_5008;
wire v_5009;
wire v_5010;
wire v_5011;
wire v_5012;
wire v_5013;
wire v_5014;
wire v_5015;
wire v_5016;
wire v_5017;
wire v_5018;
wire v_5021;
wire v_5022;
wire v_5023;
wire v_5024;
wire v_5025;
wire v_5026;
wire v_5027;
wire v_5028;
wire v_5029;
wire v_5030;
wire v_5033;
wire v_5034;
wire v_5035;
wire v_5036;
wire v_5037;
wire v_5038;
wire v_5039;
wire v_5040;
wire v_5041;
wire v_5042;
wire v_5045;
wire v_5046;
wire v_5047;
wire v_5048;
wire v_5049;
wire v_5050;
wire v_5051;
wire v_5052;
wire v_5053;
wire v_5054;
wire v_5057;
wire v_5058;
wire v_5059;
wire v_5060;
wire v_5061;
wire v_5062;
wire v_5063;
wire v_5064;
wire v_5065;
wire v_5066;
wire v_5069;
wire v_5070;
wire v_5071;
wire v_5072;
wire v_5073;
wire v_5074;
wire v_5075;
wire v_5076;
wire v_5077;
wire v_5078;
wire v_5081;
wire v_5082;
wire v_5083;
wire v_5084;
wire v_5085;
wire v_5086;
wire v_5087;
wire v_5088;
wire v_5089;
wire v_5090;
wire v_5091;
wire v_5092;
wire v_5093;
wire v_5094;
wire v_5095;
wire v_5096;
wire v_5097;
wire v_5098;
wire v_5099;
wire v_5100;
wire v_5101;
wire v_5102;
wire v_5103;
wire v_5104;
wire v_5105;
wire v_5106;
wire v_5109;
wire v_5110;
wire v_5111;
wire v_5112;
wire v_5113;
wire v_5114;
wire v_5115;
wire v_5116;
wire v_5117;
wire v_5118;
wire v_5120;
wire v_5122;
wire v_5123;
wire v_5124;
wire v_5125;
wire v_5126;
wire v_5127;
wire v_5128;
wire v_5129;
wire v_5130;
wire v_5131;
wire v_5132;
wire v_5133;
wire v_5134;
wire v_5135;
wire v_5136;
wire v_5137;
wire v_5138;
wire v_5139;
wire v_5140;
wire v_5141;
wire v_5142;
wire v_5143;
wire v_5144;
wire v_5145;
wire v_5146;
wire v_5147;
wire v_5148;
wire v_5149;
wire v_5150;
wire v_5153;
wire v_5154;
wire v_5155;
wire v_5156;
wire v_5157;
wire v_5158;
wire v_5159;
wire v_5160;
wire v_5161;
wire v_5162;
wire v_5165;
wire v_5166;
wire v_5167;
wire v_5168;
wire v_5169;
wire v_5170;
wire v_5171;
wire v_5172;
wire v_5173;
wire v_5174;
wire v_5177;
wire v_5178;
wire v_5179;
wire v_5180;
wire v_5181;
wire v_5182;
wire v_5183;
wire v_5184;
wire v_5185;
wire v_5186;
wire v_5189;
wire v_5190;
wire v_5191;
wire v_5192;
wire v_5193;
wire v_5194;
wire v_5195;
wire v_5196;
wire v_5197;
wire v_5198;
wire v_5201;
wire v_5202;
wire v_5203;
wire v_5204;
wire v_5205;
wire v_5206;
wire v_5207;
wire v_5208;
wire v_5209;
wire v_5210;
wire v_5213;
wire v_5214;
wire v_5215;
wire v_5216;
wire v_5217;
wire v_5218;
wire v_5219;
wire v_5220;
wire v_5221;
wire v_5222;
wire v_5223;
wire v_5224;
wire v_5225;
wire v_5226;
wire v_5227;
wire v_5228;
wire v_5229;
wire v_5230;
wire v_5231;
wire v_5232;
wire v_5233;
wire v_5234;
wire v_5235;
wire v_5236;
wire v_5237;
wire v_5238;
wire v_5241;
wire v_5242;
wire v_5243;
wire v_5244;
wire v_5245;
wire v_5246;
wire v_5247;
wire v_5248;
wire v_5249;
wire v_5250;
wire v_5252;
wire v_5253;
wire v_5254;
wire v_5255;
wire v_5256;
wire v_5258;
wire v_5259;
wire v_5260;
wire v_5261;
wire v_5262;
wire v_5263;
wire v_5264;
wire v_5265;
wire v_5266;
wire v_5267;
wire v_5268;
wire v_5269;
wire v_5270;
wire v_5271;
wire v_5272;
wire v_5273;
wire v_5274;
wire v_5275;
wire v_5276;
wire v_5277;
wire v_5278;
wire v_5279;
wire v_5280;
wire v_5281;
wire v_5282;
wire v_5283;
wire v_5284;
wire v_5285;
wire v_5286;
wire v_5287;
wire v_5288;
wire v_5289;
wire v_5290;
wire v_5291;
wire v_5292;
wire v_5293;
wire v_5294;
wire v_5295;
wire v_5296;
wire v_5297;
wire v_5298;
wire v_5299;
wire v_5300;
wire v_5301;
wire v_5302;
wire v_5303;
wire v_5304;
wire v_5305;
wire v_5306;
wire v_5307;
wire v_5308;
wire v_5309;
wire v_5310;
wire v_5311;
wire v_5312;
wire v_5313;
wire v_5314;
wire v_5315;
wire v_5316;
wire v_5317;
wire v_5318;
wire v_5319;
wire v_5320;
wire v_5321;
wire v_5322;
wire v_5323;
wire v_5324;
wire v_5325;
wire v_5326;
wire v_5327;
wire v_5328;
wire v_5329;
wire v_5330;
wire v_5333;
wire v_5334;
wire v_5335;
wire v_5336;
wire v_5337;
wire v_5338;
wire v_5339;
wire v_5340;
wire v_5341;
wire v_5342;
wire v_5345;
wire v_5346;
wire v_5347;
wire v_5348;
wire v_5349;
wire v_5350;
wire v_5351;
wire v_5352;
wire v_5353;
wire v_5354;
wire v_5357;
wire v_5358;
wire v_5359;
wire v_5360;
wire v_5361;
wire v_5362;
wire v_5363;
wire v_5364;
wire v_5365;
wire v_5366;
wire v_5369;
wire v_5370;
wire v_5371;
wire v_5372;
wire v_5373;
wire v_5374;
wire v_5375;
wire v_5376;
wire v_5377;
wire v_5378;
wire v_5381;
wire v_5382;
wire v_5383;
wire v_5384;
wire v_5385;
wire v_5386;
wire v_5387;
wire v_5388;
wire v_5389;
wire v_5390;
wire v_5393;
wire v_5394;
wire v_5395;
wire v_5396;
wire v_5397;
wire v_5398;
wire v_5399;
wire v_5400;
wire v_5401;
wire v_5402;
wire v_5403;
wire v_5404;
wire v_5405;
wire v_5406;
wire v_5407;
wire v_5408;
wire v_5409;
wire v_5410;
wire v_5411;
wire v_5412;
wire v_5413;
wire v_5414;
wire v_5415;
wire v_5416;
wire v_5417;
wire v_5418;
wire v_5421;
wire v_5422;
wire v_5423;
wire v_5424;
wire v_5425;
wire v_5426;
wire v_5427;
wire v_5428;
wire v_5429;
wire v_5430;
wire v_5432;
wire v_5434;
wire v_5435;
wire v_5436;
wire v_5437;
wire v_5438;
wire v_5439;
wire v_5440;
wire v_5441;
wire v_5442;
wire v_5443;
wire v_5444;
wire v_5445;
wire v_5446;
wire v_5447;
wire v_5448;
wire v_5449;
wire v_5450;
wire v_5451;
wire v_5452;
wire v_5453;
wire v_5454;
wire v_5455;
wire v_5456;
wire v_5457;
wire v_5458;
wire v_5459;
wire v_5460;
wire v_5461;
wire v_5462;
wire v_5465;
wire v_5466;
wire v_5467;
wire v_5468;
wire v_5469;
wire v_5470;
wire v_5471;
wire v_5472;
wire v_5473;
wire v_5474;
wire v_5477;
wire v_5478;
wire v_5479;
wire v_5480;
wire v_5481;
wire v_5482;
wire v_5483;
wire v_5484;
wire v_5485;
wire v_5486;
wire v_5489;
wire v_5490;
wire v_5491;
wire v_5492;
wire v_5493;
wire v_5494;
wire v_5495;
wire v_5496;
wire v_5497;
wire v_5498;
wire v_5501;
wire v_5502;
wire v_5503;
wire v_5504;
wire v_5505;
wire v_5506;
wire v_5507;
wire v_5508;
wire v_5509;
wire v_5510;
wire v_5513;
wire v_5514;
wire v_5515;
wire v_5516;
wire v_5517;
wire v_5518;
wire v_5519;
wire v_5520;
wire v_5521;
wire v_5522;
wire v_5525;
wire v_5526;
wire v_5527;
wire v_5528;
wire v_5529;
wire v_5530;
wire v_5531;
wire v_5532;
wire v_5533;
wire v_5534;
wire v_5535;
wire v_5536;
wire v_5537;
wire v_5538;
wire v_5539;
wire v_5540;
wire v_5541;
wire v_5542;
wire v_5543;
wire v_5544;
wire v_5545;
wire v_5546;
wire v_5547;
wire v_5548;
wire v_5549;
wire v_5550;
wire v_5553;
wire v_5554;
wire v_5555;
wire v_5556;
wire v_5557;
wire v_5558;
wire v_5559;
wire v_5560;
wire v_5561;
wire v_5562;
wire v_5564;
wire v_5565;
wire v_5566;
wire v_5567;
wire v_5568;
wire v_5569;
wire v_5571;
wire v_5572;
wire v_5573;
wire v_5574;
wire v_5575;
wire v_5576;
wire v_5577;
wire v_5578;
wire v_5579;
wire v_5580;
wire v_5581;
wire v_5582;
wire v_5583;
wire v_5584;
wire v_5585;
wire v_5586;
wire v_5587;
wire v_5588;
wire v_5589;
wire v_5590;
wire v_5591;
wire v_5592;
wire v_5593;
wire v_5594;
wire v_5595;
wire v_5596;
wire v_5597;
wire v_5598;
wire v_5599;
wire v_5600;
wire v_5601;
wire v_5602;
wire v_5603;
wire v_5604;
wire v_5605;
wire v_5606;
wire v_5607;
wire v_5608;
wire v_5609;
wire v_5610;
wire v_5611;
wire v_5612;
wire v_5615;
wire v_5616;
wire v_5617;
wire v_5618;
wire v_5619;
wire v_5620;
wire v_5621;
wire v_5622;
wire v_5623;
wire v_5624;
wire v_5627;
wire v_5628;
wire v_5629;
wire v_5630;
wire v_5631;
wire v_5632;
wire v_5633;
wire v_5634;
wire v_5635;
wire v_5636;
wire v_5639;
wire v_5640;
wire v_5641;
wire v_5642;
wire v_5643;
wire v_5644;
wire v_5645;
wire v_5646;
wire v_5647;
wire v_5648;
wire v_5651;
wire v_5652;
wire v_5653;
wire v_5654;
wire v_5655;
wire v_5656;
wire v_5657;
wire v_5658;
wire v_5659;
wire v_5660;
wire v_5663;
wire v_5664;
wire v_5665;
wire v_5666;
wire v_5667;
wire v_5668;
wire v_5669;
wire v_5670;
wire v_5671;
wire v_5672;
wire v_5675;
wire v_5676;
wire v_5677;
wire v_5678;
wire v_5679;
wire v_5680;
wire v_5681;
wire v_5682;
wire v_5683;
wire v_5684;
wire v_5685;
wire v_5686;
wire v_5687;
wire v_5688;
wire v_5689;
wire v_5690;
wire v_5691;
wire v_5692;
wire v_5693;
wire v_5694;
wire v_5695;
wire v_5696;
wire v_5697;
wire v_5698;
wire v_5699;
wire v_5700;
wire v_5703;
wire v_5704;
wire v_5705;
wire v_5706;
wire v_5707;
wire v_5708;
wire v_5709;
wire v_5710;
wire v_5711;
wire v_5712;
wire v_5714;
wire v_5716;
wire v_5717;
wire v_5718;
wire v_5719;
wire v_5720;
wire v_5721;
wire v_5722;
wire v_5723;
wire v_5724;
wire v_5725;
wire v_5726;
wire v_5727;
wire v_5728;
wire v_5729;
wire v_5730;
wire v_5731;
wire v_5732;
wire v_5733;
wire v_5734;
wire v_5735;
wire v_5736;
wire v_5737;
wire v_5738;
wire v_5739;
wire v_5740;
wire v_5741;
wire v_5742;
wire v_5743;
wire v_5744;
wire v_5747;
wire v_5748;
wire v_5749;
wire v_5750;
wire v_5751;
wire v_5752;
wire v_5753;
wire v_5754;
wire v_5755;
wire v_5756;
wire v_5759;
wire v_5760;
wire v_5761;
wire v_5762;
wire v_5763;
wire v_5764;
wire v_5765;
wire v_5766;
wire v_5767;
wire v_5768;
wire v_5771;
wire v_5772;
wire v_5773;
wire v_5774;
wire v_5775;
wire v_5776;
wire v_5777;
wire v_5778;
wire v_5779;
wire v_5780;
wire v_5783;
wire v_5784;
wire v_5785;
wire v_5786;
wire v_5787;
wire v_5788;
wire v_5789;
wire v_5790;
wire v_5791;
wire v_5792;
wire v_5795;
wire v_5796;
wire v_5797;
wire v_5798;
wire v_5799;
wire v_5800;
wire v_5801;
wire v_5802;
wire v_5803;
wire v_5804;
wire v_5807;
wire v_5808;
wire v_5809;
wire v_5810;
wire v_5811;
wire v_5812;
wire v_5813;
wire v_5814;
wire v_5815;
wire v_5816;
wire v_5817;
wire v_5818;
wire v_5819;
wire v_5820;
wire v_5821;
wire v_5822;
wire v_5823;
wire v_5824;
wire v_5825;
wire v_5826;
wire v_5827;
wire v_5828;
wire v_5829;
wire v_5830;
wire v_5831;
wire v_5832;
wire v_5835;
wire v_5836;
wire v_5837;
wire v_5838;
wire v_5839;
wire v_5840;
wire v_5841;
wire v_5842;
wire v_5843;
wire v_5844;
wire v_5846;
wire v_5847;
wire v_5848;
wire v_5849;
wire v_5850;
wire v_5852;
wire v_5853;
wire v_5854;
wire v_5855;
wire v_5856;
wire v_5857;
wire v_5858;
wire v_5859;
wire v_5860;
wire v_5861;
wire v_5862;
wire v_5863;
wire v_5864;
wire v_5865;
wire v_5866;
wire v_5867;
wire v_5868;
wire v_5869;
wire v_5870;
wire v_5871;
wire v_5872;
wire v_5873;
wire v_5874;
wire v_5875;
wire v_5876;
wire v_5877;
wire v_5878;
wire v_5879;
wire v_5880;
wire v_5881;
wire v_5882;
wire v_5883;
wire v_5884;
wire v_5885;
wire v_5886;
wire v_5887;
wire v_5888;
wire v_5889;
wire v_5890;
wire v_5891;
wire v_5892;
wire v_5893;
wire v_5894;
wire v_5895;
wire v_5896;
wire v_5897;
wire v_5898;
wire v_5899;
wire v_5900;
wire v_5903;
wire v_5904;
wire v_5905;
wire v_5906;
wire v_5907;
wire v_5908;
wire v_5909;
wire v_5910;
wire v_5911;
wire v_5912;
wire v_5915;
wire v_5916;
wire v_5917;
wire v_5918;
wire v_5919;
wire v_5920;
wire v_5921;
wire v_5922;
wire v_5923;
wire v_5924;
wire v_5927;
wire v_5928;
wire v_5929;
wire v_5930;
wire v_5931;
wire v_5932;
wire v_5933;
wire v_5934;
wire v_5935;
wire v_5936;
wire v_5939;
wire v_5940;
wire v_5941;
wire v_5942;
wire v_5943;
wire v_5944;
wire v_5945;
wire v_5946;
wire v_5947;
wire v_5948;
wire v_5951;
wire v_5952;
wire v_5953;
wire v_5954;
wire v_5955;
wire v_5956;
wire v_5957;
wire v_5958;
wire v_5959;
wire v_5960;
wire v_5963;
wire v_5964;
wire v_5965;
wire v_5966;
wire v_5967;
wire v_5968;
wire v_5969;
wire v_5970;
wire v_5971;
wire v_5972;
wire v_5973;
wire v_5974;
wire v_5975;
wire v_5976;
wire v_5977;
wire v_5978;
wire v_5979;
wire v_5980;
wire v_5981;
wire v_5982;
wire v_5983;
wire v_5984;
wire v_5985;
wire v_5986;
wire v_5987;
wire v_5988;
wire v_5991;
wire v_5992;
wire v_5993;
wire v_5994;
wire v_5995;
wire v_5996;
wire v_5997;
wire v_5998;
wire v_5999;
wire v_6000;
wire v_6002;
wire v_6004;
wire v_6005;
wire v_6006;
wire v_6007;
wire v_6008;
wire v_6009;
wire v_6010;
wire v_6011;
wire v_6012;
wire v_6013;
wire v_6014;
wire v_6015;
wire v_6016;
wire v_6017;
wire v_6018;
wire v_6019;
wire v_6020;
wire v_6021;
wire v_6022;
wire v_6023;
wire v_6024;
wire v_6025;
wire v_6026;
wire v_6027;
wire v_6028;
wire v_6029;
wire v_6030;
wire v_6031;
wire v_6032;
wire v_6035;
wire v_6036;
wire v_6037;
wire v_6038;
wire v_6039;
wire v_6040;
wire v_6041;
wire v_6042;
wire v_6043;
wire v_6044;
wire v_6047;
wire v_6048;
wire v_6049;
wire v_6050;
wire v_6051;
wire v_6052;
wire v_6053;
wire v_6054;
wire v_6055;
wire v_6056;
wire v_6059;
wire v_6060;
wire v_6061;
wire v_6062;
wire v_6063;
wire v_6064;
wire v_6065;
wire v_6066;
wire v_6067;
wire v_6068;
wire v_6071;
wire v_6072;
wire v_6073;
wire v_6074;
wire v_6075;
wire v_6076;
wire v_6077;
wire v_6078;
wire v_6079;
wire v_6080;
wire v_6083;
wire v_6084;
wire v_6085;
wire v_6086;
wire v_6087;
wire v_6088;
wire v_6089;
wire v_6090;
wire v_6091;
wire v_6092;
wire v_6095;
wire v_6096;
wire v_6097;
wire v_6098;
wire v_6099;
wire v_6100;
wire v_6101;
wire v_6102;
wire v_6103;
wire v_6104;
wire v_6105;
wire v_6106;
wire v_6107;
wire v_6108;
wire v_6109;
wire v_6110;
wire v_6111;
wire v_6112;
wire v_6113;
wire v_6114;
wire v_6115;
wire v_6116;
wire v_6117;
wire v_6118;
wire v_6119;
wire v_6120;
wire v_6123;
wire v_6124;
wire v_6125;
wire v_6126;
wire v_6127;
wire v_6128;
wire v_6129;
wire v_6130;
wire v_6131;
wire v_6132;
wire v_6134;
wire v_6135;
wire v_6136;
wire v_6137;
wire v_6138;
wire v_6139;
wire v_6140;
wire v_6142;
wire v_6143;
wire v_6144;
wire v_6145;
wire v_6146;
wire v_6147;
wire v_6148;
wire v_6149;
wire v_6150;
wire v_6151;
wire v_6152;
wire v_6153;
wire v_6154;
wire v_6155;
wire v_6156;
wire v_6157;
wire v_6158;
wire v_6159;
wire v_6160;
wire v_6161;
wire v_6162;
wire v_6163;
wire v_6164;
wire v_6165;
wire v_6166;
wire v_6167;
wire v_6168;
wire v_6169;
wire v_6170;
wire v_6171;
wire v_6172;
wire v_6173;
wire v_6174;
wire v_6175;
wire v_6176;
wire v_6177;
wire v_6178;
wire v_6179;
wire v_6180;
wire v_6181;
wire v_6182;
wire v_6183;
wire v_6184;
wire v_6187;
wire v_6188;
wire v_6189;
wire v_6190;
wire v_6191;
wire v_6192;
wire v_6193;
wire v_6194;
wire v_6195;
wire v_6196;
wire v_6199;
wire v_6200;
wire v_6201;
wire v_6202;
wire v_6203;
wire v_6204;
wire v_6205;
wire v_6206;
wire v_6207;
wire v_6208;
wire v_6211;
wire v_6212;
wire v_6213;
wire v_6214;
wire v_6215;
wire v_6216;
wire v_6217;
wire v_6218;
wire v_6219;
wire v_6220;
wire v_6223;
wire v_6224;
wire v_6225;
wire v_6226;
wire v_6227;
wire v_6228;
wire v_6229;
wire v_6230;
wire v_6231;
wire v_6232;
wire v_6235;
wire v_6236;
wire v_6237;
wire v_6238;
wire v_6239;
wire v_6240;
wire v_6241;
wire v_6242;
wire v_6243;
wire v_6244;
wire v_6247;
wire v_6248;
wire v_6249;
wire v_6250;
wire v_6251;
wire v_6252;
wire v_6253;
wire v_6254;
wire v_6255;
wire v_6256;
wire v_6257;
wire v_6258;
wire v_6259;
wire v_6260;
wire v_6261;
wire v_6262;
wire v_6263;
wire v_6264;
wire v_6265;
wire v_6266;
wire v_6267;
wire v_6268;
wire v_6269;
wire v_6270;
wire v_6271;
wire v_6272;
wire v_6275;
wire v_6276;
wire v_6277;
wire v_6278;
wire v_6279;
wire v_6280;
wire v_6281;
wire v_6282;
wire v_6283;
wire v_6284;
wire v_6286;
wire v_6288;
wire v_6289;
wire v_6290;
wire v_6291;
wire v_6292;
wire v_6293;
wire v_6294;
wire v_6295;
wire v_6296;
wire v_6297;
wire v_6298;
wire v_6299;
wire v_6300;
wire v_6301;
wire v_6302;
wire v_6303;
wire v_6304;
wire v_6305;
wire v_6306;
wire v_6307;
wire v_6308;
wire v_6309;
wire v_6310;
wire v_6311;
wire v_6312;
wire v_6313;
wire v_6314;
wire v_6315;
wire v_6316;
wire v_6319;
wire v_6320;
wire v_6321;
wire v_6322;
wire v_6323;
wire v_6324;
wire v_6325;
wire v_6326;
wire v_6327;
wire v_6328;
wire v_6331;
wire v_6332;
wire v_6333;
wire v_6334;
wire v_6335;
wire v_6336;
wire v_6337;
wire v_6338;
wire v_6339;
wire v_6340;
wire v_6343;
wire v_6344;
wire v_6345;
wire v_6346;
wire v_6347;
wire v_6348;
wire v_6349;
wire v_6350;
wire v_6351;
wire v_6352;
wire v_6355;
wire v_6356;
wire v_6357;
wire v_6358;
wire v_6359;
wire v_6360;
wire v_6361;
wire v_6362;
wire v_6363;
wire v_6364;
wire v_6367;
wire v_6368;
wire v_6369;
wire v_6370;
wire v_6371;
wire v_6372;
wire v_6373;
wire v_6374;
wire v_6375;
wire v_6376;
wire v_6379;
wire v_6380;
wire v_6381;
wire v_6382;
wire v_6383;
wire v_6384;
wire v_6385;
wire v_6386;
wire v_6387;
wire v_6388;
wire v_6389;
wire v_6390;
wire v_6391;
wire v_6392;
wire v_6393;
wire v_6394;
wire v_6395;
wire v_6396;
wire v_6397;
wire v_6398;
wire v_6399;
wire v_6400;
wire v_6401;
wire v_6402;
wire v_6403;
wire v_6404;
wire v_6407;
wire v_6408;
wire v_6409;
wire v_6410;
wire v_6411;
wire v_6412;
wire v_6413;
wire v_6414;
wire v_6415;
wire v_6416;
wire v_6418;
wire v_6419;
wire v_6420;
wire v_6421;
wire v_6422;
wire v_6424;
wire v_6425;
wire v_6426;
wire v_6427;
wire v_6428;
wire v_6429;
wire v_6430;
wire v_6431;
wire v_6432;
wire v_6433;
wire v_6434;
wire v_6435;
wire v_6436;
wire v_6437;
wire v_6438;
wire v_6439;
wire v_6440;
wire v_6441;
wire v_6442;
wire v_6443;
wire v_6444;
wire v_6445;
wire v_6446;
wire v_6447;
wire v_6448;
wire v_6449;
wire v_6450;
wire v_6451;
wire v_6452;
wire v_6453;
wire v_6454;
wire v_6455;
wire v_6456;
wire v_6457;
wire v_6458;
wire v_6459;
wire v_6460;
wire v_6461;
wire v_6462;
wire v_6463;
wire v_6464;
wire v_6465;
wire v_6466;
wire v_6467;
wire v_6468;
wire v_6469;
wire v_6470;
wire v_6471;
wire v_6472;
wire v_6473;
wire v_6474;
wire v_6475;
wire v_6476;
wire v_6477;
wire v_6478;
wire v_6479;
wire v_6480;
wire v_6483;
wire v_6484;
wire v_6485;
wire v_6486;
wire v_6487;
wire v_6488;
wire v_6489;
wire v_6490;
wire v_6491;
wire v_6492;
wire v_6495;
wire v_6496;
wire v_6497;
wire v_6498;
wire v_6499;
wire v_6500;
wire v_6501;
wire v_6502;
wire v_6503;
wire v_6504;
wire v_6507;
wire v_6508;
wire v_6509;
wire v_6510;
wire v_6511;
wire v_6512;
wire v_6513;
wire v_6514;
wire v_6515;
wire v_6516;
wire v_6519;
wire v_6520;
wire v_6521;
wire v_6522;
wire v_6523;
wire v_6524;
wire v_6525;
wire v_6526;
wire v_6527;
wire v_6528;
wire v_6531;
wire v_6532;
wire v_6533;
wire v_6534;
wire v_6535;
wire v_6536;
wire v_6537;
wire v_6538;
wire v_6539;
wire v_6540;
wire v_6543;
wire v_6544;
wire v_6545;
wire v_6546;
wire v_6547;
wire v_6548;
wire v_6549;
wire v_6550;
wire v_6551;
wire v_6552;
wire v_6553;
wire v_6554;
wire v_6555;
wire v_6556;
wire v_6557;
wire v_6558;
wire v_6559;
wire v_6560;
wire v_6561;
wire v_6562;
wire v_6563;
wire v_6564;
wire v_6565;
wire v_6566;
wire v_6567;
wire v_6568;
wire v_6571;
wire v_6572;
wire v_6573;
wire v_6574;
wire v_6575;
wire v_6576;
wire v_6577;
wire v_6578;
wire v_6579;
wire v_6580;
wire v_6582;
wire v_6584;
wire v_6585;
wire v_6586;
wire v_6587;
wire v_6588;
wire v_6589;
wire v_6590;
wire v_6591;
wire v_6592;
wire v_6593;
wire v_6594;
wire v_6595;
wire v_6596;
wire v_6597;
wire v_6598;
wire v_6599;
wire v_6600;
wire v_6601;
wire v_6602;
wire v_6603;
wire v_6604;
wire v_6605;
wire v_6606;
wire v_6607;
wire v_6608;
wire v_6609;
wire v_6610;
wire v_6611;
wire v_6612;
wire v_6615;
wire v_6616;
wire v_6617;
wire v_6618;
wire v_6619;
wire v_6620;
wire v_6621;
wire v_6622;
wire v_6623;
wire v_6624;
wire v_6627;
wire v_6628;
wire v_6629;
wire v_6630;
wire v_6631;
wire v_6632;
wire v_6633;
wire v_6634;
wire v_6635;
wire v_6636;
wire v_6639;
wire v_6640;
wire v_6641;
wire v_6642;
wire v_6643;
wire v_6644;
wire v_6645;
wire v_6646;
wire v_6647;
wire v_6648;
wire v_6651;
wire v_6652;
wire v_6653;
wire v_6654;
wire v_6655;
wire v_6656;
wire v_6657;
wire v_6658;
wire v_6659;
wire v_6660;
wire v_6663;
wire v_6664;
wire v_6665;
wire v_6666;
wire v_6667;
wire v_6668;
wire v_6669;
wire v_6670;
wire v_6671;
wire v_6672;
wire v_6675;
wire v_6676;
wire v_6677;
wire v_6678;
wire v_6679;
wire v_6680;
wire v_6681;
wire v_6682;
wire v_6683;
wire v_6684;
wire v_6685;
wire v_6686;
wire v_6687;
wire v_6688;
wire v_6689;
wire v_6690;
wire v_6691;
wire v_6692;
wire v_6693;
wire v_6694;
wire v_6695;
wire v_6696;
wire v_6697;
wire v_6698;
wire v_6699;
wire v_6700;
wire v_6703;
wire v_6704;
wire v_6705;
wire v_6706;
wire v_6707;
wire v_6708;
wire v_6709;
wire v_6710;
wire v_6711;
wire v_6712;
wire v_6714;
wire v_6715;
wire v_6716;
wire v_6717;
wire v_6718;
wire v_6719;
wire v_6721;
wire v_6722;
wire v_6723;
wire v_6724;
wire v_6725;
wire v_6726;
wire v_6727;
wire v_6728;
wire v_6729;
wire v_6730;
wire v_6731;
wire v_6732;
wire v_6733;
wire v_6734;
wire v_6735;
wire v_6736;
wire v_6737;
wire v_6738;
wire v_6739;
wire v_6740;
wire v_6741;
wire v_6742;
wire v_6743;
wire v_6744;
wire v_6745;
wire v_6746;
wire v_6747;
wire v_6748;
wire v_6749;
wire v_6750;
wire v_6751;
wire v_6752;
wire v_6753;
wire v_6754;
wire v_6755;
wire v_6756;
wire v_6757;
wire v_6758;
wire v_6759;
wire v_6760;
wire v_6761;
wire v_6762;
wire v_6765;
wire v_6766;
wire v_6767;
wire v_6768;
wire v_6769;
wire v_6770;
wire v_6771;
wire v_6772;
wire v_6773;
wire v_6774;
wire v_6777;
wire v_6778;
wire v_6779;
wire v_6780;
wire v_6781;
wire v_6782;
wire v_6783;
wire v_6784;
wire v_6785;
wire v_6786;
wire v_6789;
wire v_6790;
wire v_6791;
wire v_6792;
wire v_6793;
wire v_6794;
wire v_6795;
wire v_6796;
wire v_6797;
wire v_6798;
wire v_6801;
wire v_6802;
wire v_6803;
wire v_6804;
wire v_6805;
wire v_6806;
wire v_6807;
wire v_6808;
wire v_6809;
wire v_6810;
wire v_6813;
wire v_6814;
wire v_6815;
wire v_6816;
wire v_6817;
wire v_6818;
wire v_6819;
wire v_6820;
wire v_6821;
wire v_6822;
wire v_6825;
wire v_6826;
wire v_6827;
wire v_6828;
wire v_6829;
wire v_6830;
wire v_6831;
wire v_6832;
wire v_6833;
wire v_6834;
wire v_6835;
wire v_6836;
wire v_6837;
wire v_6838;
wire v_6839;
wire v_6840;
wire v_6841;
wire v_6842;
wire v_6843;
wire v_6844;
wire v_6845;
wire v_6846;
wire v_6847;
wire v_6848;
wire v_6849;
wire v_6850;
wire v_6853;
wire v_6854;
wire v_6855;
wire v_6856;
wire v_6857;
wire v_6858;
wire v_6859;
wire v_6860;
wire v_6861;
wire v_6862;
wire v_6864;
wire v_6866;
wire v_6867;
wire v_6868;
wire v_6869;
wire v_6870;
wire v_6871;
wire v_6872;
wire v_6873;
wire v_6874;
wire v_6875;
wire v_6876;
wire v_6877;
wire v_6878;
wire v_6879;
wire v_6880;
wire v_6881;
wire v_6882;
wire v_6883;
wire v_6884;
wire v_6885;
wire v_6886;
wire v_6887;
wire v_6888;
wire v_6889;
wire v_6890;
wire v_6891;
wire v_6892;
wire v_6893;
wire v_6894;
wire v_6897;
wire v_6898;
wire v_6899;
wire v_6900;
wire v_6901;
wire v_6902;
wire v_6903;
wire v_6904;
wire v_6905;
wire v_6906;
wire v_6909;
wire v_6910;
wire v_6911;
wire v_6912;
wire v_6913;
wire v_6914;
wire v_6915;
wire v_6916;
wire v_6917;
wire v_6918;
wire v_6921;
wire v_6922;
wire v_6923;
wire v_6924;
wire v_6925;
wire v_6926;
wire v_6927;
wire v_6928;
wire v_6929;
wire v_6930;
wire v_6933;
wire v_6934;
wire v_6935;
wire v_6936;
wire v_6937;
wire v_6938;
wire v_6939;
wire v_6940;
wire v_6941;
wire v_6942;
wire v_6945;
wire v_6946;
wire v_6947;
wire v_6948;
wire v_6949;
wire v_6950;
wire v_6951;
wire v_6952;
wire v_6953;
wire v_6954;
wire v_6957;
wire v_6958;
wire v_6959;
wire v_6960;
wire v_6961;
wire v_6962;
wire v_6963;
wire v_6964;
wire v_6965;
wire v_6966;
wire v_6967;
wire v_6968;
wire v_6969;
wire v_6970;
wire v_6971;
wire v_6972;
wire v_6973;
wire v_6974;
wire v_6975;
wire v_6976;
wire v_6977;
wire v_6978;
wire v_6979;
wire v_6980;
wire v_6981;
wire v_6982;
wire v_6985;
wire v_6986;
wire v_6987;
wire v_6988;
wire v_6989;
wire v_6990;
wire v_6991;
wire v_6992;
wire v_6993;
wire v_6994;
wire v_6996;
wire v_6997;
wire v_6998;
wire v_6999;
wire v_7000;
wire v_7002;
wire v_7003;
wire v_7004;
wire v_7005;
wire v_7006;
wire v_7007;
wire v_7008;
wire v_7009;
wire v_7010;
wire v_7011;
wire v_7012;
wire v_7013;
wire v_7014;
wire v_7015;
wire v_7016;
wire v_7017;
wire v_7018;
wire v_7019;
wire v_7020;
wire v_7021;
wire v_7022;
wire v_7023;
wire v_7024;
wire v_7025;
wire v_7026;
wire v_7027;
wire v_7028;
wire v_7029;
wire v_7030;
wire v_7031;
wire v_7032;
wire v_7033;
wire v_7034;
wire v_7035;
wire v_7036;
wire v_7037;
wire v_7038;
wire v_7039;
wire v_7040;
wire v_7041;
wire v_7042;
wire v_7043;
wire v_7044;
wire v_7045;
wire v_7046;
wire v_7047;
wire v_7048;
wire v_7049;
wire v_7050;
wire v_7053;
wire v_7054;
wire v_7055;
wire v_7056;
wire v_7057;
wire v_7058;
wire v_7059;
wire v_7060;
wire v_7061;
wire v_7062;
wire v_7065;
wire v_7066;
wire v_7067;
wire v_7068;
wire v_7069;
wire v_7070;
wire v_7071;
wire v_7072;
wire v_7073;
wire v_7074;
wire v_7077;
wire v_7078;
wire v_7079;
wire v_7080;
wire v_7081;
wire v_7082;
wire v_7083;
wire v_7084;
wire v_7085;
wire v_7086;
wire v_7089;
wire v_7090;
wire v_7091;
wire v_7092;
wire v_7093;
wire v_7094;
wire v_7095;
wire v_7096;
wire v_7097;
wire v_7098;
wire v_7101;
wire v_7102;
wire v_7103;
wire v_7104;
wire v_7105;
wire v_7106;
wire v_7107;
wire v_7108;
wire v_7109;
wire v_7110;
wire v_7113;
wire v_7114;
wire v_7115;
wire v_7116;
wire v_7117;
wire v_7118;
wire v_7119;
wire v_7120;
wire v_7121;
wire v_7122;
wire v_7123;
wire v_7124;
wire v_7125;
wire v_7126;
wire v_7127;
wire v_7128;
wire v_7129;
wire v_7130;
wire v_7131;
wire v_7132;
wire v_7133;
wire v_7134;
wire v_7135;
wire v_7136;
wire v_7137;
wire v_7138;
wire v_7141;
wire v_7142;
wire v_7143;
wire v_7144;
wire v_7145;
wire v_7146;
wire v_7147;
wire v_7148;
wire v_7149;
wire v_7150;
wire v_7152;
wire v_7154;
wire v_7155;
wire v_7156;
wire v_7157;
wire v_7158;
wire v_7159;
wire v_7160;
wire v_7161;
wire v_7162;
wire v_7163;
wire v_7164;
wire v_7165;
wire v_7166;
wire v_7167;
wire v_7168;
wire v_7169;
wire v_7170;
wire v_7171;
wire v_7172;
wire v_7173;
wire v_7174;
wire v_7175;
wire v_7176;
wire v_7177;
wire v_7178;
wire v_7179;
wire v_7180;
wire v_7181;
wire v_7182;
wire v_7185;
wire v_7186;
wire v_7187;
wire v_7188;
wire v_7189;
wire v_7190;
wire v_7191;
wire v_7192;
wire v_7193;
wire v_7194;
wire v_7197;
wire v_7198;
wire v_7199;
wire v_7200;
wire v_7201;
wire v_7202;
wire v_7203;
wire v_7204;
wire v_7205;
wire v_7206;
wire v_7209;
wire v_7210;
wire v_7211;
wire v_7212;
wire v_7213;
wire v_7214;
wire v_7215;
wire v_7216;
wire v_7217;
wire v_7218;
wire v_7221;
wire v_7222;
wire v_7223;
wire v_7224;
wire v_7225;
wire v_7226;
wire v_7227;
wire v_7228;
wire v_7229;
wire v_7230;
wire v_7233;
wire v_7234;
wire v_7235;
wire v_7236;
wire v_7237;
wire v_7238;
wire v_7239;
wire v_7240;
wire v_7241;
wire v_7242;
wire v_7245;
wire v_7246;
wire v_7247;
wire v_7248;
wire v_7249;
wire v_7250;
wire v_7251;
wire v_7252;
wire v_7253;
wire v_7254;
wire v_7255;
wire v_7256;
wire v_7257;
wire v_7258;
wire v_7259;
wire v_7260;
wire v_7261;
wire v_7262;
wire v_7263;
wire v_7264;
wire v_7265;
wire v_7266;
wire v_7267;
wire v_7268;
wire v_7269;
wire v_7270;
wire v_7273;
wire v_7274;
wire v_7275;
wire v_7276;
wire v_7277;
wire v_7278;
wire v_7279;
wire v_7280;
wire v_7281;
wire v_7282;
wire v_7284;
wire v_7285;
wire v_7286;
wire v_7287;
wire v_7288;
wire v_7289;
wire v_7290;
wire v_7291;
wire v_7293;
wire v_7294;
wire v_7295;
wire v_7296;
wire v_7297;
wire v_7298;
wire v_7299;
wire v_7300;
wire v_7301;
wire v_7302;
wire v_7303;
wire v_7304;
wire v_7305;
wire v_7306;
wire v_7307;
wire v_7308;
wire v_7309;
wire v_7310;
wire v_7311;
wire v_7312;
wire v_7313;
wire v_7314;
wire v_7315;
wire v_7316;
wire v_7317;
wire v_7318;
wire v_7319;
wire v_7320;
wire v_7321;
wire v_7322;
wire v_7323;
wire v_7324;
wire v_7325;
wire v_7326;
wire v_7327;
wire v_7328;
wire v_7329;
wire v_7330;
wire v_7331;
wire v_7332;
wire v_7333;
wire v_7334;
wire v_7335;
wire v_7336;
wire v_7339;
wire v_7340;
wire v_7341;
wire v_7342;
wire v_7343;
wire v_7344;
wire v_7345;
wire v_7346;
wire v_7347;
wire v_7348;
wire v_7351;
wire v_7352;
wire v_7353;
wire v_7354;
wire v_7355;
wire v_7356;
wire v_7357;
wire v_7358;
wire v_7359;
wire v_7360;
wire v_7363;
wire v_7364;
wire v_7365;
wire v_7366;
wire v_7367;
wire v_7368;
wire v_7369;
wire v_7370;
wire v_7371;
wire v_7372;
wire v_7375;
wire v_7376;
wire v_7377;
wire v_7378;
wire v_7379;
wire v_7380;
wire v_7381;
wire v_7382;
wire v_7383;
wire v_7384;
wire v_7387;
wire v_7388;
wire v_7389;
wire v_7390;
wire v_7391;
wire v_7392;
wire v_7393;
wire v_7394;
wire v_7395;
wire v_7396;
wire v_7399;
wire v_7400;
wire v_7401;
wire v_7402;
wire v_7403;
wire v_7404;
wire v_7405;
wire v_7406;
wire v_7407;
wire v_7408;
wire v_7409;
wire v_7410;
wire v_7411;
wire v_7412;
wire v_7413;
wire v_7414;
wire v_7415;
wire v_7416;
wire v_7417;
wire v_7418;
wire v_7419;
wire v_7420;
wire v_7421;
wire v_7422;
wire v_7423;
wire v_7424;
wire v_7427;
wire v_7428;
wire v_7429;
wire v_7430;
wire v_7431;
wire v_7432;
wire v_7433;
wire v_7434;
wire v_7435;
wire v_7436;
wire v_7438;
wire v_7440;
wire v_7441;
wire v_7442;
wire v_7443;
wire v_7444;
wire v_7445;
wire v_7446;
wire v_7447;
wire v_7448;
wire v_7449;
wire v_7450;
wire v_7451;
wire v_7452;
wire v_7453;
wire v_7454;
wire v_7455;
wire v_7456;
wire v_7457;
wire v_7458;
wire v_7459;
wire v_7460;
wire v_7461;
wire v_7462;
wire v_7463;
wire v_7464;
wire v_7465;
wire v_7466;
wire v_7467;
wire v_7468;
wire v_7471;
wire v_7472;
wire v_7473;
wire v_7474;
wire v_7475;
wire v_7476;
wire v_7477;
wire v_7478;
wire v_7479;
wire v_7480;
wire v_7483;
wire v_7484;
wire v_7485;
wire v_7486;
wire v_7487;
wire v_7488;
wire v_7489;
wire v_7490;
wire v_7491;
wire v_7492;
wire v_7495;
wire v_7496;
wire v_7497;
wire v_7498;
wire v_7499;
wire v_7500;
wire v_7501;
wire v_7502;
wire v_7503;
wire v_7504;
wire v_7507;
wire v_7508;
wire v_7509;
wire v_7510;
wire v_7511;
wire v_7512;
wire v_7513;
wire v_7514;
wire v_7515;
wire v_7516;
wire v_7519;
wire v_7520;
wire v_7521;
wire v_7522;
wire v_7523;
wire v_7524;
wire v_7525;
wire v_7526;
wire v_7527;
wire v_7528;
wire v_7531;
wire v_7532;
wire v_7533;
wire v_7534;
wire v_7535;
wire v_7536;
wire v_7537;
wire v_7538;
wire v_7539;
wire v_7540;
wire v_7541;
wire v_7542;
wire v_7543;
wire v_7544;
wire v_7545;
wire v_7546;
wire v_7547;
wire v_7548;
wire v_7549;
wire v_7550;
wire v_7551;
wire v_7552;
wire v_7553;
wire v_7554;
wire v_7555;
wire v_7556;
wire v_7559;
wire v_7560;
wire v_7561;
wire v_7562;
wire v_7563;
wire v_7564;
wire v_7565;
wire v_7566;
wire v_7567;
wire v_7568;
wire v_7570;
wire v_7571;
wire v_7572;
wire v_7573;
wire v_7574;
wire v_7576;
wire v_7577;
wire v_7578;
wire v_7579;
wire v_7580;
wire v_7581;
wire v_7582;
wire v_7583;
wire v_7584;
wire v_7585;
wire v_7586;
wire v_7587;
wire v_7588;
wire v_7589;
wire v_7590;
wire v_7591;
wire v_7592;
wire v_7593;
wire v_7594;
wire v_7595;
wire v_7596;
wire v_7597;
wire v_7598;
wire v_7599;
wire v_7600;
wire v_7601;
wire v_7602;
wire v_7603;
wire v_7604;
wire v_7605;
wire v_7606;
wire v_7607;
wire v_7608;
wire v_7609;
wire v_7610;
wire v_7611;
wire v_7612;
wire v_7613;
wire v_7614;
wire v_7615;
wire v_7616;
wire v_7617;
wire v_7618;
wire v_7619;
wire v_7620;
wire v_7621;
wire v_7622;
wire v_7623;
wire v_7624;
wire v_7625;
wire v_7626;
wire v_7627;
wire v_7628;
wire v_7629;
wire v_7630;
wire v_7631;
wire v_7632;
wire v_7633;
wire v_7634;
wire v_7635;
wire v_7636;
wire v_7637;
wire v_7638;
wire v_7639;
wire v_7640;
wire v_7643;
wire v_7644;
wire v_7645;
wire v_7646;
wire v_7647;
wire v_7648;
wire v_7649;
wire v_7650;
wire v_7651;
wire v_7652;
wire v_7655;
wire v_7656;
wire v_7657;
wire v_7658;
wire v_7659;
wire v_7660;
wire v_7661;
wire v_7662;
wire v_7663;
wire v_7664;
wire v_7667;
wire v_7668;
wire v_7669;
wire v_7670;
wire v_7671;
wire v_7672;
wire v_7673;
wire v_7674;
wire v_7675;
wire v_7676;
wire v_7679;
wire v_7680;
wire v_7681;
wire v_7682;
wire v_7683;
wire v_7684;
wire v_7685;
wire v_7686;
wire v_7687;
wire v_7688;
wire v_7691;
wire v_7692;
wire v_7693;
wire v_7694;
wire v_7695;
wire v_7696;
wire v_7697;
wire v_7698;
wire v_7699;
wire v_7700;
wire v_7703;
wire v_7704;
wire v_7705;
wire v_7706;
wire v_7707;
wire v_7708;
wire v_7709;
wire v_7710;
wire v_7711;
wire v_7712;
wire v_7713;
wire v_7714;
wire v_7715;
wire v_7716;
wire v_7717;
wire v_7718;
wire v_7719;
wire v_7720;
wire v_7721;
wire v_7722;
wire v_7723;
wire v_7724;
wire v_7725;
wire v_7726;
wire v_7727;
wire v_7728;
wire v_7731;
wire v_7732;
wire v_7733;
wire v_7734;
wire v_7735;
wire v_7736;
wire v_7737;
wire v_7738;
wire v_7739;
wire v_7740;
wire v_7742;
wire v_7744;
wire v_7745;
wire v_7746;
wire v_7747;
wire v_7748;
wire v_7749;
wire v_7750;
wire v_7751;
wire v_7752;
wire v_7753;
wire v_7754;
wire v_7755;
wire v_7756;
wire v_7757;
wire v_7758;
wire v_7759;
wire v_7760;
wire v_7761;
wire v_7762;
wire v_7763;
wire v_7764;
wire v_7765;
wire v_7766;
wire v_7767;
wire v_7768;
wire v_7769;
wire v_7770;
wire v_7771;
wire v_7772;
wire v_7775;
wire v_7776;
wire v_7777;
wire v_7778;
wire v_7779;
wire v_7780;
wire v_7781;
wire v_7782;
wire v_7783;
wire v_7784;
wire v_7787;
wire v_7788;
wire v_7789;
wire v_7790;
wire v_7791;
wire v_7792;
wire v_7793;
wire v_7794;
wire v_7795;
wire v_7796;
wire v_7799;
wire v_7800;
wire v_7801;
wire v_7802;
wire v_7803;
wire v_7804;
wire v_7805;
wire v_7806;
wire v_7807;
wire v_7808;
wire v_7811;
wire v_7812;
wire v_7813;
wire v_7814;
wire v_7815;
wire v_7816;
wire v_7817;
wire v_7818;
wire v_7819;
wire v_7820;
wire v_7823;
wire v_7824;
wire v_7825;
wire v_7826;
wire v_7827;
wire v_7828;
wire v_7829;
wire v_7830;
wire v_7831;
wire v_7832;
wire v_7835;
wire v_7836;
wire v_7837;
wire v_7838;
wire v_7839;
wire v_7840;
wire v_7841;
wire v_7842;
wire v_7843;
wire v_7844;
wire v_7845;
wire v_7846;
wire v_7847;
wire v_7848;
wire v_7849;
wire v_7850;
wire v_7851;
wire v_7852;
wire v_7853;
wire v_7854;
wire v_7855;
wire v_7856;
wire v_7857;
wire v_7858;
wire v_7859;
wire v_7860;
wire v_7863;
wire v_7864;
wire v_7865;
wire v_7866;
wire v_7867;
wire v_7868;
wire v_7869;
wire v_7870;
wire v_7871;
wire v_7872;
wire v_7874;
wire v_7875;
wire v_7876;
wire v_7877;
wire v_7878;
wire v_7879;
wire v_7881;
wire v_7882;
wire v_7883;
wire v_7884;
wire v_7885;
wire v_7886;
wire v_7887;
wire v_7888;
wire v_7889;
wire v_7890;
wire v_7891;
wire v_7892;
wire v_7893;
wire v_7894;
wire v_7895;
wire v_7896;
wire v_7897;
wire v_7898;
wire v_7899;
wire v_7900;
wire v_7901;
wire v_7902;
wire v_7903;
wire v_7904;
wire v_7905;
wire v_7906;
wire v_7907;
wire v_7908;
wire v_7909;
wire v_7910;
wire v_7911;
wire v_7912;
wire v_7913;
wire v_7914;
wire v_7915;
wire v_7916;
wire v_7917;
wire v_7918;
wire v_7919;
wire v_7920;
wire v_7921;
wire v_7922;
wire v_7925;
wire v_7926;
wire v_7927;
wire v_7928;
wire v_7929;
wire v_7930;
wire v_7931;
wire v_7932;
wire v_7933;
wire v_7934;
wire v_7937;
wire v_7938;
wire v_7939;
wire v_7940;
wire v_7941;
wire v_7942;
wire v_7943;
wire v_7944;
wire v_7945;
wire v_7946;
wire v_7949;
wire v_7950;
wire v_7951;
wire v_7952;
wire v_7953;
wire v_7954;
wire v_7955;
wire v_7956;
wire v_7957;
wire v_7958;
wire v_7961;
wire v_7962;
wire v_7963;
wire v_7964;
wire v_7965;
wire v_7966;
wire v_7967;
wire v_7968;
wire v_7969;
wire v_7970;
wire v_7973;
wire v_7974;
wire v_7975;
wire v_7976;
wire v_7977;
wire v_7978;
wire v_7979;
wire v_7980;
wire v_7981;
wire v_7982;
wire v_7985;
wire v_7986;
wire v_7987;
wire v_7988;
wire v_7989;
wire v_7990;
wire v_7991;
wire v_7992;
wire v_7993;
wire v_7994;
wire v_7995;
wire v_7996;
wire v_7997;
wire v_7998;
wire v_7999;
wire v_8000;
wire v_8001;
wire v_8002;
wire v_8003;
wire v_8004;
wire v_8005;
wire v_8006;
wire v_8007;
wire v_8008;
wire v_8009;
wire v_8010;
wire v_8013;
wire v_8014;
wire v_8015;
wire v_8016;
wire v_8017;
wire v_8018;
wire v_8019;
wire v_8020;
wire v_8021;
wire v_8022;
wire v_8024;
wire v_8026;
wire v_8027;
wire v_8028;
wire v_8029;
wire v_8030;
wire v_8031;
wire v_8032;
wire v_8033;
wire v_8034;
wire v_8035;
wire v_8036;
wire v_8037;
wire v_8038;
wire v_8039;
wire v_8040;
wire v_8041;
wire v_8042;
wire v_8043;
wire v_8044;
wire v_8045;
wire v_8046;
wire v_8047;
wire v_8048;
wire v_8049;
wire v_8050;
wire v_8051;
wire v_8052;
wire v_8053;
wire v_8054;
wire v_8057;
wire v_8058;
wire v_8059;
wire v_8060;
wire v_8061;
wire v_8062;
wire v_8063;
wire v_8064;
wire v_8065;
wire v_8066;
wire v_8069;
wire v_8070;
wire v_8071;
wire v_8072;
wire v_8073;
wire v_8074;
wire v_8075;
wire v_8076;
wire v_8077;
wire v_8078;
wire v_8081;
wire v_8082;
wire v_8083;
wire v_8084;
wire v_8085;
wire v_8086;
wire v_8087;
wire v_8088;
wire v_8089;
wire v_8090;
wire v_8093;
wire v_8094;
wire v_8095;
wire v_8096;
wire v_8097;
wire v_8098;
wire v_8099;
wire v_8100;
wire v_8101;
wire v_8102;
wire v_8105;
wire v_8106;
wire v_8107;
wire v_8108;
wire v_8109;
wire v_8110;
wire v_8111;
wire v_8112;
wire v_8113;
wire v_8114;
wire v_8117;
wire v_8118;
wire v_8119;
wire v_8120;
wire v_8121;
wire v_8122;
wire v_8123;
wire v_8124;
wire v_8125;
wire v_8126;
wire v_8127;
wire v_8128;
wire v_8129;
wire v_8130;
wire v_8131;
wire v_8132;
wire v_8133;
wire v_8134;
wire v_8135;
wire v_8136;
wire v_8137;
wire v_8138;
wire v_8139;
wire v_8140;
wire v_8141;
wire v_8142;
wire v_8145;
wire v_8146;
wire v_8147;
wire v_8148;
wire v_8149;
wire v_8150;
wire v_8151;
wire v_8152;
wire v_8153;
wire v_8154;
wire v_8156;
wire v_8157;
wire v_8158;
wire v_8159;
wire v_8160;
wire v_8162;
wire v_8163;
wire v_8164;
wire v_8165;
wire v_8166;
wire v_8167;
wire v_8168;
wire v_8169;
wire v_8170;
wire v_8171;
wire v_8172;
wire v_8173;
wire v_8174;
wire v_8175;
wire v_8176;
wire v_8177;
wire v_8178;
wire v_8179;
wire v_8180;
wire v_8181;
wire v_8182;
wire v_8183;
wire v_8184;
wire v_8185;
wire v_8186;
wire v_8187;
wire v_8188;
wire v_8189;
wire v_8190;
wire v_8191;
wire v_8192;
wire v_8193;
wire v_8194;
wire v_8195;
wire v_8196;
wire v_8197;
wire v_8198;
wire v_8199;
wire v_8200;
wire v_8201;
wire v_8202;
wire v_8203;
wire v_8204;
wire v_8205;
wire v_8206;
wire v_8207;
wire v_8208;
wire v_8209;
wire v_8210;
wire v_8213;
wire v_8214;
wire v_8215;
wire v_8216;
wire v_8217;
wire v_8218;
wire v_8219;
wire v_8220;
wire v_8221;
wire v_8222;
wire v_8225;
wire v_8226;
wire v_8227;
wire v_8228;
wire v_8229;
wire v_8230;
wire v_8231;
wire v_8232;
wire v_8233;
wire v_8234;
wire v_8237;
wire v_8238;
wire v_8239;
wire v_8240;
wire v_8241;
wire v_8242;
wire v_8243;
wire v_8244;
wire v_8245;
wire v_8246;
wire v_8249;
wire v_8250;
wire v_8251;
wire v_8252;
wire v_8253;
wire v_8254;
wire v_8255;
wire v_8256;
wire v_8257;
wire v_8258;
wire v_8261;
wire v_8262;
wire v_8263;
wire v_8264;
wire v_8265;
wire v_8266;
wire v_8267;
wire v_8268;
wire v_8269;
wire v_8270;
wire v_8273;
wire v_8274;
wire v_8275;
wire v_8276;
wire v_8277;
wire v_8278;
wire v_8279;
wire v_8280;
wire v_8281;
wire v_8282;
wire v_8283;
wire v_8284;
wire v_8285;
wire v_8286;
wire v_8287;
wire v_8288;
wire v_8289;
wire v_8290;
wire v_8291;
wire v_8292;
wire v_8293;
wire v_8294;
wire v_8295;
wire v_8296;
wire v_8297;
wire v_8298;
wire v_8301;
wire v_8302;
wire v_8303;
wire v_8304;
wire v_8305;
wire v_8306;
wire v_8307;
wire v_8308;
wire v_8309;
wire v_8310;
wire v_8312;
wire v_8314;
wire v_8315;
wire v_8316;
wire v_8317;
wire v_8318;
wire v_8319;
wire v_8320;
wire v_8321;
wire v_8322;
wire v_8323;
wire v_8324;
wire v_8325;
wire v_8326;
wire v_8327;
wire v_8328;
wire v_8329;
wire v_8330;
wire v_8331;
wire v_8332;
wire v_8333;
wire v_8334;
wire v_8335;
wire v_8336;
wire v_8337;
wire v_8338;
wire v_8339;
wire v_8340;
wire v_8341;
wire v_8342;
wire v_8345;
wire v_8346;
wire v_8347;
wire v_8348;
wire v_8349;
wire v_8350;
wire v_8351;
wire v_8352;
wire v_8353;
wire v_8354;
wire v_8357;
wire v_8358;
wire v_8359;
wire v_8360;
wire v_8361;
wire v_8362;
wire v_8363;
wire v_8364;
wire v_8365;
wire v_8366;
wire v_8369;
wire v_8370;
wire v_8371;
wire v_8372;
wire v_8373;
wire v_8374;
wire v_8375;
wire v_8376;
wire v_8377;
wire v_8378;
wire v_8381;
wire v_8382;
wire v_8383;
wire v_8384;
wire v_8385;
wire v_8386;
wire v_8387;
wire v_8388;
wire v_8389;
wire v_8390;
wire v_8393;
wire v_8394;
wire v_8395;
wire v_8396;
wire v_8397;
wire v_8398;
wire v_8399;
wire v_8400;
wire v_8401;
wire v_8402;
wire v_8405;
wire v_8406;
wire v_8407;
wire v_8408;
wire v_8409;
wire v_8410;
wire v_8411;
wire v_8412;
wire v_8413;
wire v_8414;
wire v_8415;
wire v_8416;
wire v_8417;
wire v_8418;
wire v_8419;
wire v_8420;
wire v_8421;
wire v_8422;
wire v_8423;
wire v_8424;
wire v_8425;
wire v_8426;
wire v_8427;
wire v_8428;
wire v_8429;
wire v_8430;
wire v_8433;
wire v_8434;
wire v_8435;
wire v_8436;
wire v_8437;
wire v_8438;
wire v_8439;
wire v_8440;
wire v_8441;
wire v_8442;
wire v_8444;
wire v_8445;
wire v_8446;
wire v_8447;
wire v_8448;
wire v_8449;
wire v_8450;
wire v_8452;
wire v_8453;
wire v_8454;
wire v_8455;
wire v_8456;
wire v_8457;
wire v_8458;
wire v_8459;
wire v_8460;
wire v_8461;
wire v_8462;
wire v_8463;
wire v_8464;
wire v_8465;
wire v_8466;
wire v_8467;
wire v_8468;
wire v_8469;
wire v_8470;
wire v_8471;
wire v_8472;
wire v_8473;
wire v_8474;
wire v_8475;
wire v_8476;
wire v_8477;
wire v_8478;
wire v_8479;
wire v_8480;
wire v_8481;
wire v_8482;
wire v_8483;
wire v_8484;
wire v_8485;
wire v_8486;
wire v_8487;
wire v_8488;
wire v_8489;
wire v_8490;
wire v_8491;
wire v_8492;
wire v_8493;
wire v_8494;
wire v_8497;
wire v_8498;
wire v_8499;
wire v_8500;
wire v_8501;
wire v_8502;
wire v_8503;
wire v_8504;
wire v_8505;
wire v_8506;
wire v_8509;
wire v_8510;
wire v_8511;
wire v_8512;
wire v_8513;
wire v_8514;
wire v_8515;
wire v_8516;
wire v_8517;
wire v_8518;
wire v_8521;
wire v_8522;
wire v_8523;
wire v_8524;
wire v_8525;
wire v_8526;
wire v_8527;
wire v_8528;
wire v_8529;
wire v_8530;
wire v_8533;
wire v_8534;
wire v_8535;
wire v_8536;
wire v_8537;
wire v_8538;
wire v_8539;
wire v_8540;
wire v_8541;
wire v_8542;
wire v_8545;
wire v_8546;
wire v_8547;
wire v_8548;
wire v_8549;
wire v_8550;
wire v_8551;
wire v_8552;
wire v_8553;
wire v_8554;
wire v_8557;
wire v_8558;
wire v_8559;
wire v_8560;
wire v_8561;
wire v_8562;
wire v_8563;
wire v_8564;
wire v_8565;
wire v_8566;
wire v_8567;
wire v_8568;
wire v_8569;
wire v_8570;
wire v_8571;
wire v_8572;
wire v_8573;
wire v_8574;
wire v_8575;
wire v_8576;
wire v_8577;
wire v_8578;
wire v_8579;
wire v_8580;
wire v_8581;
wire v_8582;
wire v_8585;
wire v_8586;
wire v_8587;
wire v_8588;
wire v_8589;
wire v_8590;
wire v_8591;
wire v_8592;
wire v_8593;
wire v_8594;
wire v_8596;
wire v_8598;
wire v_8599;
wire v_8600;
wire v_8601;
wire v_8602;
wire v_8603;
wire v_8604;
wire v_8605;
wire v_8606;
wire v_8607;
wire v_8608;
wire v_8609;
wire v_8610;
wire v_8611;
wire v_8612;
wire v_8613;
wire v_8614;
wire v_8615;
wire v_8616;
wire v_8617;
wire v_8618;
wire v_8619;
wire v_8620;
wire v_8621;
wire v_8622;
wire v_8623;
wire v_8624;
wire v_8625;
wire v_8626;
wire v_8629;
wire v_8630;
wire v_8631;
wire v_8632;
wire v_8633;
wire v_8634;
wire v_8635;
wire v_8636;
wire v_8637;
wire v_8638;
wire v_8641;
wire v_8642;
wire v_8643;
wire v_8644;
wire v_8645;
wire v_8646;
wire v_8647;
wire v_8648;
wire v_8649;
wire v_8650;
wire v_8653;
wire v_8654;
wire v_8655;
wire v_8656;
wire v_8657;
wire v_8658;
wire v_8659;
wire v_8660;
wire v_8661;
wire v_8662;
wire v_8665;
wire v_8666;
wire v_8667;
wire v_8668;
wire v_8669;
wire v_8670;
wire v_8671;
wire v_8672;
wire v_8673;
wire v_8674;
wire v_8677;
wire v_8678;
wire v_8679;
wire v_8680;
wire v_8681;
wire v_8682;
wire v_8683;
wire v_8684;
wire v_8685;
wire v_8686;
wire v_8689;
wire v_8690;
wire v_8691;
wire v_8692;
wire v_8693;
wire v_8694;
wire v_8695;
wire v_8696;
wire v_8697;
wire v_8698;
wire v_8699;
wire v_8700;
wire v_8701;
wire v_8702;
wire v_8703;
wire v_8704;
wire v_8705;
wire v_8706;
wire v_8707;
wire v_8708;
wire v_8709;
wire v_8710;
wire v_8711;
wire v_8712;
wire v_8713;
wire v_8714;
wire v_8717;
wire v_8718;
wire v_8719;
wire v_8720;
wire v_8721;
wire v_8722;
wire v_8723;
wire v_8724;
wire v_8725;
wire v_8726;
wire v_8728;
wire v_8729;
wire v_8730;
wire v_8731;
wire v_8732;
wire v_8734;
wire v_8735;
wire v_8736;
wire v_8737;
wire v_8738;
wire v_8739;
wire v_8740;
wire v_8741;
wire v_8742;
wire v_8743;
wire v_8744;
wire v_8745;
wire v_8746;
wire v_8747;
wire v_8748;
wire v_8749;
wire v_8750;
wire v_8751;
wire v_8752;
wire v_8753;
wire v_8754;
wire v_8755;
wire v_8756;
wire v_8757;
wire v_8758;
wire v_8759;
wire v_8760;
wire v_8761;
wire v_8762;
wire v_8763;
wire v_8764;
wire v_8765;
wire v_8766;
wire v_8767;
wire v_8768;
wire v_8769;
wire v_8770;
wire v_8771;
wire v_8772;
wire v_8773;
wire v_8774;
wire v_8775;
wire v_8776;
wire v_8777;
wire v_8778;
wire v_8779;
wire v_8780;
wire v_8781;
wire v_8782;
wire v_8783;
wire v_8784;
wire v_8785;
wire v_8786;
wire v_8787;
wire v_8788;
wire v_8789;
wire v_8790;
wire v_8793;
wire v_8794;
wire v_8795;
wire v_8796;
wire v_8797;
wire v_8798;
wire v_8799;
wire v_8800;
wire v_8801;
wire v_8802;
wire v_8805;
wire v_8806;
wire v_8807;
wire v_8808;
wire v_8809;
wire v_8810;
wire v_8811;
wire v_8812;
wire v_8813;
wire v_8814;
wire v_8817;
wire v_8818;
wire v_8819;
wire v_8820;
wire v_8821;
wire v_8822;
wire v_8823;
wire v_8824;
wire v_8825;
wire v_8826;
wire v_8829;
wire v_8830;
wire v_8831;
wire v_8832;
wire v_8833;
wire v_8834;
wire v_8835;
wire v_8836;
wire v_8837;
wire v_8838;
wire v_8841;
wire v_8842;
wire v_8843;
wire v_8844;
wire v_8845;
wire v_8846;
wire v_8847;
wire v_8848;
wire v_8849;
wire v_8850;
wire v_8853;
wire v_8854;
wire v_8855;
wire v_8856;
wire v_8857;
wire v_8858;
wire v_8859;
wire v_8860;
wire v_8861;
wire v_8862;
wire v_8863;
wire v_8864;
wire v_8865;
wire v_8866;
wire v_8867;
wire v_8868;
wire v_8869;
wire v_8870;
wire v_8871;
wire v_8872;
wire v_8873;
wire v_8874;
wire v_8875;
wire v_8876;
wire v_8877;
wire v_8878;
wire v_8881;
wire v_8882;
wire v_8883;
wire v_8884;
wire v_8885;
wire v_8886;
wire v_8887;
wire v_8888;
wire v_8889;
wire v_8890;
wire v_8892;
wire v_8894;
wire v_8895;
wire v_8896;
wire v_8897;
wire v_8898;
wire v_8899;
wire v_8900;
wire v_8901;
wire v_8902;
wire v_8903;
wire v_8904;
wire v_8905;
wire v_8906;
wire v_8907;
wire v_8908;
wire v_8909;
wire v_8910;
wire v_8911;
wire v_8912;
wire v_8913;
wire v_8914;
wire v_8915;
wire v_8916;
wire v_8917;
wire v_8918;
wire v_8919;
wire v_8920;
wire v_8921;
wire v_8922;
wire v_8925;
wire v_8926;
wire v_8927;
wire v_8928;
wire v_8929;
wire v_8930;
wire v_8931;
wire v_8932;
wire v_8933;
wire v_8934;
wire v_8937;
wire v_8938;
wire v_8939;
wire v_8940;
wire v_8941;
wire v_8942;
wire v_8943;
wire v_8944;
wire v_8945;
wire v_8946;
wire v_8949;
wire v_8950;
wire v_8951;
wire v_8952;
wire v_8953;
wire v_8954;
wire v_8955;
wire v_8956;
wire v_8957;
wire v_8958;
wire v_8961;
wire v_8962;
wire v_8963;
wire v_8964;
wire v_8965;
wire v_8966;
wire v_8967;
wire v_8968;
wire v_8969;
wire v_8970;
wire v_8973;
wire v_8974;
wire v_8975;
wire v_8976;
wire v_8977;
wire v_8978;
wire v_8979;
wire v_8980;
wire v_8981;
wire v_8982;
wire v_8985;
wire v_8986;
wire v_8987;
wire v_8988;
wire v_8989;
wire v_8990;
wire v_8991;
wire v_8992;
wire v_8993;
wire v_8994;
wire v_8995;
wire v_8996;
wire v_8997;
wire v_8998;
wire v_8999;
wire v_9000;
wire v_9001;
wire v_9002;
wire v_9003;
wire v_9004;
wire v_9005;
wire v_9006;
wire v_9007;
wire v_9008;
wire v_9009;
wire v_9010;
wire v_9013;
wire v_9014;
wire v_9015;
wire v_9016;
wire v_9017;
wire v_9018;
wire v_9019;
wire v_9020;
wire v_9021;
wire v_9022;
wire v_9024;
wire v_9025;
wire v_9026;
wire v_9027;
wire v_9028;
wire v_9029;
wire v_9031;
wire v_9032;
wire v_9033;
wire v_9034;
wire v_9035;
wire v_9036;
wire v_9037;
wire v_9038;
wire v_9039;
wire v_9040;
wire v_9041;
wire v_9042;
wire v_9043;
wire v_9044;
wire v_9045;
wire v_9046;
wire v_9047;
wire v_9048;
wire v_9049;
wire v_9050;
wire v_9051;
wire v_9052;
wire v_9053;
wire v_9054;
wire v_9055;
wire v_9056;
wire v_9057;
wire v_9058;
wire v_9059;
wire v_9060;
wire v_9061;
wire v_9062;
wire v_9063;
wire v_9064;
wire v_9065;
wire v_9066;
wire v_9067;
wire v_9068;
wire v_9069;
wire v_9070;
wire v_9071;
wire v_9072;
wire v_9075;
wire v_9076;
wire v_9077;
wire v_9078;
wire v_9079;
wire v_9080;
wire v_9081;
wire v_9082;
wire v_9083;
wire v_9084;
wire v_9087;
wire v_9088;
wire v_9089;
wire v_9090;
wire v_9091;
wire v_9092;
wire v_9093;
wire v_9094;
wire v_9095;
wire v_9096;
wire v_9099;
wire v_9100;
wire v_9101;
wire v_9102;
wire v_9103;
wire v_9104;
wire v_9105;
wire v_9106;
wire v_9107;
wire v_9108;
wire v_9111;
wire v_9112;
wire v_9113;
wire v_9114;
wire v_9115;
wire v_9116;
wire v_9117;
wire v_9118;
wire v_9119;
wire v_9120;
wire v_9123;
wire v_9124;
wire v_9125;
wire v_9126;
wire v_9127;
wire v_9128;
wire v_9129;
wire v_9130;
wire v_9131;
wire v_9132;
wire v_9135;
wire v_9136;
wire v_9137;
wire v_9138;
wire v_9139;
wire v_9140;
wire v_9141;
wire v_9142;
wire v_9143;
wire v_9144;
wire v_9145;
wire v_9146;
wire v_9147;
wire v_9148;
wire v_9149;
wire v_9150;
wire v_9151;
wire v_9152;
wire v_9153;
wire v_9154;
wire v_9155;
wire v_9156;
wire v_9157;
wire v_9158;
wire v_9159;
wire v_9160;
wire v_9163;
wire v_9164;
wire v_9165;
wire v_9166;
wire v_9167;
wire v_9168;
wire v_9169;
wire v_9170;
wire v_9171;
wire v_9172;
wire v_9174;
wire v_9176;
wire v_9177;
wire v_9178;
wire v_9179;
wire v_9180;
wire v_9181;
wire v_9182;
wire v_9183;
wire v_9184;
wire v_9185;
wire v_9186;
wire v_9187;
wire v_9188;
wire v_9189;
wire v_9190;
wire v_9191;
wire v_9192;
wire v_9193;
wire v_9194;
wire v_9195;
wire v_9196;
wire v_9197;
wire v_9198;
wire v_9199;
wire v_9200;
wire v_9201;
wire v_9202;
wire v_9203;
wire v_9204;
wire v_9207;
wire v_9208;
wire v_9209;
wire v_9210;
wire v_9211;
wire v_9212;
wire v_9213;
wire v_9214;
wire v_9215;
wire v_9216;
wire v_9219;
wire v_9220;
wire v_9221;
wire v_9222;
wire v_9223;
wire v_9224;
wire v_9225;
wire v_9226;
wire v_9227;
wire v_9228;
wire v_9231;
wire v_9232;
wire v_9233;
wire v_9234;
wire v_9235;
wire v_9236;
wire v_9237;
wire v_9238;
wire v_9239;
wire v_9240;
wire v_9243;
wire v_9244;
wire v_9245;
wire v_9246;
wire v_9247;
wire v_9248;
wire v_9249;
wire v_9250;
wire v_9251;
wire v_9252;
wire v_9255;
wire v_9256;
wire v_9257;
wire v_9258;
wire v_9259;
wire v_9260;
wire v_9261;
wire v_9262;
wire v_9263;
wire v_9264;
wire v_9267;
wire v_9268;
wire v_9269;
wire v_9270;
wire v_9271;
wire v_9272;
wire v_9273;
wire v_9274;
wire v_9275;
wire v_9276;
wire v_9277;
wire v_9278;
wire v_9279;
wire v_9280;
wire v_9281;
wire v_9282;
wire v_9283;
wire v_9284;
wire v_9285;
wire v_9286;
wire v_9287;
wire v_9288;
wire v_9289;
wire v_9290;
wire v_9291;
wire v_9292;
wire v_9295;
wire v_9296;
wire v_9297;
wire v_9298;
wire v_9299;
wire v_9300;
wire v_9301;
wire v_9302;
wire v_9303;
wire v_9304;
wire v_9306;
wire v_9307;
wire v_9308;
wire v_9309;
wire v_9310;
wire v_9312;
wire v_9313;
wire v_9314;
wire v_9315;
wire v_9316;
wire v_9317;
wire v_9318;
wire v_9319;
wire v_9320;
wire v_9321;
wire v_9322;
wire v_9323;
wire v_9324;
wire v_9325;
wire v_9326;
wire v_9327;
wire v_9328;
wire v_9329;
wire v_9330;
wire v_9331;
wire v_9332;
wire v_9333;
wire v_9334;
wire v_9335;
wire v_9336;
wire v_9337;
wire v_9338;
wire v_9339;
wire v_9340;
wire v_9341;
wire v_9342;
wire v_9343;
wire v_9344;
wire v_9345;
wire v_9346;
wire v_9347;
wire v_9348;
wire v_9349;
wire v_9350;
wire v_9351;
wire v_9352;
wire v_9353;
wire v_9354;
wire v_9355;
wire v_9356;
wire v_9357;
wire v_9358;
wire v_9359;
wire v_9360;
wire v_9363;
wire v_9364;
wire v_9365;
wire v_9366;
wire v_9367;
wire v_9368;
wire v_9369;
wire v_9370;
wire v_9371;
wire v_9372;
wire v_9375;
wire v_9376;
wire v_9377;
wire v_9378;
wire v_9379;
wire v_9380;
wire v_9381;
wire v_9382;
wire v_9383;
wire v_9384;
wire v_9387;
wire v_9388;
wire v_9389;
wire v_9390;
wire v_9391;
wire v_9392;
wire v_9393;
wire v_9394;
wire v_9395;
wire v_9396;
wire v_9399;
wire v_9400;
wire v_9401;
wire v_9402;
wire v_9403;
wire v_9404;
wire v_9405;
wire v_9406;
wire v_9407;
wire v_9408;
wire v_9411;
wire v_9412;
wire v_9413;
wire v_9414;
wire v_9415;
wire v_9416;
wire v_9417;
wire v_9418;
wire v_9419;
wire v_9420;
wire v_9423;
wire v_9424;
wire v_9425;
wire v_9426;
wire v_9427;
wire v_9428;
wire v_9429;
wire v_9430;
wire v_9431;
wire v_9432;
wire v_9433;
wire v_9434;
wire v_9435;
wire v_9436;
wire v_9437;
wire v_9438;
wire v_9439;
wire v_9440;
wire v_9441;
wire v_9442;
wire v_9443;
wire v_9444;
wire v_9445;
wire v_9446;
wire v_9447;
wire v_9448;
wire v_9451;
wire v_9452;
wire v_9453;
wire v_9454;
wire v_9455;
wire v_9456;
wire v_9457;
wire v_9458;
wire v_9459;
wire v_9460;
wire v_9462;
wire v_9464;
wire v_9465;
wire v_9466;
wire v_9467;
wire v_9468;
wire v_9469;
wire v_9470;
wire v_9471;
wire v_9472;
wire v_9473;
wire v_9474;
wire v_9475;
wire v_9476;
wire v_9477;
wire v_9478;
wire v_9479;
wire v_9480;
wire v_9481;
wire v_9482;
wire v_9483;
wire v_9484;
wire v_9485;
wire v_9486;
wire v_9487;
wire v_9488;
wire v_9489;
wire v_9490;
wire v_9491;
wire v_9492;
wire v_9495;
wire v_9496;
wire v_9497;
wire v_9498;
wire v_9499;
wire v_9500;
wire v_9501;
wire v_9502;
wire v_9503;
wire v_9504;
wire v_9507;
wire v_9508;
wire v_9509;
wire v_9510;
wire v_9511;
wire v_9512;
wire v_9513;
wire v_9514;
wire v_9515;
wire v_9516;
wire v_9519;
wire v_9520;
wire v_9521;
wire v_9522;
wire v_9523;
wire v_9524;
wire v_9525;
wire v_9526;
wire v_9527;
wire v_9528;
wire v_9531;
wire v_9532;
wire v_9533;
wire v_9534;
wire v_9535;
wire v_9536;
wire v_9537;
wire v_9538;
wire v_9539;
wire v_9540;
wire v_9543;
wire v_9544;
wire v_9545;
wire v_9546;
wire v_9547;
wire v_9548;
wire v_9549;
wire v_9550;
wire v_9551;
wire v_9552;
wire v_9555;
wire v_9556;
wire v_9557;
wire v_9558;
wire v_9559;
wire v_9560;
wire v_9561;
wire v_9562;
wire v_9563;
wire v_9564;
wire v_9565;
wire v_9566;
wire v_9567;
wire v_9568;
wire v_9569;
wire v_9570;
wire v_9571;
wire v_9572;
wire v_9573;
wire v_9574;
wire v_9575;
wire v_9576;
wire v_9577;
wire v_9578;
wire v_9579;
wire v_9580;
wire v_9583;
wire v_9584;
wire v_9585;
wire v_9586;
wire v_9587;
wire v_9588;
wire v_9589;
wire v_9590;
wire v_9591;
wire v_9592;
wire v_9594;
wire v_9595;
wire v_9596;
wire v_9597;
wire v_9598;
wire v_9599;
wire v_9600;
wire v_9601;
wire v_9602;
wire v_9603;
wire v_9605;
wire v_9606;
wire v_9607;
wire v_9608;
wire v_9609;
wire v_9610;
wire v_9611;
wire v_9612;
wire v_9613;
wire v_9614;
wire v_9615;
wire v_9616;
wire v_9617;
wire v_9618;
wire v_9619;
wire v_9620;
wire v_9621;
wire v_9622;
wire v_9623;
wire v_9624;
wire v_9625;
wire v_9626;
wire v_9627;
wire v_9628;
wire v_9629;
wire v_9630;
wire v_9631;
wire v_9632;
wire v_9633;
wire v_9634;
wire v_9635;
wire v_9636;
wire v_9637;
wire v_9638;
wire v_9639;
wire v_9640;
wire v_9641;
wire v_9642;
wire v_9643;
wire v_9644;
wire v_9645;
wire v_9646;
wire v_9647;
wire v_9648;
wire v_9649;
wire v_9650;
wire v_9653;
wire v_9654;
wire v_9655;
wire v_9656;
wire v_9657;
wire v_9658;
wire v_9659;
wire v_9660;
wire v_9661;
wire v_9662;
wire v_9665;
wire v_9666;
wire v_9667;
wire v_9668;
wire v_9669;
wire v_9670;
wire v_9671;
wire v_9672;
wire v_9673;
wire v_9674;
wire v_9677;
wire v_9678;
wire v_9679;
wire v_9680;
wire v_9681;
wire v_9682;
wire v_9683;
wire v_9684;
wire v_9685;
wire v_9686;
wire v_9689;
wire v_9690;
wire v_9691;
wire v_9692;
wire v_9693;
wire v_9694;
wire v_9695;
wire v_9696;
wire v_9697;
wire v_9698;
wire v_9701;
wire v_9702;
wire v_9703;
wire v_9704;
wire v_9705;
wire v_9706;
wire v_9707;
wire v_9708;
wire v_9709;
wire v_9710;
wire v_9713;
wire v_9714;
wire v_9715;
wire v_9716;
wire v_9717;
wire v_9718;
wire v_9719;
wire v_9720;
wire v_9721;
wire v_9722;
wire v_9723;
wire v_9724;
wire v_9725;
wire v_9726;
wire v_9727;
wire v_9728;
wire v_9729;
wire v_9730;
wire v_9731;
wire v_9732;
wire v_9733;
wire v_9734;
wire v_9735;
wire v_9736;
wire v_9737;
wire v_9738;
wire v_9741;
wire v_9742;
wire v_9743;
wire v_9744;
wire v_9745;
wire v_9746;
wire v_9747;
wire v_9748;
wire v_9749;
wire v_9750;
wire v_9752;
wire v_9754;
wire v_9755;
wire v_9756;
wire v_9757;
wire v_9758;
wire v_9759;
wire v_9760;
wire v_9761;
wire v_9762;
wire v_9763;
wire v_9764;
wire v_9765;
wire v_9766;
wire v_9767;
wire v_9768;
wire v_9769;
wire v_9770;
wire v_9771;
wire v_9772;
wire v_9773;
wire v_9774;
wire v_9775;
wire v_9776;
wire v_9777;
wire v_9778;
wire v_9779;
wire v_9780;
wire v_9781;
wire v_9782;
wire v_9785;
wire v_9786;
wire v_9787;
wire v_9788;
wire v_9789;
wire v_9790;
wire v_9791;
wire v_9792;
wire v_9793;
wire v_9794;
wire v_9797;
wire v_9798;
wire v_9799;
wire v_9800;
wire v_9801;
wire v_9802;
wire v_9803;
wire v_9804;
wire v_9805;
wire v_9806;
wire v_9809;
wire v_9810;
wire v_9811;
wire v_9812;
wire v_9813;
wire v_9814;
wire v_9815;
wire v_9816;
wire v_9817;
wire v_9818;
wire v_9821;
wire v_9822;
wire v_9823;
wire v_9824;
wire v_9825;
wire v_9826;
wire v_9827;
wire v_9828;
wire v_9829;
wire v_9830;
wire v_9833;
wire v_9834;
wire v_9835;
wire v_9836;
wire v_9837;
wire v_9838;
wire v_9839;
wire v_9840;
wire v_9841;
wire v_9842;
wire v_9845;
wire v_9846;
wire v_9847;
wire v_9848;
wire v_9849;
wire v_9850;
wire v_9851;
wire v_9852;
wire v_9853;
wire v_9854;
wire v_9855;
wire v_9856;
wire v_9857;
wire v_9858;
wire v_9859;
wire v_9860;
wire v_9861;
wire v_9862;
wire v_9863;
wire v_9864;
wire v_9865;
wire v_9866;
wire v_9867;
wire v_9868;
wire v_9869;
wire v_9870;
wire v_9873;
wire v_9874;
wire v_9875;
wire v_9876;
wire v_9877;
wire v_9878;
wire v_9879;
wire v_9880;
wire v_9881;
wire v_9882;
wire v_9885;
wire v_9886;
wire v_9887;
wire v_9888;
wire v_9889;
wire v_9890;
wire v_9891;
wire v_9892;
wire v_9893;
wire v_9894;
wire v_9895;
wire v_9896;
wire v_9897;
wire v_9898;
wire v_9899;
wire v_9900;
wire v_9901;
wire v_9902;
wire v_9904;
wire v_9905;
wire v_9906;
wire v_9907;
wire v_9908;
wire v_9909;
wire v_9910;
wire v_9911;
wire v_9912;
wire v_9913;
wire v_9914;
wire v_9915;
wire v_9916;
wire v_9917;
wire v_9918;
wire v_9919;
wire v_9920;
wire v_9921;
wire v_9922;
wire v_9923;
wire v_9924;
wire v_9925;
wire v_9926;
wire v_9927;
wire v_9928;
wire v_9929;
wire v_9930;
wire v_9931;
wire v_9932;
wire v_9933;
wire v_9934;
wire v_9935;
wire v_9936;
wire v_9937;
wire v_9938;
wire v_9939;
wire v_9940;
wire v_9941;
wire v_9942;
wire v_9943;
wire v_9944;
wire v_9945;
wire v_9946;
wire v_9947;
wire v_9949;
wire v_9950;
wire v_9951;
wire v_9952;
wire v_9953;
wire v_9954;
wire v_9955;
wire v_9956;
wire v_9957;
wire v_9958;
wire v_9959;
wire v_9960;
wire v_9961;
wire v_9962;
wire v_9963;
wire v_9964;
wire v_9965;
wire v_9966;
wire v_9967;
wire v_9968;
wire v_9969;
wire v_9970;
wire v_9971;
wire v_9972;
wire v_9973;
wire v_9974;
wire v_9975;
wire v_9976;
wire v_9977;
wire v_9978;
wire v_9979;
wire v_9980;
wire v_9981;
wire v_9982;
wire v_9983;
wire v_9984;
wire v_9986;
wire v_9987;
wire v_9988;
wire v_9989;
wire v_9990;
wire v_9991;
wire v_9992;
wire v_9993;
wire v_9994;
wire v_9995;
wire v_9996;
wire v_9997;
wire v_9998;
wire v_9999;
wire v_10000;
wire v_10001;
wire v_10002;
wire v_10003;
wire v_10004;
wire v_10005;
wire v_10006;
wire v_10007;
wire v_10008;
wire v_10009;
wire v_10010;
wire v_10011;
wire v_10012;
wire v_10013;
wire v_10014;
wire v_10015;
wire v_10016;
wire v_10017;
wire v_10018;
wire v_10019;
wire v_10020;
wire v_10021;
wire v_10023;
wire v_10024;
wire v_10025;
wire v_10026;
wire v_10027;
wire v_10028;
wire v_10029;
wire v_10030;
wire v_10031;
wire v_10032;
wire v_10033;
wire v_10034;
wire v_10035;
wire v_10036;
wire v_10037;
wire v_10038;
wire v_10039;
wire v_10040;
wire v_10041;
wire v_10042;
wire v_10043;
wire v_10044;
wire v_10045;
wire v_10046;
wire v_10047;
wire v_10048;
wire v_10049;
wire v_10050;
wire v_10051;
wire v_10052;
wire v_10053;
wire v_10054;
wire v_10055;
wire v_10056;
wire v_10057;
wire v_10058;
wire v_10060;
wire v_10061;
wire v_10062;
wire v_10063;
wire v_10064;
wire v_10065;
wire v_10066;
wire v_10067;
wire v_10068;
wire v_10069;
wire v_10070;
wire v_10071;
wire v_10072;
wire v_10073;
wire v_10074;
wire v_10075;
wire v_10076;
wire v_10077;
wire v_10078;
wire v_10079;
wire v_10080;
wire v_10081;
wire v_10082;
wire v_10083;
wire v_10084;
wire v_10085;
wire v_10086;
wire v_10087;
wire v_10088;
wire v_10089;
wire v_10090;
wire v_10091;
wire v_10092;
wire v_10093;
wire v_10094;
wire v_10095;
wire v_10097;
wire v_10098;
wire v_10099;
wire v_10100;
wire v_10101;
wire v_10102;
wire v_10103;
wire v_10104;
wire v_10105;
wire v_10106;
wire v_10107;
wire v_10108;
wire v_10109;
wire v_10110;
wire v_10111;
wire v_10112;
wire v_10113;
wire v_10114;
wire v_10115;
wire v_10116;
wire v_10117;
wire v_10118;
wire v_10119;
wire v_10120;
wire v_10121;
wire v_10122;
wire v_10123;
wire v_10124;
wire v_10125;
wire v_10126;
wire v_10127;
wire v_10128;
wire v_10129;
wire v_10130;
wire v_10131;
wire v_10132;
wire v_10134;
wire v_10135;
wire v_10136;
wire v_10137;
wire v_10138;
wire v_10139;
wire v_10140;
wire v_10141;
wire v_10142;
wire v_10143;
wire v_10144;
wire v_10145;
wire v_10146;
wire v_10147;
wire v_10148;
wire v_10149;
wire v_10150;
wire v_10151;
wire v_10152;
wire v_10153;
wire v_10154;
wire v_10155;
wire v_10156;
wire v_10157;
wire v_10158;
wire v_10159;
wire v_10160;
wire v_10161;
wire v_10162;
wire v_10163;
wire v_10164;
wire v_10165;
wire v_10166;
wire v_10167;
wire v_10169;
wire v_10170;
wire v_10171;
wire v_10172;
wire v_10173;
wire v_10174;
wire v_10175;
wire v_10176;
wire v_10177;
wire v_10178;
wire v_10179;
wire v_10180;
wire v_10181;
wire v_10182;
wire v_10183;
wire v_10184;
wire v_10185;
wire v_10186;
wire v_10187;
wire v_10188;
wire v_10189;
wire v_10190;
wire v_10191;
wire v_10192;
wire v_10193;
wire v_10194;
wire v_10197;
wire v_10198;
wire v_10199;
wire v_10201;
wire v_10202;
wire v_10203;
wire v_10204;
wire v_10205;
wire v_10206;
wire v_10207;
wire v_10208;
wire v_10209;
wire v_10210;
wire v_10211;
wire v_10212;
wire v_10213;
wire v_10214;
wire v_10215;
wire v_10216;
wire v_10217;
wire v_10218;
wire v_10219;
wire v_10220;
wire v_10221;
wire v_10222;
wire v_10223;
wire v_10225;
wire v_10226;
wire v_10227;
wire v_10228;
wire v_10229;
wire v_10230;
wire v_10231;
wire v_10232;
wire v_10233;
wire v_10234;
wire v_10235;
wire v_10236;
wire v_10237;
wire v_10238;
wire v_10239;
wire v_10240;
wire v_10241;
wire v_10242;
wire v_10243;
wire v_10244;
wire v_10245;
wire v_10246;
wire v_10247;
wire v_10248;
wire v_10249;
wire v_10250;
wire v_10252;
wire v_10253;
wire v_10254;
wire v_10255;
wire v_10256;
wire v_10257;
wire v_10258;
wire v_10259;
wire v_10260;
wire v_10261;
wire v_10262;
wire v_10263;
wire v_10264;
wire v_10265;
wire v_10266;
wire v_10267;
wire v_10268;
wire v_10269;
wire v_10270;
wire v_10271;
wire v_10272;
wire v_10273;
wire v_10274;
wire v_10275;
wire v_10276;
wire v_10277;
wire v_10279;
wire v_10280;
wire v_10281;
wire v_10282;
wire v_10283;
wire v_10284;
wire v_10285;
wire v_10286;
wire v_10287;
wire v_10288;
wire v_10289;
wire v_10290;
wire v_10291;
wire v_10292;
wire v_10293;
wire v_10294;
wire v_10295;
wire v_10296;
wire v_10297;
wire v_10298;
wire v_10299;
wire v_10300;
wire v_10301;
wire v_10302;
wire v_10303;
wire v_10304;
wire v_10306;
wire v_10307;
wire v_10308;
wire v_10309;
wire v_10310;
wire v_10311;
wire v_10312;
wire v_10313;
wire v_10314;
wire v_10315;
wire v_10316;
wire v_10317;
wire v_10318;
wire v_10319;
wire v_10320;
wire v_10321;
wire v_10322;
wire v_10323;
wire v_10324;
wire v_10325;
wire v_10326;
wire v_10327;
wire v_10328;
wire v_10329;
wire v_10330;
wire v_10331;
wire v_10333;
wire v_10334;
wire v_10335;
wire v_10336;
wire v_10337;
wire v_10338;
wire v_10339;
wire v_10340;
wire v_10341;
wire v_10342;
wire v_10343;
wire v_10344;
wire v_10345;
wire v_10346;
wire v_10347;
wire v_10348;
wire v_10349;
wire v_10350;
wire v_10351;
wire v_10352;
wire v_10353;
wire v_10354;
wire v_10355;
wire v_10356;
wire v_10357;
wire v_10358;
wire v_10360;
wire v_10361;
wire v_10362;
wire v_10363;
wire v_10364;
wire v_10365;
wire v_10366;
wire v_10367;
wire v_10368;
wire v_10369;
wire v_10370;
wire v_10371;
wire v_10372;
wire v_10373;
wire v_10374;
wire v_10375;
wire v_10376;
wire v_10377;
wire v_10378;
wire v_10379;
wire v_10380;
wire v_10381;
wire v_10382;
wire v_10383;
wire v_10384;
wire v_10385;
wire v_10387;
wire v_10388;
wire v_10389;
wire v_10390;
wire v_10391;
wire v_10392;
wire v_10393;
wire v_10394;
wire v_10395;
wire v_10396;
wire v_10397;
wire v_10398;
wire v_10399;
wire v_10400;
wire v_10401;
wire v_10402;
wire v_10403;
wire v_10404;
wire v_10405;
wire v_10406;
wire v_10407;
wire v_10408;
wire v_10409;
wire v_10410;
wire v_10411;
wire v_10412;
wire v_10416;
wire v_10417;
wire v_10418;
wire v_10419;
wire v_10422;
wire v_10423;
wire v_10424;
wire v_10425;
wire v_10428;
wire v_10429;
wire v_10430;
wire v_10431;
wire v_10434;
wire v_10435;
wire v_10436;
wire v_10437;
wire v_10440;
wire v_10441;
wire v_10442;
wire v_10443;
wire v_10446;
wire v_10447;
wire v_10448;
wire v_10449;
wire v_10452;
wire v_10453;
wire v_10454;
wire v_10455;
wire v_10457;
wire v_10458;
wire v_10459;
wire v_10460;
wire v_10463;
wire v_10464;
wire v_10466;
wire v_10467;
wire v_10468;
wire v_10469;
wire v_10470;
wire v_10471;
wire v_10472;
wire v_10473;
wire v_10474;
wire v_10475;
wire v_10476;
wire v_10477;
wire v_10478;
wire v_10479;
wire v_10480;
wire v_10481;
wire v_10482;
wire v_10483;
wire v_10484;
wire v_10485;
wire v_10486;
wire v_10487;
wire v_10488;
wire v_10489;
wire v_10490;
wire v_10491;
wire v_10492;
wire v_10493;
wire v_10494;
wire v_10495;
wire v_10496;
wire v_10497;
wire v_10498;
wire v_10499;
wire v_10500;
wire v_10501;
wire v_10502;
wire v_10503;
wire v_10504;
wire v_10505;
wire v_10506;
wire v_10507;
wire v_10508;
wire v_10509;
wire v_10510;
wire v_10511;
wire v_10512;
wire v_10513;
wire v_10514;
wire v_10515;
wire v_10516;
wire v_10517;
wire v_10518;
wire v_10519;
wire v_10520;
wire v_10521;
wire v_10522;
wire v_10523;
wire v_10524;
wire v_10525;
wire v_10526;
wire v_10527;
wire v_10528;
wire v_10529;
wire v_10530;
wire v_10531;
wire v_10532;
wire v_10533;
wire v_10534;
wire v_10535;
wire v_10536;
wire v_10537;
wire v_10538;
wire v_10539;
wire v_10540;
wire v_10541;
wire v_10542;
wire v_10543;
wire v_10544;
wire v_10545;
wire v_10546;
wire v_10547;
wire v_10548;
wire v_10549;
wire v_10550;
wire v_10551;
wire v_10552;
wire v_10553;
wire v_10554;
wire v_10555;
wire v_10556;
wire v_10557;
wire v_10558;
wire v_10559;
wire v_10560;
wire v_10561;
wire v_10562;
wire v_10563;
wire v_10564;
wire v_10565;
wire v_10566;
wire v_10567;
wire v_10568;
wire v_10569;
wire v_10570;
wire v_10571;
wire v_10572;
wire v_10573;
wire v_10574;
wire v_10575;
wire v_10576;
wire v_10577;
wire v_10578;
wire v_10579;
wire v_10580;
wire v_10581;
wire v_10582;
wire v_10583;
wire v_10584;
wire v_10585;
wire v_10586;
wire v_10587;
wire v_10588;
wire v_10589;
wire v_10590;
wire v_10591;
wire v_10592;
wire v_10593;
wire v_10594;
wire v_10595;
wire v_10596;
wire v_10597;
wire v_10598;
wire v_10599;
wire v_10600;
wire v_10601;
wire v_10602;
wire v_10603;
wire v_10604;
wire v_10605;
wire v_10606;
wire v_10607;
wire v_10608;
wire v_10609;
wire v_10610;
wire v_10611;
wire v_10612;
wire v_10613;
wire v_10614;
wire v_10615;
wire v_10616;
wire v_10617;
wire v_10618;
wire v_10619;
wire v_10620;
wire v_10621;
wire v_10622;
wire v_10623;
wire v_10624;
wire v_10625;
wire v_10626;
wire v_10627;
wire v_10628;
wire v_10629;
wire v_10630;
wire v_10631;
wire v_10632;
wire v_10633;
wire v_10634;
wire v_10635;
wire v_10636;
wire v_10637;
wire v_10638;
wire v_10639;
wire v_10640;
wire v_10641;
wire v_10642;
wire v_10643;
wire v_10644;
wire v_10645;
wire v_10646;
wire v_10647;
wire v_10648;
wire v_10649;
wire v_10650;
wire v_10651;
wire v_10652;
wire v_10653;
wire v_10654;
wire v_10655;
wire v_10656;
wire v_10657;
wire v_10658;
wire v_10659;
wire v_10660;
wire v_10661;
wire v_10662;
wire v_10663;
wire v_10664;
wire v_10665;
wire v_10666;
wire v_10667;
wire v_10668;
wire v_10669;
wire v_10670;
wire v_10671;
wire v_10672;
wire v_10673;
wire v_10674;
wire v_10675;
wire v_10676;
wire v_10677;
wire v_10678;
wire v_10679;
wire v_10680;
wire v_10681;
wire v_10682;
wire v_10683;
wire v_10684;
wire v_10685;
wire v_10686;
wire v_10687;
wire v_10688;
wire v_10689;
wire v_10690;
wire v_10691;
wire v_10692;
wire v_10693;
wire v_10694;
wire v_10695;
wire v_10696;
wire v_10697;
wire v_10698;
wire v_10699;
wire v_10700;
wire v_10701;
wire v_10702;
wire v_10703;
wire v_10704;
wire v_10705;
wire v_10706;
wire v_10707;
wire v_10708;
wire v_10709;
wire v_10710;
wire v_10711;
wire v_10712;
wire v_10713;
wire v_10714;
wire v_10715;
wire v_10716;
wire v_10717;
wire v_10718;
wire v_10719;
wire v_10720;
wire v_10721;
wire v_10722;
wire v_10723;
wire v_10724;
wire v_10725;
wire v_10726;
wire v_10727;
wire v_10728;
wire v_10729;
wire v_10730;
wire v_10731;
wire v_10732;
wire v_10733;
wire v_10734;
wire v_10735;
wire v_10736;
wire v_10737;
wire v_10738;
wire v_10739;
wire v_10740;
wire v_10741;
wire v_10742;
wire v_10743;
wire v_10744;
wire v_10745;
wire v_10746;
wire v_10747;
wire v_10748;
wire v_10749;
wire v_10750;
wire v_10751;
wire v_10752;
wire v_10753;
wire v_10754;
wire v_10755;
wire v_10756;
wire v_10757;
wire v_10758;
wire v_10759;
wire v_10760;
wire v_10761;
wire v_10762;
wire v_10763;
wire v_10764;
wire v_10765;
wire v_10766;
wire v_10767;
wire v_10768;
wire v_10769;
wire v_10770;
wire v_10771;
wire v_10772;
wire v_10773;
wire v_10774;
wire v_10775;
wire v_10776;
wire v_10777;
wire v_10778;
wire v_10779;
wire v_10780;
wire v_10781;
wire v_10782;
wire v_10783;
wire v_10784;
wire v_10785;
wire v_10786;
wire v_10787;
wire v_10788;
wire v_10789;
wire v_10790;
wire v_10791;
wire v_10792;
wire v_10793;
wire v_10794;
wire v_10795;
wire v_10796;
wire v_10797;
wire v_10798;
wire v_10799;
wire v_10800;
wire v_10801;
wire v_10802;
wire v_10803;
wire v_10804;
wire v_10805;
wire v_10806;
wire v_10807;
wire v_10808;
wire v_10809;
wire v_10810;
wire v_10811;
wire v_10812;
wire v_10813;
wire v_10814;
wire v_10815;
wire v_10816;
wire v_10817;
wire v_10818;
wire v_10819;
wire v_10820;
wire v_10821;
wire v_10822;
wire v_10823;
wire v_10824;
wire v_10825;
wire v_10826;
wire v_10827;
wire v_10828;
wire v_10829;
wire v_10830;
wire v_10831;
wire v_10832;
wire v_10833;
wire v_10834;
wire v_10835;
wire v_10836;
wire v_10837;
wire v_10838;
wire v_10839;
wire v_10840;
wire v_10841;
wire v_10842;
wire v_10843;
wire v_10844;
wire v_10845;
wire v_10846;
wire v_10847;
wire v_10848;
wire v_10849;
wire v_10850;
wire v_10851;
wire v_10852;
wire v_10853;
wire v_10854;
wire v_10855;
wire v_10856;
wire v_10857;
wire v_10858;
wire v_10859;
wire v_10860;
wire v_10861;
wire v_10862;
wire v_10863;
wire v_10864;
wire v_10865;
wire v_10866;
wire v_10867;
wire v_10868;
wire v_10869;
wire v_10870;
wire v_10871;
wire v_10872;
wire v_10873;
wire v_10874;
wire v_10875;
wire v_10876;
wire v_10877;
wire v_10878;
wire v_10879;
wire v_10880;
wire v_10881;
wire v_10882;
wire v_10883;
wire v_10884;
wire v_10885;
wire v_10886;
wire v_10887;
wire v_10888;
wire v_10889;
wire v_10890;
wire v_10891;
wire v_10892;
wire v_10893;
wire v_10894;
wire v_10895;
wire v_10896;
wire v_10897;
wire v_10898;
wire v_10899;
wire v_10900;
wire v_10901;
wire v_10902;
wire v_10903;
wire v_10904;
wire v_10905;
wire v_10906;
wire v_10907;
wire v_10908;
wire v_10909;
wire v_10910;
wire v_10911;
wire v_10912;
wire v_10913;
wire v_10914;
wire v_10915;
wire v_10916;
wire v_10917;
wire v_10918;
wire v_10919;
wire v_10920;
wire v_10921;
wire v_10922;
wire v_10923;
wire v_10924;
wire v_10925;
wire v_10926;
wire v_10927;
wire v_10928;
wire v_10929;
wire v_10930;
wire v_10931;
wire v_10932;
wire v_10933;
wire v_10934;
wire v_10935;
wire v_10936;
wire v_10937;
wire v_10938;
wire v_10939;
wire v_10940;
wire v_10941;
wire v_10942;
wire v_10943;
wire v_10944;
wire v_10945;
wire v_10946;
wire v_10947;
wire v_10948;
wire v_10949;
wire v_10950;
wire v_10951;
wire v_10952;
wire v_10953;
wire v_10954;
wire v_10955;
wire v_10956;
wire v_10957;
wire v_10958;
wire v_10959;
wire v_10960;
wire v_10961;
wire v_10962;
wire v_10963;
wire v_10964;
wire v_10965;
wire v_10966;
wire v_10967;
wire v_10968;
wire v_10969;
wire v_10970;
wire v_10971;
wire v_10972;
wire v_10973;
wire v_10974;
wire v_10975;
wire v_10976;
wire v_10977;
wire v_10978;
wire v_10979;
wire v_10980;
wire v_10981;
wire v_10982;
wire v_10983;
wire v_10984;
wire v_10985;
wire v_10986;
wire v_10987;
wire v_10988;
wire v_10989;
wire v_10990;
wire v_10991;
wire v_10992;
wire v_10993;
wire v_10994;
wire v_10995;
wire v_10996;
wire v_10997;
wire v_10998;
wire v_10999;
wire v_11000;
wire v_11001;
wire v_11002;
wire v_11003;
wire v_11004;
wire v_11005;
wire v_11006;
wire v_11007;
wire v_11008;
wire v_11009;
wire v_11010;
wire v_11011;
wire v_11012;
wire v_11013;
wire v_11014;
wire v_11015;
wire v_11016;
wire v_11017;
wire v_11018;
wire v_11019;
wire v_11020;
wire v_11021;
wire v_11022;
wire v_11023;
wire v_11024;
wire v_11025;
wire v_11026;
wire v_11027;
wire v_11028;
wire v_11029;
wire v_11030;
wire v_11031;
wire v_11032;
wire v_11033;
wire v_11034;
wire v_11035;
wire v_11036;
wire v_11037;
wire v_11038;
wire v_11039;
wire v_11040;
wire v_11041;
wire v_11042;
wire v_11043;
wire v_11044;
wire v_11045;
wire v_11046;
wire v_11047;
wire v_11048;
wire v_11049;
wire v_11050;
wire v_11051;
wire v_11052;
wire v_11053;
wire v_11054;
wire v_11055;
wire v_11056;
wire v_11057;
wire v_11058;
wire v_11059;
wire v_11060;
wire v_11061;
wire v_11062;
wire v_11063;
wire v_11064;
wire v_11065;
wire v_11066;
wire v_11067;
wire v_11068;
wire v_11069;
wire v_11070;
wire v_11071;
wire v_11072;
wire v_11073;
wire v_11074;
wire v_11075;
wire v_11076;
wire v_11077;
wire v_11078;
wire v_11079;
wire v_11080;
wire v_11081;
wire v_11082;
wire v_11083;
wire v_11084;
wire v_11085;
wire v_11086;
wire v_11087;
wire v_11088;
wire v_11089;
wire v_11090;
wire v_11091;
wire v_11092;
wire v_11093;
wire v_11094;
wire v_11095;
wire v_11096;
wire v_11097;
wire v_11098;
wire v_11099;
wire v_11100;
wire v_11101;
wire v_11102;
wire v_11103;
wire v_11104;
wire v_11105;
wire v_11106;
wire v_11107;
wire v_11108;
wire v_11109;
wire v_11110;
wire v_11111;
wire v_11112;
wire v_11113;
wire v_11114;
wire v_11115;
wire v_11116;
wire v_11117;
wire v_11118;
wire v_11119;
wire v_11120;
wire v_11121;
wire v_11122;
wire v_11123;
wire v_11124;
wire v_11125;
wire v_11126;
wire v_11127;
wire v_11128;
wire v_11129;
wire v_11130;
wire v_11131;
wire v_11132;
wire v_11133;
wire v_11134;
wire v_11135;
wire v_11136;
wire v_11137;
wire v_11138;
wire v_11139;
wire v_11140;
wire v_11141;
wire v_11142;
wire v_11143;
wire v_11144;
wire v_11145;
wire v_11146;
wire v_11147;
wire v_11148;
wire v_11149;
wire v_11150;
wire v_11151;
wire v_11152;
wire v_11153;
wire v_11154;
wire v_11155;
wire v_11156;
wire v_11157;
wire v_11158;
wire v_11159;
wire v_11160;
wire v_11161;
wire v_11162;
wire v_11163;
wire v_11164;
wire v_11165;
wire v_11166;
wire v_11167;
wire v_11168;
wire v_11169;
wire v_11170;
wire v_11171;
wire v_11172;
wire v_11173;
wire v_11174;
wire v_11175;
wire v_11176;
wire v_11177;
wire v_11178;
wire v_11179;
wire v_11180;
wire v_11181;
wire v_11182;
wire v_11183;
wire v_11184;
wire v_11185;
wire v_11186;
wire v_11187;
wire v_11188;
wire v_11189;
wire v_11190;
wire v_11191;
wire v_11192;
wire v_11193;
wire v_11194;
wire v_11195;
wire v_11196;
wire v_11197;
wire v_11198;
wire v_11199;
wire v_11200;
wire v_11201;
wire v_11202;
wire v_11203;
wire v_11204;
wire v_11205;
wire v_11206;
wire v_11207;
wire v_11208;
wire v_11209;
wire v_11210;
wire v_11211;
wire v_11212;
wire v_11213;
wire v_11214;
wire v_11215;
wire v_11216;
wire v_11217;
wire v_11218;
wire v_11219;
wire v_11220;
wire v_11221;
wire v_11222;
wire v_11223;
wire v_11224;
wire v_11225;
wire v_11226;
wire v_11227;
wire v_11228;
wire v_11229;
wire v_11230;
wire v_11231;
wire v_11232;
wire v_11233;
wire v_11234;
wire v_11235;
wire v_11236;
wire v_11237;
wire v_11238;
wire v_11239;
wire v_11240;
wire v_11241;
wire v_11242;
wire v_11243;
wire v_11244;
wire v_11245;
wire v_11246;
wire v_11247;
wire v_11248;
wire v_11249;
wire v_11250;
wire v_11251;
wire v_11252;
wire v_11253;
wire v_11254;
wire v_11255;
wire v_11256;
wire v_11257;
wire v_11258;
wire v_11259;
wire v_11260;
wire v_11261;
wire v_11262;
wire v_11263;
wire v_11264;
wire v_11265;
wire v_11266;
wire v_11267;
wire v_11268;
wire v_11269;
wire v_11270;
wire v_11271;
wire v_11272;
wire v_11273;
wire v_11274;
wire v_11275;
wire v_11276;
wire v_11277;
wire v_11278;
wire v_11279;
wire v_11280;
wire v_11281;
wire v_11282;
wire v_11283;
wire v_11284;
wire v_11285;
wire v_11286;
wire v_11287;
wire v_11288;
wire v_11289;
wire v_11290;
wire v_11291;
wire v_11292;
wire v_11293;
wire v_11294;
wire v_11295;
wire v_11296;
wire v_11297;
wire v_11298;
wire v_11299;
wire v_11300;
wire v_11301;
wire v_11302;
wire v_11303;
wire v_11304;
wire v_11305;
wire v_11306;
wire v_11307;
wire v_11308;
wire v_11309;
wire v_11310;
wire v_11311;
wire v_11312;
wire v_11313;
wire v_11314;
wire v_11315;
wire v_11316;
wire v_11317;
wire v_11318;
wire v_11319;
wire v_11320;
wire v_11321;
wire v_11322;
wire v_11323;
wire v_11324;
wire v_11325;
wire v_11326;
wire v_11327;
wire v_11328;
wire v_11329;
wire v_11330;
wire v_11331;
wire v_11332;
wire v_11333;
wire v_11334;
wire v_11335;
wire v_11336;
wire v_11337;
wire v_11338;
wire v_11339;
wire v_11340;
wire v_11341;
wire v_11342;
wire v_11343;
wire v_11344;
wire v_11345;
wire v_11346;
wire v_11347;
wire v_11348;
wire v_11349;
wire v_11350;
wire v_11351;
wire v_11352;
wire v_11353;
wire v_11354;
wire v_11355;
wire v_11356;
wire v_11357;
wire v_11358;
wire v_11359;
wire v_11360;
wire v_11361;
wire v_11362;
wire v_11363;
wire v_11364;
wire v_11365;
wire v_11366;
wire v_11367;
wire v_11368;
wire v_11369;
wire v_11370;
wire v_11371;
wire v_11372;
wire v_11373;
wire v_11374;
wire v_11375;
wire v_11376;
wire v_11377;
wire v_11378;
wire v_11379;
wire v_11380;
wire v_11381;
wire v_11382;
wire v_11383;
wire v_11384;
wire v_11385;
wire v_11386;
wire v_11387;
wire v_11388;
wire v_11389;
wire v_11390;
wire v_11391;
wire v_11392;
wire v_11393;
wire v_11394;
wire v_11395;
wire v_11396;
wire v_11397;
wire v_11398;
wire v_11399;
wire v_11400;
wire v_11401;
wire v_11402;
wire v_11403;
wire v_11404;
wire v_11405;
wire v_11406;
wire v_11407;
wire v_11408;
wire v_11409;
wire v_11410;
wire v_11411;
wire v_11412;
wire v_11413;
wire v_11414;
wire v_11415;
wire v_11416;
wire v_11417;
wire v_11418;
wire v_11419;
wire v_11420;
wire v_11421;
wire v_11422;
wire v_11423;
wire v_11424;
wire v_11425;
wire v_11426;
wire v_11427;
wire v_11428;
wire v_11429;
wire v_11430;
wire v_11431;
wire v_11432;
wire v_11433;
wire v_11434;
wire v_11435;
wire v_11436;
wire v_11437;
wire v_11438;
wire v_11439;
wire v_11440;
wire v_11441;
wire v_11442;
wire v_11443;
wire v_11444;
wire v_11445;
wire v_11446;
wire v_11447;
wire v_11448;
wire v_11449;
wire v_11450;
wire v_11451;
wire v_11452;
wire v_11453;
wire v_11454;
wire v_11455;
wire v_11456;
wire v_11457;
wire v_11458;
wire v_11459;
wire v_11460;
wire v_11461;
wire v_11462;
wire v_11463;
wire v_11464;
wire v_11465;
wire v_11466;
wire v_11467;
wire v_11468;
wire v_11469;
wire v_11470;
wire v_11471;
wire v_11472;
wire v_11473;
wire v_11474;
wire v_11475;
wire v_11476;
wire v_11477;
wire v_11478;
wire v_11479;
wire v_11480;
wire v_11481;
wire v_11482;
wire v_11483;
wire v_11484;
wire v_11485;
wire v_11486;
wire v_11487;
wire v_11488;
wire v_11489;
wire v_11490;
wire v_11491;
wire v_11492;
wire v_11493;
wire v_11494;
wire v_11495;
wire v_11496;
wire v_11497;
wire v_11498;
wire v_11499;
wire v_11500;
wire v_11501;
wire v_11502;
wire v_11503;
wire v_11504;
wire v_11505;
wire v_11506;
wire v_11507;
wire v_11508;
wire v_11509;
wire v_11510;
wire v_11511;
wire v_11512;
wire v_11513;
wire v_11514;
wire v_11515;
wire v_11516;
wire v_11517;
wire v_11518;
wire v_11519;
wire v_11520;
wire v_11521;
wire v_11522;
wire v_11523;
wire v_11524;
wire v_11525;
wire v_11526;
wire v_11527;
wire v_11528;
wire v_11529;
wire v_11530;
wire v_11531;
wire v_11532;
wire v_11533;
wire v_11534;
wire v_11535;
wire v_11536;
wire v_11537;
wire v_11538;
wire v_11539;
wire v_11540;
wire v_11541;
wire v_11542;
wire v_11543;
wire v_11544;
wire v_11545;
wire v_11546;
wire v_11547;
wire v_11548;
wire v_11549;
wire v_11550;
wire v_11551;
wire v_11552;
wire v_11553;
wire v_11554;
wire v_11555;
wire v_11556;
wire v_11557;
wire v_11558;
wire v_11559;
wire v_11560;
wire v_11561;
wire v_11562;
wire v_11563;
wire v_11564;
wire v_11565;
wire v_11566;
wire v_11567;
wire v_11568;
wire v_11569;
wire v_11570;
wire v_11571;
wire v_11572;
wire v_11573;
wire v_11574;
wire v_11575;
wire v_11576;
wire v_11577;
wire v_11578;
wire v_11579;
wire v_11580;
wire v_11581;
wire v_11582;
wire v_11583;
wire v_11584;
wire v_11585;
wire v_11586;
wire v_11587;
wire v_11588;
wire v_11589;
wire v_11590;
wire v_11591;
wire v_11592;
wire v_11593;
wire v_11594;
wire v_11595;
wire v_11596;
wire v_11597;
wire v_11598;
wire v_11599;
wire v_11600;
wire v_11601;
wire v_11602;
wire v_11603;
wire v_11604;
wire v_11605;
wire v_11606;
wire v_11607;
wire v_11608;
wire v_11609;
wire v_11610;
wire v_11611;
wire v_11612;
wire v_11613;
wire v_11614;
wire v_11615;
wire v_11616;
wire v_11617;
wire v_11618;
wire v_11619;
wire v_11620;
wire v_11621;
wire v_11622;
wire v_11623;
wire v_11624;
wire v_11625;
wire v_11626;
wire v_11627;
wire v_11628;
wire v_11629;
wire v_11630;
wire v_11631;
wire v_11632;
wire v_11633;
wire v_11634;
wire v_11635;
wire v_11636;
wire v_11637;
wire v_11638;
wire v_11639;
wire v_11640;
wire v_11641;
wire v_11642;
wire v_11643;
wire v_11644;
wire v_11645;
wire v_11646;
wire v_11647;
wire v_11648;
wire v_11649;
wire v_11650;
wire v_11651;
wire v_11652;
wire v_11653;
wire v_11654;
wire v_11655;
wire v_11656;
wire v_11657;
wire v_11658;
wire v_11659;
wire v_11660;
wire v_11661;
wire v_11662;
wire v_11663;
wire v_11664;
wire v_11665;
wire v_11666;
wire v_11667;
wire v_11668;
wire v_11669;
wire v_11670;
wire v_11671;
wire v_11672;
wire v_11673;
wire v_11674;
wire v_11675;
wire v_11676;
wire v_11677;
wire v_11678;
wire v_11679;
wire v_11680;
wire v_11681;
wire v_11682;
wire v_11683;
wire v_11684;
wire v_11685;
wire v_11686;
wire v_11687;
wire v_11688;
wire v_11689;
wire v_11690;
wire v_11691;
wire v_11692;
wire v_11693;
wire v_11694;
wire v_11695;
wire v_11696;
wire v_11697;
wire v_11698;
wire v_11699;
wire v_11700;
wire v_11701;
wire v_11702;
wire v_11703;
wire v_11704;
wire v_11705;
wire v_11706;
wire v_11707;
wire v_11708;
wire v_11709;
wire v_11710;
wire v_11711;
wire v_11712;
wire v_11713;
wire v_11714;
wire v_11715;
wire v_11716;
wire v_11717;
wire v_11718;
wire v_11719;
wire v_11720;
wire v_11721;
wire v_11722;
wire v_11723;
wire v_11724;
wire v_11725;
wire v_11726;
wire v_11727;
wire v_11728;
wire v_11729;
wire v_11730;
wire v_11731;
wire v_11732;
wire v_11733;
wire v_11734;
wire v_11735;
wire v_11736;
wire v_11737;
wire v_11738;
wire v_11739;
wire v_11740;
wire v_11741;
wire v_11742;
wire v_11743;
wire v_11744;
wire v_11745;
wire v_11746;
wire v_11747;
wire v_11748;
wire v_11749;
wire v_11750;
wire v_11751;
wire v_11752;
wire v_11753;
wire v_11754;
wire v_11755;
wire v_11756;
wire v_11757;
wire v_11758;
wire v_11759;
wire v_11760;
wire v_11761;
wire v_11762;
wire v_11763;
wire v_11764;
wire v_11765;
wire v_11766;
wire v_11767;
wire v_11768;
wire v_11769;
wire v_11770;
wire v_11771;
wire v_11772;
wire v_11773;
wire v_11774;
wire v_11775;
wire v_11776;
wire v_11777;
wire v_11778;
wire v_11779;
wire v_11780;
wire v_11781;
wire v_11782;
wire v_11783;
wire v_11784;
wire v_11785;
wire v_11786;
wire v_11787;
wire v_11788;
wire v_11789;
wire v_11790;
wire v_11791;
wire v_11792;
wire v_11793;
wire v_11794;
wire v_11795;
wire v_11796;
wire v_11797;
wire v_11798;
wire v_11799;
wire v_11800;
wire v_11801;
wire v_11802;
wire v_11803;
wire v_11804;
wire v_11805;
wire v_11806;
wire v_11807;
wire v_11808;
wire v_11809;
wire v_11810;
wire v_11811;
wire v_11812;
wire v_11813;
wire v_11814;
wire v_11815;
wire v_11816;
wire v_11817;
wire v_11818;
wire v_11819;
wire v_11820;
wire v_11821;
wire v_11822;
wire v_11823;
wire v_11824;
wire v_11825;
wire v_11826;
wire v_11827;
wire v_11828;
wire v_11829;
wire v_11830;
wire v_11831;
wire v_11832;
wire v_11833;
wire v_11834;
wire v_11835;
wire v_11836;
wire v_11837;
wire v_11838;
wire v_11839;
wire v_11840;
wire v_11841;
wire v_11842;
wire v_11843;
wire v_11844;
wire v_11845;
wire v_11846;
wire v_11847;
wire v_11848;
wire v_11849;
wire v_11850;
wire v_11851;
wire v_11852;
wire v_11853;
wire v_11854;
wire v_11855;
wire v_11856;
wire v_11857;
wire v_11858;
wire v_11859;
wire v_11860;
wire v_11861;
wire v_11862;
wire v_11863;
wire v_11864;
wire v_11865;
wire v_11866;
wire v_11867;
wire v_11868;
wire v_11869;
wire v_11870;
wire v_11871;
wire v_11872;
wire v_11873;
wire v_11874;
wire v_11875;
wire v_11876;
wire v_11877;
wire v_11878;
wire v_11879;
wire v_11880;
wire v_11881;
wire v_11882;
wire v_11883;
wire v_11884;
wire v_11885;
wire v_11886;
wire v_11887;
wire v_11888;
wire v_11889;
wire v_11890;
wire v_11891;
wire v_11892;
wire v_11893;
wire v_11894;
wire v_11895;
wire v_11896;
wire v_11897;
wire v_11898;
wire v_11899;
wire v_11900;
wire v_11901;
wire v_11902;
wire v_11903;
wire v_11904;
wire v_11905;
wire v_11906;
wire v_11907;
wire v_11908;
wire v_11909;
wire v_11910;
wire v_11911;
wire v_11912;
wire v_11913;
wire v_11914;
wire v_11915;
wire v_11916;
wire v_11917;
wire v_11918;
wire v_11919;
wire v_11920;
wire v_11921;
wire v_11922;
wire v_11923;
wire v_11924;
wire v_11925;
wire v_11926;
wire v_11927;
wire v_11928;
wire v_11929;
wire v_11930;
wire v_11931;
wire v_11932;
wire v_11933;
wire v_11934;
wire v_11935;
wire v_11936;
wire v_11937;
wire v_11938;
wire v_11939;
wire v_11940;
wire v_11941;
wire v_11942;
wire v_11943;
wire v_11944;
wire v_11945;
wire v_11946;
wire v_11947;
wire v_11948;
wire v_11949;
wire v_11950;
wire v_11951;
wire v_11952;
wire v_11953;
wire v_11954;
wire v_11955;
wire v_11956;
wire v_11957;
wire v_11958;
wire v_11959;
wire v_11960;
wire v_11961;
wire v_11962;
wire v_11963;
wire v_11964;
wire v_11965;
wire v_11966;
wire v_11967;
wire v_11968;
wire v_11969;
wire v_11970;
wire v_11971;
wire v_11972;
wire v_11973;
wire v_11974;
wire v_11975;
wire v_11976;
wire v_11977;
wire v_11978;
wire v_11979;
wire v_11980;
wire v_11981;
wire v_11982;
wire v_11983;
wire v_11984;
wire v_11985;
wire v_11986;
wire v_11987;
wire v_11988;
wire v_11989;
wire v_11990;
wire v_11991;
wire v_11992;
wire v_11993;
wire v_11994;
wire v_11995;
wire v_11996;
wire v_11997;
wire v_11998;
wire v_11999;
wire v_12000;
wire v_12001;
wire v_12002;
wire v_12003;
wire v_12004;
wire v_12005;
wire v_12006;
wire v_12007;
wire v_12008;
wire v_12009;
wire v_12010;
wire v_12011;
wire v_12012;
wire v_12013;
wire v_12014;
wire v_12015;
wire v_12016;
wire v_12017;
wire v_12018;
wire v_12019;
wire v_12020;
wire v_12021;
wire v_12022;
wire v_12023;
wire v_12024;
wire v_12025;
wire v_12026;
wire v_12027;
wire v_12028;
wire v_12029;
wire v_12030;
wire v_12031;
wire v_12032;
wire v_12033;
wire v_12034;
wire v_12035;
wire v_12036;
wire v_12037;
wire v_12038;
wire v_12039;
wire v_12040;
wire v_12041;
wire v_12042;
wire v_12043;
wire v_12044;
wire v_12045;
wire v_12046;
wire v_12047;
wire v_12048;
wire v_12049;
wire v_12050;
wire v_12051;
wire v_12052;
wire v_12053;
wire v_12054;
wire v_12055;
wire v_12056;
wire v_12057;
wire v_12058;
wire v_12059;
wire v_12060;
wire v_12061;
wire v_12062;
wire v_12063;
wire v_12064;
wire v_12065;
wire v_12066;
wire v_12067;
wire v_12068;
wire v_12069;
wire v_12070;
wire v_12071;
wire v_12072;
wire v_12073;
wire v_12074;
wire v_12075;
wire v_12076;
wire v_12077;
wire v_12078;
wire v_12079;
wire v_12080;
wire v_12081;
wire v_12082;
wire v_12083;
wire v_12084;
wire v_12085;
wire v_12086;
wire v_12087;
wire v_12088;
wire v_12089;
wire v_12090;
wire v_12091;
wire v_12092;
wire v_12093;
wire v_12094;
wire v_12095;
wire v_12096;
wire v_12097;
wire v_12098;
wire v_12099;
wire v_12100;
wire v_12101;
wire v_12102;
wire v_12103;
wire v_12104;
wire v_12105;
wire v_12106;
wire v_12107;
wire v_12108;
wire v_12109;
wire v_12110;
wire v_12111;
wire v_12112;
wire v_12113;
wire v_12114;
wire v_12115;
wire v_12116;
wire v_12117;
wire v_12118;
wire v_12119;
wire v_12120;
wire v_12121;
wire v_12122;
wire v_12123;
wire v_12124;
wire v_12125;
wire v_12126;
wire v_12127;
wire v_12128;
wire v_12129;
wire v_12130;
wire v_12131;
wire v_12132;
wire v_12133;
wire v_12134;
wire v_12135;
wire v_12136;
wire v_12137;
wire v_12138;
wire v_12139;
wire v_12140;
wire v_12141;
wire v_12142;
wire v_12143;
wire v_12144;
wire v_12145;
wire v_12146;
wire v_12147;
wire v_12148;
wire v_12149;
wire v_12150;
wire v_12151;
wire v_12152;
wire v_12153;
wire v_12154;
wire v_12155;
wire v_12156;
wire v_12157;
wire v_12158;
wire v_12159;
wire v_12160;
wire v_12161;
wire v_12162;
wire v_12163;
wire v_12164;
wire v_12165;
wire v_12166;
wire v_12167;
wire v_12168;
wire v_12169;
wire v_12170;
wire v_12171;
wire v_12172;
wire v_12173;
wire v_12174;
wire v_12175;
wire v_12176;
wire v_12177;
wire v_12178;
wire v_12179;
wire v_12180;
wire v_12181;
wire v_12182;
wire v_12183;
wire v_12184;
wire v_12185;
wire v_12186;
wire v_12187;
wire v_12188;
wire v_12189;
wire v_12190;
wire v_12191;
wire v_12192;
wire v_12193;
wire v_12194;
wire v_12195;
wire v_12196;
wire v_12197;
wire v_12198;
wire v_12199;
wire v_12200;
wire v_12201;
wire v_12202;
wire v_12203;
wire v_12204;
wire v_12205;
wire v_12206;
wire v_12207;
wire v_12208;
wire v_12209;
wire v_12210;
wire v_12211;
wire v_12212;
wire v_12213;
wire v_12214;
wire v_12215;
wire v_12216;
wire v_12217;
wire v_12218;
wire v_12219;
wire v_12220;
wire v_12221;
wire v_12222;
wire v_12223;
wire v_12224;
wire v_12225;
wire v_12226;
wire v_12227;
wire v_12228;
wire v_12229;
wire v_12230;
wire v_12231;
wire v_12232;
wire v_12233;
wire v_12234;
wire v_12235;
wire v_12236;
wire v_12237;
wire v_12238;
wire v_12239;
wire v_12240;
wire v_12241;
wire v_12242;
wire v_12243;
wire v_12244;
wire v_12245;
wire v_12246;
wire v_12247;
wire v_12248;
wire v_12249;
wire v_12250;
wire v_12251;
wire v_12252;
wire v_12253;
wire v_12254;
wire v_12255;
wire v_12256;
wire v_12257;
wire v_12258;
wire v_12259;
wire v_12260;
wire v_12261;
wire v_12262;
wire v_12263;
wire v_12264;
wire v_12265;
wire v_12266;
wire v_12267;
wire v_12268;
wire v_12269;
wire v_12270;
wire v_12271;
wire v_12272;
wire v_12273;
wire v_12274;
wire v_12275;
wire v_12276;
wire v_12277;
wire v_12278;
wire v_12279;
wire v_12280;
wire v_12281;
wire v_12282;
wire v_12283;
wire v_12284;
wire v_12285;
wire v_12286;
wire v_12287;
wire v_12288;
wire v_12289;
wire v_12290;
wire v_12291;
wire v_12292;
wire v_12293;
wire v_12294;
wire v_12295;
wire v_12296;
wire v_12297;
wire v_12298;
wire v_12299;
wire v_12300;
wire v_12301;
wire v_12302;
wire v_12303;
wire v_12304;
wire v_12305;
wire v_12306;
wire v_12307;
wire v_12308;
wire v_12309;
wire v_12310;
wire v_12311;
wire v_12312;
wire v_12313;
wire v_12314;
wire v_12315;
wire v_12316;
wire v_12317;
wire v_12318;
wire v_12319;
wire v_12320;
wire v_12321;
wire v_12322;
wire v_12323;
wire v_12324;
wire v_12325;
wire v_12326;
wire v_12327;
wire v_12328;
wire v_12329;
wire v_12330;
wire v_12331;
wire v_12332;
wire v_12333;
wire v_12334;
wire v_12335;
wire v_12336;
wire v_12337;
wire v_12338;
wire v_12339;
wire v_12340;
wire v_12341;
wire v_12342;
wire v_12343;
wire v_12344;
wire v_12345;
wire v_12346;
wire v_12347;
wire v_12348;
wire v_12349;
wire v_12350;
wire v_12351;
wire v_12352;
wire v_12353;
wire v_12354;
wire v_12355;
wire v_12356;
wire v_12357;
wire v_12358;
wire v_12359;
wire v_12360;
wire v_12361;
wire v_12362;
wire v_12363;
wire v_12364;
wire v_12365;
wire v_12366;
wire v_12367;
wire v_12368;
wire v_12369;
wire v_12370;
wire v_12371;
wire v_12372;
wire v_12373;
wire v_12374;
wire v_12375;
wire v_12376;
wire v_12377;
wire v_12378;
wire v_12379;
wire v_12380;
wire v_12381;
wire v_12382;
wire v_12383;
wire v_12384;
wire v_12385;
wire v_12386;
wire v_12387;
wire v_12388;
wire v_12389;
wire v_12390;
wire v_12391;
wire v_12392;
wire v_12393;
wire v_12394;
wire v_12395;
wire v_12396;
wire v_12397;
wire v_12398;
wire v_12399;
wire v_12400;
wire v_12401;
wire v_12402;
wire v_12403;
wire v_12404;
wire v_12405;
wire v_12406;
wire v_12407;
wire v_12408;
wire v_12409;
wire v_12410;
wire v_12411;
wire v_12412;
wire v_12413;
wire v_12414;
wire v_12415;
wire v_12416;
wire v_12417;
wire v_12418;
wire v_12419;
wire v_12420;
wire v_12421;
wire v_12422;
wire v_12423;
wire v_12424;
wire v_12425;
wire v_12426;
wire v_12427;
wire v_12428;
wire v_12429;
wire v_12430;
wire v_12431;
wire v_12432;
wire v_12433;
wire v_12434;
wire v_12435;
wire v_12436;
wire v_12437;
wire v_12438;
wire v_12439;
wire v_12440;
wire v_12441;
wire v_12442;
wire v_12443;
wire v_12444;
wire v_12445;
wire v_12446;
wire v_12447;
wire v_12448;
wire v_12449;
wire v_12450;
wire v_12451;
wire v_12452;
wire v_12453;
wire v_12454;
wire v_12455;
wire v_12456;
wire v_12457;
wire v_12458;
wire v_12459;
wire v_12460;
wire v_12461;
wire v_12462;
wire v_12463;
wire v_12464;
wire v_12465;
wire v_12466;
wire v_12467;
wire v_12468;
wire v_12469;
wire v_12470;
wire v_12471;
wire v_12472;
wire v_12473;
wire v_12474;
wire v_12475;
wire v_12476;
wire v_12477;
wire v_12478;
wire v_12479;
wire v_12480;
wire v_12481;
wire v_12482;
wire v_12483;
wire v_12484;
wire v_12485;
wire v_12486;
wire v_12487;
wire v_12488;
wire v_12489;
wire v_12490;
wire v_12491;
wire v_12492;
wire v_12493;
wire v_12494;
wire v_12495;
wire v_12496;
wire v_12497;
wire v_12498;
wire v_12499;
wire v_12500;
wire v_12501;
wire v_12502;
wire v_12503;
wire v_12504;
wire v_12505;
wire v_12506;
wire v_12507;
wire v_12508;
wire v_12509;
wire v_12510;
wire v_12511;
wire v_12512;
wire v_12513;
wire v_12514;
wire v_12515;
wire v_12516;
wire v_12517;
wire v_12518;
wire v_12519;
wire v_12520;
wire v_12521;
wire v_12522;
wire v_12523;
wire v_12524;
wire v_12525;
wire v_12526;
wire v_12527;
wire v_12528;
wire v_12529;
wire v_12530;
wire v_12531;
wire v_12532;
wire v_12533;
wire v_12534;
wire v_12535;
wire v_12536;
wire v_12537;
wire v_12538;
wire v_12539;
wire v_12540;
wire v_12541;
wire v_12542;
wire v_12543;
wire v_12544;
wire v_12545;
wire v_12546;
wire v_12547;
wire v_12548;
wire v_12549;
wire v_12550;
wire v_12551;
wire v_12552;
wire v_12553;
wire v_12554;
wire v_12555;
wire v_12556;
wire v_12557;
wire v_12558;
wire v_12559;
wire v_12560;
wire v_12561;
wire v_12562;
wire v_12563;
wire v_12564;
wire v_12565;
wire v_12566;
wire v_12567;
wire v_12568;
wire v_12569;
wire v_12570;
wire v_12571;
wire v_12572;
wire v_12573;
wire v_12574;
wire v_12575;
wire v_12576;
wire v_12577;
wire v_12578;
wire v_12579;
wire v_12580;
wire v_12581;
wire v_12582;
wire v_12583;
wire v_12584;
wire v_12585;
wire v_12586;
wire v_12587;
wire v_12588;
wire v_12589;
wire v_12590;
wire v_12591;
wire v_12592;
wire v_12593;
wire v_12594;
wire v_12595;
wire v_12596;
wire v_12597;
wire v_12598;
wire v_12599;
wire v_12600;
wire v_12601;
wire v_12602;
wire v_12603;
wire v_12604;
wire v_12605;
wire v_12606;
wire v_12607;
wire v_12608;
wire v_12609;
wire v_12610;
wire v_12611;
wire v_12612;
wire v_12613;
wire v_12614;
wire v_12615;
wire v_12616;
wire v_12617;
wire v_12618;
wire v_12619;
wire v_12620;
wire v_12621;
wire v_12622;
wire v_12623;
wire v_12624;
wire v_12625;
wire v_12626;
wire v_12627;
wire v_12628;
wire v_12629;
wire v_12630;
wire v_12631;
wire v_12632;
wire v_12633;
wire v_12634;
wire v_12635;
wire v_12636;
wire v_12637;
wire v_12638;
wire v_12639;
wire v_12640;
wire v_12641;
wire v_12642;
wire v_12643;
wire v_12644;
wire v_12645;
wire v_12646;
wire v_12647;
wire v_12648;
wire v_12649;
wire v_12650;
wire v_12651;
wire v_12652;
wire v_12653;
wire v_12654;
wire v_12655;
wire v_12656;
wire v_12657;
wire v_12658;
wire v_12659;
wire v_12660;
wire v_12661;
wire v_12662;
wire v_12663;
wire v_12664;
wire v_12665;
wire v_12666;
wire v_12667;
wire v_12668;
wire v_12669;
wire v_12670;
wire v_12671;
wire v_12672;
wire v_12673;
wire v_12674;
wire v_12675;
wire v_12676;
wire v_12677;
wire v_12678;
wire v_12679;
wire v_12680;
wire v_12681;
wire v_12682;
wire v_12683;
wire v_12684;
wire v_12685;
wire v_12686;
wire v_12687;
wire v_12688;
wire v_12689;
wire v_12690;
wire v_12691;
wire v_12692;
wire v_12693;
wire v_12694;
wire v_12695;
wire v_12696;
wire v_12697;
wire v_12698;
wire v_12699;
wire v_12700;
wire v_12701;
wire v_12702;
wire v_12703;
wire v_12704;
wire v_12705;
wire v_12706;
wire v_12707;
wire v_12708;
wire v_12709;
wire v_12710;
wire v_12711;
wire v_12712;
wire v_12713;
wire v_12714;
wire v_12715;
wire v_12716;
wire v_12717;
wire v_12718;
wire v_12719;
wire v_12720;
wire v_12721;
wire v_12722;
wire v_12723;
wire v_12724;
wire v_12725;
wire v_12726;
wire v_12727;
wire v_12728;
wire v_12729;
wire v_12730;
wire v_12731;
wire v_12732;
wire v_12733;
wire v_12734;
wire v_12735;
wire v_12736;
wire v_12737;
wire v_12738;
wire v_12739;
wire v_12740;
wire v_12741;
wire v_12742;
wire v_12743;
wire v_12744;
wire v_12745;
wire v_12746;
wire v_12747;
wire v_12748;
wire v_12749;
wire v_12750;
wire v_12751;
wire v_12752;
wire v_12753;
wire v_12754;
wire v_12755;
wire v_12756;
wire v_12757;
wire v_12758;
wire v_12759;
wire v_12760;
wire v_12761;
wire v_12762;
wire v_12763;
wire v_12764;
wire v_12765;
wire v_12766;
wire v_12767;
wire v_12768;
wire v_12769;
wire v_12770;
wire v_12771;
wire v_12772;
wire v_12773;
wire v_12774;
wire v_12775;
wire v_12776;
wire v_12777;
wire v_12778;
wire v_12779;
wire v_12780;
wire v_12781;
wire v_12782;
wire v_12783;
wire v_12784;
wire v_12785;
wire v_12786;
wire v_12787;
wire v_12788;
wire v_12789;
wire v_12790;
wire v_12791;
wire v_12792;
wire v_12793;
wire v_12794;
wire v_12795;
wire v_12796;
wire v_12797;
wire v_12798;
wire v_12799;
wire v_12800;
wire v_12801;
wire v_12802;
wire v_12803;
wire v_12804;
wire v_12805;
wire v_12806;
wire v_12807;
wire v_12808;
wire v_12809;
wire v_12810;
wire v_12811;
wire v_12812;
wire v_12813;
wire v_12814;
wire v_12815;
wire v_12816;
wire v_12817;
wire v_12818;
wire v_12819;
wire v_12820;
wire v_12821;
wire v_12822;
wire v_12823;
wire v_12824;
wire v_12825;
wire v_12826;
wire v_12827;
wire v_12828;
wire v_12829;
wire v_12830;
wire v_12831;
wire v_12832;
wire v_12833;
wire v_12834;
wire v_12835;
wire v_12836;
wire v_12837;
wire v_12838;
wire v_12839;
wire v_12840;
wire v_12841;
wire v_12842;
wire v_12843;
wire v_12844;
wire v_12845;
wire v_12846;
wire v_12847;
wire v_12848;
wire v_12849;
wire v_12850;
wire v_12851;
wire v_12852;
wire v_12853;
wire v_12854;
wire v_12855;
wire v_12856;
wire v_12857;
wire v_12858;
wire v_12859;
wire v_12860;
wire v_12861;
wire v_12862;
wire v_12863;
wire v_12864;
wire v_12865;
wire v_12866;
wire v_12867;
wire v_12868;
wire v_12869;
wire v_12870;
wire v_12871;
wire v_12872;
wire v_12873;
wire v_12874;
wire v_12875;
wire v_12876;
wire v_12877;
wire v_12878;
wire v_12879;
wire v_12880;
wire v_12881;
wire v_12882;
wire v_12883;
wire v_12884;
wire v_12885;
wire v_12886;
wire v_12887;
wire v_12888;
wire v_12889;
wire v_12890;
wire v_12891;
wire v_12892;
wire v_12893;
wire v_12894;
wire v_12895;
wire v_12896;
wire v_12897;
wire v_12898;
wire v_12899;
wire v_12900;
wire v_12901;
wire v_12902;
wire v_12903;
wire v_12904;
wire v_12905;
wire v_12906;
wire v_12907;
wire v_12908;
wire v_12909;
wire v_12910;
wire v_12911;
wire v_12912;
wire v_12913;
wire v_12914;
wire v_12915;
wire v_12916;
wire v_12917;
wire v_12918;
wire v_12919;
wire v_12920;
wire v_12921;
wire v_12922;
wire v_12923;
wire v_12924;
wire v_12925;
wire v_12926;
wire v_12927;
wire v_12928;
wire v_12929;
wire v_12930;
wire v_12931;
wire v_12932;
wire v_12933;
wire v_12934;
wire v_12935;
wire v_12936;
wire v_12937;
wire v_12938;
wire v_12939;
wire v_12940;
wire v_12941;
wire v_12942;
wire v_12943;
wire v_12944;
wire v_12945;
wire v_12946;
wire v_12947;
wire v_12948;
wire v_12949;
wire v_12950;
wire v_12951;
wire v_12952;
wire v_12953;
wire v_12954;
wire v_12955;
wire v_12956;
wire v_12957;
wire v_12958;
wire v_12959;
wire v_12960;
wire v_12961;
wire v_12962;
wire v_12963;
wire v_12964;
wire v_12965;
wire v_12966;
wire v_12967;
wire v_12968;
wire v_12969;
wire v_12970;
wire v_12971;
wire v_12972;
wire v_12973;
wire v_12974;
wire v_12975;
wire v_12976;
wire v_12977;
wire v_12978;
wire v_12979;
wire v_12980;
wire v_12981;
wire v_12982;
wire v_12983;
wire v_12984;
wire v_12985;
wire v_12986;
wire v_12987;
wire v_12988;
wire v_12989;
wire v_12990;
wire v_12991;
wire v_12992;
wire v_12993;
wire v_12994;
wire v_12995;
wire v_12996;
wire v_12997;
wire v_12998;
wire v_12999;
wire v_13000;
wire v_13001;
wire v_13002;
wire v_13003;
wire v_13004;
wire v_13005;
wire v_13006;
wire v_13007;
wire v_13008;
wire v_13009;
wire v_13010;
wire v_13011;
wire v_13012;
wire v_13013;
wire v_13014;
wire v_13015;
wire v_13016;
wire v_13017;
wire v_13018;
wire v_13019;
wire v_13020;
wire v_13021;
wire v_13022;
wire v_13023;
wire v_13024;
wire v_13025;
wire v_13026;
wire v_13027;
wire v_13028;
wire v_13029;
wire v_13030;
wire v_13031;
wire v_13032;
wire v_13033;
wire v_13034;
wire v_13035;
wire v_13036;
wire v_13037;
wire v_13038;
wire v_13039;
wire v_13040;
wire v_13041;
wire v_13042;
wire v_13043;
wire v_13044;
wire v_13045;
wire v_13046;
wire v_13047;
wire v_13048;
wire v_13049;
wire v_13050;
wire v_13051;
wire v_13052;
wire v_13053;
wire v_13054;
wire v_13055;
wire v_13056;
wire v_13057;
wire v_13058;
wire v_13059;
wire v_13060;
wire v_13061;
wire v_13062;
wire v_13063;
wire v_13064;
wire v_13065;
wire v_13066;
wire v_13067;
wire v_13068;
wire v_13069;
wire v_13070;
wire v_13071;
wire v_13072;
wire v_13073;
wire v_13074;
wire v_13075;
wire v_13076;
wire v_13077;
wire v_13078;
wire v_13079;
wire v_13080;
wire v_13081;
wire v_13082;
wire v_13083;
wire v_13084;
wire v_13085;
wire v_13086;
wire v_13087;
wire v_13088;
wire v_13089;
wire v_13090;
wire v_13091;
wire v_13092;
wire v_13093;
wire v_13094;
wire v_13095;
wire v_13096;
wire v_13097;
wire v_13098;
wire v_13099;
wire v_13100;
wire v_13101;
wire v_13102;
wire v_13103;
wire v_13104;
wire v_13105;
wire v_13106;
wire v_13107;
wire v_13108;
wire v_13109;
wire v_13110;
wire v_13111;
wire v_13112;
wire v_13113;
wire v_13114;
wire v_13115;
wire v_13116;
wire v_13117;
wire v_13118;
wire v_13119;
wire v_13120;
wire v_13121;
wire v_13122;
wire v_13123;
wire v_13124;
wire v_13125;
wire v_13126;
wire v_13127;
wire v_13128;
wire v_13129;
wire v_13130;
wire v_13131;
wire v_13132;
wire v_13133;
wire v_13134;
wire v_13135;
wire v_13136;
wire v_13137;
wire v_13138;
wire v_13139;
wire v_13140;
wire v_13141;
wire v_13142;
wire v_13143;
wire v_13144;
wire v_13145;
wire v_13146;
wire v_13147;
wire v_13148;
wire v_13149;
wire v_13150;
wire v_13151;
wire v_13152;
wire v_13153;
wire v_13154;
wire v_13155;
wire v_13156;
wire v_13157;
wire v_13158;
wire v_13159;
wire v_13160;
wire v_13161;
wire v_13162;
wire v_13163;
wire v_13164;
wire v_13165;
wire v_13166;
wire v_13167;
wire v_13168;
wire v_13169;
wire v_13170;
wire v_13171;
wire v_13172;
wire v_13173;
wire v_13174;
wire v_13175;
wire v_13176;
wire v_13177;
wire v_13178;
wire v_13179;
wire v_13180;
wire v_13181;
wire v_13182;
wire v_13183;
wire v_13184;
wire v_13185;
wire v_13186;
wire v_13187;
wire v_13188;
wire v_13189;
wire v_13190;
wire v_13191;
wire v_13192;
wire v_13193;
wire v_13194;
wire v_13195;
wire v_13196;
wire v_13197;
wire v_13198;
wire v_13199;
wire v_13200;
wire v_13201;
wire v_13202;
wire v_13203;
wire v_13204;
wire v_13205;
wire v_13206;
wire v_13207;
wire v_13208;
wire v_13209;
wire v_13210;
wire v_13211;
wire v_13212;
wire v_13213;
wire v_13214;
wire v_13215;
wire v_13216;
wire v_13217;
wire v_13218;
wire v_13219;
wire v_13220;
wire v_13221;
wire v_13222;
wire v_13223;
wire v_13224;
wire v_13225;
wire v_13226;
wire v_13227;
wire v_13228;
wire v_13229;
wire v_13230;
wire v_13231;
wire v_13232;
wire v_13233;
wire v_13234;
wire v_13235;
wire v_13236;
wire v_13237;
wire v_13238;
wire v_13239;
wire v_13240;
wire v_13241;
wire v_13242;
wire v_13243;
wire v_13244;
wire v_13245;
wire v_13246;
wire v_13247;
wire v_13248;
wire v_13249;
wire v_13250;
wire v_13251;
wire v_13252;
wire v_13253;
wire v_13254;
wire v_13255;
wire v_13256;
wire v_13257;
wire v_13258;
wire v_13259;
wire v_13260;
wire v_13261;
wire v_13262;
wire v_13263;
wire v_13264;
wire v_13265;
wire v_13266;
wire v_13267;
wire v_13268;
wire v_13269;
wire v_13270;
wire v_13271;
wire v_13272;
wire v_13273;
wire v_13274;
wire v_13275;
wire v_13276;
wire v_13277;
wire v_13278;
wire v_13279;
wire v_13280;
wire v_13281;
wire v_13282;
wire v_13283;
wire v_13284;
wire v_13285;
wire v_13286;
wire v_13287;
wire v_13288;
wire v_13289;
wire v_13290;
wire v_13291;
wire v_13292;
wire v_13293;
wire v_13294;
wire v_13295;
wire v_13296;
wire v_13297;
wire v_13298;
wire v_13299;
wire v_13300;
wire v_13301;
wire v_13302;
wire v_13303;
wire v_13304;
wire v_13305;
wire v_13306;
wire v_13307;
wire v_13308;
wire v_13309;
wire v_13310;
wire v_13311;
wire v_13312;
wire v_13313;
wire v_13314;
wire v_13315;
wire v_13316;
wire v_13317;
wire v_13318;
wire v_13319;
wire v_13320;
wire v_13321;
wire v_13322;
wire v_13323;
wire v_13324;
wire v_13325;
wire v_13326;
wire v_13327;
wire v_13328;
wire v_13329;
wire v_13330;
wire v_13331;
wire v_13332;
wire v_13333;
wire v_13334;
wire v_13335;
wire v_13336;
wire v_13337;
wire v_13338;
wire v_13339;
wire v_13340;
wire v_13341;
wire v_13342;
wire v_13343;
wire v_13344;
wire v_13345;
wire v_13346;
wire v_13347;
wire v_13348;
wire v_13349;
wire v_13350;
wire v_13351;
wire v_13352;
wire v_13353;
wire v_13354;
wire v_13355;
wire v_13356;
wire v_13357;
wire v_13358;
wire v_13359;
wire v_13360;
wire v_13361;
wire v_13362;
wire v_13363;
wire v_13364;
wire v_13365;
wire v_13366;
wire v_13367;
wire v_13368;
wire v_13369;
wire v_13370;
wire v_13371;
wire v_13372;
wire v_13373;
wire v_13374;
wire v_13375;
wire v_13376;
wire v_13377;
wire v_13378;
wire v_13379;
wire v_13380;
wire v_13381;
wire v_13382;
wire v_13383;
wire v_13384;
wire v_13385;
wire v_13386;
wire v_13387;
wire v_13388;
wire v_13389;
wire v_13390;
wire v_13391;
wire v_13392;
wire v_13393;
wire v_13394;
wire v_13395;
wire v_13396;
wire v_13397;
wire v_13398;
wire v_13399;
wire v_13400;
wire v_13401;
wire v_13402;
wire v_13403;
wire v_13404;
wire v_13405;
wire v_13406;
wire v_13407;
wire v_13408;
wire v_13409;
wire v_13410;
wire v_13411;
wire v_13412;
wire v_13413;
wire v_13414;
wire v_13415;
wire v_13416;
wire v_13417;
wire v_13418;
wire v_13419;
wire v_13420;
wire v_13421;
wire v_13422;
wire v_13423;
wire v_13424;
wire v_13425;
wire v_13426;
wire v_13427;
wire v_13428;
wire v_13429;
wire v_13430;
wire v_13431;
wire v_13432;
wire v_13433;
wire v_13434;
wire v_13435;
wire v_13436;
wire v_13437;
wire v_13438;
wire v_13439;
wire v_13440;
wire v_13441;
wire v_13442;
wire v_13443;
wire v_13444;
wire v_13445;
wire v_13446;
wire v_13447;
wire v_13448;
wire v_13449;
wire v_13450;
wire v_13451;
wire v_13452;
wire v_13453;
wire v_13454;
wire v_13455;
wire v_13456;
wire v_13457;
wire v_13458;
wire v_13459;
wire v_13460;
wire v_13461;
wire v_13462;
wire v_13463;
wire v_13464;
wire v_13465;
wire v_13466;
wire v_13467;
wire v_13468;
wire v_13469;
wire v_13470;
wire v_13471;
wire v_13472;
wire v_13473;
wire v_13474;
wire v_13475;
wire v_13476;
wire v_13477;
wire v_13478;
wire v_13479;
wire v_13480;
wire v_13481;
wire v_13482;
wire v_13483;
wire v_13484;
wire v_13485;
wire v_13486;
wire v_13487;
wire v_13488;
wire v_13489;
wire v_13490;
wire v_13491;
wire v_13492;
wire v_13493;
wire v_13494;
wire v_13495;
wire v_13496;
wire v_13497;
wire v_13498;
wire v_13499;
wire v_13500;
wire v_13501;
wire v_13502;
wire v_13503;
wire v_13504;
wire v_13505;
wire v_13506;
wire v_13507;
wire v_13508;
wire v_13509;
wire v_13510;
wire v_13511;
wire v_13512;
wire v_13513;
wire v_13514;
wire v_13515;
wire v_13516;
wire v_13517;
wire v_13518;
wire v_13519;
wire v_13520;
wire v_13521;
wire v_13522;
wire v_13523;
wire v_13524;
wire v_13525;
wire v_13526;
wire v_13527;
wire v_13528;
wire v_13529;
wire v_13530;
wire v_13531;
wire v_13532;
wire v_13533;
wire v_13534;
wire v_13535;
wire v_13536;
wire v_13537;
wire v_13538;
wire v_13539;
wire v_13540;
wire v_13541;
wire v_13542;
wire v_13543;
wire v_13544;
wire v_13545;
wire v_13546;
wire v_13547;
wire v_13548;
wire v_13549;
wire v_13550;
wire v_13551;
wire v_13552;
wire v_13553;
wire v_13554;
wire v_13555;
wire v_13556;
wire v_13557;
wire v_13558;
wire v_13559;
wire v_13560;
wire v_13561;
wire v_13562;
wire v_13563;
wire v_13564;
wire v_13565;
wire v_13566;
wire v_13567;
wire v_13568;
wire v_13569;
wire v_13570;
wire v_13571;
wire v_13572;
wire v_13573;
wire v_13574;
wire v_13575;
wire v_13576;
wire v_13577;
wire v_13578;
wire v_13579;
wire v_13580;
wire v_13581;
wire v_13582;
wire v_13583;
wire v_13584;
wire v_13585;
wire v_13586;
wire v_13587;
wire v_13588;
wire v_13589;
wire v_13590;
wire v_13591;
wire v_13592;
wire v_13593;
wire v_13594;
wire v_13595;
wire v_13596;
wire v_13597;
wire v_13598;
wire v_13599;
wire v_13600;
wire v_13601;
wire v_13602;
wire v_13603;
wire v_13604;
wire v_13605;
wire v_13606;
wire v_13607;
wire v_13608;
wire v_13609;
wire v_13610;
wire v_13611;
wire v_13612;
wire v_13613;
wire v_13614;
wire v_13615;
wire v_13616;
wire v_13617;
wire v_13618;
wire v_13619;
wire v_13620;
wire v_13621;
wire v_13622;
wire v_13623;
wire v_13624;
wire v_13625;
wire v_13626;
wire v_13627;
wire v_13628;
wire v_13629;
wire v_13630;
wire v_13631;
wire v_13632;
wire v_13633;
wire v_13634;
wire v_13635;
wire v_13636;
wire v_13637;
wire v_13638;
wire v_13639;
wire v_13640;
wire v_13641;
wire v_13642;
wire v_13643;
wire v_13644;
wire v_13645;
wire v_13646;
wire v_13647;
wire v_13648;
wire v_13649;
wire v_13650;
wire v_13651;
wire v_13652;
wire v_13653;
wire v_13654;
wire v_13655;
wire v_13656;
wire v_13657;
wire v_13658;
wire v_13659;
wire v_13660;
wire v_13661;
wire v_13662;
wire v_13663;
wire v_13664;
wire v_13665;
wire v_13666;
wire v_13667;
wire v_13668;
wire v_13669;
wire v_13670;
wire v_13671;
wire v_13672;
wire v_13673;
wire v_13674;
wire v_13675;
wire v_13676;
wire v_13677;
wire v_13678;
wire v_13679;
wire v_13680;
wire v_13681;
wire v_13682;
wire v_13683;
wire v_13684;
wire v_13685;
wire v_13686;
wire v_13687;
wire v_13688;
wire v_13689;
wire v_13690;
wire v_13691;
wire v_13692;
wire v_13693;
wire v_13694;
wire v_13695;
wire v_13696;
wire v_13697;
wire v_13698;
wire v_13699;
wire v_13700;
wire v_13701;
wire v_13702;
wire v_13703;
wire v_13704;
wire v_13705;
wire v_13706;
wire v_13707;
wire v_13708;
wire v_13709;
wire v_13710;
wire v_13711;
wire v_13712;
wire v_13713;
wire v_13714;
wire v_13715;
wire v_13716;
wire v_13717;
wire v_13718;
wire v_13719;
wire v_13720;
wire v_13721;
wire v_13722;
wire v_13723;
wire v_13724;
wire v_13725;
wire v_13726;
wire v_13727;
wire v_13728;
wire v_13729;
wire v_13730;
wire v_13731;
wire v_13732;
wire v_13733;
wire v_13734;
wire v_13735;
wire v_13736;
wire v_13737;
wire v_13738;
wire v_13739;
wire v_13740;
wire v_13741;
wire v_13742;
wire v_13743;
wire v_13744;
wire v_13745;
wire v_13746;
wire v_13747;
wire v_13748;
wire v_13749;
wire v_13750;
wire v_13751;
wire v_13752;
wire v_13753;
wire v_13754;
wire v_13755;
wire v_13756;
wire v_13757;
wire v_13758;
wire v_13759;
wire v_13760;
wire v_13761;
wire v_13762;
wire v_13763;
wire v_13764;
wire v_13765;
wire v_13766;
wire v_13767;
wire v_13768;
wire v_13769;
wire v_13770;
wire v_13771;
wire v_13772;
wire v_13773;
wire v_13774;
wire v_13775;
wire v_13776;
wire v_13777;
wire v_13778;
wire v_13779;
wire v_13780;
wire v_13781;
wire v_13782;
wire v_13783;
wire v_13784;
wire v_13785;
wire v_13786;
wire v_13787;
wire v_13788;
wire v_13789;
wire v_13790;
wire v_13791;
wire v_13792;
wire v_13793;
wire v_13794;
wire v_13795;
wire v_13796;
wire v_13797;
wire v_13798;
wire v_13799;
wire v_13800;
wire v_13801;
wire v_13802;
wire v_13803;
wire v_13804;
wire v_13805;
wire v_13806;
wire v_13807;
wire v_13808;
wire v_13809;
wire v_13810;
wire v_13811;
wire v_13812;
wire v_13813;
wire v_13814;
wire v_13815;
wire v_13816;
wire v_13817;
wire v_13818;
wire v_13819;
wire v_13820;
wire v_13821;
wire v_13822;
wire v_13823;
wire v_13824;
wire v_13825;
wire v_13826;
wire v_13827;
wire v_13828;
wire v_13829;
wire v_13830;
wire v_13831;
wire v_13832;
wire v_13833;
wire v_13834;
wire v_13835;
wire v_13836;
wire v_13837;
wire v_13838;
wire v_13839;
wire v_13840;
wire v_13841;
wire v_13842;
wire v_13843;
wire v_13844;
wire v_13845;
wire v_13846;
wire v_13847;
wire v_13848;
wire v_13849;
wire v_13850;
wire v_13851;
wire v_13852;
wire v_13853;
wire v_13854;
wire v_13855;
wire v_13856;
wire v_13857;
wire v_13858;
wire v_13859;
wire v_13860;
wire v_13861;
wire v_13862;
wire v_13863;
wire v_13864;
wire v_13865;
wire v_13866;
wire v_13867;
wire v_13868;
wire v_13869;
wire v_13870;
wire v_13871;
wire v_13872;
wire v_13873;
wire v_13874;
wire v_13875;
wire v_13876;
wire v_13877;
wire v_13878;
wire v_13879;
wire v_13880;
wire v_13881;
wire v_13882;
wire v_13883;
wire v_13884;
wire v_13885;
wire v_13886;
wire v_13887;
wire v_13888;
wire v_13889;
wire v_13890;
wire v_13891;
wire v_13892;
wire v_13893;
wire v_13894;
wire v_13895;
wire v_13896;
wire v_13897;
wire v_13898;
wire v_13899;
wire v_13900;
wire v_13901;
wire v_13902;
wire v_13903;
wire v_13904;
wire v_13905;
wire v_13906;
wire v_13907;
wire v_13908;
wire v_13909;
wire v_13910;
wire v_13911;
wire v_13912;
wire v_13913;
wire v_13914;
wire v_13915;
wire v_13916;
wire v_13917;
wire v_13918;
wire v_13919;
wire v_13920;
wire v_13921;
wire v_13922;
wire v_13923;
wire v_13924;
wire v_13925;
wire v_13926;
wire v_13927;
wire v_13928;
wire v_13929;
wire v_13930;
wire v_13931;
wire v_13932;
wire v_13933;
wire v_13934;
wire v_13935;
wire v_13936;
wire v_13937;
wire v_13938;
wire v_13939;
wire v_13940;
wire v_13941;
wire v_13942;
wire v_13943;
wire v_13944;
wire v_13945;
wire v_13946;
wire v_13947;
wire v_13948;
wire v_13949;
wire v_13950;
wire v_13951;
wire v_13952;
wire v_13953;
wire v_13954;
wire v_13955;
wire v_13956;
wire v_13957;
wire v_13958;
wire v_13959;
wire v_13960;
wire v_13961;
wire v_13962;
wire v_13963;
wire v_13964;
wire v_13965;
wire v_13966;
wire v_13967;
wire v_13968;
wire v_13969;
wire v_13970;
wire v_13971;
wire v_13972;
wire v_13973;
wire v_13974;
wire v_13975;
wire v_13976;
wire v_13977;
wire v_13978;
wire v_13979;
wire v_13980;
wire v_13981;
wire v_13982;
wire v_13983;
wire v_13984;
wire v_13985;
wire v_13986;
wire v_13987;
wire v_13988;
wire v_13989;
wire v_13990;
wire v_13991;
wire v_13992;
wire v_13993;
wire v_13994;
wire v_13995;
wire v_13996;
wire v_13997;
wire v_13998;
wire v_13999;
wire v_14000;
wire v_14001;
wire v_14002;
wire v_14003;
wire v_14004;
wire v_14005;
wire v_14006;
wire v_14007;
wire v_14008;
wire v_14009;
wire v_14010;
wire v_14011;
wire v_14012;
wire v_14013;
wire v_14014;
wire v_14015;
wire v_14016;
wire v_14017;
wire v_14018;
wire v_14019;
wire v_14020;
wire v_14021;
wire v_14022;
wire v_14023;
wire v_14024;
wire v_14025;
wire v_14026;
wire v_14027;
wire v_14028;
wire v_14029;
wire v_14030;
wire v_14031;
wire v_14032;
wire v_14033;
wire v_14034;
wire v_14035;
wire v_14036;
wire v_14037;
wire v_14038;
wire v_14039;
wire v_14040;
wire v_14041;
wire v_14042;
wire v_14043;
wire v_14044;
wire v_14045;
wire v_14046;
wire v_14047;
wire v_14048;
wire v_14049;
wire v_14050;
wire v_14051;
wire v_14052;
wire v_14053;
wire v_14054;
wire v_14055;
wire v_14056;
wire v_14057;
wire v_14058;
wire v_14059;
wire v_14060;
wire v_14061;
wire v_14062;
wire v_14063;
wire v_14064;
wire v_14065;
wire v_14066;
wire v_14067;
wire v_14068;
wire v_14069;
wire v_14070;
wire v_14071;
wire v_14072;
wire v_14073;
wire v_14074;
wire v_14075;
wire v_14076;
wire v_14077;
wire v_14078;
wire v_14079;
wire v_14080;
wire v_14081;
wire v_14082;
wire v_14083;
wire v_14084;
wire v_14085;
wire v_14086;
wire v_14087;
wire v_14088;
wire v_14089;
wire v_14090;
wire v_14091;
wire v_14092;
wire v_14093;
wire v_14094;
wire v_14095;
wire v_14096;
wire v_14097;
wire v_14098;
wire v_14099;
wire v_14100;
wire v_14101;
wire v_14102;
wire v_14103;
wire v_14104;
wire v_14105;
wire v_14106;
wire v_14107;
wire v_14108;
wire v_14109;
wire v_14110;
wire v_14111;
wire v_14112;
wire v_14113;
wire v_14114;
wire v_14115;
wire v_14116;
wire v_14117;
wire v_14118;
wire v_14119;
wire v_14120;
wire v_14121;
wire v_14122;
wire v_14123;
wire v_14124;
wire v_14125;
wire v_14126;
wire v_14127;
wire v_14128;
wire v_14129;
wire v_14130;
wire v_14131;
wire v_14132;
wire v_14133;
wire v_14134;
wire v_14135;
wire v_14136;
wire v_14137;
wire v_14138;
wire v_14139;
wire v_14140;
wire v_14141;
wire v_14142;
wire v_14143;
wire v_14144;
wire v_14145;
wire v_14146;
wire v_14147;
wire v_14148;
wire v_14149;
wire v_14150;
wire v_14151;
wire v_14152;
wire v_14153;
wire v_14154;
wire v_14155;
wire v_14156;
wire v_14157;
wire v_14158;
wire v_14159;
wire v_14160;
wire v_14161;
wire v_14162;
wire v_14163;
wire v_14164;
wire v_14165;
wire v_14166;
wire v_14167;
wire v_14168;
wire v_14169;
wire v_14170;
wire v_14171;
wire v_14172;
wire v_14173;
wire v_14174;
wire v_14175;
wire v_14176;
wire v_14177;
wire v_14178;
wire v_14179;
wire v_14180;
wire v_14181;
wire v_14182;
wire v_14183;
wire v_14184;
wire v_14185;
wire v_14186;
wire v_14187;
wire v_14188;
wire v_14189;
wire v_14190;
wire v_14191;
wire v_14192;
wire v_14193;
wire v_14194;
wire v_14195;
wire v_14196;
wire v_14197;
wire v_14198;
wire v_14199;
wire v_14200;
wire v_14201;
wire v_14202;
wire v_14203;
wire v_14204;
wire v_14205;
wire v_14206;
wire v_14207;
wire v_14208;
wire v_14209;
wire v_14210;
wire v_14211;
wire v_14212;
wire v_14213;
wire v_14214;
wire v_14215;
wire v_14216;
wire v_14217;
wire v_14218;
wire v_14219;
wire v_14220;
wire v_14221;
wire v_14222;
wire v_14223;
wire v_14224;
wire v_14225;
wire v_14226;
wire v_14227;
wire v_14228;
wire v_14229;
wire v_14230;
wire v_14231;
wire v_14232;
wire v_14233;
wire v_14234;
wire v_14235;
wire v_14236;
wire v_14237;
wire v_14238;
wire v_14239;
wire v_14240;
wire v_14241;
wire v_14242;
wire v_14243;
wire v_14244;
wire v_14245;
wire v_14246;
wire v_14247;
wire v_14248;
wire v_14249;
wire v_14250;
wire v_14251;
wire v_14252;
wire v_14253;
wire v_14254;
wire v_14255;
wire v_14256;
wire v_14257;
wire v_14258;
wire v_14259;
wire v_14260;
wire v_14261;
wire v_14262;
wire v_14263;
wire v_14264;
wire v_14265;
wire v_14266;
wire v_14267;
wire v_14268;
wire v_14269;
wire v_14270;
wire v_14271;
wire v_14272;
wire v_14273;
wire v_14274;
wire v_14275;
wire v_14276;
wire v_14277;
wire v_14278;
wire v_14279;
wire v_14280;
wire v_14281;
wire v_14282;
wire v_14283;
wire v_14284;
wire v_14285;
wire v_14286;
wire v_14287;
wire v_14288;
wire v_14289;
wire v_14290;
wire v_14291;
wire v_14292;
wire v_14293;
wire v_14294;
wire v_14295;
wire v_14296;
wire v_14297;
wire v_14298;
wire v_14299;
wire v_14300;
wire v_14301;
wire v_14302;
wire v_14303;
wire v_14304;
wire v_14305;
wire v_14306;
wire v_14307;
wire v_14308;
wire v_14309;
wire v_14310;
wire v_14311;
wire v_14312;
wire v_14313;
wire v_14314;
wire v_14315;
wire v_14316;
wire v_14317;
wire v_14318;
wire v_14319;
wire v_14320;
wire v_14321;
wire v_14322;
wire v_14323;
wire v_14324;
wire v_14325;
wire v_14326;
wire v_14327;
wire v_14328;
wire v_14329;
wire v_14330;
wire v_14331;
wire v_14332;
wire v_14333;
wire v_14334;
wire v_14335;
wire v_14336;
wire v_14337;
wire v_14338;
wire v_14339;
wire v_14340;
wire v_14341;
wire v_14342;
wire v_14343;
wire v_14344;
wire v_14345;
wire v_14346;
wire v_14347;
wire v_14348;
wire v_14349;
wire v_14350;
wire v_14351;
wire v_14352;
wire v_14353;
wire v_14354;
wire v_14355;
wire v_14356;
wire v_14357;
wire v_14358;
wire v_14359;
wire v_14360;
wire v_14361;
wire v_14362;
wire v_14363;
wire v_14364;
wire v_14365;
wire v_14366;
wire v_14367;
wire v_14368;
wire v_14369;
wire v_14370;
wire v_14371;
wire v_14372;
wire v_14373;
wire v_14374;
wire v_14375;
wire v_14376;
wire v_14377;
wire v_14378;
wire v_14379;
wire v_14380;
wire v_14381;
wire v_14382;
wire v_14383;
wire v_14384;
wire v_14385;
wire v_14386;
wire v_14387;
wire v_14388;
wire v_14389;
wire v_14390;
wire v_14391;
wire v_14392;
wire v_14393;
wire v_14394;
wire v_14395;
wire v_14396;
wire v_14397;
wire v_14398;
wire v_14399;
wire v_14400;
wire v_14401;
wire v_14402;
wire v_14403;
wire v_14404;
wire v_14405;
wire v_14406;
wire v_14407;
wire v_14408;
wire v_14409;
wire v_14410;
wire v_14411;
wire v_14412;
wire v_14413;
wire v_14414;
wire v_14415;
wire v_14416;
wire v_14417;
wire v_14418;
wire v_14419;
wire v_14420;
wire v_14421;
wire v_14422;
wire v_14423;
wire v_14424;
wire v_14425;
wire v_14426;
wire v_14427;
wire v_14428;
wire v_14429;
wire v_14430;
wire v_14431;
wire v_14432;
wire v_14433;
wire v_14434;
wire v_14435;
wire v_14436;
wire v_14437;
wire v_14438;
wire v_14439;
wire v_14440;
wire v_14441;
wire v_14442;
wire v_14443;
wire v_14444;
wire v_14445;
wire v_14446;
wire v_14447;
wire v_14448;
wire v_14449;
wire v_14450;
wire v_14451;
wire v_14452;
wire v_14453;
wire v_14454;
wire v_14455;
wire v_14456;
wire v_14457;
wire v_14458;
wire v_14459;
wire v_14460;
wire v_14461;
wire v_14462;
wire v_14463;
wire v_14464;
wire v_14465;
wire v_14466;
wire v_14467;
wire v_14468;
wire v_14469;
wire v_14470;
wire v_14471;
wire v_14472;
wire v_14473;
wire v_14474;
wire v_14475;
wire v_14476;
wire v_14477;
wire v_14478;
wire v_14479;
wire v_14480;
wire v_14481;
wire v_14482;
wire v_14483;
wire v_14484;
wire v_14485;
wire v_14486;
wire v_14487;
wire v_14488;
wire v_14489;
wire v_14490;
wire v_14491;
wire v_14492;
wire v_14493;
wire v_14494;
wire v_14495;
wire v_14496;
wire v_14497;
wire v_14498;
wire v_14499;
wire v_14500;
wire v_14501;
wire v_14502;
wire v_14503;
wire v_14504;
wire v_14505;
wire v_14506;
wire v_14507;
wire v_14508;
wire v_14509;
wire v_14510;
wire v_14511;
wire v_14512;
wire v_14513;
wire v_14514;
wire v_14515;
wire v_14516;
wire v_14517;
wire v_14518;
wire v_14519;
wire v_14520;
wire v_14521;
wire v_14522;
wire v_14523;
wire v_14524;
wire v_14525;
wire v_14526;
wire v_14527;
wire v_14528;
wire v_14529;
wire v_14530;
wire v_14531;
wire v_14532;
wire v_14533;
wire v_14534;
wire v_14535;
wire v_14536;
wire v_14537;
wire v_14538;
wire v_14539;
wire v_14540;
wire v_14541;
wire v_14542;
wire v_14543;
wire v_14544;
wire v_14545;
wire v_14546;
wire v_14547;
wire v_14548;
wire v_14549;
wire v_14550;
wire v_14551;
wire v_14552;
wire v_14553;
wire v_14554;
wire v_14555;
wire v_14556;
wire v_14557;
wire v_14558;
wire v_14559;
wire v_14560;
wire v_14561;
wire v_14562;
wire v_14563;
wire v_14564;
wire v_14565;
wire v_14566;
wire v_14567;
wire v_14568;
wire v_14569;
wire v_14570;
wire v_14571;
wire v_14572;
wire v_14573;
wire v_14574;
wire v_14575;
wire v_14576;
wire v_14577;
wire v_14578;
wire v_14579;
wire v_14580;
wire v_14581;
wire v_14582;
wire v_14583;
wire v_14584;
wire v_14585;
wire v_14586;
wire v_14587;
wire v_14588;
wire v_14589;
wire v_14590;
wire v_14591;
wire v_14592;
wire v_14593;
wire v_14594;
wire v_14595;
wire v_14596;
wire v_14597;
wire v_14598;
wire v_14599;
wire v_14600;
wire v_14601;
wire v_14602;
wire v_14603;
wire v_14604;
wire v_14605;
wire v_14606;
wire v_14607;
wire v_14608;
wire v_14609;
wire v_14610;
wire v_14611;
wire v_14612;
wire v_14613;
wire v_14614;
wire v_14615;
wire v_14616;
wire v_14617;
wire v_14618;
wire v_14619;
wire v_14620;
wire v_14621;
wire v_14622;
wire v_14623;
wire v_14624;
wire v_14625;
wire v_14626;
wire v_14627;
wire v_14628;
wire v_14629;
wire v_14630;
wire v_14631;
wire v_14632;
wire v_14633;
wire v_14634;
wire v_14635;
wire v_14636;
wire v_14637;
wire v_14638;
wire v_14639;
wire v_14640;
wire v_14641;
wire v_14642;
wire v_14643;
wire v_14644;
wire v_14645;
wire v_14646;
wire v_14647;
wire v_14648;
wire v_14649;
wire v_14650;
wire v_14651;
wire v_14652;
wire v_14653;
wire v_14654;
wire v_14655;
wire v_14656;
wire v_14657;
wire v_14658;
wire v_14659;
wire v_14660;
wire v_14661;
wire v_14662;
wire v_14663;
wire v_14664;
wire v_14665;
wire v_14666;
wire v_14667;
wire v_14668;
wire v_14669;
wire v_14670;
wire v_14671;
wire v_14672;
wire v_14673;
wire v_14674;
wire v_14675;
wire v_14676;
wire v_14677;
wire v_14678;
wire v_14679;
wire v_14680;
wire v_14681;
wire v_14682;
wire v_14683;
wire v_14684;
wire v_14685;
wire v_14686;
wire v_14687;
wire v_14688;
wire v_14689;
wire v_14690;
wire v_14691;
wire v_14692;
wire v_14693;
wire v_14694;
wire v_14695;
wire v_14696;
wire v_14697;
wire v_14698;
wire v_14699;
wire v_14700;
wire v_14701;
wire v_14702;
wire v_14703;
wire v_14704;
wire v_14705;
wire v_14706;
wire v_14707;
wire v_14708;
wire v_14709;
wire v_14710;
wire v_14711;
wire v_14712;
wire v_14713;
wire v_14714;
wire v_14715;
wire v_14716;
wire v_14717;
wire v_14718;
wire v_14719;
wire v_14720;
wire v_14721;
wire v_14722;
wire v_14723;
wire v_14724;
wire v_14725;
wire v_14726;
wire v_14727;
wire v_14728;
wire v_14729;
wire v_14730;
wire v_14731;
wire v_14732;
wire v_14733;
wire v_14734;
wire v_14735;
wire v_14736;
wire v_14737;
wire v_14738;
wire v_14739;
wire v_14740;
wire v_14741;
wire v_14742;
wire v_14743;
wire v_14744;
wire v_14745;
wire v_14746;
wire v_14747;
wire v_14748;
wire v_14749;
wire v_14750;
wire v_14751;
wire v_14752;
wire v_14753;
wire v_14754;
wire v_14755;
wire v_14756;
wire v_14757;
wire v_14758;
wire v_14759;
wire v_14760;
wire v_14761;
wire v_14762;
wire v_14763;
wire v_14764;
wire v_14765;
wire v_14766;
wire v_14767;
wire v_14768;
wire v_14769;
wire v_14770;
wire v_14771;
wire v_14772;
wire v_14773;
wire v_14774;
wire v_14775;
wire v_14776;
wire v_14777;
wire v_14778;
wire v_14779;
wire v_14780;
wire v_14781;
wire v_14782;
wire v_14783;
wire v_14784;
wire v_14785;
wire v_14786;
wire v_14787;
wire v_14788;
wire v_14789;
wire v_14790;
wire v_14791;
wire v_14792;
wire v_14793;
wire v_14794;
wire v_14795;
wire v_14796;
wire v_14797;
wire v_14798;
wire v_14799;
wire v_14800;
wire v_14801;
wire v_14802;
wire v_14803;
wire v_14804;
wire v_14805;
wire v_14806;
wire v_14807;
wire v_14808;
wire v_14809;
wire v_14810;
wire v_14811;
wire v_14812;
wire v_14813;
wire v_14814;
wire v_14815;
wire v_14816;
wire v_14817;
wire v_14818;
wire v_14819;
wire v_14820;
wire v_14821;
wire v_14822;
wire v_14823;
wire v_14824;
wire v_14825;
wire v_14826;
wire v_14827;
wire v_14828;
wire v_14829;
wire v_14830;
wire v_14831;
wire v_14832;
wire v_14833;
wire v_14834;
wire v_14835;
wire v_14836;
wire v_14837;
wire v_14838;
wire v_14839;
wire v_14840;
wire v_14841;
wire v_14842;
wire v_14843;
wire v_14844;
wire v_14845;
wire v_14846;
wire v_14847;
wire v_14848;
wire v_14849;
wire v_14850;
wire v_14851;
wire v_14852;
wire v_14853;
wire v_14854;
wire v_14855;
wire v_14856;
wire v_14857;
wire v_14858;
wire v_14859;
wire v_14860;
wire v_14861;
wire v_14862;
wire v_14863;
wire v_14864;
wire v_14865;
wire v_14866;
wire v_14867;
wire v_14868;
wire v_14869;
wire v_14870;
wire v_14871;
wire v_14872;
wire v_14873;
wire v_14874;
wire v_14875;
wire v_14876;
wire v_14877;
wire v_14878;
wire v_14879;
wire v_14880;
wire v_14881;
wire v_14882;
wire v_14883;
wire v_14884;
wire v_14885;
wire v_14886;
wire v_14887;
wire v_14888;
wire v_14889;
wire v_14890;
wire v_14891;
wire v_14892;
wire v_14893;
wire v_14894;
wire v_14895;
wire v_14896;
wire v_14897;
wire v_14898;
wire v_14899;
wire v_14900;
wire v_14901;
wire v_14902;
wire v_14903;
wire v_14904;
wire v_14905;
wire v_14906;
wire v_14907;
wire v_14908;
wire v_14909;
wire v_14910;
wire v_14911;
wire v_14912;
wire v_14913;
wire v_14914;
wire v_14915;
wire v_14916;
wire v_14917;
wire v_14918;
wire v_14919;
wire v_14920;
wire v_14921;
wire v_14922;
wire v_14923;
wire v_14924;
wire v_14925;
wire v_14926;
wire v_14927;
wire v_14928;
wire v_14929;
wire v_14930;
wire v_14931;
wire v_14932;
wire v_14933;
wire v_14934;
wire v_14935;
wire v_14936;
wire v_14937;
wire v_14938;
wire v_14939;
wire v_14940;
wire v_14941;
wire v_14942;
wire v_14943;
wire v_14944;
wire v_14945;
wire v_14946;
wire v_14947;
wire v_14948;
wire v_14949;
wire v_14950;
wire v_14951;
wire v_14952;
wire v_14953;
wire v_14954;
wire v_14955;
wire v_14956;
wire v_14957;
wire v_14958;
wire v_14959;
wire v_14960;
wire v_14961;
wire v_14962;
wire v_14963;
wire v_14964;
wire v_14965;
wire v_14966;
wire v_14967;
wire v_14968;
wire v_14969;
wire v_14970;
wire v_14971;
wire v_14972;
wire v_14973;
wire v_14974;
wire v_14975;
wire v_14976;
wire v_14977;
wire v_14978;
wire v_14979;
wire v_14980;
wire v_14981;
wire v_14982;
wire v_14983;
wire v_14984;
wire v_14985;
wire v_14986;
wire v_14987;
wire v_14988;
wire v_14989;
wire v_14990;
wire v_14991;
wire v_14992;
wire v_14993;
wire v_14994;
wire v_14995;
wire v_14996;
wire v_14997;
wire v_14998;
wire v_14999;
wire v_15000;
wire v_15001;
wire v_15002;
wire v_15003;
wire v_15004;
wire v_15005;
wire v_15006;
wire v_15007;
wire v_15008;
wire v_15009;
wire v_15010;
wire v_15011;
wire v_15012;
wire v_15013;
wire v_15014;
wire v_15015;
wire v_15016;
wire v_15017;
wire v_15018;
wire v_15019;
wire v_15020;
wire v_15021;
wire v_15022;
wire v_15023;
wire v_15024;
wire v_15025;
wire v_15026;
wire v_15027;
wire v_15028;
wire v_15029;
wire v_15030;
wire v_15031;
wire v_15032;
wire v_15033;
wire v_15034;
wire v_15035;
wire v_15036;
wire v_15037;
wire v_15038;
wire v_15039;
wire v_15040;
wire v_15041;
wire v_15042;
wire v_15043;
wire v_15044;
wire v_15045;
wire v_15046;
wire v_15047;
wire v_15048;
wire v_15049;
wire v_15050;
wire v_15051;
wire v_15052;
wire v_15053;
wire v_15054;
wire v_15055;
wire v_15056;
wire v_15057;
wire v_15058;
wire v_15059;
wire v_15060;
wire v_15061;
wire v_15062;
wire v_15063;
wire v_15064;
wire v_15065;
wire v_15066;
wire v_15067;
wire v_15068;
wire v_15069;
wire v_15070;
wire v_15071;
wire v_15072;
wire v_15073;
wire v_15074;
wire v_15075;
wire v_15076;
wire v_15077;
wire v_15078;
wire v_15079;
wire v_15080;
wire v_15081;
wire v_15082;
wire v_15083;
wire v_15084;
wire v_15085;
wire v_15086;
wire v_15087;
wire v_15088;
wire v_15089;
wire v_15090;
wire v_15091;
wire v_15092;
wire v_15093;
wire v_15094;
wire v_15095;
wire v_15096;
wire v_15097;
wire v_15098;
wire v_15099;
wire v_15100;
wire v_15101;
wire v_15102;
wire v_15103;
wire v_15104;
wire v_15105;
wire v_15106;
wire v_15107;
wire v_15108;
wire v_15109;
wire v_15110;
wire v_15111;
wire v_15112;
wire v_15113;
wire v_15114;
wire v_15115;
wire v_15116;
wire v_15117;
wire v_15118;
wire v_15119;
wire v_15120;
wire v_15121;
wire v_15122;
wire v_15123;
wire v_15124;
wire v_15125;
wire v_15126;
wire v_15127;
wire v_15128;
wire v_15129;
wire v_15130;
wire v_15131;
wire v_15132;
wire v_15133;
wire v_15134;
wire v_15135;
wire v_15136;
wire v_15137;
wire v_15138;
wire v_15139;
wire v_15140;
wire v_15141;
wire v_15142;
wire v_15143;
wire v_15144;
wire v_15145;
wire v_15146;
wire v_15147;
wire v_15148;
wire v_15149;
wire v_15150;
wire v_15151;
wire v_15152;
wire v_15153;
wire v_15154;
wire v_15155;
wire v_15156;
wire v_15157;
wire v_15158;
wire v_15159;
wire v_15160;
wire v_15161;
wire v_15162;
wire v_15163;
wire v_15164;
wire v_15165;
wire v_15166;
wire v_15167;
wire v_15168;
wire v_15169;
wire v_15170;
wire v_15171;
wire v_15172;
wire v_15173;
wire v_15174;
wire v_15175;
wire v_15176;
wire v_15177;
wire v_15178;
wire v_15179;
wire v_15180;
wire v_15181;
wire v_15182;
wire v_15183;
wire v_15184;
wire v_15185;
wire v_15186;
wire v_15187;
wire v_15188;
wire v_15189;
wire v_15190;
wire v_15191;
wire v_15192;
wire v_15193;
wire v_15194;
wire v_15195;
wire v_15196;
wire v_15197;
wire v_15198;
wire v_15199;
wire v_15200;
wire v_15201;
wire v_15202;
wire v_15203;
wire v_15204;
wire v_15205;
wire v_15206;
wire v_15207;
wire v_15208;
wire v_15209;
wire v_15210;
wire v_15211;
wire v_15212;
wire v_15213;
wire v_15214;
wire v_15215;
wire v_15216;
wire v_15217;
wire v_15218;
wire v_15219;
wire v_15220;
wire v_15221;
wire v_15222;
wire v_15223;
wire v_15224;
wire v_15225;
wire v_15226;
wire v_15227;
wire v_15228;
wire v_15229;
wire v_15230;
wire v_15231;
wire v_15232;
wire v_15233;
wire v_15234;
wire v_15235;
wire v_15236;
wire v_15237;
wire v_15238;
wire v_15239;
wire v_15240;
wire v_15241;
wire v_15242;
wire v_15243;
wire v_15244;
wire v_15245;
wire v_15246;
wire v_15247;
wire v_15248;
wire v_15249;
wire v_15250;
wire v_15251;
wire v_15252;
wire v_15253;
wire v_15254;
wire v_15255;
wire v_15256;
wire v_15257;
wire v_15258;
wire v_15259;
wire v_15260;
wire v_15261;
wire v_15262;
wire v_15263;
wire v_15264;
wire v_15265;
wire v_15266;
wire v_15267;
wire v_15268;
wire v_15269;
wire v_15270;
wire v_15271;
wire v_15272;
wire v_15273;
wire v_15274;
wire v_15275;
wire v_15276;
wire v_15277;
wire v_15278;
wire v_15279;
wire v_15280;
wire v_15281;
wire v_15282;
wire v_15283;
wire v_15284;
wire v_15285;
wire v_15286;
wire v_15287;
wire v_15288;
wire v_15289;
wire v_15290;
wire v_15291;
wire v_15292;
wire v_15293;
wire v_15294;
wire v_15295;
wire v_15296;
wire v_15297;
wire v_15298;
wire v_15299;
wire v_15300;
wire v_15301;
wire v_15302;
wire v_15303;
wire v_15304;
wire v_15305;
wire v_15306;
wire v_15307;
wire v_15308;
wire v_15309;
wire v_15310;
wire v_15311;
wire v_15312;
wire v_15313;
wire v_15314;
wire v_15315;
wire v_15316;
wire v_15317;
wire v_15318;
wire v_15319;
wire v_15320;
wire v_15321;
wire v_15322;
wire v_15323;
wire v_15324;
wire v_15325;
wire v_15326;
wire v_15327;
wire v_15328;
wire v_15329;
wire v_15330;
wire v_15331;
wire v_15332;
wire v_15333;
wire v_15334;
wire v_15335;
wire v_15336;
wire v_15337;
wire v_15338;
wire v_15339;
wire v_15340;
wire v_15341;
wire v_15342;
wire v_15343;
wire v_15344;
wire v_15345;
wire v_15346;
wire v_15347;
wire v_15348;
wire v_15349;
wire v_15350;
wire v_15351;
wire v_15352;
wire v_15353;
wire v_15354;
wire v_15355;
wire v_15356;
wire v_15357;
wire v_15358;
wire v_15359;
wire v_15360;
wire v_15361;
wire v_15362;
wire v_15363;
wire v_15364;
wire v_15365;
wire v_15366;
wire v_15367;
wire v_15368;
wire v_15369;
wire v_15370;
wire v_15371;
wire v_15372;
wire v_15373;
wire v_15374;
wire v_15375;
wire v_15376;
wire v_15377;
wire v_15378;
wire v_15379;
wire v_15380;
wire v_15381;
wire v_15382;
wire v_15383;
wire v_15384;
wire v_15385;
wire v_15386;
wire v_15387;
wire v_15388;
wire v_15389;
wire v_15390;
wire v_15391;
wire v_15392;
wire v_15393;
wire v_15394;
wire v_15395;
wire v_15396;
wire v_15397;
wire v_15398;
wire v_15399;
wire v_15400;
wire v_15401;
wire v_15402;
wire v_15403;
wire v_15404;
wire v_15405;
wire v_15406;
wire v_15407;
wire v_15408;
wire v_15409;
wire v_15410;
wire v_15411;
wire v_15412;
wire v_15413;
wire v_15414;
wire v_15415;
wire v_15416;
wire v_15417;
wire v_15418;
wire v_15419;
wire v_15420;
wire v_15421;
wire v_15422;
wire v_15423;
wire v_15424;
wire v_15425;
wire v_15426;
wire v_15427;
wire v_15428;
wire v_15429;
wire v_15430;
wire v_15431;
wire v_15432;
wire v_15433;
wire v_15434;
wire v_15435;
wire v_15436;
wire v_15437;
wire v_15438;
wire v_15439;
wire v_15440;
wire v_15441;
wire v_15442;
wire v_15443;
wire v_15444;
wire v_15445;
wire v_15446;
wire v_15447;
wire v_15448;
wire v_15449;
wire v_15450;
wire v_15451;
wire v_15452;
wire v_15453;
wire v_15454;
wire v_15455;
wire v_15456;
wire v_15457;
wire v_15458;
wire v_15459;
wire v_15460;
wire v_15461;
wire v_15462;
wire v_15463;
wire v_15464;
wire v_15465;
wire v_15466;
wire v_15467;
wire v_15468;
wire v_15469;
wire v_15470;
wire v_15471;
wire v_15472;
wire v_15473;
wire v_15474;
wire v_15475;
wire v_15476;
wire v_15477;
wire v_15478;
wire v_15479;
wire v_15480;
wire v_15481;
wire v_15482;
wire v_15483;
wire v_15484;
wire v_15485;
wire v_15486;
wire v_15487;
wire v_15488;
wire v_15489;
wire v_15490;
wire v_15491;
wire v_15492;
wire v_15493;
wire v_15494;
wire v_15495;
wire v_15496;
wire v_15497;
wire v_15498;
wire v_15499;
wire v_15500;
wire v_15501;
wire v_15502;
wire v_15503;
wire v_15504;
wire v_15505;
wire v_15506;
wire v_15507;
wire v_15508;
wire v_15509;
wire v_15510;
wire v_15511;
wire v_15512;
wire v_15513;
wire v_15514;
wire v_15515;
wire v_15516;
wire v_15517;
wire v_15518;
wire v_15519;
wire v_15520;
wire v_15521;
wire v_15522;
wire v_15523;
wire v_15524;
wire v_15525;
wire v_15526;
wire v_15527;
wire v_15528;
wire v_15529;
wire v_15530;
wire v_15531;
wire v_15532;
wire v_15533;
wire v_15534;
wire v_15535;
wire v_15536;
wire v_15537;
wire v_15538;
wire v_15539;
wire v_15540;
wire v_15541;
wire v_15542;
wire v_15543;
wire v_15544;
wire v_15545;
wire v_15546;
wire v_15547;
wire v_15548;
wire v_15549;
wire v_15550;
wire v_15551;
wire v_15552;
wire v_15553;
wire v_15554;
wire v_15555;
wire v_15556;
wire v_15557;
wire v_15558;
wire v_15559;
wire v_15560;
wire v_15561;
wire v_15562;
wire v_15563;
wire v_15564;
wire v_15565;
wire v_15566;
wire v_15567;
wire v_15568;
wire v_15569;
wire v_15570;
wire v_15571;
wire v_15572;
wire v_15573;
wire v_15574;
wire v_15575;
wire v_15576;
wire v_15577;
wire v_15578;
wire v_15579;
wire v_15580;
wire v_15581;
wire v_15582;
wire v_15583;
wire v_15584;
wire v_15585;
wire v_15586;
wire v_15587;
wire v_15588;
wire v_15589;
wire v_15590;
wire v_15591;
wire v_15592;
wire v_15593;
wire v_15594;
wire v_15595;
wire v_15596;
wire v_15597;
wire v_15598;
wire v_15599;
wire v_15600;
wire v_15601;
wire v_15602;
wire v_15603;
wire v_15604;
wire v_15605;
wire v_15606;
wire v_15607;
wire v_15608;
wire v_15609;
wire v_15610;
wire v_15611;
wire v_15612;
wire v_15613;
wire v_15614;
wire v_15615;
wire v_15616;
wire v_15617;
wire v_15618;
wire v_15619;
wire v_15620;
wire v_15621;
wire v_15622;
wire v_15623;
wire v_15624;
wire v_15625;
wire v_15626;
wire v_15627;
wire v_15628;
wire v_15629;
wire v_15630;
wire v_15631;
wire v_15632;
wire v_15633;
wire v_15634;
wire v_15635;
wire v_15636;
wire v_15637;
wire v_15638;
wire v_15639;
wire v_15640;
wire v_15641;
wire v_15642;
wire v_15643;
wire v_15644;
wire v_15645;
wire v_15646;
wire v_15647;
wire v_15648;
wire v_15649;
wire v_15650;
wire v_15651;
wire v_15652;
wire v_15653;
wire v_15654;
wire v_15655;
wire v_15656;
wire v_15657;
wire v_15658;
wire v_15659;
wire v_15660;
wire v_15661;
wire v_15662;
wire v_15663;
wire v_15664;
wire v_15665;
wire v_15666;
wire v_15667;
wire v_15668;
wire v_15669;
wire v_15670;
wire v_15671;
wire v_15672;
wire v_15673;
wire v_15674;
wire v_15675;
wire v_15676;
wire v_15677;
wire v_15678;
wire v_15679;
wire v_15680;
wire v_15681;
wire v_15682;
wire v_15683;
wire v_15684;
wire v_15685;
wire v_15686;
wire v_15687;
wire v_15688;
wire v_15689;
wire v_15690;
wire v_15691;
wire v_15692;
wire v_15693;
wire v_15694;
wire v_15695;
wire v_15696;
wire v_15697;
wire v_15698;
wire v_15699;
wire v_15700;
wire v_15701;
wire v_15702;
wire v_15703;
wire v_15704;
wire v_15705;
wire v_15706;
wire v_15707;
wire v_15708;
wire v_15709;
wire v_15710;
wire v_15711;
wire v_15712;
wire v_15713;
wire v_15714;
wire v_15715;
wire v_15716;
wire v_15717;
wire v_15718;
wire v_15719;
wire v_15720;
wire v_15721;
wire v_15722;
wire v_15723;
wire v_15724;
wire v_15725;
wire v_15726;
wire v_15727;
wire v_15728;
wire v_15729;
wire v_15730;
wire v_15731;
wire v_15732;
wire v_15733;
wire v_15734;
wire v_15735;
wire v_15736;
wire v_15737;
wire v_15738;
wire v_15739;
wire v_15740;
wire v_15741;
wire v_15742;
wire v_15743;
wire v_15744;
wire v_15745;
wire v_15746;
wire v_15747;
wire v_15748;
wire v_15749;
wire v_15750;
wire v_15751;
wire v_15752;
wire v_15753;
wire v_15754;
wire v_15755;
wire v_15756;
wire v_15757;
wire v_15758;
wire v_15759;
wire v_15760;
wire v_15761;
wire v_15762;
wire v_15763;
wire v_15764;
wire v_15765;
wire v_15766;
wire v_15767;
wire v_15768;
wire v_15769;
wire v_15770;
wire v_15771;
wire v_15772;
wire v_15773;
wire v_15774;
wire v_15775;
wire v_15776;
wire v_15777;
wire v_15778;
wire v_15779;
wire v_15780;
wire v_15781;
wire v_15782;
wire v_15783;
wire v_15784;
wire v_15785;
wire v_15786;
wire v_15787;
wire v_15788;
wire v_15789;
wire v_15790;
wire v_15791;
wire v_15792;
wire v_15793;
wire v_15794;
wire v_15795;
wire v_15796;
wire v_15797;
wire v_15798;
wire v_15799;
wire v_15800;
wire v_15801;
wire v_15802;
wire v_15803;
wire v_15804;
wire v_15805;
wire v_15806;
wire v_15807;
wire v_15808;
wire v_15809;
wire v_15810;
wire v_15811;
wire v_15812;
wire v_15813;
wire v_15814;
wire v_15815;
wire v_15816;
wire v_15817;
wire v_15818;
wire v_15819;
wire v_15820;
wire v_15821;
wire v_15822;
wire v_15823;
wire v_15824;
wire v_15825;
wire v_15826;
wire v_15827;
wire v_15828;
wire v_15829;
wire v_15830;
wire v_15831;
wire v_15832;
wire v_15833;
wire v_15834;
wire v_15835;
wire v_15836;
wire v_15837;
wire v_15838;
wire v_15839;
wire v_15840;
wire v_15841;
wire v_15842;
wire v_15843;
wire v_15844;
wire v_15845;
wire v_15846;
wire v_15847;
wire v_15848;
wire v_15849;
wire v_15850;
wire v_15851;
wire v_15852;
wire v_15853;
wire v_15854;
wire v_15855;
wire v_15856;
wire v_15857;
wire v_15858;
wire v_15859;
wire v_15860;
wire v_15861;
wire v_15862;
wire v_15863;
wire v_15864;
wire v_15865;
wire v_15866;
wire v_15867;
wire v_15868;
wire v_15869;
wire v_15870;
wire v_15871;
wire v_15872;
wire v_15873;
wire v_15874;
wire v_15875;
wire v_15876;
wire v_15877;
wire v_15878;
wire v_15879;
wire v_15880;
wire v_15881;
wire v_15882;
wire v_15883;
wire v_15884;
wire v_15885;
wire v_15886;
wire v_15887;
wire v_15888;
wire v_15889;
wire v_15890;
wire v_15891;
wire v_15892;
wire v_15893;
wire v_15894;
wire v_15895;
wire v_15896;
wire v_15897;
wire v_15898;
wire v_15899;
wire v_15900;
wire v_15901;
wire v_15902;
wire v_15903;
wire v_15904;
wire v_15905;
wire v_15906;
wire v_15907;
wire v_15908;
wire v_15909;
wire v_15910;
wire v_15911;
wire v_15912;
wire v_15913;
wire v_15914;
wire v_15915;
wire v_15916;
wire v_15917;
wire v_15918;
wire v_15919;
wire v_15920;
wire v_15921;
wire v_15922;
wire v_15923;
wire v_15924;
wire v_15925;
wire v_15926;
wire v_15927;
wire v_15928;
wire v_15929;
wire v_15930;
wire v_15931;
wire v_15932;
wire v_15933;
wire v_15934;
wire v_15935;
wire v_15936;
wire v_15937;
wire v_15938;
wire v_15939;
wire v_15940;
wire v_15941;
wire v_15942;
wire v_15943;
wire v_15944;
wire v_15945;
wire v_15946;
wire v_15947;
wire v_15948;
wire v_15949;
wire v_15950;
wire v_15951;
wire v_15952;
wire v_15953;
wire v_15954;
wire v_15955;
wire v_15956;
wire v_15957;
wire v_15958;
wire v_15959;
wire v_15960;
wire v_15961;
wire v_15962;
wire v_15963;
wire v_15964;
wire v_15965;
wire v_15966;
wire v_15967;
wire v_15968;
wire v_15969;
wire v_15970;
wire v_15971;
wire v_15972;
wire v_15973;
wire v_15974;
wire v_15975;
wire v_15976;
wire v_15977;
wire v_15978;
wire v_15979;
wire v_15980;
wire v_15981;
wire v_15982;
wire v_15983;
wire v_15984;
wire v_15985;
wire v_15986;
wire v_15987;
wire v_15988;
wire v_15989;
wire v_15990;
wire v_15991;
wire v_15992;
wire v_15993;
wire v_15994;
wire v_15995;
wire v_15996;
wire v_15997;
wire v_15998;
wire v_15999;
wire v_16000;
wire v_16001;
wire v_16002;
wire v_16003;
wire v_16004;
wire v_16005;
wire v_16006;
wire v_16007;
wire v_16008;
wire v_16009;
wire v_16010;
wire v_16011;
wire v_16012;
wire v_16013;
wire v_16014;
wire v_16015;
wire v_16016;
wire v_16017;
wire v_16018;
wire v_16019;
wire v_16020;
wire v_16021;
wire v_16022;
wire v_16023;
wire v_16024;
wire v_16025;
wire v_16026;
wire v_16027;
wire v_16028;
wire v_16029;
wire v_16030;
wire v_16031;
wire v_16032;
wire v_16033;
wire v_16034;
wire v_16035;
wire v_16036;
wire v_16037;
wire v_16038;
wire v_16039;
wire v_16040;
wire v_16041;
wire v_16042;
wire v_16043;
wire v_16044;
wire v_16045;
wire v_16046;
wire v_16047;
wire v_16048;
wire v_16049;
wire v_16050;
wire v_16051;
wire v_16052;
wire v_16053;
wire v_16054;
wire v_16055;
wire v_16056;
wire v_16057;
wire v_16058;
wire v_16059;
wire v_16060;
wire v_16061;
wire v_16062;
wire v_16063;
wire v_16064;
wire v_16065;
wire v_16066;
wire v_16067;
wire v_16068;
wire v_16069;
wire v_16070;
wire v_16071;
wire v_16072;
wire v_16073;
wire v_16074;
wire v_16075;
wire v_16076;
wire v_16077;
wire v_16078;
wire v_16079;
wire v_16080;
wire v_16081;
wire v_16082;
wire v_16083;
wire v_16084;
wire v_16085;
wire v_16086;
wire v_16087;
wire v_16088;
wire v_16089;
wire v_16090;
wire v_16091;
wire v_16092;
wire v_16093;
wire v_16094;
wire v_16095;
wire v_16096;
wire v_16097;
wire v_16098;
wire v_16099;
wire v_16100;
wire v_16101;
wire v_16102;
wire v_16103;
wire v_16104;
wire v_16105;
wire v_16106;
wire v_16107;
wire v_16108;
wire v_16109;
wire v_16110;
wire v_16111;
wire v_16112;
wire v_16113;
wire v_16114;
wire v_16115;
wire v_16116;
wire v_16117;
wire v_16118;
wire v_16119;
wire v_16120;
wire v_16121;
wire v_16122;
wire v_16123;
wire v_16124;
wire v_16125;
wire v_16126;
wire v_16127;
wire v_16128;
wire v_16129;
wire v_16130;
wire v_16131;
wire v_16132;
wire v_16133;
wire v_16134;
wire v_16135;
wire v_16136;
wire v_16137;
wire v_16138;
wire v_16139;
wire v_16140;
wire v_16141;
wire v_16142;
wire v_16143;
wire v_16144;
wire v_16145;
wire v_16146;
wire v_16147;
wire v_16148;
wire v_16149;
wire v_16150;
wire v_16151;
wire v_16152;
wire v_16153;
wire v_16154;
wire v_16155;
wire v_16156;
wire v_16157;
wire v_16158;
wire v_16159;
wire v_16160;
wire v_16161;
wire v_16162;
wire v_16163;
wire v_16164;
wire v_16165;
wire v_16166;
wire v_16167;
wire v_16168;
wire v_16169;
wire v_16170;
wire v_16171;
wire v_16172;
wire v_16173;
wire v_16174;
wire v_16175;
wire v_16176;
wire v_16177;
wire v_16178;
wire v_16179;
wire v_16180;
wire v_16181;
wire v_16182;
wire v_16183;
wire v_16184;
wire v_16185;
wire v_16186;
wire v_16187;
wire v_16188;
wire v_16189;
wire v_16190;
wire v_16191;
wire v_16192;
wire v_16193;
wire v_16194;
wire v_16195;
wire v_16196;
wire v_16197;
wire v_16198;
wire v_16199;
wire v_16200;
wire v_16201;
wire v_16202;
wire v_16203;
wire v_16204;
wire v_16205;
wire v_16206;
wire v_16207;
wire v_16208;
wire v_16209;
wire v_16210;
wire v_16211;
wire v_16212;
wire v_16213;
wire v_16214;
wire v_16215;
wire v_16216;
wire v_16217;
wire v_16218;
wire v_16219;
wire v_16220;
wire v_16221;
wire v_16222;
wire v_16223;
wire v_16224;
wire v_16225;
wire v_16226;
wire v_16227;
wire v_16228;
wire v_16229;
wire v_16230;
wire v_16231;
wire v_16232;
wire v_16233;
wire v_16234;
wire v_16235;
wire v_16236;
wire v_16237;
wire v_16238;
wire v_16239;
wire v_16240;
wire v_16241;
wire v_16242;
wire v_16243;
wire v_16244;
wire v_16245;
wire v_16246;
wire v_16247;
wire v_16248;
wire v_16249;
wire v_16250;
wire v_16251;
wire v_16252;
wire v_16253;
wire v_16254;
wire v_16255;
wire v_16256;
wire v_16257;
wire v_16258;
wire v_16259;
wire v_16260;
wire v_16261;
wire v_16262;
wire v_16263;
wire v_16264;
wire v_16265;
wire v_16266;
wire v_16267;
wire v_16268;
wire v_16269;
wire v_16270;
wire v_16271;
wire v_16272;
wire v_16273;
wire v_16274;
wire v_16275;
wire v_16276;
wire v_16277;
wire v_16278;
wire v_16279;
wire v_16280;
wire v_16281;
wire v_16282;
wire v_16283;
wire v_16284;
wire v_16285;
wire v_16286;
wire v_16287;
wire v_16288;
wire v_16289;
wire v_16290;
wire v_16291;
wire v_16292;
wire v_16293;
wire v_16294;
wire v_16295;
wire v_16296;
wire v_16297;
wire v_16298;
wire v_16299;
wire v_16300;
wire v_16301;
wire v_16302;
wire v_16303;
wire v_16304;
wire v_16305;
wire v_16306;
wire v_16307;
wire v_16308;
wire v_16309;
wire v_16310;
wire v_16311;
wire v_16312;
wire v_16313;
wire v_16314;
wire v_16315;
wire v_16316;
wire v_16317;
wire v_16318;
wire v_16319;
wire v_16320;
wire v_16321;
wire v_16322;
wire v_16323;
wire v_16324;
wire v_16325;
wire v_16326;
wire v_16327;
wire v_16328;
wire v_16329;
wire v_16330;
wire v_16331;
wire v_16332;
wire v_16333;
wire v_16334;
wire v_16335;
wire v_16336;
wire v_16337;
wire v_16338;
wire v_16339;
wire v_16340;
wire v_16341;
wire v_16342;
wire v_16343;
wire v_16344;
wire v_16345;
wire v_16346;
wire v_16347;
wire v_16348;
wire v_16349;
wire v_16350;
wire v_16351;
wire v_16352;
wire v_16353;
wire v_16354;
wire v_16355;
wire v_16356;
wire v_16357;
wire v_16358;
wire v_16359;
wire v_16360;
wire v_16361;
wire v_16362;
wire v_16363;
wire v_16364;
wire v_16365;
wire v_16366;
wire v_16367;
wire v_16368;
wire v_16369;
wire v_16370;
wire v_16371;
wire v_16372;
wire v_16373;
wire v_16374;
wire v_16375;
wire v_16376;
wire v_16377;
wire v_16378;
wire v_16379;
wire v_16380;
wire v_16381;
wire v_16382;
wire v_16383;
wire v_16384;
wire v_16385;
wire v_16386;
wire v_16387;
wire v_16388;
wire v_16389;
wire v_16390;
wire v_16391;
wire v_16392;
wire v_16393;
wire v_16394;
wire v_16395;
wire v_16396;
wire v_16397;
wire v_16398;
wire v_16399;
wire v_16400;
wire v_16401;
wire v_16402;
wire v_16403;
wire v_16404;
wire v_16405;
wire v_16406;
wire v_16407;
wire v_16408;
wire v_16409;
wire v_16410;
wire v_16411;
wire v_16412;
wire v_16413;
wire v_16414;
wire v_16415;
wire v_16416;
wire v_16417;
wire v_16418;
wire v_16419;
wire v_16420;
wire v_16421;
wire v_16422;
wire v_16423;
wire v_16424;
wire v_16425;
wire v_16426;
wire v_16427;
wire v_16428;
wire v_16429;
wire v_16430;
wire v_16431;
wire v_16432;
wire v_16433;
wire v_16434;
wire v_16435;
wire v_16436;
wire v_16437;
wire v_16438;
wire v_16439;
wire v_16440;
wire v_16441;
wire v_16442;
wire v_16443;
wire v_16444;
wire v_16445;
wire v_16446;
wire v_16447;
wire v_16448;
wire v_16449;
wire v_16450;
wire v_16451;
wire v_16452;
wire v_16453;
wire v_16454;
wire v_16455;
wire v_16456;
wire v_16457;
wire v_16458;
wire v_16459;
wire v_16460;
wire v_16461;
wire v_16462;
wire v_16463;
wire v_16464;
wire v_16465;
wire v_16466;
wire v_16467;
wire v_16468;
wire v_16469;
wire v_16470;
wire v_16471;
wire v_16472;
wire v_16473;
wire v_16474;
wire v_16475;
wire v_16476;
wire v_16477;
wire v_16478;
wire v_16479;
wire v_16480;
wire v_16481;
wire v_16482;
wire v_16483;
wire v_16484;
wire v_16485;
wire v_16486;
wire v_16487;
wire v_16488;
wire v_16489;
wire v_16490;
wire v_16491;
wire v_16492;
wire v_16493;
wire v_16494;
wire v_16495;
wire v_16496;
wire v_16497;
wire v_16498;
wire v_16499;
wire v_16500;
wire v_16501;
wire v_16502;
wire v_16503;
wire v_16504;
wire v_16505;
wire v_16506;
wire v_16507;
wire v_16508;
wire v_16509;
wire v_16510;
wire v_16511;
wire v_16512;
wire v_16513;
wire v_16514;
wire v_16515;
wire v_16516;
wire v_16517;
wire v_16518;
wire v_16519;
wire v_16520;
wire v_16521;
wire v_16522;
wire v_16523;
wire v_16524;
wire v_16525;
wire v_16526;
wire v_16527;
wire v_16528;
wire v_16529;
wire v_16530;
wire v_16531;
wire v_16532;
wire v_16533;
wire v_16534;
wire v_16535;
wire v_16536;
wire v_16537;
wire v_16538;
wire v_16539;
wire v_16540;
wire v_16541;
wire v_16542;
wire v_16543;
wire v_16544;
wire v_16545;
wire v_16546;
wire v_16547;
wire v_16548;
wire v_16549;
wire v_16550;
wire v_16551;
wire v_16552;
wire v_16553;
wire v_16554;
wire v_16555;
wire v_16556;
wire v_16557;
wire v_16558;
wire v_16559;
wire v_16560;
wire v_16561;
wire v_16562;
wire v_16563;
wire v_16564;
wire v_16565;
wire v_16566;
wire v_16567;
wire v_16568;
wire v_16569;
wire v_16570;
wire v_16571;
wire v_16572;
wire v_16573;
wire v_16574;
wire v_16575;
wire v_16576;
wire v_16577;
wire v_16578;
wire v_16579;
wire v_16580;
wire v_16581;
wire v_16582;
wire v_16583;
wire v_16584;
wire v_16585;
wire v_16586;
wire v_16587;
wire v_16588;
wire v_16589;
wire v_16590;
wire v_16591;
wire v_16592;
wire v_16593;
wire v_16594;
wire v_16595;
wire v_16596;
wire v_16597;
wire v_16598;
wire v_16599;
wire v_16600;
wire v_16601;
wire v_16602;
wire v_16603;
wire v_16604;
wire v_16605;
wire v_16606;
wire v_16607;
wire v_16608;
wire v_16609;
wire v_16610;
wire v_16611;
wire v_16612;
wire v_16613;
wire v_16614;
wire v_16615;
wire v_16616;
wire v_16617;
wire v_16618;
wire v_16619;
wire v_16620;
wire v_16621;
wire v_16622;
wire v_16623;
wire v_16624;
wire v_16625;
wire v_16626;
wire v_16627;
wire v_16628;
wire v_16629;
wire v_16630;
wire v_16631;
wire v_16632;
wire v_16633;
wire v_16634;
wire v_16635;
wire v_16636;
wire v_16637;
wire v_16638;
wire v_16639;
wire v_16640;
wire v_16641;
wire v_16642;
wire v_16643;
wire v_16644;
wire v_16645;
wire v_16646;
wire v_16647;
wire v_16648;
wire v_16649;
wire v_16650;
wire v_16651;
wire v_16652;
wire v_16653;
wire v_16654;
wire v_16655;
wire v_16656;
wire v_16657;
wire v_16658;
wire v_16659;
wire v_16660;
wire v_16661;
wire v_16662;
wire v_16663;
wire v_16664;
wire v_16665;
wire v_16666;
wire v_16667;
wire v_16668;
wire v_16669;
wire v_16670;
wire v_16671;
wire v_16672;
wire v_16673;
wire v_16674;
wire v_16675;
wire v_16676;
wire v_16677;
wire v_16678;
wire v_16679;
wire v_16680;
wire v_16681;
wire v_16682;
wire v_16683;
wire v_16684;
wire v_16685;
wire v_16686;
wire v_16687;
wire v_16688;
wire v_16689;
wire v_16690;
wire v_16691;
wire v_16692;
wire v_16693;
wire v_16694;
wire v_16695;
wire v_16696;
wire v_16697;
wire v_16698;
wire v_16699;
wire v_16700;
wire v_16701;
wire v_16702;
wire v_16703;
wire v_16704;
wire v_16705;
wire v_16706;
wire v_16707;
wire v_16708;
wire v_16709;
wire v_16710;
wire v_16711;
wire v_16712;
wire v_16713;
wire v_16714;
wire v_16715;
wire v_16716;
wire v_16717;
wire v_16718;
wire v_16719;
wire v_16720;
wire v_16721;
wire v_16722;
wire v_16723;
wire v_16724;
wire v_16725;
wire v_16726;
wire v_16727;
wire v_16728;
wire v_16729;
wire v_16730;
wire v_16731;
wire v_16732;
wire v_16733;
wire v_16734;
wire v_16735;
wire v_16736;
wire v_16737;
wire v_16738;
wire v_16739;
wire v_16740;
wire v_16741;
wire v_16742;
wire v_16743;
wire v_16744;
wire v_16745;
wire v_16746;
wire v_16747;
wire v_16748;
wire v_16749;
wire v_16750;
wire v_16751;
wire v_16752;
wire v_16753;
wire v_16754;
wire v_16755;
wire v_16756;
wire v_16757;
wire v_16758;
wire v_16759;
wire v_16760;
wire v_16761;
wire v_16762;
wire v_16763;
wire v_16764;
wire v_16765;
wire v_16766;
wire v_16767;
wire v_16768;
wire v_16769;
wire v_16770;
wire v_16771;
wire v_16772;
wire v_16773;
wire v_16774;
wire v_16775;
wire v_16776;
wire v_16777;
wire v_16778;
wire v_16779;
wire v_16780;
wire v_16781;
wire v_16782;
wire v_16783;
wire v_16784;
wire v_16785;
wire v_16786;
wire v_16787;
wire v_16788;
wire v_16789;
wire v_16790;
wire v_16791;
wire v_16792;
wire v_16793;
wire v_16794;
wire v_16795;
wire v_16796;
wire v_16797;
wire v_16798;
wire v_16799;
wire v_16800;
wire v_16801;
wire v_16802;
wire v_16803;
wire v_16804;
wire v_16805;
wire v_16806;
wire v_16807;
wire v_16808;
wire v_16809;
wire v_16810;
wire v_16811;
wire v_16812;
wire v_16813;
wire v_16814;
wire v_16815;
wire v_16816;
wire v_16817;
wire v_16818;
wire v_16819;
wire v_16820;
wire v_16821;
wire v_16822;
wire v_16823;
wire v_16824;
wire v_16825;
wire v_16826;
wire v_16827;
wire v_16828;
wire v_16829;
wire v_16830;
wire v_16831;
wire v_16832;
wire v_16833;
wire v_16834;
wire v_16835;
wire v_16836;
wire v_16837;
wire v_16838;
wire v_16839;
wire v_16840;
wire v_16841;
wire v_16842;
wire v_16843;
wire v_16844;
wire v_16845;
wire v_16846;
wire v_16847;
wire v_16848;
wire v_16849;
wire v_16850;
wire v_16851;
wire v_16852;
wire v_16853;
wire v_16854;
wire v_16855;
wire v_16856;
wire v_16857;
wire v_16858;
wire v_16859;
wire v_16860;
wire v_16861;
wire v_16862;
wire v_16863;
wire v_16864;
wire v_16865;
wire v_16866;
wire v_16867;
wire v_16868;
wire v_16869;
wire v_16870;
wire v_16871;
wire v_16872;
wire v_16873;
wire v_16874;
wire v_16875;
wire v_16876;
wire v_16877;
wire v_16878;
wire v_16879;
wire v_16880;
wire v_16881;
wire v_16882;
wire v_16883;
wire v_16884;
wire v_16885;
wire v_16886;
wire v_16887;
wire v_16888;
wire v_16889;
wire v_16890;
wire v_16891;
wire v_16892;
wire v_16893;
wire v_16894;
wire v_16895;
wire v_16896;
wire v_16897;
wire v_16898;
wire v_16899;
wire v_16900;
wire v_16901;
wire v_16902;
wire v_16903;
wire v_16904;
wire v_16905;
wire v_16906;
wire v_16907;
wire v_16908;
wire v_16909;
wire v_16910;
wire v_16911;
wire v_16912;
wire v_16913;
wire v_16914;
wire v_16915;
wire v_16916;
wire v_16917;
wire v_16918;
wire v_16919;
wire v_16920;
wire v_16921;
wire v_16922;
wire v_16923;
wire v_16924;
wire v_16925;
wire v_16926;
wire v_16927;
wire v_16928;
wire v_16929;
wire v_16930;
wire v_16931;
wire v_16932;
wire v_16933;
wire v_16934;
wire v_16935;
wire v_16936;
wire v_16937;
wire v_16938;
wire v_16939;
wire v_16940;
wire v_16941;
wire v_16942;
wire v_16943;
wire v_16944;
wire v_16945;
wire v_16946;
wire v_16947;
wire v_16948;
wire v_16949;
wire v_16950;
wire v_16951;
wire v_16952;
wire v_16953;
wire v_16954;
wire v_16955;
wire v_16956;
wire v_16957;
wire v_16958;
wire v_16959;
wire v_16960;
wire v_16961;
wire v_16962;
wire v_16963;
wire v_16964;
wire v_16965;
wire v_16966;
wire v_16967;
wire v_16968;
wire v_16969;
wire v_16970;
wire v_16971;
wire v_16972;
wire v_16973;
wire v_16974;
wire v_16975;
wire v_16976;
wire v_16977;
wire v_16978;
wire v_16979;
wire v_16980;
wire v_16981;
wire v_16982;
wire v_16983;
wire v_16984;
wire v_16985;
wire v_16986;
wire v_16987;
wire v_16988;
wire v_16989;
wire v_16990;
wire v_16991;
wire v_16992;
wire v_16993;
wire v_16994;
wire v_16995;
wire v_16996;
wire v_16997;
wire v_16998;
wire v_16999;
wire v_17000;
wire v_17001;
wire v_17002;
wire v_17003;
wire v_17004;
wire v_17005;
wire v_17006;
wire v_17007;
wire v_17008;
wire v_17009;
wire v_17010;
wire v_17011;
wire v_17012;
wire v_17013;
wire v_17014;
wire v_17015;
wire v_17016;
wire v_17017;
wire v_17018;
wire v_17019;
wire v_17020;
wire v_17021;
wire v_17022;
wire v_17023;
wire v_17024;
wire v_17025;
wire v_17026;
wire v_17027;
wire v_17028;
wire v_17029;
wire v_17030;
wire v_17031;
wire v_17032;
wire v_17033;
wire v_17034;
wire v_17035;
wire v_17036;
wire v_17037;
wire v_17038;
wire v_17039;
wire v_17040;
wire v_17041;
wire v_17042;
wire v_17043;
wire v_17044;
wire v_17045;
wire v_17046;
wire v_17047;
wire v_17048;
wire v_17049;
wire v_17050;
wire v_17051;
wire v_17052;
wire v_17053;
wire v_17054;
wire v_17055;
wire v_17056;
wire v_17057;
wire v_17058;
wire v_17059;
wire v_17060;
wire v_17061;
wire v_17062;
wire v_17063;
wire v_17064;
wire v_17065;
wire v_17066;
wire v_17067;
wire v_17068;
wire v_17069;
wire v_17070;
wire v_17071;
wire v_17072;
wire v_17073;
wire v_17074;
wire v_17075;
wire v_17076;
wire v_17077;
wire v_17078;
wire v_17079;
wire v_17080;
wire v_17081;
wire v_17082;
wire v_17083;
wire v_17084;
wire v_17085;
wire v_17086;
wire v_17087;
wire v_17088;
wire v_17089;
wire v_17090;
wire v_17091;
wire v_17092;
wire v_17093;
wire v_17094;
wire v_17095;
wire v_17096;
wire v_17097;
wire v_17098;
wire v_17099;
wire v_17100;
wire v_17101;
wire v_17102;
wire v_17103;
wire v_17104;
wire v_17105;
wire v_17106;
wire v_17107;
wire v_17108;
wire v_17109;
wire v_17110;
wire v_17111;
wire v_17112;
wire v_17113;
wire v_17114;
wire v_17115;
wire v_17116;
wire v_17117;
wire v_17118;
wire v_17119;
wire v_17120;
wire v_17121;
wire v_17122;
wire v_17123;
wire v_17124;
wire v_17125;
wire v_17126;
wire v_17127;
wire v_17128;
wire v_17129;
wire v_17130;
wire v_17131;
wire v_17132;
wire v_17133;
wire v_17134;
wire v_17135;
wire v_17136;
wire v_17137;
wire v_17138;
wire v_17139;
wire v_17140;
wire v_17141;
wire v_17142;
wire v_17143;
wire v_17144;
wire v_17145;
wire v_17146;
wire v_17147;
wire v_17148;
wire v_17149;
wire v_17150;
wire v_17151;
wire v_17152;
wire v_17153;
wire v_17154;
wire v_17155;
wire v_17156;
wire v_17157;
wire v_17158;
wire v_17159;
wire v_17160;
wire v_17161;
wire v_17162;
wire v_17163;
wire v_17164;
wire v_17165;
wire v_17166;
wire v_17167;
wire v_17168;
wire v_17169;
wire v_17170;
wire v_17171;
wire v_17172;
wire v_17173;
wire v_17174;
wire v_17175;
wire v_17176;
wire v_17177;
wire v_17178;
wire v_17179;
wire v_17180;
wire v_17181;
wire v_17182;
wire v_17183;
wire v_17184;
wire v_17185;
wire v_17186;
wire v_17187;
wire v_17188;
wire v_17189;
wire v_17190;
wire v_17191;
wire v_17192;
wire v_17193;
wire v_17194;
wire v_17195;
wire v_17196;
wire v_17197;
wire v_17198;
wire v_17199;
wire v_17200;
wire v_17201;
wire v_17202;
wire v_17203;
wire v_17204;
wire v_17205;
wire v_17206;
wire v_17207;
wire v_17208;
wire v_17209;
wire v_17210;
wire v_17211;
wire v_17212;
wire v_17213;
wire v_17214;
wire v_17215;
wire v_17216;
wire v_17217;
wire v_17218;
wire v_17219;
wire v_17220;
wire v_17221;
wire v_17222;
wire v_17223;
wire v_17224;
wire v_17225;
wire v_17226;
wire v_17227;
wire v_17228;
wire v_17229;
wire v_17230;
wire v_17231;
wire v_17232;
wire v_17233;
wire v_17234;
wire v_17235;
wire v_17236;
wire v_17237;
wire v_17238;
wire v_17239;
wire v_17240;
wire v_17241;
wire v_17242;
wire v_17243;
wire v_17244;
wire v_17245;
wire v_17246;
wire v_17247;
wire v_17248;
wire v_17249;
wire v_17250;
wire v_17251;
wire v_17252;
wire v_17253;
wire v_17254;
wire v_17255;
wire v_17256;
wire v_17257;
wire v_17258;
wire v_17259;
wire v_17260;
wire v_17261;
wire v_17262;
wire v_17263;
wire v_17264;
wire v_17265;
wire v_17266;
wire v_17267;
wire v_17268;
wire v_17269;
wire v_17270;
wire v_17271;
wire v_17272;
wire v_17273;
wire v_17274;
wire v_17275;
wire v_17276;
wire v_17277;
wire v_17278;
wire v_17279;
wire v_17280;
wire v_17281;
wire v_17282;
wire v_17283;
wire v_17284;
wire v_17285;
wire v_17286;
wire v_17287;
wire v_17288;
wire v_17289;
wire v_17290;
wire v_17291;
wire v_17292;
wire v_17293;
wire v_17294;
wire v_17295;
wire v_17296;
wire v_17297;
wire v_17298;
wire v_17299;
wire v_17300;
wire v_17301;
wire v_17302;
wire v_17303;
wire v_17304;
wire v_17305;
wire v_17306;
wire v_17307;
wire v_17308;
wire v_17309;
wire v_17310;
wire v_17311;
wire v_17312;
wire v_17313;
wire v_17314;
wire v_17315;
wire v_17316;
wire v_17317;
wire v_17318;
wire v_17319;
wire v_17320;
wire v_17321;
wire v_17322;
wire v_17323;
wire v_17324;
wire v_17325;
wire v_17326;
wire v_17327;
wire v_17328;
wire v_17329;
wire v_17330;
wire v_17331;
wire v_17332;
wire v_17333;
wire v_17334;
wire v_17335;
wire v_17336;
wire v_17337;
wire v_17338;
wire v_17339;
wire v_17340;
wire v_17341;
wire v_17342;
wire v_17343;
wire v_17344;
wire v_17345;
wire v_17346;
wire v_17347;
wire v_17348;
wire v_17349;
wire v_17350;
wire v_17351;
wire v_17352;
wire v_17353;
wire v_17354;
wire v_17355;
wire v_17356;
wire v_17357;
wire v_17358;
wire v_17359;
wire v_17360;
wire v_17361;
wire v_17362;
wire v_17363;
wire v_17364;
wire v_17365;
wire v_17366;
wire v_17367;
wire v_17368;
wire v_17369;
wire v_17370;
wire v_17371;
wire v_17372;
wire v_17373;
wire v_17374;
wire v_17375;
wire v_17376;
wire v_17377;
wire v_17378;
wire v_17379;
wire v_17380;
wire v_17381;
wire v_17382;
wire v_17383;
wire v_17384;
wire v_17385;
wire v_17386;
wire v_17387;
wire v_17388;
wire v_17389;
wire v_17390;
wire v_17391;
wire v_17392;
wire v_17393;
wire v_17394;
wire v_17395;
wire v_17396;
wire v_17397;
wire v_17398;
wire v_17399;
wire v_17400;
wire v_17401;
wire v_17402;
wire v_17403;
wire v_17404;
wire v_17405;
wire v_17406;
wire v_17407;
wire v_17408;
wire v_17409;
wire v_17410;
wire v_17411;
wire v_17412;
wire v_17413;
wire v_17414;
wire v_17415;
wire v_17416;
wire v_17417;
wire v_17418;
wire v_17419;
wire v_17420;
wire v_17421;
wire v_17422;
wire v_17423;
wire v_17424;
wire v_17425;
wire v_17426;
wire v_17427;
wire v_17428;
wire v_17429;
wire v_17430;
wire v_17431;
wire v_17432;
wire v_17433;
wire v_17434;
wire v_17435;
wire v_17436;
wire v_17437;
wire v_17438;
wire v_17439;
wire v_17440;
wire v_17441;
wire v_17442;
wire v_17443;
wire v_17444;
wire v_17445;
wire v_17446;
wire v_17447;
wire v_17448;
wire v_17449;
wire v_17450;
wire v_17451;
wire v_17452;
wire v_17453;
wire v_17454;
wire v_17455;
wire v_17456;
wire v_17457;
wire v_17458;
wire v_17459;
wire v_17460;
wire v_17461;
wire v_17462;
wire v_17463;
wire v_17464;
wire v_17465;
wire v_17466;
wire v_17467;
wire v_17468;
wire v_17469;
wire v_17470;
wire v_17471;
wire v_17472;
wire v_17473;
wire v_17474;
wire v_17475;
wire v_17476;
wire v_17477;
wire v_17478;
wire v_17479;
wire v_17480;
wire v_17481;
wire v_17482;
wire v_17483;
wire v_17484;
wire v_17485;
wire v_17486;
wire v_17487;
wire v_17488;
wire v_17489;
wire v_17490;
wire v_17491;
wire v_17492;
wire v_17493;
wire v_17494;
wire v_17495;
wire v_17496;
wire v_17497;
wire v_17498;
wire v_17499;
wire v_17500;
wire v_17501;
wire v_17502;
wire v_17503;
wire v_17504;
wire v_17505;
wire v_17506;
wire v_17507;
wire v_17508;
wire v_17509;
wire v_17510;
wire v_17511;
wire v_17512;
wire v_17513;
wire v_17514;
wire v_17515;
wire v_17516;
wire v_17517;
wire v_17518;
wire v_17519;
wire v_17520;
wire v_17521;
wire v_17522;
wire v_17523;
wire v_17524;
wire v_17525;
wire v_17526;
wire v_17527;
wire v_17528;
wire v_17529;
wire v_17530;
wire v_17531;
wire v_17532;
wire v_17533;
wire v_17534;
wire v_17535;
wire v_17536;
wire v_17537;
wire v_17538;
wire v_17539;
wire v_17540;
wire v_17541;
wire v_17542;
wire v_17543;
wire v_17544;
wire v_17545;
wire v_17546;
wire v_17547;
wire v_17548;
wire v_17549;
wire v_17550;
wire v_17551;
wire v_17552;
wire v_17553;
wire v_17554;
wire v_17555;
wire v_17556;
wire v_17557;
wire v_17558;
wire v_17559;
wire v_17560;
wire v_17561;
wire v_17562;
wire v_17563;
wire v_17564;
wire v_17565;
wire v_17566;
wire v_17567;
wire v_17568;
wire v_17569;
wire v_17570;
wire v_17571;
wire v_17572;
wire v_17573;
wire v_17574;
wire v_17575;
wire v_17576;
wire v_17577;
wire v_17578;
wire v_17579;
wire v_17580;
wire v_17581;
wire v_17582;
wire v_17583;
wire v_17584;
wire v_17585;
wire v_17586;
wire v_17587;
wire v_17588;
wire v_17589;
wire v_17590;
wire v_17591;
wire v_17592;
wire v_17593;
wire v_17594;
wire v_17595;
wire v_17596;
wire v_17597;
wire v_17598;
wire v_17599;
wire v_17600;
wire v_17601;
wire v_17602;
wire v_17603;
wire v_17604;
wire v_17605;
wire v_17606;
wire v_17607;
wire v_17608;
wire v_17609;
wire v_17610;
wire v_17611;
wire v_17612;
wire v_17613;
wire v_17614;
wire v_17615;
wire v_17616;
wire v_17617;
wire v_17618;
wire v_17619;
wire v_17620;
wire v_17621;
wire v_17622;
wire v_17623;
wire v_17624;
wire v_17625;
wire v_17626;
wire v_17627;
wire v_17628;
wire v_17629;
wire v_17630;
wire v_17631;
wire v_17632;
wire v_17633;
wire v_17634;
wire v_17635;
wire v_17636;
wire v_17637;
wire v_17638;
wire v_17639;
wire v_17640;
wire v_17641;
wire v_17642;
wire v_17643;
wire v_17644;
wire v_17645;
wire v_17646;
wire v_17647;
wire v_17648;
wire v_17649;
wire v_17650;
wire v_17651;
wire v_17652;
wire v_17653;
wire v_17654;
wire v_17655;
wire v_17656;
wire v_17657;
wire v_17658;
wire v_17659;
wire v_17660;
wire v_17661;
wire v_17662;
wire v_17663;
wire v_17664;
wire v_17665;
wire v_17666;
wire v_17667;
wire v_17668;
wire v_17669;
wire v_17670;
wire v_17671;
wire v_17672;
wire v_17673;
wire v_17674;
wire v_17675;
wire v_17676;
wire v_17677;
wire v_17678;
wire v_17679;
wire v_17680;
wire v_17681;
wire v_17682;
wire v_17683;
wire v_17684;
wire v_17685;
wire v_17686;
wire v_17687;
wire v_17688;
wire v_17689;
wire v_17690;
wire v_17691;
wire v_17692;
wire v_17693;
wire v_17694;
wire v_17695;
wire v_17696;
wire v_17697;
wire v_17698;
wire v_17699;
wire v_17700;
wire v_17701;
wire v_17702;
wire v_17703;
wire v_17704;
wire v_17705;
wire v_17706;
wire v_17707;
wire v_17708;
wire v_17709;
wire v_17710;
wire v_17711;
wire v_17712;
wire v_17713;
wire v_17714;
wire v_17715;
wire v_17716;
wire v_17717;
wire v_17718;
wire v_17719;
wire v_17720;
wire v_17721;
wire v_17722;
wire v_17723;
wire v_17724;
wire v_17725;
wire v_17726;
wire v_17727;
wire v_17728;
wire v_17729;
wire v_17730;
wire v_17731;
wire v_17732;
wire v_17733;
wire v_17734;
wire v_17735;
wire v_17736;
wire v_17737;
wire v_17738;
wire v_17739;
wire v_17740;
wire v_17741;
wire v_17742;
wire v_17743;
wire v_17744;
wire v_17745;
wire v_17746;
wire v_17747;
wire v_17748;
wire v_17749;
wire v_17750;
wire v_17751;
wire v_17752;
wire v_17753;
wire v_17754;
wire v_17755;
wire v_17756;
wire v_17757;
wire v_17758;
wire v_17759;
wire v_17760;
wire v_17761;
wire v_17762;
wire v_17763;
wire v_17764;
wire v_17765;
wire v_17766;
wire v_17767;
wire v_17768;
wire v_17769;
wire v_17770;
wire v_17771;
wire v_17772;
wire v_17773;
wire v_17774;
wire v_17775;
wire v_17776;
wire v_17777;
wire v_17778;
wire v_17779;
wire v_17780;
wire v_17781;
wire v_17782;
wire v_17783;
wire v_17784;
wire v_17785;
wire v_17786;
wire v_17787;
wire v_17788;
wire v_17789;
wire v_17790;
wire v_17791;
wire v_17792;
wire v_17793;
wire v_17794;
wire v_17795;
wire v_17796;
wire v_17797;
wire v_17798;
wire v_17799;
wire v_17800;
wire v_17801;
wire v_17802;
wire v_17803;
wire v_17804;
wire v_17805;
wire v_17806;
wire v_17807;
wire v_17808;
wire v_17809;
wire v_17810;
wire v_17811;
wire v_17812;
wire v_17813;
wire v_17814;
wire v_17815;
wire v_17816;
wire v_17817;
wire v_17818;
wire v_17819;
wire v_17820;
wire v_17821;
wire v_17822;
wire v_17823;
wire v_17824;
wire v_17825;
wire v_17826;
wire v_17827;
wire v_17828;
wire v_17829;
wire v_17830;
wire v_17831;
wire v_17832;
wire v_17833;
wire v_17834;
wire v_17835;
wire v_17836;
wire v_17837;
wire v_17838;
wire v_17839;
wire v_17840;
wire v_17841;
wire v_17842;
wire v_17843;
wire v_17844;
wire v_17845;
wire v_17846;
wire v_17847;
wire v_17848;
wire v_17849;
wire v_17850;
wire v_17851;
wire v_17852;
wire v_17853;
wire v_17854;
wire v_17855;
wire v_17856;
wire v_17857;
wire v_17858;
wire v_17859;
wire v_17860;
wire v_17861;
wire v_17862;
wire v_17863;
wire v_17864;
wire v_17865;
wire v_17866;
wire v_17867;
wire v_17868;
wire v_17869;
wire v_17870;
wire v_17871;
wire v_17872;
wire v_17873;
wire v_17874;
wire v_17875;
wire v_17876;
wire v_17877;
wire v_17878;
wire v_17879;
wire v_17880;
wire v_17881;
wire v_17882;
wire v_17883;
wire v_17884;
wire v_17885;
wire v_17886;
wire v_17887;
wire v_17888;
wire v_17889;
wire v_17890;
wire v_17891;
wire v_17892;
wire v_17893;
wire v_17894;
wire v_17895;
wire v_17896;
wire v_17897;
wire v_17898;
wire v_17899;
wire v_17900;
wire v_17901;
wire v_17902;
wire v_17903;
wire v_17904;
wire v_17905;
wire v_17906;
wire v_17907;
wire v_17908;
wire v_17909;
wire v_17910;
wire v_17911;
wire v_17912;
wire v_17913;
wire v_17914;
wire v_17915;
wire v_17916;
wire v_17917;
wire v_17918;
wire v_17919;
wire v_17920;
wire v_17921;
wire v_17922;
wire v_17923;
wire v_17924;
wire v_17925;
wire v_17926;
wire v_17927;
wire v_17928;
wire v_17929;
wire v_17930;
wire v_17931;
wire v_17932;
wire v_17933;
wire v_17934;
wire v_17935;
wire v_17936;
wire v_17937;
wire v_17938;
wire v_17939;
wire v_17940;
wire v_17941;
wire v_17942;
wire v_17943;
wire v_17944;
wire v_17945;
wire v_17946;
wire v_17947;
wire v_17948;
wire v_17949;
wire v_17950;
wire v_17951;
wire v_17952;
wire v_17953;
wire v_17954;
wire v_17955;
wire v_17956;
wire v_17957;
wire v_17958;
wire v_17959;
wire v_17960;
wire v_17961;
wire v_17962;
wire v_17963;
wire v_17964;
wire v_17965;
wire v_17966;
wire v_17967;
wire v_17968;
wire v_17969;
wire v_17970;
wire v_17971;
wire v_17972;
wire v_17973;
wire v_17974;
wire v_17975;
wire v_17976;
wire v_17977;
wire v_17978;
wire v_17979;
wire v_17980;
wire v_17981;
wire v_17982;
wire v_17983;
wire v_17984;
wire v_17985;
wire v_17986;
wire v_17987;
wire v_17988;
wire v_17989;
wire v_17990;
wire v_17991;
wire v_17992;
wire v_17993;
wire v_17994;
wire v_17995;
wire v_17996;
wire v_17997;
wire v_17998;
wire v_17999;
wire v_18000;
wire v_18001;
wire v_18002;
wire v_18003;
wire v_18004;
wire v_18005;
wire v_18006;
wire v_18007;
wire v_18008;
wire v_18009;
wire v_18010;
wire v_18011;
wire v_18012;
wire v_18013;
wire v_18014;
wire v_18015;
wire v_18016;
wire v_18017;
wire v_18018;
wire v_18019;
wire v_18020;
wire v_18021;
wire v_18022;
wire v_18023;
wire v_18024;
wire v_18025;
wire v_18026;
wire v_18027;
wire v_18028;
wire v_18029;
wire v_18030;
wire v_18031;
wire v_18032;
wire v_18033;
wire v_18034;
wire v_18035;
wire v_18036;
wire v_18037;
wire v_18038;
wire v_18039;
wire v_18040;
wire v_18041;
wire v_18042;
wire v_18043;
wire v_18044;
wire v_18045;
wire v_18046;
wire v_18047;
wire v_18048;
wire v_18049;
wire v_18050;
wire v_18051;
wire v_18052;
wire v_18053;
wire v_18054;
wire v_18055;
wire v_18056;
wire v_18057;
wire v_18058;
wire v_18059;
wire v_18060;
wire v_18061;
wire v_18062;
wire v_18063;
wire v_18064;
wire v_18065;
wire v_18066;
wire v_18067;
wire v_18068;
wire v_18069;
wire v_18070;
wire v_18071;
wire v_18072;
wire v_18073;
wire v_18074;
wire v_18075;
wire v_18076;
wire v_18077;
wire v_18078;
wire v_18079;
wire v_18080;
wire v_18081;
wire v_18082;
wire v_18083;
wire v_18084;
wire v_18085;
wire v_18086;
wire v_18087;
wire v_18088;
wire v_18089;
wire v_18090;
wire v_18091;
wire v_18092;
wire v_18093;
wire v_18094;
wire v_18095;
wire v_18096;
wire v_18097;
wire v_18098;
wire v_18099;
wire v_18100;
wire v_18101;
wire v_18102;
wire v_18103;
wire v_18104;
wire v_18105;
wire v_18106;
wire v_18107;
wire v_18108;
wire v_18109;
wire v_18110;
wire v_18111;
wire v_18112;
wire v_18113;
wire v_18114;
wire v_18115;
wire v_18116;
wire v_18117;
wire v_18118;
wire v_18119;
wire v_18120;
wire v_18121;
wire v_18122;
wire v_18123;
wire v_18124;
wire v_18125;
wire v_18126;
wire v_18127;
wire v_18128;
wire v_18129;
wire v_18130;
wire v_18131;
wire v_18132;
wire v_18133;
wire v_18134;
wire v_18135;
wire v_18136;
wire v_18137;
wire v_18138;
wire v_18139;
wire v_18140;
wire v_18141;
wire v_18142;
wire v_18143;
wire v_18144;
wire v_18145;
wire v_18146;
wire v_18147;
wire v_18148;
wire v_18149;
wire v_18150;
wire v_18151;
wire v_18152;
wire v_18153;
wire v_18154;
wire v_18155;
wire v_18156;
wire v_18157;
wire v_18158;
wire v_18159;
wire v_18160;
wire v_18161;
wire v_18162;
wire v_18163;
wire v_18164;
wire v_18165;
wire v_18166;
wire v_18167;
wire v_18168;
wire v_18169;
wire v_18170;
wire v_18171;
wire v_18172;
wire v_18173;
wire v_18174;
wire v_18175;
wire v_18176;
wire v_18177;
wire v_18178;
wire v_18179;
wire v_18180;
wire v_18181;
wire v_18182;
wire v_18183;
wire v_18184;
wire v_18185;
wire v_18186;
wire v_18187;
wire v_18188;
wire v_18189;
wire v_18190;
wire v_18191;
wire v_18192;
wire v_18193;
wire v_18194;
wire v_18195;
wire v_18196;
wire v_18197;
wire v_18198;
wire v_18199;
wire v_18200;
wire v_18201;
wire v_18202;
wire v_18203;
wire v_18204;
wire v_18205;
wire v_18206;
wire v_18207;
wire v_18208;
wire v_18209;
wire v_18210;
wire v_18211;
wire v_18212;
wire v_18213;
wire v_18214;
wire v_18215;
wire v_18216;
wire v_18217;
wire v_18218;
wire v_18219;
wire v_18220;
wire v_18221;
wire v_18222;
wire v_18223;
wire v_18224;
wire v_18225;
wire v_18226;
wire v_18227;
wire v_18228;
wire v_18229;
wire v_18230;
wire v_18231;
wire v_18232;
wire v_18233;
wire v_18234;
wire v_18235;
wire v_18236;
wire v_18237;
wire v_18238;
wire v_18239;
wire v_18240;
wire v_18241;
wire v_18242;
wire v_18243;
wire v_18244;
wire v_18245;
wire v_18246;
wire v_18247;
wire v_18248;
wire v_18249;
wire v_18250;
wire v_18251;
wire v_18252;
wire v_18253;
wire v_18254;
wire v_18255;
wire v_18256;
wire v_18257;
wire v_18258;
wire v_18259;
wire v_18260;
wire v_18261;
wire v_18262;
wire v_18263;
wire v_18264;
wire v_18265;
wire v_18266;
wire v_18267;
wire v_18268;
wire v_18269;
wire v_18270;
wire v_18271;
wire v_18272;
wire v_18273;
wire v_18274;
wire v_18275;
wire v_18276;
wire v_18277;
wire v_18278;
wire v_18279;
wire v_18280;
wire v_18281;
wire v_18282;
wire v_18283;
wire v_18284;
wire v_18285;
wire v_18286;
wire v_18287;
wire v_18288;
wire v_18289;
wire v_18290;
wire v_18291;
wire v_18292;
wire v_18293;
wire v_18294;
wire v_18295;
wire v_18296;
wire v_18297;
wire v_18298;
wire v_18299;
wire v_18300;
wire v_18301;
wire v_18302;
wire v_18303;
wire v_18304;
wire v_18305;
wire v_18306;
wire v_18307;
wire v_18308;
wire v_18309;
wire v_18310;
wire v_18311;
wire v_18312;
wire v_18313;
wire v_18314;
wire v_18315;
wire v_18316;
wire v_18317;
wire v_18318;
wire v_18319;
wire v_18320;
wire v_18321;
wire v_18322;
wire v_18323;
wire v_18324;
wire v_18325;
wire v_18326;
wire v_18327;
wire v_18328;
wire v_18329;
wire v_18330;
wire v_18331;
wire v_18332;
wire v_18333;
wire v_18334;
wire v_18335;
wire v_18336;
wire v_18337;
wire v_18338;
wire v_18339;
wire v_18340;
wire v_18341;
wire v_18342;
wire v_18343;
wire v_18344;
wire v_18345;
wire v_18346;
wire v_18347;
wire v_18348;
wire v_18349;
wire v_18350;
wire v_18351;
wire v_18352;
wire v_18353;
wire v_18354;
wire v_18355;
wire v_18356;
wire v_18357;
wire v_18358;
wire v_18359;
wire v_18360;
wire v_18361;
wire v_18362;
wire v_18363;
wire v_18364;
wire v_18365;
wire v_18366;
wire v_18367;
wire v_18368;
wire v_18369;
wire v_18370;
wire v_18371;
wire v_18372;
wire v_18373;
wire v_18374;
wire v_18375;
wire v_18376;
wire v_18377;
wire v_18378;
wire v_18379;
wire v_18380;
wire v_18381;
wire v_18382;
wire v_18383;
wire v_18384;
wire v_18385;
wire v_18386;
wire v_18387;
wire v_18388;
wire v_18389;
wire v_18390;
wire v_18391;
wire v_18392;
wire v_18393;
wire v_18394;
wire v_18395;
wire v_18396;
wire v_18397;
wire v_18398;
wire v_18399;
wire v_18400;
wire v_18401;
wire v_18402;
wire v_18403;
wire v_18404;
wire v_18405;
wire v_18406;
wire v_18407;
wire v_18408;
wire v_18409;
wire v_18410;
wire v_18411;
wire v_18412;
wire v_18413;
wire v_18414;
wire v_18415;
wire v_18416;
wire v_18417;
wire v_18418;
wire v_18419;
wire v_18420;
wire v_18421;
wire v_18422;
wire v_18423;
wire v_18424;
wire v_18425;
wire v_18426;
wire v_18427;
wire v_18428;
wire v_18429;
wire v_18430;
wire v_18431;
wire v_18432;
wire v_18433;
wire v_18434;
wire v_18435;
wire v_18436;
wire v_18437;
wire v_18438;
wire v_18439;
wire v_18440;
wire v_18441;
wire v_18442;
wire v_18443;
wire v_18444;
wire v_18445;
wire v_18446;
wire v_18447;
wire v_18448;
wire v_18449;
wire v_18450;
wire v_18451;
wire v_18452;
wire v_18453;
wire v_18454;
wire v_18455;
wire v_18456;
wire v_18457;
wire v_18458;
wire v_18459;
wire v_18460;
wire v_18461;
wire v_18462;
wire v_18463;
wire v_18464;
wire v_18465;
wire v_18466;
wire v_18467;
wire v_18468;
wire v_18469;
wire v_18470;
wire v_18471;
wire v_18472;
wire v_18473;
wire v_18474;
wire v_18475;
wire v_18476;
wire v_18477;
wire v_18478;
wire v_18479;
wire v_18480;
wire v_18481;
wire v_18482;
wire v_18483;
wire v_18484;
wire v_18485;
wire v_18486;
wire v_18487;
wire v_18488;
wire v_18489;
wire v_18490;
wire v_18491;
wire v_18492;
wire v_18493;
wire v_18494;
wire v_18495;
wire v_18496;
wire v_18497;
wire v_18498;
wire v_18499;
wire v_18500;
wire v_18501;
wire v_18502;
wire v_18503;
wire v_18504;
wire v_18505;
wire v_18506;
wire v_18507;
wire v_18508;
wire v_18509;
wire v_18510;
wire v_18511;
wire v_18512;
wire v_18513;
wire v_18514;
wire v_18515;
wire v_18516;
wire v_18517;
wire v_18518;
wire v_18519;
wire v_18520;
wire v_18521;
wire v_18522;
wire v_18523;
wire v_18524;
wire v_18525;
wire v_18526;
wire v_18527;
wire v_18528;
wire v_18529;
wire v_18530;
wire v_18531;
wire v_18532;
wire v_18533;
wire v_18534;
wire v_18535;
wire v_18536;
wire v_18537;
wire v_18538;
wire v_18539;
wire v_18540;
wire v_18541;
wire v_18542;
wire v_18543;
wire v_18544;
wire v_18545;
wire v_18546;
wire v_18547;
wire v_18548;
wire v_18549;
wire v_18550;
wire v_18551;
wire v_18552;
wire v_18553;
wire v_18554;
wire v_18555;
wire v_18556;
wire v_18557;
wire v_18558;
wire v_18559;
wire v_18560;
wire v_18561;
wire v_18562;
wire v_18563;
wire v_18564;
wire v_18565;
wire v_18566;
wire v_18567;
wire v_18568;
wire v_18569;
wire v_18570;
wire v_18571;
wire v_18572;
wire v_18573;
wire v_18574;
wire v_18575;
wire v_18576;
wire v_18577;
wire v_18578;
wire v_18579;
wire v_18580;
wire v_18581;
wire v_18582;
wire v_18583;
wire v_18584;
wire v_18585;
wire v_18586;
wire v_18587;
wire v_18588;
wire v_18589;
wire v_18590;
wire v_18591;
wire v_18592;
wire v_18593;
wire v_18594;
wire v_18595;
wire v_18596;
wire v_18597;
wire v_18598;
wire v_18599;
wire v_18600;
wire v_18601;
wire v_18602;
wire v_18603;
wire v_18604;
wire v_18605;
wire v_18606;
wire v_18607;
wire v_18608;
wire v_18609;
wire v_18610;
wire v_18611;
wire v_18612;
wire v_18613;
wire v_18614;
wire v_18615;
wire v_18616;
wire v_18617;
wire v_18618;
wire v_18619;
wire v_18620;
wire v_18621;
wire v_18622;
wire v_18623;
wire v_18624;
wire v_18625;
wire v_18626;
wire v_18627;
wire v_18628;
wire v_18629;
wire v_18630;
wire v_18631;
wire v_18632;
wire v_18633;
wire v_18634;
wire v_18635;
wire v_18636;
wire v_18637;
wire v_18638;
wire v_18639;
wire v_18640;
wire v_18641;
wire v_18642;
wire v_18643;
wire v_18644;
wire v_18645;
wire v_18646;
wire v_18647;
wire v_18648;
wire v_18649;
wire v_18650;
wire v_18651;
wire v_18652;
wire v_18653;
wire v_18654;
wire v_18655;
wire v_18656;
wire v_18657;
wire v_18658;
wire v_18659;
wire v_18660;
wire v_18661;
wire v_18662;
wire v_18663;
wire v_18664;
wire v_18665;
wire v_18666;
wire v_18667;
wire v_18668;
wire v_18669;
wire v_18670;
wire v_18671;
wire v_18672;
wire v_18673;
wire v_18674;
wire v_18675;
wire v_18676;
wire v_18677;
wire v_18678;
wire v_18679;
wire v_18680;
wire v_18681;
wire v_18682;
wire v_18683;
wire v_18684;
wire v_18685;
wire v_18686;
wire v_18687;
wire v_18688;
wire v_18689;
wire v_18690;
wire v_18691;
wire v_18692;
wire v_18693;
wire v_18694;
wire v_18695;
wire v_18696;
wire v_18697;
wire v_18698;
wire v_18699;
wire v_18700;
wire v_18701;
wire v_18702;
wire v_18703;
wire v_18704;
wire v_18705;
wire v_18706;
wire v_18707;
wire v_18708;
wire v_18709;
wire v_18710;
wire v_18711;
wire v_18712;
wire v_18713;
wire v_18714;
wire v_18715;
wire v_18716;
wire v_18717;
wire v_18718;
wire v_18719;
wire v_18720;
wire v_18721;
wire v_18722;
wire v_18723;
wire v_18724;
wire v_18725;
wire v_18726;
wire v_18727;
wire v_18728;
wire v_18729;
wire v_18730;
wire v_18731;
wire v_18732;
wire v_18733;
wire v_18734;
wire v_18735;
wire v_18736;
wire v_18737;
wire v_18738;
wire v_18739;
wire v_18740;
wire v_18741;
wire v_18742;
wire v_18743;
wire v_18744;
wire v_18745;
wire v_18746;
wire v_18747;
wire v_18748;
wire v_18749;
wire v_18750;
wire v_18751;
wire v_18752;
wire v_18753;
wire v_18754;
wire v_18755;
wire v_18756;
wire v_18757;
wire v_18758;
wire v_18759;
wire v_18760;
wire v_18761;
wire v_18762;
wire v_18763;
wire v_18764;
wire v_18765;
wire v_18766;
wire v_18767;
wire v_18768;
wire v_18769;
wire v_18770;
wire v_18771;
wire v_18772;
wire v_18773;
wire v_18774;
wire v_18775;
wire v_18776;
wire v_18777;
wire v_18778;
wire v_18779;
wire v_18780;
wire v_18781;
wire v_18782;
wire v_18783;
wire v_18784;
wire v_18785;
wire v_18786;
wire v_18787;
wire v_18788;
wire v_18789;
wire v_18790;
wire v_18791;
wire v_18792;
wire v_18793;
wire v_18794;
wire v_18795;
wire v_18796;
wire v_18797;
wire v_18798;
wire v_18799;
wire v_18800;
wire v_18801;
wire v_18802;
wire v_18803;
wire v_18804;
wire v_18805;
wire v_18806;
wire v_18807;
wire v_18808;
wire v_18809;
wire v_18810;
wire v_18811;
wire v_18812;
wire v_18813;
wire v_18814;
wire v_18815;
wire v_18816;
wire v_18817;
wire v_18818;
wire v_18819;
wire v_18820;
wire v_18821;
wire v_18822;
wire v_18823;
wire v_18824;
wire v_18825;
wire v_18826;
wire v_18827;
wire v_18828;
wire v_18829;
wire v_18830;
wire v_18831;
wire v_18832;
wire v_18833;
wire v_18834;
wire v_18835;
wire v_18836;
wire v_18837;
wire v_18838;
wire v_18839;
wire v_18840;
wire v_18841;
wire v_18842;
wire v_18843;
wire v_18844;
wire v_18845;
wire v_18846;
wire v_18847;
wire v_18848;
wire v_18849;
wire v_18850;
wire v_18851;
wire v_18852;
wire v_18853;
wire v_18854;
wire v_18855;
wire v_18856;
wire v_18857;
wire v_18858;
wire v_18859;
wire v_18860;
wire v_18861;
wire v_18862;
wire v_18863;
wire v_18864;
wire v_18865;
wire v_18866;
wire v_18867;
wire v_18868;
wire v_18869;
wire v_18870;
wire v_18871;
wire v_18872;
wire v_18873;
wire v_18874;
wire v_18875;
wire v_18876;
wire v_18877;
wire v_18878;
wire v_18879;
wire v_18880;
wire v_18881;
wire v_18882;
wire v_18883;
wire v_18884;
wire v_18885;
wire v_18886;
wire v_18887;
wire v_18888;
wire v_18889;
wire v_18890;
wire v_18891;
wire v_18892;
wire v_18893;
wire v_18894;
wire v_18895;
wire v_18896;
wire v_18897;
wire v_18898;
wire v_18899;
wire v_18900;
wire v_18901;
wire v_18902;
wire v_18903;
wire v_18904;
wire v_18905;
wire v_18906;
wire v_18907;
wire v_18908;
wire v_18909;
wire v_18910;
wire v_18911;
wire v_18912;
wire v_18913;
wire v_18914;
wire v_18915;
wire v_18916;
wire v_18917;
wire v_18918;
wire v_18919;
wire v_18920;
wire v_18921;
wire v_18922;
wire v_18923;
wire v_18924;
wire v_18925;
wire v_18926;
wire v_18927;
wire v_18928;
wire v_18929;
wire v_18930;
wire v_18931;
wire v_18932;
wire v_18933;
wire v_18934;
wire v_18935;
wire v_18936;
wire v_18937;
wire v_18938;
wire v_18939;
wire v_18940;
wire v_18941;
wire v_18942;
wire v_18943;
wire v_18944;
wire v_18945;
wire v_18946;
wire v_18947;
wire v_18948;
wire v_18949;
wire v_18950;
wire v_18951;
wire v_18952;
wire v_18953;
wire v_18954;
wire v_18955;
wire v_18956;
wire v_18957;
wire v_18958;
wire v_18959;
wire v_18960;
wire v_18961;
wire v_18962;
wire v_18963;
wire v_18964;
wire v_18965;
wire v_18966;
wire v_18967;
wire v_18968;
wire v_18969;
wire v_18970;
wire v_18971;
wire v_18972;
wire v_18973;
wire v_18974;
wire v_18975;
wire v_18976;
wire v_18977;
wire v_18978;
wire v_18979;
wire v_18980;
wire v_18981;
wire v_18982;
wire v_18983;
wire v_18984;
wire v_18985;
wire v_18986;
wire v_18987;
wire v_18988;
wire v_18989;
wire v_18990;
wire v_18991;
wire v_18992;
wire v_18993;
wire v_18994;
wire v_18995;
wire v_18996;
wire v_18997;
wire v_18998;
wire v_18999;
wire v_19000;
wire v_19001;
wire v_19002;
wire v_19003;
wire v_19004;
wire v_19005;
wire v_19006;
wire v_19007;
wire v_19008;
wire v_19009;
wire v_19010;
wire v_19011;
wire v_19012;
wire v_19013;
wire v_19014;
wire v_19015;
wire v_19016;
wire v_19017;
wire v_19018;
wire v_19019;
wire v_19020;
wire v_19021;
wire v_19022;
wire v_19023;
wire v_19024;
wire v_19025;
wire v_19026;
wire v_19027;
wire v_19028;
wire v_19029;
wire v_19030;
wire v_19031;
wire v_19032;
wire v_19033;
wire v_19034;
wire v_19035;
wire v_19036;
wire v_19037;
wire v_19038;
wire v_19039;
wire v_19040;
wire v_19041;
wire v_19042;
wire v_19043;
wire v_19044;
wire v_19045;
wire v_19046;
wire v_19047;
wire v_19048;
wire v_19049;
wire v_19050;
wire v_19051;
wire v_19052;
wire v_19053;
wire v_19054;
wire v_19055;
wire v_19056;
wire v_19057;
wire v_19058;
wire v_19059;
wire v_19060;
wire v_19061;
wire v_19062;
wire v_19063;
wire v_19064;
wire v_19065;
wire v_19066;
wire v_19067;
wire v_19068;
wire v_19069;
wire v_19070;
wire v_19071;
wire v_19072;
wire v_19073;
wire v_19074;
wire v_19075;
wire v_19076;
wire v_19077;
wire v_19078;
wire v_19079;
wire v_19080;
wire v_19081;
wire v_19082;
wire v_19083;
wire v_19084;
wire v_19085;
wire v_19086;
wire v_19087;
wire v_19088;
wire v_19089;
wire v_19090;
wire v_19091;
wire v_19092;
wire v_19093;
wire v_19094;
wire v_19095;
wire v_19096;
wire v_19097;
wire v_19098;
wire v_19099;
wire v_19100;
wire v_19101;
wire v_19102;
wire v_19103;
wire v_19104;
wire v_19105;
wire v_19106;
wire v_19107;
wire v_19108;
wire v_19109;
wire v_19110;
wire v_19111;
wire v_19112;
wire v_19113;
wire v_19114;
wire v_19115;
wire v_19116;
wire v_19117;
wire v_19118;
wire v_19119;
wire v_19120;
wire v_19121;
wire v_19122;
wire v_19123;
wire v_19124;
wire v_19125;
wire v_19126;
wire v_19127;
wire v_19128;
wire v_19129;
wire v_19130;
wire v_19131;
wire v_19132;
wire v_19133;
wire v_19134;
wire v_19135;
wire v_19136;
wire v_19137;
wire v_19138;
wire v_19139;
wire v_19140;
wire v_19141;
wire v_19142;
wire v_19143;
wire v_19144;
wire v_19145;
wire v_19146;
wire v_19147;
wire v_19148;
wire v_19149;
wire v_19150;
wire v_19151;
wire v_19152;
wire v_19153;
wire v_19154;
wire v_19155;
wire v_19156;
wire v_19157;
wire v_19158;
wire v_19159;
wire v_19160;
wire v_19161;
wire v_19162;
wire v_19163;
wire v_19164;
wire v_19165;
wire v_19166;
wire v_19167;
wire v_19168;
wire v_19169;
wire v_19170;
wire v_19171;
wire v_19172;
wire v_19173;
wire v_19174;
wire v_19175;
wire v_19176;
wire v_19177;
wire v_19178;
wire v_19179;
wire v_19180;
wire v_19181;
wire v_19182;
wire v_19183;
wire v_19184;
wire v_19185;
wire v_19186;
wire v_19187;
wire v_19188;
wire v_19189;
wire v_19190;
wire v_19191;
wire v_19192;
wire v_19193;
wire v_19194;
wire v_19195;
wire v_19196;
wire v_19197;
wire v_19198;
wire v_19199;
wire v_19200;
wire v_19201;
wire v_19202;
wire v_19203;
wire v_19204;
wire v_19205;
wire v_19206;
wire v_19207;
wire v_19208;
wire v_19209;
wire v_19210;
wire v_19211;
wire v_19212;
wire v_19213;
wire v_19214;
wire v_19215;
wire v_19216;
wire v_19217;
wire v_19218;
wire v_19219;
wire v_19220;
wire v_19221;
wire v_19222;
wire v_19223;
wire v_19224;
wire v_19225;
wire v_19226;
wire v_19227;
wire v_19228;
wire v_19229;
wire v_19230;
wire v_19231;
wire v_19232;
wire v_19233;
wire v_19234;
wire v_19235;
wire v_19236;
wire v_19237;
wire v_19238;
wire v_19239;
wire v_19240;
wire v_19241;
wire v_19242;
wire v_19243;
wire v_19244;
wire v_19245;
wire v_19246;
wire v_19247;
wire v_19248;
wire v_19249;
wire v_19250;
wire v_19251;
wire v_19252;
wire v_19253;
wire v_19254;
wire v_19255;
wire v_19256;
wire v_19257;
wire v_19258;
wire v_19259;
wire v_19260;
wire v_19261;
wire v_19262;
wire v_19263;
wire v_19264;
wire v_19265;
wire v_19266;
wire v_19267;
wire v_19268;
wire v_19269;
wire v_19270;
wire v_19271;
wire v_19272;
wire v_19273;
wire v_19274;
wire v_19275;
wire v_19276;
wire v_19277;
wire v_19278;
wire v_19279;
wire v_19280;
wire v_19281;
wire v_19282;
wire v_19283;
wire v_19284;
wire v_19285;
wire v_19286;
wire v_19287;
wire v_19288;
wire v_19289;
wire v_19290;
wire v_19291;
wire v_19292;
wire v_19293;
wire v_19294;
wire v_19295;
wire v_19296;
wire v_19297;
wire v_19298;
wire v_19299;
wire v_19300;
wire v_19301;
wire v_19302;
wire v_19303;
wire v_19304;
wire v_19305;
wire v_19306;
wire v_19307;
wire v_19308;
wire v_19309;
wire v_19310;
wire v_19311;
wire v_19312;
wire v_19313;
wire v_19314;
wire v_19315;
wire v_19316;
wire v_19317;
wire v_19318;
wire v_19319;
wire v_19320;
wire v_19321;
wire v_19322;
wire v_19323;
wire v_19324;
wire v_19325;
wire v_19326;
wire v_19327;
wire v_19328;
wire v_19329;
wire v_19330;
wire v_19331;
wire v_19332;
wire v_19333;
wire v_19334;
wire v_19335;
wire v_19336;
wire v_19337;
wire v_19338;
wire v_19339;
wire v_19340;
wire v_19341;
wire v_19342;
wire v_19343;
wire v_19344;
wire v_19345;
wire v_19346;
wire v_19347;
wire v_19348;
wire v_19349;
wire v_19350;
wire v_19351;
wire v_19352;
wire v_19353;
wire v_19354;
wire v_19355;
wire v_19356;
wire v_19357;
wire v_19358;
wire v_19359;
wire v_19360;
wire v_19361;
wire v_19362;
wire v_19363;
wire v_19364;
wire v_19365;
wire v_19366;
wire v_19367;
wire v_19368;
wire v_19369;
wire v_19370;
wire v_19371;
wire v_19372;
wire v_19373;
wire v_19374;
wire v_19375;
wire v_19376;
wire v_19377;
wire v_19378;
wire v_19379;
wire v_19380;
wire v_19381;
wire v_19382;
wire v_19383;
wire v_19384;
wire v_19385;
wire v_19386;
wire v_19387;
wire v_19388;
wire v_19389;
wire v_19390;
wire v_19391;
wire v_19392;
wire v_19393;
wire v_19394;
wire v_19395;
wire v_19396;
wire v_19397;
wire v_19398;
wire v_19399;
wire v_19400;
wire v_19401;
wire v_19402;
wire v_19403;
wire v_19404;
wire v_19405;
wire v_19406;
wire v_19407;
wire v_19408;
wire v_19409;
wire v_19410;
wire v_19411;
wire v_19412;
wire v_19413;
wire v_19414;
wire v_19415;
wire v_19416;
wire v_19417;
wire v_19418;
wire v_19419;
wire v_19420;
wire v_19421;
wire v_19422;
wire v_19423;
wire v_19424;
wire v_19425;
wire v_19426;
wire v_19427;
wire v_19428;
wire v_19429;
wire v_19430;
wire v_19431;
wire v_19432;
wire v_19433;
wire v_19434;
wire v_19435;
wire v_19436;
wire v_19437;
wire v_19438;
wire v_19439;
wire v_19440;
wire v_19441;
wire v_19442;
wire v_19443;
wire v_19444;
wire v_19445;
wire v_19446;
wire v_19447;
wire v_19448;
wire v_19449;
wire v_19450;
wire v_19451;
wire v_19452;
wire v_19453;
wire v_19454;
wire v_19455;
wire v_19456;
wire v_19457;
wire v_19458;
wire v_19459;
wire v_19460;
wire v_19461;
wire v_19462;
wire v_19463;
wire v_19464;
wire v_19465;
wire v_19466;
wire v_19467;
wire v_19468;
wire v_19469;
wire v_19470;
wire v_19471;
wire v_19472;
wire v_19473;
wire v_19474;
wire v_19475;
wire v_19476;
wire v_19477;
wire v_19478;
wire v_19479;
wire v_19480;
wire v_19481;
wire v_19482;
wire v_19483;
wire v_19484;
wire v_19485;
wire v_19486;
wire v_19487;
wire v_19488;
wire v_19489;
wire v_19490;
wire v_19491;
wire v_19492;
wire v_19493;
wire v_19494;
wire v_19495;
wire v_19496;
wire v_19497;
wire v_19498;
wire v_19499;
wire v_19500;
wire v_19501;
wire v_19502;
wire v_19503;
wire v_19504;
wire v_19505;
wire v_19506;
wire v_19507;
wire v_19508;
wire v_19509;
wire v_19510;
wire v_19511;
wire v_19512;
wire v_19513;
wire v_19514;
wire v_19515;
wire v_19516;
wire v_19517;
wire v_19518;
wire v_19519;
wire v_19520;
wire v_19521;
wire v_19522;
wire v_19523;
wire v_19524;
wire v_19525;
wire v_19526;
wire v_19527;
wire v_19528;
wire v_19529;
wire v_19530;
wire v_19531;
wire v_19532;
wire v_19533;
wire v_19534;
wire v_19535;
wire v_19536;
wire v_19537;
wire v_19538;
wire v_19539;
wire v_19540;
wire v_19541;
wire v_19542;
wire v_19543;
wire v_19544;
wire v_19545;
wire v_19546;
wire v_19547;
wire v_19548;
wire v_19549;
wire v_19550;
wire v_19551;
wire v_19552;
wire v_19553;
wire v_19554;
wire v_19555;
wire v_19556;
wire v_19557;
wire v_19558;
wire v_19559;
wire v_19560;
wire v_19561;
wire v_19562;
wire v_19563;
wire v_19564;
wire v_19565;
wire v_19566;
wire v_19567;
wire v_19568;
wire v_19569;
wire v_19570;
wire v_19571;
wire v_19572;
wire v_19573;
wire v_19574;
wire v_19575;
wire v_19576;
wire v_19577;
wire v_19578;
wire v_19579;
wire v_19580;
wire v_19581;
wire v_19582;
wire v_19583;
wire v_19584;
wire v_19585;
wire v_19586;
wire v_19587;
wire v_19588;
wire v_19589;
wire v_19590;
wire v_19591;
wire v_19592;
wire v_19593;
wire v_19594;
wire v_19595;
wire v_19596;
wire v_19597;
wire v_19598;
wire v_19599;
wire v_19600;
wire v_19601;
wire v_19602;
wire v_19603;
wire v_19604;
wire v_19605;
wire v_19606;
wire v_19607;
wire v_19608;
wire v_19609;
wire v_19610;
wire v_19611;
wire v_19612;
wire v_19613;
wire v_19614;
wire v_19615;
wire v_19616;
wire v_19617;
wire v_19618;
wire v_19619;
wire v_19620;
wire v_19621;
wire v_19622;
wire v_19623;
wire v_19624;
wire v_19625;
wire v_19626;
wire v_19627;
wire v_19628;
wire v_19629;
wire v_19630;
wire v_19631;
wire v_19632;
wire v_19633;
wire v_19634;
wire v_19635;
wire v_19636;
wire v_19637;
wire v_19638;
wire v_19639;
wire v_19640;
wire v_19641;
wire v_19642;
wire v_19643;
wire v_19644;
wire v_19645;
wire v_19646;
wire v_19647;
wire v_19648;
wire v_19649;
wire v_19650;
wire v_19651;
wire v_19652;
wire v_19653;
wire v_19654;
wire v_19655;
wire v_19656;
wire v_19657;
wire v_19658;
wire v_19659;
wire v_19660;
wire v_19661;
wire v_19662;
wire v_19663;
wire v_19664;
wire v_19665;
wire v_19666;
wire v_19667;
wire v_19668;
wire v_19669;
wire v_19670;
wire v_19671;
wire v_19672;
wire v_19673;
wire v_19674;
wire v_19675;
wire v_19676;
wire v_19677;
wire v_19678;
wire v_19679;
wire v_19680;
wire v_19681;
wire v_19682;
wire v_19683;
wire v_19684;
wire v_19685;
wire v_19686;
wire v_19687;
wire v_19688;
wire v_19689;
wire v_19690;
wire v_19691;
wire v_19692;
wire v_19693;
wire v_19694;
wire v_19695;
wire v_19696;
wire v_19697;
wire v_19698;
wire v_19699;
wire v_19700;
wire v_19701;
wire v_19702;
wire v_19703;
wire v_19704;
wire v_19705;
wire v_19706;
wire v_19707;
wire v_19708;
wire v_19709;
wire v_19710;
wire v_19711;
wire v_19712;
wire v_19713;
wire v_19714;
wire v_19715;
wire v_19716;
wire v_19717;
wire v_19718;
wire v_19719;
wire v_19720;
wire v_19721;
wire v_19722;
wire v_19723;
wire v_19724;
wire v_19725;
wire v_19726;
wire v_19727;
wire v_19728;
wire v_19729;
wire v_19730;
wire v_19731;
wire v_19732;
wire v_19733;
wire v_19734;
wire v_19735;
wire v_19736;
wire v_19737;
wire v_19738;
wire v_19739;
wire v_19740;
wire v_19741;
wire v_19742;
wire v_19743;
wire v_19744;
wire v_19745;
wire v_19746;
wire v_19747;
wire v_19748;
wire v_19749;
wire v_19750;
wire v_19751;
wire v_19752;
wire v_19753;
wire v_19754;
wire v_19755;
wire v_19756;
wire v_19757;
wire v_19758;
wire v_19759;
wire v_19760;
wire v_19761;
wire v_19762;
wire v_19763;
wire v_19764;
wire v_19765;
wire v_19766;
wire v_19767;
wire v_19768;
wire v_19769;
wire v_19770;
wire v_19771;
wire v_19772;
wire v_19773;
wire v_19774;
wire v_19775;
wire v_19776;
wire v_19777;
wire v_19778;
wire v_19779;
wire v_19780;
wire v_19781;
wire v_19782;
wire v_19783;
wire v_19784;
wire v_19785;
wire v_19786;
wire v_19787;
wire v_19788;
wire v_19789;
wire v_19790;
wire v_19791;
wire v_19792;
wire v_19793;
wire v_19794;
wire v_19795;
wire v_19796;
wire v_19797;
wire v_19798;
wire v_19799;
wire v_19800;
wire v_19801;
wire v_19802;
wire v_19803;
wire v_19804;
wire v_19805;
wire v_19806;
wire v_19807;
wire v_19808;
wire v_19809;
wire v_19810;
wire v_19811;
wire v_19812;
wire v_19813;
wire v_19814;
wire v_19815;
wire v_19816;
wire v_19817;
wire v_19818;
wire v_19819;
wire v_19820;
wire v_19821;
wire v_19822;
wire v_19823;
wire v_19824;
wire v_19825;
wire v_19826;
wire v_19827;
wire v_19828;
wire v_19829;
wire v_19830;
wire v_19831;
wire v_19832;
wire v_19833;
wire v_19834;
wire v_19835;
wire v_19836;
wire v_19837;
wire v_19838;
wire v_19839;
wire v_19840;
wire v_19841;
wire v_19842;
wire v_19843;
wire v_19844;
wire v_19845;
wire v_19846;
wire v_19847;
wire v_19848;
wire v_19849;
wire v_19850;
wire v_19851;
wire v_19852;
wire v_19853;
wire v_19854;
wire v_19855;
wire v_19856;
wire v_19857;
wire v_19858;
wire v_19859;
wire v_19860;
wire v_19861;
wire v_19862;
wire v_19863;
wire v_19864;
wire v_19865;
wire v_19866;
wire v_19867;
wire v_19868;
wire v_19869;
wire v_19870;
wire v_19871;
wire v_19872;
wire v_19873;
wire v_19874;
wire v_19875;
wire v_19876;
wire v_19877;
wire v_19878;
wire v_19879;
wire v_19880;
wire v_19881;
wire v_19882;
wire v_19883;
wire v_19884;
wire v_19885;
wire v_19886;
wire v_19887;
wire v_19888;
wire v_19889;
wire v_19890;
wire v_19891;
wire v_19892;
wire v_19893;
wire v_19894;
wire v_19895;
wire v_19896;
wire v_19897;
wire v_19898;
wire v_19899;
wire v_19900;
wire v_19901;
wire v_19902;
wire v_19903;
wire v_19904;
wire v_19905;
wire v_19906;
wire v_19907;
wire v_19908;
wire v_19909;
wire v_19910;
wire v_19911;
wire v_19912;
wire v_19913;
wire v_19914;
wire v_19915;
wire v_19916;
wire v_19917;
wire v_19918;
wire v_19919;
wire v_19920;
wire v_19921;
wire v_19922;
wire v_19923;
wire v_19924;
wire v_19925;
wire v_19926;
wire v_19927;
wire v_19928;
wire v_19929;
wire v_19930;
wire v_19931;
wire v_19932;
wire v_19933;
wire v_19934;
wire v_19935;
wire v_19936;
wire v_19937;
wire v_19938;
wire v_19939;
wire v_19940;
wire v_19941;
wire v_19942;
wire v_19943;
wire v_19944;
wire v_19945;
wire v_19946;
wire v_19947;
wire v_19948;
wire v_19949;
wire v_19950;
wire v_19951;
wire v_19952;
wire v_19953;
wire v_19954;
wire v_19955;
wire v_19956;
wire v_19957;
wire v_19958;
wire v_19959;
wire v_19960;
wire v_19961;
wire v_19962;
wire v_19963;
wire v_19964;
wire v_19965;
wire v_19966;
wire v_19967;
wire v_19968;
wire v_19969;
wire v_19970;
wire v_19971;
wire v_19972;
wire v_19973;
wire v_19974;
wire v_19975;
wire v_19976;
wire v_19977;
wire v_19978;
wire v_19979;
wire v_19980;
wire v_19981;
wire v_19982;
wire v_19983;
wire v_19984;
wire v_19985;
wire v_19986;
wire v_19987;
wire v_19988;
wire v_19989;
wire v_19990;
wire v_19991;
wire v_19992;
wire v_19993;
wire v_19994;
wire v_19995;
wire v_19996;
wire v_19997;
wire v_19998;
wire v_19999;
wire v_20000;
wire v_20001;
wire v_20002;
wire v_20003;
wire v_20004;
wire v_20005;
wire v_20006;
wire v_20007;
wire v_20008;
wire v_20009;
wire v_20010;
wire v_20011;
wire v_20012;
wire v_20013;
wire v_20014;
wire v_20015;
wire v_20016;
wire v_20017;
wire v_20018;
wire v_20019;
wire v_20020;
wire v_20021;
wire v_20022;
wire v_20023;
wire v_20024;
wire v_20025;
wire v_20026;
wire v_20027;
wire v_20028;
wire v_20029;
wire v_20030;
wire v_20031;
wire v_20032;
wire v_20033;
wire v_20034;
wire v_20035;
wire v_20036;
wire v_20037;
wire v_20038;
wire v_20039;
wire v_20040;
wire v_20041;
wire v_20042;
wire v_20043;
wire v_20044;
wire v_20045;
wire v_20046;
wire v_20047;
wire v_20048;
wire v_20049;
wire v_20050;
wire v_20051;
wire v_20052;
wire v_20053;
wire v_20054;
wire v_20055;
wire v_20056;
wire v_20057;
wire v_20058;
wire v_20059;
wire v_20060;
wire v_20061;
wire v_20062;
wire v_20063;
wire v_20064;
wire v_20065;
wire v_20066;
wire v_20067;
wire v_20068;
wire v_20069;
wire v_20070;
wire v_20071;
wire v_20072;
wire v_20073;
wire v_20074;
wire v_20075;
wire v_20076;
wire v_20077;
wire v_20078;
wire v_20079;
wire v_20080;
wire v_20081;
wire v_20082;
wire v_20083;
wire v_20084;
wire v_20085;
wire v_20086;
wire v_20087;
wire v_20088;
wire v_20089;
wire v_20090;
wire v_20091;
wire v_20092;
wire v_20093;
wire v_20094;
wire v_20095;
wire v_20096;
wire v_20097;
wire v_20098;
wire v_20099;
wire v_20100;
wire v_20101;
wire v_20102;
wire v_20103;
wire v_20104;
wire v_20105;
wire v_20106;
wire v_20107;
wire v_20108;
wire v_20109;
wire v_20110;
wire v_20111;
wire v_20112;
wire v_20113;
wire v_20114;
wire v_20115;
wire v_20116;
wire v_20117;
wire v_20118;
wire v_20119;
wire v_20120;
wire v_20121;
wire v_20122;
wire v_20123;
wire v_20124;
wire v_20125;
wire v_20126;
wire v_20127;
wire v_20128;
wire v_20129;
wire v_20130;
wire v_20131;
wire v_20132;
wire v_20133;
wire v_20134;
wire v_20135;
wire v_20136;
wire v_20137;
wire v_20138;
wire v_20139;
wire v_20140;
wire v_20141;
wire v_20142;
wire v_20143;
wire v_20144;
wire v_20145;
wire v_20146;
wire v_20147;
wire v_20148;
wire v_20149;
wire v_20150;
wire v_20151;
wire v_20152;
wire v_20153;
wire v_20154;
wire v_20155;
wire v_20156;
wire v_20157;
wire v_20158;
wire v_20159;
wire v_20160;
wire v_20161;
wire v_20162;
wire v_20163;
wire v_20164;
wire v_20165;
wire v_20166;
wire v_20167;
wire v_20168;
wire v_20169;
wire v_20170;
wire v_20171;
wire v_20172;
wire v_20173;
wire v_20174;
wire v_20175;
wire v_20176;
wire v_20177;
wire v_20178;
wire v_20179;
wire v_20180;
wire v_20181;
wire v_20182;
wire v_20183;
wire v_20184;
wire v_20185;
wire v_20186;
wire v_20187;
wire v_20188;
wire v_20189;
wire v_20190;
wire v_20191;
wire v_20192;
wire v_20193;
wire v_20194;
wire v_20195;
wire v_20196;
wire v_20197;
wire v_20198;
wire v_20199;
wire v_20200;
wire v_20201;
wire v_20202;
wire v_20203;
wire v_20204;
wire v_20205;
wire v_20206;
wire v_20207;
wire v_20208;
wire v_20209;
wire v_20210;
wire v_20211;
wire v_20212;
wire v_20213;
wire v_20214;
wire v_20215;
wire v_20216;
wire v_20217;
wire v_20218;
wire v_20219;
wire v_20220;
wire v_20221;
wire v_20222;
wire v_20223;
wire v_20224;
wire v_20225;
wire v_20226;
wire v_20227;
wire v_20228;
wire v_20229;
wire v_20230;
wire v_20231;
wire v_20232;
wire v_20233;
wire v_20234;
wire v_20235;
wire v_20236;
wire v_20237;
wire v_20238;
wire v_20239;
wire v_20240;
wire v_20241;
wire v_20242;
wire v_20243;
wire v_20244;
wire v_20245;
wire v_20246;
wire v_20247;
wire v_20248;
wire v_20249;
wire v_20250;
wire v_20251;
wire v_20252;
wire v_20253;
wire v_20254;
wire v_20255;
wire v_20256;
wire v_20257;
wire v_20258;
wire v_20259;
wire v_20260;
wire v_20261;
wire v_20262;
wire v_20263;
wire v_20264;
wire v_20265;
wire v_20266;
wire v_20267;
wire v_20268;
wire v_20269;
wire v_20270;
wire v_20271;
wire v_20272;
wire v_20273;
wire v_20274;
wire v_20275;
wire v_20276;
wire v_20277;
wire v_20278;
wire v_20279;
wire v_20280;
wire v_20281;
wire v_20282;
wire v_20283;
wire v_20284;
wire v_20285;
wire v_20286;
wire v_20287;
wire v_20288;
wire v_20289;
wire v_20290;
wire v_20291;
wire v_20292;
wire v_20293;
wire v_20294;
wire v_20295;
wire v_20296;
wire v_20297;
wire v_20298;
wire v_20299;
wire v_20300;
wire v_20301;
wire v_20302;
wire v_20303;
wire v_20304;
wire v_20305;
wire v_20306;
wire v_20307;
wire v_20308;
wire v_20309;
wire v_20310;
wire v_20311;
wire v_20312;
wire v_20313;
wire v_20314;
wire v_20315;
wire v_20316;
wire v_20317;
wire v_20318;
wire v_20319;
wire v_20320;
wire v_20321;
wire v_20322;
wire v_20323;
wire v_20324;
wire v_20325;
wire v_20326;
wire v_20327;
wire v_20328;
wire v_20329;
wire v_20330;
wire v_20331;
wire v_20332;
wire v_20333;
wire v_20334;
wire v_20335;
wire v_20336;
wire v_20337;
wire v_20338;
wire v_20339;
wire v_20340;
wire v_20341;
wire v_20342;
wire v_20343;
wire v_20344;
wire v_20345;
wire v_20346;
wire v_20347;
wire v_20348;
wire v_20349;
wire v_20350;
wire v_20351;
wire v_20352;
wire v_20353;
wire v_20354;
wire v_20355;
wire v_20356;
wire v_20357;
wire v_20358;
wire v_20359;
wire v_20360;
wire v_20361;
wire v_20362;
wire v_20363;
wire v_20364;
wire v_20365;
wire v_20366;
wire v_20367;
wire v_20368;
wire v_20369;
wire v_20370;
wire v_20371;
wire v_20372;
wire v_20373;
wire v_20374;
wire v_20375;
wire v_20376;
wire v_20377;
wire v_20378;
wire v_20379;
wire v_20380;
wire v_20381;
wire v_20382;
wire v_20383;
wire v_20384;
wire v_20385;
wire v_20386;
wire v_20387;
wire v_20388;
wire v_20389;
wire v_20390;
wire v_20391;
wire v_20392;
wire v_20393;
wire v_20394;
wire v_20395;
wire v_20396;
wire v_20397;
wire v_20398;
wire v_20399;
wire v_20400;
wire v_20401;
wire v_20402;
wire v_20403;
wire v_20404;
wire v_20405;
wire v_20406;
wire v_20407;
wire v_20408;
wire v_20409;
wire v_20410;
wire v_20411;
wire v_20412;
wire v_20413;
wire v_20414;
wire v_20415;
wire v_20416;
wire v_20417;
wire v_20418;
wire v_20419;
wire v_20420;
wire v_20421;
wire v_20422;
wire v_20423;
wire v_20424;
wire v_20425;
wire v_20426;
wire v_20427;
wire v_20428;
wire v_20429;
wire v_20430;
wire v_20431;
wire v_20432;
wire v_20433;
wire v_20434;
wire v_20435;
wire v_20436;
wire v_20437;
wire v_20438;
wire v_20439;
wire v_20440;
wire v_20441;
wire v_20442;
wire v_20443;
wire v_20444;
wire v_20445;
wire v_20446;
wire v_20447;
wire v_20448;
wire v_20449;
wire v_20450;
wire v_20451;
wire v_20452;
wire v_20453;
wire v_20454;
wire v_20455;
wire v_20456;
wire v_20457;
wire v_20458;
wire v_20459;
wire v_20460;
wire v_20461;
wire v_20462;
wire v_20463;
wire v_20464;
wire v_20465;
wire v_20466;
wire v_20467;
wire v_20468;
wire v_20469;
wire v_20470;
wire v_20471;
wire v_20472;
wire v_20473;
wire v_20474;
wire v_20475;
wire v_20476;
wire v_20477;
wire v_20478;
wire v_20479;
wire v_20480;
wire v_20481;
wire v_20482;
wire v_20483;
wire v_20484;
wire v_20485;
wire v_20486;
wire v_20487;
wire v_20488;
wire v_20489;
wire v_20490;
wire v_20491;
wire v_20492;
wire v_20493;
wire v_20494;
wire v_20495;
wire v_20496;
wire v_20497;
wire v_20498;
wire v_20499;
wire v_20500;
wire v_20501;
wire v_20502;
wire v_20503;
wire v_20504;
wire v_20505;
wire v_20506;
wire v_20507;
wire v_20508;
wire v_20509;
wire v_20510;
wire v_20511;
wire v_20512;
wire v_20513;
wire v_20514;
wire v_20515;
wire v_20516;
wire v_20517;
wire v_20518;
wire v_20519;
wire v_20520;
wire v_20521;
wire v_20522;
wire v_20523;
wire v_20524;
wire v_20525;
wire v_20526;
wire v_20527;
wire v_20528;
wire v_20529;
wire v_20530;
wire v_20531;
wire v_20532;
wire v_20533;
wire v_20534;
wire v_20535;
wire v_20536;
wire v_20537;
wire v_20538;
wire v_20539;
wire v_20540;
wire v_20541;
wire v_20542;
wire v_20543;
wire v_20544;
wire v_20545;
wire v_20546;
wire v_20547;
wire v_20548;
wire v_20549;
wire v_20550;
wire v_20551;
wire v_20552;
wire v_20553;
wire v_20554;
wire v_20555;
wire v_20556;
wire v_20557;
wire v_20558;
wire v_20559;
wire v_20560;
wire v_20561;
wire v_20562;
wire v_20563;
wire v_20564;
wire v_20565;
wire v_20566;
wire v_20567;
wire v_20568;
wire v_20569;
wire v_20570;
wire v_20571;
wire v_20572;
wire v_20573;
wire v_20574;
wire v_20575;
wire v_20576;
wire v_20577;
wire v_20578;
wire v_20579;
wire v_20580;
wire v_20581;
wire v_20582;
wire v_20583;
wire v_20584;
wire v_20585;
wire v_20586;
wire v_20587;
wire v_20588;
wire v_20589;
wire v_20590;
wire v_20591;
wire v_20592;
wire v_20593;
wire v_20594;
wire v_20595;
wire v_20596;
wire v_20597;
wire v_20598;
wire v_20599;
wire v_20600;
wire v_20601;
wire v_20602;
wire v_20603;
wire v_20604;
wire v_20605;
wire v_20606;
wire v_20607;
wire v_20608;
wire v_20609;
wire v_20610;
wire v_20611;
wire v_20612;
wire v_20613;
wire v_20614;
wire v_20615;
wire v_20616;
wire v_20617;
wire v_20618;
wire v_20619;
wire v_20620;
wire v_20621;
wire v_20622;
wire v_20623;
wire v_20624;
wire v_20625;
wire v_20626;
wire v_20627;
wire v_20628;
wire v_20629;
wire v_20630;
wire v_20631;
wire v_20632;
wire v_20633;
wire v_20634;
wire v_20635;
wire v_20636;
wire v_20637;
wire v_20638;
wire v_20639;
wire v_20640;
wire v_20641;
wire v_20642;
wire v_20643;
wire v_20644;
wire v_20645;
wire v_20646;
wire v_20647;
wire v_20648;
wire v_20649;
wire v_20650;
wire v_20651;
wire v_20652;
wire v_20653;
wire v_20654;
wire v_20655;
wire v_20656;
wire v_20657;
wire v_20658;
wire v_20659;
wire v_20660;
wire v_20661;
wire v_20662;
wire v_20663;
wire v_20664;
wire v_20665;
wire v_20666;
wire v_20667;
wire v_20668;
wire v_20669;
wire v_20670;
wire v_20671;
wire v_20672;
wire v_20673;
wire v_20674;
wire v_20675;
wire v_20676;
wire v_20677;
wire v_20678;
wire v_20679;
wire v_20680;
wire v_20681;
wire v_20682;
wire v_20683;
wire v_20684;
wire v_20685;
wire v_20686;
wire v_20687;
wire v_20688;
wire v_20689;
wire v_20690;
wire v_20691;
wire v_20692;
wire v_20693;
wire v_20694;
wire v_20695;
wire v_20696;
wire v_20697;
wire v_20698;
wire v_20699;
wire v_20700;
wire v_20701;
wire v_20702;
wire v_20703;
wire v_20704;
wire v_20705;
wire v_20706;
wire v_20707;
wire v_20708;
wire v_20709;
wire v_20710;
wire v_20711;
wire v_20712;
wire v_20713;
wire v_20714;
wire v_20715;
wire v_20716;
wire v_20717;
wire v_20718;
wire v_20719;
wire v_20720;
wire v_20721;
wire v_20722;
wire v_20723;
wire v_20724;
wire v_20725;
wire v_20726;
wire v_20727;
wire v_20728;
wire v_20729;
wire v_20730;
wire v_20731;
wire v_20732;
wire v_20733;
wire v_20734;
wire v_20735;
wire v_20736;
wire v_20737;
wire v_20738;
wire v_20739;
wire v_20740;
wire v_20741;
wire v_20742;
wire v_20743;
wire v_20744;
wire v_20745;
wire v_20746;
wire v_20747;
wire v_20748;
wire v_20749;
wire v_20750;
wire v_20751;
wire v_20752;
wire v_20753;
wire v_20754;
wire v_20755;
wire v_20756;
wire v_20757;
wire v_20758;
wire v_20759;
wire v_20760;
wire v_20761;
wire v_20762;
wire v_20763;
wire v_20764;
wire v_20765;
wire v_20766;
wire v_20767;
wire v_20768;
wire v_20769;
wire v_20770;
wire v_20771;
wire v_20772;
wire v_20773;
wire v_20774;
wire v_20775;
wire v_20776;
wire v_20777;
wire v_20778;
wire v_20779;
wire v_20780;
wire v_20781;
wire v_20782;
wire v_20783;
wire v_20784;
wire v_20785;
wire v_20786;
wire v_20787;
wire v_20788;
wire v_20789;
wire v_20790;
wire v_20791;
wire v_20792;
wire v_20793;
wire v_20794;
wire v_20795;
wire v_20796;
wire v_20797;
wire v_20798;
wire v_20799;
wire v_20800;
wire v_20801;
wire v_20802;
wire v_20803;
wire v_20804;
wire v_20805;
wire v_20806;
wire v_20807;
wire v_20808;
wire v_20809;
wire v_20810;
wire v_20811;
wire v_20812;
wire v_20813;
wire v_20814;
wire v_20815;
wire v_20816;
wire v_20817;
wire v_20818;
wire v_20819;
wire v_20820;
wire v_20821;
wire v_20822;
wire v_20823;
wire v_20824;
wire v_20825;
wire v_20826;
wire v_20827;
wire v_20828;
wire v_20829;
wire v_20830;
wire v_20831;
wire v_20832;
wire v_20833;
wire v_20834;
wire v_20835;
wire v_20836;
wire v_20837;
wire v_20838;
wire v_20839;
wire v_20840;
wire v_20841;
wire v_20842;
wire v_20843;
wire v_20844;
wire v_20845;
wire v_20846;
wire v_20847;
wire v_20848;
wire v_20849;
wire v_20850;
wire v_20851;
wire v_20852;
wire v_20853;
wire v_20854;
wire v_20855;
wire v_20856;
wire v_20857;
wire v_20858;
wire v_20859;
wire v_20860;
wire v_20861;
wire v_20862;
wire v_20863;
wire v_20864;
wire v_20865;
wire v_20866;
wire v_20867;
wire v_20868;
wire v_20869;
wire v_20870;
wire v_20871;
wire v_20872;
wire v_20873;
wire v_20874;
wire v_20875;
wire v_20876;
wire v_20877;
wire v_20878;
wire v_20879;
wire v_20880;
wire v_20881;
wire v_20882;
wire v_20883;
wire v_20884;
wire v_20885;
wire v_20886;
wire v_20887;
wire v_20888;
wire v_20889;
wire v_20890;
wire v_20891;
wire v_20892;
wire v_20893;
wire v_20894;
wire v_20895;
wire v_20896;
wire v_20897;
wire v_20898;
wire v_20899;
wire v_20900;
wire v_20901;
wire v_20902;
wire v_20903;
wire v_20904;
wire v_20905;
wire v_20906;
wire v_20907;
wire v_20908;
wire v_20909;
wire v_20910;
wire v_20911;
wire v_20912;
wire v_20913;
wire v_20914;
wire v_20915;
wire v_20916;
wire v_20917;
wire v_20918;
wire v_20919;
wire v_20920;
wire v_20921;
wire v_20922;
wire v_20923;
wire v_20924;
wire v_20925;
wire v_20926;
wire v_20927;
wire v_20928;
wire v_20929;
wire v_20930;
wire v_20931;
wire v_20932;
wire v_20933;
wire v_20934;
wire v_20935;
wire v_20936;
wire v_20937;
wire v_20938;
wire v_20939;
wire v_20940;
wire v_20941;
wire v_20942;
wire v_20943;
wire v_20944;
wire v_20945;
wire v_20946;
wire v_20947;
wire v_20948;
wire v_20949;
wire v_20950;
wire v_20951;
wire v_20952;
wire v_20953;
wire v_20954;
wire v_20955;
wire v_20956;
wire v_20957;
wire v_20958;
wire v_20959;
wire v_20960;
wire v_20961;
wire v_20962;
wire v_20963;
wire v_20964;
wire v_20965;
wire v_20966;
wire v_20967;
wire v_20968;
wire v_20969;
wire v_20970;
wire v_20971;
wire v_20972;
wire v_20973;
wire v_20974;
wire v_20975;
wire v_20976;
wire v_20977;
wire v_20978;
wire v_20979;
wire v_20980;
wire v_20981;
wire v_20982;
wire v_20983;
wire v_20984;
wire v_20985;
wire v_20986;
wire v_20987;
wire v_20988;
wire v_20989;
wire v_20990;
wire v_20991;
wire v_20992;
wire v_20993;
wire v_20994;
wire v_20995;
wire v_20996;
wire v_20997;
wire v_20998;
wire v_20999;
wire v_21000;
wire v_21001;
wire v_21002;
wire v_21003;
wire v_21004;
wire v_21005;
wire v_21006;
wire v_21007;
wire v_21008;
wire v_21009;
wire v_21010;
wire v_21011;
wire v_21012;
wire v_21013;
wire v_21014;
wire v_21015;
wire v_21016;
wire v_21017;
wire v_21018;
wire v_21019;
wire v_21020;
wire v_21021;
wire v_21022;
wire v_21023;
wire v_21024;
wire v_21025;
wire v_21026;
wire v_21027;
wire v_21028;
wire v_21029;
wire v_21030;
wire v_21031;
wire v_21032;
wire v_21033;
wire v_21034;
wire v_21035;
wire v_21036;
wire v_21037;
wire v_21038;
wire v_21039;
wire v_21040;
wire v_21041;
wire v_21042;
wire v_21043;
wire v_21044;
wire v_21045;
wire v_21046;
wire v_21047;
wire v_21048;
wire v_21049;
wire v_21050;
wire v_21051;
wire v_21052;
wire v_21053;
wire v_21054;
wire v_21055;
wire v_21056;
wire v_21057;
wire v_21058;
wire v_21059;
wire v_21060;
wire v_21061;
wire v_21062;
wire v_21063;
wire v_21064;
wire v_21065;
wire v_21066;
wire v_21067;
wire v_21068;
wire v_21069;
wire v_21070;
wire v_21071;
wire v_21072;
wire v_21073;
wire v_21074;
wire v_21075;
wire v_21076;
wire v_21077;
wire v_21078;
wire v_21079;
wire v_21080;
wire v_21081;
wire v_21082;
wire v_21083;
wire v_21084;
wire v_21085;
wire v_21086;
wire v_21087;
wire v_21088;
wire v_21089;
wire v_21090;
wire v_21091;
wire v_21092;
wire v_21093;
wire v_21094;
wire v_21095;
wire v_21096;
wire v_21097;
wire v_21098;
wire v_21099;
wire v_21100;
wire v_21101;
wire v_21102;
wire v_21103;
wire v_21104;
wire v_21105;
wire v_21106;
wire v_21107;
wire v_21108;
wire v_21109;
wire v_21110;
wire v_21111;
wire v_21112;
wire v_21113;
wire v_21114;
wire v_21115;
wire v_21116;
wire v_21117;
wire v_21118;
wire v_21119;
wire v_21120;
wire v_21121;
wire v_21122;
wire v_21123;
wire v_21124;
wire v_21125;
wire v_21126;
wire v_21127;
wire v_21128;
wire v_21129;
wire v_21130;
wire v_21131;
wire v_21132;
wire v_21133;
wire v_21134;
wire v_21135;
wire v_21136;
wire v_21137;
wire v_21138;
wire v_21139;
wire v_21140;
wire v_21141;
wire v_21142;
wire v_21143;
wire v_21144;
wire v_21145;
wire v_21146;
wire v_21147;
wire v_21148;
wire v_21149;
wire v_21150;
wire v_21151;
wire v_21152;
wire v_21153;
wire v_21154;
wire v_21155;
wire v_21156;
wire v_21157;
wire v_21158;
wire v_21159;
wire v_21160;
wire v_21161;
wire v_21162;
wire v_21163;
wire v_21164;
wire v_21165;
wire v_21166;
wire v_21167;
wire v_21168;
wire v_21169;
wire v_21170;
wire v_21171;
wire v_21172;
wire v_21173;
wire v_21174;
wire v_21175;
wire v_21176;
wire v_21177;
wire v_21178;
wire v_21179;
wire v_21180;
wire v_21181;
wire v_21182;
wire v_21183;
wire v_21184;
wire v_21185;
wire v_21186;
wire v_21187;
wire v_21188;
wire v_21189;
wire v_21190;
wire v_21191;
wire v_21192;
wire v_21193;
wire v_21194;
wire v_21195;
wire v_21196;
wire v_21197;
wire v_21198;
wire v_21199;
wire v_21200;
wire v_21201;
wire v_21202;
wire v_21203;
wire v_21204;
wire v_21205;
wire v_21206;
wire v_21207;
wire v_21208;
wire v_21209;
wire v_21210;
wire v_21211;
wire v_21212;
wire v_21213;
wire v_21214;
wire v_21215;
wire v_21216;
wire v_21217;
wire v_21218;
wire v_21219;
wire v_21220;
wire v_21221;
wire v_21222;
wire v_21223;
wire v_21224;
wire v_21225;
wire v_21226;
wire v_21227;
wire v_21228;
wire v_21229;
wire v_21230;
wire v_21231;
wire v_21232;
wire v_21233;
wire v_21234;
wire v_21235;
wire v_21236;
wire v_21237;
wire v_21238;
wire v_21239;
wire v_21240;
wire v_21241;
wire v_21242;
wire v_21243;
wire v_21244;
wire v_21245;
wire v_21246;
wire v_21247;
wire v_21248;
wire v_21249;
wire v_21250;
wire v_21251;
wire v_21252;
wire v_21253;
wire v_21254;
wire v_21255;
wire v_21256;
wire v_21257;
wire v_21258;
wire v_21259;
wire v_21260;
wire v_21261;
wire v_21262;
wire v_21263;
wire v_21264;
wire v_21265;
wire v_21266;
wire v_21267;
wire v_21268;
wire v_21269;
wire v_21270;
wire v_21271;
wire v_21272;
wire v_21273;
wire v_21274;
wire v_21275;
wire v_21276;
wire v_21277;
wire v_21278;
wire v_21279;
wire v_21280;
wire v_21281;
wire v_21282;
wire v_21283;
wire v_21284;
wire v_21285;
wire v_21286;
wire v_21287;
wire v_21288;
wire v_21289;
wire v_21290;
wire v_21291;
wire v_21292;
wire v_21293;
wire v_21294;
wire v_21295;
wire v_21296;
wire v_21297;
wire v_21298;
wire v_21299;
wire v_21300;
wire v_21301;
wire v_21302;
wire v_21303;
wire v_21304;
wire v_21305;
wire v_21306;
wire v_21307;
wire v_21308;
wire v_21309;
wire v_21310;
wire v_21311;
wire v_21312;
wire v_21313;
wire v_21314;
wire v_21315;
wire v_21316;
wire v_21317;
wire v_21318;
wire v_21319;
wire v_21320;
wire v_21321;
wire v_21322;
wire v_21323;
wire v_21324;
wire v_21325;
wire v_21326;
wire v_21327;
wire v_21328;
wire v_21329;
wire v_21330;
wire v_21331;
wire v_21332;
wire v_21333;
wire v_21334;
wire v_21335;
wire v_21336;
wire v_21337;
wire v_21338;
wire v_21339;
wire v_21340;
wire v_21341;
wire v_21342;
wire v_21343;
wire v_21344;
wire v_21345;
wire v_21346;
wire v_21347;
wire v_21348;
wire v_21349;
wire v_21350;
wire v_21351;
wire v_21352;
wire v_21353;
wire v_21354;
wire v_21355;
wire v_21356;
wire v_21357;
wire v_21358;
wire v_21359;
wire v_21360;
wire v_21361;
wire v_21362;
wire v_21363;
wire v_21364;
wire v_21365;
wire v_21366;
wire v_21367;
wire v_21368;
wire v_21369;
wire v_21370;
wire v_21371;
wire v_21372;
wire v_21373;
wire v_21374;
wire v_21375;
wire v_21376;
wire v_21377;
wire v_21378;
wire v_21379;
wire v_21380;
wire v_21381;
wire v_21382;
wire v_21383;
wire v_21384;
wire v_21385;
wire v_21386;
wire v_21387;
wire v_21388;
wire v_21389;
wire v_21390;
wire v_21391;
wire v_21392;
wire v_21393;
wire v_21394;
wire v_21395;
wire v_21396;
wire v_21397;
wire v_21398;
wire v_21399;
wire v_21400;
wire v_21401;
wire v_21402;
wire v_21403;
wire v_21404;
wire v_21405;
wire v_21406;
wire v_21407;
wire v_21408;
wire v_21409;
wire v_21410;
wire v_21411;
wire v_21412;
wire v_21413;
wire v_21414;
wire v_21415;
wire v_21416;
wire v_21417;
wire v_21418;
wire v_21419;
wire v_21420;
wire v_21421;
wire v_21422;
wire v_21423;
wire v_21424;
wire v_21425;
wire v_21426;
wire v_21427;
wire v_21428;
wire v_21429;
wire v_21430;
wire v_21431;
wire v_21432;
wire v_21433;
wire v_21434;
wire v_21435;
wire v_21436;
wire v_21437;
wire v_21438;
wire v_21439;
wire v_21440;
wire v_21441;
wire v_21442;
wire v_21443;
wire v_21444;
wire v_21445;
wire v_21446;
wire v_21447;
wire v_21448;
wire v_21449;
wire v_21450;
wire v_21451;
wire v_21452;
wire v_21453;
wire v_21454;
wire v_21455;
wire v_21456;
wire v_21457;
wire v_21458;
wire v_21459;
wire v_21460;
wire v_21461;
wire v_21462;
wire v_21463;
wire v_21464;
wire v_21465;
wire v_21466;
wire v_21467;
wire v_21468;
wire v_21469;
wire v_21470;
wire v_21471;
wire v_21472;
wire v_21473;
wire v_21474;
wire v_21475;
wire v_21476;
wire v_21477;
wire v_21478;
wire v_21479;
wire v_21480;
wire v_21481;
wire v_21482;
wire v_21483;
wire v_21484;
wire v_21485;
wire v_21486;
wire v_21487;
wire v_21488;
wire v_21489;
wire v_21490;
wire v_21491;
wire v_21492;
wire v_21493;
wire v_21494;
wire v_21495;
wire v_21496;
wire v_21497;
wire v_21498;
wire v_21499;
wire v_21500;
wire v_21501;
wire v_21502;
wire v_21503;
wire v_21504;
wire v_21505;
wire v_21506;
wire v_21507;
wire v_21508;
wire v_21509;
wire v_21510;
wire v_21511;
wire v_21512;
wire v_21513;
wire v_21514;
wire v_21515;
wire v_21516;
wire v_21517;
wire v_21518;
wire v_21519;
wire v_21520;
wire v_21521;
wire v_21522;
wire v_21523;
wire v_21524;
wire v_21525;
wire v_21526;
wire v_21527;
wire v_21528;
wire v_21529;
wire v_21530;
wire v_21531;
wire v_21532;
wire v_21533;
wire v_21534;
wire v_21535;
wire v_21536;
wire v_21537;
wire v_21538;
wire v_21539;
wire v_21540;
wire v_21541;
wire v_21542;
wire v_21543;
wire v_21544;
wire v_21545;
wire v_21546;
wire v_21547;
wire v_21548;
wire v_21549;
wire v_21550;
wire v_21551;
wire v_21552;
wire v_21553;
wire v_21554;
wire v_21555;
wire v_21556;
wire v_21557;
wire v_21558;
wire v_21559;
wire v_21560;
wire v_21561;
wire v_21562;
wire v_21563;
wire v_21564;
wire v_21565;
wire v_21566;
wire v_21567;
wire v_21568;
wire v_21569;
wire v_21570;
wire v_21571;
wire v_21572;
wire v_21573;
wire v_21574;
wire v_21575;
wire v_21576;
wire v_21577;
wire v_21578;
wire v_21579;
wire v_21580;
wire v_21581;
wire v_21582;
wire v_21583;
wire v_21584;
wire v_21585;
wire v_21586;
wire v_21587;
wire v_21588;
wire v_21589;
wire v_21590;
wire v_21591;
wire v_21592;
wire v_21593;
wire v_21594;
wire v_21595;
wire v_21596;
wire v_21597;
wire v_21598;
wire v_21599;
wire v_21600;
wire v_21601;
wire v_21602;
wire v_21603;
wire v_21604;
wire v_21605;
wire v_21606;
wire v_21607;
wire v_21608;
wire v_21609;
wire v_21610;
wire v_21611;
wire v_21612;
wire v_21613;
wire v_21614;
wire v_21615;
wire v_21616;
wire v_21617;
wire v_21618;
wire v_21619;
wire v_21620;
wire v_21621;
wire v_21622;
wire v_21623;
wire v_21624;
wire v_21625;
wire v_21626;
wire v_21627;
wire v_21628;
wire v_21629;
wire v_21630;
wire v_21631;
wire v_21632;
wire v_21633;
wire v_21634;
wire v_21635;
wire v_21636;
wire v_21637;
wire v_21638;
wire v_21639;
wire v_21640;
wire v_21641;
wire v_21642;
wire v_21643;
wire v_21644;
wire v_21645;
wire v_21646;
wire v_21647;
wire v_21648;
wire v_21649;
wire v_21650;
wire v_21651;
wire v_21652;
wire v_21653;
wire v_21654;
wire v_21655;
wire v_21656;
wire v_21657;
wire v_21658;
wire v_21659;
wire v_21660;
wire v_21661;
wire v_21662;
wire v_21663;
wire v_21664;
wire v_21665;
wire v_21666;
wire v_21667;
wire v_21668;
wire v_21669;
wire v_21670;
wire v_21671;
wire v_21672;
wire v_21673;
wire v_21674;
wire v_21675;
wire v_21676;
wire v_21677;
wire v_21678;
wire v_21679;
wire v_21680;
wire v_21681;
wire v_21682;
wire v_21683;
wire v_21684;
wire v_21685;
wire v_21686;
wire v_21687;
wire v_21688;
wire v_21689;
wire v_21690;
wire v_21691;
wire v_21692;
wire v_21693;
wire v_21694;
wire v_21695;
wire v_21696;
wire v_21697;
wire v_21698;
wire v_21699;
wire v_21700;
wire v_21701;
wire v_21702;
wire v_21703;
wire v_21704;
wire v_21705;
wire v_21706;
wire v_21707;
wire v_21708;
wire v_21709;
wire v_21710;
wire v_21711;
wire v_21712;
wire v_21713;
wire v_21714;
wire v_21715;
wire v_21716;
wire v_21717;
wire v_21718;
wire v_21719;
wire v_21720;
wire v_21721;
wire v_21722;
wire v_21723;
wire v_21724;
wire v_21725;
wire v_21726;
wire v_21727;
wire v_21728;
wire v_21729;
wire v_21730;
wire v_21731;
wire v_21732;
wire v_21733;
wire v_21734;
wire v_21735;
wire v_21736;
wire v_21737;
wire v_21738;
wire v_21739;
wire v_21740;
wire v_21741;
wire v_21742;
wire v_21743;
wire v_21744;
wire v_21745;
wire v_21746;
wire v_21747;
wire v_21748;
wire v_21749;
wire v_21750;
wire v_21751;
wire v_21752;
wire v_21753;
wire v_21754;
wire v_21755;
wire v_21756;
wire v_21757;
wire v_21758;
wire v_21759;
wire v_21760;
wire v_21761;
wire v_21762;
wire v_21763;
wire v_21764;
wire v_21765;
wire v_21766;
wire v_21767;
wire v_21768;
wire v_21769;
wire v_21770;
wire v_21771;
wire v_21772;
wire v_21773;
wire v_21774;
wire v_21775;
wire v_21776;
wire v_21777;
wire v_21778;
wire v_21779;
wire v_21780;
wire v_21781;
wire v_21782;
wire v_21783;
wire v_21784;
wire v_21785;
wire v_21786;
wire v_21787;
wire v_21788;
wire v_21789;
wire v_21790;
wire v_21791;
wire v_21792;
wire v_21793;
wire v_21794;
wire v_21795;
wire v_21796;
wire v_21797;
wire v_21798;
wire v_21799;
wire v_21800;
wire v_21801;
wire v_21802;
wire v_21803;
wire v_21804;
wire v_21805;
wire v_21806;
wire v_21807;
wire v_21808;
wire v_21809;
wire v_21810;
wire v_21811;
wire v_21812;
wire v_21813;
wire v_21814;
wire v_21815;
wire v_21816;
wire v_21817;
wire v_21818;
wire v_21819;
wire v_21820;
wire v_21821;
wire v_21822;
wire v_21823;
wire v_21824;
wire v_21825;
wire v_21826;
wire v_21827;
wire v_21828;
wire v_21829;
wire v_21830;
wire v_21831;
wire v_21832;
wire v_21833;
wire v_21834;
wire v_21835;
wire v_21836;
wire v_21837;
wire v_21838;
wire v_21839;
wire v_21840;
wire v_21841;
wire v_21842;
wire v_21843;
wire v_21844;
wire v_21845;
wire v_21846;
wire v_21847;
wire v_21848;
wire v_21849;
wire v_21850;
wire v_21851;
wire v_21852;
wire v_21853;
wire v_21854;
wire v_21855;
wire v_21856;
wire v_21857;
wire v_21858;
wire v_21859;
wire v_21860;
wire v_21861;
wire v_21862;
wire v_21863;
wire v_21864;
wire v_21865;
wire v_21866;
wire v_21867;
wire v_21868;
wire v_21869;
wire v_21870;
wire v_21871;
wire v_21872;
wire v_21873;
wire v_21874;
wire v_21875;
wire v_21876;
wire v_21877;
wire v_21878;
wire v_21879;
wire v_21880;
wire v_21881;
wire v_21882;
wire v_21883;
wire v_21884;
wire v_21885;
wire v_21886;
wire v_21887;
wire v_21888;
wire v_21889;
wire v_21890;
wire v_21891;
wire v_21892;
wire v_21893;
wire v_21894;
wire v_21895;
wire v_21896;
wire v_21897;
wire v_21898;
wire v_21899;
wire v_21900;
wire v_21901;
wire v_21902;
wire v_21903;
wire v_21904;
wire v_21905;
wire v_21906;
wire v_21907;
wire v_21908;
wire v_21909;
wire v_21910;
wire v_21911;
wire v_21912;
wire v_21913;
wire v_21914;
wire v_21915;
wire v_21916;
wire v_21917;
wire v_21918;
wire v_21919;
wire v_21920;
wire v_21921;
wire v_21922;
wire v_21923;
wire v_21924;
wire v_21925;
wire v_21926;
wire v_21927;
wire v_21928;
wire v_21929;
wire v_21930;
wire v_21931;
wire v_21932;
wire v_21933;
wire v_21934;
wire v_21935;
wire v_21936;
wire v_21937;
wire v_21938;
wire v_21939;
wire v_21940;
wire v_21941;
wire v_21942;
wire v_21943;
wire v_21944;
wire v_21945;
wire v_21946;
wire v_21947;
wire v_21948;
wire v_21949;
wire v_21950;
wire v_21951;
wire v_21952;
wire v_21953;
wire v_21954;
wire v_21955;
wire v_21956;
wire v_21957;
wire v_21958;
wire v_21959;
wire v_21960;
wire v_21961;
wire v_21962;
wire v_21963;
wire v_21964;
wire v_21965;
wire v_21966;
wire v_21967;
wire v_21968;
wire v_21969;
wire v_21970;
wire v_21971;
wire v_21972;
wire v_21973;
wire v_21974;
wire v_21975;
wire v_21976;
wire v_21977;
wire v_21978;
wire v_21979;
wire v_21980;
wire v_21981;
wire v_21982;
wire v_21983;
wire v_21984;
wire v_21985;
wire v_21986;
wire v_21987;
wire v_21988;
wire v_21989;
wire v_21990;
wire v_21991;
wire v_21992;
wire v_21993;
wire v_21994;
wire v_21995;
wire v_21996;
wire v_21997;
wire v_21998;
wire v_21999;
wire v_22000;
wire v_22001;
wire v_22002;
wire v_22003;
wire v_22004;
wire v_22005;
wire v_22006;
wire v_22007;
wire v_22008;
wire v_22009;
wire v_22010;
wire v_22011;
wire v_22012;
wire v_22013;
wire v_22014;
wire v_22015;
wire v_22016;
wire v_22017;
wire v_22018;
wire v_22019;
wire v_22020;
wire v_22021;
wire v_22022;
wire v_22023;
wire v_22024;
wire v_22025;
wire v_22026;
wire v_22027;
wire v_22028;
wire v_22029;
wire v_22030;
wire v_22031;
wire v_22032;
wire v_22033;
wire v_22034;
wire v_22035;
wire v_22036;
wire v_22037;
wire v_22038;
wire v_22039;
wire v_22040;
wire v_22041;
wire v_22042;
wire v_22043;
wire v_22044;
wire v_22045;
wire v_22046;
wire v_22047;
wire v_22048;
wire v_22049;
wire v_22050;
wire v_22051;
wire v_22052;
wire v_22053;
wire v_22054;
wire v_22055;
wire v_22056;
wire v_22057;
wire v_22058;
wire v_22059;
wire v_22060;
wire v_22061;
wire v_22062;
wire v_22063;
wire v_22064;
wire v_22065;
wire v_22066;
wire v_22067;
wire v_22068;
wire v_22069;
wire v_22070;
wire v_22071;
wire v_22072;
wire v_22073;
wire v_22074;
wire v_22075;
wire v_22076;
wire v_22077;
wire v_22078;
wire v_22079;
wire v_22080;
wire v_22081;
wire v_22082;
wire v_22083;
wire v_22084;
wire v_22085;
wire v_22086;
wire v_22087;
wire v_22088;
wire v_22089;
wire v_22090;
wire v_22091;
wire v_22092;
wire v_22093;
wire v_22094;
wire v_22095;
wire v_22096;
wire v_22097;
wire v_22098;
wire v_22099;
wire v_22100;
wire v_22101;
wire v_22102;
wire v_22103;
wire v_22104;
wire v_22105;
wire v_22106;
wire v_22107;
wire v_22108;
wire v_22109;
wire v_22110;
wire v_22111;
wire v_22112;
wire v_22113;
wire v_22114;
wire v_22115;
wire v_22116;
wire v_22117;
wire v_22118;
wire v_22119;
wire v_22120;
wire v_22121;
wire v_22122;
wire v_22123;
wire v_22124;
wire v_22125;
wire v_22126;
wire v_22127;
wire v_22128;
wire v_22129;
wire v_22130;
wire v_22131;
wire v_22132;
wire v_22133;
wire v_22134;
wire v_22135;
wire v_22136;
wire v_22137;
wire v_22138;
wire v_22139;
wire v_22140;
wire v_22141;
wire v_22142;
wire v_22143;
wire v_22144;
wire v_22145;
wire v_22146;
wire v_22147;
wire v_22148;
wire v_22149;
wire v_22150;
wire v_22151;
wire v_22152;
wire v_22153;
wire v_22154;
wire v_22155;
wire v_22156;
wire v_22157;
wire v_22158;
wire v_22159;
wire v_22160;
wire v_22161;
wire v_22162;
wire v_22163;
wire v_22164;
wire v_22165;
wire v_22166;
wire v_22167;
wire v_22168;
wire v_22169;
wire v_22170;
wire v_22171;
wire v_22172;
wire v_22173;
wire v_22174;
wire v_22175;
wire v_22176;
wire v_22177;
wire v_22178;
wire v_22179;
wire v_22180;
wire v_22181;
wire v_22182;
wire v_22183;
wire v_22184;
wire v_22185;
wire v_22186;
wire v_22187;
wire v_22188;
wire v_22189;
wire v_22190;
wire v_22191;
wire v_22192;
wire v_22193;
wire v_22194;
wire v_22195;
wire v_22196;
wire v_22197;
wire v_22198;
wire v_22199;
wire v_22200;
wire v_22201;
wire v_22202;
wire v_22203;
wire v_22204;
wire v_22205;
wire v_22206;
wire v_22207;
wire v_22208;
wire v_22209;
wire v_22210;
wire v_22211;
wire v_22212;
wire v_22213;
wire v_22214;
wire v_22215;
wire v_22216;
wire v_22217;
wire v_22218;
wire v_22219;
wire v_22220;
wire v_22221;
wire v_22222;
wire v_22223;
wire v_22224;
wire v_22225;
wire v_22226;
wire v_22227;
wire v_22228;
wire v_22229;
wire v_22230;
wire v_22231;
wire v_22232;
wire v_22233;
wire v_22234;
wire v_22235;
wire v_22236;
wire v_22237;
wire v_22238;
wire v_22239;
wire v_22240;
wire v_22241;
wire v_22242;
wire v_22243;
wire v_22244;
wire v_22245;
wire v_22246;
wire v_22247;
wire v_22248;
wire v_22249;
wire v_22250;
wire v_22251;
wire v_22252;
wire v_22253;
wire v_22254;
wire v_22255;
wire v_22256;
wire v_22257;
wire v_22258;
wire v_22259;
wire v_22260;
wire v_22261;
wire v_22262;
wire v_22263;
wire v_22264;
wire v_22265;
wire v_22266;
wire v_22267;
wire v_22268;
wire v_22269;
wire v_22270;
wire v_22271;
wire v_22272;
wire v_22273;
wire v_22274;
wire v_22275;
wire v_22276;
wire v_22277;
wire v_22278;
wire v_22279;
wire v_22280;
wire v_22281;
wire v_22282;
wire v_22283;
wire v_22284;
wire v_22285;
wire v_22286;
wire v_22287;
wire v_22288;
wire v_22289;
wire v_22290;
wire v_22291;
wire v_22292;
wire v_22293;
wire v_22294;
wire v_22295;
wire v_22296;
wire v_22297;
wire v_22298;
wire v_22299;
wire v_22300;
wire v_22301;
wire v_22302;
wire v_22303;
wire v_22304;
wire v_22305;
wire v_22306;
wire v_22307;
wire v_22308;
wire v_22309;
wire v_22310;
wire v_22311;
wire v_22312;
wire v_22313;
wire v_22314;
wire v_22315;
wire v_22316;
wire v_22317;
wire v_22318;
wire v_22319;
wire v_22320;
wire v_22321;
wire v_22322;
wire v_22323;
wire v_22324;
wire v_22325;
wire v_22326;
wire v_22327;
wire v_22328;
wire v_22329;
wire v_22330;
wire v_22331;
wire v_22332;
wire v_22333;
wire v_22334;
wire v_22335;
wire v_22336;
wire v_22337;
wire v_22338;
wire v_22339;
wire v_22340;
wire v_22341;
wire v_22342;
wire v_22343;
wire v_22344;
wire v_22345;
wire v_22346;
wire v_22347;
wire v_22348;
wire v_22349;
wire v_22350;
wire v_22351;
wire v_22352;
wire v_22353;
wire v_22354;
wire v_22355;
wire v_22356;
wire v_22357;
wire v_22358;
wire v_22359;
wire v_22360;
wire v_22361;
wire v_22362;
wire v_22363;
wire v_22364;
wire v_22365;
wire v_22366;
wire v_22367;
wire v_22368;
wire v_22369;
wire v_22370;
wire v_22371;
wire v_22372;
wire v_22373;
wire v_22374;
wire v_22375;
wire v_22376;
wire v_22377;
wire v_22378;
wire v_22379;
wire v_22380;
wire v_22381;
wire v_22382;
wire v_22383;
wire v_22384;
wire v_22385;
wire v_22386;
wire v_22387;
wire v_22388;
wire v_22389;
wire v_22390;
wire v_22391;
wire v_22392;
wire v_22393;
wire v_22394;
wire v_22395;
wire v_22396;
wire v_22397;
wire v_22398;
wire v_22399;
wire v_22400;
wire v_22401;
wire v_22402;
wire v_22403;
wire v_22404;
wire v_22405;
wire v_22406;
wire v_22407;
wire v_22408;
wire v_22409;
wire v_22410;
wire v_22411;
wire v_22412;
wire v_22413;
wire v_22414;
wire v_22415;
wire v_22416;
wire v_22417;
wire v_22418;
wire v_22419;
wire v_22420;
wire v_22421;
wire v_22422;
wire v_22423;
wire v_22424;
wire v_22425;
wire v_22426;
wire v_22427;
wire v_22428;
wire v_22429;
wire v_22430;
wire v_22431;
wire v_22432;
wire v_22433;
wire v_22434;
wire v_22435;
wire v_22436;
wire v_22437;
wire v_22438;
wire v_22439;
wire v_22440;
wire v_22441;
wire v_22442;
wire v_22443;
wire v_22444;
wire v_22445;
wire v_22446;
wire v_22447;
wire v_22448;
wire v_22449;
wire v_22450;
wire v_22451;
wire v_22452;
wire v_22453;
wire v_22454;
wire v_22455;
wire v_22456;
wire v_22457;
wire v_22458;
wire v_22459;
wire v_22460;
wire v_22461;
wire v_22462;
wire v_22463;
wire v_22464;
wire v_22465;
wire v_22466;
wire v_22467;
wire v_22468;
wire v_22469;
wire v_22470;
wire v_22471;
wire v_22472;
wire v_22473;
wire v_22474;
wire v_22475;
wire v_22476;
wire v_22477;
wire v_22478;
wire v_22479;
wire v_22480;
wire v_22481;
wire v_22482;
wire v_22483;
wire v_22484;
wire v_22485;
wire v_22486;
wire v_22487;
wire v_22488;
wire v_22489;
wire v_22490;
wire v_22491;
wire v_22492;
wire v_22493;
wire v_22494;
wire v_22495;
wire v_22496;
wire v_22497;
wire v_22498;
wire v_22499;
wire v_22500;
wire v_22501;
wire v_22502;
wire v_22503;
wire v_22504;
wire v_22505;
wire v_22506;
wire v_22507;
wire v_22508;
wire v_22509;
wire v_22510;
wire v_22511;
wire v_22512;
wire v_22513;
wire v_22514;
wire v_22515;
wire v_22516;
wire v_22517;
wire v_22518;
wire v_22519;
wire v_22520;
wire v_22521;
wire v_22522;
wire v_22523;
wire v_22524;
wire v_22525;
wire v_22526;
wire v_22527;
wire v_22528;
wire v_22529;
wire v_22530;
wire v_22531;
wire v_22532;
wire v_22533;
wire v_22534;
wire v_22535;
wire v_22536;
wire v_22537;
wire v_22538;
wire v_22539;
wire v_22540;
wire v_22541;
wire v_22542;
wire v_22543;
wire v_22544;
wire v_22545;
wire v_22546;
wire v_22547;
wire v_22548;
wire v_22549;
wire v_22550;
wire v_22551;
wire v_22552;
wire v_22553;
wire v_22554;
wire v_22555;
wire v_22556;
wire v_22557;
wire v_22558;
wire v_22559;
wire v_22560;
wire v_22561;
wire v_22562;
wire v_22563;
wire v_22564;
wire v_22565;
wire v_22566;
wire v_22567;
wire v_22568;
wire v_22569;
wire v_22570;
wire v_22571;
wire v_22572;
wire v_22573;
wire v_22574;
wire v_22575;
wire v_22576;
wire v_22577;
wire v_22578;
wire v_22579;
wire v_22580;
wire v_22581;
wire v_22582;
wire v_22583;
wire v_22584;
wire v_22585;
wire v_22586;
wire v_22587;
wire v_22588;
wire v_22589;
wire v_22590;
wire v_22591;
wire v_22592;
wire v_22593;
wire v_22594;
wire v_22595;
wire v_22596;
wire v_22597;
wire v_22598;
wire v_22599;
wire v_22600;
wire v_22601;
wire v_22602;
wire v_22603;
wire v_22604;
wire v_22605;
wire v_22606;
wire v_22607;
wire v_22608;
wire v_22609;
wire v_22610;
wire v_22611;
wire v_22612;
wire v_22613;
wire v_22614;
wire v_22615;
wire v_22616;
wire v_22617;
wire v_22618;
wire v_22619;
wire v_22620;
wire v_22621;
wire v_22622;
wire v_22623;
wire v_22624;
wire v_22625;
wire v_22626;
wire v_22627;
wire v_22628;
wire v_22629;
wire v_22630;
wire v_22631;
wire v_22632;
wire v_22633;
wire v_22634;
wire v_22635;
wire v_22636;
wire v_22637;
wire v_22638;
wire v_22639;
wire v_22640;
wire v_22641;
wire v_22642;
wire v_22643;
wire v_22644;
wire v_22645;
wire v_22646;
wire v_22647;
wire v_22648;
wire v_22649;
wire v_22650;
wire v_22651;
wire v_22652;
wire v_22653;
wire v_22654;
wire v_22655;
wire v_22656;
wire v_22657;
wire v_22658;
wire v_22659;
wire v_22660;
wire v_22661;
wire v_22662;
wire v_22663;
wire v_22664;
wire v_22665;
wire v_22666;
wire v_22667;
wire v_22668;
wire v_22669;
wire v_22670;
wire v_22671;
wire v_22672;
wire v_22673;
wire v_22674;
wire v_22675;
wire v_22676;
wire v_22677;
wire v_22678;
wire v_22679;
wire v_22680;
wire v_22681;
wire v_22682;
wire v_22683;
wire v_22684;
wire v_22685;
wire v_22686;
wire v_22687;
wire v_22688;
wire v_22689;
wire v_22690;
wire v_22691;
wire v_22692;
wire v_22693;
wire v_22694;
wire v_22695;
wire v_22696;
wire v_22697;
wire v_22698;
wire v_22699;
wire v_22700;
wire v_22701;
wire v_22702;
wire v_22703;
wire v_22704;
wire v_22705;
wire v_22706;
wire v_22707;
wire v_22708;
wire v_22709;
wire v_22710;
wire v_22711;
wire v_22712;
wire v_22713;
wire v_22714;
wire v_22715;
wire v_22716;
wire v_22717;
wire v_22718;
wire v_22719;
wire v_22720;
wire v_22721;
wire v_22722;
wire v_22723;
wire v_22724;
wire v_22725;
wire v_22726;
wire v_22727;
wire v_22728;
wire v_22729;
wire v_22730;
wire v_22731;
wire v_22732;
wire v_22733;
wire v_22734;
wire v_22735;
wire v_22736;
wire v_22737;
wire v_22738;
wire v_22739;
wire v_22740;
wire v_22741;
wire v_22742;
wire v_22743;
wire v_22744;
wire v_22745;
wire v_22746;
wire v_22747;
wire v_22748;
wire v_22749;
wire v_22750;
wire v_22751;
wire v_22752;
wire v_22753;
wire v_22754;
wire v_22755;
wire v_22756;
wire v_22757;
wire v_22758;
wire v_22759;
wire v_22760;
wire v_22761;
wire v_22762;
wire v_22763;
wire v_22764;
wire v_22765;
wire v_22766;
wire v_22767;
wire v_22768;
wire v_22769;
wire v_22770;
wire v_22771;
wire v_22772;
wire v_22773;
wire v_22774;
wire v_22775;
wire v_22776;
wire v_22777;
wire v_22778;
wire v_22779;
wire v_22780;
wire v_22781;
wire v_22782;
wire v_22783;
wire v_22784;
wire v_22785;
wire v_22786;
wire v_22787;
wire v_22788;
wire v_22789;
wire v_22790;
wire v_22791;
wire v_22792;
wire v_22793;
wire v_22794;
wire v_22795;
wire v_22796;
wire v_22797;
wire v_22798;
wire v_22799;
wire v_22800;
wire v_22801;
wire v_22802;
wire v_22803;
wire v_22804;
wire v_22805;
wire v_22806;
wire v_22807;
wire v_22808;
wire v_22809;
wire v_22810;
wire v_22811;
wire v_22812;
wire v_22813;
wire v_22814;
wire v_22815;
wire v_22816;
wire v_22817;
wire v_22818;
wire v_22819;
wire v_22820;
wire v_22821;
wire v_22822;
wire v_22823;
wire v_22824;
wire v_22825;
wire v_22826;
wire v_22827;
wire v_22828;
wire v_22829;
wire v_22830;
wire v_22831;
wire v_22832;
wire v_22833;
wire v_22834;
wire v_22835;
wire v_22836;
wire v_22837;
wire v_22838;
wire v_22839;
wire v_22840;
wire v_22841;
wire v_22842;
wire v_22843;
wire v_22844;
wire v_22845;
wire v_22846;
wire v_22847;
wire v_22848;
wire v_22849;
wire v_22850;
wire v_22851;
wire v_22852;
wire v_22853;
wire v_22854;
wire v_22855;
wire v_22856;
wire v_22857;
wire v_22858;
wire v_22859;
wire v_22860;
wire v_22861;
wire v_22862;
wire v_22863;
wire v_22864;
wire v_22865;
wire v_22866;
wire v_22867;
wire v_22868;
wire v_22869;
wire v_22870;
wire v_22871;
wire v_22872;
wire v_22873;
wire v_22874;
wire v_22875;
wire v_22876;
wire v_22877;
wire v_22878;
wire v_22879;
wire v_22880;
wire v_22881;
wire v_22882;
wire v_22883;
wire v_22884;
wire v_22885;
wire v_22886;
wire v_22887;
wire v_22888;
wire v_22889;
wire v_22890;
wire v_22891;
wire v_22892;
wire v_22893;
wire v_22894;
wire v_22895;
wire v_22896;
wire v_22897;
wire v_22898;
wire v_22899;
wire v_22900;
wire v_22901;
wire v_22902;
wire v_22903;
wire v_22904;
wire v_22905;
wire v_22906;
wire v_22907;
wire v_22908;
wire v_22909;
wire v_22910;
wire v_22911;
wire v_22912;
wire v_22913;
wire v_22914;
wire v_22915;
wire v_22916;
wire v_22917;
wire v_22918;
wire v_22919;
wire v_22920;
wire v_22921;
wire v_22922;
wire v_22923;
wire v_22924;
wire v_22925;
wire v_22926;
wire v_22927;
wire v_22928;
wire v_22929;
wire v_22930;
wire v_22931;
wire v_22932;
wire v_22933;
wire v_22934;
wire v_22935;
wire v_22936;
wire v_22937;
wire v_22938;
wire v_22939;
wire v_22940;
wire v_22941;
wire v_22942;
wire v_22943;
wire v_22944;
wire v_22945;
wire v_22946;
wire v_22947;
wire v_22948;
wire v_22949;
wire v_22950;
wire v_22951;
wire v_22952;
wire v_22953;
wire v_22954;
wire v_22955;
wire v_22956;
wire v_22957;
wire v_22958;
wire v_22959;
wire v_22960;
wire v_22961;
wire v_22962;
wire v_22963;
wire v_22964;
wire v_22965;
wire v_22966;
wire v_22967;
wire v_22968;
wire v_22969;
wire v_22970;
wire v_22971;
wire v_22972;
wire v_22973;
wire v_22974;
wire v_22975;
wire v_22976;
wire v_22977;
wire v_22978;
wire v_22979;
wire v_22980;
wire v_22981;
wire v_22982;
wire v_22983;
wire v_22984;
wire v_22985;
wire v_22986;
wire v_22987;
wire v_22988;
wire v_22989;
wire v_22990;
wire v_22991;
wire v_22992;
wire v_22993;
wire v_22994;
wire v_22995;
wire v_22996;
wire v_22997;
wire v_22998;
wire v_22999;
wire v_23000;
wire v_23001;
wire v_23002;
wire v_23003;
wire v_23004;
wire v_23005;
wire v_23006;
wire v_23007;
wire v_23008;
wire v_23009;
wire v_23010;
wire v_23011;
wire v_23012;
wire v_23013;
wire v_23014;
wire v_23015;
wire v_23016;
wire v_23017;
wire v_23018;
wire v_23019;
wire v_23020;
wire v_23021;
wire v_23022;
wire v_23023;
wire v_23024;
wire v_23025;
wire v_23026;
wire v_23027;
wire v_23028;
wire v_23029;
wire v_23030;
wire v_23031;
wire v_23032;
wire v_23033;
wire v_23034;
wire v_23035;
wire v_23036;
wire v_23037;
wire v_23038;
wire v_23039;
wire v_23040;
wire v_23041;
wire v_23042;
wire v_23043;
wire v_23044;
wire v_23045;
wire v_23046;
wire v_23047;
wire v_23048;
wire v_23049;
wire v_23050;
wire v_23051;
wire v_23052;
wire v_23053;
wire v_23054;
wire v_23055;
wire v_23056;
wire v_23057;
wire v_23058;
wire v_23059;
wire v_23060;
wire v_23061;
wire v_23062;
wire v_23063;
wire v_23064;
wire v_23065;
wire v_23066;
wire v_23067;
wire v_23068;
wire v_23069;
wire v_23070;
wire v_23071;
wire v_23072;
wire v_23073;
wire v_23074;
wire v_23075;
wire v_23076;
wire v_23077;
wire v_23078;
wire v_23079;
wire v_23080;
wire v_23081;
wire v_23082;
wire v_23083;
wire v_23084;
wire v_23085;
wire v_23086;
wire v_23087;
wire v_23088;
wire v_23089;
wire v_23090;
wire v_23091;
wire v_23092;
wire v_23093;
wire v_23094;
wire v_23095;
wire v_23096;
wire v_23097;
wire v_23098;
wire v_23099;
wire v_23100;
wire v_23101;
wire v_23102;
wire v_23103;
wire v_23104;
wire v_23105;
wire v_23106;
wire v_23107;
wire v_23108;
wire v_23109;
wire v_23110;
wire v_23111;
wire v_23112;
wire v_23113;
wire v_23114;
wire v_23115;
wire v_23116;
wire v_23117;
wire v_23118;
wire v_23119;
wire v_23120;
wire v_23121;
wire v_23122;
wire v_23123;
wire v_23124;
wire v_23125;
wire v_23126;
wire v_23127;
wire v_23128;
wire v_23129;
wire v_23130;
wire v_23131;
wire v_23132;
wire v_23133;
wire v_23134;
wire v_23135;
wire v_23136;
wire v_23137;
wire v_23138;
wire v_23139;
wire v_23140;
wire v_23141;
wire v_23142;
wire v_23143;
wire v_23144;
wire v_23145;
wire v_23146;
wire v_23147;
wire v_23148;
wire v_23149;
wire v_23150;
wire v_23151;
wire v_23152;
wire v_23153;
wire v_23154;
wire v_23155;
wire v_23156;
wire v_23157;
wire v_23158;
wire v_23159;
wire v_23160;
wire v_23161;
wire v_23162;
wire v_23163;
wire v_23164;
wire v_23165;
wire v_23166;
wire v_23167;
wire v_23168;
wire v_23169;
wire v_23170;
wire v_23171;
wire v_23172;
wire v_23173;
wire v_23174;
wire v_23175;
wire v_23176;
wire v_23177;
wire v_23178;
wire v_23179;
wire v_23180;
wire v_23181;
wire v_23182;
wire v_23183;
wire v_23184;
wire v_23185;
wire v_23186;
wire v_23187;
wire v_23188;
wire v_23189;
wire v_23190;
wire v_23191;
wire v_23192;
wire v_23193;
wire v_23194;
wire v_23195;
wire v_23196;
wire v_23197;
wire v_23198;
wire v_23199;
wire v_23200;
wire v_23201;
wire v_23202;
wire v_23203;
wire v_23204;
wire v_23205;
wire v_23206;
wire v_23207;
wire v_23208;
wire v_23209;
wire v_23210;
wire v_23211;
wire v_23212;
wire v_23213;
wire v_23214;
wire v_23215;
wire v_23216;
wire v_23217;
wire v_23218;
wire v_23219;
wire v_23220;
wire v_23221;
wire v_23222;
wire v_23223;
wire v_23224;
wire v_23225;
wire v_23226;
wire v_23227;
wire v_23228;
wire v_23229;
wire v_23230;
wire v_23231;
wire v_23232;
wire v_23233;
wire v_23234;
wire v_23235;
wire v_23236;
wire v_23237;
wire v_23238;
wire v_23239;
wire v_23240;
wire v_23241;
wire v_23242;
wire v_23243;
wire v_23244;
wire v_23245;
wire v_23246;
wire v_23247;
wire v_23248;
wire v_23249;
wire v_23250;
wire v_23251;
wire v_23252;
wire v_23253;
wire v_23254;
wire v_23255;
wire v_23256;
wire v_23257;
wire v_23258;
wire v_23259;
wire v_23260;
wire v_23261;
wire v_23262;
wire v_23263;
wire v_23264;
wire v_23265;
wire v_23266;
wire v_23267;
wire v_23268;
wire v_23269;
wire v_23270;
wire v_23271;
wire v_23272;
wire v_23273;
wire v_23274;
wire v_23275;
wire v_23276;
wire v_23277;
wire v_23278;
wire v_23279;
wire v_23280;
wire v_23281;
wire v_23282;
wire v_23283;
wire v_23284;
wire v_23285;
wire v_23286;
wire v_23287;
wire v_23288;
wire v_23289;
wire v_23290;
wire v_23291;
wire v_23292;
wire v_23293;
wire v_23294;
wire v_23295;
wire v_23296;
wire v_23297;
wire v_23298;
wire v_23299;
wire v_23300;
wire v_23301;
wire v_23302;
wire v_23303;
wire v_23304;
wire v_23305;
wire v_23306;
wire v_23307;
wire v_23308;
wire v_23309;
wire v_23310;
wire v_23311;
wire v_23312;
wire v_23313;
wire v_23314;
wire v_23315;
wire v_23316;
wire v_23317;
wire v_23318;
wire v_23319;
wire v_23320;
wire v_23321;
wire v_23322;
wire v_23323;
wire v_23324;
wire v_23325;
wire v_23326;
wire v_23327;
wire v_23328;
wire v_23329;
wire v_23330;
wire v_23331;
wire v_23332;
wire v_23333;
wire v_23334;
wire v_23335;
wire v_23336;
wire v_23337;
wire v_23338;
wire v_23339;
wire v_23340;
wire v_23341;
wire v_23342;
wire v_23343;
wire v_23344;
wire v_23345;
wire v_23346;
wire v_23347;
wire v_23348;
wire v_23349;
wire v_23350;
wire v_23351;
wire v_23352;
wire v_23353;
wire v_23354;
wire v_23355;
wire v_23356;
wire v_23357;
wire v_23358;
wire v_23359;
wire v_23360;
wire v_23361;
wire v_23362;
wire v_23363;
wire v_23364;
wire v_23365;
wire v_23366;
wire v_23367;
wire v_23368;
wire v_23369;
wire v_23370;
wire v_23371;
wire v_23372;
wire v_23373;
wire v_23374;
wire v_23375;
wire v_23376;
wire v_23377;
wire v_23378;
wire v_23379;
wire v_23380;
wire v_23381;
wire v_23382;
wire v_23383;
wire v_23384;
wire v_23385;
wire v_23386;
wire v_23387;
wire v_23388;
wire v_23389;
wire v_23390;
wire v_23391;
wire v_23392;
wire v_23393;
wire v_23394;
wire v_23395;
wire v_23396;
wire v_23397;
wire v_23398;
wire v_23399;
wire v_23400;
wire v_23401;
wire v_23402;
wire v_23403;
wire v_23404;
wire v_23405;
wire v_23406;
wire v_23407;
wire v_23408;
wire v_23409;
wire v_23410;
wire v_23411;
wire v_23412;
wire v_23413;
wire v_23414;
wire v_23415;
wire v_23416;
wire v_23417;
wire v_23418;
wire v_23419;
wire v_23420;
wire v_23421;
wire v_23422;
wire v_23423;
wire v_23424;
wire v_23425;
wire v_23426;
wire v_23427;
wire v_23428;
wire v_23429;
wire v_23430;
wire v_23431;
wire v_23432;
wire v_23433;
wire v_23434;
wire v_23435;
wire v_23436;
wire v_23437;
wire v_23438;
wire v_23439;
wire v_23440;
wire v_23441;
wire v_23442;
wire v_23443;
wire v_23444;
wire v_23445;
wire v_23446;
wire v_23447;
wire v_23448;
wire v_23449;
wire v_23450;
wire v_23451;
wire v_23452;
wire v_23453;
wire v_23454;
wire v_23455;
wire v_23456;
wire v_23457;
wire v_23458;
wire v_23459;
wire v_23460;
wire v_23461;
wire v_23462;
wire v_23463;
wire v_23464;
wire v_23465;
wire v_23466;
wire v_23467;
wire v_23468;
wire v_23469;
wire v_23470;
wire v_23471;
wire v_23472;
wire v_23473;
wire v_23474;
wire v_23475;
wire v_23476;
wire v_23477;
wire v_23478;
wire v_23479;
wire v_23480;
wire v_23481;
wire v_23482;
wire v_23483;
wire v_23484;
wire v_23485;
wire v_23486;
wire v_23487;
wire v_23488;
wire v_23489;
wire v_23490;
wire v_23491;
wire v_23492;
wire v_23493;
wire v_23494;
wire v_23495;
wire v_23496;
wire v_23497;
wire v_23498;
wire v_23499;
wire v_23500;
wire v_23501;
wire v_23502;
wire v_23503;
wire v_23504;
wire v_23505;
wire v_23506;
wire v_23507;
wire v_23508;
wire v_23509;
wire v_23510;
wire v_23511;
wire v_23512;
wire v_23513;
wire v_23514;
wire v_23515;
wire v_23516;
wire v_23517;
wire v_23518;
wire v_23519;
wire v_23520;
wire v_23521;
wire v_23522;
wire v_23523;
wire v_23524;
wire v_23525;
wire v_23526;
wire v_23527;
wire v_23528;
wire v_23529;
wire v_23530;
wire v_23531;
wire v_23532;
wire v_23533;
wire v_23534;
wire v_23535;
wire v_23536;
wire v_23537;
wire v_23538;
wire v_23539;
wire v_23540;
wire v_23541;
wire v_23542;
wire v_23543;
wire v_23544;
wire v_23545;
wire v_23546;
wire v_23547;
wire v_23548;
wire v_23549;
wire v_23550;
wire v_23551;
wire v_23552;
wire v_23553;
wire v_23554;
wire v_23555;
wire v_23556;
wire v_23557;
wire v_23558;
wire v_23559;
wire v_23560;
wire v_23561;
wire v_23562;
wire v_23563;
wire v_23564;
wire v_23565;
wire v_23566;
wire v_23567;
wire v_23568;
wire v_23569;
wire v_23570;
wire v_23571;
wire v_23572;
wire v_23573;
wire v_23574;
wire v_23575;
wire v_23576;
wire v_23577;
wire v_23578;
wire v_23579;
wire v_23580;
wire v_23581;
wire v_23582;
wire v_23583;
wire v_23584;
wire v_23585;
wire v_23586;
wire v_23587;
wire v_23588;
wire v_23589;
wire v_23590;
wire v_23591;
wire v_23592;
wire v_23593;
wire v_23594;
wire v_23595;
wire v_23596;
wire v_23597;
wire v_23598;
wire v_23599;
wire v_23600;
wire v_23601;
wire v_23602;
wire v_23603;
wire v_23604;
wire v_23605;
wire v_23606;
wire v_23607;
wire v_23608;
wire v_23609;
wire v_23610;
wire v_23611;
wire v_23612;
wire v_23613;
wire v_23614;
wire v_23615;
wire v_23616;
wire v_23617;
wire v_23618;
wire v_23619;
wire v_23620;
wire v_23621;
wire v_23622;
wire v_23623;
wire v_23624;
wire v_23625;
wire v_23626;
wire v_23627;
wire v_23628;
wire v_23629;
wire v_23630;
wire v_23631;
wire v_23632;
wire v_23633;
wire v_23634;
wire v_23635;
wire v_23636;
wire v_23637;
wire v_23638;
wire v_23639;
wire v_23640;
wire v_23641;
wire v_23642;
wire v_23643;
wire v_23644;
wire v_23645;
wire v_23646;
wire v_23647;
wire v_23648;
wire v_23649;
wire v_23650;
wire v_23651;
wire v_23652;
wire v_23653;
wire v_23654;
wire v_23655;
wire v_23656;
wire v_23657;
wire v_23658;
wire v_23659;
wire v_23660;
wire v_23661;
wire v_23662;
wire v_23663;
wire v_23664;
wire v_23665;
wire v_23666;
wire v_23667;
wire v_23668;
wire v_23669;
wire v_23670;
wire v_23671;
wire v_23672;
wire v_23673;
wire v_23674;
wire v_23675;
wire v_23676;
wire v_23677;
wire v_23678;
wire v_23679;
wire v_23680;
wire v_23681;
wire v_23682;
wire v_23683;
wire v_23684;
wire v_23685;
wire v_23686;
wire v_23687;
wire v_23688;
wire v_23689;
wire v_23690;
wire v_23691;
wire v_23692;
wire v_23693;
wire v_23694;
wire v_23695;
wire v_23696;
wire v_23697;
wire v_23698;
wire v_23699;
wire v_23700;
wire v_23701;
wire v_23702;
wire v_23703;
wire v_23704;
wire v_23705;
wire v_23706;
wire v_23707;
wire v_23708;
wire v_23709;
wire v_23710;
wire v_23711;
wire v_23712;
wire v_23713;
wire v_23714;
wire v_23715;
wire v_23716;
wire v_23717;
wire v_23718;
wire v_23719;
wire v_23720;
wire v_23721;
wire v_23722;
wire v_23723;
wire v_23724;
wire v_23725;
wire v_23726;
wire v_23727;
wire v_23728;
wire v_23729;
wire v_23730;
wire v_23731;
wire v_23732;
wire v_23733;
wire v_23734;
wire v_23735;
wire v_23736;
wire v_23737;
wire v_23738;
wire v_23739;
wire v_23740;
wire v_23741;
wire v_23742;
wire v_23743;
wire v_23744;
wire v_23745;
wire v_23746;
wire v_23747;
wire v_23748;
wire v_23749;
wire v_23750;
wire v_23751;
wire v_23752;
wire v_23753;
wire v_23754;
wire v_23755;
wire v_23756;
wire v_23757;
wire v_23758;
wire v_23759;
wire v_23760;
wire v_23761;
wire v_23762;
wire v_23763;
wire v_23764;
wire v_23765;
wire v_23766;
wire v_23767;
wire v_23768;
wire v_23769;
wire v_23770;
wire v_23771;
wire v_23772;
wire v_23773;
wire v_23774;
wire v_23775;
wire v_23776;
wire v_23777;
wire v_23778;
wire v_23779;
wire v_23780;
wire v_23781;
wire v_23782;
wire v_23783;
wire v_23784;
wire v_23785;
wire v_23786;
wire v_23787;
wire v_23788;
wire v_23789;
wire v_23790;
wire v_23791;
wire v_23792;
wire v_23793;
wire v_23794;
wire v_23795;
wire v_23796;
wire v_23797;
wire v_23798;
wire v_23799;
wire v_23800;
wire v_23801;
wire v_23802;
wire v_23803;
wire v_23804;
wire v_23805;
wire v_23806;
wire v_23807;
wire v_23808;
wire v_23809;
wire v_23810;
wire v_23811;
wire v_23812;
wire v_23813;
wire v_23814;
wire v_23815;
wire v_23816;
wire v_23817;
wire v_23818;
wire v_23819;
wire v_23820;
wire v_23821;
wire v_23822;
wire v_23823;
wire v_23824;
wire v_23825;
wire v_23826;
wire v_23827;
wire v_23828;
wire v_23829;
wire v_23830;
wire v_23831;
wire v_23832;
wire v_23833;
wire v_23834;
wire v_23835;
wire v_23836;
wire v_23837;
wire v_23838;
wire v_23839;
wire v_23840;
wire v_23841;
wire v_23842;
wire v_23843;
wire v_23844;
wire v_23845;
wire v_23846;
wire v_23847;
wire v_23848;
wire v_23849;
wire v_23850;
wire v_23851;
wire v_23852;
wire v_23853;
wire v_23854;
wire v_23855;
wire v_23856;
wire v_23857;
wire v_23858;
wire v_23859;
wire v_23860;
wire v_23861;
wire v_23862;
wire v_23863;
wire v_23864;
wire v_23865;
wire v_23866;
wire v_23867;
wire v_23868;
wire v_23869;
wire v_23870;
wire v_23871;
wire v_23872;
wire v_23873;
wire v_23874;
wire v_23875;
wire v_23876;
wire v_23877;
wire v_23878;
wire v_23879;
wire v_23880;
wire v_23881;
wire v_23882;
wire v_23883;
wire v_23884;
wire v_23885;
wire v_23886;
wire v_23887;
wire v_23888;
wire v_23889;
wire v_23890;
wire v_23891;
wire v_23892;
wire v_23893;
wire v_23894;
wire v_23895;
wire v_23896;
wire v_23897;
wire v_23898;
wire v_23899;
wire v_23900;
wire v_23901;
wire v_23902;
wire v_23903;
wire v_23904;
wire v_23905;
wire v_23906;
wire v_23907;
wire v_23908;
wire v_23909;
wire v_23910;
wire v_23911;
wire v_23912;
wire v_23913;
wire v_23914;
wire v_23915;
wire v_23916;
wire v_23917;
wire v_23918;
wire v_23919;
wire v_23920;
wire v_23921;
wire v_23922;
wire v_23923;
wire v_23924;
wire v_23925;
wire v_23926;
wire v_23927;
wire v_23928;
wire v_23929;
wire v_23930;
wire v_23931;
wire v_23932;
wire v_23933;
wire v_23934;
wire v_23935;
wire v_23936;
wire v_23937;
wire v_23938;
wire v_23939;
wire v_23940;
wire v_23941;
wire v_23942;
wire v_23943;
wire v_23944;
wire v_23945;
wire v_23946;
wire v_23947;
wire v_23948;
wire v_23949;
wire v_23950;
wire v_23951;
wire v_23952;
wire v_23953;
wire v_23954;
wire v_23955;
wire v_23956;
wire v_23957;
wire v_23958;
wire v_23959;
wire v_23960;
wire v_23961;
wire v_23962;
wire v_23963;
wire v_23964;
wire v_23965;
wire v_23966;
wire v_23967;
wire v_23968;
wire v_23969;
wire v_23970;
wire v_23971;
wire v_23972;
wire v_23973;
wire v_23974;
wire v_23975;
wire v_23976;
wire v_23977;
wire v_23978;
wire v_23979;
wire v_23980;
wire v_23981;
wire v_23982;
wire v_23983;
wire v_23984;
wire v_23985;
wire v_23986;
wire v_23987;
wire v_23988;
wire v_23989;
wire v_23990;
wire v_23991;
wire v_23992;
wire v_23993;
wire v_23994;
wire v_23995;
wire v_23996;
wire v_23997;
wire v_23998;
wire v_23999;
wire v_24000;
wire v_24001;
wire v_24002;
wire v_24003;
wire v_24004;
wire v_24005;
wire v_24006;
wire v_24007;
wire v_24008;
wire v_24009;
wire v_24010;
wire v_24011;
wire v_24012;
wire v_24013;
wire v_24014;
wire v_24015;
wire v_24016;
wire v_24017;
wire v_24018;
wire v_24019;
wire v_24020;
wire v_24021;
wire v_24022;
wire v_24023;
wire v_24024;
wire v_24025;
wire v_24026;
wire v_24027;
wire v_24028;
wire v_24029;
wire v_24030;
wire v_24031;
wire v_24032;
wire v_24033;
wire v_24034;
wire v_24035;
wire v_24036;
wire v_24037;
wire v_24038;
wire v_24039;
wire v_24040;
wire v_24041;
wire v_24042;
wire v_24043;
wire v_24044;
wire v_24045;
wire v_24046;
wire v_24047;
wire v_24048;
wire v_24049;
wire v_24050;
wire v_24051;
wire v_24052;
wire v_24053;
wire v_24054;
wire v_24055;
wire v_24056;
wire v_24057;
wire v_24058;
wire v_24059;
wire v_24060;
wire v_24061;
wire v_24062;
wire v_24063;
wire v_24064;
wire v_24065;
wire v_24066;
wire v_24067;
wire v_24068;
wire v_24069;
wire v_24070;
wire v_24071;
wire v_24072;
wire v_24073;
wire v_24074;
wire v_24075;
wire v_24076;
wire v_24077;
wire v_24078;
wire v_24079;
wire v_24080;
wire v_24081;
wire v_24082;
wire v_24083;
wire v_24084;
wire v_24085;
wire v_24086;
wire v_24087;
wire v_24088;
wire v_24089;
wire v_24090;
wire v_24091;
wire v_24092;
wire v_24093;
wire v_24094;
wire v_24095;
wire v_24096;
wire v_24097;
wire v_24098;
wire v_24099;
wire v_24100;
wire v_24101;
wire v_24102;
wire v_24103;
wire v_24104;
wire v_24105;
wire v_24106;
wire v_24107;
wire v_24108;
wire v_24109;
wire v_24110;
wire v_24111;
wire v_24112;
wire v_24113;
wire v_24114;
wire v_24115;
wire v_24116;
wire v_24117;
wire v_24118;
wire v_24119;
wire v_24120;
wire v_24121;
wire v_24122;
wire v_24123;
wire v_24124;
wire v_24125;
wire v_24126;
wire v_24127;
wire v_24128;
wire v_24129;
wire v_24130;
wire v_24131;
wire v_24132;
wire v_24133;
wire v_24134;
wire v_24135;
wire v_24136;
wire v_24137;
wire v_24138;
wire v_24139;
wire v_24140;
wire v_24141;
wire v_24142;
wire v_24143;
wire v_24144;
wire v_24145;
wire v_24146;
wire v_24147;
wire v_24148;
wire v_24149;
wire v_24150;
wire v_24151;
wire v_24152;
wire v_24153;
wire v_24154;
wire v_24155;
wire v_24156;
wire v_24157;
wire v_24158;
wire v_24159;
wire v_24160;
wire v_24161;
wire v_24162;
wire v_24163;
wire v_24164;
wire v_24165;
wire v_24166;
wire v_24167;
wire v_24168;
wire v_24169;
wire v_24170;
wire v_24171;
wire v_24172;
wire v_24173;
wire v_24174;
wire v_24175;
wire v_24176;
wire v_24177;
wire v_24178;
wire v_24179;
wire v_24180;
wire v_24181;
wire v_24182;
wire v_24183;
wire v_24184;
wire v_24185;
wire v_24186;
wire v_24187;
wire v_24188;
wire v_24189;
wire v_24190;
wire v_24191;
wire v_24192;
wire v_24193;
wire v_24194;
wire v_24195;
wire v_24196;
wire v_24197;
wire v_24198;
wire v_24199;
wire v_24200;
wire v_24201;
wire v_24202;
wire v_24203;
wire v_24204;
wire v_24205;
wire v_24206;
wire v_24207;
wire v_24208;
wire v_24209;
wire v_24210;
wire v_24211;
wire v_24212;
wire v_24213;
wire v_24214;
wire v_24215;
wire v_24216;
wire v_24217;
wire v_24218;
wire v_24219;
wire v_24220;
wire v_24221;
wire v_24222;
wire v_24223;
wire v_24224;
wire v_24225;
wire v_24226;
wire v_24227;
wire v_24228;
wire v_24229;
wire v_24230;
wire v_24231;
wire v_24232;
wire v_24233;
wire v_24234;
wire v_24235;
wire v_24236;
wire v_24237;
wire v_24238;
wire v_24239;
wire v_24240;
wire v_24241;
wire v_24242;
wire v_24243;
wire v_24244;
wire v_24245;
wire v_24246;
wire v_24247;
wire v_24248;
wire v_24249;
wire v_24250;
wire v_24251;
wire v_24252;
wire v_24253;
wire v_24254;
wire v_24255;
wire v_24256;
wire v_24257;
wire v_24258;
wire v_24259;
wire v_24260;
wire v_24261;
wire v_24262;
wire v_24263;
wire v_24264;
wire v_24265;
wire v_24266;
wire v_24267;
wire v_24268;
wire v_24269;
wire v_24270;
wire v_24271;
wire v_24272;
wire v_24273;
wire v_24274;
wire v_24275;
wire v_24276;
wire v_24277;
wire v_24278;
wire v_24279;
wire v_24280;
wire v_24281;
wire v_24282;
wire v_24283;
wire v_24284;
wire v_24285;
wire v_24286;
wire v_24287;
wire v_24288;
wire v_24289;
wire v_24290;
wire v_24291;
wire v_24292;
wire v_24293;
wire v_24294;
wire v_24295;
wire v_24296;
wire v_24297;
wire v_24298;
wire v_24299;
wire v_24300;
wire v_24301;
wire v_24302;
wire v_24303;
wire v_24304;
wire v_24305;
wire v_24306;
wire v_24307;
wire v_24308;
wire v_24309;
wire v_24310;
wire v_24311;
wire v_24312;
wire v_24313;
wire v_24314;
wire v_24315;
wire v_24316;
wire v_24317;
wire v_24318;
wire v_24319;
wire v_24320;
wire v_24321;
wire v_24322;
wire v_24323;
wire v_24324;
wire v_24325;
wire v_24326;
wire v_24327;
wire v_24328;
wire v_24329;
wire v_24330;
wire v_24331;
wire v_24332;
wire v_24333;
wire v_24334;
wire v_24335;
wire v_24336;
wire v_24337;
wire v_24338;
wire v_24339;
wire v_24340;
wire v_24341;
wire v_24342;
wire v_24343;
wire v_24344;
wire v_24345;
wire v_24346;
wire v_24347;
wire v_24348;
wire v_24349;
wire v_24350;
wire v_24351;
wire v_24352;
wire v_24353;
wire v_24354;
wire v_24355;
wire v_24356;
wire v_24357;
wire v_24358;
wire v_24359;
wire v_24360;
wire v_24361;
wire v_24362;
wire v_24363;
wire v_24364;
wire v_24365;
wire v_24366;
wire v_24367;
wire v_24368;
wire v_24369;
wire v_24370;
wire v_24371;
wire v_24372;
wire v_24373;
wire v_24374;
wire v_24375;
wire v_24376;
wire v_24377;
wire v_24378;
wire v_24379;
wire v_24380;
wire v_24381;
wire v_24382;
wire v_24383;
wire v_24384;
wire v_24385;
wire v_24386;
wire v_24387;
wire v_24388;
wire v_24389;
wire v_24390;
wire v_24391;
wire v_24392;
wire v_24393;
wire v_24394;
wire v_24395;
wire v_24396;
wire v_24397;
wire v_24398;
wire v_24399;
wire v_24400;
wire v_24401;
wire v_24402;
wire v_24403;
wire v_24404;
wire v_24405;
wire v_24406;
wire v_24407;
wire v_24408;
wire v_24409;
wire v_24410;
wire v_24411;
wire v_24412;
wire v_24413;
wire v_24414;
wire v_24415;
wire v_24416;
wire v_24417;
wire v_24418;
wire v_24419;
wire v_24420;
wire v_24421;
wire v_24422;
wire v_24423;
wire v_24424;
wire v_24425;
wire v_24426;
wire v_24427;
wire v_24428;
wire v_24429;
wire v_24430;
wire v_24431;
wire v_24432;
wire v_24433;
wire v_24434;
wire v_24435;
wire v_24436;
wire v_24437;
wire v_24438;
wire v_24439;
wire v_24440;
wire v_24441;
wire v_24442;
wire v_24443;
wire v_24444;
wire v_24445;
wire v_24446;
wire v_24447;
wire v_24448;
wire v_24449;
wire v_24450;
wire v_24451;
wire v_24452;
wire v_24453;
wire v_24454;
wire v_24455;
wire v_24456;
wire v_24457;
wire v_24458;
wire v_24459;
wire v_24460;
wire v_24461;
wire v_24462;
wire v_24463;
wire v_24464;
wire v_24465;
wire v_24466;
wire v_24467;
wire v_24468;
wire v_24469;
wire v_24470;
wire v_24471;
wire v_24472;
wire v_24473;
wire v_24474;
wire v_24475;
wire v_24476;
wire v_24477;
wire v_24478;
wire v_24479;
wire v_24480;
wire v_24481;
wire v_24482;
wire v_24483;
wire v_24484;
wire v_24485;
wire v_24486;
wire v_24487;
wire v_24488;
wire v_24489;
wire v_24490;
wire v_24491;
wire v_24492;
wire v_24493;
wire v_24494;
wire v_24495;
wire v_24496;
wire v_24497;
wire v_24498;
wire v_24499;
wire v_24500;
wire v_24501;
wire v_24502;
wire v_24503;
wire v_24504;
wire v_24505;
wire v_24506;
wire v_24507;
wire v_24508;
wire v_24509;
wire v_24510;
wire v_24511;
wire v_24512;
wire v_24513;
wire v_24514;
wire v_24515;
wire v_24516;
wire v_24517;
wire v_24518;
wire v_24519;
wire v_24520;
wire v_24521;
wire v_24522;
wire v_24523;
wire v_24524;
wire v_24525;
wire v_24526;
wire v_24527;
wire v_24528;
wire v_24529;
wire v_24530;
wire v_24531;
wire v_24532;
wire v_24533;
wire v_24534;
wire v_24535;
wire v_24536;
wire v_24537;
wire v_24538;
wire v_24539;
wire v_24540;
wire v_24541;
wire v_24542;
wire v_24543;
wire v_24544;
wire v_24545;
wire v_24546;
wire v_24547;
wire v_24548;
wire v_24549;
wire v_24550;
wire v_24551;
wire v_24552;
wire v_24553;
wire v_24554;
wire v_24555;
wire v_24556;
wire v_24557;
wire v_24558;
wire v_24559;
wire v_24560;
wire v_24561;
wire v_24562;
wire v_24563;
wire v_24564;
wire v_24565;
wire v_24566;
wire v_24567;
wire v_24568;
wire v_24569;
wire v_24570;
wire v_24571;
wire v_24572;
wire v_24573;
wire v_24574;
wire v_24575;
wire v_24576;
wire v_24577;
wire v_24578;
wire v_24579;
wire v_24580;
wire v_24581;
wire v_24582;
wire v_24583;
wire v_24584;
wire v_24585;
wire v_24586;
wire v_24587;
wire v_24588;
wire v_24589;
wire v_24590;
wire v_24591;
wire v_24592;
wire v_24593;
wire v_24594;
wire v_24595;
wire v_24596;
wire v_24597;
wire v_24598;
wire v_24599;
wire v_24600;
wire v_24601;
wire v_24602;
wire v_24603;
wire v_24604;
wire v_24605;
wire v_24606;
wire v_24607;
wire v_24608;
wire v_24609;
wire v_24610;
wire v_24611;
wire v_24612;
wire v_24613;
wire v_24614;
wire v_24615;
wire v_24616;
wire v_24617;
wire v_24618;
wire v_24619;
wire v_24620;
wire v_24621;
wire v_24622;
wire v_24623;
wire v_24624;
wire v_24625;
wire v_24626;
wire v_24627;
wire v_24628;
wire v_24629;
wire v_24630;
wire v_24631;
wire v_24632;
wire v_24633;
wire v_24634;
wire v_24635;
wire v_24636;
wire v_24637;
wire v_24638;
wire v_24639;
wire v_24640;
wire v_24641;
wire v_24642;
wire v_24643;
wire v_24644;
wire v_24645;
wire v_24646;
wire v_24647;
wire v_24648;
wire v_24649;
wire v_24650;
wire v_24651;
wire v_24652;
wire v_24653;
wire v_24654;
wire v_24655;
wire v_24656;
wire v_24657;
wire v_24658;
wire v_24659;
wire v_24660;
wire v_24661;
wire v_24662;
wire v_24663;
wire v_24664;
wire v_24665;
wire v_24666;
wire v_24667;
wire v_24668;
wire v_24669;
wire v_24670;
wire v_24671;
wire v_24672;
wire v_24673;
wire v_24674;
wire v_24675;
wire v_24676;
wire v_24677;
wire v_24678;
wire v_24679;
wire v_24680;
wire v_24681;
wire v_24682;
wire v_24683;
wire v_24684;
wire v_24685;
wire v_24686;
wire v_24687;
wire v_24688;
wire v_24689;
wire v_24690;
wire v_24691;
wire v_24692;
wire v_24693;
wire v_24694;
wire v_24695;
wire v_24696;
wire v_24697;
wire v_24698;
wire v_24699;
wire v_24700;
wire v_24701;
wire v_24702;
wire v_24703;
wire v_24704;
wire v_24705;
wire v_24706;
wire v_24707;
wire v_24708;
wire v_24709;
wire v_24710;
wire v_24711;
wire v_24712;
wire v_24713;
wire v_24714;
wire v_24715;
wire v_24716;
wire v_24717;
wire v_24718;
wire v_24719;
wire v_24720;
wire v_24721;
wire v_24722;
wire v_24723;
wire v_24724;
wire v_24725;
wire v_24726;
wire v_24727;
wire v_24728;
wire v_24729;
wire v_24730;
wire v_24731;
wire v_24732;
wire v_24733;
wire v_24734;
wire v_24735;
wire v_24736;
wire v_24737;
wire v_24738;
wire v_24739;
wire v_24740;
wire v_24741;
wire v_24742;
wire v_24743;
wire v_24744;
wire v_24745;
wire v_24746;
wire v_24747;
wire v_24748;
wire v_24749;
wire v_24750;
wire v_24751;
wire v_24752;
wire v_24753;
wire v_24754;
wire v_24755;
wire v_24756;
wire v_24757;
wire v_24758;
wire v_24759;
wire v_24760;
wire v_24761;
wire v_24762;
wire v_24763;
wire v_24764;
wire v_24765;
wire v_24766;
wire v_24767;
wire v_24768;
wire v_24769;
wire v_24770;
wire v_24771;
wire v_24772;
wire v_24773;
wire v_24774;
wire v_24775;
wire v_24776;
wire v_24777;
wire v_24778;
wire v_24779;
wire v_24780;
wire v_24781;
wire v_24782;
wire v_24783;
wire v_24784;
wire v_24785;
wire v_24786;
wire v_24787;
wire v_24788;
wire v_24789;
wire v_24790;
wire v_24791;
wire v_24792;
wire v_24793;
wire v_24794;
wire v_24795;
wire v_24796;
wire v_24797;
wire v_24798;
wire v_24799;
wire v_24800;
wire v_24801;
wire v_24802;
wire v_24803;
wire v_24804;
wire v_24805;
wire v_24806;
wire v_24807;
wire v_24808;
wire v_24809;
wire v_24810;
wire v_24811;
wire v_24812;
wire v_24813;
wire v_24814;
wire v_24815;
wire v_24816;
wire v_24817;
wire v_24818;
wire v_24819;
wire v_24820;
wire v_24821;
wire v_24822;
wire v_24823;
wire v_24824;
wire v_24825;
wire v_24826;
wire v_24827;
wire v_24828;
wire v_24829;
wire v_24830;
wire v_24831;
wire v_24832;
wire v_24833;
wire v_24834;
wire v_24835;
wire v_24836;
wire v_24837;
wire v_24838;
wire v_24839;
wire v_24840;
wire v_24841;
wire v_24842;
wire v_24843;
wire v_24844;
wire v_24845;
wire v_24846;
wire v_24847;
wire v_24848;
wire v_24849;
wire v_24850;
wire v_24851;
wire v_24852;
wire v_24853;
wire v_24854;
wire v_24855;
wire v_24856;
wire v_24857;
wire v_24858;
wire v_24859;
wire v_24860;
wire v_24861;
wire v_24862;
wire v_24863;
wire v_24864;
wire v_24865;
wire v_24866;
wire v_24867;
wire v_24868;
wire v_24869;
wire v_24870;
wire v_24871;
wire v_24872;
wire v_24873;
wire v_24874;
wire v_24875;
wire v_24876;
wire v_24877;
wire v_24878;
wire v_24879;
wire v_24880;
wire v_24881;
wire v_24882;
wire v_24883;
wire v_24884;
wire v_24885;
wire v_24886;
wire v_24887;
wire v_24888;
wire v_24889;
wire v_24890;
wire v_24891;
wire v_24892;
wire v_24893;
wire v_24894;
wire v_24895;
wire v_24896;
wire v_24897;
wire v_24898;
wire v_24899;
wire v_24900;
wire v_24901;
wire v_24902;
wire v_24903;
wire v_24904;
wire v_24905;
wire v_24906;
wire v_24907;
wire v_24908;
wire v_24909;
wire v_24910;
wire v_24911;
wire v_24912;
wire v_24913;
wire v_24914;
wire v_24915;
wire v_24916;
wire v_24917;
wire v_24918;
wire v_24919;
wire v_24920;
wire v_24921;
wire v_24922;
wire v_24923;
wire v_24924;
wire v_24925;
wire v_24926;
wire v_24927;
wire v_24928;
wire v_24929;
wire v_24930;
wire v_24931;
wire v_24932;
wire v_24933;
wire v_24934;
wire v_24935;
wire v_24936;
wire v_24937;
wire v_24938;
wire v_24939;
wire v_24940;
wire v_24941;
wire v_24942;
wire v_24943;
wire v_24944;
wire v_24945;
wire v_24946;
wire v_24947;
wire v_24948;
wire v_24949;
wire v_24950;
wire v_24951;
wire v_24952;
wire v_24953;
wire v_24954;
wire v_24955;
wire v_24956;
wire v_24957;
wire v_24958;
wire v_24959;
wire v_24960;
wire v_24961;
wire v_24962;
wire v_24963;
wire v_24964;
wire v_24965;
wire v_24966;
wire v_24967;
wire v_24968;
wire v_24969;
wire v_24970;
wire v_24971;
wire v_24972;
wire v_24973;
wire v_24974;
wire v_24975;
wire v_24976;
wire v_24977;
wire v_24978;
wire v_24979;
wire v_24980;
wire v_24981;
wire v_24982;
wire v_24983;
wire v_24984;
wire v_24985;
wire v_24986;
wire v_24987;
wire v_24988;
wire v_24989;
wire v_24990;
wire v_24991;
wire v_24992;
wire v_24993;
wire v_24994;
wire v_24995;
wire v_24996;
wire v_24997;
wire v_24998;
wire v_24999;
wire v_25000;
wire v_25001;
wire v_25002;
wire v_25003;
wire v_25004;
wire v_25005;
wire v_25006;
wire v_25007;
wire v_25008;
wire v_25009;
wire v_25010;
wire v_25011;
wire v_25012;
wire v_25013;
wire v_25014;
wire v_25015;
wire v_25016;
wire v_25017;
wire v_25018;
wire v_25019;
wire v_25020;
wire v_25021;
wire v_25022;
wire v_25023;
wire v_25024;
wire v_25025;
wire v_25026;
wire v_25027;
wire v_25028;
wire v_25029;
wire v_25030;
wire v_25031;
wire v_25032;
wire v_25033;
wire v_25034;
wire v_25035;
wire v_25036;
wire v_25037;
wire v_25038;
wire v_25039;
wire v_25040;
wire v_25041;
wire v_25042;
wire v_25043;
wire v_25044;
wire v_25045;
wire v_25046;
wire v_25047;
wire v_25048;
wire v_25049;
wire v_25050;
wire v_25051;
wire v_25052;
wire v_25053;
wire v_25054;
wire v_25055;
wire v_25056;
wire v_25057;
wire v_25058;
wire v_25059;
wire v_25060;
wire v_25061;
wire v_25062;
wire v_25063;
wire v_25064;
wire v_25065;
wire v_25066;
wire v_25067;
wire v_25068;
wire v_25069;
wire v_25070;
wire v_25071;
wire v_25072;
wire v_25073;
wire v_25074;
wire v_25075;
wire v_25076;
wire v_25077;
wire v_25078;
wire v_25079;
wire v_25080;
wire v_25081;
wire v_25082;
wire v_25083;
wire v_25084;
wire v_25085;
wire v_25086;
wire v_25087;
wire v_25088;
wire v_25089;
wire v_25090;
wire v_25091;
wire v_25092;
wire v_25093;
wire v_25094;
wire v_25095;
wire v_25096;
wire v_25097;
wire v_25098;
wire v_25099;
wire v_25100;
wire v_25101;
wire v_25102;
wire v_25103;
wire v_25104;
wire v_25105;
wire v_25106;
wire v_25107;
wire v_25108;
wire v_25109;
wire v_25110;
wire v_25111;
wire v_25112;
wire v_25113;
wire v_25114;
wire v_25115;
wire v_25116;
wire v_25117;
wire v_25118;
wire v_25119;
wire v_25120;
wire v_25121;
wire v_25122;
wire v_25123;
wire v_25124;
wire v_25125;
wire v_25126;
wire v_25127;
wire v_25128;
wire v_25129;
wire v_25130;
wire v_25131;
wire v_25132;
wire v_25133;
wire v_25134;
wire v_25135;
wire v_25136;
wire v_25137;
wire v_25138;
wire v_25139;
wire v_25140;
wire v_25141;
wire v_25142;
wire v_25143;
wire v_25144;
wire v_25145;
wire v_25146;
wire v_25147;
wire v_25148;
wire v_25149;
wire v_25150;
wire v_25151;
wire v_25152;
wire v_25153;
wire v_25154;
wire v_25155;
wire v_25156;
wire v_25157;
wire v_25158;
wire v_25159;
wire v_25160;
wire v_25161;
wire v_25162;
wire v_25163;
wire v_25164;
wire v_25165;
wire v_25166;
wire v_25167;
wire v_25168;
wire v_25169;
wire v_25170;
wire v_25171;
wire v_25172;
wire v_25173;
wire v_25174;
wire v_25175;
wire v_25176;
wire v_25177;
wire v_25178;
wire v_25179;
wire v_25180;
wire v_25181;
wire v_25182;
wire v_25183;
wire v_25184;
wire v_25185;
wire v_25186;
wire v_25187;
wire v_25188;
wire v_25189;
wire v_25190;
wire v_25191;
wire v_25192;
wire v_25193;
wire v_25194;
wire v_25195;
wire v_25196;
wire v_25197;
wire v_25198;
wire v_25199;
wire v_25200;
wire v_25201;
wire v_25202;
wire v_25203;
wire v_25204;
wire v_25205;
wire v_25206;
wire v_25207;
wire v_25208;
wire v_25209;
wire v_25210;
wire v_25211;
wire v_25212;
wire v_25213;
wire v_25214;
wire v_25215;
wire v_25216;
wire v_25217;
wire v_25218;
wire v_25219;
wire v_25220;
wire v_25221;
wire v_25222;
wire v_25223;
wire v_25224;
wire v_25225;
wire v_25226;
wire v_25227;
wire v_25228;
wire v_25229;
wire v_25230;
wire v_25231;
wire v_25232;
wire v_25233;
wire v_25234;
wire v_25235;
wire v_25236;
wire v_25237;
wire v_25238;
wire v_25239;
wire v_25240;
wire v_25241;
wire v_25242;
wire v_25243;
wire v_25244;
wire v_25245;
wire v_25246;
wire v_25247;
wire v_25248;
wire v_25249;
wire v_25250;
wire v_25251;
wire v_25252;
wire v_25253;
wire v_25254;
wire v_25255;
wire v_25256;
wire v_25257;
wire v_25258;
wire v_25259;
wire v_25260;
wire v_25261;
wire v_25262;
wire v_25263;
wire v_25264;
wire v_25265;
wire v_25266;
wire v_25267;
wire v_25268;
wire v_25269;
wire v_25270;
wire v_25271;
wire v_25272;
wire v_25273;
wire v_25274;
wire v_25275;
wire v_25276;
wire v_25277;
wire v_25278;
wire v_25279;
wire v_25280;
wire v_25281;
wire v_25282;
wire v_25283;
wire v_25284;
wire v_25285;
wire v_25286;
wire v_25287;
wire v_25288;
wire v_25289;
wire v_25290;
wire v_25291;
wire v_25292;
wire v_25293;
wire v_25294;
wire v_25295;
wire v_25296;
wire v_25297;
wire v_25298;
wire v_25299;
wire v_25300;
wire v_25301;
wire v_25302;
wire v_25303;
wire v_25304;
wire v_25305;
wire v_25306;
wire v_25307;
wire v_25308;
wire v_25309;
wire v_25310;
wire v_25311;
wire v_25312;
wire v_25313;
wire v_25314;
wire v_25315;
wire v_25316;
wire v_25317;
wire v_25318;
wire v_25319;
wire v_25320;
wire v_25321;
wire v_25322;
wire v_25323;
wire v_25324;
wire v_25325;
wire v_25326;
wire v_25327;
wire v_25328;
wire v_25329;
wire v_25330;
wire v_25331;
wire v_25332;
wire v_25333;
wire v_25334;
wire v_25335;
wire v_25336;
wire v_25337;
wire v_25338;
wire v_25339;
wire v_25340;
wire v_25341;
wire v_25342;
wire v_25343;
wire v_25344;
wire v_25345;
wire v_25346;
wire v_25347;
wire v_25348;
wire v_25349;
wire v_25350;
wire v_25351;
wire v_25352;
wire v_25353;
wire v_25354;
wire v_25355;
wire v_25356;
wire v_25357;
wire v_25358;
wire v_25359;
wire v_25360;
wire v_25361;
wire v_25362;
wire v_25363;
wire v_25364;
wire v_25365;
wire v_25366;
wire v_25367;
wire v_25368;
wire v_25369;
wire v_25370;
wire v_25371;
wire v_25372;
wire v_25373;
wire v_25374;
wire v_25375;
wire v_25376;
wire v_25377;
wire v_25378;
wire v_25379;
wire v_25380;
wire v_25381;
wire v_25382;
wire v_25383;
wire v_25384;
wire v_25385;
wire v_25386;
wire v_25387;
wire v_25388;
wire v_25389;
wire v_25390;
wire v_25391;
wire v_25392;
wire v_25393;
wire v_25394;
wire v_25395;
wire v_25396;
wire v_25397;
wire v_25398;
wire v_25399;
wire v_25400;
wire v_25401;
wire v_25402;
wire v_25403;
wire v_25404;
wire v_25405;
wire v_25406;
wire v_25407;
wire v_25408;
wire v_25409;
wire v_25410;
wire v_25411;
wire v_25412;
wire v_25413;
wire v_25414;
wire v_25415;
wire v_25416;
wire v_25417;
wire v_25418;
wire v_25419;
wire v_25420;
wire v_25421;
wire v_25422;
wire v_25423;
wire v_25424;
wire v_25425;
wire v_25426;
wire v_25427;
wire v_25428;
wire v_25429;
wire v_25430;
wire v_25431;
wire v_25432;
wire v_25433;
wire v_25434;
wire v_25435;
wire v_25436;
wire v_25437;
wire v_25438;
wire v_25439;
wire v_25440;
wire v_25441;
wire v_25442;
wire v_25443;
wire v_25444;
wire v_25445;
wire v_25446;
wire v_25447;
wire v_25448;
wire v_25449;
wire v_25450;
wire v_25451;
wire v_25452;
wire v_25453;
wire v_25454;
wire v_25455;
wire v_25456;
wire v_25457;
wire v_25458;
wire v_25459;
wire v_25460;
wire v_25461;
wire v_25462;
wire v_25463;
wire v_25464;
wire v_25465;
wire v_25466;
wire v_25467;
wire v_25468;
wire v_25469;
wire v_25470;
wire v_25471;
wire v_25472;
wire v_25473;
wire v_25474;
wire v_25475;
wire v_25476;
wire v_25477;
wire v_25478;
wire v_25479;
wire v_25480;
wire v_25481;
wire v_25482;
wire v_25483;
wire v_25484;
wire v_25485;
wire v_25486;
wire v_25487;
wire v_25488;
wire v_25489;
wire v_25490;
wire v_25491;
wire v_25492;
wire v_25493;
wire v_25494;
wire v_25495;
wire v_25496;
wire v_25497;
wire v_25498;
wire v_25499;
wire v_25500;
wire v_25501;
wire v_25502;
wire v_25503;
wire v_25504;
wire v_25505;
wire v_25506;
wire v_25507;
wire v_25508;
wire v_25509;
wire v_25510;
wire v_25511;
wire v_25512;
wire v_25513;
wire v_25514;
wire v_25515;
wire v_25516;
wire v_25517;
wire v_25518;
wire v_25519;
wire v_25520;
wire v_25521;
wire v_25522;
wire v_25523;
wire v_25524;
wire v_25525;
wire v_25526;
wire v_25527;
wire v_25528;
wire v_25529;
wire v_25530;
wire v_25531;
wire v_25532;
wire v_25533;
wire v_25534;
wire v_25535;
wire v_25536;
wire v_25537;
wire v_25538;
wire v_25539;
wire v_25540;
wire v_25541;
wire v_25542;
wire v_25543;
wire v_25544;
wire v_25545;
wire v_25546;
wire v_25547;
wire v_25548;
wire v_25549;
wire v_25550;
wire v_25551;
wire v_25552;
wire v_25553;
wire v_25554;
wire v_25555;
wire v_25556;
wire v_25557;
wire v_25558;
wire v_25559;
wire v_25560;
wire v_25561;
wire v_25562;
wire v_25563;
wire v_25564;
wire v_25565;
wire v_25566;
wire v_25567;
wire v_25568;
wire v_25569;
wire v_25570;
wire v_25571;
wire v_25572;
wire v_25573;
wire v_25574;
wire v_25575;
wire v_25576;
wire v_25577;
wire v_25578;
wire v_25579;
wire v_25580;
wire v_25581;
wire v_25582;
wire v_25583;
wire v_25584;
wire v_25585;
wire v_25586;
wire v_25587;
wire v_25588;
wire v_25589;
wire v_25590;
wire v_25591;
wire v_25592;
wire v_25593;
wire v_25594;
wire v_25595;
wire v_25596;
wire v_25597;
wire v_25598;
wire v_25599;
wire v_25600;
wire v_25601;
wire v_25602;
wire v_25603;
wire v_25604;
wire v_25605;
wire v_25606;
wire v_25607;
wire v_25608;
wire v_25609;
wire v_25610;
wire v_25611;
wire v_25612;
wire v_25613;
wire v_25614;
wire v_25615;
wire v_25616;
wire v_25617;
wire v_25618;
wire v_25619;
wire v_25620;
wire v_25621;
wire v_25622;
wire v_25623;
wire v_25624;
wire v_25625;
wire v_25626;
wire v_25627;
wire v_25628;
wire v_25629;
wire v_25630;
wire v_25631;
wire v_25632;
wire v_25633;
wire v_25634;
wire v_25635;
wire v_25636;
wire v_25637;
wire v_25638;
wire v_25639;
wire v_25640;
wire v_25641;
wire v_25642;
wire v_25643;
wire v_25644;
wire v_25645;
wire v_25646;
wire v_25647;
wire v_25648;
wire v_25649;
wire v_25650;
wire v_25651;
wire v_25652;
wire v_25653;
wire v_25654;
wire v_25655;
wire v_25656;
wire v_25657;
wire v_25658;
wire v_25659;
wire v_25660;
wire v_25661;
wire v_25662;
wire v_25663;
wire v_25664;
wire v_25665;
wire v_25666;
wire v_25667;
wire v_25668;
wire v_25669;
wire v_25670;
wire v_25671;
wire v_25672;
wire v_25673;
wire v_25674;
wire v_25675;
wire v_25676;
wire v_25677;
wire v_25678;
wire v_25679;
wire v_25680;
wire v_25681;
wire v_25682;
wire v_25683;
wire v_25684;
wire v_25685;
wire v_25686;
wire v_25687;
wire v_25688;
wire v_25689;
wire v_25690;
wire v_25691;
wire v_25692;
wire v_25693;
wire v_25694;
wire v_25695;
wire v_25696;
wire v_25697;
wire v_25698;
wire v_25699;
wire v_25700;
wire v_25701;
wire v_25702;
wire v_25703;
wire v_25704;
wire v_25705;
wire v_25706;
wire v_25707;
wire v_25708;
wire v_25709;
wire v_25710;
wire v_25711;
wire v_25712;
wire v_25713;
wire v_25714;
wire v_25715;
wire v_25716;
wire v_25717;
wire v_25718;
wire v_25719;
wire v_25720;
wire v_25721;
wire v_25722;
wire v_25723;
wire v_25724;
wire v_25725;
wire v_25726;
wire v_25727;
wire v_25728;
wire v_25729;
wire v_25730;
wire v_25731;
wire v_25732;
wire v_25733;
wire v_25734;
wire v_25735;
wire v_25736;
wire v_25737;
wire v_25738;
wire v_25739;
wire v_25740;
wire v_25741;
wire v_25742;
wire v_25743;
wire v_25744;
wire v_25745;
wire v_25746;
wire v_25747;
wire v_25748;
wire v_25749;
wire v_25750;
wire v_25751;
wire v_25752;
wire v_25753;
wire v_25754;
wire v_25755;
wire v_25756;
wire v_25757;
wire v_25758;
wire v_25759;
wire v_25760;
wire v_25761;
wire v_25762;
wire v_25763;
wire v_25764;
wire v_25765;
wire v_25766;
wire v_25767;
wire v_25768;
wire v_25769;
wire v_25770;
wire v_25771;
wire v_25772;
wire v_25773;
wire v_25774;
wire v_25775;
wire v_25776;
wire v_25777;
wire v_25778;
wire v_25779;
wire v_25780;
wire v_25781;
wire v_25782;
wire v_25783;
wire v_25784;
wire v_25785;
wire v_25786;
wire v_25787;
wire v_25788;
wire v_25789;
wire v_25790;
wire v_25791;
wire v_25792;
wire v_25793;
wire v_25794;
wire v_25795;
wire v_25796;
wire v_25797;
wire v_25798;
wire v_25799;
wire v_25800;
wire v_25801;
wire v_25802;
wire v_25803;
wire v_25804;
wire v_25805;
wire v_25806;
wire v_25807;
wire v_25808;
wire v_25809;
wire v_25810;
wire v_25811;
wire v_25812;
wire v_25813;
wire v_25814;
wire v_25815;
wire v_25816;
wire v_25817;
wire v_25818;
wire v_25819;
wire v_25820;
wire v_25821;
wire v_25822;
wire v_25823;
wire v_25824;
wire v_25825;
wire v_25826;
wire v_25827;
wire v_25828;
wire v_25829;
wire v_25830;
wire v_25831;
wire v_25832;
wire v_25833;
wire v_25834;
wire v_25835;
wire v_25836;
wire v_25837;
wire v_25838;
wire v_25839;
wire v_25840;
wire v_25841;
wire v_25842;
wire v_25843;
wire v_25844;
wire v_25845;
wire v_25846;
wire v_25847;
wire v_25848;
wire v_25849;
wire v_25850;
wire v_25851;
wire v_25852;
wire v_25853;
wire v_25854;
wire v_25855;
wire v_25856;
wire v_25857;
wire v_25858;
wire v_25859;
wire v_25860;
wire v_25861;
wire v_25862;
wire v_25863;
wire v_25864;
wire v_25865;
wire v_25866;
wire v_25867;
wire v_25868;
wire v_25869;
wire v_25870;
wire v_25871;
wire v_25872;
wire v_25873;
wire v_25874;
wire v_25875;
wire v_25876;
wire v_25877;
wire v_25878;
wire v_25879;
wire v_25880;
wire v_25881;
wire v_25882;
wire v_25883;
wire v_25884;
wire v_25885;
wire v_25886;
wire v_25887;
wire v_25888;
wire v_25889;
wire v_25890;
wire v_25891;
wire v_25892;
wire v_25893;
wire v_25894;
wire v_25895;
wire v_25896;
wire v_25897;
wire v_25898;
wire v_25899;
wire v_25900;
wire v_25901;
wire v_25902;
wire v_25903;
wire v_25904;
wire v_25905;
wire v_25906;
wire v_25907;
wire v_25908;
wire v_25909;
wire v_25910;
wire v_25911;
wire v_25912;
wire v_25913;
wire v_25914;
wire v_25915;
wire v_25916;
wire v_25917;
wire v_25918;
wire v_25919;
wire v_25920;
wire v_25921;
wire v_25922;
wire v_25923;
wire v_25924;
wire v_25925;
wire v_25926;
wire v_25927;
wire v_25928;
wire v_25929;
wire v_25930;
wire v_25931;
wire v_25932;
wire v_25933;
wire v_25934;
wire v_25935;
wire v_25936;
wire v_25937;
wire v_25938;
wire v_25939;
wire v_25940;
wire v_25941;
wire v_25942;
wire v_25943;
wire v_25944;
wire v_25945;
wire v_25946;
wire v_25947;
wire v_25948;
wire v_25949;
wire v_25950;
wire v_25951;
wire v_25952;
wire v_25953;
wire v_25954;
wire v_25955;
wire v_25956;
wire v_25957;
wire v_25958;
wire v_25959;
wire v_25960;
wire v_25961;
wire v_25962;
wire v_25963;
wire v_25964;
wire v_25965;
wire v_25966;
wire v_25967;
wire v_25968;
wire v_25969;
wire v_25970;
wire v_25971;
wire v_25972;
wire v_25973;
wire v_25974;
wire v_25975;
wire v_25976;
wire v_25977;
wire v_25978;
wire v_25979;
wire v_25980;
wire v_25981;
wire v_25982;
wire v_25983;
wire v_25984;
wire v_25985;
wire v_25986;
wire v_25987;
wire v_25988;
wire v_25989;
wire v_25990;
wire v_25991;
wire v_25992;
wire v_25993;
wire v_25994;
wire v_25995;
wire v_25996;
wire v_25997;
wire v_25998;
wire v_25999;
wire v_26000;
wire v_26001;
wire v_26002;
wire v_26003;
wire v_26004;
wire v_26005;
wire v_26006;
wire v_26007;
wire v_26008;
wire v_26009;
wire v_26010;
wire v_26011;
wire v_26012;
wire v_26013;
wire v_26014;
wire v_26015;
wire v_26016;
wire v_26017;
wire v_26018;
wire v_26019;
wire v_26020;
wire v_26021;
wire v_26022;
wire v_26023;
wire v_26024;
wire v_26025;
wire v_26026;
wire v_26027;
wire v_26028;
wire v_26029;
wire v_26030;
wire v_26031;
wire v_26032;
wire v_26033;
wire v_26034;
wire v_26035;
wire v_26036;
wire v_26037;
wire v_26038;
wire v_26039;
wire v_26040;
wire v_26041;
wire v_26042;
wire v_26043;
wire v_26044;
wire v_26045;
wire v_26046;
wire v_26047;
wire v_26048;
wire v_26049;
wire v_26050;
wire v_26051;
wire v_26052;
wire v_26053;
wire v_26054;
wire v_26055;
wire v_26056;
wire v_26057;
wire v_26058;
wire v_26059;
wire v_26060;
wire v_26061;
wire v_26062;
wire v_26063;
wire v_26064;
wire v_26065;
wire v_26066;
wire v_26067;
wire v_26068;
wire v_26069;
wire v_26070;
wire v_26071;
wire v_26072;
wire v_26073;
wire v_26074;
wire v_26075;
wire v_26076;
wire v_26077;
wire v_26078;
wire v_26079;
wire v_26080;
wire v_26081;
wire v_26082;
wire v_26083;
wire v_26084;
wire v_26085;
wire v_26086;
wire v_26087;
wire v_26088;
wire v_26089;
wire v_26090;
wire v_26091;
wire v_26092;
wire v_26093;
wire v_26094;
wire v_26095;
wire v_26096;
wire v_26097;
wire v_26098;
wire v_26099;
wire v_26100;
wire v_26101;
wire v_26102;
wire v_26103;
wire v_26104;
wire v_26105;
wire v_26106;
wire v_26107;
wire v_26108;
wire v_26109;
wire v_26110;
wire v_26111;
wire v_26112;
wire v_26113;
wire v_26114;
wire v_26115;
wire v_26116;
wire v_26117;
wire v_26118;
wire v_26119;
wire v_26120;
wire v_26121;
wire v_26122;
wire v_26123;
wire v_26124;
wire v_26125;
wire v_26126;
wire v_26127;
wire v_26128;
wire v_26129;
wire v_26130;
wire v_26131;
wire v_26132;
wire v_26133;
wire v_26134;
wire v_26135;
wire v_26136;
wire v_26137;
wire v_26138;
wire v_26139;
wire v_26140;
wire v_26141;
wire v_26142;
wire v_26143;
wire v_26144;
wire v_26145;
wire v_26146;
wire v_26147;
wire v_26148;
wire v_26149;
wire v_26150;
wire v_26151;
wire v_26152;
wire v_26153;
wire v_26154;
wire v_26155;
wire v_26156;
wire v_26157;
wire v_26158;
wire v_26159;
wire v_26160;
wire v_26161;
wire v_26162;
wire v_26163;
wire v_26164;
wire v_26165;
wire v_26166;
wire v_26167;
wire v_26168;
wire v_26169;
wire v_26170;
wire v_26171;
wire v_26172;
wire v_26173;
wire v_26174;
wire v_26175;
wire v_26176;
wire v_26177;
wire v_26178;
wire v_26179;
wire v_26180;
wire v_26181;
wire v_26182;
wire v_26183;
wire v_26184;
wire v_26185;
wire v_26186;
wire v_26187;
wire v_26188;
wire v_26189;
wire v_26190;
wire v_26191;
wire v_26192;
wire v_26193;
wire v_26194;
wire v_26195;
wire v_26196;
wire v_26197;
wire v_26198;
wire v_26199;
wire v_26200;
wire v_26201;
wire v_26202;
wire v_26203;
wire v_26204;
wire v_26205;
wire v_26206;
wire v_26207;
wire v_26208;
wire v_26209;
wire v_26210;
wire v_26211;
wire v_26212;
wire v_26213;
wire v_26214;
wire v_26215;
wire v_26216;
wire v_26217;
wire v_26218;
wire v_26219;
wire v_26220;
wire v_26221;
wire v_26222;
wire v_26223;
wire v_26224;
wire v_26225;
wire v_26226;
wire v_26227;
wire v_26228;
wire v_26229;
wire v_26230;
wire v_26231;
wire v_26232;
wire v_26233;
wire v_26234;
wire v_26235;
wire v_26236;
wire v_26237;
wire v_26238;
wire v_26239;
wire v_26240;
wire v_26241;
wire v_26242;
wire v_26243;
wire v_26244;
wire v_26245;
wire v_26246;
wire v_26247;
wire v_26248;
wire v_26249;
wire v_26250;
wire v_26251;
wire v_26252;
wire v_26253;
wire v_26254;
wire v_26255;
wire v_26256;
wire v_26257;
wire v_26258;
wire v_26259;
wire v_26260;
wire v_26261;
wire v_26262;
wire v_26263;
wire v_26264;
wire v_26265;
wire v_26266;
wire v_26267;
wire v_26268;
wire v_26269;
wire v_26270;
wire v_26271;
wire v_26272;
wire v_26273;
wire v_26274;
wire v_26275;
wire v_26276;
wire v_26277;
wire v_26278;
wire v_26279;
wire v_26280;
wire v_26281;
wire v_26282;
wire v_26283;
wire v_26284;
wire v_26285;
wire v_26286;
wire v_26287;
wire v_26288;
wire v_26289;
wire v_26290;
wire v_26291;
wire v_26292;
wire v_26293;
wire v_26294;
wire v_26295;
wire v_26296;
wire v_26297;
wire v_26298;
wire v_26299;
wire v_26300;
wire v_26301;
wire v_26302;
wire v_26303;
wire v_26304;
wire v_26305;
wire v_26306;
wire v_26307;
wire v_26308;
wire v_26309;
wire v_26310;
wire v_26311;
wire v_26312;
wire v_26313;
wire v_26314;
wire v_26315;
wire v_26316;
wire v_26317;
wire v_26318;
wire v_26319;
wire v_26320;
wire v_26321;
wire v_26322;
wire v_26323;
wire v_26324;
wire v_26325;
wire v_26326;
wire v_26327;
wire v_26328;
wire v_26329;
wire v_26330;
wire v_26331;
wire v_26332;
wire v_26333;
wire v_26334;
wire v_26335;
wire v_26336;
wire v_26337;
wire v_26338;
wire v_26339;
wire v_26340;
wire v_26341;
wire v_26342;
wire v_26343;
wire v_26344;
wire v_26345;
wire v_26346;
wire v_26347;
wire v_26348;
wire v_26349;
wire v_26350;
wire v_26351;
wire v_26352;
wire v_26353;
wire v_26354;
wire v_26355;
wire v_26356;
wire v_26357;
wire v_26358;
wire v_26359;
wire v_26360;
wire v_26361;
wire v_26362;
wire v_26363;
wire v_26364;
wire v_26365;
wire v_26366;
wire v_26367;
wire v_26368;
wire v_26369;
wire v_26370;
wire v_26371;
wire v_26372;
wire v_26373;
wire v_26374;
wire v_26375;
wire v_26376;
wire v_26377;
wire v_26378;
wire v_26379;
wire v_26380;
wire v_26381;
wire v_26382;
wire v_26383;
wire v_26384;
wire v_26385;
wire v_26386;
wire v_26387;
wire v_26388;
wire v_26389;
wire v_26390;
wire v_26391;
wire v_26392;
wire v_26393;
wire v_26394;
wire v_26395;
wire v_26396;
wire v_26397;
wire v_26398;
wire v_26399;
wire v_26400;
wire v_26401;
wire v_26402;
wire v_26403;
wire v_26404;
wire v_26405;
wire v_26406;
wire v_26407;
wire v_26408;
wire v_26409;
wire v_26410;
wire v_26411;
wire v_26412;
wire v_26413;
wire v_26414;
wire v_26415;
wire v_26416;
wire v_26417;
wire v_26418;
wire v_26419;
wire v_26420;
wire v_26421;
wire v_26422;
wire v_26423;
wire v_26424;
wire v_26425;
wire v_26426;
wire v_26427;
wire v_26428;
wire v_26429;
wire v_26430;
wire v_26431;
wire v_26432;
wire v_26433;
wire v_26434;
wire v_26435;
wire v_26436;
wire v_26437;
wire v_26438;
wire v_26439;
wire v_26440;
wire v_26441;
wire v_26442;
wire v_26443;
wire v_26444;
wire v_26445;
wire v_26446;
wire v_26447;
wire v_26448;
wire v_26449;
wire v_26450;
wire v_26451;
wire v_26452;
wire v_26453;
wire v_26454;
wire v_26455;
wire v_26456;
wire v_26457;
wire v_26458;
wire v_26459;
wire v_26460;
wire v_26461;
wire v_26462;
wire v_26463;
wire v_26464;
wire v_26465;
wire v_26466;
wire v_26467;
wire v_26468;
wire v_26469;
wire v_26470;
wire v_26471;
wire v_26472;
wire v_26473;
wire v_26474;
wire v_26475;
wire v_26476;
wire v_26477;
wire v_26478;
wire v_26479;
wire v_26480;
wire v_26481;
wire v_26482;
wire v_26483;
wire v_26484;
wire v_26485;
wire v_26486;
wire v_26487;
wire v_26488;
wire v_26489;
wire v_26490;
wire v_26491;
wire v_26492;
wire v_26493;
wire v_26494;
wire v_26495;
wire v_26496;
wire v_26497;
wire v_26498;
wire v_26499;
wire v_26500;
wire v_26501;
wire v_26502;
wire v_26503;
wire v_26504;
wire v_26505;
wire v_26506;
wire v_26507;
wire v_26508;
wire v_26509;
wire v_26510;
wire v_26511;
wire v_26512;
wire v_26513;
wire v_26514;
wire v_26515;
wire v_26516;
wire v_26517;
wire v_26518;
wire v_26519;
wire v_26520;
wire v_26521;
wire v_26522;
wire v_26523;
wire v_26524;
wire v_26525;
wire v_26526;
wire v_26527;
wire v_26528;
wire v_26529;
wire v_26530;
wire v_26531;
wire v_26532;
wire v_26533;
wire v_26534;
wire v_26535;
wire v_26536;
wire v_26537;
wire v_26538;
wire v_26539;
wire v_26540;
wire v_26541;
wire v_26542;
wire v_26543;
wire v_26544;
wire v_26545;
wire v_26546;
wire v_26547;
wire v_26548;
wire v_26549;
wire v_26550;
wire v_26551;
wire v_26552;
wire v_26553;
wire v_26554;
wire v_26555;
wire v_26556;
wire v_26557;
wire v_26558;
wire v_26559;
wire v_26560;
wire v_26561;
wire v_26562;
wire v_26563;
wire v_26564;
wire v_26565;
wire v_26566;
wire v_26567;
wire v_26568;
wire v_26569;
wire v_26570;
wire v_26571;
wire v_26572;
wire v_26573;
wire v_26574;
wire v_26575;
wire v_26576;
wire v_26577;
wire v_26578;
wire v_26579;
wire v_26580;
wire v_26581;
wire v_26582;
wire v_26583;
wire v_26584;
wire v_26585;
wire v_26586;
wire v_26587;
wire v_26588;
wire v_26589;
wire v_26590;
wire v_26591;
wire v_26592;
wire v_26593;
wire v_26594;
wire v_26595;
wire v_26596;
wire v_26597;
wire v_26598;
wire v_26599;
wire v_26600;
wire v_26601;
wire v_26602;
wire v_26603;
wire v_26604;
wire v_26605;
wire v_26606;
wire v_26607;
wire v_26608;
wire v_26609;
wire v_26610;
wire v_26611;
wire v_26612;
wire v_26613;
wire v_26614;
wire v_26615;
wire v_26616;
wire v_26617;
wire v_26618;
wire v_26619;
wire v_26620;
wire v_26621;
wire v_26622;
wire v_26623;
wire v_26624;
wire v_26625;
wire v_26626;
wire v_26627;
wire v_26628;
wire v_26629;
wire v_26630;
wire v_26631;
wire v_26632;
wire v_26633;
wire v_26634;
wire v_26635;
wire v_26636;
wire v_26637;
wire v_26638;
wire v_26639;
wire v_26640;
wire v_26641;
wire v_26642;
wire v_26643;
wire v_26644;
wire v_26645;
wire v_26646;
wire v_26647;
wire v_26648;
wire v_26649;
wire v_26650;
wire v_26651;
wire v_26652;
wire v_26653;
wire v_26654;
wire v_26655;
wire v_26656;
wire v_26657;
wire v_26658;
wire v_26659;
wire v_26660;
wire v_26661;
wire v_26662;
wire v_26663;
wire v_26664;
wire v_26665;
wire v_26666;
wire v_26667;
wire v_26668;
wire v_26669;
wire v_26670;
wire v_26671;
wire v_26672;
wire v_26673;
wire v_26674;
wire v_26675;
wire v_26676;
wire v_26677;
wire v_26678;
wire v_26679;
wire v_26680;
wire v_26681;
wire v_26682;
wire v_26683;
wire v_26684;
wire v_26685;
wire v_26686;
wire v_26687;
wire v_26688;
wire v_26689;
wire v_26690;
wire v_26691;
wire v_26692;
wire v_26693;
wire v_26694;
wire v_26695;
wire v_26696;
wire v_26697;
wire v_26698;
wire v_26699;
wire v_26700;
wire v_26701;
wire v_26702;
wire v_26703;
wire v_26704;
wire v_26705;
wire v_26706;
wire v_26707;
wire v_26708;
wire v_26709;
wire v_26710;
wire v_26711;
wire v_26712;
wire v_26713;
wire v_26714;
wire v_26715;
wire v_26716;
wire v_26717;
wire v_26718;
wire v_26719;
wire v_26720;
wire v_26721;
wire v_26722;
wire v_26723;
wire v_26724;
wire v_26725;
wire v_26726;
wire v_26727;
wire v_26728;
wire v_26729;
wire v_26730;
wire v_26731;
wire v_26732;
wire v_26733;
wire v_26734;
wire v_26735;
wire v_26736;
wire v_26737;
wire v_26738;
wire v_26739;
wire v_26740;
wire v_26741;
wire v_26742;
wire v_26743;
wire v_26744;
wire v_26745;
wire v_26746;
wire v_26747;
wire v_26748;
wire v_26749;
wire v_26750;
wire v_26751;
wire v_26752;
wire v_26753;
wire v_26754;
wire v_26755;
wire v_26756;
wire v_26757;
wire v_26758;
wire v_26759;
wire v_26760;
wire v_26761;
wire v_26762;
wire v_26763;
wire v_26764;
wire v_26765;
wire v_26766;
wire v_26767;
wire v_26768;
wire v_26769;
wire v_26770;
wire v_26771;
wire v_26772;
wire v_26773;
wire v_26774;
wire v_26775;
wire v_26776;
wire v_26777;
wire v_26778;
wire v_26779;
wire v_26780;
wire v_26781;
wire v_26782;
wire v_26783;
wire v_26784;
wire v_26785;
wire v_26786;
wire v_26787;
wire v_26788;
wire v_26789;
wire v_26790;
wire v_26791;
wire v_26792;
wire v_26793;
wire v_26794;
wire v_26795;
wire v_26796;
wire v_26797;
wire v_26798;
wire v_26799;
wire v_26800;
wire v_26801;
wire v_26802;
wire v_26803;
wire v_26804;
wire v_26805;
wire v_26806;
wire v_26807;
wire v_26808;
wire v_26809;
wire v_26810;
wire v_26811;
wire v_26812;
wire v_26813;
wire v_26814;
wire v_26815;
wire v_26816;
wire v_26817;
wire v_26818;
wire v_26819;
wire v_26820;
wire v_26821;
wire v_26822;
wire v_26823;
wire v_26824;
wire v_26825;
wire v_26826;
wire v_26827;
wire v_26828;
wire v_26829;
wire v_26830;
wire v_26831;
wire v_26832;
wire v_26833;
wire v_26834;
wire v_26835;
wire v_26836;
wire v_26837;
wire v_26838;
wire v_26839;
wire v_26840;
wire v_26841;
wire v_26842;
wire v_26843;
wire v_26844;
wire v_26845;
wire v_26846;
wire v_26847;
wire v_26848;
wire v_26849;
wire v_26850;
wire v_26851;
wire v_26852;
wire v_26853;
wire v_26854;
wire v_26855;
wire v_26856;
wire v_26857;
wire v_26858;
wire v_26859;
wire v_26860;
wire v_26861;
wire v_26862;
wire v_26863;
wire v_26864;
wire v_26865;
wire v_26866;
wire v_26867;
wire v_26868;
wire v_26869;
wire v_26870;
wire v_26871;
wire v_26872;
wire v_26873;
wire v_26874;
wire v_26875;
wire v_26876;
wire v_26877;
wire v_26878;
wire v_26879;
wire v_26880;
wire v_26881;
wire v_26882;
wire v_26883;
wire v_26884;
wire v_26885;
wire v_26886;
wire v_26887;
wire v_26888;
wire v_26889;
wire v_26890;
wire v_26891;
wire v_26892;
wire v_26893;
wire v_26894;
wire v_26895;
wire v_26896;
wire v_26897;
wire v_26898;
wire v_26899;
wire v_26900;
wire v_26901;
wire v_26902;
wire v_26903;
wire v_26904;
wire v_26905;
wire v_26906;
wire v_26907;
wire v_26908;
wire v_26909;
wire v_26910;
wire v_26911;
wire v_26912;
wire v_26913;
wire v_26914;
wire v_26915;
wire v_26916;
wire v_26917;
wire v_26918;
wire v_26919;
wire v_26920;
wire v_26921;
wire v_26922;
wire v_26923;
wire v_26924;
wire v_26925;
wire v_26926;
wire v_26927;
wire v_26928;
wire v_26929;
wire v_26930;
wire v_26931;
wire v_26932;
wire v_26933;
wire v_26934;
wire v_26935;
wire v_26936;
wire v_26937;
wire v_26938;
wire v_26939;
wire v_26940;
wire v_26941;
wire v_26942;
wire v_26943;
wire v_26944;
wire v_26945;
wire v_26946;
wire v_26947;
wire v_26948;
wire v_26949;
wire v_26950;
wire v_26951;
wire v_26952;
wire v_26953;
wire v_26954;
wire v_26955;
wire v_26956;
wire v_26957;
wire v_26958;
wire v_26959;
wire v_26960;
wire v_26961;
wire v_26962;
wire v_26963;
wire v_26964;
wire v_26965;
wire v_26966;
wire v_26967;
wire v_26968;
wire v_26969;
wire v_26970;
wire v_26971;
wire v_26972;
wire v_26973;
wire v_26974;
wire v_26975;
wire v_26976;
wire v_26977;
wire v_26978;
wire v_26979;
wire v_26980;
wire v_26981;
wire v_26982;
wire v_26983;
wire v_26984;
wire v_26985;
wire v_26986;
wire v_26987;
wire v_26988;
wire v_26989;
wire v_26990;
wire v_26991;
wire v_26992;
wire v_26993;
wire v_26994;
wire v_26995;
wire v_26996;
wire v_26997;
wire v_26998;
wire v_26999;
wire v_27000;
wire v_27001;
wire v_27002;
wire v_27003;
wire v_27004;
wire v_27005;
wire v_27006;
wire v_27007;
wire v_27008;
wire v_27009;
wire v_27010;
wire v_27011;
wire v_27012;
wire v_27013;
wire v_27014;
wire v_27015;
wire v_27016;
wire v_27017;
wire v_27018;
wire v_27019;
wire v_27020;
wire v_27021;
wire v_27022;
wire v_27023;
wire v_27024;
wire v_27025;
wire v_27026;
wire v_27027;
wire v_27028;
wire v_27029;
wire v_27030;
wire v_27031;
wire v_27032;
wire v_27033;
wire v_27034;
wire v_27035;
wire v_27036;
wire v_27037;
wire v_27038;
wire v_27039;
wire v_27040;
wire v_27041;
wire v_27042;
wire v_27043;
wire v_27044;
wire v_27045;
wire v_27046;
wire v_27047;
wire v_27048;
wire v_27049;
wire v_27050;
wire v_27051;
wire v_27052;
wire v_27053;
wire v_27054;
wire v_27055;
wire v_27056;
wire v_27057;
wire v_27058;
wire v_27059;
wire v_27060;
wire v_27061;
wire v_27062;
wire v_27063;
wire v_27064;
wire v_27065;
wire v_27066;
wire v_27067;
wire v_27068;
wire v_27069;
wire v_27070;
wire v_27071;
wire v_27072;
wire v_27073;
wire v_27074;
wire v_27075;
wire v_27076;
wire v_27077;
wire v_27078;
wire v_27079;
wire v_27080;
wire v_27081;
wire v_27082;
wire v_27083;
wire v_27084;
wire v_27085;
wire v_27086;
wire v_27087;
wire v_27088;
wire v_27089;
wire v_27090;
wire v_27091;
wire v_27092;
wire v_27093;
wire v_27094;
wire v_27095;
wire v_27096;
wire v_27097;
wire v_27098;
wire v_27099;
wire v_27100;
wire v_27101;
wire v_27102;
wire v_27103;
wire v_27104;
wire v_27105;
wire v_27106;
wire v_27107;
wire v_27108;
wire v_27109;
wire v_27110;
wire v_27111;
wire v_27112;
wire v_27113;
wire v_27114;
wire v_27115;
wire v_27116;
wire v_27117;
wire v_27118;
wire v_27119;
wire v_27120;
wire v_27121;
wire v_27122;
wire v_27123;
wire v_27124;
wire v_27125;
wire v_27126;
wire v_27127;
wire v_27128;
wire v_27129;
wire v_27130;
wire v_27131;
wire v_27132;
wire v_27133;
wire v_27134;
wire v_27135;
wire v_27136;
wire v_27137;
wire v_27138;
wire v_27139;
wire v_27140;
wire v_27141;
wire v_27142;
wire v_27143;
wire v_27144;
wire v_27145;
wire v_27146;
wire v_27147;
wire v_27148;
wire v_27149;
wire v_27150;
wire v_27151;
wire v_27152;
wire v_27153;
wire v_27154;
wire v_27155;
wire v_27156;
wire v_27157;
wire v_27158;
wire v_27159;
wire v_27160;
wire v_27161;
wire v_27162;
wire v_27163;
wire v_27164;
wire v_27165;
wire v_27166;
wire v_27167;
wire v_27168;
wire v_27169;
wire v_27170;
wire v_27171;
wire v_27172;
wire v_27173;
wire v_27174;
wire v_27175;
wire v_27176;
wire v_27177;
wire v_27178;
wire v_27179;
wire v_27180;
wire v_27181;
wire v_27182;
wire v_27183;
wire v_27184;
wire v_27185;
wire v_27186;
wire v_27187;
wire v_27188;
wire v_27189;
wire v_27190;
wire v_27191;
wire v_27192;
wire v_27193;
wire v_27194;
wire v_27195;
wire v_27196;
wire v_27197;
wire v_27198;
wire v_27199;
wire v_27200;
wire v_27201;
wire v_27202;
wire v_27203;
wire v_27204;
wire v_27205;
wire v_27206;
wire v_27207;
wire v_27208;
wire v_27209;
wire v_27210;
wire v_27211;
wire v_27212;
wire v_27213;
wire v_27214;
wire v_27215;
wire v_27216;
wire v_27217;
wire v_27218;
wire v_27219;
wire v_27220;
wire v_27221;
wire v_27222;
wire v_27223;
wire v_27224;
wire v_27225;
wire v_27226;
wire v_27227;
wire v_27228;
wire v_27229;
wire v_27230;
wire v_27231;
wire v_27232;
wire v_27233;
wire v_27234;
wire v_27235;
wire v_27236;
wire v_27237;
wire v_27238;
wire v_27239;
wire v_27240;
wire v_27241;
wire v_27242;
wire v_27243;
wire v_27244;
wire v_27245;
wire v_27246;
wire v_27247;
wire v_27248;
wire v_27249;
wire v_27250;
wire v_27251;
wire v_27252;
wire v_27253;
wire v_27254;
wire v_27255;
wire v_27256;
wire v_27257;
wire v_27258;
wire v_27259;
wire v_27260;
wire v_27261;
wire v_27262;
wire v_27263;
wire v_27264;
wire v_27265;
wire v_27266;
wire v_27267;
wire v_27268;
wire v_27269;
wire v_27270;
wire v_27271;
wire v_27272;
wire v_27273;
wire v_27274;
wire v_27275;
wire v_27276;
wire v_27277;
wire v_27278;
wire v_27279;
wire v_27280;
wire v_27281;
wire v_27282;
wire v_27283;
wire v_27284;
wire v_27285;
wire v_27286;
wire v_27287;
wire v_27288;
wire v_27289;
wire v_27290;
wire v_27291;
wire v_27292;
wire v_27293;
wire v_27294;
wire v_27295;
wire v_27296;
wire v_27297;
wire v_27298;
wire v_27299;
wire v_27300;
wire v_27301;
wire v_27302;
wire v_27303;
wire v_27304;
wire v_27305;
wire v_27306;
wire v_27307;
wire v_27308;
wire v_27309;
wire v_27310;
wire v_27311;
wire v_27312;
wire v_27313;
wire v_27314;
wire v_27315;
wire v_27316;
wire v_27317;
wire v_27318;
wire v_27319;
wire v_27320;
wire v_27321;
wire v_27322;
wire v_27323;
wire v_27324;
wire v_27325;
wire v_27326;
wire v_27327;
wire v_27328;
wire v_27329;
wire v_27330;
wire v_27331;
wire v_27332;
wire v_27333;
wire v_27334;
wire v_27335;
wire v_27336;
wire v_27337;
wire v_27338;
wire v_27339;
wire v_27340;
wire v_27341;
wire v_27342;
wire v_27343;
wire v_27344;
wire v_27345;
wire v_27346;
wire v_27347;
wire v_27348;
wire v_27349;
wire v_27350;
wire v_27351;
wire v_27352;
wire v_27353;
wire v_27354;
wire v_27355;
wire v_27356;
wire v_27357;
wire v_27358;
wire v_27359;
wire v_27360;
wire v_27361;
wire v_27362;
wire v_27363;
wire v_27364;
wire v_27365;
wire v_27366;
wire v_27367;
wire v_27368;
wire v_27369;
wire v_27370;
wire v_27371;
wire v_27372;
wire v_27373;
wire v_27374;
wire v_27375;
wire v_27376;
wire v_27377;
wire v_27378;
wire v_27379;
wire v_27380;
wire v_27381;
wire v_27382;
wire v_27383;
wire v_27384;
wire v_27385;
wire v_27386;
wire v_27387;
wire v_27388;
wire v_27389;
wire v_27390;
wire v_27391;
wire v_27392;
wire v_27393;
wire v_27394;
wire v_27395;
wire v_27396;
wire v_27397;
wire v_27398;
wire v_27399;
wire v_27400;
wire v_27401;
wire v_27402;
wire v_27403;
wire v_27404;
wire v_27405;
wire v_27406;
wire v_27407;
wire v_27408;
wire v_27409;
wire v_27410;
wire v_27411;
wire v_27412;
wire v_27413;
wire v_27414;
wire v_27415;
wire v_27416;
wire v_27417;
wire v_27418;
wire v_27419;
wire v_27420;
wire v_27421;
wire v_27422;
wire v_27423;
wire v_27424;
wire v_27425;
wire v_27426;
wire v_27427;
wire v_27428;
wire v_27429;
wire v_27430;
wire v_27431;
wire v_27432;
wire v_27433;
wire v_27434;
wire v_27435;
wire v_27436;
wire v_27437;
wire v_27438;
wire v_27439;
wire v_27440;
wire v_27441;
wire v_27442;
wire v_27443;
wire v_27444;
wire v_27445;
wire v_27446;
wire v_27447;
wire v_27448;
wire v_27449;
wire v_27450;
wire v_27451;
wire v_27452;
wire v_27453;
wire v_27454;
wire v_27455;
wire v_27456;
wire v_27457;
wire v_27458;
wire v_27459;
wire v_27460;
wire v_27461;
wire v_27462;
wire v_27463;
wire v_27464;
wire v_27465;
wire v_27466;
wire v_27467;
wire v_27468;
wire v_27469;
wire v_27470;
wire v_27471;
wire v_27472;
wire v_27473;
wire v_27474;
wire v_27475;
wire v_27476;
wire v_27477;
wire v_27478;
wire v_27479;
wire v_27480;
wire v_27481;
wire v_27482;
wire v_27483;
wire v_27484;
wire v_27485;
wire v_27486;
wire v_27487;
wire v_27488;
wire v_27489;
wire v_27490;
wire v_27491;
wire v_27492;
wire v_27493;
wire v_27494;
wire v_27495;
wire v_27496;
wire v_27497;
wire v_27498;
wire v_27499;
wire v_27500;
wire v_27501;
wire v_27502;
wire v_27503;
wire v_27504;
wire v_27505;
wire v_27506;
wire v_27507;
wire v_27508;
wire v_27509;
wire v_27510;
wire v_27511;
wire v_27512;
wire v_27513;
wire v_27514;
wire v_27515;
wire v_27516;
wire v_27517;
wire v_27518;
wire v_27519;
wire v_27520;
wire v_27521;
wire v_27522;
wire v_27523;
wire v_27524;
wire v_27525;
wire v_27526;
wire v_27527;
wire v_27528;
wire v_27529;
wire v_27530;
wire v_27531;
wire v_27532;
wire v_27533;
wire v_27534;
wire v_27535;
wire v_27536;
wire v_27537;
wire v_27538;
wire v_27539;
wire v_27540;
wire v_27541;
wire v_27542;
wire v_27543;
wire v_27544;
wire v_27545;
wire v_27546;
wire v_27547;
wire v_27548;
wire v_27549;
wire v_27550;
wire v_27551;
wire v_27552;
wire v_27553;
wire v_27554;
wire v_27555;
wire v_27556;
wire v_27557;
wire v_27558;
wire v_27559;
wire v_27560;
wire v_27561;
wire v_27562;
wire v_27563;
wire v_27564;
wire v_27565;
wire v_27566;
wire v_27567;
wire v_27568;
wire v_27569;
wire v_27570;
wire v_27571;
wire v_27572;
wire v_27573;
wire v_27574;
wire v_27575;
wire v_27576;
wire v_27577;
wire v_27578;
wire v_27579;
wire v_27580;
wire v_27581;
wire v_27582;
wire v_27583;
wire v_27584;
wire v_27585;
wire v_27586;
wire v_27587;
wire v_27588;
wire v_27589;
wire v_27590;
wire v_27591;
wire v_27592;
wire v_27593;
wire v_27594;
wire v_27595;
wire v_27596;
wire v_27597;
wire v_27598;
wire v_27599;
wire v_27600;
wire v_27601;
wire v_27602;
wire v_27603;
wire v_27604;
wire v_27605;
wire v_27606;
wire v_27607;
wire v_27608;
wire v_27609;
wire v_27610;
wire v_27611;
wire v_27612;
wire v_27613;
wire v_27614;
wire v_27615;
wire v_27616;
wire v_27617;
wire v_27618;
wire v_27619;
wire v_27620;
wire v_27621;
wire v_27622;
wire v_27623;
wire v_27624;
wire v_27625;
wire v_27626;
wire v_27627;
wire v_27628;
wire v_27629;
wire v_27630;
wire v_27631;
wire v_27632;
wire v_27633;
wire v_27634;
wire v_27635;
wire v_27636;
wire v_27637;
wire v_27638;
wire v_27639;
wire v_27640;
wire v_27641;
wire v_27642;
wire v_27643;
wire v_27644;
wire v_27645;
wire v_27646;
wire v_27647;
wire v_27648;
wire v_27649;
wire v_27650;
wire v_27651;
wire v_27652;
wire v_27653;
wire v_27654;
wire v_27655;
wire v_27656;
wire v_27657;
wire v_27658;
wire v_27659;
wire v_27660;
wire v_27661;
wire v_27662;
wire v_27663;
wire v_27664;
wire v_27665;
wire v_27666;
wire v_27667;
wire v_27668;
wire v_27669;
wire v_27670;
wire v_27671;
wire v_27672;
wire v_27673;
wire v_27674;
wire v_27675;
wire v_27676;
wire v_27677;
wire v_27678;
wire v_27679;
wire v_27680;
wire v_27681;
wire v_27682;
wire v_27683;
wire v_27684;
wire v_27685;
wire v_27686;
wire v_27687;
wire v_27688;
wire v_27689;
wire v_27690;
wire v_27691;
wire v_27692;
wire v_27693;
wire v_27694;
wire v_27695;
wire v_27696;
wire v_27697;
wire v_27698;
wire v_27699;
wire v_27700;
wire v_27701;
wire v_27702;
wire v_27703;
wire v_27704;
wire v_27705;
wire v_27706;
wire v_27707;
wire v_27708;
wire v_27709;
wire v_27710;
wire v_27711;
wire v_27712;
wire v_27713;
wire v_27714;
wire v_27715;
wire v_27716;
wire v_27717;
wire v_27718;
wire v_27719;
wire v_27720;
wire v_27721;
wire v_27722;
wire v_27723;
wire v_27724;
wire v_27725;
wire v_27726;
wire v_27727;
wire v_27728;
wire v_27729;
wire v_27730;
wire v_27731;
wire v_27732;
wire v_27733;
wire v_27734;
wire v_27735;
wire v_27736;
wire v_27737;
wire v_27738;
wire v_27739;
wire v_27740;
wire v_27741;
wire v_27742;
wire v_27743;
wire v_27744;
wire v_27745;
wire v_27746;
wire v_27747;
wire v_27748;
wire v_27749;
wire v_27750;
wire v_27751;
wire v_27752;
wire v_27753;
wire v_27754;
wire v_27755;
wire v_27756;
wire v_27757;
wire v_27758;
wire v_27759;
wire v_27760;
wire v_27761;
wire v_27762;
wire v_27763;
wire v_27764;
wire v_27765;
wire v_27766;
wire v_27767;
wire v_27768;
wire v_27769;
wire v_27770;
wire v_27771;
wire v_27772;
wire v_27773;
wire v_27774;
wire v_27775;
wire v_27776;
wire v_27777;
wire v_27778;
wire v_27779;
wire v_27780;
wire v_27781;
wire v_27782;
wire v_27783;
wire v_27784;
wire v_27785;
wire v_27786;
wire v_27787;
wire v_27788;
wire v_27789;
wire v_27790;
wire v_27791;
wire v_27792;
wire v_27793;
wire v_27794;
wire v_27795;
wire v_27796;
wire v_27797;
wire v_27798;
wire v_27799;
wire v_27800;
wire v_27801;
wire v_27802;
wire v_27803;
wire v_27804;
wire v_27805;
wire v_27806;
wire v_27807;
wire v_27808;
wire v_27809;
wire v_27810;
wire v_27811;
wire v_27812;
wire v_27813;
wire v_27814;
wire v_27815;
wire v_27816;
wire v_27817;
wire v_27818;
wire v_27819;
wire v_27820;
wire v_27821;
wire v_27822;
wire v_27823;
wire v_27824;
wire v_27825;
wire v_27826;
wire v_27827;
wire v_27828;
wire v_27829;
wire v_27830;
wire v_27831;
wire v_27832;
wire v_27833;
wire v_27834;
wire v_27835;
wire v_27836;
wire v_27837;
wire v_27838;
wire v_27839;
wire v_27840;
wire v_27841;
wire v_27842;
wire v_27843;
wire v_27844;
wire v_27845;
wire v_27846;
wire v_27847;
wire v_27848;
wire v_27849;
wire v_27850;
wire v_27851;
wire v_27852;
wire v_27853;
wire v_27854;
wire v_27855;
wire v_27856;
wire v_27857;
wire v_27858;
wire v_27859;
wire v_27860;
wire v_27861;
wire v_27862;
wire v_27863;
wire v_27864;
wire v_27865;
wire v_27866;
wire v_27867;
wire v_27868;
wire v_27869;
wire v_27870;
wire v_27871;
wire v_27872;
wire v_27873;
wire v_27874;
wire v_27875;
wire v_27876;
wire v_27877;
wire v_27878;
wire v_27879;
wire v_27880;
wire v_27881;
wire v_27882;
wire v_27883;
wire v_27884;
wire v_27885;
wire v_27886;
wire v_27887;
wire v_27888;
wire v_27889;
wire v_27890;
wire v_27891;
wire v_27892;
wire v_27893;
wire v_27894;
wire v_27895;
wire v_27896;
wire v_27897;
wire v_27898;
wire v_27899;
wire v_27900;
wire v_27901;
wire v_27902;
wire v_27903;
wire v_27904;
wire v_27905;
wire v_27906;
wire v_27907;
wire v_27908;
wire v_27909;
wire v_27910;
wire v_27911;
wire v_27912;
wire v_27913;
wire v_27914;
wire v_27915;
wire v_27916;
wire v_27917;
wire v_27918;
wire v_27919;
wire v_27920;
wire v_27921;
wire v_27922;
wire v_27923;
wire v_27924;
wire v_27925;
wire v_27926;
wire v_27927;
wire v_27928;
wire v_27929;
wire v_27930;
wire v_27931;
wire v_27932;
wire v_27933;
wire v_27934;
wire v_27935;
wire v_27936;
wire v_27937;
wire v_27938;
wire v_27939;
wire v_27940;
wire v_27941;
wire v_27942;
wire v_27943;
wire v_27944;
wire v_27945;
wire v_27946;
wire v_27947;
wire v_27948;
wire v_27949;
wire v_27950;
wire v_27951;
wire v_27952;
wire v_27953;
wire v_27954;
wire v_27955;
wire v_27956;
wire v_27957;
wire v_27958;
wire v_27959;
wire v_27960;
wire v_27961;
wire v_27962;
wire v_27963;
wire v_27964;
wire v_27965;
wire v_27966;
wire v_27967;
wire v_27968;
wire v_27969;
wire v_27970;
wire v_27971;
wire v_27972;
wire v_27973;
wire v_27974;
wire v_27975;
wire v_27976;
wire v_27977;
wire v_27978;
wire v_27979;
wire v_27980;
wire v_27981;
wire v_27982;
wire v_27983;
wire v_27984;
wire v_27985;
wire v_27986;
wire v_27987;
wire v_27988;
wire v_27989;
wire v_27990;
wire v_27991;
wire v_27992;
wire v_27993;
wire v_27994;
wire v_27995;
wire v_27996;
wire v_27997;
wire v_27998;
wire v_27999;
wire v_28000;
wire v_28001;
wire v_28002;
wire v_28003;
wire v_28004;
wire v_28005;
wire v_28006;
wire v_28007;
wire v_28008;
wire v_28009;
wire v_28010;
wire v_28011;
wire v_28012;
wire v_28013;
wire v_28014;
wire v_28015;
wire v_28016;
wire v_28017;
wire v_28018;
wire v_28019;
wire v_28020;
wire v_28021;
wire v_28022;
wire v_28023;
wire v_28024;
wire v_28025;
wire v_28026;
wire v_28027;
wire v_28028;
wire v_28029;
wire v_28030;
wire v_28031;
wire v_28032;
wire v_28033;
wire v_28034;
wire v_28035;
wire v_28036;
wire v_28037;
wire v_28038;
wire v_28039;
wire v_28040;
wire v_28041;
wire v_28042;
wire v_28043;
wire v_28044;
wire v_28045;
wire v_28046;
wire v_28047;
wire v_28048;
wire v_28049;
wire v_28050;
wire v_28051;
wire v_28052;
wire v_28053;
wire v_28054;
wire v_28055;
wire v_28056;
wire v_28057;
wire v_28058;
wire v_28059;
wire v_28060;
wire v_28061;
wire v_28062;
wire v_28063;
wire v_28064;
wire v_28065;
wire v_28066;
wire v_28067;
wire v_28068;
wire v_28069;
wire v_28070;
wire v_28071;
wire v_28072;
wire v_28073;
wire v_28074;
wire v_28075;
wire v_28076;
wire v_28077;
wire v_28078;
wire v_28079;
wire v_28080;
wire v_28081;
wire v_28082;
wire v_28083;
wire v_28084;
wire v_28085;
wire v_28086;
wire v_28087;
wire v_28088;
wire v_28089;
wire v_28090;
wire v_28091;
wire v_28092;
wire v_28093;
wire v_28094;
wire v_28095;
wire v_28096;
wire v_28097;
wire v_28098;
wire v_28099;
wire v_28100;
wire v_28101;
wire v_28102;
wire v_28103;
wire v_28104;
wire v_28105;
wire v_28106;
wire v_28107;
wire v_28108;
wire v_28109;
wire v_28110;
wire v_28111;
wire v_28112;
wire v_28113;
wire v_28114;
wire v_28115;
wire v_28116;
wire v_28117;
wire v_28118;
wire v_28119;
wire v_28120;
wire v_28121;
wire v_28122;
wire v_28123;
wire v_28124;
wire v_28125;
wire v_28126;
wire v_28127;
wire v_28128;
wire v_28129;
wire v_28130;
wire v_28131;
wire v_28132;
wire v_28133;
wire v_28134;
wire v_28135;
wire v_28136;
wire v_28137;
wire v_28138;
wire v_28139;
wire v_28140;
wire v_28141;
wire v_28142;
wire v_28143;
wire v_28144;
wire v_28145;
wire v_28146;
wire v_28147;
wire v_28148;
wire v_28149;
wire v_28150;
wire v_28151;
wire v_28152;
wire v_28153;
wire v_28154;
wire v_28155;
wire v_28156;
wire v_28157;
wire v_28158;
wire v_28159;
wire v_28160;
wire v_28161;
wire v_28162;
wire v_28163;
wire v_28164;
wire v_28165;
wire v_28166;
wire v_28167;
wire v_28168;
wire v_28169;
wire v_28170;
wire v_28171;
wire v_28172;
wire v_28173;
wire v_28174;
wire v_28175;
wire v_28176;
wire v_28177;
wire v_28178;
wire v_28179;
wire v_28180;
wire v_28181;
wire v_28182;
wire v_28183;
wire v_28184;
wire v_28185;
wire v_28186;
wire v_28187;
wire v_28188;
wire v_28189;
wire v_28190;
wire v_28191;
wire v_28192;
wire v_28193;
wire v_28194;
wire v_28195;
wire v_28196;
wire v_28197;
wire v_28198;
wire v_28199;
wire v_28200;
wire v_28201;
wire v_28202;
wire v_28203;
wire v_28204;
wire v_28205;
wire v_28206;
wire v_28207;
wire v_28208;
wire v_28209;
wire v_28210;
wire v_28211;
wire v_28212;
wire v_28213;
wire v_28214;
wire v_28215;
wire v_28216;
wire v_28217;
wire v_28218;
wire v_28219;
wire v_28220;
wire v_28221;
wire v_28222;
wire v_28223;
wire v_28224;
wire v_28225;
wire v_28226;
wire v_28227;
wire v_28228;
wire v_28229;
wire v_28230;
wire v_28231;
wire v_28232;
wire v_28233;
wire v_28234;
wire v_28235;
wire v_28236;
wire v_28237;
wire v_28238;
wire v_28239;
wire v_28240;
wire v_28241;
wire v_28242;
wire v_28243;
wire v_28244;
wire v_28245;
wire v_28246;
wire v_28247;
wire v_28248;
wire v_28249;
wire v_28250;
wire v_28251;
wire v_28252;
wire v_28253;
wire v_28254;
wire v_28255;
wire v_28256;
wire v_28257;
wire v_28258;
wire v_28259;
wire v_28260;
wire v_28261;
wire v_28262;
wire v_28263;
wire v_28264;
wire v_28265;
wire v_28266;
wire v_28267;
wire v_28268;
wire v_28269;
wire v_28270;
wire v_28271;
wire v_28272;
wire v_28273;
wire v_28274;
wire v_28275;
wire v_28276;
wire v_28277;
wire v_28278;
wire v_28279;
wire v_28280;
wire v_28281;
wire v_28282;
wire v_28283;
wire v_28284;
wire v_28285;
wire v_28286;
wire v_28287;
wire v_28288;
wire v_28289;
wire v_28290;
wire v_28291;
wire v_28292;
wire v_28293;
wire v_28294;
wire v_28295;
wire v_28296;
wire v_28297;
wire v_28298;
wire v_28299;
wire v_28300;
wire v_28301;
wire v_28302;
wire v_28303;
wire v_28304;
wire v_28305;
wire v_28306;
wire v_28307;
wire v_28308;
wire v_28309;
wire v_28310;
wire v_28311;
wire v_28312;
wire v_28313;
wire v_28314;
wire v_28315;
wire v_28316;
wire v_28317;
wire v_28318;
wire v_28319;
wire v_28320;
wire v_28321;
wire v_28322;
wire v_28323;
wire v_28324;
wire v_28325;
wire v_28326;
wire v_28327;
wire v_28328;
wire v_28329;
wire v_28330;
wire v_28331;
wire v_28332;
wire v_28333;
wire v_28334;
wire v_28335;
wire v_28336;
wire v_28337;
wire v_28338;
wire v_28339;
wire v_28340;
wire v_28341;
wire v_28342;
wire v_28343;
wire v_28344;
wire v_28345;
wire v_28346;
wire v_28347;
wire v_28348;
wire v_28349;
wire v_28350;
wire v_28351;
wire v_28352;
wire v_28353;
wire v_28354;
wire v_28355;
wire v_28356;
wire v_28357;
wire v_28358;
wire v_28359;
wire v_28360;
wire v_28361;
wire v_28362;
wire v_28363;
wire v_28364;
wire v_28365;
wire v_28366;
wire v_28367;
wire v_28368;
wire v_28369;
wire v_28370;
wire v_28371;
wire v_28372;
wire v_28373;
wire v_28374;
wire v_28375;
wire v_28376;
wire v_28377;
wire v_28378;
wire v_28379;
wire v_28380;
wire v_28381;
wire v_28382;
wire v_28383;
wire v_28384;
wire v_28385;
wire v_28386;
wire v_28387;
wire v_28388;
wire v_28389;
wire v_28390;
wire v_28391;
wire v_28392;
wire v_28393;
wire v_28394;
wire v_28395;
wire v_28396;
wire v_28397;
wire v_28398;
wire v_28399;
wire v_28400;
wire v_28401;
wire v_28402;
wire v_28403;
wire v_28404;
wire v_28405;
wire v_28406;
wire v_28407;
wire v_28408;
wire v_28409;
wire v_28410;
wire v_28411;
wire v_28412;
wire v_28413;
wire v_28414;
wire v_28415;
wire v_28416;
wire v_28417;
wire v_28418;
wire v_28419;
wire v_28420;
wire v_28421;
wire v_28422;
wire v_28423;
wire v_28424;
wire v_28425;
wire v_28426;
wire v_28427;
wire v_28428;
wire v_28429;
wire v_28430;
wire v_28431;
wire v_28432;
wire v_28433;
wire v_28434;
wire v_28435;
wire v_28436;
wire v_28437;
wire v_28438;
wire v_28439;
wire v_28440;
wire v_28441;
wire v_28442;
wire v_28443;
wire v_28444;
wire v_28445;
wire v_28446;
wire v_28447;
wire v_28448;
wire v_28449;
wire v_28450;
wire v_28451;
wire v_28452;
wire v_28453;
wire v_28454;
wire v_28455;
wire v_28456;
wire v_28457;
wire v_28458;
wire v_28459;
wire v_28460;
wire v_28461;
wire v_28462;
wire v_28463;
wire v_28464;
wire v_28465;
wire v_28466;
wire v_28467;
wire v_28468;
wire v_28469;
wire v_28470;
wire v_28471;
wire v_28472;
wire v_28473;
wire v_28474;
wire v_28475;
wire v_28476;
wire v_28477;
wire v_28478;
wire v_28479;
wire v_28480;
wire v_28481;
wire v_28482;
wire v_28483;
wire v_28484;
wire v_28485;
wire v_28486;
wire v_28487;
wire v_28488;
wire v_28489;
wire v_28490;
wire v_28491;
wire v_28492;
wire v_28493;
wire v_28494;
wire v_28495;
wire v_28496;
wire v_28497;
wire v_28498;
wire v_28499;
wire v_28500;
wire v_28501;
wire v_28502;
wire v_28503;
wire v_28504;
wire v_28505;
wire v_28506;
wire v_28507;
wire v_28508;
wire v_28509;
wire v_28510;
wire v_28511;
wire v_28512;
wire v_28513;
wire v_28514;
wire v_28515;
wire v_28516;
wire v_28517;
wire v_28518;
wire v_28519;
wire v_28520;
wire v_28521;
wire v_28522;
wire v_28523;
wire v_28524;
wire v_28525;
wire v_28526;
wire v_28527;
wire v_28528;
wire v_28529;
wire v_28530;
wire v_28531;
wire v_28532;
wire v_28533;
wire v_28534;
wire v_28535;
wire v_28536;
wire v_28537;
wire v_28538;
wire v_28539;
wire v_28540;
wire v_28541;
wire v_28542;
wire v_28543;
wire v_28544;
wire v_28545;
wire v_28546;
wire v_28547;
wire v_28548;
wire v_28549;
wire v_28550;
wire v_28551;
wire v_28552;
wire v_28553;
wire v_28554;
wire v_28555;
wire v_28556;
wire v_28557;
wire v_28558;
wire v_28559;
wire v_28560;
wire v_28561;
wire v_28562;
wire v_28563;
wire v_28564;
wire v_28565;
wire v_28566;
wire v_28567;
wire v_28568;
wire v_28569;
wire v_28570;
wire v_28571;
wire v_28572;
wire v_28573;
wire v_28574;
wire v_28575;
wire v_28576;
wire v_28577;
wire v_28578;
wire v_28579;
wire v_28580;
wire v_28581;
wire v_28582;
wire v_28583;
wire v_28584;
wire v_28585;
wire v_28586;
wire v_28587;
wire v_28588;
wire v_28589;
wire v_28590;
wire v_28591;
wire v_28592;
wire v_28593;
wire v_28594;
wire v_28595;
wire v_28596;
wire v_28597;
wire v_28598;
wire v_28599;
wire v_28600;
wire v_28601;
wire v_28602;
wire v_28603;
wire v_28604;
wire v_28605;
wire v_28606;
wire v_28607;
wire v_28608;
wire v_28609;
wire v_28610;
wire v_28611;
wire v_28612;
wire v_28613;
wire v_28614;
wire v_28615;
wire v_28616;
wire v_28617;
wire v_28618;
wire v_28619;
wire v_28620;
wire v_28621;
wire v_28622;
wire v_28623;
wire v_28624;
wire v_28625;
wire v_28626;
wire v_28627;
wire v_28628;
wire v_28629;
wire v_28630;
wire v_28631;
wire v_28632;
wire v_28633;
wire v_28634;
wire v_28635;
wire v_28636;
wire v_28637;
wire v_28638;
wire v_28639;
wire v_28640;
wire v_28641;
wire v_28642;
wire v_28643;
wire v_28644;
wire v_28645;
wire v_28646;
wire v_28647;
wire v_28648;
wire v_28649;
wire v_28650;
wire v_28651;
wire v_28652;
wire v_28653;
wire v_28654;
wire v_28655;
wire v_28656;
wire v_28657;
wire v_28658;
wire v_28659;
wire v_28660;
wire v_28661;
wire v_28662;
wire v_28663;
wire v_28664;
wire v_28665;
wire v_28666;
wire v_28667;
wire v_28668;
wire v_28669;
wire v_28670;
wire v_28671;
wire v_28672;
wire v_28673;
wire v_28674;
wire v_28675;
wire v_28676;
wire v_28677;
wire v_28678;
wire v_28679;
wire v_28680;
wire v_28681;
wire v_28682;
wire v_28683;
wire v_28684;
wire v_28685;
wire v_28686;
wire v_28687;
wire v_28688;
wire v_28689;
wire v_28690;
wire v_28691;
wire v_28692;
wire v_28693;
wire v_28694;
wire v_28695;
wire v_28696;
wire v_28697;
wire v_28698;
wire v_28699;
wire v_28700;
wire v_28701;
wire v_28702;
wire v_28703;
wire v_28704;
wire v_28705;
wire v_28706;
wire v_28707;
wire v_28708;
wire v_28709;
wire v_28710;
wire v_28711;
wire v_28712;
wire v_28713;
wire v_28714;
wire v_28715;
wire v_28716;
wire v_28717;
wire v_28718;
wire v_28719;
wire v_28720;
wire v_28721;
wire v_28722;
wire v_28723;
wire v_28724;
wire v_28725;
wire v_28726;
wire v_28727;
wire v_28728;
wire v_28729;
wire v_28730;
wire v_28731;
wire v_28732;
wire v_28733;
wire v_28734;
wire v_28735;
wire v_28736;
wire v_28737;
wire v_28738;
wire v_28739;
wire v_28740;
wire v_28741;
wire v_28742;
wire v_28743;
wire v_28744;
wire v_28745;
wire v_28746;
wire v_28747;
wire v_28748;
wire v_28749;
wire v_28750;
wire v_28751;
wire v_28752;
wire v_28753;
wire v_28754;
wire v_28755;
wire v_28756;
wire v_28757;
wire v_28758;
wire v_28759;
wire v_28760;
wire v_28761;
wire v_28762;
wire v_28763;
wire v_28764;
wire v_28765;
wire v_28766;
wire v_28767;
wire v_28768;
wire v_28769;
wire v_28770;
wire v_28771;
wire v_28772;
wire v_28773;
wire v_28774;
wire v_28775;
wire v_28776;
wire v_28777;
wire v_28778;
wire v_28779;
wire v_28780;
wire v_28781;
wire v_28782;
wire v_28783;
wire v_28784;
wire v_28785;
wire v_28786;
wire v_28787;
wire v_28788;
wire v_28789;
wire v_28790;
wire v_28791;
wire v_28792;
wire v_28793;
wire v_28794;
wire v_28795;
wire v_28796;
wire v_28797;
wire v_28798;
wire v_28799;
wire v_28800;
wire v_28801;
wire v_28802;
wire v_28803;
wire v_28804;
wire v_28805;
wire v_28806;
wire v_28807;
wire v_28808;
wire v_28809;
wire v_28810;
wire v_28811;
wire v_28812;
wire v_28813;
wire v_28814;
wire v_28815;
wire v_28816;
wire v_28817;
wire v_28818;
wire v_28819;
wire v_28820;
wire v_28821;
wire v_28822;
wire v_28823;
wire v_28824;
wire v_28825;
wire v_28826;
wire v_28827;
wire v_28828;
wire v_28829;
wire v_28830;
wire v_28831;
wire v_28832;
wire v_28833;
wire v_28834;
wire v_28835;
wire v_28836;
wire v_28837;
wire v_28838;
wire v_28839;
wire v_28840;
wire v_28841;
wire v_28842;
wire v_28843;
wire v_28844;
wire v_28845;
wire v_28846;
wire v_28847;
wire v_28848;
wire v_28849;
wire v_28850;
wire v_28851;
wire v_28852;
wire v_28853;
wire v_28854;
wire v_28855;
wire v_28856;
wire v_28857;
wire v_28858;
wire v_28859;
wire v_28860;
wire v_28861;
wire v_28862;
wire v_28863;
wire v_28864;
wire v_28865;
wire v_28866;
wire v_28867;
wire v_28868;
wire v_28869;
wire v_28870;
wire v_28871;
wire v_28872;
wire v_28873;
wire v_28874;
wire v_28875;
wire v_28876;
wire v_28877;
wire v_28878;
wire v_28879;
wire v_28880;
wire v_28881;
wire v_28882;
wire v_28883;
wire v_28884;
wire v_28885;
wire v_28886;
wire v_28887;
wire v_28888;
wire v_28889;
wire v_28890;
wire v_28891;
wire v_28892;
wire v_28893;
wire v_28894;
wire v_28895;
wire v_28896;
wire v_28897;
wire v_28898;
wire v_28899;
wire v_28900;
wire v_28901;
wire v_28902;
wire v_28903;
wire v_28904;
wire v_28905;
wire v_28906;
wire v_28907;
wire v_28908;
wire v_28909;
wire v_28910;
wire v_28911;
wire v_28912;
wire v_28913;
wire v_28914;
wire v_28915;
wire v_28916;
wire v_28917;
wire v_28918;
wire v_28919;
wire v_28920;
wire v_28921;
wire v_28922;
wire v_28923;
wire v_28924;
wire v_28925;
wire v_28926;
wire v_28927;
wire v_28928;
wire v_28929;
wire v_28930;
wire v_28931;
wire v_28932;
wire v_28933;
wire v_28934;
wire v_28935;
wire v_28936;
wire v_28937;
wire v_28938;
wire v_28939;
wire v_28940;
wire v_28941;
wire v_28942;
wire v_28943;
wire v_28944;
wire v_28945;
wire v_28946;
wire v_28947;
wire v_28948;
wire v_28949;
wire v_28950;
wire v_28951;
wire v_28952;
wire v_28953;
wire v_28954;
wire v_28955;
wire v_28956;
wire v_28957;
wire v_28958;
wire v_28959;
wire v_28960;
wire v_28961;
wire v_28962;
wire v_28963;
wire v_28964;
wire v_28965;
wire v_28966;
wire v_28967;
wire v_28968;
wire v_28969;
wire v_28970;
wire v_28971;
wire v_28972;
wire v_28973;
wire v_28974;
wire v_28975;
wire v_28976;
wire v_28977;
wire v_28978;
wire v_28979;
wire v_28980;
wire v_28981;
wire v_28982;
wire v_28983;
wire v_28984;
wire v_28985;
wire v_28986;
wire v_28987;
wire v_28988;
wire v_28989;
wire v_28990;
wire v_28991;
wire v_28992;
wire v_28993;
wire v_28994;
wire v_28995;
wire v_28996;
wire v_28997;
wire v_28998;
wire v_28999;
wire v_29000;
wire v_29001;
wire v_29002;
wire v_29003;
wire v_29004;
wire v_29005;
wire v_29006;
wire v_29007;
wire v_29008;
wire v_29009;
wire v_29010;
wire v_29011;
wire v_29012;
wire v_29013;
wire v_29014;
wire v_29015;
wire v_29016;
wire v_29017;
wire v_29018;
wire v_29019;
wire v_29020;
wire v_29021;
wire v_29022;
wire v_29023;
wire v_29024;
wire v_29025;
wire v_29026;
wire v_29027;
wire v_29028;
wire v_29029;
wire v_29030;
wire v_29031;
wire v_29032;
wire v_29033;
wire v_29034;
wire v_29035;
wire v_29036;
wire v_29037;
wire v_29038;
wire v_29039;
wire v_29040;
wire v_29041;
wire v_29042;
wire v_29043;
wire v_29044;
wire v_29045;
wire v_29046;
wire v_29047;
wire v_29048;
wire v_29049;
wire v_29050;
wire v_29051;
wire v_29052;
wire v_29053;
wire v_29054;
wire v_29055;
wire v_29056;
wire v_29057;
wire v_29058;
wire v_29059;
wire v_29060;
wire v_29061;
wire v_29062;
wire v_29063;
wire v_29064;
wire v_29065;
wire v_29066;
wire v_29067;
wire v_29068;
wire v_29069;
wire v_29070;
wire v_29071;
wire v_29072;
wire v_29073;
wire v_29074;
wire v_29075;
wire v_29076;
wire v_29077;
wire v_29078;
wire v_29079;
wire v_29080;
wire v_29081;
wire v_29082;
wire v_29083;
wire v_29084;
wire v_29085;
wire v_29086;
wire v_29087;
wire v_29088;
wire v_29089;
wire v_29090;
wire v_29091;
wire v_29092;
wire v_29093;
wire v_29094;
wire v_29095;
wire v_29096;
wire v_29097;
wire v_29098;
wire v_29099;
wire v_29100;
wire v_29101;
wire v_29102;
wire v_29103;
wire v_29104;
wire v_29105;
wire v_29106;
wire v_29107;
wire v_29108;
wire v_29109;
wire v_29110;
wire v_29111;
wire v_29112;
wire v_29113;
wire v_29114;
wire v_29115;
wire v_29116;
wire v_29117;
wire v_29118;
wire v_29119;
wire v_29120;
wire v_29121;
wire v_29122;
wire v_29123;
wire v_29124;
wire v_29125;
wire v_29126;
wire v_29127;
wire v_29128;
wire v_29129;
wire v_29130;
wire v_29131;
wire v_29132;
wire v_29133;
wire v_29134;
wire v_29135;
wire v_29136;
wire v_29137;
wire v_29138;
wire v_29139;
wire v_29140;
wire v_29141;
wire v_29142;
wire v_29143;
wire v_29144;
wire v_29145;
wire v_29146;
wire v_29147;
wire v_29148;
wire v_29149;
wire v_29150;
wire v_29151;
wire v_29152;
wire v_29153;
wire v_29154;
wire v_29155;
wire v_29156;
wire v_29157;
wire v_29158;
wire v_29159;
wire v_29160;
wire v_29161;
wire v_29162;
wire v_29163;
wire v_29164;
wire v_29165;
wire v_29166;
wire v_29167;
wire v_29168;
wire v_29169;
wire v_29170;
wire v_29171;
wire v_29172;
wire v_29173;
wire v_29174;
wire v_29175;
wire v_29176;
wire v_29177;
wire v_29178;
wire v_29179;
wire v_29180;
wire v_29181;
wire v_29182;
wire v_29183;
wire v_29184;
wire v_29185;
wire v_29186;
wire v_29187;
wire v_29188;
wire v_29189;
wire v_29190;
wire v_29191;
wire v_29192;
wire v_29193;
wire v_29194;
wire v_29195;
wire v_29196;
wire v_29197;
wire v_29198;
wire v_29199;
wire v_29200;
wire v_29201;
wire v_29202;
wire v_29203;
wire v_29204;
wire v_29205;
wire v_29206;
wire v_29207;
wire v_29208;
wire v_29209;
wire v_29210;
wire v_29211;
wire v_29212;
wire v_29213;
wire v_29214;
wire v_29215;
wire v_29216;
wire v_29217;
wire v_29218;
wire v_29219;
wire v_29220;
wire v_29221;
wire v_29222;
wire v_29223;
wire v_29224;
wire v_29225;
wire v_29226;
wire v_29227;
wire v_29228;
wire v_29229;
wire v_29230;
wire v_29231;
wire v_29232;
wire v_29233;
wire v_29234;
wire v_29235;
wire v_29236;
wire v_29237;
wire v_29238;
wire v_29239;
wire v_29240;
wire v_29241;
wire v_29242;
wire v_29243;
wire v_29244;
wire v_29245;
wire v_29246;
wire v_29247;
wire v_29248;
wire v_29249;
wire v_29250;
wire v_29251;
wire v_29252;
wire v_29253;
wire v_29254;
wire v_29255;
wire v_29256;
wire v_29257;
wire v_29258;
wire v_29259;
wire v_29260;
wire v_29261;
wire v_29262;
wire v_29263;
wire v_29264;
wire v_29265;
wire v_29266;
wire v_29267;
wire v_29268;
wire v_29269;
wire v_29270;
wire v_29271;
wire v_29272;
wire v_29273;
wire v_29274;
wire v_29275;
wire v_29276;
wire v_29277;
wire v_29278;
wire v_29279;
wire v_29280;
wire v_29281;
wire v_29282;
wire v_29283;
wire v_29284;
wire v_29285;
wire v_29286;
wire v_29287;
wire v_29288;
wire v_29289;
wire v_29290;
wire v_29291;
wire v_29292;
wire v_29293;
wire v_29294;
wire v_29295;
wire v_29296;
wire v_29297;
wire v_29298;
wire v_29299;
wire v_29300;
wire v_29301;
wire v_29302;
wire v_29303;
wire v_29304;
wire v_29305;
wire v_29306;
wire v_29307;
wire v_29308;
wire v_29309;
wire v_29310;
wire v_29311;
wire v_29312;
wire v_29313;
wire v_29314;
wire v_29315;
wire v_29316;
wire v_29317;
wire v_29318;
wire v_29319;
wire v_29320;
wire v_29321;
wire v_29322;
wire v_29323;
wire v_29324;
wire v_29325;
wire v_29326;
wire v_29327;
wire v_29328;
wire v_29329;
wire v_29330;
wire v_29331;
wire v_29332;
wire v_29333;
wire v_29334;
wire v_29335;
wire v_29336;
wire v_29337;
wire v_29338;
wire v_29339;
wire v_29340;
wire v_29341;
wire v_29342;
wire v_29343;
wire v_29344;
wire v_29345;
wire v_29346;
wire v_29347;
wire v_29348;
wire v_29349;
wire v_29350;
wire v_29351;
wire v_29352;
wire v_29353;
wire v_29354;
wire v_29355;
wire v_29356;
wire v_29357;
wire v_29358;
wire v_29359;
wire v_29360;
wire v_29361;
wire v_29362;
wire v_29363;
wire v_29364;
wire v_29365;
wire v_29366;
wire v_29367;
wire v_29368;
wire v_29369;
wire v_29370;
wire v_29371;
wire v_29372;
wire v_29373;
wire v_29374;
wire v_29375;
wire v_29376;
wire v_29377;
wire v_29378;
wire v_29379;
wire v_29380;
wire v_29381;
wire v_29382;
wire v_29383;
wire v_29384;
wire v_29385;
wire v_29386;
wire v_29387;
wire v_29388;
wire v_29389;
wire v_29390;
wire v_29391;
wire v_29392;
wire v_29393;
wire v_29394;
wire v_29395;
wire v_29396;
wire v_29397;
wire v_29398;
wire v_29399;
wire v_29400;
wire v_29401;
wire v_29402;
wire v_29403;
wire v_29404;
wire v_29405;
wire v_29406;
wire v_29407;
wire v_29408;
wire v_29409;
wire v_29410;
wire v_29411;
wire v_29412;
wire v_29413;
wire v_29414;
wire v_29415;
wire v_29416;
wire v_29417;
wire v_29418;
wire v_29419;
wire v_29420;
wire v_29421;
wire v_29422;
wire v_29423;
wire v_29424;
wire v_29425;
wire v_29426;
wire v_29427;
wire v_29428;
wire v_29429;
wire v_29430;
wire v_29431;
wire v_29432;
wire v_29433;
wire v_29434;
wire v_29435;
wire v_29436;
wire v_29437;
wire v_29438;
wire v_29439;
wire v_29440;
wire v_29441;
wire v_29442;
wire v_29443;
wire v_29444;
wire v_29445;
wire v_29446;
wire v_29447;
wire v_29448;
wire v_29449;
wire v_29450;
wire v_29451;
wire v_29452;
wire v_29453;
wire v_29454;
wire v_29455;
wire v_29456;
wire v_29457;
wire v_29458;
wire v_29459;
wire v_29460;
wire v_29461;
wire v_29462;
wire v_29463;
wire v_29464;
wire v_29465;
wire v_29466;
wire v_29467;
wire v_29468;
wire v_29469;
wire v_29470;
wire v_29471;
wire v_29472;
wire v_29473;
wire v_29474;
wire v_29475;
wire v_29476;
wire v_29477;
wire v_29478;
wire v_29479;
wire v_29480;
wire v_29481;
wire v_29482;
wire v_29483;
wire v_29484;
wire v_29485;
wire v_29486;
wire v_29487;
wire v_29488;
wire v_29489;
wire v_29490;
wire v_29491;
wire v_29492;
wire v_29493;
wire v_29494;
wire v_29495;
wire v_29496;
wire v_29497;
wire v_29498;
wire v_29499;
wire v_29500;
wire v_29501;
wire v_29502;
wire v_29503;
wire v_29504;
wire v_29505;
wire v_29506;
wire v_29507;
wire v_29508;
wire v_29509;
wire v_29510;
wire v_29511;
wire v_29512;
wire v_29513;
wire v_29514;
wire v_29515;
wire v_29516;
wire v_29517;
wire v_29518;
wire v_29519;
wire v_29520;
wire v_29521;
wire v_29522;
wire v_29523;
wire v_29524;
wire v_29525;
wire v_29526;
wire v_29527;
wire v_29528;
wire v_29529;
wire v_29530;
wire v_29531;
wire v_29532;
wire v_29533;
wire v_29534;
wire v_29535;
wire v_29536;
wire v_29537;
wire v_29538;
wire v_29539;
wire v_29540;
wire v_29541;
wire v_29542;
wire v_29543;
wire v_29544;
wire v_29545;
wire v_29546;
wire v_29547;
wire v_29548;
wire v_29549;
wire v_29550;
wire v_29551;
wire v_29552;
wire v_29553;
wire v_29554;
wire v_29555;
wire v_29556;
wire v_29557;
wire v_29558;
wire v_29559;
wire v_29560;
wire v_29561;
wire v_29562;
wire v_29563;
wire v_29564;
wire v_29565;
wire v_29566;
wire v_29567;
wire v_29568;
wire v_29569;
wire v_29570;
wire v_29571;
wire v_29572;
wire v_29573;
wire v_29574;
wire v_29575;
wire v_29576;
wire v_29577;
wire v_29578;
wire v_29579;
wire v_29580;
wire v_29581;
wire v_29582;
wire v_29583;
wire v_29584;
wire v_29585;
wire v_29586;
wire v_29587;
wire v_29588;
wire v_29589;
wire v_29590;
wire v_29591;
wire v_29592;
wire v_29593;
wire v_29594;
wire v_29595;
wire v_29596;
wire v_29597;
wire v_29598;
wire v_29599;
wire v_29600;
wire v_29601;
wire v_29602;
wire v_29603;
wire v_29604;
wire v_29605;
wire v_29606;
wire v_29607;
wire v_29608;
wire v_29609;
wire v_29610;
wire v_29611;
wire v_29612;
wire v_29613;
wire v_29614;
wire v_29615;
wire v_29616;
wire v_29617;
wire v_29618;
wire v_29619;
wire v_29620;
wire v_29621;
wire v_29622;
wire v_29623;
wire v_29624;
wire v_29625;
wire v_29626;
wire v_29627;
wire v_29628;
wire v_29629;
wire v_29630;
wire v_29631;
wire v_29632;
wire v_29633;
wire v_29634;
wire v_29635;
wire v_29636;
wire v_29637;
wire v_29638;
wire v_29639;
wire v_29640;
wire v_29641;
wire v_29642;
wire v_29643;
wire v_29644;
wire v_29645;
wire v_29646;
wire v_29647;
wire v_29648;
wire v_29649;
wire v_29650;
wire v_29651;
wire v_29652;
wire v_29653;
wire v_29654;
wire v_29655;
wire v_29656;
wire v_29657;
wire v_29658;
wire v_29659;
wire v_29660;
wire v_29661;
wire v_29662;
wire v_29663;
wire v_29664;
wire v_29665;
wire v_29666;
wire v_29667;
wire v_29668;
wire v_29669;
wire v_29670;
wire v_29671;
wire v_29672;
wire v_29673;
wire v_29674;
wire v_29675;
wire v_29676;
wire v_29677;
wire v_29678;
wire v_29679;
wire v_29680;
wire v_29681;
wire v_29682;
wire v_29683;
wire v_29684;
wire v_29685;
wire v_29686;
wire v_29687;
wire v_29688;
wire v_29689;
wire v_29690;
wire v_29691;
wire v_29692;
wire v_29693;
wire v_29694;
wire v_29695;
wire v_29696;
wire v_29697;
wire v_29698;
wire v_29699;
wire v_29700;
wire v_29701;
wire v_29702;
wire v_29703;
wire v_29704;
wire v_29705;
wire v_29706;
wire v_29707;
wire v_29708;
wire v_29709;
wire v_29710;
wire v_29711;
wire v_29712;
wire v_29713;
wire v_29714;
wire v_29715;
wire v_29716;
wire v_29717;
wire v_29718;
wire v_29719;
wire v_29720;
wire v_29721;
wire v_29722;
wire v_29723;
wire v_29724;
wire v_29725;
wire v_29726;
wire v_29727;
wire v_29728;
wire v_29729;
wire v_29730;
wire v_29731;
wire v_29732;
wire v_29733;
wire v_29734;
wire v_29735;
wire v_29736;
wire v_29737;
wire v_29738;
wire v_29739;
wire v_29740;
wire v_29741;
wire v_29742;
wire v_29743;
wire v_29744;
wire v_29745;
wire v_29746;
wire v_29747;
wire v_29748;
wire v_29749;
wire v_29750;
wire v_29751;
wire v_29752;
wire v_29753;
wire v_29754;
wire v_29755;
wire v_29756;
wire v_29757;
wire v_29758;
wire v_29759;
wire v_29760;
wire v_29761;
wire v_29762;
wire v_29763;
wire v_29764;
wire v_29765;
wire v_29766;
wire v_29767;
wire v_29768;
wire v_29769;
wire v_29770;
wire v_29771;
wire v_29772;
wire v_29773;
wire v_29774;
wire v_29775;
wire v_29776;
wire v_29777;
wire v_29778;
wire v_29779;
wire v_29780;
wire v_29781;
wire v_29782;
wire v_29783;
wire v_29784;
wire v_29785;
wire v_29786;
wire v_29787;
wire v_29788;
wire v_29789;
wire v_29790;
wire v_29791;
wire v_29792;
wire v_29793;
wire v_29794;
wire v_29795;
wire v_29796;
wire v_29797;
wire v_29798;
wire v_29799;
wire v_29800;
wire v_29801;
wire v_29802;
wire v_29803;
wire v_29804;
wire v_29805;
wire v_29806;
wire v_29807;
wire v_29808;
wire v_29809;
wire v_29810;
wire v_29811;
wire v_29812;
wire v_29813;
wire v_29814;
wire v_29815;
wire v_29816;
wire v_29817;
wire v_29818;
wire v_29819;
wire v_29820;
wire v_29821;
wire v_29822;
wire v_29823;
wire v_29824;
wire v_29825;
wire v_29826;
wire v_29827;
wire v_29828;
wire v_29829;
wire v_29830;
wire v_29831;
wire v_29832;
wire v_29833;
wire v_29834;
wire v_29835;
wire v_29836;
wire v_29837;
wire v_29838;
wire v_29839;
wire v_29840;
wire v_29841;
wire v_29842;
wire v_29843;
wire v_29844;
wire v_29845;
wire v_29846;
wire v_29847;
wire v_29848;
wire v_29849;
wire v_29850;
wire v_29851;
wire v_29852;
wire v_29853;
wire v_29854;
wire v_29855;
wire v_29856;
wire v_29857;
wire v_29858;
wire v_29859;
wire v_29860;
wire v_29861;
wire v_29862;
wire v_29863;
wire v_29864;
wire v_29865;
wire v_29866;
wire v_29867;
wire v_29868;
wire v_29869;
wire v_29870;
wire v_29871;
wire v_29872;
wire v_29873;
wire v_29874;
wire v_29875;
wire v_29876;
wire v_29877;
wire v_29878;
wire v_29879;
wire v_29880;
wire v_29881;
wire v_29882;
wire v_29883;
wire v_29884;
wire v_29885;
wire v_29886;
wire v_29887;
wire v_29888;
wire v_29889;
wire v_29890;
wire v_29891;
wire v_29892;
wire v_29893;
wire v_29894;
wire v_29895;
wire v_29896;
wire v_29897;
wire v_29898;
wire v_29899;
wire v_29900;
wire v_29901;
wire v_29902;
wire v_29903;
wire v_29904;
wire v_29905;
wire v_29906;
wire v_29907;
wire v_29908;
wire v_29909;
wire v_29910;
wire v_29911;
wire v_29912;
wire v_29913;
wire v_29914;
wire v_29915;
wire v_29916;
wire v_29917;
wire v_29918;
wire v_29919;
wire v_29920;
wire v_29921;
wire v_29922;
wire v_29923;
wire v_29924;
wire v_29925;
wire v_29926;
wire v_29927;
wire v_29928;
wire v_29929;
wire v_29930;
wire v_29931;
wire v_29932;
wire v_29933;
wire v_29934;
wire v_29935;
wire v_29936;
wire v_29937;
wire v_29938;
wire v_29939;
wire v_29940;
wire v_29941;
wire v_29942;
wire v_29943;
wire v_29944;
wire v_29945;
wire v_29946;
wire v_29947;
wire v_29948;
wire v_29949;
wire v_29950;
wire v_29951;
wire v_29952;
wire v_29953;
wire v_29954;
wire v_29955;
wire v_29956;
wire v_29957;
wire v_29958;
wire v_29959;
wire v_29960;
wire v_29961;
wire v_29962;
wire v_29963;
wire v_29964;
wire v_29965;
wire v_29966;
wire v_29967;
wire v_29968;
wire v_29969;
wire v_29970;
wire v_29971;
wire v_29972;
wire v_29973;
wire v_29974;
wire v_29975;
wire v_29976;
wire v_29977;
wire v_29978;
wire v_29979;
wire v_29980;
wire v_29981;
wire v_29982;
wire v_29983;
wire v_29984;
wire v_29985;
wire v_29986;
wire v_29987;
wire v_29988;
wire v_29989;
wire v_29990;
wire v_29991;
wire v_29992;
wire v_29993;
wire v_29994;
wire v_29995;
wire v_29996;
wire v_29997;
wire v_29998;
wire v_29999;
wire v_30000;
wire v_30001;
wire v_30002;
wire v_30003;
wire v_30004;
wire v_30005;
wire v_30006;
wire v_30007;
wire v_30008;
wire v_30009;
wire v_30010;
wire v_30011;
wire v_30012;
wire v_30013;
wire v_30014;
wire v_30015;
wire v_30016;
wire v_30017;
wire v_30018;
wire v_30019;
wire v_30020;
wire v_30021;
wire v_30022;
wire v_30023;
wire v_30024;
wire v_30025;
wire v_30026;
wire v_30027;
wire v_30028;
wire v_30029;
wire v_30030;
wire v_30031;
wire v_30032;
wire v_30033;
wire v_30034;
wire v_30035;
wire v_30036;
wire v_30037;
wire v_30038;
wire v_30039;
wire v_30040;
wire v_30041;
wire v_30042;
wire v_30043;
wire v_30044;
wire v_30045;
wire v_30046;
wire v_30047;
wire v_30048;
wire v_30049;
wire v_30050;
wire v_30051;
wire v_30052;
wire v_30053;
wire v_30054;
wire v_30055;
wire v_30056;
wire v_30057;
wire v_30058;
wire v_30059;
wire v_30060;
wire v_30061;
wire v_30062;
wire v_30063;
wire v_30064;
wire v_30065;
wire v_30066;
wire v_30067;
wire v_30068;
wire v_30069;
wire v_30070;
wire v_30071;
wire v_30072;
wire v_30073;
wire v_30074;
wire v_30075;
wire v_30076;
wire v_30077;
wire v_30078;
wire v_30079;
wire v_30080;
wire v_30081;
wire v_30082;
wire v_30083;
wire v_30084;
wire v_30085;
wire v_30086;
wire v_30087;
wire v_30088;
wire v_30089;
wire v_30090;
wire v_30091;
wire v_30092;
wire v_30093;
wire v_30094;
wire v_30095;
wire v_30096;
wire v_30097;
wire v_30098;
wire v_30099;
wire v_30100;
wire v_30101;
wire v_30102;
wire v_30103;
wire v_30104;
wire v_30105;
wire v_30106;
wire v_30107;
wire v_30108;
wire v_30109;
wire v_30110;
wire v_30111;
wire v_30112;
wire v_30113;
wire v_30114;
wire v_30115;
wire v_30116;
wire v_30117;
wire v_30118;
wire v_30119;
wire v_30120;
wire v_30121;
wire v_30122;
wire v_30123;
wire v_30124;
wire v_30125;
wire v_30126;
wire v_30127;
wire v_30128;
wire v_30129;
wire v_30130;
wire v_30131;
wire v_30132;
wire v_30133;
wire v_30134;
wire v_30135;
wire v_30136;
wire v_30137;
wire v_30138;
wire v_30139;
wire v_30140;
wire v_30141;
wire v_30142;
wire v_30143;
wire v_30144;
wire v_30145;
wire v_30146;
wire v_30147;
wire v_30148;
wire v_30149;
wire v_30150;
wire v_30151;
wire v_30152;
wire v_30153;
wire v_30154;
wire v_30155;
wire v_30156;
wire v_30157;
wire v_30158;
wire v_30159;
wire v_30160;
wire v_30161;
wire v_30162;
wire v_30163;
wire v_30164;
wire v_30165;
wire v_30166;
wire v_30167;
wire v_30168;
wire v_30169;
wire v_30170;
wire v_30171;
wire v_30172;
wire v_30173;
wire v_30174;
wire v_30175;
wire v_30176;
wire v_30177;
wire v_30178;
wire v_30179;
wire v_30180;
wire v_30181;
wire v_30182;
wire v_30183;
wire v_30184;
wire v_30185;
wire v_30186;
wire v_30187;
wire v_30188;
wire v_30189;
wire v_30190;
wire v_30191;
wire v_30192;
wire v_30193;
wire v_30194;
wire v_30195;
wire v_30196;
wire v_30197;
wire v_30198;
wire v_30199;
wire v_30200;
wire v_30201;
wire v_30202;
wire v_30203;
wire v_30204;
wire v_30205;
wire v_30206;
wire v_30207;
wire v_30208;
wire v_30209;
wire v_30210;
wire v_30211;
wire v_30212;
wire v_30213;
wire v_30214;
wire v_30215;
wire v_30216;
wire v_30217;
wire v_30218;
wire v_30219;
wire v_30220;
wire v_30221;
wire v_30222;
wire v_30223;
wire v_30224;
wire v_30225;
wire v_30226;
wire v_30227;
wire v_30228;
wire v_30229;
wire v_30230;
wire v_30231;
wire v_30232;
wire v_30233;
wire v_30234;
wire v_30235;
wire v_30236;
wire v_30237;
wire v_30238;
wire v_30239;
wire v_30240;
wire v_30241;
wire v_30242;
wire v_30243;
wire v_30244;
wire v_30245;
wire v_30246;
wire v_30247;
wire v_30248;
wire v_30249;
wire v_30250;
wire v_30251;
wire v_30252;
wire v_30253;
wire v_30254;
wire v_30255;
wire v_30256;
wire v_30257;
wire v_30258;
wire v_30259;
wire v_30260;
wire v_30261;
wire v_30262;
wire v_30263;
wire v_30264;
wire v_30265;
wire v_30266;
wire v_30267;
wire v_30268;
wire v_30269;
wire v_30270;
wire v_30271;
wire v_30272;
wire v_30273;
wire v_30274;
wire v_30275;
wire v_30276;
wire v_30277;
wire v_30278;
wire v_30279;
wire v_30280;
wire v_30281;
wire v_30282;
wire v_30283;
wire v_30284;
wire v_30285;
wire v_30286;
wire v_30287;
wire v_30288;
wire v_30289;
wire v_30290;
wire v_30291;
wire v_30292;
wire v_30293;
wire v_30294;
wire v_30295;
wire v_30296;
wire v_30297;
wire v_30298;
wire v_30299;
wire v_30300;
wire v_30301;
wire v_30302;
wire v_30303;
wire v_30304;
wire v_30305;
wire v_30306;
wire v_30307;
wire v_30308;
wire v_30309;
wire v_30310;
wire v_30311;
wire v_30312;
wire v_30313;
wire v_30314;
wire v_30315;
wire v_30316;
wire v_30317;
wire v_30318;
wire v_30319;
wire v_30320;
wire v_30321;
wire v_30322;
wire v_30323;
wire v_30324;
wire v_30325;
wire v_30326;
wire v_30327;
wire v_30328;
wire v_30329;
wire v_30330;
wire v_30331;
wire v_30332;
wire v_30333;
wire v_30334;
wire v_30335;
wire v_30336;
wire v_30337;
wire v_30338;
wire v_30339;
wire v_30340;
wire v_30341;
wire v_30342;
wire v_30343;
wire v_30344;
wire v_30345;
wire v_30346;
wire v_30347;
wire v_30348;
wire v_30349;
wire v_30350;
wire v_30351;
wire v_30352;
wire v_30353;
wire v_30354;
wire v_30355;
wire v_30356;
wire v_30357;
wire v_30358;
wire v_30359;
wire v_30360;
wire v_30361;
wire v_30362;
wire v_30363;
wire v_30364;
wire v_30365;
wire v_30366;
wire v_30367;
wire v_30368;
wire v_30369;
wire v_30370;
wire v_30371;
wire v_30372;
wire v_30373;
wire v_30374;
wire v_30375;
wire v_30376;
wire v_30377;
wire v_30378;
wire v_30379;
wire v_30380;
wire v_30381;
wire v_30382;
wire v_30383;
wire v_30384;
wire v_30385;
wire v_30386;
wire v_30387;
wire v_30388;
wire v_30389;
wire v_30390;
wire v_30391;
wire v_30392;
wire v_30393;
wire v_30394;
wire v_30395;
wire v_30396;
wire v_30397;
wire v_30398;
wire v_30399;
wire v_30400;
wire v_30401;
wire v_30402;
wire v_30403;
wire v_30404;
wire v_30405;
wire v_30406;
wire v_30407;
wire v_30408;
wire v_30409;
wire v_30410;
wire v_30411;
wire v_30412;
wire v_30413;
wire v_30414;
wire v_30415;
wire v_30416;
wire v_30417;
wire v_30418;
wire v_30419;
wire v_30420;
wire v_30421;
wire v_30422;
wire v_30423;
wire v_30424;
wire v_30425;
wire v_30426;
wire v_30427;
wire v_30428;
wire v_30429;
wire v_30430;
wire v_30431;
wire v_30432;
wire v_30433;
wire v_30434;
wire v_30435;
wire v_30436;
wire v_30437;
wire v_30438;
wire v_30439;
wire v_30440;
wire v_30441;
wire v_30442;
wire v_30443;
wire v_30444;
wire v_30445;
wire v_30446;
wire v_30447;
wire v_30448;
wire v_30449;
wire v_30450;
wire v_30451;
wire v_30452;
wire v_30453;
wire v_30454;
wire v_30455;
wire v_30456;
wire v_30457;
wire v_30458;
wire v_30459;
wire v_30460;
wire v_30461;
wire v_30462;
wire v_30463;
wire v_30464;
wire v_30465;
wire v_30466;
wire v_30467;
wire v_30468;
wire v_30469;
wire v_30470;
wire v_30471;
wire v_30472;
wire v_30473;
wire v_30474;
wire v_30475;
wire v_30476;
wire v_30477;
wire v_30478;
wire v_30479;
wire v_30480;
wire v_30481;
wire v_30482;
wire v_30483;
wire v_30484;
wire v_30485;
wire v_30486;
wire v_30487;
wire v_30488;
wire v_30489;
wire v_30490;
wire v_30491;
wire v_30492;
wire v_30493;
wire v_30494;
wire v_30495;
wire v_30496;
wire v_30497;
wire v_30498;
wire v_30499;
wire v_30500;
wire v_30501;
wire v_30502;
wire v_30503;
wire v_30504;
wire v_30505;
wire v_30506;
wire v_30507;
wire v_30508;
wire v_30509;
wire v_30510;
wire v_30511;
wire v_30512;
wire v_30513;
wire v_30514;
wire v_30515;
wire v_30516;
wire v_30517;
wire v_30518;
wire v_30519;
wire v_30520;
wire v_30521;
wire v_30522;
wire v_30523;
wire v_30524;
wire v_30525;
wire v_30526;
wire v_30527;
wire v_30528;
wire v_30529;
wire v_30530;
wire v_30531;
wire v_30532;
wire v_30533;
wire v_30534;
wire v_30535;
wire v_30536;
wire v_30537;
wire v_30538;
wire v_30539;
wire v_30540;
wire v_30541;
wire v_30542;
wire v_30543;
wire v_30544;
wire v_30545;
wire v_30546;
wire v_30547;
wire v_30548;
wire v_30549;
wire v_30550;
wire v_30551;
wire v_30552;
wire v_30553;
wire v_30554;
wire v_30555;
wire v_30556;
wire v_30557;
wire v_30558;
wire v_30559;
wire v_30560;
wire v_30561;
wire v_30562;
wire v_30563;
wire v_30564;
wire v_30565;
wire v_30566;
wire v_30567;
wire v_30568;
wire v_30569;
wire v_30570;
wire v_30571;
wire v_30572;
wire v_30573;
wire v_30574;
wire v_30575;
wire v_30576;
wire v_30577;
wire v_30578;
wire v_30579;
wire v_30580;
wire v_30581;
wire v_30582;
wire v_30583;
wire v_30584;
wire v_30585;
wire v_30586;
wire v_30587;
wire v_30588;
wire v_30589;
wire v_30590;
wire v_30591;
wire v_30592;
wire v_30593;
wire v_30594;
wire v_30595;
wire v_30596;
wire v_30597;
wire v_30598;
wire v_30599;
wire v_30600;
wire v_30601;
wire v_30602;
wire v_30603;
wire v_30604;
wire v_30605;
wire v_30606;
wire v_30607;
wire v_30608;
wire v_30609;
wire v_30610;
wire v_30611;
wire v_30612;
wire v_30613;
wire v_30614;
wire v_30615;
wire v_30616;
wire v_30617;
wire v_30618;
wire v_30619;
wire v_30620;
wire v_30621;
wire v_30622;
wire v_30623;
wire v_30624;
wire v_30625;
wire v_30626;
wire v_30627;
wire v_30628;
wire v_30629;
wire v_30630;
wire v_30631;
wire v_30632;
wire v_30633;
wire v_30634;
wire v_30635;
wire v_30636;
wire v_30637;
wire v_30638;
wire v_30639;
wire v_30640;
wire v_30641;
wire v_30642;
wire v_30643;
wire v_30644;
wire v_30645;
wire v_30646;
wire v_30647;
wire v_30648;
wire v_30649;
wire v_30650;
wire v_30651;
wire v_30652;
wire v_30653;
wire v_30654;
wire v_30655;
wire v_30656;
wire v_30657;
wire v_30658;
wire v_30659;
wire v_30660;
wire v_30661;
wire v_30662;
wire v_30663;
wire v_30664;
wire v_30665;
wire v_30666;
wire v_30667;
wire v_30668;
wire v_30669;
wire v_30670;
wire v_30671;
wire v_30672;
wire v_30673;
wire v_30674;
wire v_30675;
wire v_30676;
wire v_30677;
wire v_30678;
wire v_30679;
wire v_30680;
wire v_30681;
wire v_30682;
wire v_30683;
wire v_30684;
wire v_30685;
wire v_30686;
wire v_30687;
wire v_30688;
wire v_30689;
wire v_30690;
wire v_30691;
wire v_30692;
wire v_30693;
wire v_30694;
wire v_30695;
wire v_30696;
wire v_30697;
wire v_30698;
wire v_30699;
wire v_30700;
wire v_30701;
wire v_30702;
wire v_30703;
wire v_30704;
wire v_30705;
wire v_30706;
wire v_30707;
wire v_30708;
wire v_30709;
wire v_30710;
wire v_30711;
wire v_30712;
wire v_30713;
wire v_30714;
wire v_30715;
wire v_30716;
wire v_30717;
wire v_30718;
wire v_30719;
wire v_30720;
wire v_30721;
wire v_30722;
wire v_30723;
wire v_30724;
wire v_30725;
wire v_30726;
wire v_30727;
wire v_30728;
wire v_30729;
wire v_30730;
wire v_30731;
wire v_30732;
wire v_30733;
wire v_30734;
wire v_30735;
wire v_30736;
wire v_30737;
wire v_30738;
wire v_30739;
wire v_30740;
wire v_30741;
wire v_30742;
wire v_30743;
wire v_30744;
wire v_30745;
wire v_30746;
wire v_30747;
wire v_30748;
wire v_30749;
wire v_30750;
wire v_30751;
wire v_30752;
wire v_30753;
wire v_30754;
wire v_30755;
wire v_30756;
wire v_30757;
wire v_30758;
wire v_30759;
wire v_30760;
wire v_30761;
wire v_30762;
wire v_30763;
wire v_30764;
wire v_30765;
wire v_30766;
wire v_30767;
wire v_30768;
wire v_30769;
wire v_30770;
wire v_30771;
wire v_30772;
wire v_30773;
wire v_30774;
wire v_30775;
wire v_30776;
wire v_30777;
wire v_30778;
wire v_30779;
wire v_30780;
wire v_30781;
wire v_30782;
wire v_30783;
wire v_30784;
wire v_30785;
wire v_30786;
wire v_30787;
wire v_30788;
wire v_30789;
wire v_30790;
wire v_30791;
wire v_30792;
wire v_30793;
wire v_30794;
wire v_30795;
wire v_30796;
wire v_30797;
wire v_30798;
wire v_30799;
wire v_30800;
wire v_30801;
wire v_30802;
wire v_30803;
wire v_30804;
wire v_30805;
wire v_30806;
wire v_30807;
wire v_30808;
wire v_30809;
wire v_30810;
wire v_30811;
wire v_30812;
wire v_30813;
wire v_30814;
wire v_30815;
wire v_30816;
wire v_30817;
wire v_30818;
wire v_30819;
wire v_30820;
wire v_30821;
wire v_30822;
wire v_30823;
wire v_30824;
wire v_30825;
wire v_30826;
wire v_30827;
wire v_30828;
wire v_30829;
wire v_30830;
wire v_30831;
wire v_30832;
wire v_30833;
wire v_30834;
wire v_30835;
wire v_30836;
wire v_30837;
wire v_30838;
wire v_30839;
wire v_30840;
wire v_30841;
wire v_30842;
wire v_30843;
wire v_30844;
wire v_30845;
wire v_30846;
wire v_30847;
wire v_30848;
wire v_30849;
wire v_30850;
wire v_30851;
wire v_30852;
wire v_30853;
wire v_30854;
wire v_30855;
wire v_30856;
wire v_30857;
wire v_30858;
wire v_30859;
wire v_30860;
wire v_30861;
wire v_30862;
wire v_30863;
wire v_30864;
wire v_30865;
wire v_30866;
wire v_30867;
wire v_30868;
wire v_30869;
wire v_30870;
wire v_30871;
wire v_30872;
wire v_30873;
wire v_30874;
wire v_30875;
wire v_30876;
wire v_30877;
wire v_30878;
wire v_30879;
wire v_30880;
wire v_30881;
wire v_30882;
wire v_30883;
wire v_30884;
wire v_30885;
wire v_30886;
wire v_30887;
wire v_30888;
wire v_30889;
wire v_30890;
wire v_30891;
wire v_30892;
wire v_30893;
wire v_30894;
wire v_30895;
wire v_30896;
wire v_30897;
wire v_30898;
wire v_30899;
wire v_30900;
wire v_30901;
wire v_30902;
wire v_30903;
wire v_30904;
wire v_30905;
wire v_30906;
wire v_30907;
wire v_30908;
wire v_30909;
wire v_30910;
wire v_30911;
wire v_30912;
wire v_30913;
wire v_30914;
wire v_30915;
wire v_30916;
wire v_30917;
wire v_30918;
wire v_30919;
wire v_30920;
wire v_30921;
wire v_30922;
wire v_30923;
wire v_30924;
wire v_30925;
wire v_30926;
wire v_30927;
wire v_30928;
wire v_30929;
wire v_30930;
wire v_30931;
wire v_30932;
wire v_30933;
wire v_30934;
wire v_30935;
wire v_30936;
wire v_30937;
wire v_30938;
wire v_30939;
wire v_30940;
wire v_30941;
wire v_30942;
wire v_30943;
wire v_30944;
wire v_30945;
wire v_30946;
wire v_30947;
wire v_30948;
wire v_30949;
wire v_30950;
wire v_30951;
wire v_30952;
wire v_30953;
wire v_30954;
wire v_30955;
wire v_30956;
wire v_30957;
wire v_30958;
wire v_30959;
wire v_30960;
wire v_30961;
wire v_30962;
wire v_30963;
wire v_30964;
wire v_30965;
wire v_30966;
wire v_30967;
wire v_30968;
wire v_30969;
wire v_30970;
wire v_30971;
wire v_30972;
wire v_30973;
wire v_30974;
wire v_30975;
wire v_30976;
wire v_30977;
wire v_30978;
wire v_30979;
wire v_30980;
wire v_30981;
wire v_30982;
wire v_30983;
wire v_30984;
wire v_30985;
wire v_30986;
wire v_30987;
wire v_30988;
wire v_30989;
wire v_30990;
wire v_30991;
wire v_30992;
wire v_30993;
wire v_30994;
wire v_30995;
wire v_30996;
wire v_30997;
wire v_30998;
wire v_30999;
wire v_31000;
wire v_31001;
wire v_31002;
wire v_31003;
wire v_31004;
wire v_31005;
wire v_31006;
wire v_31007;
wire v_31008;
wire v_31009;
wire v_31010;
wire v_31011;
wire v_31012;
wire v_31013;
wire v_31014;
wire v_31015;
wire v_31016;
wire v_31017;
wire v_31018;
wire v_31019;
wire v_31020;
wire v_31021;
wire v_31022;
wire v_31023;
wire v_31024;
wire v_31025;
wire v_31026;
wire v_31027;
wire v_31028;
wire v_31029;
wire v_31030;
wire v_31031;
wire v_31032;
wire v_31033;
wire v_31034;
wire v_31035;
wire v_31036;
wire v_31037;
wire v_31038;
wire v_31039;
wire v_31040;
wire v_31041;
wire v_31042;
wire v_31043;
wire v_31044;
wire v_31045;
wire v_31046;
wire v_31047;
wire v_31048;
wire v_31049;
wire v_31050;
wire v_31051;
wire v_31052;
wire v_31053;
wire v_31054;
wire v_31055;
wire v_31056;
wire v_31057;
wire v_31058;
wire v_31059;
wire v_31060;
wire v_31061;
wire v_31062;
wire v_31063;
wire v_31064;
wire v_31065;
wire v_31066;
wire v_31067;
wire v_31068;
wire v_31069;
wire v_31070;
wire v_31071;
wire v_31072;
wire v_31073;
wire v_31074;
wire v_31075;
wire v_31076;
wire v_31077;
wire v_31078;
wire v_31079;
wire v_31080;
wire v_31081;
wire v_31082;
wire v_31083;
wire v_31084;
wire v_31085;
wire v_31086;
wire v_31087;
wire v_31088;
wire v_31089;
wire v_31090;
wire v_31091;
wire v_31092;
wire v_31093;
wire v_31094;
wire v_31095;
wire v_31096;
wire v_31097;
wire v_31098;
wire v_31099;
wire v_31100;
wire v_31101;
wire v_31102;
wire v_31103;
wire v_31104;
wire v_31105;
wire v_31106;
wire v_31107;
wire v_31108;
wire v_31109;
wire v_31110;
wire v_31111;
wire v_31112;
wire v_31113;
wire v_31114;
wire v_31115;
wire v_31116;
wire v_31117;
wire v_31118;
wire v_31119;
wire v_31120;
wire v_31121;
wire v_31122;
wire v_31123;
wire v_31124;
wire v_31125;
wire v_31126;
wire v_31127;
wire v_31128;
wire v_31129;
wire v_31130;
wire v_31131;
wire v_31132;
wire v_31133;
wire v_31134;
wire v_31135;
wire v_31136;
wire v_31137;
wire v_31138;
wire v_31139;
wire v_31140;
wire v_31141;
wire v_31142;
wire v_31143;
wire v_31144;
wire v_31145;
wire v_31146;
wire v_31147;
wire v_31148;
wire v_31149;
wire v_31150;
wire v_31151;
wire v_31152;
wire v_31153;
wire v_31154;
wire v_31155;
wire v_31156;
wire v_31157;
wire v_31158;
wire v_31159;
wire v_31160;
wire v_31161;
wire v_31162;
wire v_31163;
wire v_31164;
wire v_31165;
wire v_31166;
wire v_31167;
wire v_31168;
wire v_31169;
wire v_31170;
wire v_31171;
wire v_31172;
wire v_31173;
wire v_31174;
wire v_31175;
wire v_31176;
wire v_31177;
wire v_31178;
wire v_31179;
wire v_31180;
wire v_31181;
wire v_31182;
wire v_31183;
wire v_31184;
wire v_31185;
wire v_31186;
wire v_31187;
wire v_31188;
wire v_31189;
wire v_31190;
wire v_31191;
wire v_31192;
wire v_31193;
wire v_31194;
wire v_31195;
wire v_31196;
wire v_31197;
wire v_31198;
wire v_31199;
wire v_31200;
wire v_31201;
wire v_31202;
wire v_31203;
wire v_31204;
wire v_31205;
wire v_31206;
wire v_31207;
wire v_31208;
wire v_31209;
wire v_31210;
wire v_31211;
wire v_31212;
wire v_31213;
wire v_31214;
wire v_31215;
wire v_31216;
wire v_31217;
wire v_31218;
wire v_31219;
wire v_31220;
wire v_31221;
wire v_31222;
wire v_31223;
wire v_31224;
wire v_31225;
wire v_31226;
wire v_31227;
wire v_31228;
wire v_31229;
wire v_31230;
wire v_31231;
wire v_31232;
wire v_31233;
wire v_31234;
wire v_31235;
wire v_31236;
wire v_31237;
wire v_31238;
wire v_31239;
wire v_31240;
wire v_31241;
wire v_31242;
wire v_31243;
wire v_31244;
wire v_31245;
wire v_31246;
wire v_31247;
wire v_31248;
wire v_31249;
wire v_31250;
wire v_31251;
wire v_31252;
wire v_31253;
wire v_31254;
wire v_31255;
wire v_31256;
wire v_31257;
wire v_31258;
wire v_31259;
wire v_31260;
wire v_31261;
wire v_31262;
wire v_31263;
wire v_31264;
wire v_31265;
wire v_31266;
wire v_31267;
wire v_31268;
wire v_31269;
wire v_31270;
wire v_31271;
wire v_31272;
wire v_31273;
wire v_31274;
wire v_31275;
wire v_31276;
wire v_31277;
wire v_31278;
wire v_31279;
wire v_31280;
wire v_31281;
wire v_31282;
wire v_31283;
wire v_31284;
wire v_31285;
wire v_31286;
wire v_31287;
wire v_31288;
wire v_31289;
wire v_31290;
wire v_31291;
wire v_31292;
wire v_31293;
wire v_31294;
wire v_31295;
wire v_31296;
wire v_31297;
wire v_31298;
wire v_31299;
wire v_31300;
wire v_31301;
wire v_31302;
wire v_31303;
wire v_31304;
wire v_31305;
wire v_31306;
wire v_31307;
wire v_31308;
wire v_31309;
wire v_31310;
wire v_31311;
wire v_31312;
wire v_31313;
wire v_31314;
wire v_31315;
wire v_31316;
wire v_31317;
wire v_31318;
wire v_31319;
wire v_31320;
wire v_31321;
wire v_31322;
wire v_31323;
wire v_31324;
wire v_31325;
wire v_31326;
wire v_31327;
wire v_31328;
wire v_31329;
wire v_31330;
wire v_31331;
wire v_31332;
wire v_31333;
wire v_31334;
wire v_31335;
wire v_31336;
wire v_31337;
wire v_31338;
wire v_31339;
wire v_31340;
wire v_31341;
wire v_31342;
wire v_31343;
wire v_31344;
wire v_31345;
wire v_31346;
wire v_31347;
wire v_31348;
wire v_31349;
wire v_31350;
wire v_31351;
wire v_31352;
wire v_31353;
wire v_31354;
wire v_31355;
wire v_31356;
wire v_31357;
wire v_31358;
wire v_31359;
wire v_31360;
wire v_31361;
wire v_31362;
wire v_31363;
wire v_31364;
wire v_31365;
wire v_31366;
wire v_31367;
wire v_31368;
wire v_31369;
wire v_31370;
wire v_31371;
wire v_31372;
wire v_31373;
wire v_31374;
wire v_31375;
wire v_31376;
wire v_31377;
wire v_31378;
wire v_31379;
wire v_31380;
wire v_31381;
wire v_31382;
wire v_31383;
wire v_31384;
wire v_31385;
wire v_31386;
wire v_31387;
wire v_31388;
wire v_31389;
wire v_31390;
wire v_31391;
wire v_31392;
wire v_31393;
wire v_31394;
wire v_31395;
wire v_31396;
wire v_31397;
wire v_31398;
wire v_31399;
wire v_31400;
wire v_31401;
wire v_31402;
wire v_31403;
wire v_31404;
wire v_31405;
wire v_31406;
wire v_31407;
wire v_31408;
wire v_31409;
wire v_31410;
wire v_31411;
wire v_31412;
wire v_31413;
wire v_31414;
wire v_31415;
wire v_31416;
wire v_31417;
wire v_31418;
wire v_31419;
wire v_31420;
wire v_31421;
wire v_31422;
wire v_31423;
wire v_31424;
wire v_31425;
wire v_31426;
wire v_31427;
wire v_31428;
wire v_31429;
wire v_31430;
wire v_31431;
wire v_31432;
wire v_31433;
wire v_31434;
wire v_31435;
wire v_31436;
wire v_31437;
wire v_31438;
wire v_31439;
wire v_31440;
wire v_31441;
wire v_31442;
wire v_31443;
wire v_31444;
wire v_31445;
wire v_31446;
wire v_31447;
wire v_31448;
wire v_31449;
wire v_31450;
wire v_31451;
wire v_31452;
wire v_31453;
wire v_31454;
wire v_31455;
wire v_31456;
wire v_31457;
wire v_31458;
wire v_31459;
wire v_31460;
wire v_31461;
wire v_31462;
wire v_31463;
wire v_31464;
wire v_31465;
wire v_31466;
wire v_31467;
wire v_31468;
wire v_31469;
wire v_31470;
wire v_31471;
wire v_31472;
wire v_31473;
wire v_31474;
wire v_31475;
wire v_31476;
wire v_31477;
wire v_31478;
wire v_31479;
wire v_31480;
wire v_31481;
wire v_31482;
wire v_31483;
wire v_31484;
wire v_31485;
wire v_31486;
wire v_31487;
wire v_31488;
wire v_31489;
wire v_31490;
wire v_31491;
wire v_31492;
wire v_31493;
wire v_31494;
wire v_31495;
wire v_31496;
wire v_31497;
wire v_31498;
wire v_31499;
wire v_31500;
wire v_31501;
wire v_31502;
wire v_31503;
wire v_31504;
wire v_31505;
wire v_31506;
wire v_31507;
wire v_31508;
wire v_31509;
wire v_31510;
wire v_31511;
wire v_31512;
wire v_31513;
wire v_31514;
wire v_31515;
wire v_31516;
wire v_31517;
wire v_31518;
wire v_31519;
wire v_31520;
wire v_31521;
wire v_31522;
wire v_31523;
wire v_31524;
wire v_31525;
wire v_31526;
wire v_31527;
wire v_31528;
wire v_31529;
wire v_31530;
wire v_31531;
wire v_31532;
wire v_31533;
wire v_31534;
wire v_31535;
wire v_31536;
wire v_31537;
wire v_31538;
wire v_31539;
wire v_31540;
wire v_31541;
wire v_31542;
wire v_31543;
wire v_31544;
wire v_31545;
wire v_31546;
wire v_31547;
wire v_31548;
wire v_31549;
wire v_31550;
wire v_31551;
wire v_31552;
wire v_31553;
wire v_31554;
wire v_31555;
wire v_31556;
wire v_31557;
wire v_31558;
wire v_31559;
wire v_31560;
wire v_31561;
wire v_31562;
wire v_31563;
wire v_31564;
wire v_31565;
wire v_31566;
wire v_31567;
wire v_31568;
wire v_31569;
wire v_31570;
wire v_31571;
wire v_31572;
wire v_31573;
wire v_31574;
wire v_31575;
wire v_31576;
wire v_31577;
wire v_31578;
wire v_31579;
wire v_31580;
wire v_31581;
wire v_31582;
wire v_31583;
wire v_31584;
wire v_31585;
wire v_31586;
wire v_31587;
wire v_31588;
wire v_31589;
wire v_31590;
wire v_31591;
wire v_31592;
wire v_31593;
wire v_31594;
wire v_31595;
wire v_31596;
wire v_31597;
wire v_31598;
wire v_31599;
wire v_31600;
wire v_31601;
wire v_31602;
wire v_31603;
wire v_31604;
wire v_31605;
wire v_31606;
wire v_31607;
wire v_31608;
wire v_31609;
wire v_31610;
wire v_31611;
wire v_31612;
wire v_31613;
wire v_31614;
wire v_31615;
wire v_31616;
wire v_31617;
wire v_31618;
wire v_31619;
wire v_31620;
wire v_31621;
wire v_31622;
wire v_31623;
wire v_31624;
wire v_31625;
wire v_31626;
wire v_31627;
wire v_31628;
wire v_31629;
wire v_31630;
wire v_31631;
wire v_31632;
wire v_31633;
wire v_31634;
wire v_31635;
wire v_31636;
wire v_31637;
wire v_31638;
wire v_31639;
wire v_31640;
wire v_31641;
wire v_31642;
wire v_31643;
wire v_31644;
wire v_31645;
wire v_31646;
wire v_31647;
wire v_31648;
wire v_31649;
wire v_31650;
wire v_31651;
wire v_31652;
wire v_31653;
wire v_31654;
wire v_31655;
wire v_31656;
wire v_31657;
wire v_31658;
wire v_31659;
wire v_31660;
wire v_31661;
wire v_31662;
wire v_31663;
wire v_31664;
wire v_31665;
wire v_31666;
wire v_31667;
wire v_31668;
wire v_31669;
wire v_31670;
wire v_31671;
wire v_31672;
wire v_31673;
wire v_31674;
wire v_31675;
wire v_31676;
wire v_31677;
wire v_31678;
wire v_31679;
wire v_31680;
wire v_31681;
wire v_31682;
wire v_31683;
wire v_31684;
wire v_31685;
wire v_31686;
wire v_31687;
wire v_31688;
wire v_31689;
wire v_31690;
wire v_31691;
wire v_31692;
wire v_31693;
wire v_31694;
wire v_31695;
wire v_31696;
wire v_31697;
wire v_31698;
wire v_31699;
wire v_31700;
wire v_31701;
wire v_31702;
wire v_31703;
wire v_31704;
wire v_31705;
wire v_31706;
wire v_31707;
wire v_31708;
wire v_31709;
wire v_31710;
wire v_31711;
wire v_31712;
wire v_31713;
wire v_31714;
wire v_31715;
wire v_31716;
wire v_31717;
wire v_31718;
wire v_31719;
wire v_31720;
wire v_31721;
wire v_31722;
wire v_31723;
wire v_31724;
wire v_31725;
wire v_31726;
wire v_31727;
wire v_31728;
wire v_31729;
wire v_31730;
wire v_31731;
wire v_31732;
wire v_31733;
wire v_31734;
wire v_31735;
wire v_31736;
wire v_31737;
wire v_31738;
wire v_31739;
wire v_31740;
wire v_31741;
wire v_31742;
wire v_31743;
wire v_31744;
wire v_31745;
wire v_31746;
wire v_31747;
wire v_31748;
wire v_31749;
wire v_31750;
wire v_31751;
wire v_31752;
wire v_31753;
wire v_31754;
wire v_31755;
wire v_31756;
wire v_31757;
wire v_31758;
wire v_31759;
wire v_31760;
wire v_31761;
wire v_31762;
wire v_31763;
wire v_31764;
wire v_31765;
wire v_31766;
wire v_31767;
wire v_31768;
wire v_31769;
wire v_31770;
wire v_31771;
wire v_31772;
wire v_31773;
wire v_31774;
wire v_31775;
wire v_31776;
wire v_31777;
wire v_31778;
wire v_31779;
wire v_31780;
wire v_31781;
wire v_31782;
wire v_31783;
wire v_31784;
wire v_31785;
wire v_31786;
wire v_31787;
wire v_31788;
wire v_31789;
wire v_31790;
wire v_31791;
wire v_31792;
wire v_31793;
wire v_31794;
wire v_31795;
wire v_31796;
wire v_31797;
wire v_31798;
wire v_31799;
wire v_31800;
wire v_31801;
wire v_31802;
wire v_31803;
wire v_31804;
wire v_31805;
wire v_31806;
wire v_31807;
wire v_31808;
wire v_31809;
wire v_31810;
wire v_31811;
wire v_31812;
wire v_31813;
wire v_31814;
wire v_31815;
wire v_31816;
wire v_31817;
wire v_31818;
wire v_31819;
wire v_31820;
wire v_31821;
wire v_31822;
wire v_31823;
wire v_31824;
wire v_31825;
wire v_31826;
wire v_31827;
wire v_31828;
wire v_31829;
wire v_31830;
wire v_31831;
wire v_31832;
wire v_31833;
wire v_31834;
wire v_31835;
wire v_31836;
wire v_31837;
wire v_31838;
wire v_31839;
wire v_31840;
wire v_31841;
wire v_31842;
wire v_31843;
wire v_31844;
wire v_31845;
wire v_31846;
wire v_31847;
wire v_31848;
wire v_31849;
wire v_31850;
wire v_31851;
wire v_31852;
wire v_31853;
wire v_31854;
wire v_31855;
wire v_31856;
wire v_31857;
wire v_31858;
wire v_31859;
wire v_31860;
wire v_31861;
wire v_31862;
wire v_31863;
wire v_31864;
wire v_31865;
wire v_31866;
wire v_31867;
wire v_31868;
wire v_31869;
wire v_31870;
wire v_31871;
wire v_31872;
wire v_31873;
wire v_31874;
wire v_31875;
wire v_31876;
wire v_31877;
wire v_31878;
wire v_31879;
wire v_31880;
wire v_31881;
wire v_31882;
wire v_31883;
wire v_31884;
wire v_31885;
wire v_31886;
wire v_31887;
wire v_31888;
wire v_31889;
wire v_31890;
wire v_31891;
wire v_31892;
wire v_31893;
wire v_31894;
wire v_31895;
wire v_31896;
wire v_31897;
wire v_31898;
wire v_31899;
wire v_31900;
wire v_31901;
wire v_31902;
wire v_31903;
wire v_31904;
wire v_31905;
wire v_31906;
wire v_31907;
wire v_31908;
wire v_31909;
wire v_31910;
wire v_31911;
wire v_31912;
wire v_31913;
wire v_31914;
wire v_31915;
wire v_31916;
wire v_31917;
wire v_31918;
wire v_31919;
wire v_31920;
wire v_31921;
wire v_31922;
wire v_31923;
wire v_31924;
wire v_31925;
wire v_31926;
wire v_31927;
wire v_31928;
wire v_31929;
wire v_31930;
wire v_31931;
wire v_31932;
wire v_31933;
wire v_31934;
wire v_31935;
wire v_31936;
wire v_31937;
wire v_31938;
wire v_31939;
wire v_31940;
wire v_31941;
wire v_31942;
wire v_31943;
wire v_31944;
wire v_31945;
wire v_31946;
wire v_31947;
wire v_31948;
wire v_31949;
wire v_31950;
wire v_31951;
wire v_31952;
wire v_31953;
wire v_31954;
wire v_31955;
wire v_31956;
wire v_31957;
wire v_31958;
wire v_31959;
wire v_31960;
wire v_31961;
wire v_31962;
wire v_31963;
wire v_31964;
wire v_31965;
wire v_31966;
wire v_31967;
wire v_31968;
wire v_31969;
wire v_31970;
wire v_31971;
wire v_31972;
wire v_31973;
wire v_31974;
wire v_31975;
wire v_31976;
wire v_31977;
wire v_31978;
wire v_31979;
wire v_31980;
wire v_31981;
wire v_31982;
wire v_31983;
wire v_31984;
wire v_31985;
wire v_31986;
wire v_31987;
wire v_31988;
wire v_31989;
wire v_31990;
wire v_31991;
wire v_31992;
wire v_31993;
wire v_31994;
wire v_31995;
wire v_31996;
wire v_31997;
wire v_31998;
wire v_31999;
wire v_32000;
wire v_32001;
wire v_32002;
wire v_32003;
wire v_32004;
wire v_32005;
wire v_32006;
wire v_32007;
wire v_32008;
wire v_32009;
wire v_32010;
wire v_32011;
wire v_32012;
wire v_32013;
wire v_32014;
wire v_32015;
wire v_32016;
wire v_32017;
wire v_32018;
wire v_32019;
wire v_32020;
wire v_32021;
wire v_32022;
wire v_32023;
wire v_32024;
wire v_32025;
wire v_32026;
wire v_32027;
wire v_32028;
wire v_32029;
wire v_32030;
wire v_32031;
wire v_32032;
wire v_32033;
wire v_32034;
wire v_32035;
wire v_32036;
wire v_32037;
wire v_32038;
wire v_32039;
wire v_32040;
wire v_32041;
wire v_32042;
wire v_32043;
wire v_32044;
wire v_32045;
wire v_32046;
wire v_32047;
wire v_32048;
wire v_32049;
wire v_32050;
wire v_32051;
wire v_32052;
wire v_32053;
wire v_32054;
wire v_32055;
wire v_32056;
wire v_32057;
wire v_32058;
wire v_32059;
wire v_32060;
wire v_32061;
wire v_32062;
wire v_32063;
wire v_32064;
wire v_32065;
wire v_32066;
wire v_32067;
wire v_32068;
wire v_32069;
wire v_32070;
wire v_32071;
wire v_32072;
wire v_32073;
wire v_32074;
wire v_32075;
wire v_32076;
wire v_32077;
wire v_32078;
wire v_32079;
wire v_32080;
wire v_32081;
wire v_32082;
wire v_32083;
wire v_32084;
wire v_32085;
wire v_32086;
wire v_32087;
wire v_32088;
wire v_32089;
wire v_32090;
wire v_32091;
wire v_32092;
wire v_32093;
wire v_32094;
wire v_32095;
wire v_32096;
wire v_32097;
wire v_32098;
wire v_32099;
wire v_32100;
wire v_32101;
wire v_32102;
wire v_32103;
wire v_32104;
wire v_32105;
wire v_32106;
wire v_32107;
wire v_32108;
wire v_32109;
wire v_32110;
wire v_32111;
wire v_32112;
wire v_32113;
wire v_32114;
wire v_32115;
wire v_32116;
wire v_32117;
wire v_32118;
wire v_32119;
wire v_32120;
wire v_32121;
wire v_32122;
wire v_32123;
wire v_32124;
wire v_32125;
wire v_32126;
wire v_32127;
wire v_32128;
wire v_32129;
wire v_32130;
wire v_32131;
wire v_32132;
wire v_32133;
wire v_32134;
wire v_32135;
wire v_32136;
wire v_32137;
wire v_32138;
wire v_32139;
wire v_32140;
wire v_32141;
wire v_32142;
wire v_32143;
wire v_32144;
wire v_32145;
wire v_32146;
wire v_32147;
wire v_32148;
wire v_32149;
wire v_32150;
wire v_32151;
wire v_32152;
wire v_32153;
wire v_32154;
wire v_32155;
wire v_32156;
wire v_32157;
wire v_32158;
wire v_32159;
wire v_32160;
wire v_32161;
wire v_32162;
wire v_32163;
wire v_32164;
wire v_32165;
wire v_32166;
wire v_32167;
wire v_32168;
wire v_32169;
wire v_32170;
wire v_32171;
wire v_32172;
wire v_32173;
wire v_32174;
wire v_32175;
wire v_32176;
wire v_32177;
wire v_32178;
wire v_32179;
wire v_32180;
wire v_32181;
wire v_32182;
wire v_32183;
wire v_32184;
wire v_32185;
wire v_32186;
wire v_32187;
wire v_32188;
wire v_32189;
wire v_32190;
wire v_32191;
wire v_32192;
wire v_32193;
wire v_32194;
wire v_32195;
wire v_32196;
wire v_32197;
wire v_32198;
wire v_32199;
wire v_32200;
wire v_32201;
wire v_32202;
wire v_32203;
wire v_32204;
wire v_32205;
wire v_32206;
wire v_32207;
wire v_32208;
wire v_32209;
wire v_32210;
wire v_32211;
wire v_32212;
wire v_32213;
wire v_32214;
wire v_32215;
wire v_32216;
wire v_32217;
wire v_32218;
wire v_32219;
wire v_32220;
wire v_32221;
wire v_32222;
wire v_32223;
wire v_32224;
wire v_32225;
wire v_32226;
wire v_32227;
wire v_32228;
wire v_32229;
wire v_32230;
wire v_32231;
wire v_32232;
wire v_32233;
wire v_32234;
wire v_32235;
wire v_32236;
wire v_32237;
wire v_32238;
wire v_32239;
wire v_32240;
wire v_32241;
wire v_32242;
wire v_32243;
wire v_32244;
wire v_32245;
wire v_32246;
wire v_32247;
wire v_32248;
wire v_32249;
wire v_32250;
wire v_32251;
wire v_32252;
wire v_32253;
wire v_32254;
wire v_32255;
wire v_32256;
wire v_32257;
wire v_32258;
wire v_32259;
wire v_32260;
wire v_32261;
wire v_32262;
wire v_32263;
wire v_32264;
wire v_32265;
wire v_32266;
wire v_32267;
wire v_32268;
wire v_32269;
wire v_32270;
wire v_32271;
wire v_32272;
wire v_32273;
wire v_32274;
wire v_32275;
wire v_32276;
wire v_32277;
wire v_32278;
wire v_32279;
wire v_32280;
wire v_32281;
wire v_32282;
wire v_32283;
wire v_32284;
wire v_32285;
wire v_32286;
wire v_32287;
wire v_32288;
wire v_32289;
wire v_32290;
wire v_32291;
wire v_32292;
wire v_32293;
wire v_32294;
wire v_32295;
wire v_32296;
wire v_32297;
wire v_32298;
wire v_32299;
wire v_32300;
wire v_32301;
wire v_32302;
wire v_32303;
wire v_32304;
wire v_32305;
wire v_32306;
wire v_32307;
wire v_32308;
wire v_32309;
wire v_32310;
wire v_32311;
wire v_32312;
wire v_32313;
wire v_32314;
wire v_32315;
wire v_32316;
wire v_32317;
wire v_32318;
wire v_32319;
wire v_32320;
wire v_32321;
wire v_32322;
wire v_32323;
wire v_32324;
wire v_32325;
wire v_32326;
wire v_32327;
wire v_32328;
wire v_32329;
wire v_32330;
wire v_32331;
wire v_32332;
wire v_32333;
wire v_32334;
wire v_32335;
wire v_32336;
wire v_32337;
wire v_32338;
wire v_32339;
wire v_32340;
wire v_32341;
wire v_32342;
wire v_32343;
wire v_32344;
wire v_32345;
wire v_32346;
wire v_32347;
wire v_32348;
wire v_32349;
wire v_32350;
wire v_32351;
wire v_32352;
wire v_32353;
wire v_32354;
wire v_32355;
wire v_32356;
wire v_32357;
wire v_32358;
wire v_32359;
wire v_32360;
wire v_32361;
wire v_32362;
wire v_32363;
wire v_32364;
wire v_32365;
wire v_32366;
wire v_32367;
wire v_32368;
wire v_32369;
wire v_32370;
wire v_32371;
wire v_32372;
wire v_32373;
wire v_32374;
wire v_32375;
wire v_32376;
wire v_32377;
wire v_32378;
wire v_32379;
wire v_32380;
wire v_32381;
wire v_32382;
wire v_32383;
wire v_32384;
wire v_32385;
wire v_32386;
wire v_32387;
wire v_32388;
wire v_32389;
wire v_32390;
wire v_32391;
wire v_32392;
wire v_32393;
wire v_32394;
wire v_32395;
wire v_32396;
wire v_32397;
wire v_32398;
wire v_32399;
wire v_32400;
wire v_32401;
wire v_32402;
wire v_32403;
wire v_32404;
wire v_32405;
wire v_32406;
wire v_32407;
wire v_32408;
wire v_32409;
wire v_32410;
wire v_32411;
wire v_32412;
wire v_32413;
wire v_32414;
wire v_32415;
wire v_32416;
wire v_32417;
wire v_32418;
wire v_32419;
wire v_32420;
wire v_32421;
wire v_32422;
wire v_32423;
wire v_32424;
wire v_32425;
wire v_32426;
wire v_32427;
wire v_32428;
wire v_32429;
wire v_32430;
wire v_32431;
wire v_32432;
wire v_32433;
wire v_32434;
wire v_32435;
wire v_32436;
wire v_32437;
wire v_32438;
wire v_32439;
wire v_32440;
wire v_32441;
wire v_32442;
wire v_32443;
wire v_32444;
wire v_32445;
wire v_32446;
wire v_32447;
wire v_32448;
wire v_32449;
wire v_32450;
wire v_32451;
wire v_32452;
wire v_32453;
wire v_32454;
wire v_32455;
wire v_32456;
wire v_32457;
wire v_32458;
wire v_32459;
wire v_32460;
wire v_32461;
wire v_32462;
wire v_32463;
wire v_32464;
wire v_32465;
wire v_32466;
wire v_32467;
wire v_32468;
wire v_32469;
wire v_32470;
wire v_32471;
wire v_32472;
wire v_32473;
wire v_32474;
wire v_32475;
wire v_32476;
wire v_32477;
wire v_32478;
wire v_32479;
wire v_32480;
wire v_32481;
wire v_32482;
wire v_32483;
wire v_32484;
wire v_32485;
wire v_32486;
wire v_32487;
wire v_32488;
wire v_32489;
wire v_32490;
wire v_32491;
wire v_32492;
wire v_32493;
wire v_32494;
wire v_32495;
wire v_32496;
wire v_32497;
wire v_32498;
wire v_32499;
wire v_32500;
wire v_32501;
wire v_32502;
wire v_32503;
wire v_32504;
wire v_32505;
wire v_32506;
wire v_32507;
wire v_32508;
wire v_32509;
wire v_32510;
wire v_32511;
wire v_32512;
wire v_32513;
wire v_32514;
wire v_32515;
wire v_32516;
wire v_32517;
wire v_32518;
wire v_32519;
wire v_32520;
wire v_32521;
wire v_32522;
wire v_32523;
wire v_32524;
wire v_32525;
wire v_32526;
wire v_32527;
wire v_32528;
wire v_32529;
wire v_32530;
wire v_32531;
wire v_32532;
wire v_32533;
wire v_32534;
wire v_32535;
wire v_32536;
wire v_32537;
wire v_32538;
wire v_32539;
wire v_32540;
wire v_32541;
wire v_32542;
wire v_32543;
wire v_32544;
wire v_32545;
wire v_32546;
wire v_32547;
wire v_32548;
wire v_32549;
wire v_32550;
wire v_32551;
wire v_32552;
wire v_32553;
wire v_32554;
wire v_32555;
wire v_32556;
wire v_32557;
wire v_32558;
wire v_32559;
wire v_32560;
wire v_32561;
wire v_32562;
wire v_32563;
wire v_32564;
wire v_32565;
wire v_32566;
wire v_32567;
wire v_32568;
wire v_32569;
wire v_32570;
wire v_32571;
wire v_32572;
wire v_32573;
wire v_32574;
wire v_32575;
wire v_32576;
wire v_32577;
wire v_32578;
wire v_32579;
wire v_32580;
wire v_32581;
wire v_32582;
wire v_32583;
wire v_32584;
wire v_32585;
wire v_32586;
wire v_32587;
wire v_32588;
wire v_32589;
wire v_32590;
wire v_32591;
wire v_32592;
wire v_32593;
wire v_32594;
wire v_32595;
wire v_32596;
wire v_32597;
wire v_32598;
wire v_32599;
wire v_32600;
wire v_32601;
wire v_32602;
wire v_32603;
wire v_32604;
wire v_32605;
wire v_32606;
wire v_32607;
wire v_32608;
wire v_32609;
wire v_32610;
wire v_32611;
wire v_32612;
wire v_32613;
wire v_32614;
wire v_32615;
wire v_32616;
wire v_32617;
wire v_32618;
wire v_32619;
wire v_32620;
wire v_32621;
wire v_32622;
wire v_32623;
wire v_32624;
wire v_32625;
wire v_32626;
wire v_32627;
wire v_32628;
wire v_32629;
wire v_32630;
wire v_32631;
wire v_32632;
wire v_32633;
wire v_32634;
wire v_32635;
wire v_32636;
wire v_32637;
wire v_32638;
wire v_32639;
wire v_32640;
wire v_32641;
wire v_32642;
wire v_32643;
wire v_32644;
wire v_32645;
wire v_32646;
wire v_32647;
wire v_32648;
wire v_32649;
wire v_32650;
wire v_32651;
wire v_32652;
wire v_32653;
wire v_32654;
wire v_32655;
wire v_32656;
wire v_32657;
wire v_32658;
wire v_32659;
wire v_32660;
wire v_32661;
wire v_32662;
wire v_32663;
wire v_32664;
wire v_32665;
wire v_32666;
wire v_32667;
wire v_32668;
wire v_32669;
wire v_32670;
wire v_32671;
wire v_32672;
wire v_32673;
wire v_32674;
wire v_32675;
wire v_32676;
wire v_32677;
wire v_32678;
wire v_32679;
wire v_32680;
wire v_32681;
wire v_32682;
wire v_32683;
wire v_32684;
wire v_32685;
wire v_32686;
wire v_32687;
wire v_32688;
wire v_32689;
wire v_32690;
wire v_32691;
wire v_32692;
wire v_32693;
wire v_32694;
wire v_32695;
wire v_32696;
wire v_32697;
wire v_32698;
wire v_32699;
wire v_32700;
wire v_32701;
wire v_32702;
wire v_32703;
wire v_32704;
wire v_32705;
wire v_32706;
wire v_32707;
wire v_32708;
wire v_32709;
wire v_32710;
wire v_32711;
wire v_32712;
wire v_32713;
wire v_32714;
wire v_32715;
wire v_32716;
wire v_32717;
wire v_32718;
wire v_32719;
wire v_32720;
wire v_32721;
wire v_32722;
wire v_32723;
wire v_32724;
wire v_32725;
wire v_32726;
wire v_32727;
wire v_32728;
wire v_32729;
wire v_32730;
wire v_32731;
wire v_32732;
wire v_32733;
wire v_32734;
wire v_32735;
wire v_32736;
wire v_32737;
wire v_32738;
wire v_32739;
wire v_32740;
wire v_32741;
wire v_32742;
wire v_32743;
wire v_32744;
wire v_32745;
wire v_32746;
wire v_32747;
wire v_32748;
wire v_32749;
wire v_32750;
wire v_32751;
wire v_32752;
wire v_32753;
wire v_32754;
wire v_32755;
wire v_32756;
wire v_32757;
wire v_32758;
wire v_32759;
wire v_32760;
wire v_32761;
wire v_32762;
wire v_32763;
wire v_32764;
wire v_32765;
wire v_32766;
wire v_32767;
wire v_32768;
wire v_32769;
wire v_32770;
wire v_32771;
wire v_32772;
wire v_32773;
wire v_32774;
wire v_32775;
wire v_32776;
wire v_32777;
wire v_32778;
wire v_32779;
wire v_32780;
wire v_32781;
wire v_32782;
wire v_32783;
wire v_32784;
wire v_32785;
wire v_32786;
wire v_32787;
wire v_32788;
wire v_32789;
wire v_32790;
wire v_32791;
wire v_32792;
wire v_32793;
wire v_32794;
wire v_32795;
wire v_32796;
wire v_32797;
wire v_32798;
wire v_32799;
wire v_32800;
wire v_32801;
wire v_32802;
wire v_32803;
wire v_32804;
wire v_32805;
wire v_32806;
wire v_32807;
wire v_32808;
wire v_32809;
wire v_32810;
wire v_32811;
wire v_32812;
wire v_32813;
wire v_32814;
wire v_32815;
wire v_32816;
wire v_32817;
wire v_32818;
wire v_32819;
wire v_32820;
wire v_32821;
wire v_32822;
wire v_32823;
wire v_32824;
wire v_32825;
wire v_32826;
wire v_32827;
wire v_32828;
wire v_32829;
wire v_32830;
wire v_32831;
wire v_32832;
wire v_32833;
wire v_32834;
wire v_32835;
wire v_32836;
wire v_32837;
wire v_32838;
wire v_32839;
wire v_32840;
wire v_32841;
wire v_32842;
wire v_32843;
wire v_32844;
wire v_32845;
wire v_32846;
wire v_32847;
wire v_32848;
wire v_32849;
wire v_32850;
wire v_32851;
wire v_32852;
wire v_32853;
wire v_32854;
wire v_32855;
wire v_32856;
wire v_32857;
wire v_32858;
wire v_32859;
wire v_32860;
wire v_32861;
wire v_32862;
wire v_32863;
wire v_32864;
wire v_32865;
wire v_32866;
wire v_32867;
wire v_32868;
wire v_32869;
wire v_32870;
wire v_32871;
wire v_32872;
wire v_32873;
wire v_32874;
wire v_32875;
wire v_32876;
wire v_32877;
wire v_32878;
wire v_32879;
wire v_32880;
wire v_32881;
wire v_32882;
wire v_32883;
wire v_32884;
wire v_32885;
wire v_32886;
wire v_32887;
wire v_32888;
wire v_32889;
wire v_32890;
wire v_32891;
wire v_32892;
wire v_32893;
wire v_32894;
wire v_32895;
wire v_32896;
wire v_32897;
wire v_32898;
wire v_32899;
wire v_32900;
wire v_32901;
wire v_32902;
wire v_32903;
wire v_32904;
wire v_32905;
wire v_32906;
wire v_32907;
wire v_32908;
wire v_32909;
wire v_32910;
wire v_32911;
wire v_32912;
wire v_32913;
wire v_32914;
wire v_32915;
wire v_32916;
wire v_32917;
wire v_32918;
wire v_32919;
wire v_32920;
wire v_32921;
wire v_32922;
wire v_32923;
wire v_32924;
wire v_32925;
wire v_32926;
wire v_32927;
wire v_32928;
wire v_32929;
wire v_32930;
wire v_32931;
wire v_32932;
wire v_32933;
wire v_32934;
wire v_32935;
wire v_32936;
wire v_32937;
wire v_32938;
wire v_32939;
wire v_32940;
wire v_32941;
wire v_32942;
wire v_32943;
wire v_32944;
wire v_32945;
wire v_32946;
wire v_32947;
wire v_32948;
wire v_32949;
wire v_32950;
wire v_32951;
wire v_32952;
wire v_32953;
wire v_32954;
wire v_32955;
wire v_32956;
wire v_32957;
wire v_32958;
wire v_32959;
wire v_32960;
wire v_32961;
wire v_32962;
wire v_32963;
wire v_32964;
wire v_32965;
wire v_32966;
wire v_32967;
wire v_32968;
wire v_32969;
wire v_32970;
wire v_32971;
wire v_32972;
wire v_32973;
wire v_32974;
wire v_32975;
wire v_32976;
wire v_32977;
wire v_32978;
wire v_32979;
wire v_32980;
wire v_32981;
wire v_32982;
wire v_32983;
wire v_32984;
wire v_32985;
wire v_32986;
wire v_32987;
wire v_32988;
wire v_32989;
wire v_32990;
wire v_32991;
wire v_32992;
wire v_32993;
wire v_32994;
wire v_32995;
wire v_32996;
wire v_32997;
wire v_32998;
wire v_32999;
wire v_33000;
wire v_33001;
wire v_33002;
wire v_33003;
wire v_33004;
wire v_33005;
wire v_33006;
wire v_33007;
wire v_33008;
wire v_33009;
wire v_33010;
wire v_33011;
wire v_33012;
wire v_33013;
wire v_33014;
wire v_33015;
wire v_33016;
wire v_33017;
wire v_33018;
wire v_33019;
wire v_33020;
wire v_33021;
wire v_33022;
wire v_33023;
wire v_33024;
wire v_33025;
wire v_33026;
wire v_33027;
wire v_33028;
wire v_33029;
wire v_33030;
wire v_33031;
wire v_33032;
wire v_33033;
wire v_33034;
wire v_33035;
wire v_33036;
wire v_33037;
wire v_33038;
wire v_33039;
wire v_33040;
wire v_33041;
wire v_33042;
wire v_33043;
wire v_33044;
wire v_33045;
wire v_33046;
wire v_33047;
wire v_33048;
wire v_33049;
wire v_33050;
wire v_33051;
wire v_33052;
wire v_33053;
wire v_33054;
wire v_33055;
wire v_33056;
wire v_33057;
wire v_33058;
wire v_33059;
wire v_33060;
wire v_33061;
wire v_33062;
wire v_33063;
wire v_33064;
wire v_33065;
wire v_33066;
wire v_33067;
wire v_33068;
wire v_33069;
wire v_33070;
wire v_33071;
wire v_33072;
wire v_33073;
wire v_33074;
wire v_33075;
wire v_33076;
wire v_33077;
wire v_33078;
wire v_33079;
wire v_33080;
wire v_33081;
wire v_33082;
wire v_33083;
wire v_33084;
wire v_33085;
wire v_33086;
wire v_33087;
wire v_33088;
wire v_33089;
wire v_33090;
wire v_33091;
wire v_33092;
wire v_33093;
wire v_33094;
wire v_33095;
wire v_33096;
wire v_33097;
wire v_33098;
wire v_33099;
wire v_33100;
wire v_33101;
wire v_33102;
wire v_33103;
wire v_33104;
wire v_33105;
wire v_33106;
wire v_33107;
wire v_33108;
wire v_33109;
wire v_33110;
wire v_33111;
wire v_33112;
wire v_33113;
wire v_33114;
wire v_33115;
wire v_33116;
wire v_33117;
wire v_33118;
wire v_33119;
wire v_33120;
wire v_33121;
wire v_33122;
wire v_33123;
wire v_33124;
wire v_33125;
wire v_33126;
wire v_33127;
wire v_33128;
wire v_33129;
wire v_33130;
wire v_33131;
wire v_33132;
wire v_33133;
wire v_33134;
wire v_33135;
wire v_33136;
wire v_33137;
wire v_33138;
wire v_33139;
wire v_33140;
wire v_33141;
wire v_33142;
wire v_33143;
wire v_33144;
wire v_33145;
wire v_33146;
wire v_33147;
wire v_33148;
wire v_33149;
wire v_33150;
wire v_33151;
wire v_33152;
wire v_33153;
wire v_33154;
wire v_33155;
wire v_33156;
wire v_33157;
wire v_33158;
wire v_33159;
wire v_33160;
wire v_33161;
wire v_33162;
wire v_33163;
wire v_33164;
wire v_33165;
wire v_33166;
wire v_33167;
wire v_33168;
wire v_33169;
wire v_33170;
wire v_33171;
wire v_33172;
wire v_33173;
wire v_33174;
wire v_33175;
wire v_33176;
wire v_33177;
wire v_33178;
wire v_33179;
wire v_33180;
wire v_33181;
wire v_33182;
wire v_33183;
wire v_33184;
wire v_33185;
wire v_33186;
wire v_33187;
wire v_33188;
wire v_33189;
wire v_33190;
wire v_33191;
wire v_33192;
wire v_33193;
wire v_33194;
wire v_33195;
wire v_33196;
wire v_33197;
wire v_33198;
wire v_33199;
wire v_33200;
wire v_33201;
wire v_33202;
wire v_33203;
wire v_33204;
wire v_33205;
wire v_33206;
wire v_33207;
wire v_33208;
wire v_33209;
wire v_33210;
wire v_33211;
wire v_33212;
wire v_33213;
wire v_33214;
wire v_33215;
wire v_33216;
wire v_33217;
wire v_33218;
wire v_33219;
wire v_33220;
wire v_33221;
wire v_33222;
wire v_33223;
wire v_33224;
wire v_33225;
wire v_33226;
wire v_33227;
wire v_33228;
wire v_33229;
wire v_33230;
wire v_33231;
wire v_33232;
wire v_33233;
wire v_33234;
wire v_33235;
wire v_33236;
wire v_33237;
wire v_33238;
wire v_33239;
wire v_33240;
wire v_33241;
wire v_33242;
wire v_33243;
wire v_33244;
wire v_33245;
wire v_33246;
wire v_33247;
wire v_33248;
wire v_33249;
wire v_33250;
wire v_33251;
wire v_33252;
wire v_33253;
wire v_33254;
wire v_33255;
wire v_33256;
wire v_33257;
wire v_33258;
wire v_33259;
wire v_33260;
wire v_33261;
wire v_33262;
wire v_33263;
wire v_33264;
wire v_33265;
wire v_33266;
wire v_33267;
wire v_33268;
wire v_33269;
wire v_33270;
wire v_33271;
wire v_33272;
wire v_33273;
wire v_33274;
wire v_33275;
wire v_33276;
wire v_33277;
wire v_33278;
wire v_33279;
wire v_33280;
wire v_33281;
wire v_33282;
wire v_33283;
wire v_33284;
wire v_33285;
wire v_33286;
wire v_33287;
wire v_33288;
wire v_33289;
wire v_33290;
wire v_33291;
wire v_33292;
wire v_33293;
wire v_33294;
wire v_33295;
wire v_33296;
wire v_33297;
wire v_33298;
wire v_33299;
wire v_33300;
wire v_33301;
wire v_33302;
wire v_33303;
wire v_33304;
wire v_33305;
wire v_33306;
wire v_33307;
wire v_33308;
wire v_33309;
wire v_33310;
wire v_33311;
wire v_33312;
wire v_33313;
wire v_33314;
wire v_33315;
wire v_33316;
wire v_33317;
wire v_33318;
wire v_33319;
wire v_33320;
wire v_33321;
wire v_33322;
wire v_33323;
wire v_33324;
wire v_33325;
wire v_33326;
wire v_33327;
wire v_33328;
wire v_33329;
wire v_33330;
wire v_33331;
wire v_33332;
wire v_33333;
wire v_33334;
wire v_33335;
wire v_33336;
wire v_33337;
wire v_33338;
wire v_33339;
wire v_33340;
wire v_33341;
wire v_33342;
wire v_33343;
wire v_33344;
wire v_33345;
wire v_33346;
wire v_33347;
wire v_33348;
wire v_33349;
wire v_33350;
wire v_33351;
wire v_33352;
wire v_33353;
wire v_33354;
wire v_33355;
wire v_33356;
wire v_33357;
wire v_33358;
wire v_33359;
wire v_33360;
wire v_33361;
wire v_33362;
wire v_33363;
wire v_33364;
wire v_33365;
wire v_33366;
wire v_33367;
wire v_33368;
wire v_33369;
wire v_33370;
wire v_33371;
wire v_33372;
wire v_33373;
wire v_33374;
wire v_33375;
wire v_33376;
wire v_33377;
wire v_33378;
wire v_33379;
wire v_33380;
wire v_33381;
wire v_33382;
wire v_33383;
wire v_33384;
wire v_33385;
wire v_33386;
wire v_33387;
wire v_33388;
wire v_33389;
wire v_33390;
wire v_33391;
wire v_33392;
wire v_33393;
wire v_33394;
wire v_33395;
wire v_33396;
wire v_33397;
wire v_33398;
wire v_33399;
wire v_33400;
wire v_33401;
wire v_33402;
wire v_33403;
wire v_33404;
wire v_33405;
wire v_33406;
wire v_33407;
wire v_33408;
wire v_33409;
wire v_33410;
wire v_33411;
wire v_33412;
wire v_33413;
wire v_33414;
wire v_33415;
wire v_33416;
wire v_33417;
wire v_33418;
wire v_33419;
wire v_33420;
wire v_33421;
wire v_33422;
wire v_33423;
wire v_33424;
wire v_33425;
wire v_33426;
wire v_33427;
wire v_33428;
wire v_33429;
wire v_33430;
wire v_33431;
wire v_33432;
wire v_33433;
wire v_33434;
wire v_33435;
wire v_33436;
wire v_33437;
wire v_33438;
wire v_33439;
wire v_33440;
wire v_33441;
wire v_33442;
wire v_33443;
wire v_33444;
wire v_33445;
wire v_33446;
wire v_33447;
wire v_33448;
wire v_33449;
wire v_33450;
wire v_33451;
wire v_33452;
wire v_33453;
wire v_33454;
wire v_33455;
wire v_33456;
wire v_33457;
wire v_33458;
wire v_33459;
wire v_33460;
wire v_33461;
wire v_33462;
wire v_33463;
wire v_33464;
wire v_33465;
wire v_33466;
wire v_33467;
wire v_33468;
wire v_33469;
wire v_33470;
wire v_33471;
wire v_33472;
wire v_33473;
wire v_33474;
wire v_33475;
wire v_33476;
wire v_33477;
wire v_33478;
wire v_33479;
wire v_33480;
wire v_33481;
wire v_33482;
wire v_33483;
wire v_33484;
wire v_33485;
wire v_33486;
wire v_33487;
wire v_33488;
wire v_33489;
wire v_33490;
wire v_33491;
wire v_33492;
wire v_33493;
wire v_33494;
wire v_33495;
wire v_33496;
wire v_33497;
wire v_33498;
wire v_33499;
wire v_33500;
wire v_33501;
wire v_33502;
wire v_33503;
wire v_33504;
wire v_33505;
wire v_33506;
wire v_33507;
wire v_33508;
wire v_33509;
wire v_33510;
wire v_33511;
wire v_33512;
wire v_33513;
wire v_33514;
wire v_33515;
wire v_33516;
wire v_33517;
wire v_33518;
wire v_33519;
wire v_33520;
wire v_33521;
wire v_33522;
wire v_33523;
wire v_33524;
wire v_33525;
wire v_33526;
wire v_33527;
wire v_33528;
wire v_33529;
wire v_33530;
wire v_33531;
wire v_33532;
wire v_33533;
wire v_33534;
wire v_33535;
wire v_33536;
wire v_33537;
wire v_33538;
wire v_33539;
wire v_33540;
wire v_33541;
wire v_33542;
wire v_33543;
wire v_33544;
wire v_33545;
wire v_33546;
wire v_33547;
wire v_33548;
wire v_33549;
wire v_33550;
wire v_33551;
wire v_33552;
wire v_33553;
wire v_33554;
wire v_33555;
wire v_33556;
wire v_33557;
wire v_33558;
wire v_33559;
wire v_33560;
wire v_33561;
wire v_33562;
wire v_33563;
wire v_33564;
wire v_33565;
wire v_33566;
wire v_33567;
wire v_33568;
wire v_33569;
wire v_33570;
wire v_33571;
wire v_33572;
wire v_33573;
wire v_33574;
wire v_33575;
wire v_33576;
wire v_33577;
wire v_33578;
wire v_33579;
wire v_33580;
wire v_33581;
wire v_33582;
wire v_33583;
wire v_33584;
wire v_33585;
wire v_33586;
wire v_33587;
wire v_33588;
wire v_33589;
wire v_33590;
wire v_33591;
wire v_33592;
wire v_33593;
wire v_33594;
wire v_33595;
wire v_33596;
wire v_33597;
wire v_33598;
wire v_33599;
wire v_33600;
wire v_33601;
wire v_33602;
wire v_33603;
wire v_33604;
wire v_33605;
wire v_33606;
wire v_33607;
wire v_33608;
wire v_33609;
wire v_33610;
wire v_33611;
wire v_33612;
wire v_33613;
wire v_33614;
wire v_33615;
wire v_33616;
wire v_33617;
wire v_33618;
wire v_33619;
wire v_33620;
wire v_33621;
wire v_33622;
wire v_33623;
wire v_33624;
wire v_33625;
wire v_33626;
wire v_33627;
wire v_33628;
wire v_33629;
wire v_33630;
wire v_33631;
wire v_33632;
wire v_33633;
wire v_33634;
wire v_33635;
wire v_33636;
wire v_33637;
wire v_33638;
wire v_33639;
wire v_33640;
wire v_33641;
wire v_33642;
wire v_33643;
wire v_33644;
wire v_33645;
wire v_33646;
wire v_33647;
wire v_33648;
wire v_33649;
wire v_33650;
wire v_33651;
wire v_33652;
wire v_33653;
wire v_33654;
wire v_33655;
wire v_33656;
wire v_33657;
wire v_33658;
wire v_33659;
wire v_33660;
wire v_33661;
wire v_33662;
wire v_33663;
wire v_33664;
wire v_33665;
wire v_33666;
wire v_33667;
wire v_33668;
wire v_33669;
wire v_33670;
wire v_33671;
wire v_33672;
wire v_33673;
wire v_33674;
wire v_33675;
wire v_33676;
wire v_33677;
wire v_33678;
wire v_33679;
wire v_33680;
wire v_33681;
wire v_33682;
wire v_33683;
wire v_33684;
wire v_33685;
wire v_33686;
wire v_33687;
wire v_33688;
wire v_33689;
wire v_33690;
wire v_33691;
wire v_33692;
wire v_33693;
wire v_33694;
wire v_33695;
wire v_33696;
wire v_33697;
wire v_33698;
wire v_33699;
wire v_33700;
wire v_33701;
wire v_33702;
wire v_33703;
wire v_33704;
wire v_33705;
wire v_33706;
wire v_33707;
wire v_33708;
wire v_33709;
wire v_33710;
wire v_33711;
wire v_33712;
wire v_33713;
wire v_33714;
wire v_33715;
wire v_33716;
wire v_33717;
wire v_33718;
wire v_33719;
wire v_33720;
wire v_33721;
wire v_33722;
wire v_33723;
wire v_33724;
wire v_33725;
wire v_33726;
wire v_33727;
wire v_33728;
wire v_33729;
wire v_33730;
wire v_33731;
wire v_33732;
wire v_33733;
wire v_33734;
wire v_33735;
wire v_33736;
wire v_33737;
wire v_33738;
wire v_33739;
wire v_33740;
wire v_33741;
wire v_33742;
wire v_33743;
wire v_33744;
wire v_33745;
wire v_33746;
wire v_33747;
wire v_33748;
wire v_33749;
wire v_33750;
wire v_33751;
wire v_33752;
wire v_33753;
wire v_33754;
wire v_33755;
wire v_33756;
wire v_33757;
wire v_33758;
wire v_33759;
wire v_33760;
wire v_33761;
wire v_33762;
wire v_33763;
wire v_33764;
wire v_33765;
wire v_33766;
wire v_33767;
wire v_33768;
wire v_33769;
wire v_33770;
wire v_33771;
wire v_33772;
wire v_33773;
wire v_33774;
wire v_33775;
wire v_33776;
wire v_33777;
wire v_33778;
wire v_33779;
wire v_33780;
wire v_33781;
wire v_33782;
wire v_33783;
wire v_33784;
wire v_33785;
wire v_33786;
wire v_33787;
wire v_33788;
wire v_33789;
wire v_33790;
wire v_33791;
wire v_33792;
wire v_33793;
wire v_33794;
wire v_33795;
wire v_33796;
wire v_33797;
wire v_33798;
wire v_33799;
wire v_33800;
wire v_33801;
wire v_33802;
wire v_33803;
wire v_33804;
wire v_33805;
wire v_33806;
wire v_33807;
wire v_33808;
wire v_33809;
wire v_33810;
wire v_33811;
wire v_33812;
wire v_33813;
wire v_33814;
wire v_33815;
wire v_33816;
wire v_33817;
wire v_33818;
wire v_33819;
wire v_33820;
wire v_33821;
wire v_33822;
wire v_33823;
wire v_33824;
wire v_33825;
wire v_33826;
wire v_33827;
wire v_33828;
wire v_33829;
wire v_33830;
wire v_33831;
wire v_33832;
wire v_33833;
wire v_33834;
wire v_33835;
wire v_33836;
wire v_33837;
wire v_33838;
wire v_33839;
wire v_33840;
wire v_33841;
wire v_33842;
wire v_33843;
wire v_33844;
wire v_33845;
wire v_33846;
wire v_33847;
wire v_33848;
wire v_33849;
wire v_33850;
wire v_33851;
wire v_33852;
wire v_33853;
wire v_33854;
wire v_33855;
wire v_33856;
wire v_33857;
wire v_33858;
wire v_33859;
wire v_33860;
wire v_33861;
wire v_33862;
wire v_33863;
wire v_33864;
wire v_33865;
wire v_33866;
wire v_33867;
wire v_33868;
wire v_33869;
wire v_33870;
wire v_33871;
wire v_33872;
wire v_33873;
wire v_33874;
wire v_33875;
wire v_33876;
wire v_33877;
wire v_33878;
wire v_33879;
wire v_33880;
wire v_33881;
wire v_33882;
wire v_33883;
wire v_33884;
wire v_33885;
wire v_33886;
wire v_33887;
wire v_33888;
wire v_33889;
wire v_33890;
wire v_33891;
wire v_33892;
wire v_33893;
wire v_33894;
wire v_33895;
wire v_33896;
wire v_33897;
wire v_33898;
wire v_33899;
wire v_33900;
wire v_33901;
wire v_33902;
wire v_33903;
wire v_33904;
wire v_33905;
wire v_33906;
wire v_33907;
wire v_33908;
wire v_33909;
wire v_33910;
wire v_33911;
wire v_33912;
wire v_33913;
wire v_33914;
wire v_33915;
wire v_33916;
wire v_33917;
wire v_33918;
wire v_33919;
wire v_33920;
wire v_33921;
wire v_33922;
wire v_33923;
wire v_33924;
wire v_33925;
wire v_33926;
wire v_33927;
wire v_33928;
wire v_33929;
wire v_33930;
wire v_33931;
wire v_33932;
wire v_33933;
wire v_33934;
wire v_33935;
wire v_33936;
wire v_33937;
wire v_33938;
wire v_33939;
wire v_33940;
wire v_33941;
wire v_33942;
wire v_33943;
wire v_33944;
wire v_33945;
wire v_33946;
wire v_33947;
wire v_33948;
wire v_33949;
wire v_33950;
wire v_33951;
wire v_33952;
wire v_33953;
wire v_33954;
wire v_33955;
wire v_33956;
wire v_33957;
wire v_33958;
wire v_33959;
wire v_33960;
wire v_33961;
wire v_33962;
wire v_33963;
wire v_33964;
wire v_33965;
wire v_33966;
wire v_33967;
wire v_33968;
wire v_33969;
wire v_33970;
wire v_33971;
wire v_33972;
wire v_33973;
wire v_33974;
wire v_33975;
wire v_33976;
wire v_33977;
wire v_33978;
wire v_33979;
wire v_33980;
wire v_33981;
wire v_33982;
wire v_33983;
wire v_33984;
wire v_33985;
wire v_33986;
wire v_33987;
wire v_33988;
wire v_33989;
wire v_33990;
wire v_33991;
wire v_33992;
wire v_33993;
wire v_33994;
wire v_33995;
wire v_33996;
wire v_33997;
wire v_33998;
wire v_33999;
wire v_34000;
wire v_34001;
wire v_34002;
wire v_34003;
wire v_34004;
wire v_34005;
wire v_34006;
wire v_34007;
wire v_34008;
wire v_34009;
wire v_34010;
wire v_34011;
wire v_34012;
wire v_34013;
wire v_34014;
wire v_34015;
wire v_34016;
wire v_34017;
wire v_34018;
wire v_34019;
wire v_34020;
wire v_34021;
wire v_34022;
wire v_34023;
wire v_34024;
wire v_34025;
wire v_34026;
wire v_34027;
wire v_34028;
wire v_34029;
wire v_34030;
wire v_34031;
wire v_34032;
wire v_34033;
wire v_34034;
wire v_34035;
wire v_34036;
wire v_34037;
wire v_34038;
wire v_34039;
wire v_34040;
wire v_34041;
wire v_34042;
wire v_34043;
wire v_34044;
wire v_34045;
wire v_34046;
wire v_34047;
wire v_34048;
wire v_34049;
wire v_34050;
wire v_34051;
wire v_34052;
wire v_34053;
wire v_34054;
wire v_34055;
wire v_34056;
wire v_34057;
wire v_34058;
wire v_34059;
wire v_34060;
wire v_34061;
wire v_34062;
wire v_34063;
wire v_34064;
wire v_34065;
wire v_34066;
wire v_34067;
wire v_34068;
wire v_34069;
wire v_34070;
wire v_34071;
wire v_34072;
wire v_34073;
wire v_34074;
wire v_34075;
wire v_34076;
wire v_34077;
wire v_34078;
wire v_34079;
wire v_34080;
wire v_34081;
wire v_34082;
wire v_34083;
wire v_34084;
wire v_34085;
wire v_34086;
wire v_34087;
wire v_34088;
wire v_34089;
wire v_34090;
wire v_34091;
wire v_34092;
wire v_34093;
wire v_34094;
wire v_34095;
wire v_34096;
wire v_34097;
wire v_34098;
wire v_34099;
wire v_34100;
wire v_34101;
wire v_34102;
wire v_34103;
wire v_34104;
wire v_34105;
wire v_34106;
wire v_34107;
wire v_34108;
wire v_34109;
wire v_34110;
wire v_34111;
wire v_34112;
wire v_34113;
wire v_34114;
wire v_34115;
wire v_34116;
wire v_34117;
wire v_34118;
wire v_34119;
wire v_34120;
wire v_34121;
wire v_34122;
wire v_34123;
wire v_34124;
wire v_34125;
wire v_34126;
wire v_34127;
wire v_34128;
wire v_34129;
wire v_34130;
wire v_34131;
wire v_34132;
wire v_34133;
wire v_34134;
wire v_34135;
wire v_34136;
wire v_34137;
wire v_34138;
wire v_34139;
wire v_34140;
wire v_34141;
wire v_34142;
wire v_34143;
wire v_34144;
wire v_34145;
wire v_34146;
wire v_34147;
wire v_34148;
wire v_34149;
wire v_34150;
wire v_34151;
wire v_34152;
wire v_34153;
wire v_34154;
wire v_34155;
wire v_34156;
wire v_34157;
wire v_34158;
wire v_34159;
wire v_34160;
wire v_34161;
wire v_34162;
wire v_34163;
wire v_34164;
wire v_34165;
wire v_34166;
wire v_34167;
wire v_34168;
wire v_34169;
wire v_34170;
wire v_34171;
wire v_34172;
wire v_34173;
wire v_34174;
wire v_34175;
wire v_34176;
wire v_34177;
wire v_34178;
wire v_34179;
wire v_34180;
wire v_34181;
wire v_34182;
wire v_34183;
wire v_34184;
wire v_34185;
wire v_34186;
wire v_34187;
wire v_34188;
wire v_34189;
wire v_34190;
wire v_34191;
wire v_34192;
wire v_34193;
wire v_34194;
wire v_34195;
wire v_34196;
wire v_34197;
wire v_34198;
wire v_34199;
wire v_34200;
wire v_34201;
wire v_34202;
wire v_34203;
wire v_34204;
wire v_34205;
wire v_34206;
wire v_34207;
wire v_34208;
wire v_34209;
wire v_34210;
wire v_34211;
wire v_34212;
wire v_34213;
wire v_34214;
wire v_34215;
wire v_34216;
wire v_34217;
wire v_34218;
wire v_34219;
wire v_34220;
wire v_34221;
wire v_34222;
wire v_34223;
wire v_34224;
wire v_34225;
wire v_34226;
wire v_34227;
wire v_34228;
wire v_34229;
wire v_34230;
wire v_34231;
wire v_34232;
wire v_34233;
wire v_34234;
wire v_34235;
wire v_34236;
wire v_34237;
wire v_34238;
wire v_34239;
wire v_34240;
wire v_34241;
wire v_34242;
wire v_34243;
wire v_34244;
wire v_34245;
wire v_34246;
wire v_34247;
wire v_34248;
wire v_34249;
wire v_34250;
wire v_34251;
wire v_34252;
wire v_34253;
wire v_34254;
wire v_34255;
wire v_34256;
wire v_34257;
wire v_34258;
wire v_34259;
wire v_34260;
wire v_34261;
wire v_34262;
wire v_34263;
wire v_34264;
wire v_34265;
wire v_34266;
wire v_34267;
wire v_34268;
wire v_34269;
wire v_34270;
wire v_34271;
wire v_34272;
wire v_34273;
wire v_34274;
wire v_34275;
wire v_34276;
wire v_34277;
wire v_34278;
wire v_34279;
wire v_34280;
wire v_34281;
wire v_34282;
wire v_34283;
wire v_34284;
wire v_34285;
wire v_34286;
wire v_34287;
wire v_34288;
wire v_34289;
wire v_34290;
wire v_34291;
wire v_34292;
wire v_34293;
wire v_34294;
wire v_34295;
wire v_34296;
wire v_34297;
wire v_34298;
wire v_34299;
wire v_34300;
wire v_34301;
wire v_34302;
wire v_34303;
wire v_34304;
wire v_34305;
wire v_34306;
wire v_34307;
wire v_34308;
wire v_34309;
wire v_34310;
wire v_34311;
wire v_34312;
wire v_34313;
wire v_34314;
wire v_34315;
wire v_34316;
wire v_34317;
wire v_34318;
wire v_34319;
wire v_34320;
wire v_34321;
wire v_34322;
wire v_34323;
wire v_34324;
wire v_34325;
wire v_34326;
wire v_34327;
wire v_34328;
wire v_34329;
wire v_34330;
wire v_34331;
wire v_34332;
wire v_34333;
wire v_34334;
wire v_34335;
wire v_34336;
wire v_34337;
wire v_34338;
wire v_34339;
wire v_34340;
wire v_34341;
wire v_34342;
wire v_34343;
wire v_34344;
wire v_34345;
wire v_34346;
wire v_34347;
wire v_34348;
wire v_34349;
wire v_34350;
wire v_34351;
wire v_34352;
wire v_34353;
wire v_34354;
wire v_34355;
wire v_34356;
wire v_34357;
wire v_34358;
wire v_34359;
wire v_34360;
wire v_34361;
wire v_34362;
wire v_34363;
wire v_34364;
wire v_34365;
wire v_34366;
wire v_34367;
wire v_34368;
wire v_34369;
wire v_34370;
wire v_34371;
wire v_34372;
wire v_34373;
wire v_34374;
wire v_34375;
wire v_34376;
wire v_34377;
wire v_34378;
wire v_34379;
wire v_34380;
wire v_34381;
wire v_34382;
wire v_34383;
wire v_34384;
wire v_34385;
wire v_34386;
wire v_34387;
wire v_34388;
wire v_34389;
wire v_34390;
wire v_34391;
wire v_34392;
wire v_34393;
wire v_34394;
wire v_34395;
wire v_34396;
wire v_34397;
wire v_34398;
wire v_34399;
wire v_34400;
wire v_34401;
wire v_34402;
wire v_34403;
wire v_34404;
wire v_34405;
wire v_34406;
wire v_34407;
wire v_34408;
wire v_34409;
wire v_34410;
wire v_34411;
wire v_34412;
wire v_34413;
wire v_34414;
wire v_34415;
wire v_34416;
wire v_34417;
wire v_34418;
wire v_34419;
wire v_34420;
wire v_34421;
wire v_34422;
wire v_34423;
wire v_34424;
wire v_34425;
wire v_34426;
wire v_34427;
wire v_34428;
wire v_34429;
wire v_34430;
wire v_34431;
wire v_34432;
wire v_34433;
wire v_34434;
wire v_34435;
wire v_34436;
wire v_34437;
wire v_34438;
wire v_34439;
wire v_34440;
wire v_34441;
wire v_34442;
wire v_34443;
wire v_34444;
wire v_34445;
wire v_34446;
wire v_34447;
wire v_34448;
wire v_34449;
wire v_34450;
wire v_34451;
wire v_34452;
wire v_34453;
wire v_34454;
wire v_34455;
wire v_34456;
wire v_34457;
wire v_34458;
wire v_34459;
wire v_34460;
wire v_34461;
wire v_34462;
wire v_34463;
wire v_34464;
wire v_34465;
wire v_34466;
wire v_34467;
wire v_34468;
wire v_34469;
wire v_34470;
wire v_34471;
wire v_34472;
wire v_34473;
wire v_34474;
wire v_34475;
wire v_34476;
wire v_34477;
wire v_34478;
wire v_34479;
wire v_34480;
wire v_34481;
wire v_34482;
wire v_34483;
wire v_34484;
wire v_34485;
wire v_34486;
wire v_34487;
wire v_34488;
wire v_34489;
wire v_34490;
wire v_34491;
wire v_34492;
wire v_34493;
wire v_34494;
wire v_34495;
wire v_34496;
wire v_34497;
wire v_34498;
wire v_34499;
wire v_34500;
wire v_34501;
wire v_34502;
wire v_34503;
wire v_34504;
wire v_34505;
wire v_34506;
wire v_34507;
wire v_34508;
wire v_34509;
wire v_34510;
wire v_34511;
wire v_34512;
wire v_34513;
wire v_34514;
wire v_34515;
wire v_34516;
wire v_34517;
wire v_34518;
wire v_34519;
wire v_34520;
wire v_34521;
wire v_34522;
wire v_34523;
wire v_34524;
wire v_34525;
wire v_34526;
wire v_34527;
wire v_34528;
wire v_34529;
wire v_34530;
wire v_34531;
wire v_34532;
wire v_34533;
wire v_34534;
wire v_34535;
wire v_34536;
wire v_34537;
wire v_34538;
wire v_34539;
wire v_34540;
wire v_34541;
wire v_34542;
wire v_34543;
wire v_34544;
wire v_34545;
wire v_34546;
wire v_34547;
wire v_34548;
wire v_34549;
wire v_34550;
wire v_34551;
wire v_34552;
wire v_34553;
wire v_34554;
wire v_34555;
wire v_34556;
wire v_34557;
wire v_34558;
wire v_34559;
wire v_34560;
wire v_34561;
wire v_34562;
wire v_34563;
wire v_34564;
wire v_34565;
wire v_34566;
wire v_34567;
wire v_34568;
wire v_34569;
wire v_34570;
wire v_34571;
wire v_34572;
wire v_34573;
wire v_34574;
wire v_34575;
wire v_34576;
wire v_34577;
wire v_34578;
wire v_34579;
wire v_34580;
wire v_34581;
wire v_34582;
wire v_34583;
wire v_34584;
wire v_34585;
wire v_34586;
wire v_34587;
wire v_34588;
wire v_34589;
wire v_34590;
wire v_34591;
wire v_34592;
wire v_34593;
wire v_34594;
wire v_34595;
wire v_34596;
wire v_34597;
wire v_34598;
wire v_34599;
wire v_34600;
wire v_34601;
wire v_34602;
wire v_34603;
wire v_34604;
wire v_34605;
wire v_34606;
wire v_34607;
wire v_34608;
wire v_34609;
wire v_34610;
wire v_34611;
wire v_34612;
wire v_34613;
wire v_34614;
wire v_34615;
wire v_34616;
wire v_34617;
wire v_34618;
wire v_34619;
wire v_34620;
wire v_34621;
wire v_34622;
wire v_34623;
wire v_34624;
wire v_34625;
wire v_34626;
wire v_34627;
wire v_34628;
wire v_34629;
wire v_34630;
wire v_34631;
wire v_34632;
wire v_34633;
wire v_34634;
wire v_34635;
wire v_34636;
wire v_34637;
wire v_34638;
wire v_34639;
wire v_34640;
wire v_34641;
wire v_34642;
wire v_34643;
wire v_34644;
wire v_34645;
wire v_34646;
wire v_34647;
wire v_34648;
wire v_34649;
wire v_34650;
wire v_34651;
wire v_34652;
wire v_34653;
wire v_34654;
wire v_34655;
wire v_34656;
wire v_34657;
wire v_34658;
wire v_34659;
wire v_34660;
wire v_34661;
wire v_34662;
wire v_34663;
wire v_34664;
wire v_34665;
wire v_34666;
wire v_34667;
wire v_34668;
wire v_34669;
wire v_34670;
wire v_34671;
wire v_34672;
wire v_34673;
wire v_34674;
wire v_34675;
wire v_34676;
wire v_34677;
wire v_34678;
wire v_34679;
wire v_34680;
wire v_34681;
wire v_34682;
wire v_34683;
wire v_34684;
wire v_34685;
wire v_34686;
wire v_34687;
wire v_34688;
wire v_34689;
wire v_34690;
wire v_34691;
wire v_34692;
wire v_34693;
wire v_34694;
wire v_34695;
wire v_34696;
wire v_34697;
wire v_34698;
wire v_34699;
wire v_34700;
wire v_34701;
wire v_34702;
wire v_34703;
wire v_34704;
wire v_34705;
wire v_34706;
wire v_34707;
wire v_34708;
wire v_34709;
wire v_34710;
wire v_34711;
wire v_34712;
wire v_34713;
wire v_34714;
wire v_34715;
wire v_34716;
wire v_34717;
wire v_34718;
wire v_34719;
wire v_34720;
wire v_34721;
wire v_34722;
wire v_34723;
wire v_34724;
wire v_34725;
wire v_34726;
wire v_34727;
wire v_34728;
wire v_34729;
wire v_34730;
wire v_34731;
wire v_34732;
wire v_34733;
wire v_34734;
wire v_34735;
wire v_34736;
wire v_34737;
wire v_34738;
wire v_34739;
wire v_34740;
wire v_34741;
wire v_34742;
wire v_34743;
wire v_34744;
wire v_34745;
wire v_34746;
wire v_34747;
wire v_34748;
wire v_34749;
wire v_34750;
wire v_34751;
wire v_34752;
wire v_34753;
wire v_34754;
wire v_34755;
wire v_34756;
wire v_34757;
wire v_34758;
wire v_34759;
wire v_34760;
wire v_34761;
wire v_34762;
wire v_34763;
wire v_34764;
wire v_34765;
wire v_34766;
wire v_34767;
wire v_34768;
wire v_34769;
wire v_34770;
wire v_34771;
wire v_34772;
wire v_34773;
wire v_34774;
wire v_34775;
wire v_34776;
wire v_34777;
wire v_34778;
wire v_34779;
wire v_34780;
wire v_34781;
wire v_34782;
wire v_34783;
wire v_34784;
wire v_34785;
wire v_34786;
wire v_34787;
wire v_34788;
wire v_34789;
wire v_34790;
wire v_34791;
wire v_34792;
wire v_34793;
wire v_34794;
wire v_34795;
wire v_34796;
wire v_34797;
wire v_34798;
wire v_34799;
wire v_34800;
wire v_34801;
wire v_34802;
wire v_34803;
wire v_34804;
wire v_34805;
wire v_34806;
wire v_34807;
wire v_34808;
wire v_34809;
wire v_34810;
wire v_34811;
wire v_34812;
wire v_34813;
wire v_34814;
wire v_34815;
wire v_34816;
wire v_34817;
wire v_34818;
wire v_34819;
wire v_34820;
wire v_34821;
wire v_34822;
wire v_34823;
wire v_34824;
wire v_34825;
wire v_34826;
wire v_34827;
wire v_34828;
wire v_34829;
wire v_34830;
wire v_34831;
wire v_34832;
wire v_34833;
wire v_34834;
wire v_34835;
wire v_34836;
wire v_34837;
wire v_34838;
wire v_34839;
wire v_34840;
wire v_34841;
wire v_34842;
wire v_34843;
wire v_34844;
wire v_34845;
wire v_34846;
wire v_34847;
wire v_34848;
wire v_34849;
wire v_34850;
wire v_34851;
wire v_34853;
wire v_34854;
wire v_34855;
wire v_34856;
wire v_34857;
wire v_34858;
wire v_34859;
wire v_34860;
wire v_34861;
wire v_34862;
wire v_34863;
wire v_34864;
wire v_34865;
wire v_34866;
wire v_34867;
wire v_34868;
wire v_34869;
wire v_34870;
wire v_34871;
wire v_34872;
wire v_34873;
wire v_34874;
wire v_34875;
wire v_34876;
wire v_34877;
wire v_34878;
wire v_34879;
wire v_34880;
wire v_34881;
wire v_34882;
wire v_34883;
wire v_34884;
wire v_34885;
wire v_34886;
wire v_34887;
wire v_34888;
wire v_34889;
wire v_34890;
wire v_34891;
wire v_34892;
wire v_34893;
wire v_34894;
wire v_34895;
wire v_34896;
wire v_34897;
wire v_34898;
wire v_34899;
wire v_34900;
wire v_34901;
wire v_34902;
wire v_34903;
wire v_34904;
wire v_34905;
wire v_34906;
wire v_34907;
wire v_34908;
wire v_34909;
wire v_34910;
wire v_34911;
wire v_34912;
wire v_34913;
wire v_34914;
wire v_34915;
wire v_34916;
wire v_34917;
wire v_34918;
wire v_34919;
wire v_34920;
wire v_34921;
wire v_34922;
wire v_34923;
wire v_34924;
wire v_34925;
wire v_34926;
wire v_34927;
wire v_34928;
wire v_34929;
wire v_34930;
wire v_34931;
wire v_34932;
wire v_34933;
wire v_34934;
wire v_34935;
wire v_34936;
wire v_34937;
wire v_34938;
wire v_34939;
wire v_34940;
wire v_34941;
wire v_34942;
wire v_34943;
wire v_34944;
wire v_34945;
wire v_34946;
wire v_34947;
wire v_34948;
wire v_34949;
wire v_34950;
wire v_34951;
wire v_34952;
wire v_34953;
wire v_34954;
wire v_34955;
wire v_34956;
wire v_34957;
wire v_34958;
wire v_34959;
wire v_34960;
wire v_34961;
wire v_34962;
wire v_34963;
wire v_34964;
wire v_34965;
wire v_34966;
wire v_34967;
wire v_34968;
wire v_34969;
wire v_34970;
wire v_34971;
wire v_34972;
wire v_34973;
wire v_34974;
wire v_34975;
wire v_34976;
wire v_34977;
wire v_34978;
wire v_34979;
wire v_34980;
wire v_34981;
wire v_34982;
wire v_34983;
wire v_34984;
wire v_34985;
wire v_34986;
wire v_34987;
wire v_34988;
wire v_34989;
wire v_34990;
wire v_34991;
wire v_34992;
wire v_34993;
wire v_34994;
wire v_34995;
wire v_34996;
wire v_34997;
wire v_34998;
wire v_34999;
wire v_35000;
wire v_35001;
wire v_35002;
wire v_35003;
wire v_35004;
wire v_35005;
wire v_35006;
wire v_35007;
wire v_35008;
wire v_35009;
wire v_35010;
wire v_35011;
wire v_35012;
wire v_35013;
wire v_35014;
wire v_35015;
wire v_35016;
wire v_35017;
wire v_35018;
wire v_35019;
wire v_35020;
wire v_35021;
wire v_35022;
wire v_35023;
wire v_35024;
wire v_35025;
wire v_35026;
wire v_35027;
wire v_35028;
wire v_35029;
wire v_35030;
wire v_35031;
wire v_35032;
wire v_35033;
wire v_35034;
wire v_35035;
wire v_35036;
wire v_35037;
wire v_35038;
wire v_35039;
wire v_35040;
wire v_35041;
wire v_35042;
wire v_35043;
wire v_35044;
wire v_35045;
wire v_35046;
wire v_35047;
wire v_35048;
wire v_35049;
wire v_35050;
wire v_35051;
wire v_35052;
wire v_35053;
wire v_35054;
wire v_35055;
wire v_35056;
wire v_35057;
wire v_35058;
wire v_35059;
wire v_35060;
wire v_35061;
wire v_35062;
wire v_35063;
wire v_35064;
wire v_35065;
wire v_35066;
wire v_35067;
wire v_35068;
wire v_35069;
wire v_35070;
wire v_35071;
wire v_35072;
wire v_35073;
wire v_35074;
wire v_35075;
wire v_35076;
wire v_35077;
wire v_35078;
wire v_35079;
wire v_35080;
wire v_35081;
wire v_35082;
wire v_35083;
wire v_35084;
wire v_35085;
wire v_35086;
wire v_35087;
wire v_35088;
wire v_35089;
wire v_35090;
wire v_35091;
wire v_35092;
wire v_35093;
wire v_35094;
wire v_35095;
wire v_35096;
wire v_35097;
wire v_35098;
wire v_35099;
wire v_35100;
wire v_35101;
wire v_35102;
wire v_35103;
wire v_35104;
wire v_35105;
wire v_35106;
wire v_35107;
wire v_35108;
wire v_35109;
wire v_35110;
wire v_35111;
wire v_35112;
wire v_35113;
wire v_35114;
wire v_35115;
wire v_35116;
wire v_35117;
wire v_35118;
wire v_35119;
wire v_35120;
wire v_35121;
wire v_35122;
wire v_35123;
wire v_35124;
wire v_35125;
wire v_35126;
wire v_35127;
wire v_35128;
wire v_35129;
wire v_35130;
wire v_35131;
wire v_35132;
wire v_35133;
wire v_35134;
wire x_1;
assign v_34863 = 1;
assign v_2 = v_1;
assign v_5 = ~v_3 & v_4;
assign v_12 = v_10 & v_11;
assign v_17 = v_15 & v_16;
assign v_22 = v_20 & v_21;
assign v_27 = v_25 & v_26;
assign v_30 = v_28 & v_29;
assign v_31 = v_27 & v_30;
assign v_32 = ~v_23 & v_24;
assign v_34 = v_22 & v_33;
assign v_35 = ~v_18 & v_19;
assign v_37 = v_17 & v_36;
assign v_38 = v_13 & v_14;
assign v_40 = v_12 & v_39;
assign v_41 = v_8 & v_9;
assign v_44 = v_42 & v_43;
assign v_46 = v_44 & v_45;
assign v_52 = ~v_8 & ~v_9;
assign v_54 = ~v_13 & ~v_14;
assign v_56 = v_18 & ~v_19;
assign v_58 = v_23 & ~v_24;
assign v_62 = v_26 & v_61;
assign v_64 = v_21 & v_63;
assign v_66 = v_16 & v_65;
assign v_68 = v_11 & v_67;
assign v_70 = v_51 & v_69;
assign v_73 = v_67 & v_72;
assign v_76 = v_65 & v_75;
assign v_79 = v_63 & v_78;
assign v_82 = v_61 & v_81;
assign v_85 = v_60 & v_84;
assign v_95 = v_92 & v_94;
assign v_99 = v_97 & v_98;
assign v_100 = v_18 & v_23;
assign v_101 = ~v_13 & v_100;
assign v_102 = ~v_8 & v_101;
assign v_103 = ~v_43 & v_102;
assign v_104 = ~v_45 & v_103;
assign v_105 = ~v_47 & v_104;
assign v_106 = v_47 & v_104;
assign v_112 = ~v_47 & v_111;
assign v_114 = v_45 & v_103;
assign v_115 = ~v_45 & v_110;
assign v_117 = v_8 & v_101;
assign v_118 = ~v_8 & v_108;
assign v_120 = ~v_9 & v_119;
assign v_123 = v_121 & v_122;
assign v_124 = v_9 & v_123;
assign v_126 = v_13 & v_100;
assign v_127 = ~v_13 & v_107;
assign v_129 = ~v_14 & v_128;
assign v_132 = v_130 & v_131;
assign v_133 = v_14 & v_132;
assign v_135 = ~v_18 & v_23;
assign v_136 = v_18 & ~v_23;
assign v_138 = ~v_19 & v_137;
assign v_141 = v_139 & v_140;
assign v_142 = v_19 & v_141;
assign v_144 = ~v_23 & ~v_24;
assign v_145 = v_23 & v_24;
assign v_149 = v_147 & v_148;
assign v_152 = v_150 & v_151;
assign v_155 = v_153 & v_154;
assign v_158 = v_156 & v_157;
assign v_159 = v_43 & v_102;
assign v_160 = ~v_43 & v_109;
assign v_165 = v_105 & v_164;
assign v_168 = v_166 & v_167;
assign v_171 = v_169 & v_170;
assign v_173 = v_157 & v_172;
assign v_175 = v_154 & v_174;
assign v_177 = v_151 & v_176;
assign v_179 = v_148 & v_178;
assign v_180 = v_30 & v_179;
assign v_182 = v_177 & v_181;
assign v_184 = v_175 & v_183;
assign v_186 = v_173 & v_185;
assign v_190 = v_188 & v_189;
assign v_191 = v_187 & v_190;
assign v_192 = v_171 & v_191;
assign v_193 = v_168 & v_192;
assign v_197 = v_194 & v_196;
assign v_200 = v_164 & v_199;
assign v_203 = v_163 & v_202;
assign v_206 = v_162 & v_205;
assign v_209 = v_156 & v_208;
assign v_212 = v_153 & v_211;
assign v_215 = v_150 & v_214;
assign v_218 = v_147 & v_217;
assign v_224 = v_23 & ~v_28;
assign v_225 = v_18 & v_224;
assign v_226 = ~v_13 & v_225;
assign v_227 = ~v_8 & v_226;
assign v_228 = ~v_43 & v_227;
assign v_229 = ~v_45 & v_228;
assign v_230 = ~v_47 & v_229;
assign v_231 = v_47 & v_229;
assign v_238 = ~v_47 & v_237;
assign v_240 = v_45 & v_228;
assign v_241 = ~v_45 & v_236;
assign v_243 = v_8 & v_226;
assign v_244 = ~v_8 & v_234;
assign v_246 = ~v_9 & v_245;
assign v_249 = v_247 & v_248;
assign v_250 = v_9 & v_249;
assign v_252 = v_13 & v_225;
assign v_253 = ~v_13 & v_233;
assign v_255 = ~v_14 & v_254;
assign v_258 = v_256 & v_257;
assign v_259 = v_14 & v_258;
assign v_261 = ~v_18 & v_224;
assign v_262 = v_18 & v_232;
assign v_264 = ~v_19 & v_263;
assign v_267 = v_265 & v_266;
assign v_268 = v_19 & v_267;
assign v_270 = ~v_23 & ~v_28;
assign v_271 = v_23 & v_28;
assign v_273 = ~v_24 & v_272;
assign v_276 = v_274 & v_275;
assign v_277 = v_24 & v_276;
assign v_282 = v_280 & v_281;
assign v_285 = v_283 & v_284;
assign v_288 = v_286 & v_287;
assign v_291 = v_289 & v_290;
assign v_292 = v_43 & v_227;
assign v_293 = ~v_43 & v_235;
assign v_298 = v_230 & v_297;
assign v_301 = v_299 & v_300;
assign v_304 = v_302 & v_303;
assign v_306 = v_290 & v_305;
assign v_308 = v_287 & v_307;
assign v_310 = v_284 & v_309;
assign v_312 = v_281 & v_311;
assign v_313 = ~v_28 & v_29;
assign v_314 = v_312 & v_313;
assign v_316 = v_310 & v_315;
assign v_318 = v_308 & v_317;
assign v_320 = v_306 & v_319;
assign v_324 = v_322 & v_323;
assign v_325 = v_321 & v_324;
assign v_326 = v_304 & v_325;
assign v_327 = v_301 & v_326;
assign v_331 = v_328 & v_330;
assign v_334 = v_297 & v_333;
assign v_337 = v_296 & v_336;
assign v_340 = v_295 & v_339;
assign v_343 = v_289 & v_342;
assign v_346 = v_286 & v_345;
assign v_349 = v_283 & v_348;
assign v_352 = v_280 & v_351;
assign v_355 = v_279 & v_354;
assign v_360 = v_223 & v_359;
assign v_363 = v_99 & v_362;
assign v_364 = ~v_18 & ~v_23;
assign v_365 = v_13 & v_364;
assign v_366 = v_8 & v_365;
assign v_367 = v_43 & v_366;
assign v_368 = v_45 & v_367;
assign v_376 = v_369 & v_375;
assign v_378 = v_374 & v_377;
assign v_380 = v_372 & v_379;
assign v_382 = ~v_8 & v_371;
assign v_385 = v_381 & v_384;
assign v_387 = v_371 & v_386;
assign v_389 = ~v_13 & v_370;
assign v_392 = v_388 & v_391;
assign v_393 = v_107 & v_370;
assign v_397 = v_394 & v_396;
assign v_398 = v_181 & v_397;
assign v_399 = v_19 & v_393;
assign v_401 = v_392 & v_400;
assign v_402 = v_14 & v_387;
assign v_404 = v_385 & v_403;
assign v_405 = v_9 & v_380;
assign v_408 = v_373 & v_407;
assign v_409 = v_406 & v_408;
assign v_410 = v_378 & v_409;
assign v_411 = v_376 & v_410;
assign v_412 = v_47 & v_368;
assign v_417 = ~v_45 & v_373;
assign v_419 = ~v_9 & v_383;
assign v_421 = ~v_14 & v_390;
assign v_423 = ~v_19 & v_395;
assign v_426 = v_396 & v_425;
assign v_428 = v_391 & v_427;
assign v_430 = v_384 & v_429;
assign v_431 = ~v_43 & v_372;
assign v_435 = v_416 & v_434;
assign v_438 = v_433 & v_437;
assign v_441 = v_429 & v_440;
assign v_444 = v_427 & v_443;
assign v_447 = v_425 & v_446;
assign v_454 = ~v_23 & v_28;
assign v_455 = ~v_18 & v_454;
assign v_456 = v_13 & v_455;
assign v_457 = v_8 & v_456;
assign v_458 = v_43 & v_457;
assign v_459 = v_45 & v_458;
assign v_468 = v_460 & v_467;
assign v_470 = v_466 & v_469;
assign v_472 = v_464 & v_471;
assign v_474 = ~v_8 & v_463;
assign v_477 = v_473 & v_476;
assign v_479 = v_463 & v_478;
assign v_481 = ~v_13 & v_462;
assign v_484 = v_480 & v_483;
assign v_486 = v_462 & v_485;
assign v_488 = v_18 & v_461;
assign v_491 = v_487 & v_490;
assign v_492 = v_232 & v_461;
assign v_496 = v_493 & v_495;
assign v_497 = v_313 & v_496;
assign v_498 = v_24 & v_492;
assign v_500 = v_491 & v_499;
assign v_501 = v_19 & v_486;
assign v_503 = v_484 & v_502;
assign v_504 = v_14 & v_479;
assign v_506 = v_477 & v_505;
assign v_507 = v_9 & v_472;
assign v_510 = v_465 & v_509;
assign v_511 = v_508 & v_510;
assign v_512 = v_470 & v_511;
assign v_513 = v_468 & v_512;
assign v_514 = v_47 & v_459;
assign v_519 = ~v_45 & v_465;
assign v_521 = ~v_9 & v_475;
assign v_523 = ~v_14 & v_482;
assign v_525 = ~v_19 & v_489;
assign v_527 = ~v_24 & v_494;
assign v_530 = v_495 & v_529;
assign v_532 = v_490 & v_531;
assign v_534 = v_483 & v_533;
assign v_536 = v_476 & v_535;
assign v_537 = ~v_43 & v_464;
assign v_541 = v_518 & v_540;
assign v_544 = v_539 & v_543;
assign v_547 = v_535 & v_546;
assign v_550 = v_533 & v_549;
assign v_553 = v_531 & v_552;
assign v_556 = v_529 & v_555;
assign v_562 = v_453 & v_561;
assign v_565 = v_363 & v_564;
assign v_568 = ~v_47 & v_567;
assign v_569 = ~v_45 & v_69;
assign v_570 = v_568 & v_569;
assign v_571 = ~v_43 & v_68;
assign v_573 = v_570 & v_572;
assign v_574 = v_53 & v_66;
assign v_576 = v_573 & v_575;
assign v_577 = v_55 & v_64;
assign v_579 = v_576 & v_578;
assign v_580 = v_57 & v_62;
assign v_582 = v_579 & v_581;
assign v_583 = v_59 & v_60;
assign v_585 = v_582 & v_584;
assign v_586 = ~v_28 & ~v_29;
assign v_588 = v_585 & v_587;
assign v_589 = v_87 & v_588;
assign v_590 = v_89 & v_589;
assign v_591 = ~v_91 & v_590;
assign v_592 = ~v_89 & v_589;
assign v_593 = v_91 & v_592;
assign v_595 = v_96 & v_594;
assign v_598 = v_164 & v_195;
assign v_599 = v_105 & v_193;
assign v_601 = v_597 & v_600;
assign v_602 = v_113 & v_163;
assign v_604 = v_601 & v_603;
assign v_605 = v_116 & v_162;
assign v_607 = v_604 & v_606;
assign v_608 = v_158 & v_161;
assign v_610 = v_607 & v_609;
assign v_611 = v_125 & v_155;
assign v_613 = v_610 & v_612;
assign v_614 = v_134 & v_152;
assign v_616 = v_613 & v_615;
assign v_617 = v_143 & v_149;
assign v_619 = v_616 & v_618;
assign v_620 = v_60 & v_146;
assign v_622 = v_619 & v_621;
assign v_623 = v_587 & v_622;
assign v_624 = v_87 & v_623;
assign v_625 = ~v_89 & v_624;
assign v_626 = ~v_91 & v_625;
assign v_628 = v_297 & v_329;
assign v_629 = v_230 & v_327;
assign v_631 = v_627 & v_630;
assign v_632 = v_239 & v_296;
assign v_634 = v_631 & v_633;
assign v_635 = v_242 & v_295;
assign v_637 = v_634 & v_636;
assign v_638 = v_291 & v_294;
assign v_640 = v_637 & v_639;
assign v_641 = v_251 & v_288;
assign v_643 = v_640 & v_642;
assign v_644 = v_260 & v_285;
assign v_646 = v_643 & v_645;
assign v_647 = v_269 & v_282;
assign v_649 = v_646 & v_648;
assign v_650 = v_278 & v_279;
assign v_652 = v_649 & v_651;
assign v_653 = v_28 & ~v_29;
assign v_655 = v_652 & v_654;
assign v_656 = v_87 & v_655;
assign v_657 = ~v_89 & v_656;
assign v_658 = ~v_91 & v_657;
assign v_660 = v_361 & v_659;
assign v_662 = ~v_47 & v_374;
assign v_665 = v_375 & v_664;
assign v_666 = v_434 & v_663;
assign v_667 = v_665 & v_666;
assign v_668 = v_418 & v_433;
assign v_670 = v_667 & v_669;
assign v_671 = v_430 & v_432;
assign v_673 = v_670 & v_672;
assign v_674 = v_420 & v_428;
assign v_676 = v_673 & v_675;
assign v_677 = v_422 & v_426;
assign v_679 = v_676 & v_678;
assign v_680 = v_149 & v_424;
assign v_682 = v_679 & v_681;
assign v_683 = v_621 & v_682;
assign v_684 = v_587 & v_683;
assign v_685 = v_87 & v_684;
assign v_686 = ~v_89 & v_685;
assign v_687 = ~v_91 & v_686;
assign v_688 = ~v_47 & v_466;
assign v_691 = v_467 & v_690;
assign v_692 = v_540 & v_689;
assign v_693 = v_691 & v_692;
assign v_694 = v_520 & v_539;
assign v_696 = v_693 & v_695;
assign v_697 = v_536 & v_538;
assign v_699 = v_696 & v_698;
assign v_700 = v_522 & v_534;
assign v_702 = v_699 & v_701;
assign v_703 = v_524 & v_532;
assign v_705 = v_702 & v_704;
assign v_706 = v_526 & v_530;
assign v_708 = v_705 & v_707;
assign v_709 = v_279 & v_528;
assign v_711 = v_708 & v_710;
assign v_712 = v_654 & v_711;
assign v_713 = v_87 & v_712;
assign v_714 = ~v_89 & v_713;
assign v_715 = ~v_91 & v_714;
assign v_717 = v_563 & v_716;
assign v_722 = v_97 & v_721;
assign v_723 = v_362 & v_722;
assign v_724 = v_564 & v_723;
assign v_732 = v_97 & v_731;
assign v_733 = v_362 & v_732;
assign v_734 = v_564 & v_733;
assign v_742 = v_97 & v_741;
assign v_743 = v_362 & v_742;
assign v_744 = v_564 & v_743;
assign v_752 = v_97 & v_751;
assign v_753 = v_362 & v_752;
assign v_754 = v_564 & v_753;
assign v_762 = v_97 & v_761;
assign v_763 = v_362 & v_762;
assign v_764 = v_564 & v_763;
assign v_772 = v_97 & v_771;
assign v_773 = v_94 & v_595;
assign v_775 = v_362 & v_774;
assign v_776 = v_359 & v_660;
assign v_778 = v_564 & v_777;
assign v_779 = v_561 & v_717;
assign v_784 = v_782 & v_783;
assign v_787 = v_785 & v_786;
assign v_790 = v_788 & v_789;
assign v_798 = v_97 & ~v_793;
assign v_799 = v_362 & v_798;
assign v_800 = v_564 & v_799;
assign v_805 = v_803 & v_804;
assign v_809 = v_805 & v_808;
assign v_812 = v_810 & v_811;
assign v_814 = v_809 & v_813;
assign v_817 = v_815 & v_816;
assign v_819 = v_814 & v_818;
assign v_821 = v_96 & v_590;
assign v_823 = ~v_91 & v_592;
assign v_824 = v_807 & v_823;
assign v_826 = v_91 & v_625;
assign v_827 = v_91 & v_657;
assign v_829 = v_361 & v_828;
assign v_831 = v_91 & v_686;
assign v_832 = v_91 & v_714;
assign v_834 = v_563 & v_833;
assign v_839 = v_803 & v_838;
assign v_840 = v_808 & v_839;
assign v_841 = v_813 & v_840;
assign v_842 = v_818 & v_841;
assign v_851 = v_803 & v_850;
assign v_852 = v_808 & v_851;
assign v_853 = v_813 & v_852;
assign v_854 = v_818 & v_853;
assign v_863 = v_803 & v_862;
assign v_864 = v_808 & v_863;
assign v_865 = v_813 & v_864;
assign v_866 = v_818 & v_865;
assign v_875 = v_803 & v_874;
assign v_876 = v_808 & v_875;
assign v_877 = v_813 & v_876;
assign v_878 = v_818 & v_877;
assign v_887 = v_803 & v_886;
assign v_888 = v_808 & v_887;
assign v_889 = v_813 & v_888;
assign v_890 = v_818 & v_889;
assign v_899 = v_803 & v_898;
assign v_900 = v_91 & v_821;
assign v_902 = v_808 & v_901;
assign v_903 = v_813 & v_902;
assign v_904 = v_811 & v_829;
assign v_906 = v_818 & v_905;
assign v_907 = v_816 & v_834;
assign v_912 = v_910 & v_911;
assign v_916 = v_914 & v_915;
assign v_919 = v_917 & v_918;
assign v_928 = v_803 & ~v_922;
assign v_929 = v_808 & v_928;
assign v_930 = v_813 & v_929;
assign v_931 = v_818 & v_930;
assign v_938 = v_936 & v_937;
assign v_941 = v_939 & v_940;
assign v_943 = v_941 & v_942;
assign v_948 = v_945 & v_947;
assign v_950 = v_943 & v_949;
assign v_955 = v_952 & v_954;
assign v_957 = v_950 & v_956;
assign v_959 = ~v_87 & v_588;
assign v_960 = ~v_89 & v_959;
assign v_961 = ~v_91 & v_960;
assign v_962 = v_91 & v_590;
assign v_964 = v_96 & v_963;
assign v_966 = v_592 & v_807;
assign v_968 = v_89 & v_624;
assign v_969 = ~v_91 & v_968;
assign v_970 = v_89 & v_656;
assign v_971 = ~v_91 & v_970;
assign v_973 = v_361 & v_972;
assign v_975 = v_89 & v_685;
assign v_976 = ~v_91 & v_975;
assign v_977 = v_89 & v_713;
assign v_978 = ~v_91 & v_977;
assign v_980 = v_563 & v_979;
assign v_985 = v_939 & v_984;
assign v_986 = v_942 & v_985;
assign v_987 = v_949 & v_986;
assign v_988 = v_956 & v_987;
assign v_997 = v_939 & v_996;
assign v_998 = v_942 & v_997;
assign v_999 = v_949 & v_998;
assign v_1000 = v_956 & v_999;
assign v_1009 = v_939 & v_1008;
assign v_1010 = v_942 & v_1009;
assign v_1011 = v_949 & v_1010;
assign v_1012 = v_956 & v_1011;
assign v_1021 = v_939 & v_1020;
assign v_1022 = v_942 & v_1021;
assign v_1023 = v_949 & v_1022;
assign v_1024 = v_956 & v_1023;
assign v_1033 = v_939 & v_1032;
assign v_1034 = v_942 & v_1033;
assign v_1035 = v_949 & v_1034;
assign v_1036 = v_956 & v_1035;
assign v_1045 = v_939 & v_1044;
assign v_1046 = v_937 & v_964;
assign v_1048 = v_942 & v_1047;
assign v_1049 = ~v_91 & v_966;
assign v_1051 = v_949 & v_1050;
assign v_1052 = v_947 & v_973;
assign v_1054 = v_956 & v_1053;
assign v_1055 = v_954 & v_980;
assign v_1060 = v_1058 & v_1059;
assign v_1063 = v_1061 & v_1062;
assign v_1066 = v_1064 & v_1065;
assign v_1069 = v_1067 & v_1068;
assign v_1078 = v_939 & ~v_1072;
assign v_1079 = v_942 & v_1078;
assign v_1080 = v_949 & v_1079;
assign v_1081 = v_956 & v_1080;
assign v_1086 = v_1084 & v_1085;
assign v_1088 = v_1086 & v_1087;
assign v_1091 = v_1089 & v_1090;
assign v_1093 = v_1088 & v_1092;
assign v_1096 = v_1094 & v_1095;
assign v_1098 = v_1093 & v_1097;
assign v_1100 = v_96 & v_960;
assign v_1102 = v_594 & v_807;
assign v_1104 = v_91 & v_968;
assign v_1105 = v_91 & v_970;
assign v_1107 = v_361 & v_1106;
assign v_1109 = v_91 & v_975;
assign v_1110 = v_91 & v_977;
assign v_1112 = v_563 & v_1111;
assign v_1117 = v_1084 & v_1116;
assign v_1118 = v_1087 & v_1117;
assign v_1119 = v_1092 & v_1118;
assign v_1120 = v_1097 & v_1119;
assign v_1129 = v_1084 & v_1128;
assign v_1130 = v_1087 & v_1129;
assign v_1131 = v_1092 & v_1130;
assign v_1132 = v_1097 & v_1131;
assign v_1141 = v_1084 & v_1140;
assign v_1142 = v_1087 & v_1141;
assign v_1143 = v_1092 & v_1142;
assign v_1144 = v_1097 & v_1143;
assign v_1153 = v_1084 & v_1152;
assign v_1154 = v_1087 & v_1153;
assign v_1155 = v_1092 & v_1154;
assign v_1156 = v_1097 & v_1155;
assign v_1165 = v_1084 & v_1164;
assign v_1166 = v_1087 & v_1165;
assign v_1167 = v_1092 & v_1166;
assign v_1168 = v_1097 & v_1167;
assign v_1177 = v_1084 & v_1176;
assign v_1178 = v_91 & v_1100;
assign v_1180 = v_1087 & v_1179;
assign v_1181 = v_92 & v_1102;
assign v_1183 = v_1092 & v_1182;
assign v_1184 = v_1090 & v_1107;
assign v_1186 = v_1097 & v_1185;
assign v_1187 = v_1095 & v_1112;
assign v_1192 = v_1190 & v_1191;
assign v_1195 = v_1193 & v_1194;
assign v_1198 = v_1196 & v_1197;
assign v_1201 = v_1199 & v_1200;
assign v_1210 = v_1084 & ~v_1204;
assign v_1211 = v_1087 & v_1210;
assign v_1212 = v_1092 & v_1211;
assign v_1213 = v_1097 & v_1212;
assign v_1219 = v_1217 & v_1218;
assign v_1222 = v_1220 & v_1221;
assign v_1224 = v_1222 & v_1223;
assign v_1231 = v_1227 & v_1230;
assign v_1233 = v_1224 & v_1232;
assign v_1240 = v_1236 & v_1239;
assign v_1242 = v_1233 & v_1241;
assign v_1244 = v_89 & v_959;
assign v_1245 = ~v_91 & v_1244;
assign v_1246 = v_91 & v_960;
assign v_1248 = v_96 & v_1247;
assign v_1250 = v_590 & v_807;
assign v_1252 = ~v_87 & v_623;
assign v_1253 = ~v_89 & v_1252;
assign v_1254 = ~v_91 & v_1253;
assign v_1255 = ~v_87 & v_655;
assign v_1256 = ~v_89 & v_1255;
assign v_1257 = ~v_91 & v_1256;
assign v_1259 = v_361 & v_1258;
assign v_1261 = ~v_87 & v_684;
assign v_1262 = ~v_89 & v_1261;
assign v_1263 = ~v_91 & v_1262;
assign v_1264 = ~v_87 & v_712;
assign v_1265 = ~v_89 & v_1264;
assign v_1266 = ~v_91 & v_1265;
assign v_1268 = v_563 & v_1267;
assign v_1273 = v_1220 & v_1272;
assign v_1274 = v_1223 & v_1273;
assign v_1275 = v_1232 & v_1274;
assign v_1276 = v_1241 & v_1275;
assign v_1285 = v_1220 & v_1284;
assign v_1286 = v_1223 & v_1285;
assign v_1287 = v_1232 & v_1286;
assign v_1288 = v_1241 & v_1287;
assign v_1297 = v_1220 & v_1296;
assign v_1298 = v_1223 & v_1297;
assign v_1299 = v_1232 & v_1298;
assign v_1300 = v_1241 & v_1299;
assign v_1309 = v_1220 & v_1308;
assign v_1310 = v_1223 & v_1309;
assign v_1311 = v_1232 & v_1310;
assign v_1312 = v_1241 & v_1311;
assign v_1321 = v_1220 & v_1320;
assign v_1322 = v_1223 & v_1321;
assign v_1323 = v_1232 & v_1322;
assign v_1324 = v_1241 & v_1323;
assign v_1333 = v_1220 & v_1332;
assign v_1334 = v_1218 & v_1248;
assign v_1336 = v_1223 & v_1335;
assign v_1337 = ~v_91 & v_1250;
assign v_1339 = v_1232 & v_1338;
assign v_1340 = v_1230 & v_1259;
assign v_1342 = v_1241 & v_1341;
assign v_1343 = v_1239 & v_1268;
assign v_1348 = v_1346 & v_1347;
assign v_1351 = v_1349 & v_1350;
assign v_1354 = v_1352 & v_1353;
assign v_1357 = v_1355 & v_1356;
assign v_1366 = v_1220 & ~v_1360;
assign v_1367 = v_1223 & v_1366;
assign v_1368 = v_1232 & v_1367;
assign v_1369 = v_1241 & v_1368;
assign v_1374 = v_1372 & v_1373;
assign v_1376 = v_1374 & v_1375;
assign v_1379 = v_1377 & v_1378;
assign v_1381 = v_1376 & v_1380;
assign v_1384 = v_1382 & v_1383;
assign v_1386 = v_1381 & v_1385;
assign v_1388 = v_96 & v_1244;
assign v_1390 = v_807 & v_963;
assign v_1392 = v_91 & v_1253;
assign v_1393 = v_91 & v_1256;
assign v_1395 = v_361 & v_1394;
assign v_1397 = v_91 & v_1262;
assign v_1398 = v_91 & v_1265;
assign v_1400 = v_563 & v_1399;
assign v_1405 = v_1372 & v_1404;
assign v_1406 = v_1375 & v_1405;
assign v_1407 = v_1380 & v_1406;
assign v_1408 = v_1385 & v_1407;
assign v_1417 = v_1372 & v_1416;
assign v_1418 = v_1375 & v_1417;
assign v_1419 = v_1380 & v_1418;
assign v_1420 = v_1385 & v_1419;
assign v_1429 = v_1372 & v_1428;
assign v_1430 = v_1375 & v_1429;
assign v_1431 = v_1380 & v_1430;
assign v_1432 = v_1385 & v_1431;
assign v_1441 = v_1372 & v_1440;
assign v_1442 = v_1375 & v_1441;
assign v_1443 = v_1380 & v_1442;
assign v_1444 = v_1385 & v_1443;
assign v_1453 = v_1372 & v_1452;
assign v_1454 = v_1375 & v_1453;
assign v_1455 = v_1380 & v_1454;
assign v_1456 = v_1385 & v_1455;
assign v_1465 = v_1372 & v_1464;
assign v_1466 = v_91 & v_1388;
assign v_1468 = v_1375 & v_1467;
assign v_1469 = v_936 & v_1390;
assign v_1471 = v_1380 & v_1470;
assign v_1472 = v_1378 & v_1395;
assign v_1474 = v_1385 & v_1473;
assign v_1475 = v_1383 & v_1400;
assign v_1480 = v_1478 & v_1479;
assign v_1483 = v_1481 & v_1482;
assign v_1486 = v_1484 & v_1485;
assign v_1489 = v_1487 & v_1488;
assign v_1498 = v_1372 & ~v_1492;
assign v_1499 = v_1375 & v_1498;
assign v_1500 = v_1380 & v_1499;
assign v_1501 = v_1385 & v_1500;
assign v_1509 = v_1507 & v_1508;
assign v_1512 = v_1510 & v_1511;
assign v_1514 = v_1512 & v_1513;
assign v_1519 = v_1516 & v_1518;
assign v_1521 = v_1514 & v_1520;
assign v_1526 = v_1523 & v_1525;
assign v_1528 = v_1521 & v_1527;
assign v_1530 = v_85 & v_585;
assign v_1531 = v_87 & v_1530;
assign v_1532 = ~v_89 & v_1531;
assign v_1533 = ~v_91 & v_1532;
assign v_1534 = v_91 & v_1244;
assign v_1536 = v_96 & v_1535;
assign v_1538 = v_807 & v_960;
assign v_1540 = v_89 & v_1252;
assign v_1541 = ~v_91 & v_1540;
assign v_1542 = v_89 & v_1255;
assign v_1543 = ~v_91 & v_1542;
assign v_1545 = v_361 & v_1544;
assign v_1547 = v_89 & v_1261;
assign v_1548 = ~v_91 & v_1547;
assign v_1549 = v_89 & v_1264;
assign v_1550 = ~v_91 & v_1549;
assign v_1552 = v_563 & v_1551;
assign v_1557 = v_1510 & v_1556;
assign v_1558 = v_1513 & v_1557;
assign v_1559 = v_1520 & v_1558;
assign v_1560 = v_1527 & v_1559;
assign v_1569 = v_1510 & v_1568;
assign v_1570 = v_1513 & v_1569;
assign v_1571 = v_1520 & v_1570;
assign v_1572 = v_1527 & v_1571;
assign v_1581 = v_1510 & v_1580;
assign v_1582 = v_1513 & v_1581;
assign v_1583 = v_1520 & v_1582;
assign v_1584 = v_1527 & v_1583;
assign v_1593 = v_1510 & v_1592;
assign v_1594 = v_1513 & v_1593;
assign v_1595 = v_1520 & v_1594;
assign v_1596 = v_1527 & v_1595;
assign v_1605 = v_1510 & v_1604;
assign v_1606 = v_1513 & v_1605;
assign v_1607 = v_1520 & v_1606;
assign v_1608 = v_1527 & v_1607;
assign v_1617 = v_1510 & v_1616;
assign v_1618 = v_1508 & v_1536;
assign v_1620 = v_1513 & v_1619;
assign v_1621 = ~v_91 & v_1538;
assign v_1623 = v_1520 & v_1622;
assign v_1624 = v_1518 & v_1545;
assign v_1626 = v_1527 & v_1625;
assign v_1627 = v_1525 & v_1552;
assign v_1632 = v_1630 & v_1631;
assign v_1635 = v_1633 & v_1634;
assign v_1638 = v_1636 & v_1637;
assign v_1641 = v_1639 & v_1640;
assign v_1650 = v_1510 & ~v_1644;
assign v_1651 = v_1513 & v_1650;
assign v_1652 = v_1520 & v_1651;
assign v_1653 = v_1527 & v_1652;
assign v_1658 = v_1656 & v_1657;
assign v_1660 = v_1658 & v_1659;
assign v_1663 = v_1661 & v_1662;
assign v_1665 = v_1660 & v_1664;
assign v_1668 = v_1666 & v_1667;
assign v_1670 = v_1665 & v_1669;
assign v_1672 = v_96 & v_1532;
assign v_1674 = v_807 & v_1247;
assign v_1676 = v_91 & v_1540;
assign v_1677 = v_91 & v_1542;
assign v_1679 = v_361 & v_1678;
assign v_1681 = v_91 & v_1547;
assign v_1682 = v_91 & v_1549;
assign v_1684 = v_563 & v_1683;
assign v_1689 = v_1656 & v_1688;
assign v_1690 = v_1659 & v_1689;
assign v_1691 = v_1664 & v_1690;
assign v_1692 = v_1669 & v_1691;
assign v_1701 = v_1656 & v_1700;
assign v_1702 = v_1659 & v_1701;
assign v_1703 = v_1664 & v_1702;
assign v_1704 = v_1669 & v_1703;
assign v_1713 = v_1656 & v_1712;
assign v_1714 = v_1659 & v_1713;
assign v_1715 = v_1664 & v_1714;
assign v_1716 = v_1669 & v_1715;
assign v_1725 = v_1656 & v_1724;
assign v_1726 = v_1659 & v_1725;
assign v_1727 = v_1664 & v_1726;
assign v_1728 = v_1669 & v_1727;
assign v_1737 = v_1656 & v_1736;
assign v_1738 = v_1659 & v_1737;
assign v_1739 = v_1664 & v_1738;
assign v_1740 = v_1669 & v_1739;
assign v_1749 = v_1656 & v_1748;
assign v_1750 = v_91 & v_1672;
assign v_1752 = v_1659 & v_1751;
assign v_1753 = v_1217 & v_1674;
assign v_1755 = v_1664 & v_1754;
assign v_1756 = v_1662 & v_1679;
assign v_1758 = v_1669 & v_1757;
assign v_1759 = v_1667 & v_1684;
assign v_1764 = v_1762 & v_1763;
assign v_1767 = v_1765 & v_1766;
assign v_1770 = v_1768 & v_1769;
assign v_1773 = v_1771 & v_1772;
assign v_1782 = v_1656 & ~v_1776;
assign v_1783 = v_1659 & v_1782;
assign v_1784 = v_1664 & v_1783;
assign v_1785 = v_1669 & v_1784;
assign v_1791 = v_1789 & v_1790;
assign v_1794 = v_1792 & v_1793;
assign v_1796 = v_1794 & v_1795;
assign v_1805 = v_1800 & v_1804;
assign v_1807 = v_1796 & v_1806;
assign v_1816 = v_1811 & v_1815;
assign v_1818 = v_1807 & v_1817;
assign v_1820 = v_89 & v_1531;
assign v_1821 = ~v_91 & v_1820;
assign v_1822 = v_91 & v_1532;
assign v_1824 = v_96 & v_1823;
assign v_1826 = v_807 & v_1244;
assign v_1828 = v_85 & v_622;
assign v_1829 = v_87 & v_1828;
assign v_1830 = ~v_89 & v_1829;
assign v_1831 = ~v_91 & v_1830;
assign v_1832 = v_355 & v_652;
assign v_1833 = v_87 & v_1832;
assign v_1834 = ~v_89 & v_1833;
assign v_1835 = ~v_91 & v_1834;
assign v_1837 = v_361 & v_1836;
assign v_1839 = v_85 & v_683;
assign v_1840 = v_87 & v_1839;
assign v_1841 = ~v_89 & v_1840;
assign v_1842 = ~v_91 & v_1841;
assign v_1843 = v_355 & v_711;
assign v_1844 = v_87 & v_1843;
assign v_1845 = ~v_89 & v_1844;
assign v_1846 = ~v_91 & v_1845;
assign v_1848 = v_563 & v_1847;
assign v_1853 = v_1792 & v_1852;
assign v_1854 = v_1795 & v_1853;
assign v_1855 = v_1806 & v_1854;
assign v_1856 = v_1817 & v_1855;
assign v_1865 = v_1792 & v_1864;
assign v_1866 = v_1795 & v_1865;
assign v_1867 = v_1806 & v_1866;
assign v_1868 = v_1817 & v_1867;
assign v_1877 = v_1792 & v_1876;
assign v_1878 = v_1795 & v_1877;
assign v_1879 = v_1806 & v_1878;
assign v_1880 = v_1817 & v_1879;
assign v_1889 = v_1792 & v_1888;
assign v_1890 = v_1795 & v_1889;
assign v_1891 = v_1806 & v_1890;
assign v_1892 = v_1817 & v_1891;
assign v_1901 = v_1792 & v_1900;
assign v_1902 = v_1795 & v_1901;
assign v_1903 = v_1806 & v_1902;
assign v_1904 = v_1817 & v_1903;
assign v_1913 = v_1792 & v_1912;
assign v_1914 = v_1790 & v_1824;
assign v_1916 = v_1795 & v_1915;
assign v_1917 = ~v_91 & v_1826;
assign v_1919 = v_1806 & v_1918;
assign v_1920 = v_1804 & v_1837;
assign v_1922 = v_1817 & v_1921;
assign v_1923 = v_1815 & v_1848;
assign v_1928 = v_1926 & v_1927;
assign v_1931 = v_1929 & v_1930;
assign v_1934 = v_1932 & v_1933;
assign v_1937 = v_1935 & v_1936;
assign v_1946 = v_1792 & ~v_1940;
assign v_1947 = v_1795 & v_1946;
assign v_1948 = v_1806 & v_1947;
assign v_1949 = v_1817 & v_1948;
assign v_1954 = v_1952 & v_1953;
assign v_1956 = v_1954 & v_1955;
assign v_1959 = v_1957 & v_1958;
assign v_1961 = v_1956 & v_1960;
assign v_1964 = v_1962 & v_1963;
assign v_1966 = v_1961 & v_1965;
assign v_1968 = v_96 & v_1820;
assign v_1970 = v_807 & v_1535;
assign v_1972 = v_91 & v_1830;
assign v_1973 = v_91 & v_1834;
assign v_1975 = v_361 & v_1974;
assign v_1977 = v_91 & v_1841;
assign v_1978 = v_91 & v_1845;
assign v_1980 = v_563 & v_1979;
assign v_1985 = v_1952 & v_1984;
assign v_1986 = v_1955 & v_1985;
assign v_1987 = v_1960 & v_1986;
assign v_1988 = v_1965 & v_1987;
assign v_1997 = v_1952 & v_1996;
assign v_1998 = v_1955 & v_1997;
assign v_1999 = v_1960 & v_1998;
assign v_2000 = v_1965 & v_1999;
assign v_2009 = v_1952 & v_2008;
assign v_2010 = v_1955 & v_2009;
assign v_2011 = v_1960 & v_2010;
assign v_2012 = v_1965 & v_2011;
assign v_2021 = v_1952 & v_2020;
assign v_2022 = v_1955 & v_2021;
assign v_2023 = v_1960 & v_2022;
assign v_2024 = v_1965 & v_2023;
assign v_2033 = v_1952 & v_2032;
assign v_2034 = v_1955 & v_2033;
assign v_2035 = v_1960 & v_2034;
assign v_2036 = v_1965 & v_2035;
assign v_2045 = v_1952 & v_2044;
assign v_2046 = v_91 & v_1968;
assign v_2048 = v_1955 & v_2047;
assign v_2049 = v_1507 & v_1970;
assign v_2051 = v_1960 & v_2050;
assign v_2052 = v_1958 & v_1975;
assign v_2054 = v_1965 & v_2053;
assign v_2055 = v_1963 & v_1980;
assign v_2060 = v_2058 & v_2059;
assign v_2063 = v_2061 & v_2062;
assign v_2066 = v_2064 & v_2065;
assign v_2069 = v_2067 & v_2068;
assign v_2073 = v_1952 & v_2072;
assign v_2074 = v_1955 & v_2073;
assign v_2075 = v_1960 & v_2074;
assign v_2076 = v_1965 & v_2075;
assign v_2088 = v_2086 & v_2087;
assign v_2091 = v_2089 & v_2090;
assign v_2093 = v_2091 & v_2092;
assign v_2098 = v_2095 & v_2097;
assign v_2100 = v_2093 & v_2099;
assign v_2105 = v_2102 & v_2104;
assign v_2107 = v_2100 & v_2106;
assign v_2109 = ~v_87 & v_1530;
assign v_2110 = ~v_89 & v_2109;
assign v_2111 = ~v_91 & v_2110;
assign v_2112 = v_91 & v_1820;
assign v_2114 = v_96 & v_2113;
assign v_2116 = v_807 & v_1532;
assign v_2118 = v_89 & v_1829;
assign v_2119 = ~v_91 & v_2118;
assign v_2120 = v_89 & v_1833;
assign v_2121 = ~v_91 & v_2120;
assign v_2123 = v_361 & v_2122;
assign v_2125 = v_89 & v_1840;
assign v_2126 = ~v_91 & v_2125;
assign v_2127 = v_89 & v_1844;
assign v_2128 = ~v_91 & v_2127;
assign v_2130 = v_563 & v_2129;
assign v_2135 = v_2089 & v_2134;
assign v_2136 = v_2092 & v_2135;
assign v_2137 = v_2099 & v_2136;
assign v_2138 = v_2106 & v_2137;
assign v_2147 = v_2089 & v_2146;
assign v_2148 = v_2092 & v_2147;
assign v_2149 = v_2099 & v_2148;
assign v_2150 = v_2106 & v_2149;
assign v_2159 = v_2089 & v_2158;
assign v_2160 = v_2092 & v_2159;
assign v_2161 = v_2099 & v_2160;
assign v_2162 = v_2106 & v_2161;
assign v_2171 = v_2089 & v_2170;
assign v_2172 = v_2092 & v_2171;
assign v_2173 = v_2099 & v_2172;
assign v_2174 = v_2106 & v_2173;
assign v_2183 = v_2089 & v_2182;
assign v_2184 = v_2092 & v_2183;
assign v_2185 = v_2099 & v_2184;
assign v_2186 = v_2106 & v_2185;
assign v_2195 = v_2089 & v_2194;
assign v_2196 = v_2087 & v_2114;
assign v_2198 = v_2092 & v_2197;
assign v_2199 = ~v_91 & v_2116;
assign v_2201 = v_2099 & v_2200;
assign v_2202 = v_2097 & v_2123;
assign v_2204 = v_2106 & v_2203;
assign v_2205 = v_2104 & v_2130;
assign v_2210 = v_2208 & v_2209;
assign v_2213 = v_2211 & v_2212;
assign v_2216 = v_2214 & v_2215;
assign v_2219 = v_2217 & v_2218;
assign v_2223 = v_2089 & v_2222;
assign v_2224 = v_2092 & v_2223;
assign v_2225 = v_2099 & v_2224;
assign v_2226 = v_2106 & v_2225;
assign v_2236 = v_2234 & v_2235;
assign v_2238 = v_2236 & v_2237;
assign v_2241 = v_2239 & v_2240;
assign v_2243 = v_2238 & v_2242;
assign v_2246 = v_2244 & v_2245;
assign v_2248 = v_2243 & v_2247;
assign v_2250 = v_96 & v_2110;
assign v_2252 = v_807 & v_1823;
assign v_2254 = v_91 & v_2118;
assign v_2255 = v_91 & v_2120;
assign v_2257 = v_361 & v_2256;
assign v_2259 = v_91 & v_2125;
assign v_2260 = v_91 & v_2127;
assign v_2262 = v_563 & v_2261;
assign v_2267 = v_2234 & v_2266;
assign v_2268 = v_2237 & v_2267;
assign v_2269 = v_2242 & v_2268;
assign v_2270 = v_2247 & v_2269;
assign v_2279 = v_2234 & v_2278;
assign v_2280 = v_2237 & v_2279;
assign v_2281 = v_2242 & v_2280;
assign v_2282 = v_2247 & v_2281;
assign v_2291 = v_2234 & v_2290;
assign v_2292 = v_2237 & v_2291;
assign v_2293 = v_2242 & v_2292;
assign v_2294 = v_2247 & v_2293;
assign v_2303 = v_2234 & v_2302;
assign v_2304 = v_2237 & v_2303;
assign v_2305 = v_2242 & v_2304;
assign v_2306 = v_2247 & v_2305;
assign v_2315 = v_2234 & v_2314;
assign v_2316 = v_2237 & v_2315;
assign v_2317 = v_2242 & v_2316;
assign v_2318 = v_2247 & v_2317;
assign v_2327 = v_2234 & v_2326;
assign v_2328 = v_91 & v_2250;
assign v_2330 = v_2237 & v_2329;
assign v_2331 = v_1789 & v_2252;
assign v_2333 = v_2242 & v_2332;
assign v_2334 = v_2240 & v_2257;
assign v_2336 = v_2247 & v_2335;
assign v_2337 = v_2245 & v_2262;
assign v_2342 = v_2340 & v_2341;
assign v_2345 = v_2343 & v_2344;
assign v_2348 = v_2346 & v_2347;
assign v_2351 = v_2349 & v_2350;
assign v_2355 = v_2234 & v_2354;
assign v_2356 = v_2237 & v_2355;
assign v_2357 = v_2242 & v_2356;
assign v_2358 = v_2247 & v_2357;
assign v_2369 = v_2367 & v_2368;
assign v_2372 = v_2370 & v_2371;
assign v_2374 = v_2372 & v_2373;
assign v_2381 = v_2377 & v_2380;
assign v_2383 = v_2374 & v_2382;
assign v_2390 = v_2386 & v_2389;
assign v_2392 = v_2383 & v_2391;
assign v_2394 = v_89 & v_2109;
assign v_2395 = ~v_91 & v_2394;
assign v_2396 = v_91 & v_2110;
assign v_2398 = v_96 & v_2397;
assign v_2400 = v_807 & v_1820;
assign v_2402 = ~v_87 & v_1828;
assign v_2403 = ~v_89 & v_2402;
assign v_2404 = ~v_91 & v_2403;
assign v_2405 = ~v_87 & v_1832;
assign v_2406 = ~v_89 & v_2405;
assign v_2407 = ~v_91 & v_2406;
assign v_2409 = v_361 & v_2408;
assign v_2411 = ~v_87 & v_1839;
assign v_2412 = ~v_89 & v_2411;
assign v_2413 = ~v_91 & v_2412;
assign v_2414 = ~v_87 & v_1843;
assign v_2415 = ~v_89 & v_2414;
assign v_2416 = ~v_91 & v_2415;
assign v_2418 = v_563 & v_2417;
assign v_2423 = v_2370 & v_2422;
assign v_2424 = v_2373 & v_2423;
assign v_2425 = v_2382 & v_2424;
assign v_2426 = v_2391 & v_2425;
assign v_2435 = v_2370 & v_2434;
assign v_2436 = v_2373 & v_2435;
assign v_2437 = v_2382 & v_2436;
assign v_2438 = v_2391 & v_2437;
assign v_2447 = v_2370 & v_2446;
assign v_2448 = v_2373 & v_2447;
assign v_2449 = v_2382 & v_2448;
assign v_2450 = v_2391 & v_2449;
assign v_2459 = v_2370 & v_2458;
assign v_2460 = v_2373 & v_2459;
assign v_2461 = v_2382 & v_2460;
assign v_2462 = v_2391 & v_2461;
assign v_2471 = v_2370 & v_2470;
assign v_2472 = v_2373 & v_2471;
assign v_2473 = v_2382 & v_2472;
assign v_2474 = v_2391 & v_2473;
assign v_2483 = v_2370 & v_2482;
assign v_2484 = v_2368 & v_2398;
assign v_2486 = v_2373 & v_2485;
assign v_2487 = ~v_91 & v_2400;
assign v_2489 = v_2382 & v_2488;
assign v_2490 = v_2380 & v_2409;
assign v_2492 = v_2391 & v_2491;
assign v_2493 = v_2389 & v_2418;
assign v_2498 = v_2496 & v_2497;
assign v_2501 = v_2499 & v_2500;
assign v_2504 = v_2502 & v_2503;
assign v_2507 = v_2505 & v_2506;
assign v_2516 = v_2370 & ~v_2510;
assign v_2517 = v_2373 & v_2516;
assign v_2518 = v_2382 & v_2517;
assign v_2519 = v_2391 & v_2518;
assign v_2524 = v_2522 & v_2523;
assign v_2526 = v_2524 & v_2525;
assign v_2529 = v_2527 & v_2528;
assign v_2531 = v_2526 & v_2530;
assign v_2534 = v_2532 & v_2533;
assign v_2536 = v_2531 & v_2535;
assign v_2538 = v_96 & v_2394;
assign v_2540 = v_807 & v_2113;
assign v_2542 = v_91 & v_2403;
assign v_2543 = v_91 & v_2406;
assign v_2545 = v_361 & v_2544;
assign v_2547 = v_91 & v_2412;
assign v_2548 = v_91 & v_2415;
assign v_2550 = v_563 & v_2549;
assign v_2555 = v_2522 & v_2554;
assign v_2556 = v_2525 & v_2555;
assign v_2557 = v_2530 & v_2556;
assign v_2558 = v_2535 & v_2557;
assign v_2567 = v_2522 & v_2566;
assign v_2568 = v_2525 & v_2567;
assign v_2569 = v_2530 & v_2568;
assign v_2570 = v_2535 & v_2569;
assign v_2579 = v_2522 & v_2578;
assign v_2580 = v_2525 & v_2579;
assign v_2581 = v_2530 & v_2580;
assign v_2582 = v_2535 & v_2581;
assign v_2591 = v_2522 & v_2590;
assign v_2592 = v_2525 & v_2591;
assign v_2593 = v_2530 & v_2592;
assign v_2594 = v_2535 & v_2593;
assign v_2603 = v_2522 & v_2602;
assign v_2604 = v_2525 & v_2603;
assign v_2605 = v_2530 & v_2604;
assign v_2606 = v_2535 & v_2605;
assign v_2615 = v_2522 & v_2614;
assign v_2616 = v_91 & v_2538;
assign v_2618 = v_2525 & v_2617;
assign v_2619 = v_2086 & v_2540;
assign v_2621 = v_2530 & v_2620;
assign v_2622 = v_2528 & v_2545;
assign v_2624 = v_2535 & v_2623;
assign v_2625 = v_2533 & v_2550;
assign v_2630 = v_2628 & v_2629;
assign v_2633 = v_2631 & v_2632;
assign v_2636 = v_2634 & v_2635;
assign v_2639 = v_2637 & v_2638;
assign v_2648 = v_2522 & ~v_2642;
assign v_2649 = v_2525 & v_2648;
assign v_2650 = v_2530 & v_2649;
assign v_2651 = v_2535 & v_2650;
assign v_2660 = v_2658 & v_2659;
assign v_2663 = v_2661 & v_2662;
assign v_2665 = v_2663 & v_2664;
assign v_2670 = v_2667 & v_2669;
assign v_2672 = v_2665 & v_2671;
assign v_2677 = v_2674 & v_2676;
assign v_2679 = v_2672 & v_2678;
assign v_2681 = v_82 & v_582;
assign v_2682 = v_587 & v_2681;
assign v_2683 = v_87 & v_2682;
assign v_2684 = ~v_89 & v_2683;
assign v_2685 = ~v_91 & v_2684;
assign v_2686 = v_91 & v_2394;
assign v_2688 = v_96 & v_2687;
assign v_2690 = v_807 & v_2110;
assign v_2692 = v_89 & v_2402;
assign v_2693 = ~v_91 & v_2692;
assign v_2694 = v_89 & v_2405;
assign v_2695 = ~v_91 & v_2694;
assign v_2697 = v_361 & v_2696;
assign v_2699 = v_89 & v_2411;
assign v_2700 = ~v_91 & v_2699;
assign v_2701 = v_89 & v_2414;
assign v_2702 = ~v_91 & v_2701;
assign v_2704 = v_563 & v_2703;
assign v_2709 = v_2661 & v_2708;
assign v_2710 = v_2664 & v_2709;
assign v_2711 = v_2671 & v_2710;
assign v_2712 = v_2678 & v_2711;
assign v_2721 = v_2661 & v_2720;
assign v_2722 = v_2664 & v_2721;
assign v_2723 = v_2671 & v_2722;
assign v_2724 = v_2678 & v_2723;
assign v_2733 = v_2661 & v_2732;
assign v_2734 = v_2664 & v_2733;
assign v_2735 = v_2671 & v_2734;
assign v_2736 = v_2678 & v_2735;
assign v_2745 = v_2661 & v_2744;
assign v_2746 = v_2664 & v_2745;
assign v_2747 = v_2671 & v_2746;
assign v_2748 = v_2678 & v_2747;
assign v_2757 = v_2661 & v_2756;
assign v_2758 = v_2664 & v_2757;
assign v_2759 = v_2671 & v_2758;
assign v_2760 = v_2678 & v_2759;
assign v_2769 = v_2661 & v_2768;
assign v_2770 = v_2659 & v_2688;
assign v_2772 = v_2664 & v_2771;
assign v_2773 = ~v_91 & v_2690;
assign v_2775 = v_2671 & v_2774;
assign v_2776 = v_2669 & v_2697;
assign v_2778 = v_2678 & v_2777;
assign v_2779 = v_2676 & v_2704;
assign v_2784 = v_2782 & v_2783;
assign v_2787 = v_2785 & v_2786;
assign v_2790 = v_2788 & v_2789;
assign v_2793 = v_2791 & v_2792;
assign v_2802 = v_2661 & ~v_2796;
assign v_2803 = v_2664 & v_2802;
assign v_2804 = v_2671 & v_2803;
assign v_2805 = v_2678 & v_2804;
assign v_2810 = v_2808 & v_2809;
assign v_2812 = v_2810 & v_2811;
assign v_2815 = v_2813 & v_2814;
assign v_2817 = v_2812 & v_2816;
assign v_2820 = v_2818 & v_2819;
assign v_2822 = v_2817 & v_2821;
assign v_2824 = v_96 & v_2684;
assign v_2826 = v_807 & v_2397;
assign v_2828 = v_91 & v_2692;
assign v_2829 = v_91 & v_2694;
assign v_2831 = v_361 & v_2830;
assign v_2833 = v_91 & v_2699;
assign v_2834 = v_91 & v_2701;
assign v_2836 = v_563 & v_2835;
assign v_2841 = v_2808 & v_2840;
assign v_2842 = v_2811 & v_2841;
assign v_2843 = v_2816 & v_2842;
assign v_2844 = v_2821 & v_2843;
assign v_2853 = v_2808 & v_2852;
assign v_2854 = v_2811 & v_2853;
assign v_2855 = v_2816 & v_2854;
assign v_2856 = v_2821 & v_2855;
assign v_2865 = v_2808 & v_2864;
assign v_2866 = v_2811 & v_2865;
assign v_2867 = v_2816 & v_2866;
assign v_2868 = v_2821 & v_2867;
assign v_2877 = v_2808 & v_2876;
assign v_2878 = v_2811 & v_2877;
assign v_2879 = v_2816 & v_2878;
assign v_2880 = v_2821 & v_2879;
assign v_2889 = v_2808 & v_2888;
assign v_2890 = v_2811 & v_2889;
assign v_2891 = v_2816 & v_2890;
assign v_2892 = v_2821 & v_2891;
assign v_2901 = v_2808 & v_2900;
assign v_2902 = v_91 & v_2824;
assign v_2904 = v_2811 & v_2903;
assign v_2905 = v_2367 & v_2826;
assign v_2907 = v_2816 & v_2906;
assign v_2908 = v_2814 & v_2831;
assign v_2910 = v_2821 & v_2909;
assign v_2911 = v_2819 & v_2836;
assign v_2916 = v_2914 & v_2915;
assign v_2919 = v_2917 & v_2918;
assign v_2922 = v_2920 & v_2921;
assign v_2925 = v_2923 & v_2924;
assign v_2934 = v_2808 & ~v_2928;
assign v_2935 = v_2811 & v_2934;
assign v_2936 = v_2816 & v_2935;
assign v_2937 = v_2821 & v_2936;
assign v_2943 = v_2941 & v_2942;
assign v_2946 = v_2944 & v_2945;
assign v_2948 = v_2946 & v_2947;
assign v_2959 = v_2953 & v_2958;
assign v_2961 = v_2948 & v_2960;
assign v_2972 = v_2966 & v_2971;
assign v_2974 = v_2961 & v_2973;
assign v_2976 = v_89 & v_2683;
assign v_2977 = ~v_91 & v_2976;
assign v_2978 = v_91 & v_2684;
assign v_2980 = v_96 & v_2979;
assign v_2982 = v_807 & v_2394;
assign v_2984 = v_218 & v_619;
assign v_2985 = v_587 & v_2984;
assign v_2986 = v_87 & v_2985;
assign v_2987 = ~v_89 & v_2986;
assign v_2988 = ~v_91 & v_2987;
assign v_2989 = v_352 & v_649;
assign v_2990 = v_654 & v_2989;
assign v_2991 = v_87 & v_2990;
assign v_2992 = ~v_89 & v_2991;
assign v_2993 = ~v_91 & v_2992;
assign v_2995 = v_361 & v_2994;
assign v_2997 = v_218 & v_682;
assign v_2998 = v_587 & v_2997;
assign v_2999 = v_87 & v_2998;
assign v_3000 = ~v_89 & v_2999;
assign v_3001 = ~v_91 & v_3000;
assign v_3002 = v_556 & v_708;
assign v_3003 = v_654 & v_3002;
assign v_3004 = v_87 & v_3003;
assign v_3005 = ~v_89 & v_3004;
assign v_3006 = ~v_91 & v_3005;
assign v_3008 = v_563 & v_3007;
assign v_3013 = v_2944 & v_3012;
assign v_3014 = v_2947 & v_3013;
assign v_3015 = v_2960 & v_3014;
assign v_3016 = v_2973 & v_3015;
assign v_3025 = v_2944 & v_3024;
assign v_3026 = v_2947 & v_3025;
assign v_3027 = v_2960 & v_3026;
assign v_3028 = v_2973 & v_3027;
assign v_3037 = v_2944 & v_3036;
assign v_3038 = v_2947 & v_3037;
assign v_3039 = v_2960 & v_3038;
assign v_3040 = v_2973 & v_3039;
assign v_3049 = v_2944 & v_3048;
assign v_3050 = v_2947 & v_3049;
assign v_3051 = v_2960 & v_3050;
assign v_3052 = v_2973 & v_3051;
assign v_3061 = v_2944 & v_3060;
assign v_3062 = v_2947 & v_3061;
assign v_3063 = v_2960 & v_3062;
assign v_3064 = v_2973 & v_3063;
assign v_3073 = v_2944 & v_3072;
assign v_3074 = v_2942 & v_2980;
assign v_3076 = v_2947 & v_3075;
assign v_3077 = ~v_91 & v_2982;
assign v_3079 = v_2960 & v_3078;
assign v_3080 = v_2958 & v_2995;
assign v_3082 = v_2973 & v_3081;
assign v_3083 = v_2971 & v_3008;
assign v_3088 = v_3086 & v_3087;
assign v_3091 = v_3089 & v_3090;
assign v_3094 = v_3092 & v_3093;
assign v_3097 = v_3095 & v_3096;
assign v_3106 = v_2944 & ~v_3100;
assign v_3107 = v_2947 & v_3106;
assign v_3108 = v_2960 & v_3107;
assign v_3109 = v_2973 & v_3108;
assign v_3114 = v_3112 & v_3113;
assign v_3116 = v_3114 & v_3115;
assign v_3119 = v_3117 & v_3118;
assign v_3121 = v_3116 & v_3120;
assign v_3124 = v_3122 & v_3123;
assign v_3126 = v_3121 & v_3125;
assign v_3128 = v_96 & v_2976;
assign v_3130 = v_807 & v_2687;
assign v_3132 = v_91 & v_2987;
assign v_3133 = v_91 & v_2992;
assign v_3135 = v_361 & v_3134;
assign v_3137 = v_91 & v_3000;
assign v_3138 = v_91 & v_3005;
assign v_3140 = v_563 & v_3139;
assign v_3145 = v_3112 & v_3144;
assign v_3146 = v_3115 & v_3145;
assign v_3147 = v_3120 & v_3146;
assign v_3148 = v_3125 & v_3147;
assign v_3157 = v_3112 & v_3156;
assign v_3158 = v_3115 & v_3157;
assign v_3159 = v_3120 & v_3158;
assign v_3160 = v_3125 & v_3159;
assign v_3169 = v_3112 & v_3168;
assign v_3170 = v_3115 & v_3169;
assign v_3171 = v_3120 & v_3170;
assign v_3172 = v_3125 & v_3171;
assign v_3181 = v_3112 & v_3180;
assign v_3182 = v_3115 & v_3181;
assign v_3183 = v_3120 & v_3182;
assign v_3184 = v_3125 & v_3183;
assign v_3193 = v_3112 & v_3192;
assign v_3194 = v_3115 & v_3193;
assign v_3195 = v_3120 & v_3194;
assign v_3196 = v_3125 & v_3195;
assign v_3207 = v_3205 & v_3206;
assign v_3210 = v_3208 & v_3209;
assign v_3213 = v_3211 & v_3212;
assign v_3216 = v_3214 & v_3215;
assign v_3218 = v_3112 & ~v_3204;
assign v_3219 = v_91 & v_3128;
assign v_3221 = v_3115 & v_3220;
assign v_3222 = v_2658 & v_3130;
assign v_3224 = v_3120 & v_3223;
assign v_3225 = v_3118 & v_3135;
assign v_3227 = v_3125 & v_3226;
assign v_3228 = v_3123 & v_3140;
assign v_3233 = v_3112 & v_3232;
assign v_3234 = v_3115 & v_3233;
assign v_3235 = v_3120 & v_3234;
assign v_3236 = v_3125 & v_3235;
assign v_3248 = v_3246 & v_3247;
assign v_3251 = v_3249 & v_3250;
assign v_3253 = v_3251 & v_3252;
assign v_3258 = v_3255 & v_3257;
assign v_3260 = v_3253 & v_3259;
assign v_3265 = v_3262 & v_3264;
assign v_3267 = v_3260 & v_3266;
assign v_3269 = ~v_87 & v_2682;
assign v_3270 = ~v_89 & v_3269;
assign v_3271 = ~v_91 & v_3270;
assign v_3272 = v_91 & v_2976;
assign v_3274 = v_96 & v_3273;
assign v_3276 = v_807 & v_2684;
assign v_3278 = v_89 & v_2986;
assign v_3279 = ~v_91 & v_3278;
assign v_3280 = v_89 & v_2991;
assign v_3281 = ~v_91 & v_3280;
assign v_3283 = v_361 & v_3282;
assign v_3285 = v_89 & v_2999;
assign v_3286 = ~v_91 & v_3285;
assign v_3287 = v_89 & v_3004;
assign v_3288 = ~v_91 & v_3287;
assign v_3290 = v_563 & v_3289;
assign v_3295 = v_3249 & v_3294;
assign v_3296 = v_3252 & v_3295;
assign v_3297 = v_3259 & v_3296;
assign v_3298 = v_3266 & v_3297;
assign v_3307 = v_3249 & v_3306;
assign v_3308 = v_3252 & v_3307;
assign v_3309 = v_3259 & v_3308;
assign v_3310 = v_3266 & v_3309;
assign v_3319 = v_3249 & v_3318;
assign v_3320 = v_3252 & v_3319;
assign v_3321 = v_3259 & v_3320;
assign v_3322 = v_3266 & v_3321;
assign v_3331 = v_3249 & v_3330;
assign v_3332 = v_3252 & v_3331;
assign v_3333 = v_3259 & v_3332;
assign v_3334 = v_3266 & v_3333;
assign v_3343 = v_3249 & v_3342;
assign v_3344 = v_3252 & v_3343;
assign v_3345 = v_3259 & v_3344;
assign v_3346 = v_3266 & v_3345;
assign v_3355 = v_3249 & v_3354;
assign v_3356 = v_3247 & v_3274;
assign v_3358 = v_3252 & v_3357;
assign v_3359 = ~v_91 & v_3276;
assign v_3361 = v_3259 & v_3360;
assign v_3362 = v_3257 & v_3283;
assign v_3364 = v_3266 & v_3363;
assign v_3365 = v_3264 & v_3290;
assign v_3370 = v_3368 & v_3369;
assign v_3373 = v_3371 & v_3372;
assign v_3376 = v_3374 & v_3375;
assign v_3379 = v_3377 & v_3378;
assign v_3388 = v_3249 & ~v_3382;
assign v_3389 = v_3252 & v_3388;
assign v_3390 = v_3259 & v_3389;
assign v_3391 = v_3266 & v_3390;
assign v_3396 = v_3394 & v_3395;
assign v_3398 = v_3396 & v_3397;
assign v_3401 = v_3399 & v_3400;
assign v_3403 = v_3398 & v_3402;
assign v_3406 = v_3404 & v_3405;
assign v_3408 = v_3403 & v_3407;
assign v_3410 = v_96 & v_3270;
assign v_3412 = v_807 & v_2979;
assign v_3414 = v_91 & v_3278;
assign v_3415 = v_91 & v_3280;
assign v_3417 = v_361 & v_3416;
assign v_3419 = v_91 & v_3285;
assign v_3420 = v_91 & v_3287;
assign v_3422 = v_563 & v_3421;
assign v_3427 = v_3394 & v_3426;
assign v_3428 = v_3397 & v_3427;
assign v_3429 = v_3402 & v_3428;
assign v_3430 = v_3407 & v_3429;
assign v_3439 = v_3394 & v_3438;
assign v_3440 = v_3397 & v_3439;
assign v_3441 = v_3402 & v_3440;
assign v_3442 = v_3407 & v_3441;
assign v_3451 = v_3394 & v_3450;
assign v_3452 = v_3397 & v_3451;
assign v_3453 = v_3402 & v_3452;
assign v_3454 = v_3407 & v_3453;
assign v_3463 = v_3394 & v_3462;
assign v_3464 = v_3397 & v_3463;
assign v_3465 = v_3402 & v_3464;
assign v_3466 = v_3407 & v_3465;
assign v_3475 = v_3394 & v_3474;
assign v_3476 = v_3397 & v_3475;
assign v_3477 = v_3402 & v_3476;
assign v_3478 = v_3407 & v_3477;
assign v_3487 = v_3394 & v_3486;
assign v_3488 = v_91 & v_3410;
assign v_3490 = v_3397 & v_3489;
assign v_3491 = v_2941 & v_3412;
assign v_3493 = v_3402 & v_3492;
assign v_3494 = v_3400 & v_3417;
assign v_3496 = v_3407 & v_3495;
assign v_3497 = v_3405 & v_3422;
assign v_3502 = v_3500 & v_3501;
assign v_3505 = v_3503 & v_3504;
assign v_3508 = v_3506 & v_3507;
assign v_3511 = v_3509 & v_3510;
assign v_3515 = v_3394 & v_3514;
assign v_3516 = v_3397 & v_3515;
assign v_3517 = v_3402 & v_3516;
assign v_3518 = v_3407 & v_3517;
assign v_3529 = v_3527 & v_3528;
assign v_3532 = v_3530 & v_3531;
assign v_3534 = v_3532 & v_3533;
assign v_3541 = v_3537 & v_3540;
assign v_3543 = v_3534 & v_3542;
assign v_3550 = v_3546 & v_3549;
assign v_3552 = v_3543 & v_3551;
assign v_3554 = v_89 & v_3269;
assign v_3555 = ~v_91 & v_3554;
assign v_3556 = v_91 & v_3270;
assign v_3558 = v_96 & v_3557;
assign v_3560 = v_807 & v_2976;
assign v_3562 = ~v_87 & v_2985;
assign v_3563 = ~v_89 & v_3562;
assign v_3564 = ~v_91 & v_3563;
assign v_3565 = ~v_87 & v_2990;
assign v_3566 = ~v_89 & v_3565;
assign v_3567 = ~v_91 & v_3566;
assign v_3569 = v_361 & v_3568;
assign v_3571 = ~v_87 & v_2998;
assign v_3572 = ~v_89 & v_3571;
assign v_3573 = ~v_91 & v_3572;
assign v_3574 = ~v_87 & v_3003;
assign v_3575 = ~v_89 & v_3574;
assign v_3576 = ~v_91 & v_3575;
assign v_3578 = v_563 & v_3577;
assign v_3583 = v_3530 & v_3582;
assign v_3584 = v_3533 & v_3583;
assign v_3585 = v_3542 & v_3584;
assign v_3586 = v_3551 & v_3585;
assign v_3595 = v_3530 & v_3594;
assign v_3596 = v_3533 & v_3595;
assign v_3597 = v_3542 & v_3596;
assign v_3598 = v_3551 & v_3597;
assign v_3607 = v_3530 & v_3606;
assign v_3608 = v_3533 & v_3607;
assign v_3609 = v_3542 & v_3608;
assign v_3610 = v_3551 & v_3609;
assign v_3619 = v_3530 & v_3618;
assign v_3620 = v_3533 & v_3619;
assign v_3621 = v_3542 & v_3620;
assign v_3622 = v_3551 & v_3621;
assign v_3631 = v_3530 & v_3630;
assign v_3632 = v_3533 & v_3631;
assign v_3633 = v_3542 & v_3632;
assign v_3634 = v_3551 & v_3633;
assign v_3643 = v_3530 & v_3642;
assign v_3644 = v_3528 & v_3558;
assign v_3646 = v_3533 & v_3645;
assign v_3647 = ~v_91 & v_3560;
assign v_3649 = v_3542 & v_3648;
assign v_3650 = v_3540 & v_3569;
assign v_3652 = v_3551 & v_3651;
assign v_3653 = v_3549 & v_3578;
assign v_3658 = v_3656 & v_3657;
assign v_3661 = v_3659 & v_3660;
assign v_3664 = v_3662 & v_3663;
assign v_3667 = v_3665 & v_3666;
assign v_3676 = v_3530 & ~v_3670;
assign v_3677 = v_3533 & v_3676;
assign v_3678 = v_3542 & v_3677;
assign v_3679 = v_3551 & v_3678;
assign v_3684 = v_3682 & v_3683;
assign v_3686 = v_3684 & v_3685;
assign v_3689 = v_3687 & v_3688;
assign v_3691 = v_3686 & v_3690;
assign v_3694 = v_3692 & v_3693;
assign v_3696 = v_3691 & v_3695;
assign v_3698 = v_96 & v_3554;
assign v_3700 = v_807 & v_3273;
assign v_3702 = v_91 & v_3563;
assign v_3703 = v_91 & v_3566;
assign v_3705 = v_361 & v_3704;
assign v_3707 = v_91 & v_3572;
assign v_3708 = v_91 & v_3575;
assign v_3710 = v_563 & v_3709;
assign v_3715 = v_3682 & v_3714;
assign v_3716 = v_3685 & v_3715;
assign v_3717 = v_3690 & v_3716;
assign v_3718 = v_3695 & v_3717;
assign v_3727 = v_3682 & v_3726;
assign v_3728 = v_3685 & v_3727;
assign v_3729 = v_3690 & v_3728;
assign v_3730 = v_3695 & v_3729;
assign v_3739 = v_3682 & v_3738;
assign v_3740 = v_3685 & v_3739;
assign v_3741 = v_3690 & v_3740;
assign v_3742 = v_3695 & v_3741;
assign v_3751 = v_3682 & v_3750;
assign v_3752 = v_3685 & v_3751;
assign v_3753 = v_3690 & v_3752;
assign v_3754 = v_3695 & v_3753;
assign v_3763 = v_3682 & v_3762;
assign v_3764 = v_3685 & v_3763;
assign v_3765 = v_3690 & v_3764;
assign v_3766 = v_3695 & v_3765;
assign v_3775 = v_3682 & v_3774;
assign v_3776 = v_91 & v_3698;
assign v_3778 = v_3685 & v_3777;
assign v_3779 = v_3246 & v_3700;
assign v_3781 = v_3690 & v_3780;
assign v_3782 = v_3688 & v_3705;
assign v_3784 = v_3695 & v_3783;
assign v_3785 = v_3693 & v_3710;
assign v_3790 = v_3788 & v_3789;
assign v_3793 = v_3791 & v_3792;
assign v_3796 = v_3794 & v_3795;
assign v_3799 = v_3797 & v_3798;
assign v_3808 = v_3682 & ~v_3802;
assign v_3809 = v_3685 & v_3808;
assign v_3810 = v_3690 & v_3809;
assign v_3811 = v_3695 & v_3810;
assign v_3819 = v_3817 & v_3818;
assign v_3822 = v_3820 & v_3821;
assign v_3824 = v_3822 & v_3823;
assign v_3829 = v_3826 & v_3828;
assign v_3831 = v_3824 & v_3830;
assign v_3836 = v_3833 & v_3835;
assign v_3838 = v_3831 & v_3837;
assign v_3840 = v_85 & v_2681;
assign v_3841 = v_87 & v_3840;
assign v_3842 = ~v_89 & v_3841;
assign v_3843 = ~v_91 & v_3842;
assign v_3844 = v_91 & v_3554;
assign v_3846 = v_96 & v_3845;
assign v_3848 = v_807 & v_3270;
assign v_3850 = v_89 & v_3562;
assign v_3851 = ~v_91 & v_3850;
assign v_3852 = v_89 & v_3565;
assign v_3853 = ~v_91 & v_3852;
assign v_3855 = v_361 & v_3854;
assign v_3857 = v_89 & v_3571;
assign v_3858 = ~v_91 & v_3857;
assign v_3859 = v_89 & v_3574;
assign v_3860 = ~v_91 & v_3859;
assign v_3862 = v_563 & v_3861;
assign v_3867 = v_3820 & v_3866;
assign v_3868 = v_3823 & v_3867;
assign v_3869 = v_3830 & v_3868;
assign v_3870 = v_3837 & v_3869;
assign v_3879 = v_3820 & v_3878;
assign v_3880 = v_3823 & v_3879;
assign v_3881 = v_3830 & v_3880;
assign v_3882 = v_3837 & v_3881;
assign v_3891 = v_3820 & v_3890;
assign v_3892 = v_3823 & v_3891;
assign v_3893 = v_3830 & v_3892;
assign v_3894 = v_3837 & v_3893;
assign v_3903 = v_3820 & v_3902;
assign v_3904 = v_3823 & v_3903;
assign v_3905 = v_3830 & v_3904;
assign v_3906 = v_3837 & v_3905;
assign v_3915 = v_3820 & v_3914;
assign v_3916 = v_3823 & v_3915;
assign v_3917 = v_3830 & v_3916;
assign v_3918 = v_3837 & v_3917;
assign v_3927 = v_3820 & v_3926;
assign v_3928 = v_3818 & v_3846;
assign v_3930 = v_3823 & v_3929;
assign v_3931 = ~v_91 & v_3848;
assign v_3933 = v_3830 & v_3932;
assign v_3934 = v_3828 & v_3855;
assign v_3936 = v_3837 & v_3935;
assign v_3937 = v_3835 & v_3862;
assign v_3942 = v_3940 & v_3941;
assign v_3945 = v_3943 & v_3944;
assign v_3948 = v_3946 & v_3947;
assign v_3951 = v_3949 & v_3950;
assign v_3960 = v_3820 & ~v_3954;
assign v_3961 = v_3823 & v_3960;
assign v_3962 = v_3830 & v_3961;
assign v_3963 = v_3837 & v_3962;
assign v_3968 = v_3966 & v_3967;
assign v_3970 = v_3968 & v_3969;
assign v_3973 = v_3971 & v_3972;
assign v_3975 = v_3970 & v_3974;
assign v_3978 = v_3976 & v_3977;
assign v_3980 = v_3975 & v_3979;
assign v_3982 = v_96 & v_3842;
assign v_3984 = v_807 & v_3557;
assign v_3986 = v_91 & v_3850;
assign v_3987 = v_91 & v_3852;
assign v_3989 = v_361 & v_3988;
assign v_3991 = v_91 & v_3857;
assign v_3992 = v_91 & v_3859;
assign v_3994 = v_563 & v_3993;
assign v_3999 = v_3966 & v_3998;
assign v_4000 = v_3969 & v_3999;
assign v_4001 = v_3974 & v_4000;
assign v_4002 = v_3979 & v_4001;
assign v_4011 = v_3966 & v_4010;
assign v_4012 = v_3969 & v_4011;
assign v_4013 = v_3974 & v_4012;
assign v_4014 = v_3979 & v_4013;
assign v_4023 = v_3966 & v_4022;
assign v_4024 = v_3969 & v_4023;
assign v_4025 = v_3974 & v_4024;
assign v_4026 = v_3979 & v_4025;
assign v_4035 = v_3966 & v_4034;
assign v_4036 = v_3969 & v_4035;
assign v_4037 = v_3974 & v_4036;
assign v_4038 = v_3979 & v_4037;
assign v_4047 = v_3966 & v_4046;
assign v_4048 = v_3969 & v_4047;
assign v_4049 = v_3974 & v_4048;
assign v_4050 = v_3979 & v_4049;
assign v_4059 = v_3966 & v_4058;
assign v_4060 = v_91 & v_3982;
assign v_4062 = v_3969 & v_4061;
assign v_4063 = v_3527 & v_3984;
assign v_4065 = v_3974 & v_4064;
assign v_4066 = v_3972 & v_3989;
assign v_4068 = v_3979 & v_4067;
assign v_4069 = v_3977 & v_3994;
assign v_4074 = v_4072 & v_4073;
assign v_4077 = v_4075 & v_4076;
assign v_4080 = v_4078 & v_4079;
assign v_4083 = v_4081 & v_4082;
assign v_4092 = v_3966 & ~v_4086;
assign v_4093 = v_3969 & v_4092;
assign v_4094 = v_3974 & v_4093;
assign v_4095 = v_3979 & v_4094;
assign v_4101 = v_4099 & v_4100;
assign v_4104 = v_4102 & v_4103;
assign v_4106 = v_4104 & v_4105;
assign v_4115 = v_4110 & v_4114;
assign v_4117 = v_4106 & v_4116;
assign v_4126 = v_4121 & v_4125;
assign v_4128 = v_4117 & v_4127;
assign v_4130 = v_89 & v_3841;
assign v_4131 = ~v_91 & v_4130;
assign v_4132 = v_91 & v_3842;
assign v_4134 = v_96 & v_4133;
assign v_4136 = v_807 & v_3554;
assign v_4138 = v_85 & v_2984;
assign v_4139 = v_87 & v_4138;
assign v_4140 = ~v_89 & v_4139;
assign v_4141 = ~v_91 & v_4140;
assign v_4142 = v_355 & v_2989;
assign v_4143 = v_87 & v_4142;
assign v_4144 = ~v_89 & v_4143;
assign v_4145 = ~v_91 & v_4144;
assign v_4147 = v_361 & v_4146;
assign v_4149 = v_85 & v_2997;
assign v_4150 = v_87 & v_4149;
assign v_4151 = ~v_89 & v_4150;
assign v_4152 = ~v_91 & v_4151;
assign v_4153 = v_355 & v_3002;
assign v_4154 = v_87 & v_4153;
assign v_4155 = ~v_89 & v_4154;
assign v_4156 = ~v_91 & v_4155;
assign v_4158 = v_563 & v_4157;
assign v_4163 = v_4102 & v_4162;
assign v_4164 = v_4105 & v_4163;
assign v_4165 = v_4116 & v_4164;
assign v_4166 = v_4127 & v_4165;
assign v_4175 = v_4102 & v_4174;
assign v_4176 = v_4105 & v_4175;
assign v_4177 = v_4116 & v_4176;
assign v_4178 = v_4127 & v_4177;
assign v_4187 = v_4102 & v_4186;
assign v_4188 = v_4105 & v_4187;
assign v_4189 = v_4116 & v_4188;
assign v_4190 = v_4127 & v_4189;
assign v_4199 = v_4102 & v_4198;
assign v_4200 = v_4105 & v_4199;
assign v_4201 = v_4116 & v_4200;
assign v_4202 = v_4127 & v_4201;
assign v_4211 = v_4102 & v_4210;
assign v_4212 = v_4105 & v_4211;
assign v_4213 = v_4116 & v_4212;
assign v_4214 = v_4127 & v_4213;
assign v_4223 = v_4102 & v_4222;
assign v_4224 = v_4100 & v_4134;
assign v_4226 = v_4105 & v_4225;
assign v_4227 = ~v_91 & v_4136;
assign v_4229 = v_4116 & v_4228;
assign v_4230 = v_4114 & v_4147;
assign v_4232 = v_4127 & v_4231;
assign v_4233 = v_4125 & v_4158;
assign v_4238 = v_4236 & v_4237;
assign v_4241 = v_4239 & v_4240;
assign v_4244 = v_4242 & v_4243;
assign v_4247 = v_4245 & v_4246;
assign v_4256 = v_4102 & ~v_4250;
assign v_4257 = v_4105 & v_4256;
assign v_4258 = v_4116 & v_4257;
assign v_4259 = v_4127 & v_4258;
assign v_4264 = v_4262 & v_4263;
assign v_4266 = v_4264 & v_4265;
assign v_4269 = v_4267 & v_4268;
assign v_4271 = v_4266 & v_4270;
assign v_4274 = v_4272 & v_4273;
assign v_4276 = v_4271 & v_4275;
assign v_4278 = v_96 & v_4130;
assign v_4280 = v_807 & v_3845;
assign v_4282 = v_91 & v_4140;
assign v_4283 = v_91 & v_4144;
assign v_4285 = v_361 & v_4284;
assign v_4287 = v_91 & v_4151;
assign v_4288 = v_91 & v_4155;
assign v_4290 = v_563 & v_4289;
assign v_4295 = v_4262 & v_4294;
assign v_4296 = v_4265 & v_4295;
assign v_4297 = v_4270 & v_4296;
assign v_4298 = v_4275 & v_4297;
assign v_4307 = v_4262 & v_4306;
assign v_4308 = v_4265 & v_4307;
assign v_4309 = v_4270 & v_4308;
assign v_4310 = v_4275 & v_4309;
assign v_4319 = v_4262 & v_4318;
assign v_4320 = v_4265 & v_4319;
assign v_4321 = v_4270 & v_4320;
assign v_4322 = v_4275 & v_4321;
assign v_4331 = v_4262 & v_4330;
assign v_4332 = v_4265 & v_4331;
assign v_4333 = v_4270 & v_4332;
assign v_4334 = v_4275 & v_4333;
assign v_4343 = v_4262 & v_4342;
assign v_4344 = v_4265 & v_4343;
assign v_4345 = v_4270 & v_4344;
assign v_4346 = v_4275 & v_4345;
assign v_4355 = v_4262 & v_4354;
assign v_4356 = v_91 & v_4278;
assign v_4358 = v_4265 & v_4357;
assign v_4359 = v_3817 & v_4280;
assign v_4361 = v_4270 & v_4360;
assign v_4362 = v_4268 & v_4285;
assign v_4364 = v_4275 & v_4363;
assign v_4365 = v_4273 & v_4290;
assign v_4370 = v_4368 & v_4369;
assign v_4373 = v_4371 & v_4372;
assign v_4376 = v_4374 & v_4375;
assign v_4379 = v_4377 & v_4378;
assign v_4383 = v_4262 & v_4382;
assign v_4384 = v_4265 & v_4383;
assign v_4385 = v_4270 & v_4384;
assign v_4386 = v_4275 & v_4385;
assign v_4398 = v_4396 & v_4397;
assign v_4401 = v_4399 & v_4400;
assign v_4403 = v_4401 & v_4402;
assign v_4408 = v_4405 & v_4407;
assign v_4410 = v_4403 & v_4409;
assign v_4415 = v_4412 & v_4414;
assign v_4417 = v_4410 & v_4416;
assign v_4419 = ~v_87 & v_3840;
assign v_4420 = ~v_89 & v_4419;
assign v_4421 = ~v_91 & v_4420;
assign v_4422 = v_91 & v_4130;
assign v_4424 = v_96 & v_4423;
assign v_4426 = v_807 & v_3842;
assign v_4428 = v_89 & v_4139;
assign v_4429 = ~v_91 & v_4428;
assign v_4430 = v_89 & v_4143;
assign v_4431 = ~v_91 & v_4430;
assign v_4433 = v_361 & v_4432;
assign v_4435 = v_89 & v_4150;
assign v_4436 = ~v_91 & v_4435;
assign v_4437 = v_89 & v_4154;
assign v_4438 = ~v_91 & v_4437;
assign v_4440 = v_563 & v_4439;
assign v_4445 = v_4399 & v_4444;
assign v_4446 = v_4402 & v_4445;
assign v_4447 = v_4409 & v_4446;
assign v_4448 = v_4416 & v_4447;
assign v_4457 = v_4399 & v_4456;
assign v_4458 = v_4402 & v_4457;
assign v_4459 = v_4409 & v_4458;
assign v_4460 = v_4416 & v_4459;
assign v_4469 = v_4399 & v_4468;
assign v_4470 = v_4402 & v_4469;
assign v_4471 = v_4409 & v_4470;
assign v_4472 = v_4416 & v_4471;
assign v_4481 = v_4399 & v_4480;
assign v_4482 = v_4402 & v_4481;
assign v_4483 = v_4409 & v_4482;
assign v_4484 = v_4416 & v_4483;
assign v_4493 = v_4399 & v_4492;
assign v_4494 = v_4402 & v_4493;
assign v_4495 = v_4409 & v_4494;
assign v_4496 = v_4416 & v_4495;
assign v_4505 = v_4399 & v_4504;
assign v_4506 = v_4397 & v_4424;
assign v_4508 = v_4402 & v_4507;
assign v_4509 = ~v_91 & v_4426;
assign v_4511 = v_4409 & v_4510;
assign v_4512 = v_4407 & v_4433;
assign v_4514 = v_4416 & v_4513;
assign v_4515 = v_4414 & v_4440;
assign v_4520 = v_4518 & v_4519;
assign v_4523 = v_4521 & v_4522;
assign v_4526 = v_4524 & v_4525;
assign v_4529 = v_4527 & v_4528;
assign v_4533 = v_4399 & v_4532;
assign v_4534 = v_4402 & v_4533;
assign v_4535 = v_4409 & v_4534;
assign v_4536 = v_4416 & v_4535;
assign v_4546 = v_4544 & v_4545;
assign v_4548 = v_4546 & v_4547;
assign v_4551 = v_4549 & v_4550;
assign v_4553 = v_4548 & v_4552;
assign v_4556 = v_4554 & v_4555;
assign v_4558 = v_4553 & v_4557;
assign v_4560 = v_96 & v_4420;
assign v_4562 = v_807 & v_4133;
assign v_4564 = v_91 & v_4428;
assign v_4565 = v_91 & v_4430;
assign v_4567 = v_361 & v_4566;
assign v_4569 = v_91 & v_4435;
assign v_4570 = v_91 & v_4437;
assign v_4572 = v_563 & v_4571;
assign v_4577 = v_4544 & v_4576;
assign v_4578 = v_4547 & v_4577;
assign v_4579 = v_4552 & v_4578;
assign v_4580 = v_4557 & v_4579;
assign v_4589 = v_4544 & v_4588;
assign v_4590 = v_4547 & v_4589;
assign v_4591 = v_4552 & v_4590;
assign v_4592 = v_4557 & v_4591;
assign v_4601 = v_4544 & v_4600;
assign v_4602 = v_4547 & v_4601;
assign v_4603 = v_4552 & v_4602;
assign v_4604 = v_4557 & v_4603;
assign v_4613 = v_4544 & v_4612;
assign v_4614 = v_4547 & v_4613;
assign v_4615 = v_4552 & v_4614;
assign v_4616 = v_4557 & v_4615;
assign v_4625 = v_4544 & v_4624;
assign v_4626 = v_4547 & v_4625;
assign v_4627 = v_4552 & v_4626;
assign v_4628 = v_4557 & v_4627;
assign v_4637 = v_4544 & v_4636;
assign v_4638 = v_91 & v_4560;
assign v_4640 = v_4547 & v_4639;
assign v_4641 = v_4099 & v_4562;
assign v_4643 = v_4552 & v_4642;
assign v_4644 = v_4550 & v_4567;
assign v_4646 = v_4557 & v_4645;
assign v_4647 = v_4555 & v_4572;
assign v_4652 = v_4650 & v_4651;
assign v_4655 = v_4653 & v_4654;
assign v_4658 = v_4656 & v_4657;
assign v_4661 = v_4659 & v_4660;
assign v_4665 = v_4544 & v_4664;
assign v_4666 = v_4547 & v_4665;
assign v_4667 = v_4552 & v_4666;
assign v_4668 = v_4557 & v_4667;
assign v_4679 = v_4677 & v_4678;
assign v_4682 = v_4680 & v_4681;
assign v_4684 = v_4682 & v_4683;
assign v_4691 = v_4687 & v_4690;
assign v_4693 = v_4684 & v_4692;
assign v_4700 = v_4696 & v_4699;
assign v_4702 = v_4693 & v_4701;
assign v_4704 = v_89 & v_4419;
assign v_4705 = ~v_91 & v_4704;
assign v_4706 = v_91 & v_4420;
assign v_4708 = v_96 & v_4707;
assign v_4710 = v_807 & v_4130;
assign v_4712 = ~v_87 & v_4138;
assign v_4713 = ~v_89 & v_4712;
assign v_4714 = ~v_91 & v_4713;
assign v_4715 = ~v_87 & v_4142;
assign v_4716 = ~v_89 & v_4715;
assign v_4717 = ~v_91 & v_4716;
assign v_4719 = v_361 & v_4718;
assign v_4721 = ~v_87 & v_4149;
assign v_4722 = ~v_89 & v_4721;
assign v_4723 = ~v_91 & v_4722;
assign v_4724 = ~v_87 & v_4153;
assign v_4725 = ~v_89 & v_4724;
assign v_4726 = ~v_91 & v_4725;
assign v_4728 = v_563 & v_4727;
assign v_4733 = v_4680 & v_4732;
assign v_4734 = v_4683 & v_4733;
assign v_4735 = v_4692 & v_4734;
assign v_4736 = v_4701 & v_4735;
assign v_4745 = v_4680 & v_4744;
assign v_4746 = v_4683 & v_4745;
assign v_4747 = v_4692 & v_4746;
assign v_4748 = v_4701 & v_4747;
assign v_4757 = v_4680 & v_4756;
assign v_4758 = v_4683 & v_4757;
assign v_4759 = v_4692 & v_4758;
assign v_4760 = v_4701 & v_4759;
assign v_4769 = v_4680 & v_4768;
assign v_4770 = v_4683 & v_4769;
assign v_4771 = v_4692 & v_4770;
assign v_4772 = v_4701 & v_4771;
assign v_4781 = v_4680 & v_4780;
assign v_4782 = v_4683 & v_4781;
assign v_4783 = v_4692 & v_4782;
assign v_4784 = v_4701 & v_4783;
assign v_4793 = v_4680 & v_4792;
assign v_4794 = v_4678 & v_4708;
assign v_4796 = v_4683 & v_4795;
assign v_4797 = ~v_91 & v_4710;
assign v_4799 = v_4692 & v_4798;
assign v_4800 = v_4690 & v_4719;
assign v_4802 = v_4701 & v_4801;
assign v_4803 = v_4699 & v_4728;
assign v_4808 = v_4806 & v_4807;
assign v_4811 = v_4809 & v_4810;
assign v_4814 = v_4812 & v_4813;
assign v_4817 = v_4815 & v_4816;
assign v_4821 = v_4680 & v_4820;
assign v_4822 = v_4683 & v_4821;
assign v_4823 = v_4692 & v_4822;
assign v_4824 = v_4701 & v_4823;
assign v_4834 = v_4832 & v_4833;
assign v_4836 = v_4834 & v_4835;
assign v_4839 = v_4837 & v_4838;
assign v_4841 = v_4836 & v_4840;
assign v_4844 = v_4842 & v_4843;
assign v_4846 = v_4841 & v_4845;
assign v_4848 = v_96 & v_4704;
assign v_4850 = v_807 & v_4423;
assign v_4852 = v_91 & v_4713;
assign v_4853 = v_91 & v_4716;
assign v_4855 = v_361 & v_4854;
assign v_4857 = v_91 & v_4722;
assign v_4858 = v_91 & v_4725;
assign v_4860 = v_563 & v_4859;
assign v_4865 = v_4832 & v_4864;
assign v_4866 = v_4835 & v_4865;
assign v_4867 = v_4840 & v_4866;
assign v_4868 = v_4845 & v_4867;
assign v_4877 = v_4832 & v_4876;
assign v_4878 = v_4835 & v_4877;
assign v_4879 = v_4840 & v_4878;
assign v_4880 = v_4845 & v_4879;
assign v_4889 = v_4832 & v_4888;
assign v_4890 = v_4835 & v_4889;
assign v_4891 = v_4840 & v_4890;
assign v_4892 = v_4845 & v_4891;
assign v_4901 = v_4832 & v_4900;
assign v_4902 = v_4835 & v_4901;
assign v_4903 = v_4840 & v_4902;
assign v_4904 = v_4845 & v_4903;
assign v_4913 = v_4832 & v_4912;
assign v_4914 = v_4835 & v_4913;
assign v_4915 = v_4840 & v_4914;
assign v_4916 = v_4845 & v_4915;
assign v_4925 = v_4832 & v_4924;
assign v_4926 = v_91 & v_4848;
assign v_4928 = v_4835 & v_4927;
assign v_4929 = v_4396 & v_4850;
assign v_4931 = v_4840 & v_4930;
assign v_4932 = v_4838 & v_4855;
assign v_4934 = v_4845 & v_4933;
assign v_4935 = v_4843 & v_4860;
assign v_4940 = v_4938 & v_4939;
assign v_4943 = v_4941 & v_4942;
assign v_4946 = v_4944 & v_4945;
assign v_4949 = v_4947 & v_4948;
assign v_4953 = v_4832 & v_4952;
assign v_4954 = v_4835 & v_4953;
assign v_4955 = v_4840 & v_4954;
assign v_4956 = v_4845 & v_4955;
assign v_4971 = v_4969 & v_4970;
assign v_4974 = v_4972 & v_4973;
assign v_4976 = v_4974 & v_4975;
assign v_4981 = v_4978 & v_4980;
assign v_4983 = v_4976 & v_4982;
assign v_4988 = v_4985 & v_4987;
assign v_4990 = v_4983 & v_4989;
assign v_4992 = v_79 & v_579;
assign v_4993 = v_584 & v_4992;
assign v_4994 = v_587 & v_4993;
assign v_4995 = v_87 & v_4994;
assign v_4996 = ~v_89 & v_4995;
assign v_4997 = ~v_91 & v_4996;
assign v_4998 = v_91 & v_4704;
assign v_5000 = v_96 & v_4999;
assign v_5002 = v_807 & v_4420;
assign v_5004 = v_89 & v_4712;
assign v_5005 = ~v_91 & v_5004;
assign v_5006 = v_89 & v_4715;
assign v_5007 = ~v_91 & v_5006;
assign v_5009 = v_361 & v_5008;
assign v_5011 = v_89 & v_4721;
assign v_5012 = ~v_91 & v_5011;
assign v_5013 = v_89 & v_4724;
assign v_5014 = ~v_91 & v_5013;
assign v_5016 = v_563 & v_5015;
assign v_5021 = v_4972 & v_5020;
assign v_5022 = v_4975 & v_5021;
assign v_5023 = v_4982 & v_5022;
assign v_5024 = v_4989 & v_5023;
assign v_5033 = v_4972 & v_5032;
assign v_5034 = v_4975 & v_5033;
assign v_5035 = v_4982 & v_5034;
assign v_5036 = v_4989 & v_5035;
assign v_5045 = v_4972 & v_5044;
assign v_5046 = v_4975 & v_5045;
assign v_5047 = v_4982 & v_5046;
assign v_5048 = v_4989 & v_5047;
assign v_5057 = v_4972 & v_5056;
assign v_5058 = v_4975 & v_5057;
assign v_5059 = v_4982 & v_5058;
assign v_5060 = v_4989 & v_5059;
assign v_5069 = v_4972 & v_5068;
assign v_5070 = v_4975 & v_5069;
assign v_5071 = v_4982 & v_5070;
assign v_5072 = v_4989 & v_5071;
assign v_5081 = v_4972 & v_5080;
assign v_5082 = v_4970 & v_5000;
assign v_5084 = v_4975 & v_5083;
assign v_5085 = ~v_91 & v_5002;
assign v_5087 = v_4982 & v_5086;
assign v_5088 = v_4980 & v_5009;
assign v_5090 = v_4989 & v_5089;
assign v_5091 = v_4987 & v_5016;
assign v_5096 = v_5094 & v_5095;
assign v_5099 = v_5097 & v_5098;
assign v_5102 = v_5100 & v_5101;
assign v_5105 = v_5103 & v_5104;
assign v_5109 = v_4972 & v_5108;
assign v_5110 = v_4975 & v_5109;
assign v_5111 = v_4982 & v_5110;
assign v_5112 = v_4989 & v_5111;
assign v_5122 = v_5120 & v_5121;
assign v_5124 = v_5122 & v_5123;
assign v_5127 = v_5125 & v_5126;
assign v_5129 = v_5124 & v_5128;
assign v_5132 = v_5130 & v_5131;
assign v_5134 = v_5129 & v_5133;
assign v_5136 = v_96 & v_4996;
assign v_5138 = v_807 & v_4707;
assign v_5140 = v_91 & v_5004;
assign v_5141 = v_91 & v_5006;
assign v_5143 = v_361 & v_5142;
assign v_5145 = v_91 & v_5011;
assign v_5146 = v_91 & v_5013;
assign v_5148 = v_563 & v_5147;
assign v_5153 = v_5120 & v_5152;
assign v_5154 = v_5123 & v_5153;
assign v_5155 = v_5128 & v_5154;
assign v_5156 = v_5133 & v_5155;
assign v_5165 = v_5120 & v_5164;
assign v_5166 = v_5123 & v_5165;
assign v_5167 = v_5128 & v_5166;
assign v_5168 = v_5133 & v_5167;
assign v_5177 = v_5120 & v_5176;
assign v_5178 = v_5123 & v_5177;
assign v_5179 = v_5128 & v_5178;
assign v_5180 = v_5133 & v_5179;
assign v_5189 = v_5120 & v_5188;
assign v_5190 = v_5123 & v_5189;
assign v_5191 = v_5128 & v_5190;
assign v_5192 = v_5133 & v_5191;
assign v_5201 = v_5120 & v_5200;
assign v_5202 = v_5123 & v_5201;
assign v_5203 = v_5128 & v_5202;
assign v_5204 = v_5133 & v_5203;
assign v_5213 = v_5120 & v_5212;
assign v_5214 = v_91 & v_5136;
assign v_5216 = v_5123 & v_5215;
assign v_5217 = v_4677 & v_5138;
assign v_5219 = v_5128 & v_5218;
assign v_5220 = v_5126 & v_5143;
assign v_5222 = v_5133 & v_5221;
assign v_5223 = v_5131 & v_5148;
assign v_5228 = v_5226 & v_5227;
assign v_5231 = v_5229 & v_5230;
assign v_5234 = v_5232 & v_5233;
assign v_5237 = v_5235 & v_5236;
assign v_5246 = v_5120 & ~v_5240;
assign v_5247 = v_5123 & v_5246;
assign v_5248 = v_5128 & v_5247;
assign v_5249 = v_5133 & v_5248;
assign v_5255 = v_5253 & v_5254;
assign v_5258 = v_5256 & v_5257;
assign v_5260 = v_5258 & v_5259;
assign v_5273 = v_5266 & v_5272;
assign v_5275 = v_5260 & v_5274;
assign v_5288 = v_5281 & v_5287;
assign v_5290 = v_5275 & v_5289;
assign v_5292 = v_89 & v_4995;
assign v_5293 = ~v_91 & v_5292;
assign v_5294 = v_91 & v_4996;
assign v_5296 = v_96 & v_5295;
assign v_5298 = v_807 & v_4704;
assign v_5300 = v_215 & v_616;
assign v_5301 = v_621 & v_5300;
assign v_5302 = v_587 & v_5301;
assign v_5303 = v_87 & v_5302;
assign v_5304 = ~v_89 & v_5303;
assign v_5305 = ~v_91 & v_5304;
assign v_5306 = v_349 & v_646;
assign v_5307 = v_651 & v_5306;
assign v_5308 = v_654 & v_5307;
assign v_5309 = v_87 & v_5308;
assign v_5310 = ~v_89 & v_5309;
assign v_5311 = ~v_91 & v_5310;
assign v_5313 = v_361 & v_5312;
assign v_5315 = v_447 & v_679;
assign v_5316 = v_621 & v_5315;
assign v_5317 = v_587 & v_5316;
assign v_5318 = v_87 & v_5317;
assign v_5319 = ~v_89 & v_5318;
assign v_5320 = ~v_91 & v_5319;
assign v_5321 = v_553 & v_705;
assign v_5322 = v_710 & v_5321;
assign v_5323 = v_654 & v_5322;
assign v_5324 = v_87 & v_5323;
assign v_5325 = ~v_89 & v_5324;
assign v_5326 = ~v_91 & v_5325;
assign v_5328 = v_563 & v_5327;
assign v_5333 = v_5256 & v_5332;
assign v_5334 = v_5259 & v_5333;
assign v_5335 = v_5274 & v_5334;
assign v_5336 = v_5289 & v_5335;
assign v_5345 = v_5256 & v_5344;
assign v_5346 = v_5259 & v_5345;
assign v_5347 = v_5274 & v_5346;
assign v_5348 = v_5289 & v_5347;
assign v_5357 = v_5256 & v_5356;
assign v_5358 = v_5259 & v_5357;
assign v_5359 = v_5274 & v_5358;
assign v_5360 = v_5289 & v_5359;
assign v_5369 = v_5256 & v_5368;
assign v_5370 = v_5259 & v_5369;
assign v_5371 = v_5274 & v_5370;
assign v_5372 = v_5289 & v_5371;
assign v_5381 = v_5256 & v_5380;
assign v_5382 = v_5259 & v_5381;
assign v_5383 = v_5274 & v_5382;
assign v_5384 = v_5289 & v_5383;
assign v_5393 = v_5256 & v_5392;
assign v_5394 = v_5254 & v_5296;
assign v_5396 = v_5259 & v_5395;
assign v_5397 = ~v_91 & v_5298;
assign v_5399 = v_5274 & v_5398;
assign v_5400 = v_5272 & v_5313;
assign v_5402 = v_5289 & v_5401;
assign v_5403 = v_5287 & v_5328;
assign v_5408 = v_5406 & v_5407;
assign v_5411 = v_5409 & v_5410;
assign v_5414 = v_5412 & v_5413;
assign v_5417 = v_5415 & v_5416;
assign v_5426 = v_5256 & ~v_5420;
assign v_5427 = v_5259 & v_5426;
assign v_5428 = v_5274 & v_5427;
assign v_5429 = v_5289 & v_5428;
assign v_5434 = v_5432 & v_5433;
assign v_5436 = v_5434 & v_5435;
assign v_5439 = v_5437 & v_5438;
assign v_5441 = v_5436 & v_5440;
assign v_5444 = v_5442 & v_5443;
assign v_5446 = v_5441 & v_5445;
assign v_5448 = v_96 & v_5292;
assign v_5450 = v_807 & v_4999;
assign v_5452 = v_91 & v_5304;
assign v_5453 = v_91 & v_5310;
assign v_5455 = v_361 & v_5454;
assign v_5457 = v_91 & v_5319;
assign v_5458 = v_91 & v_5325;
assign v_5460 = v_563 & v_5459;
assign v_5465 = v_5432 & v_5464;
assign v_5466 = v_5435 & v_5465;
assign v_5467 = v_5440 & v_5466;
assign v_5468 = v_5445 & v_5467;
assign v_5477 = v_5432 & v_5476;
assign v_5478 = v_5435 & v_5477;
assign v_5479 = v_5440 & v_5478;
assign v_5480 = v_5445 & v_5479;
assign v_5489 = v_5432 & v_5488;
assign v_5490 = v_5435 & v_5489;
assign v_5491 = v_5440 & v_5490;
assign v_5492 = v_5445 & v_5491;
assign v_5501 = v_5432 & v_5500;
assign v_5502 = v_5435 & v_5501;
assign v_5503 = v_5440 & v_5502;
assign v_5504 = v_5445 & v_5503;
assign v_5513 = v_5432 & v_5512;
assign v_5514 = v_5435 & v_5513;
assign v_5515 = v_5440 & v_5514;
assign v_5516 = v_5445 & v_5515;
assign v_5525 = v_5432 & v_5524;
assign v_5526 = v_91 & v_5448;
assign v_5528 = v_5435 & v_5527;
assign v_5529 = v_4969 & v_5450;
assign v_5531 = v_5440 & v_5530;
assign v_5532 = v_5438 & v_5455;
assign v_5534 = v_5445 & v_5533;
assign v_5535 = v_5443 & v_5460;
assign v_5540 = v_5538 & v_5539;
assign v_5543 = v_5541 & v_5542;
assign v_5546 = v_5544 & v_5545;
assign v_5549 = v_5547 & v_5548;
assign v_5553 = v_5432 & v_5552;
assign v_5554 = v_5435 & v_5553;
assign v_5555 = v_5440 & v_5554;
assign v_5556 = v_5445 & v_5555;
assign v_5568 = v_5566 & v_5567;
assign v_5571 = v_5569 & v_5570;
assign v_5573 = v_5571 & v_5572;
assign v_5578 = v_5575 & v_5577;
assign v_5580 = v_5573 & v_5579;
assign v_5585 = v_5582 & v_5584;
assign v_5587 = v_5580 & v_5586;
assign v_5589 = ~v_87 & v_4994;
assign v_5590 = ~v_89 & v_5589;
assign v_5591 = ~v_91 & v_5590;
assign v_5592 = v_91 & v_5292;
assign v_5594 = v_96 & v_5593;
assign v_5596 = v_807 & v_4996;
assign v_5598 = v_89 & v_5303;
assign v_5599 = ~v_91 & v_5598;
assign v_5600 = v_89 & v_5309;
assign v_5601 = ~v_91 & v_5600;
assign v_5603 = v_361 & v_5602;
assign v_5605 = v_89 & v_5318;
assign v_5606 = ~v_91 & v_5605;
assign v_5607 = v_89 & v_5324;
assign v_5608 = ~v_91 & v_5607;
assign v_5610 = v_563 & v_5609;
assign v_5615 = v_5569 & v_5614;
assign v_5616 = v_5572 & v_5615;
assign v_5617 = v_5579 & v_5616;
assign v_5618 = v_5586 & v_5617;
assign v_5627 = v_5569 & v_5626;
assign v_5628 = v_5572 & v_5627;
assign v_5629 = v_5579 & v_5628;
assign v_5630 = v_5586 & v_5629;
assign v_5639 = v_5569 & v_5638;
assign v_5640 = v_5572 & v_5639;
assign v_5641 = v_5579 & v_5640;
assign v_5642 = v_5586 & v_5641;
assign v_5651 = v_5569 & v_5650;
assign v_5652 = v_5572 & v_5651;
assign v_5653 = v_5579 & v_5652;
assign v_5654 = v_5586 & v_5653;
assign v_5663 = v_5569 & v_5662;
assign v_5664 = v_5572 & v_5663;
assign v_5665 = v_5579 & v_5664;
assign v_5666 = v_5586 & v_5665;
assign v_5675 = v_5569 & v_5674;
assign v_5676 = v_5567 & v_5594;
assign v_5678 = v_5572 & v_5677;
assign v_5679 = ~v_91 & v_5596;
assign v_5681 = v_5579 & v_5680;
assign v_5682 = v_5577 & v_5603;
assign v_5684 = v_5586 & v_5683;
assign v_5685 = v_5584 & v_5610;
assign v_5690 = v_5688 & v_5689;
assign v_5693 = v_5691 & v_5692;
assign v_5696 = v_5694 & v_5695;
assign v_5699 = v_5697 & v_5698;
assign v_5703 = v_5569 & v_5702;
assign v_5704 = v_5572 & v_5703;
assign v_5705 = v_5579 & v_5704;
assign v_5706 = v_5586 & v_5705;
assign v_5716 = v_5714 & v_5715;
assign v_5718 = v_5716 & v_5717;
assign v_5721 = v_5719 & v_5720;
assign v_5723 = v_5718 & v_5722;
assign v_5726 = v_5724 & v_5725;
assign v_5728 = v_5723 & v_5727;
assign v_5730 = v_96 & v_5590;
assign v_5732 = v_807 & v_5295;
assign v_5734 = v_91 & v_5598;
assign v_5735 = v_91 & v_5600;
assign v_5737 = v_361 & v_5736;
assign v_5739 = v_91 & v_5605;
assign v_5740 = v_91 & v_5607;
assign v_5742 = v_563 & v_5741;
assign v_5747 = v_5714 & v_5746;
assign v_5748 = v_5717 & v_5747;
assign v_5749 = v_5722 & v_5748;
assign v_5750 = v_5727 & v_5749;
assign v_5759 = v_5714 & v_5758;
assign v_5760 = v_5717 & v_5759;
assign v_5761 = v_5722 & v_5760;
assign v_5762 = v_5727 & v_5761;
assign v_5771 = v_5714 & v_5770;
assign v_5772 = v_5717 & v_5771;
assign v_5773 = v_5722 & v_5772;
assign v_5774 = v_5727 & v_5773;
assign v_5783 = v_5714 & v_5782;
assign v_5784 = v_5717 & v_5783;
assign v_5785 = v_5722 & v_5784;
assign v_5786 = v_5727 & v_5785;
assign v_5795 = v_5714 & v_5794;
assign v_5796 = v_5717 & v_5795;
assign v_5797 = v_5722 & v_5796;
assign v_5798 = v_5727 & v_5797;
assign v_5809 = v_5807 & v_5808;
assign v_5812 = v_5810 & v_5811;
assign v_5815 = v_5813 & v_5814;
assign v_5818 = v_5816 & v_5817;
assign v_5820 = v_5714 & ~v_5806;
assign v_5821 = v_91 & v_5730;
assign v_5823 = v_5717 & v_5822;
assign v_5824 = v_5253 & v_5732;
assign v_5826 = v_5722 & v_5825;
assign v_5827 = v_5720 & v_5737;
assign v_5829 = v_5727 & v_5828;
assign v_5830 = v_5725 & v_5742;
assign v_5835 = v_5714 & v_5834;
assign v_5836 = v_5717 & v_5835;
assign v_5837 = v_5722 & v_5836;
assign v_5838 = v_5727 & v_5837;
assign v_5849 = v_5847 & v_5848;
assign v_5852 = v_5850 & v_5851;
assign v_5854 = v_5852 & v_5853;
assign v_5861 = v_5857 & v_5860;
assign v_5863 = v_5854 & v_5862;
assign v_5870 = v_5866 & v_5869;
assign v_5872 = v_5863 & v_5871;
assign v_5874 = v_89 & v_5589;
assign v_5875 = ~v_91 & v_5874;
assign v_5876 = v_91 & v_5590;
assign v_5878 = v_96 & v_5877;
assign v_5880 = v_807 & v_5292;
assign v_5882 = ~v_87 & v_5302;
assign v_5883 = ~v_89 & v_5882;
assign v_5884 = ~v_91 & v_5883;
assign v_5885 = ~v_87 & v_5308;
assign v_5886 = ~v_89 & v_5885;
assign v_5887 = ~v_91 & v_5886;
assign v_5889 = v_361 & v_5888;
assign v_5891 = ~v_87 & v_5317;
assign v_5892 = ~v_89 & v_5891;
assign v_5893 = ~v_91 & v_5892;
assign v_5894 = ~v_87 & v_5323;
assign v_5895 = ~v_89 & v_5894;
assign v_5896 = ~v_91 & v_5895;
assign v_5898 = v_563 & v_5897;
assign v_5903 = v_5850 & v_5902;
assign v_5904 = v_5853 & v_5903;
assign v_5905 = v_5862 & v_5904;
assign v_5906 = v_5871 & v_5905;
assign v_5915 = v_5850 & v_5914;
assign v_5916 = v_5853 & v_5915;
assign v_5917 = v_5862 & v_5916;
assign v_5918 = v_5871 & v_5917;
assign v_5927 = v_5850 & v_5926;
assign v_5928 = v_5853 & v_5927;
assign v_5929 = v_5862 & v_5928;
assign v_5930 = v_5871 & v_5929;
assign v_5939 = v_5850 & v_5938;
assign v_5940 = v_5853 & v_5939;
assign v_5941 = v_5862 & v_5940;
assign v_5942 = v_5871 & v_5941;
assign v_5951 = v_5850 & v_5950;
assign v_5952 = v_5853 & v_5951;
assign v_5953 = v_5862 & v_5952;
assign v_5954 = v_5871 & v_5953;
assign v_5963 = v_5850 & v_5962;
assign v_5964 = v_5848 & v_5878;
assign v_5966 = v_5853 & v_5965;
assign v_5967 = ~v_91 & v_5880;
assign v_5969 = v_5862 & v_5968;
assign v_5970 = v_5860 & v_5889;
assign v_5972 = v_5871 & v_5971;
assign v_5973 = v_5869 & v_5898;
assign v_5978 = v_5976 & v_5977;
assign v_5981 = v_5979 & v_5980;
assign v_5984 = v_5982 & v_5983;
assign v_5987 = v_5985 & v_5986;
assign v_5991 = v_5850 & v_5990;
assign v_5992 = v_5853 & v_5991;
assign v_5993 = v_5862 & v_5992;
assign v_5994 = v_5871 & v_5993;
assign v_6004 = v_6002 & v_6003;
assign v_6006 = v_6004 & v_6005;
assign v_6009 = v_6007 & v_6008;
assign v_6011 = v_6006 & v_6010;
assign v_6014 = v_6012 & v_6013;
assign v_6016 = v_6011 & v_6015;
assign v_6018 = v_96 & v_5874;
assign v_6020 = v_807 & v_5593;
assign v_6022 = v_91 & v_5883;
assign v_6023 = v_91 & v_5886;
assign v_6025 = v_361 & v_6024;
assign v_6027 = v_91 & v_5892;
assign v_6028 = v_91 & v_5895;
assign v_6030 = v_563 & v_6029;
assign v_6035 = v_6002 & v_6034;
assign v_6036 = v_6005 & v_6035;
assign v_6037 = v_6010 & v_6036;
assign v_6038 = v_6015 & v_6037;
assign v_6047 = v_6002 & v_6046;
assign v_6048 = v_6005 & v_6047;
assign v_6049 = v_6010 & v_6048;
assign v_6050 = v_6015 & v_6049;
assign v_6059 = v_6002 & v_6058;
assign v_6060 = v_6005 & v_6059;
assign v_6061 = v_6010 & v_6060;
assign v_6062 = v_6015 & v_6061;
assign v_6071 = v_6002 & v_6070;
assign v_6072 = v_6005 & v_6071;
assign v_6073 = v_6010 & v_6072;
assign v_6074 = v_6015 & v_6073;
assign v_6083 = v_6002 & v_6082;
assign v_6084 = v_6005 & v_6083;
assign v_6085 = v_6010 & v_6084;
assign v_6086 = v_6015 & v_6085;
assign v_6097 = v_6095 & v_6096;
assign v_6100 = v_6098 & v_6099;
assign v_6103 = v_6101 & v_6102;
assign v_6106 = v_6104 & v_6105;
assign v_6108 = v_6002 & ~v_6094;
assign v_6109 = v_91 & v_6018;
assign v_6111 = v_6005 & v_6110;
assign v_6112 = v_5566 & v_6020;
assign v_6114 = v_6010 & v_6113;
assign v_6115 = v_6008 & v_6025;
assign v_6117 = v_6015 & v_6116;
assign v_6118 = v_6013 & v_6030;
assign v_6123 = v_6002 & v_6122;
assign v_6124 = v_6005 & v_6123;
assign v_6125 = v_6010 & v_6124;
assign v_6126 = v_6015 & v_6125;
assign v_6139 = v_6137 & v_6138;
assign v_6142 = v_6140 & v_6141;
assign v_6144 = v_6142 & v_6143;
assign v_6149 = v_6146 & v_6148;
assign v_6151 = v_6144 & v_6150;
assign v_6156 = v_6153 & v_6155;
assign v_6158 = v_6151 & v_6157;
assign v_6160 = v_85 & v_4993;
assign v_6161 = v_87 & v_6160;
assign v_6162 = ~v_89 & v_6161;
assign v_6163 = ~v_91 & v_6162;
assign v_6164 = v_91 & v_5874;
assign v_6166 = v_96 & v_6165;
assign v_6168 = v_807 & v_5590;
assign v_6170 = v_89 & v_5882;
assign v_6171 = ~v_91 & v_6170;
assign v_6172 = v_89 & v_5885;
assign v_6173 = ~v_91 & v_6172;
assign v_6175 = v_361 & v_6174;
assign v_6177 = v_89 & v_5891;
assign v_6178 = ~v_91 & v_6177;
assign v_6179 = v_89 & v_5894;
assign v_6180 = ~v_91 & v_6179;
assign v_6182 = v_563 & v_6181;
assign v_6187 = v_6140 & v_6186;
assign v_6188 = v_6143 & v_6187;
assign v_6189 = v_6150 & v_6188;
assign v_6190 = v_6157 & v_6189;
assign v_6199 = v_6140 & v_6198;
assign v_6200 = v_6143 & v_6199;
assign v_6201 = v_6150 & v_6200;
assign v_6202 = v_6157 & v_6201;
assign v_6211 = v_6140 & v_6210;
assign v_6212 = v_6143 & v_6211;
assign v_6213 = v_6150 & v_6212;
assign v_6214 = v_6157 & v_6213;
assign v_6223 = v_6140 & v_6222;
assign v_6224 = v_6143 & v_6223;
assign v_6225 = v_6150 & v_6224;
assign v_6226 = v_6157 & v_6225;
assign v_6235 = v_6140 & v_6234;
assign v_6236 = v_6143 & v_6235;
assign v_6237 = v_6150 & v_6236;
assign v_6238 = v_6157 & v_6237;
assign v_6247 = v_6140 & v_6246;
assign v_6248 = v_6138 & v_6166;
assign v_6250 = v_6143 & v_6249;
assign v_6251 = ~v_91 & v_6168;
assign v_6253 = v_6150 & v_6252;
assign v_6254 = v_6148 & v_6175;
assign v_6256 = v_6157 & v_6255;
assign v_6257 = v_6155 & v_6182;
assign v_6262 = v_6260 & v_6261;
assign v_6265 = v_6263 & v_6264;
assign v_6268 = v_6266 & v_6267;
assign v_6271 = v_6269 & v_6270;
assign v_6275 = v_6140 & v_6274;
assign v_6276 = v_6143 & v_6275;
assign v_6277 = v_6150 & v_6276;
assign v_6278 = v_6157 & v_6277;
assign v_6288 = v_6286 & v_6287;
assign v_6290 = v_6288 & v_6289;
assign v_6293 = v_6291 & v_6292;
assign v_6295 = v_6290 & v_6294;
assign v_6298 = v_6296 & v_6297;
assign v_6300 = v_6295 & v_6299;
assign v_6302 = v_96 & v_6162;
assign v_6304 = v_807 & v_5877;
assign v_6306 = v_91 & v_6170;
assign v_6307 = v_91 & v_6172;
assign v_6309 = v_361 & v_6308;
assign v_6311 = v_91 & v_6177;
assign v_6312 = v_91 & v_6179;
assign v_6314 = v_563 & v_6313;
assign v_6319 = v_6286 & v_6318;
assign v_6320 = v_6289 & v_6319;
assign v_6321 = v_6294 & v_6320;
assign v_6322 = v_6299 & v_6321;
assign v_6331 = v_6286 & v_6330;
assign v_6332 = v_6289 & v_6331;
assign v_6333 = v_6294 & v_6332;
assign v_6334 = v_6299 & v_6333;
assign v_6343 = v_6286 & v_6342;
assign v_6344 = v_6289 & v_6343;
assign v_6345 = v_6294 & v_6344;
assign v_6346 = v_6299 & v_6345;
assign v_6355 = v_6286 & v_6354;
assign v_6356 = v_6289 & v_6355;
assign v_6357 = v_6294 & v_6356;
assign v_6358 = v_6299 & v_6357;
assign v_6367 = v_6286 & v_6366;
assign v_6368 = v_6289 & v_6367;
assign v_6369 = v_6294 & v_6368;
assign v_6370 = v_6299 & v_6369;
assign v_6379 = v_6286 & v_6378;
assign v_6380 = v_91 & v_6302;
assign v_6382 = v_6289 & v_6381;
assign v_6383 = v_5847 & v_6304;
assign v_6385 = v_6294 & v_6384;
assign v_6386 = v_6292 & v_6309;
assign v_6388 = v_6299 & v_6387;
assign v_6389 = v_6297 & v_6314;
assign v_6394 = v_6392 & v_6393;
assign v_6397 = v_6395 & v_6396;
assign v_6400 = v_6398 & v_6399;
assign v_6403 = v_6401 & v_6402;
assign v_6412 = v_6286 & ~v_6406;
assign v_6413 = v_6289 & v_6412;
assign v_6414 = v_6294 & v_6413;
assign v_6415 = v_6299 & v_6414;
assign v_6421 = v_6419 & v_6420;
assign v_6424 = v_6422 & v_6423;
assign v_6426 = v_6424 & v_6425;
assign v_6435 = v_6430 & v_6434;
assign v_6437 = v_6426 & v_6436;
assign v_6446 = v_6441 & v_6445;
assign v_6448 = v_6437 & v_6447;
assign v_6450 = v_89 & v_6161;
assign v_6451 = ~v_91 & v_6450;
assign v_6452 = v_91 & v_6162;
assign v_6454 = v_96 & v_6453;
assign v_6456 = v_807 & v_5874;
assign v_6458 = v_85 & v_5301;
assign v_6459 = v_87 & v_6458;
assign v_6460 = ~v_89 & v_6459;
assign v_6461 = ~v_91 & v_6460;
assign v_6462 = v_355 & v_5307;
assign v_6463 = v_87 & v_6462;
assign v_6464 = ~v_89 & v_6463;
assign v_6465 = ~v_91 & v_6464;
assign v_6467 = v_361 & v_6466;
assign v_6469 = v_85 & v_5316;
assign v_6470 = v_87 & v_6469;
assign v_6471 = ~v_89 & v_6470;
assign v_6472 = ~v_91 & v_6471;
assign v_6473 = v_355 & v_5322;
assign v_6474 = v_87 & v_6473;
assign v_6475 = ~v_89 & v_6474;
assign v_6476 = ~v_91 & v_6475;
assign v_6478 = v_563 & v_6477;
assign v_6483 = v_6422 & v_6482;
assign v_6484 = v_6425 & v_6483;
assign v_6485 = v_6436 & v_6484;
assign v_6486 = v_6447 & v_6485;
assign v_6495 = v_6422 & v_6494;
assign v_6496 = v_6425 & v_6495;
assign v_6497 = v_6436 & v_6496;
assign v_6498 = v_6447 & v_6497;
assign v_6507 = v_6422 & v_6506;
assign v_6508 = v_6425 & v_6507;
assign v_6509 = v_6436 & v_6508;
assign v_6510 = v_6447 & v_6509;
assign v_6519 = v_6422 & v_6518;
assign v_6520 = v_6425 & v_6519;
assign v_6521 = v_6436 & v_6520;
assign v_6522 = v_6447 & v_6521;
assign v_6531 = v_6422 & v_6530;
assign v_6532 = v_6425 & v_6531;
assign v_6533 = v_6436 & v_6532;
assign v_6534 = v_6447 & v_6533;
assign v_6543 = v_6422 & v_6542;
assign v_6544 = v_6420 & v_6454;
assign v_6546 = v_6425 & v_6545;
assign v_6547 = ~v_91 & v_6456;
assign v_6549 = v_6436 & v_6548;
assign v_6550 = v_6434 & v_6467;
assign v_6552 = v_6447 & v_6551;
assign v_6553 = v_6445 & v_6478;
assign v_6558 = v_6556 & v_6557;
assign v_6561 = v_6559 & v_6560;
assign v_6564 = v_6562 & v_6563;
assign v_6567 = v_6565 & v_6566;
assign v_6576 = v_6422 & ~v_6570;
assign v_6577 = v_6425 & v_6576;
assign v_6578 = v_6436 & v_6577;
assign v_6579 = v_6447 & v_6578;
assign v_6584 = v_6582 & v_6583;
assign v_6586 = v_6584 & v_6585;
assign v_6589 = v_6587 & v_6588;
assign v_6591 = v_6586 & v_6590;
assign v_6594 = v_6592 & v_6593;
assign v_6596 = v_6591 & v_6595;
assign v_6598 = v_96 & v_6450;
assign v_6600 = v_807 & v_6165;
assign v_6602 = v_91 & v_6460;
assign v_6603 = v_91 & v_6464;
assign v_6605 = v_361 & v_6604;
assign v_6607 = v_91 & v_6471;
assign v_6608 = v_91 & v_6475;
assign v_6610 = v_563 & v_6609;
assign v_6615 = v_6582 & v_6614;
assign v_6616 = v_6585 & v_6615;
assign v_6617 = v_6590 & v_6616;
assign v_6618 = v_6595 & v_6617;
assign v_6627 = v_6582 & v_6626;
assign v_6628 = v_6585 & v_6627;
assign v_6629 = v_6590 & v_6628;
assign v_6630 = v_6595 & v_6629;
assign v_6639 = v_6582 & v_6638;
assign v_6640 = v_6585 & v_6639;
assign v_6641 = v_6590 & v_6640;
assign v_6642 = v_6595 & v_6641;
assign v_6651 = v_6582 & v_6650;
assign v_6652 = v_6585 & v_6651;
assign v_6653 = v_6590 & v_6652;
assign v_6654 = v_6595 & v_6653;
assign v_6663 = v_6582 & v_6662;
assign v_6664 = v_6585 & v_6663;
assign v_6665 = v_6590 & v_6664;
assign v_6666 = v_6595 & v_6665;
assign v_6675 = v_6582 & v_6674;
assign v_6676 = v_91 & v_6598;
assign v_6678 = v_6585 & v_6677;
assign v_6679 = v_6137 & v_6600;
assign v_6681 = v_6590 & v_6680;
assign v_6682 = v_6588 & v_6605;
assign v_6684 = v_6595 & v_6683;
assign v_6685 = v_6593 & v_6610;
assign v_6690 = v_6688 & v_6689;
assign v_6693 = v_6691 & v_6692;
assign v_6696 = v_6694 & v_6695;
assign v_6699 = v_6697 & v_6698;
assign v_6703 = v_6582 & v_6702;
assign v_6704 = v_6585 & v_6703;
assign v_6705 = v_6590 & v_6704;
assign v_6706 = v_6595 & v_6705;
assign v_6718 = v_6716 & v_6717;
assign v_6721 = v_6719 & v_6720;
assign v_6723 = v_6721 & v_6722;
assign v_6728 = v_6725 & v_6727;
assign v_6730 = v_6723 & v_6729;
assign v_6735 = v_6732 & v_6734;
assign v_6737 = v_6730 & v_6736;
assign v_6739 = ~v_87 & v_6160;
assign v_6740 = ~v_89 & v_6739;
assign v_6741 = ~v_91 & v_6740;
assign v_6742 = v_91 & v_6450;
assign v_6744 = v_96 & v_6743;
assign v_6746 = v_807 & v_6162;
assign v_6748 = v_89 & v_6459;
assign v_6749 = ~v_91 & v_6748;
assign v_6750 = v_89 & v_6463;
assign v_6751 = ~v_91 & v_6750;
assign v_6753 = v_361 & v_6752;
assign v_6755 = v_89 & v_6470;
assign v_6756 = ~v_91 & v_6755;
assign v_6757 = v_89 & v_6474;
assign v_6758 = ~v_91 & v_6757;
assign v_6760 = v_563 & v_6759;
assign v_6765 = v_6719 & v_6764;
assign v_6766 = v_6722 & v_6765;
assign v_6767 = v_6729 & v_6766;
assign v_6768 = v_6736 & v_6767;
assign v_6777 = v_6719 & v_6776;
assign v_6778 = v_6722 & v_6777;
assign v_6779 = v_6729 & v_6778;
assign v_6780 = v_6736 & v_6779;
assign v_6789 = v_6719 & v_6788;
assign v_6790 = v_6722 & v_6789;
assign v_6791 = v_6729 & v_6790;
assign v_6792 = v_6736 & v_6791;
assign v_6801 = v_6719 & v_6800;
assign v_6802 = v_6722 & v_6801;
assign v_6803 = v_6729 & v_6802;
assign v_6804 = v_6736 & v_6803;
assign v_6813 = v_6719 & v_6812;
assign v_6814 = v_6722 & v_6813;
assign v_6815 = v_6729 & v_6814;
assign v_6816 = v_6736 & v_6815;
assign v_6827 = v_6825 & v_6826;
assign v_6830 = v_6828 & v_6829;
assign v_6833 = v_6831 & v_6832;
assign v_6836 = v_6834 & v_6835;
assign v_6838 = v_6719 & ~v_6824;
assign v_6839 = v_6717 & v_6744;
assign v_6841 = v_6722 & v_6840;
assign v_6842 = ~v_91 & v_6746;
assign v_6844 = v_6729 & v_6843;
assign v_6845 = v_6727 & v_6753;
assign v_6847 = v_6736 & v_6846;
assign v_6848 = v_6734 & v_6760;
assign v_6853 = v_6719 & v_6852;
assign v_6854 = v_6722 & v_6853;
assign v_6855 = v_6729 & v_6854;
assign v_6856 = v_6736 & v_6855;
assign v_6866 = v_6864 & v_6865;
assign v_6868 = v_6866 & v_6867;
assign v_6871 = v_6869 & v_6870;
assign v_6873 = v_6868 & v_6872;
assign v_6876 = v_6874 & v_6875;
assign v_6878 = v_6873 & v_6877;
assign v_6880 = v_96 & v_6740;
assign v_6882 = v_807 & v_6453;
assign v_6884 = v_91 & v_6748;
assign v_6885 = v_91 & v_6750;
assign v_6887 = v_361 & v_6886;
assign v_6889 = v_91 & v_6755;
assign v_6890 = v_91 & v_6757;
assign v_6892 = v_563 & v_6891;
assign v_6897 = v_6864 & v_6896;
assign v_6898 = v_6867 & v_6897;
assign v_6899 = v_6872 & v_6898;
assign v_6900 = v_6877 & v_6899;
assign v_6909 = v_6864 & v_6908;
assign v_6910 = v_6867 & v_6909;
assign v_6911 = v_6872 & v_6910;
assign v_6912 = v_6877 & v_6911;
assign v_6921 = v_6864 & v_6920;
assign v_6922 = v_6867 & v_6921;
assign v_6923 = v_6872 & v_6922;
assign v_6924 = v_6877 & v_6923;
assign v_6933 = v_6864 & v_6932;
assign v_6934 = v_6867 & v_6933;
assign v_6935 = v_6872 & v_6934;
assign v_6936 = v_6877 & v_6935;
assign v_6945 = v_6864 & v_6944;
assign v_6946 = v_6867 & v_6945;
assign v_6947 = v_6872 & v_6946;
assign v_6948 = v_6877 & v_6947;
assign v_6957 = v_6864 & v_6956;
assign v_6958 = v_91 & v_6880;
assign v_6960 = v_6867 & v_6959;
assign v_6961 = v_6419 & v_6882;
assign v_6963 = v_6872 & v_6962;
assign v_6964 = v_6870 & v_6887;
assign v_6966 = v_6877 & v_6965;
assign v_6967 = v_6875 & v_6892;
assign v_6972 = v_6970 & v_6971;
assign v_6975 = v_6973 & v_6974;
assign v_6978 = v_6976 & v_6977;
assign v_6981 = v_6979 & v_6980;
assign v_6985 = v_6864 & v_6984;
assign v_6986 = v_6867 & v_6985;
assign v_6987 = v_6872 & v_6986;
assign v_6988 = v_6877 & v_6987;
assign v_6999 = v_6997 & v_6998;
assign v_7002 = v_7000 & v_7001;
assign v_7004 = v_7002 & v_7003;
assign v_7011 = v_7007 & v_7010;
assign v_7013 = v_7004 & v_7012;
assign v_7020 = v_7016 & v_7019;
assign v_7022 = v_7013 & v_7021;
assign v_7024 = v_89 & v_6739;
assign v_7025 = ~v_91 & v_7024;
assign v_7026 = v_91 & v_6740;
assign v_7028 = v_96 & v_7027;
assign v_7030 = v_807 & v_6450;
assign v_7032 = ~v_87 & v_6458;
assign v_7033 = ~v_89 & v_7032;
assign v_7034 = ~v_91 & v_7033;
assign v_7035 = ~v_87 & v_6462;
assign v_7036 = ~v_89 & v_7035;
assign v_7037 = ~v_91 & v_7036;
assign v_7039 = v_361 & v_7038;
assign v_7041 = ~v_87 & v_6469;
assign v_7042 = ~v_89 & v_7041;
assign v_7043 = ~v_91 & v_7042;
assign v_7044 = ~v_87 & v_6473;
assign v_7045 = ~v_89 & v_7044;
assign v_7046 = ~v_91 & v_7045;
assign v_7048 = v_563 & v_7047;
assign v_7053 = v_7000 & v_7052;
assign v_7054 = v_7003 & v_7053;
assign v_7055 = v_7012 & v_7054;
assign v_7056 = v_7021 & v_7055;
assign v_7065 = v_7000 & v_7064;
assign v_7066 = v_7003 & v_7065;
assign v_7067 = v_7012 & v_7066;
assign v_7068 = v_7021 & v_7067;
assign v_7077 = v_7000 & v_7076;
assign v_7078 = v_7003 & v_7077;
assign v_7079 = v_7012 & v_7078;
assign v_7080 = v_7021 & v_7079;
assign v_7089 = v_7000 & v_7088;
assign v_7090 = v_7003 & v_7089;
assign v_7091 = v_7012 & v_7090;
assign v_7092 = v_7021 & v_7091;
assign v_7101 = v_7000 & v_7100;
assign v_7102 = v_7003 & v_7101;
assign v_7103 = v_7012 & v_7102;
assign v_7104 = v_7021 & v_7103;
assign v_7113 = v_7000 & v_7112;
assign v_7114 = v_6998 & v_7028;
assign v_7116 = v_7003 & v_7115;
assign v_7117 = ~v_91 & v_7030;
assign v_7119 = v_7012 & v_7118;
assign v_7120 = v_7010 & v_7039;
assign v_7122 = v_7021 & v_7121;
assign v_7123 = v_7019 & v_7048;
assign v_7128 = v_7126 & v_7127;
assign v_7131 = v_7129 & v_7130;
assign v_7134 = v_7132 & v_7133;
assign v_7137 = v_7135 & v_7136;
assign v_7146 = v_7000 & ~v_7140;
assign v_7147 = v_7003 & v_7146;
assign v_7148 = v_7012 & v_7147;
assign v_7149 = v_7021 & v_7148;
assign v_7154 = v_7152 & v_7153;
assign v_7156 = v_7154 & v_7155;
assign v_7159 = v_7157 & v_7158;
assign v_7161 = v_7156 & v_7160;
assign v_7164 = v_7162 & v_7163;
assign v_7166 = v_7161 & v_7165;
assign v_7168 = v_96 & v_7024;
assign v_7170 = v_807 & v_6743;
assign v_7172 = v_91 & v_7033;
assign v_7173 = v_91 & v_7036;
assign v_7175 = v_361 & v_7174;
assign v_7177 = v_91 & v_7042;
assign v_7178 = v_91 & v_7045;
assign v_7180 = v_563 & v_7179;
assign v_7185 = v_7152 & v_7184;
assign v_7186 = v_7155 & v_7185;
assign v_7187 = v_7160 & v_7186;
assign v_7188 = v_7165 & v_7187;
assign v_7197 = v_7152 & v_7196;
assign v_7198 = v_7155 & v_7197;
assign v_7199 = v_7160 & v_7198;
assign v_7200 = v_7165 & v_7199;
assign v_7209 = v_7152 & v_7208;
assign v_7210 = v_7155 & v_7209;
assign v_7211 = v_7160 & v_7210;
assign v_7212 = v_7165 & v_7211;
assign v_7221 = v_7152 & v_7220;
assign v_7222 = v_7155 & v_7221;
assign v_7223 = v_7160 & v_7222;
assign v_7224 = v_7165 & v_7223;
assign v_7233 = v_7152 & v_7232;
assign v_7234 = v_7155 & v_7233;
assign v_7235 = v_7160 & v_7234;
assign v_7236 = v_7165 & v_7235;
assign v_7245 = v_7152 & v_7244;
assign v_7246 = v_91 & v_7168;
assign v_7248 = v_7155 & v_7247;
assign v_7249 = v_6716 & v_7170;
assign v_7251 = v_7160 & v_7250;
assign v_7252 = v_7158 & v_7175;
assign v_7254 = v_7165 & v_7253;
assign v_7255 = v_7163 & v_7180;
assign v_7260 = v_7258 & v_7259;
assign v_7263 = v_7261 & v_7262;
assign v_7266 = v_7264 & v_7265;
assign v_7269 = v_7267 & v_7268;
assign v_7273 = v_7152 & v_7272;
assign v_7274 = v_7155 & v_7273;
assign v_7275 = v_7160 & v_7274;
assign v_7276 = v_7165 & v_7275;
assign v_7290 = v_7288 & v_7289;
assign v_7293 = v_7291 & v_7292;
assign v_7295 = v_7293 & v_7294;
assign v_7300 = v_7297 & v_7299;
assign v_7302 = v_7295 & v_7301;
assign v_7307 = v_7304 & v_7306;
assign v_7309 = v_7302 & v_7308;
assign v_7311 = v_82 & v_4992;
assign v_7312 = v_587 & v_7311;
assign v_7313 = v_87 & v_7312;
assign v_7314 = ~v_89 & v_7313;
assign v_7315 = ~v_91 & v_7314;
assign v_7316 = v_91 & v_7024;
assign v_7318 = v_96 & v_7317;
assign v_7320 = v_807 & v_6740;
assign v_7322 = v_89 & v_7032;
assign v_7323 = ~v_91 & v_7322;
assign v_7324 = v_89 & v_7035;
assign v_7325 = ~v_91 & v_7324;
assign v_7327 = v_361 & v_7326;
assign v_7329 = v_89 & v_7041;
assign v_7330 = ~v_91 & v_7329;
assign v_7331 = v_89 & v_7044;
assign v_7332 = ~v_91 & v_7331;
assign v_7334 = v_563 & v_7333;
assign v_7339 = v_7291 & v_7338;
assign v_7340 = v_7294 & v_7339;
assign v_7341 = v_7301 & v_7340;
assign v_7342 = v_7308 & v_7341;
assign v_7351 = v_7291 & v_7350;
assign v_7352 = v_7294 & v_7351;
assign v_7353 = v_7301 & v_7352;
assign v_7354 = v_7308 & v_7353;
assign v_7363 = v_7291 & v_7362;
assign v_7364 = v_7294 & v_7363;
assign v_7365 = v_7301 & v_7364;
assign v_7366 = v_7308 & v_7365;
assign v_7375 = v_7291 & v_7374;
assign v_7376 = v_7294 & v_7375;
assign v_7377 = v_7301 & v_7376;
assign v_7378 = v_7308 & v_7377;
assign v_7387 = v_7291 & v_7386;
assign v_7388 = v_7294 & v_7387;
assign v_7389 = v_7301 & v_7388;
assign v_7390 = v_7308 & v_7389;
assign v_7399 = v_7291 & v_7398;
assign v_7400 = v_7289 & v_7318;
assign v_7402 = v_7294 & v_7401;
assign v_7403 = ~v_91 & v_7320;
assign v_7405 = v_7301 & v_7404;
assign v_7406 = v_7299 & v_7327;
assign v_7408 = v_7308 & v_7407;
assign v_7409 = v_7306 & v_7334;
assign v_7414 = v_7412 & v_7413;
assign v_7417 = v_7415 & v_7416;
assign v_7420 = v_7418 & v_7419;
assign v_7423 = v_7421 & v_7422;
assign v_7432 = v_7291 & ~v_7426;
assign v_7433 = v_7294 & v_7432;
assign v_7434 = v_7301 & v_7433;
assign v_7435 = v_7308 & v_7434;
assign v_7440 = v_7438 & v_7439;
assign v_7442 = v_7440 & v_7441;
assign v_7445 = v_7443 & v_7444;
assign v_7447 = v_7442 & v_7446;
assign v_7450 = v_7448 & v_7449;
assign v_7452 = v_7447 & v_7451;
assign v_7454 = v_96 & v_7314;
assign v_7456 = v_807 & v_7027;
assign v_7458 = v_91 & v_7322;
assign v_7459 = v_91 & v_7324;
assign v_7461 = v_361 & v_7460;
assign v_7463 = v_91 & v_7329;
assign v_7464 = v_91 & v_7331;
assign v_7466 = v_563 & v_7465;
assign v_7471 = v_7438 & v_7470;
assign v_7472 = v_7441 & v_7471;
assign v_7473 = v_7446 & v_7472;
assign v_7474 = v_7451 & v_7473;
assign v_7483 = v_7438 & v_7482;
assign v_7484 = v_7441 & v_7483;
assign v_7485 = v_7446 & v_7484;
assign v_7486 = v_7451 & v_7485;
assign v_7495 = v_7438 & v_7494;
assign v_7496 = v_7441 & v_7495;
assign v_7497 = v_7446 & v_7496;
assign v_7498 = v_7451 & v_7497;
assign v_7507 = v_7438 & v_7506;
assign v_7508 = v_7441 & v_7507;
assign v_7509 = v_7446 & v_7508;
assign v_7510 = v_7451 & v_7509;
assign v_7519 = v_7438 & v_7518;
assign v_7520 = v_7441 & v_7519;
assign v_7521 = v_7446 & v_7520;
assign v_7522 = v_7451 & v_7521;
assign v_7531 = v_7438 & v_7530;
assign v_7532 = v_91 & v_7454;
assign v_7534 = v_7441 & v_7533;
assign v_7535 = v_6997 & v_7456;
assign v_7537 = v_7446 & v_7536;
assign v_7538 = v_7444 & v_7461;
assign v_7540 = v_7451 & v_7539;
assign v_7541 = v_7449 & v_7466;
assign v_7546 = v_7544 & v_7545;
assign v_7549 = v_7547 & v_7548;
assign v_7552 = v_7550 & v_7551;
assign v_7555 = v_7553 & v_7554;
assign v_7564 = v_7438 & ~v_7558;
assign v_7565 = v_7441 & v_7564;
assign v_7566 = v_7446 & v_7565;
assign v_7567 = v_7451 & v_7566;
assign v_7573 = v_7571 & v_7572;
assign v_7576 = v_7574 & v_7575;
assign v_7578 = v_7576 & v_7577;
assign v_7589 = v_7583 & v_7588;
assign v_7591 = v_7578 & v_7590;
assign v_7602 = v_7596 & v_7601;
assign v_7604 = v_7591 & v_7603;
assign v_7606 = v_89 & v_7313;
assign v_7607 = ~v_91 & v_7606;
assign v_7608 = v_91 & v_7314;
assign v_7610 = v_96 & v_7609;
assign v_7612 = v_807 & v_7024;
assign v_7614 = v_218 & v_5300;
assign v_7615 = v_587 & v_7614;
assign v_7616 = v_87 & v_7615;
assign v_7617 = ~v_89 & v_7616;
assign v_7618 = ~v_91 & v_7617;
assign v_7619 = v_352 & v_5306;
assign v_7620 = v_654 & v_7619;
assign v_7621 = v_87 & v_7620;
assign v_7622 = ~v_89 & v_7621;
assign v_7623 = ~v_91 & v_7622;
assign v_7625 = v_361 & v_7624;
assign v_7627 = v_218 & v_5315;
assign v_7628 = v_587 & v_7627;
assign v_7629 = v_87 & v_7628;
assign v_7630 = ~v_89 & v_7629;
assign v_7631 = ~v_91 & v_7630;
assign v_7632 = v_556 & v_5321;
assign v_7633 = v_654 & v_7632;
assign v_7634 = v_87 & v_7633;
assign v_7635 = ~v_89 & v_7634;
assign v_7636 = ~v_91 & v_7635;
assign v_7638 = v_563 & v_7637;
assign v_7643 = v_7574 & v_7642;
assign v_7644 = v_7577 & v_7643;
assign v_7645 = v_7590 & v_7644;
assign v_7646 = v_7603 & v_7645;
assign v_7655 = v_7574 & v_7654;
assign v_7656 = v_7577 & v_7655;
assign v_7657 = v_7590 & v_7656;
assign v_7658 = v_7603 & v_7657;
assign v_7667 = v_7574 & v_7666;
assign v_7668 = v_7577 & v_7667;
assign v_7669 = v_7590 & v_7668;
assign v_7670 = v_7603 & v_7669;
assign v_7679 = v_7574 & v_7678;
assign v_7680 = v_7577 & v_7679;
assign v_7681 = v_7590 & v_7680;
assign v_7682 = v_7603 & v_7681;
assign v_7691 = v_7574 & v_7690;
assign v_7692 = v_7577 & v_7691;
assign v_7693 = v_7590 & v_7692;
assign v_7694 = v_7603 & v_7693;
assign v_7703 = v_7574 & v_7702;
assign v_7704 = v_7572 & v_7610;
assign v_7706 = v_7577 & v_7705;
assign v_7707 = ~v_91 & v_7612;
assign v_7709 = v_7590 & v_7708;
assign v_7710 = v_7588 & v_7625;
assign v_7712 = v_7603 & v_7711;
assign v_7713 = v_7601 & v_7638;
assign v_7718 = v_7716 & v_7717;
assign v_7721 = v_7719 & v_7720;
assign v_7724 = v_7722 & v_7723;
assign v_7727 = v_7725 & v_7726;
assign v_7736 = v_7574 & ~v_7730;
assign v_7737 = v_7577 & v_7736;
assign v_7738 = v_7590 & v_7737;
assign v_7739 = v_7603 & v_7738;
assign v_7744 = v_7742 & v_7743;
assign v_7746 = v_7744 & v_7745;
assign v_7749 = v_7747 & v_7748;
assign v_7751 = v_7746 & v_7750;
assign v_7754 = v_7752 & v_7753;
assign v_7756 = v_7751 & v_7755;
assign v_7758 = v_96 & v_7606;
assign v_7760 = v_807 & v_7317;
assign v_7762 = v_91 & v_7617;
assign v_7763 = v_91 & v_7622;
assign v_7765 = v_361 & v_7764;
assign v_7767 = v_91 & v_7630;
assign v_7768 = v_91 & v_7635;
assign v_7770 = v_563 & v_7769;
assign v_7775 = v_7742 & v_7774;
assign v_7776 = v_7745 & v_7775;
assign v_7777 = v_7750 & v_7776;
assign v_7778 = v_7755 & v_7777;
assign v_7787 = v_7742 & v_7786;
assign v_7788 = v_7745 & v_7787;
assign v_7789 = v_7750 & v_7788;
assign v_7790 = v_7755 & v_7789;
assign v_7799 = v_7742 & v_7798;
assign v_7800 = v_7745 & v_7799;
assign v_7801 = v_7750 & v_7800;
assign v_7802 = v_7755 & v_7801;
assign v_7811 = v_7742 & v_7810;
assign v_7812 = v_7745 & v_7811;
assign v_7813 = v_7750 & v_7812;
assign v_7814 = v_7755 & v_7813;
assign v_7823 = v_7742 & v_7822;
assign v_7824 = v_7745 & v_7823;
assign v_7825 = v_7750 & v_7824;
assign v_7826 = v_7755 & v_7825;
assign v_7835 = v_7742 & v_7834;
assign v_7836 = v_91 & v_7758;
assign v_7838 = v_7745 & v_7837;
assign v_7839 = v_7288 & v_7760;
assign v_7841 = v_7750 & v_7840;
assign v_7842 = v_7748 & v_7765;
assign v_7844 = v_7755 & v_7843;
assign v_7845 = v_7753 & v_7770;
assign v_7850 = v_7848 & v_7849;
assign v_7853 = v_7851 & v_7852;
assign v_7856 = v_7854 & v_7855;
assign v_7859 = v_7857 & v_7858;
assign v_7868 = v_7742 & ~v_7862;
assign v_7869 = v_7745 & v_7868;
assign v_7870 = v_7750 & v_7869;
assign v_7871 = v_7755 & v_7870;
assign v_7878 = v_7876 & v_7877;
assign v_7881 = v_7879 & v_7880;
assign v_7883 = v_7881 & v_7882;
assign v_7888 = v_7885 & v_7887;
assign v_7890 = v_7883 & v_7889;
assign v_7895 = v_7892 & v_7894;
assign v_7897 = v_7890 & v_7896;
assign v_7899 = ~v_87 & v_7312;
assign v_7900 = ~v_89 & v_7899;
assign v_7901 = ~v_91 & v_7900;
assign v_7902 = v_91 & v_7606;
assign v_7904 = v_96 & v_7903;
assign v_7906 = v_807 & v_7314;
assign v_7908 = v_89 & v_7616;
assign v_7909 = ~v_91 & v_7908;
assign v_7910 = v_89 & v_7621;
assign v_7911 = ~v_91 & v_7910;
assign v_7913 = v_361 & v_7912;
assign v_7915 = v_89 & v_7629;
assign v_7916 = ~v_91 & v_7915;
assign v_7917 = v_89 & v_7634;
assign v_7918 = ~v_91 & v_7917;
assign v_7920 = v_563 & v_7919;
assign v_7925 = v_7879 & v_7924;
assign v_7926 = v_7882 & v_7925;
assign v_7927 = v_7889 & v_7926;
assign v_7928 = v_7896 & v_7927;
assign v_7937 = v_7879 & v_7936;
assign v_7938 = v_7882 & v_7937;
assign v_7939 = v_7889 & v_7938;
assign v_7940 = v_7896 & v_7939;
assign v_7949 = v_7879 & v_7948;
assign v_7950 = v_7882 & v_7949;
assign v_7951 = v_7889 & v_7950;
assign v_7952 = v_7896 & v_7951;
assign v_7961 = v_7879 & v_7960;
assign v_7962 = v_7882 & v_7961;
assign v_7963 = v_7889 & v_7962;
assign v_7964 = v_7896 & v_7963;
assign v_7973 = v_7879 & v_7972;
assign v_7974 = v_7882 & v_7973;
assign v_7975 = v_7889 & v_7974;
assign v_7976 = v_7896 & v_7975;
assign v_7985 = v_7879 & v_7984;
assign v_7986 = v_7877 & v_7904;
assign v_7988 = v_7882 & v_7987;
assign v_7989 = ~v_91 & v_7906;
assign v_7991 = v_7889 & v_7990;
assign v_7992 = v_7887 & v_7913;
assign v_7994 = v_7896 & v_7993;
assign v_7995 = v_7894 & v_7920;
assign v_8000 = v_7998 & v_7999;
assign v_8003 = v_8001 & v_8002;
assign v_8006 = v_8004 & v_8005;
assign v_8009 = v_8007 & v_8008;
assign v_8018 = v_7879 & ~v_8012;
assign v_8019 = v_7882 & v_8018;
assign v_8020 = v_7889 & v_8019;
assign v_8021 = v_7896 & v_8020;
assign v_8026 = v_8024 & v_8025;
assign v_8028 = v_8026 & v_8027;
assign v_8031 = v_8029 & v_8030;
assign v_8033 = v_8028 & v_8032;
assign v_8036 = v_8034 & v_8035;
assign v_8038 = v_8033 & v_8037;
assign v_8040 = v_96 & v_7900;
assign v_8042 = v_807 & v_7609;
assign v_8044 = v_91 & v_7908;
assign v_8045 = v_91 & v_7910;
assign v_8047 = v_361 & v_8046;
assign v_8049 = v_91 & v_7915;
assign v_8050 = v_91 & v_7917;
assign v_8052 = v_563 & v_8051;
assign v_8057 = v_8024 & v_8056;
assign v_8058 = v_8027 & v_8057;
assign v_8059 = v_8032 & v_8058;
assign v_8060 = v_8037 & v_8059;
assign v_8069 = v_8024 & v_8068;
assign v_8070 = v_8027 & v_8069;
assign v_8071 = v_8032 & v_8070;
assign v_8072 = v_8037 & v_8071;
assign v_8081 = v_8024 & v_8080;
assign v_8082 = v_8027 & v_8081;
assign v_8083 = v_8032 & v_8082;
assign v_8084 = v_8037 & v_8083;
assign v_8093 = v_8024 & v_8092;
assign v_8094 = v_8027 & v_8093;
assign v_8095 = v_8032 & v_8094;
assign v_8096 = v_8037 & v_8095;
assign v_8105 = v_8024 & v_8104;
assign v_8106 = v_8027 & v_8105;
assign v_8107 = v_8032 & v_8106;
assign v_8108 = v_8037 & v_8107;
assign v_8117 = v_8024 & v_8116;
assign v_8118 = v_91 & v_8040;
assign v_8120 = v_8027 & v_8119;
assign v_8121 = v_7571 & v_8042;
assign v_8123 = v_8032 & v_8122;
assign v_8124 = v_8030 & v_8047;
assign v_8126 = v_8037 & v_8125;
assign v_8127 = v_8035 & v_8052;
assign v_8132 = v_8130 & v_8131;
assign v_8135 = v_8133 & v_8134;
assign v_8138 = v_8136 & v_8137;
assign v_8141 = v_8139 & v_8140;
assign v_8145 = v_8024 & v_8144;
assign v_8146 = v_8027 & v_8145;
assign v_8147 = v_8032 & v_8146;
assign v_8148 = v_8037 & v_8147;
assign v_8159 = v_8157 & v_8158;
assign v_8162 = v_8160 & v_8161;
assign v_8164 = v_8162 & v_8163;
assign v_8171 = v_8167 & v_8170;
assign v_8173 = v_8164 & v_8172;
assign v_8180 = v_8176 & v_8179;
assign v_8182 = v_8173 & v_8181;
assign v_8184 = v_89 & v_7899;
assign v_8185 = ~v_91 & v_8184;
assign v_8186 = v_91 & v_7900;
assign v_8188 = v_96 & v_8187;
assign v_8190 = v_807 & v_7606;
assign v_8192 = ~v_87 & v_7615;
assign v_8193 = ~v_89 & v_8192;
assign v_8194 = ~v_91 & v_8193;
assign v_8195 = ~v_87 & v_7620;
assign v_8196 = ~v_89 & v_8195;
assign v_8197 = ~v_91 & v_8196;
assign v_8199 = v_361 & v_8198;
assign v_8201 = ~v_87 & v_7628;
assign v_8202 = ~v_89 & v_8201;
assign v_8203 = ~v_91 & v_8202;
assign v_8204 = ~v_87 & v_7633;
assign v_8205 = ~v_89 & v_8204;
assign v_8206 = ~v_91 & v_8205;
assign v_8208 = v_563 & v_8207;
assign v_8213 = v_8160 & v_8212;
assign v_8214 = v_8163 & v_8213;
assign v_8215 = v_8172 & v_8214;
assign v_8216 = v_8181 & v_8215;
assign v_8225 = v_8160 & v_8224;
assign v_8226 = v_8163 & v_8225;
assign v_8227 = v_8172 & v_8226;
assign v_8228 = v_8181 & v_8227;
assign v_8237 = v_8160 & v_8236;
assign v_8238 = v_8163 & v_8237;
assign v_8239 = v_8172 & v_8238;
assign v_8240 = v_8181 & v_8239;
assign v_8249 = v_8160 & v_8248;
assign v_8250 = v_8163 & v_8249;
assign v_8251 = v_8172 & v_8250;
assign v_8252 = v_8181 & v_8251;
assign v_8261 = v_8160 & v_8260;
assign v_8262 = v_8163 & v_8261;
assign v_8263 = v_8172 & v_8262;
assign v_8264 = v_8181 & v_8263;
assign v_8273 = v_8160 & v_8272;
assign v_8274 = v_8158 & v_8188;
assign v_8276 = v_8163 & v_8275;
assign v_8277 = ~v_91 & v_8190;
assign v_8279 = v_8172 & v_8278;
assign v_8280 = v_8170 & v_8199;
assign v_8282 = v_8181 & v_8281;
assign v_8283 = v_8179 & v_8208;
assign v_8288 = v_8286 & v_8287;
assign v_8291 = v_8289 & v_8290;
assign v_8294 = v_8292 & v_8293;
assign v_8297 = v_8295 & v_8296;
assign v_8301 = v_8160 & v_8300;
assign v_8302 = v_8163 & v_8301;
assign v_8303 = v_8172 & v_8302;
assign v_8304 = v_8181 & v_8303;
assign v_8314 = v_8312 & v_8313;
assign v_8316 = v_8314 & v_8315;
assign v_8319 = v_8317 & v_8318;
assign v_8321 = v_8316 & v_8320;
assign v_8324 = v_8322 & v_8323;
assign v_8326 = v_8321 & v_8325;
assign v_8328 = v_96 & v_8184;
assign v_8330 = v_807 & v_7903;
assign v_8332 = v_91 & v_8193;
assign v_8333 = v_91 & v_8196;
assign v_8335 = v_361 & v_8334;
assign v_8337 = v_91 & v_8202;
assign v_8338 = v_91 & v_8205;
assign v_8340 = v_563 & v_8339;
assign v_8345 = v_8312 & v_8344;
assign v_8346 = v_8315 & v_8345;
assign v_8347 = v_8320 & v_8346;
assign v_8348 = v_8325 & v_8347;
assign v_8357 = v_8312 & v_8356;
assign v_8358 = v_8315 & v_8357;
assign v_8359 = v_8320 & v_8358;
assign v_8360 = v_8325 & v_8359;
assign v_8369 = v_8312 & v_8368;
assign v_8370 = v_8315 & v_8369;
assign v_8371 = v_8320 & v_8370;
assign v_8372 = v_8325 & v_8371;
assign v_8381 = v_8312 & v_8380;
assign v_8382 = v_8315 & v_8381;
assign v_8383 = v_8320 & v_8382;
assign v_8384 = v_8325 & v_8383;
assign v_8393 = v_8312 & v_8392;
assign v_8394 = v_8315 & v_8393;
assign v_8395 = v_8320 & v_8394;
assign v_8396 = v_8325 & v_8395;
assign v_8405 = v_8312 & v_8404;
assign v_8406 = v_91 & v_8328;
assign v_8408 = v_8315 & v_8407;
assign v_8409 = v_7876 & v_8330;
assign v_8411 = v_8320 & v_8410;
assign v_8412 = v_8318 & v_8335;
assign v_8414 = v_8325 & v_8413;
assign v_8415 = v_8323 & v_8340;
assign v_8420 = v_8418 & v_8419;
assign v_8423 = v_8421 & v_8422;
assign v_8426 = v_8424 & v_8425;
assign v_8429 = v_8427 & v_8428;
assign v_8433 = v_8312 & v_8432;
assign v_8434 = v_8315 & v_8433;
assign v_8435 = v_8320 & v_8434;
assign v_8436 = v_8325 & v_8435;
assign v_8449 = v_8447 & v_8448;
assign v_8452 = v_8450 & v_8451;
assign v_8454 = v_8452 & v_8453;
assign v_8459 = v_8456 & v_8458;
assign v_8461 = v_8454 & v_8460;
assign v_8466 = v_8463 & v_8465;
assign v_8468 = v_8461 & v_8467;
assign v_8470 = v_85 & v_7311;
assign v_8471 = v_87 & v_8470;
assign v_8472 = ~v_89 & v_8471;
assign v_8473 = ~v_91 & v_8472;
assign v_8474 = v_91 & v_8184;
assign v_8476 = v_96 & v_8475;
assign v_8478 = v_807 & v_7900;
assign v_8480 = v_89 & v_8192;
assign v_8481 = ~v_91 & v_8480;
assign v_8482 = v_89 & v_8195;
assign v_8483 = ~v_91 & v_8482;
assign v_8485 = v_361 & v_8484;
assign v_8487 = v_89 & v_8201;
assign v_8488 = ~v_91 & v_8487;
assign v_8489 = v_89 & v_8204;
assign v_8490 = ~v_91 & v_8489;
assign v_8492 = v_563 & v_8491;
assign v_8497 = v_8450 & v_8496;
assign v_8498 = v_8453 & v_8497;
assign v_8499 = v_8460 & v_8498;
assign v_8500 = v_8467 & v_8499;
assign v_8509 = v_8450 & v_8508;
assign v_8510 = v_8453 & v_8509;
assign v_8511 = v_8460 & v_8510;
assign v_8512 = v_8467 & v_8511;
assign v_8521 = v_8450 & v_8520;
assign v_8522 = v_8453 & v_8521;
assign v_8523 = v_8460 & v_8522;
assign v_8524 = v_8467 & v_8523;
assign v_8533 = v_8450 & v_8532;
assign v_8534 = v_8453 & v_8533;
assign v_8535 = v_8460 & v_8534;
assign v_8536 = v_8467 & v_8535;
assign v_8545 = v_8450 & v_8544;
assign v_8546 = v_8453 & v_8545;
assign v_8547 = v_8460 & v_8546;
assign v_8548 = v_8467 & v_8547;
assign v_8557 = v_8450 & v_8556;
assign v_8558 = v_8448 & v_8476;
assign v_8560 = v_8453 & v_8559;
assign v_8561 = ~v_91 & v_8478;
assign v_8563 = v_8460 & v_8562;
assign v_8564 = v_8458 & v_8485;
assign v_8566 = v_8467 & v_8565;
assign v_8567 = v_8465 & v_8492;
assign v_8572 = v_8570 & v_8571;
assign v_8575 = v_8573 & v_8574;
assign v_8578 = v_8576 & v_8577;
assign v_8581 = v_8579 & v_8580;
assign v_8590 = v_8450 & ~v_8584;
assign v_8591 = v_8453 & v_8590;
assign v_8592 = v_8460 & v_8591;
assign v_8593 = v_8467 & v_8592;
assign v_8598 = v_8596 & v_8597;
assign v_8600 = v_8598 & v_8599;
assign v_8603 = v_8601 & v_8602;
assign v_8605 = v_8600 & v_8604;
assign v_8608 = v_8606 & v_8607;
assign v_8610 = v_8605 & v_8609;
assign v_8612 = v_96 & v_8472;
assign v_8614 = v_807 & v_8187;
assign v_8616 = v_91 & v_8480;
assign v_8617 = v_91 & v_8482;
assign v_8619 = v_361 & v_8618;
assign v_8621 = v_91 & v_8487;
assign v_8622 = v_91 & v_8489;
assign v_8624 = v_563 & v_8623;
assign v_8629 = v_8596 & v_8628;
assign v_8630 = v_8599 & v_8629;
assign v_8631 = v_8604 & v_8630;
assign v_8632 = v_8609 & v_8631;
assign v_8641 = v_8596 & v_8640;
assign v_8642 = v_8599 & v_8641;
assign v_8643 = v_8604 & v_8642;
assign v_8644 = v_8609 & v_8643;
assign v_8653 = v_8596 & v_8652;
assign v_8654 = v_8599 & v_8653;
assign v_8655 = v_8604 & v_8654;
assign v_8656 = v_8609 & v_8655;
assign v_8665 = v_8596 & v_8664;
assign v_8666 = v_8599 & v_8665;
assign v_8667 = v_8604 & v_8666;
assign v_8668 = v_8609 & v_8667;
assign v_8677 = v_8596 & v_8676;
assign v_8678 = v_8599 & v_8677;
assign v_8679 = v_8604 & v_8678;
assign v_8680 = v_8609 & v_8679;
assign v_8689 = v_8596 & v_8688;
assign v_8690 = v_91 & v_8612;
assign v_8692 = v_8599 & v_8691;
assign v_8693 = v_8157 & v_8614;
assign v_8695 = v_8604 & v_8694;
assign v_8696 = v_8602 & v_8619;
assign v_8698 = v_8609 & v_8697;
assign v_8699 = v_8607 & v_8624;
assign v_8704 = v_8702 & v_8703;
assign v_8707 = v_8705 & v_8706;
assign v_8710 = v_8708 & v_8709;
assign v_8713 = v_8711 & v_8712;
assign v_8722 = v_8596 & ~v_8716;
assign v_8723 = v_8599 & v_8722;
assign v_8724 = v_8604 & v_8723;
assign v_8725 = v_8609 & v_8724;
assign v_8731 = v_8729 & v_8730;
assign v_8734 = v_8732 & v_8733;
assign v_8736 = v_8734 & v_8735;
assign v_8745 = v_8740 & v_8744;
assign v_8747 = v_8736 & v_8746;
assign v_8756 = v_8751 & v_8755;
assign v_8758 = v_8747 & v_8757;
assign v_8760 = v_89 & v_8471;
assign v_8761 = ~v_91 & v_8760;
assign v_8762 = v_91 & v_8472;
assign v_8764 = v_96 & v_8763;
assign v_8766 = v_807 & v_8184;
assign v_8768 = v_85 & v_7614;
assign v_8769 = v_87 & v_8768;
assign v_8770 = ~v_89 & v_8769;
assign v_8771 = ~v_91 & v_8770;
assign v_8772 = v_355 & v_7619;
assign v_8773 = v_87 & v_8772;
assign v_8774 = ~v_89 & v_8773;
assign v_8775 = ~v_91 & v_8774;
assign v_8777 = v_361 & v_8776;
assign v_8779 = v_85 & v_7627;
assign v_8780 = v_87 & v_8779;
assign v_8781 = ~v_89 & v_8780;
assign v_8782 = ~v_91 & v_8781;
assign v_8783 = v_355 & v_7632;
assign v_8784 = v_87 & v_8783;
assign v_8785 = ~v_89 & v_8784;
assign v_8786 = ~v_91 & v_8785;
assign v_8788 = v_563 & v_8787;
assign v_8793 = v_8732 & v_8792;
assign v_8794 = v_8735 & v_8793;
assign v_8795 = v_8746 & v_8794;
assign v_8796 = v_8757 & v_8795;
assign v_8805 = v_8732 & v_8804;
assign v_8806 = v_8735 & v_8805;
assign v_8807 = v_8746 & v_8806;
assign v_8808 = v_8757 & v_8807;
assign v_8817 = v_8732 & v_8816;
assign v_8818 = v_8735 & v_8817;
assign v_8819 = v_8746 & v_8818;
assign v_8820 = v_8757 & v_8819;
assign v_8829 = v_8732 & v_8828;
assign v_8830 = v_8735 & v_8829;
assign v_8831 = v_8746 & v_8830;
assign v_8832 = v_8757 & v_8831;
assign v_8841 = v_8732 & v_8840;
assign v_8842 = v_8735 & v_8841;
assign v_8843 = v_8746 & v_8842;
assign v_8844 = v_8757 & v_8843;
assign v_8853 = v_8732 & v_8852;
assign v_8854 = v_8730 & v_8764;
assign v_8856 = v_8735 & v_8855;
assign v_8857 = ~v_91 & v_8766;
assign v_8859 = v_8746 & v_8858;
assign v_8860 = v_8744 & v_8777;
assign v_8862 = v_8757 & v_8861;
assign v_8863 = v_8755 & v_8788;
assign v_8868 = v_8866 & v_8867;
assign v_8871 = v_8869 & v_8870;
assign v_8874 = v_8872 & v_8873;
assign v_8877 = v_8875 & v_8876;
assign v_8886 = v_8732 & ~v_8880;
assign v_8887 = v_8735 & v_8886;
assign v_8888 = v_8746 & v_8887;
assign v_8889 = v_8757 & v_8888;
assign v_8894 = v_8892 & v_8893;
assign v_8896 = v_8894 & v_8895;
assign v_8899 = v_8897 & v_8898;
assign v_8901 = v_8896 & v_8900;
assign v_8904 = v_8902 & v_8903;
assign v_8906 = v_8901 & v_8905;
assign v_8908 = v_96 & v_8760;
assign v_8910 = v_807 & v_8475;
assign v_8912 = v_91 & v_8770;
assign v_8913 = v_91 & v_8774;
assign v_8915 = v_361 & v_8914;
assign v_8917 = v_91 & v_8781;
assign v_8918 = v_91 & v_8785;
assign v_8920 = v_563 & v_8919;
assign v_8925 = v_8892 & v_8924;
assign v_8926 = v_8895 & v_8925;
assign v_8927 = v_8900 & v_8926;
assign v_8928 = v_8905 & v_8927;
assign v_8937 = v_8892 & v_8936;
assign v_8938 = v_8895 & v_8937;
assign v_8939 = v_8900 & v_8938;
assign v_8940 = v_8905 & v_8939;
assign v_8949 = v_8892 & v_8948;
assign v_8950 = v_8895 & v_8949;
assign v_8951 = v_8900 & v_8950;
assign v_8952 = v_8905 & v_8951;
assign v_8961 = v_8892 & v_8960;
assign v_8962 = v_8895 & v_8961;
assign v_8963 = v_8900 & v_8962;
assign v_8964 = v_8905 & v_8963;
assign v_8973 = v_8892 & v_8972;
assign v_8974 = v_8895 & v_8973;
assign v_8975 = v_8900 & v_8974;
assign v_8976 = v_8905 & v_8975;
assign v_8985 = v_8892 & v_8984;
assign v_8986 = v_91 & v_8908;
assign v_8988 = v_8895 & v_8987;
assign v_8989 = v_8447 & v_8910;
assign v_8991 = v_8900 & v_8990;
assign v_8992 = v_8898 & v_8915;
assign v_8994 = v_8905 & v_8993;
assign v_8995 = v_8903 & v_8920;
assign v_9000 = v_8998 & v_8999;
assign v_9003 = v_9001 & v_9002;
assign v_9006 = v_9004 & v_9005;
assign v_9009 = v_9007 & v_9008;
assign v_9018 = v_8892 & ~v_9012;
assign v_9019 = v_8895 & v_9018;
assign v_9020 = v_8900 & v_9019;
assign v_9021 = v_8905 & v_9020;
assign v_9028 = v_9026 & v_9027;
assign v_9031 = v_9029 & v_9030;
assign v_9033 = v_9031 & v_9032;
assign v_9038 = v_9035 & v_9037;
assign v_9040 = v_9033 & v_9039;
assign v_9045 = v_9042 & v_9044;
assign v_9047 = v_9040 & v_9046;
assign v_9049 = ~v_87 & v_8470;
assign v_9050 = ~v_89 & v_9049;
assign v_9051 = ~v_91 & v_9050;
assign v_9052 = v_91 & v_8760;
assign v_9054 = v_96 & v_9053;
assign v_9056 = v_807 & v_8472;
assign v_9058 = v_89 & v_8769;
assign v_9059 = ~v_91 & v_9058;
assign v_9060 = v_89 & v_8773;
assign v_9061 = ~v_91 & v_9060;
assign v_9063 = v_361 & v_9062;
assign v_9065 = v_89 & v_8780;
assign v_9066 = ~v_91 & v_9065;
assign v_9067 = v_89 & v_8784;
assign v_9068 = ~v_91 & v_9067;
assign v_9070 = v_563 & v_9069;
assign v_9075 = v_9029 & v_9074;
assign v_9076 = v_9032 & v_9075;
assign v_9077 = v_9039 & v_9076;
assign v_9078 = v_9046 & v_9077;
assign v_9087 = v_9029 & v_9086;
assign v_9088 = v_9032 & v_9087;
assign v_9089 = v_9039 & v_9088;
assign v_9090 = v_9046 & v_9089;
assign v_9099 = v_9029 & v_9098;
assign v_9100 = v_9032 & v_9099;
assign v_9101 = v_9039 & v_9100;
assign v_9102 = v_9046 & v_9101;
assign v_9111 = v_9029 & v_9110;
assign v_9112 = v_9032 & v_9111;
assign v_9113 = v_9039 & v_9112;
assign v_9114 = v_9046 & v_9113;
assign v_9123 = v_9029 & v_9122;
assign v_9124 = v_9032 & v_9123;
assign v_9125 = v_9039 & v_9124;
assign v_9126 = v_9046 & v_9125;
assign v_9135 = v_9029 & v_9134;
assign v_9136 = v_9027 & v_9054;
assign v_9138 = v_9032 & v_9137;
assign v_9139 = ~v_91 & v_9056;
assign v_9141 = v_9039 & v_9140;
assign v_9142 = v_9037 & v_9063;
assign v_9144 = v_9046 & v_9143;
assign v_9145 = v_9044 & v_9070;
assign v_9150 = v_9148 & v_9149;
assign v_9153 = v_9151 & v_9152;
assign v_9156 = v_9154 & v_9155;
assign v_9159 = v_9157 & v_9158;
assign v_9168 = v_9029 & ~v_9162;
assign v_9169 = v_9032 & v_9168;
assign v_9170 = v_9039 & v_9169;
assign v_9171 = v_9046 & v_9170;
assign v_9176 = v_9174 & v_9175;
assign v_9178 = v_9176 & v_9177;
assign v_9181 = v_9179 & v_9180;
assign v_9183 = v_9178 & v_9182;
assign v_9186 = v_9184 & v_9185;
assign v_9188 = v_9183 & v_9187;
assign v_9190 = v_96 & v_9050;
assign v_9192 = v_807 & v_8763;
assign v_9194 = v_91 & v_9058;
assign v_9195 = v_91 & v_9060;
assign v_9197 = v_361 & v_9196;
assign v_9199 = v_91 & v_9065;
assign v_9200 = v_91 & v_9067;
assign v_9202 = v_563 & v_9201;
assign v_9207 = v_9174 & v_9206;
assign v_9208 = v_9177 & v_9207;
assign v_9209 = v_9182 & v_9208;
assign v_9210 = v_9187 & v_9209;
assign v_9219 = v_9174 & v_9218;
assign v_9220 = v_9177 & v_9219;
assign v_9221 = v_9182 & v_9220;
assign v_9222 = v_9187 & v_9221;
assign v_9231 = v_9174 & v_9230;
assign v_9232 = v_9177 & v_9231;
assign v_9233 = v_9182 & v_9232;
assign v_9234 = v_9187 & v_9233;
assign v_9243 = v_9174 & v_9242;
assign v_9244 = v_9177 & v_9243;
assign v_9245 = v_9182 & v_9244;
assign v_9246 = v_9187 & v_9245;
assign v_9255 = v_9174 & v_9254;
assign v_9256 = v_9177 & v_9255;
assign v_9257 = v_9182 & v_9256;
assign v_9258 = v_9187 & v_9257;
assign v_9267 = v_9174 & v_9266;
assign v_9268 = v_91 & v_9190;
assign v_9270 = v_9177 & v_9269;
assign v_9271 = v_8729 & v_9192;
assign v_9273 = v_9182 & v_9272;
assign v_9274 = v_9180 & v_9197;
assign v_9276 = v_9187 & v_9275;
assign v_9277 = v_9185 & v_9202;
assign v_9282 = v_9280 & v_9281;
assign v_9285 = v_9283 & v_9284;
assign v_9288 = v_9286 & v_9287;
assign v_9291 = v_9289 & v_9290;
assign v_9300 = v_9174 & ~v_9294;
assign v_9301 = v_9177 & v_9300;
assign v_9302 = v_9182 & v_9301;
assign v_9303 = v_9187 & v_9302;
assign v_9309 = v_9307 & v_9308;
assign v_9312 = v_9310 & v_9311;
assign v_9314 = v_9312 & v_9313;
assign v_9321 = v_9317 & v_9320;
assign v_9323 = v_9314 & v_9322;
assign v_9330 = v_9326 & v_9329;
assign v_9332 = v_9323 & v_9331;
assign v_9334 = v_89 & v_9049;
assign v_9335 = ~v_91 & v_9334;
assign v_9336 = v_91 & v_9050;
assign v_9338 = v_96 & v_9337;
assign v_9340 = v_807 & v_8760;
assign v_9342 = ~v_87 & v_8768;
assign v_9343 = ~v_89 & v_9342;
assign v_9344 = ~v_91 & v_9343;
assign v_9345 = ~v_87 & v_8772;
assign v_9346 = ~v_89 & v_9345;
assign v_9347 = ~v_91 & v_9346;
assign v_9349 = v_361 & v_9348;
assign v_9351 = ~v_87 & v_8779;
assign v_9352 = ~v_89 & v_9351;
assign v_9353 = ~v_91 & v_9352;
assign v_9354 = ~v_87 & v_8783;
assign v_9355 = ~v_89 & v_9354;
assign v_9356 = ~v_91 & v_9355;
assign v_9358 = v_563 & v_9357;
assign v_9363 = v_9310 & v_9362;
assign v_9364 = v_9313 & v_9363;
assign v_9365 = v_9322 & v_9364;
assign v_9366 = v_9331 & v_9365;
assign v_9375 = v_9310 & v_9374;
assign v_9376 = v_9313 & v_9375;
assign v_9377 = v_9322 & v_9376;
assign v_9378 = v_9331 & v_9377;
assign v_9387 = v_9310 & v_9386;
assign v_9388 = v_9313 & v_9387;
assign v_9389 = v_9322 & v_9388;
assign v_9390 = v_9331 & v_9389;
assign v_9399 = v_9310 & v_9398;
assign v_9400 = v_9313 & v_9399;
assign v_9401 = v_9322 & v_9400;
assign v_9402 = v_9331 & v_9401;
assign v_9411 = v_9310 & v_9410;
assign v_9412 = v_9313 & v_9411;
assign v_9413 = v_9322 & v_9412;
assign v_9414 = v_9331 & v_9413;
assign v_9423 = v_9310 & v_9422;
assign v_9424 = v_9308 & v_9338;
assign v_9426 = v_9313 & v_9425;
assign v_9427 = ~v_91 & v_9340;
assign v_9429 = v_9322 & v_9428;
assign v_9430 = v_9320 & v_9349;
assign v_9432 = v_9331 & v_9431;
assign v_9433 = v_9329 & v_9358;
assign v_9438 = v_9436 & v_9437;
assign v_9441 = v_9439 & v_9440;
assign v_9444 = v_9442 & v_9443;
assign v_9447 = v_9445 & v_9446;
assign v_9456 = v_9310 & ~v_9450;
assign v_9457 = v_9313 & v_9456;
assign v_9458 = v_9322 & v_9457;
assign v_9459 = v_9331 & v_9458;
assign v_9464 = v_9462 & v_9463;
assign v_9466 = v_9464 & v_9465;
assign v_9469 = v_9467 & v_9468;
assign v_9471 = v_9466 & v_9470;
assign v_9474 = v_9472 & v_9473;
assign v_9476 = v_9471 & v_9475;
assign v_9478 = v_96 & v_9334;
assign v_9480 = v_807 & v_9053;
assign v_9482 = v_91 & v_9343;
assign v_9483 = v_91 & v_9346;
assign v_9485 = v_361 & v_9484;
assign v_9487 = v_91 & v_9352;
assign v_9488 = v_91 & v_9355;
assign v_9490 = v_563 & v_9489;
assign v_9495 = v_9462 & v_9494;
assign v_9496 = v_9465 & v_9495;
assign v_9497 = v_9470 & v_9496;
assign v_9498 = v_9475 & v_9497;
assign v_9507 = v_9462 & v_9506;
assign v_9508 = v_9465 & v_9507;
assign v_9509 = v_9470 & v_9508;
assign v_9510 = v_9475 & v_9509;
assign v_9519 = v_9462 & v_9518;
assign v_9520 = v_9465 & v_9519;
assign v_9521 = v_9470 & v_9520;
assign v_9522 = v_9475 & v_9521;
assign v_9531 = v_9462 & v_9530;
assign v_9532 = v_9465 & v_9531;
assign v_9533 = v_9470 & v_9532;
assign v_9534 = v_9475 & v_9533;
assign v_9543 = v_9462 & v_9542;
assign v_9544 = v_9465 & v_9543;
assign v_9545 = v_9470 & v_9544;
assign v_9546 = v_9475 & v_9545;
assign v_9555 = v_9462 & v_9554;
assign v_9556 = v_91 & v_9478;
assign v_9558 = v_9465 & v_9557;
assign v_9559 = v_9026 & v_9480;
assign v_9561 = v_9470 & v_9560;
assign v_9562 = v_9468 & v_9485;
assign v_9564 = v_9475 & v_9563;
assign v_9565 = v_9473 & v_9490;
assign v_9570 = v_9568 & v_9569;
assign v_9573 = v_9571 & v_9572;
assign v_9576 = v_9574 & v_9575;
assign v_9579 = v_9577 & v_9578;
assign v_9588 = v_9462 & ~v_9582;
assign v_9589 = v_9465 & v_9588;
assign v_9590 = v_9470 & v_9589;
assign v_9591 = v_9475 & v_9590;
assign v_9602 = v_9600 & v_9601;
assign v_9605 = v_9603 & v_9604;
assign v_9607 = v_9605 & v_9606;
assign v_9612 = v_9609 & v_9611;
assign v_9614 = v_9607 & v_9613;
assign v_9619 = v_9616 & v_9618;
assign v_9621 = v_9614 & v_9620;
assign v_9623 = v_76 & v_576;
assign v_9624 = v_581 & v_9623;
assign v_9625 = v_584 & v_9624;
assign v_9626 = v_587 & v_9625;
assign v_9627 = v_87 & v_9626;
assign v_9628 = ~v_89 & v_9627;
assign v_9629 = ~v_91 & v_9628;
assign v_9630 = v_91 & v_9334;
assign v_9632 = v_96 & v_9631;
assign v_9634 = v_807 & v_9050;
assign v_9636 = v_89 & v_9342;
assign v_9637 = ~v_91 & v_9636;
assign v_9638 = v_89 & v_9345;
assign v_9639 = ~v_91 & v_9638;
assign v_9641 = v_361 & v_9640;
assign v_9643 = v_89 & v_9351;
assign v_9644 = ~v_91 & v_9643;
assign v_9645 = v_89 & v_9354;
assign v_9646 = ~v_91 & v_9645;
assign v_9648 = v_563 & v_9647;
assign v_9653 = v_9603 & v_9652;
assign v_9654 = v_9606 & v_9653;
assign v_9655 = v_9613 & v_9654;
assign v_9656 = v_9620 & v_9655;
assign v_9665 = v_9603 & v_9664;
assign v_9666 = v_9606 & v_9665;
assign v_9667 = v_9613 & v_9666;
assign v_9668 = v_9620 & v_9667;
assign v_9677 = v_9603 & v_9676;
assign v_9678 = v_9606 & v_9677;
assign v_9679 = v_9613 & v_9678;
assign v_9680 = v_9620 & v_9679;
assign v_9689 = v_9603 & v_9688;
assign v_9690 = v_9606 & v_9689;
assign v_9691 = v_9613 & v_9690;
assign v_9692 = v_9620 & v_9691;
assign v_9701 = v_9603 & v_9700;
assign v_9702 = v_9606 & v_9701;
assign v_9703 = v_9613 & v_9702;
assign v_9704 = v_9620 & v_9703;
assign v_9713 = v_9603 & v_9712;
assign v_9714 = v_9601 & v_9632;
assign v_9716 = v_9606 & v_9715;
assign v_9717 = ~v_91 & v_9634;
assign v_9719 = v_9613 & v_9718;
assign v_9720 = v_9611 & v_9641;
assign v_9722 = v_9620 & v_9721;
assign v_9723 = v_9618 & v_9648;
assign v_9728 = v_9726 & v_9727;
assign v_9731 = v_9729 & v_9730;
assign v_9734 = v_9732 & v_9733;
assign v_9737 = v_9735 & v_9736;
assign v_9746 = v_9603 & ~v_9740;
assign v_9747 = v_9606 & v_9746;
assign v_9748 = v_9613 & v_9747;
assign v_9749 = v_9620 & v_9748;
assign v_9754 = v_9752 & v_9753;
assign v_9756 = v_9754 & v_9755;
assign v_9759 = v_9757 & v_9758;
assign v_9761 = v_9756 & v_9760;
assign v_9764 = v_9762 & v_9763;
assign v_9766 = v_9761 & v_9765;
assign v_9768 = v_96 & v_9628;
assign v_9770 = v_807 & v_9337;
assign v_9772 = v_91 & v_9636;
assign v_9773 = v_91 & v_9638;
assign v_9775 = v_361 & v_9774;
assign v_9777 = v_91 & v_9643;
assign v_9778 = v_91 & v_9645;
assign v_9780 = v_563 & v_9779;
assign v_9785 = v_9752 & v_9784;
assign v_9786 = v_9755 & v_9785;
assign v_9787 = v_9760 & v_9786;
assign v_9788 = v_9765 & v_9787;
assign v_9797 = v_9752 & v_9796;
assign v_9798 = v_9755 & v_9797;
assign v_9799 = v_9760 & v_9798;
assign v_9800 = v_9765 & v_9799;
assign v_9809 = v_9752 & v_9808;
assign v_9810 = v_9755 & v_9809;
assign v_9811 = v_9760 & v_9810;
assign v_9812 = v_9765 & v_9811;
assign v_9821 = v_9752 & v_9820;
assign v_9822 = v_9755 & v_9821;
assign v_9823 = v_9760 & v_9822;
assign v_9824 = v_9765 & v_9823;
assign v_9833 = v_9752 & v_9832;
assign v_9834 = v_9755 & v_9833;
assign v_9835 = v_9760 & v_9834;
assign v_9836 = v_9765 & v_9835;
assign v_9845 = v_9752 & v_9844;
assign v_9846 = v_91 & v_9768;
assign v_9848 = v_9755 & v_9847;
assign v_9849 = v_9307 & v_9770;
assign v_9851 = v_9760 & v_9850;
assign v_9852 = v_9758 & v_9775;
assign v_9854 = v_9765 & v_9853;
assign v_9855 = v_9763 & v_9780;
assign v_9860 = v_9858 & v_9859;
assign v_9863 = v_9861 & v_9862;
assign v_9866 = v_9864 & v_9865;
assign v_9869 = v_9867 & v_9868;
assign v_9878 = v_9752 & ~v_9872;
assign v_9879 = v_9755 & v_9878;
assign v_9880 = v_9760 & v_9879;
assign v_9881 = v_9765 & v_9880;
assign v_9885 = v_9 & ~v_9884;
assign v_9893 = ~v_89 & ~v_91;
assign v_9894 = v_87 & v_9893;
assign v_9895 = ~v_29 & v_9894;
assign v_9896 = ~v_24 & v_9895;
assign v_9897 = ~v_19 & v_9896;
assign v_9898 = ~v_14 & v_9897;
assign v_9900 = v_9892 & v_9899;
assign v_9901 = v_9884 & v_9900;
assign v_9904 = v_9902 & ~v_9903;
assign v_9905 = v_89 & v_91;
assign v_9906 = ~v_87 & v_9905;
assign v_9907 = v_29 & v_9906;
assign v_9908 = v_24 & v_9907;
assign v_9909 = v_19 & v_9908;
assign v_9910 = v_14 & v_9909;
assign v_9919 = v_9911 & v_9918;
assign v_9920 = v_9903 & v_9919;
assign v_9922 = ~v_96 & v_9921;
assign v_9923 = v_96 & v_9900;
assign v_9925 = ~v_807 & v_9924;
assign v_9926 = v_807 & v_9919;
assign v_9930 = v_9 & v_9898;
assign v_9931 = ~v_9 & v_9891;
assign v_9934 = v_9929 & v_9933;
assign v_9936 = ~v_9 & v_9917;
assign v_9937 = v_9 & v_9910;
assign v_9940 = v_9935 & v_9939;
assign v_9943 = v_9941 & v_9942;
assign v_9946 = v_9944 & v_9945;
assign v_9949 = v_14 & ~v_9884;
assign v_9952 = v_9950 & v_9951;
assign v_9953 = v_9884 & v_9952;
assign v_9955 = ~v_9903 & v_9954;
assign v_9957 = v_9917 & v_9956;
assign v_9958 = v_9903 & v_9957;
assign v_9960 = ~v_96 & v_9959;
assign v_9961 = v_96 & v_9952;
assign v_9963 = ~v_807 & v_9962;
assign v_9964 = v_807 & v_9957;
assign v_9968 = v_14 & v_9897;
assign v_9969 = ~v_14 & v_9890;
assign v_9972 = v_9967 & v_9971;
assign v_9974 = ~v_14 & v_9916;
assign v_9977 = v_9973 & v_9976;
assign v_9980 = v_9978 & v_9979;
assign v_9983 = v_9981 & v_9982;
assign v_9986 = v_19 & ~v_9884;
assign v_9989 = v_9987 & v_9988;
assign v_9990 = v_9884 & v_9989;
assign v_9992 = ~v_9903 & v_9991;
assign v_9994 = v_9916 & v_9993;
assign v_9995 = v_9903 & v_9994;
assign v_9997 = ~v_96 & v_9996;
assign v_9998 = v_96 & v_9989;
assign v_10000 = ~v_807 & v_9999;
assign v_10001 = v_807 & v_9994;
assign v_10005 = v_19 & v_9896;
assign v_10006 = ~v_19 & v_9889;
assign v_10009 = v_10004 & v_10008;
assign v_10011 = ~v_19 & v_9915;
assign v_10014 = v_10010 & v_10013;
assign v_10017 = v_10015 & v_10016;
assign v_10020 = v_10018 & v_10019;
assign v_10023 = v_24 & ~v_9884;
assign v_10026 = v_10024 & v_10025;
assign v_10027 = v_9884 & v_10026;
assign v_10029 = ~v_9903 & v_10028;
assign v_10031 = v_9915 & v_10030;
assign v_10032 = v_9903 & v_10031;
assign v_10034 = ~v_96 & v_10033;
assign v_10035 = v_96 & v_10026;
assign v_10037 = ~v_807 & v_10036;
assign v_10038 = v_807 & v_10031;
assign v_10042 = v_24 & v_9895;
assign v_10043 = ~v_24 & v_9888;
assign v_10046 = v_10041 & v_10045;
assign v_10048 = ~v_24 & v_9914;
assign v_10051 = v_10047 & v_10050;
assign v_10054 = v_10052 & v_10053;
assign v_10057 = v_10055 & v_10056;
assign v_10060 = v_29 & ~v_9884;
assign v_10063 = v_10061 & v_10062;
assign v_10064 = v_9884 & v_10063;
assign v_10066 = ~v_9903 & v_10065;
assign v_10068 = v_9914 & v_10067;
assign v_10069 = v_9903 & v_10068;
assign v_10071 = ~v_96 & v_10070;
assign v_10072 = v_96 & v_10063;
assign v_10074 = ~v_807 & v_10073;
assign v_10075 = v_807 & v_10068;
assign v_10079 = v_29 & v_9894;
assign v_10080 = ~v_29 & v_9887;
assign v_10083 = v_10078 & v_10082;
assign v_10085 = ~v_29 & v_9913;
assign v_10088 = v_10084 & v_10087;
assign v_10091 = v_10089 & v_10090;
assign v_10094 = v_10092 & v_10093;
assign v_10098 = ~v_87 & v_9893;
assign v_10099 = v_87 & v_9886;
assign v_10102 = v_10097 & v_10101;
assign v_10104 = v_87 & v_9912;
assign v_10107 = v_10103 & v_10106;
assign v_10110 = v_10108 & v_10109;
assign v_10113 = v_10111 & v_10112;
assign v_10115 = ~v_87 & ~v_9884;
assign v_10118 = v_10116 & v_10117;
assign v_10119 = v_9884 & v_10118;
assign v_10121 = ~v_9903 & v_10120;
assign v_10123 = v_9913 & v_10122;
assign v_10124 = v_9903 & v_10123;
assign v_10126 = ~v_96 & v_10125;
assign v_10127 = v_96 & v_10118;
assign v_10129 = ~v_807 & v_10128;
assign v_10130 = v_807 & v_10123;
assign v_10134 = v_89 & ~v_9884;
assign v_10137 = v_10135 & v_10136;
assign v_10138 = v_9884 & v_10137;
assign v_10140 = ~v_9903 & v_10139;
assign v_10141 = v_9886 & v_9912;
assign v_10142 = v_9903 & v_10141;
assign v_10144 = ~v_96 & v_10143;
assign v_10145 = v_96 & v_10137;
assign v_10147 = ~v_807 & v_10146;
assign v_10148 = v_807 & v_10141;
assign v_10152 = v_89 & ~v_91;
assign v_10153 = ~v_89 & v_91;
assign v_10156 = v_10151 & v_10155;
assign v_10160 = v_10157 & v_10159;
assign v_10163 = v_10161 & v_10162;
assign v_10166 = v_10164 & v_10165;
assign v_10169 = v_91 & ~v_9884;
assign v_10170 = ~v_91 & v_9884;
assign v_10172 = ~v_9903 & v_10171;
assign v_10173 = ~v_91 & v_9903;
assign v_10175 = ~v_96 & v_10174;
assign v_10176 = ~v_91 & v_96;
assign v_10178 = ~v_807 & v_10177;
assign v_10179 = ~v_91 & v_807;
assign v_10184 = v_10182 & v_10183;
assign v_10187 = v_10185 & v_10186;
assign v_10190 = v_10188 & v_10189;
assign v_10193 = v_10191 & v_10192;
assign v_10197 = v_47 & ~v_10196;
assign v_10198 = v_301 & v_10196;
assign v_10201 = v_10199 & ~v_10200;
assign v_10202 = v_468 & v_10200;
assign v_10204 = ~v_361 & v_10203;
assign v_10205 = v_301 & v_361;
assign v_10207 = ~v_563 & v_10206;
assign v_10208 = v_468 & v_563;
assign v_10213 = v_10211 & v_10212;
assign v_10216 = v_10214 & v_10215;
assign v_10219 = v_10217 & v_10218;
assign v_10222 = v_10220 & v_10221;
assign v_10225 = v_45 & ~v_10196;
assign v_10226 = v_304 & v_10196;
assign v_10228 = ~v_10200 & v_10227;
assign v_10229 = v_470 & v_10200;
assign v_10231 = ~v_361 & v_10230;
assign v_10232 = v_304 & v_361;
assign v_10234 = ~v_563 & v_10233;
assign v_10235 = v_470 & v_563;
assign v_10240 = v_10238 & v_10239;
assign v_10243 = v_10241 & v_10242;
assign v_10246 = v_10244 & v_10245;
assign v_10249 = v_10247 & v_10248;
assign v_10252 = v_43 & ~v_10196;
assign v_10253 = v_324 & v_10196;
assign v_10255 = ~v_10200 & v_10254;
assign v_10256 = v_510 & v_10200;
assign v_10258 = ~v_361 & v_10257;
assign v_10259 = v_324 & v_361;
assign v_10261 = ~v_563 & v_10260;
assign v_10262 = v_510 & v_563;
assign v_10267 = v_10265 & v_10266;
assign v_10270 = v_10268 & v_10269;
assign v_10273 = v_10271 & v_10272;
assign v_10276 = v_10274 & v_10275;
assign v_10279 = v_8 & ~v_10196;
assign v_10280 = v_249 & v_10196;
assign v_10282 = ~v_10200 & v_10281;
assign v_10283 = v_472 & v_10200;
assign v_10285 = ~v_361 & v_10284;
assign v_10286 = v_249 & v_361;
assign v_10288 = ~v_563 & v_10287;
assign v_10289 = v_472 & v_563;
assign v_10294 = v_10292 & v_10293;
assign v_10297 = v_10295 & v_10296;
assign v_10300 = v_10298 & v_10299;
assign v_10303 = v_10301 & v_10302;
assign v_10306 = v_13 & ~v_10196;
assign v_10307 = v_258 & v_10196;
assign v_10309 = ~v_10200 & v_10308;
assign v_10310 = v_479 & v_10200;
assign v_10312 = ~v_361 & v_10311;
assign v_10313 = v_258 & v_361;
assign v_10315 = ~v_563 & v_10314;
assign v_10316 = v_479 & v_563;
assign v_10321 = v_10319 & v_10320;
assign v_10324 = v_10322 & v_10323;
assign v_10327 = v_10325 & v_10326;
assign v_10330 = v_10328 & v_10329;
assign v_10335 = v_10333 & v_10334;
assign v_10338 = v_10336 & v_10337;
assign v_10341 = v_10339 & v_10340;
assign v_10344 = v_10342 & v_10343;
assign v_10346 = ~v_18 & ~v_10196;
assign v_10347 = v_267 & v_10196;
assign v_10349 = ~v_10200 & v_10348;
assign v_10350 = v_486 & v_10200;
assign v_10352 = ~v_361 & v_10351;
assign v_10353 = v_267 & v_361;
assign v_10355 = ~v_563 & v_10354;
assign v_10356 = v_486 & v_563;
assign v_10362 = v_10360 & v_10361;
assign v_10365 = v_10363 & v_10364;
assign v_10368 = v_10366 & v_10367;
assign v_10371 = v_10369 & v_10370;
assign v_10373 = ~v_23 & ~v_10196;
assign v_10374 = v_276 & v_10196;
assign v_10376 = ~v_10200 & v_10375;
assign v_10377 = v_492 & v_10200;
assign v_10379 = ~v_361 & v_10378;
assign v_10380 = v_276 & v_361;
assign v_10382 = ~v_563 & v_10381;
assign v_10383 = v_492 & v_563;
assign v_10387 = v_28 & ~v_10196;
assign v_10388 = ~v_28 & v_10196;
assign v_10390 = ~v_10200 & v_10389;
assign v_10391 = ~v_28 & v_10200;
assign v_10393 = ~v_361 & v_10392;
assign v_10394 = ~v_28 & v_361;
assign v_10396 = ~v_563 & v_10395;
assign v_10397 = ~v_28 & v_563;
assign v_10402 = v_10400 & v_10401;
assign v_10405 = v_10403 & v_10404;
assign v_10408 = v_10406 & v_10407;
assign v_10411 = v_10409 & v_10410;
assign v_10416 = v_10414 & ~v_10415;
assign v_10422 = ~v_10415 & v_10421;
assign v_10428 = ~v_10415 & v_10427;
assign v_10434 = ~v_10415 & v_10433;
assign v_10440 = ~v_10415 & v_10439;
assign v_10446 = ~v_10415 & v_10445;
assign v_10452 = ~v_10415 & v_10451;
assign v_10459 = ~v_4 & ~v_10415;
assign v_10473 = v_563 & v_10472;
assign v_10474 = v_361 & v_10471;
assign v_10475 = v_807 & v_10470;
assign v_10476 = v_96 & v_10469;
assign v_10477 = v_10200 & v_10468;
assign v_10478 = v_10196 & v_10467;
assign v_10479 = v_9903 & v_10466;
assign v_10480 = v_9884 & v_10415;
assign v_10488 = ~v_9884 & ~v_10415;
assign v_10489 = ~v_9903 & v_10488;
assign v_10490 = ~v_10196 & v_10489;
assign v_10491 = ~v_10200 & v_10490;
assign v_10492 = ~v_96 & v_10491;
assign v_10493 = ~v_807 & v_10492;
assign v_10494 = ~v_361 & v_10493;
assign v_10495 = ~v_563 & v_10494;
assign v_10496 = v_9616 & v_9784;
assign v_10497 = v_9644 & v_9652;
assign v_10499 = v_9472 & v_10498;
assign v_10500 = v_9487 & v_9494;
assign v_10502 = v_9326 & v_10501;
assign v_10503 = v_9353 & v_9362;
assign v_10505 = v_9184 & v_10504;
assign v_10506 = v_9199 & v_9206;
assign v_10508 = v_9042 & v_10507;
assign v_10509 = v_9066 & v_9074;
assign v_10511 = v_8902 & v_10510;
assign v_10512 = v_8917 & v_8924;
assign v_10514 = v_8751 & v_10513;
assign v_10515 = v_8782 & v_8792;
assign v_10517 = v_8606 & v_10516;
assign v_10518 = v_8621 & v_8628;
assign v_10520 = v_8463 & v_10519;
assign v_10521 = v_8488 & v_8496;
assign v_10523 = v_8322 & v_10522;
assign v_10524 = v_8337 & v_8344;
assign v_10526 = v_8176 & v_10525;
assign v_10527 = v_8203 & v_8212;
assign v_10529 = v_8034 & v_10528;
assign v_10530 = v_8049 & v_8056;
assign v_10532 = v_7892 & v_10531;
assign v_10533 = v_7916 & v_7924;
assign v_10535 = v_7752 & v_10534;
assign v_10536 = v_7767 & v_7774;
assign v_10538 = v_7596 & v_10537;
assign v_10539 = v_7631 & v_7642;
assign v_10541 = v_7448 & v_10540;
assign v_10542 = v_7463 & v_7470;
assign v_10544 = v_7304 & v_10543;
assign v_10545 = v_7330 & v_7338;
assign v_10547 = v_7162 & v_10546;
assign v_10548 = v_7177 & v_7184;
assign v_10550 = v_7016 & v_10549;
assign v_10551 = v_7043 & v_7052;
assign v_10553 = v_6874 & v_10552;
assign v_10554 = v_6889 & v_6896;
assign v_10556 = v_6732 & v_10555;
assign v_10557 = v_6756 & v_6764;
assign v_10559 = v_6592 & v_10558;
assign v_10560 = v_6607 & v_6614;
assign v_10562 = v_6441 & v_10561;
assign v_10563 = v_6472 & v_6482;
assign v_10565 = v_6296 & v_10564;
assign v_10566 = v_6311 & v_6318;
assign v_10568 = v_6153 & v_10567;
assign v_10569 = v_6178 & v_6186;
assign v_10571 = v_6012 & v_10570;
assign v_10572 = v_6027 & v_6034;
assign v_10574 = v_5866 & v_10573;
assign v_10575 = v_5893 & v_5902;
assign v_10577 = v_5724 & v_10576;
assign v_10578 = v_5739 & v_5746;
assign v_10580 = v_5582 & v_10579;
assign v_10581 = v_5606 & v_5614;
assign v_10583 = v_5442 & v_10582;
assign v_10584 = v_5457 & v_5464;
assign v_10586 = v_5281 & v_10585;
assign v_10587 = v_5320 & v_5332;
assign v_10589 = v_5130 & v_10588;
assign v_10590 = v_5145 & v_5152;
assign v_10592 = v_4985 & v_10591;
assign v_10593 = v_5012 & v_5020;
assign v_10595 = v_4842 & v_10594;
assign v_10596 = v_4857 & v_4864;
assign v_10598 = v_4696 & v_10597;
assign v_10599 = v_4723 & v_4732;
assign v_10601 = v_4554 & v_10600;
assign v_10602 = v_4569 & v_4576;
assign v_10604 = v_4412 & v_10603;
assign v_10605 = v_4436 & v_4444;
assign v_10607 = v_4272 & v_10606;
assign v_10608 = v_4287 & v_4294;
assign v_10610 = v_4121 & v_10609;
assign v_10611 = v_4152 & v_4162;
assign v_10613 = v_3976 & v_10612;
assign v_10614 = v_3991 & v_3998;
assign v_10616 = v_3833 & v_10615;
assign v_10617 = v_3858 & v_3866;
assign v_10619 = v_3692 & v_10618;
assign v_10620 = v_3707 & v_3714;
assign v_10622 = v_3546 & v_10621;
assign v_10623 = v_3573 & v_3582;
assign v_10625 = v_3404 & v_10624;
assign v_10626 = v_3419 & v_3426;
assign v_10628 = v_3262 & v_10627;
assign v_10629 = v_3286 & v_3294;
assign v_10631 = v_3122 & v_10630;
assign v_10632 = v_3137 & v_3144;
assign v_10634 = v_2966 & v_10633;
assign v_10635 = v_3001 & v_3012;
assign v_10637 = v_2818 & v_10636;
assign v_10638 = v_2833 & v_2840;
assign v_10640 = v_2674 & v_10639;
assign v_10641 = v_2700 & v_2708;
assign v_10643 = v_2532 & v_10642;
assign v_10644 = v_2547 & v_2554;
assign v_10646 = v_2386 & v_10645;
assign v_10647 = v_2413 & v_2422;
assign v_10649 = v_2244 & v_10648;
assign v_10650 = v_2259 & v_2266;
assign v_10652 = v_2102 & v_10651;
assign v_10653 = v_2126 & v_2134;
assign v_10655 = v_1962 & v_10654;
assign v_10656 = v_1977 & v_1984;
assign v_10658 = v_1811 & v_10657;
assign v_10659 = v_1842 & v_1852;
assign v_10661 = v_1666 & v_10660;
assign v_10662 = v_1681 & v_1688;
assign v_10664 = v_1523 & v_10663;
assign v_10665 = v_1548 & v_1556;
assign v_10667 = v_1382 & v_10666;
assign v_10668 = v_1397 & v_1404;
assign v_10670 = v_1236 & v_10669;
assign v_10671 = v_1263 & v_1272;
assign v_10673 = v_1094 & v_10672;
assign v_10674 = v_1109 & v_1116;
assign v_10676 = v_952 & v_10675;
assign v_10677 = v_976 & v_984;
assign v_10679 = v_815 & v_10678;
assign v_10680 = v_831 & v_838;
assign v_10682 = v_453 & v_10681;
assign v_10683 = v_687 & v_721;
assign v_10685 = v_9616 & v_9753;
assign v_10686 = v_9604 & v_9644;
assign v_10688 = v_9472 & v_10687;
assign v_10689 = v_9463 & v_9487;
assign v_10691 = v_9326 & v_10690;
assign v_10692 = v_9311 & v_9353;
assign v_10694 = v_9184 & v_10693;
assign v_10695 = v_9175 & v_9199;
assign v_10697 = v_9042 & v_10696;
assign v_10698 = v_9030 & v_9066;
assign v_10700 = v_8902 & v_10699;
assign v_10701 = v_8893 & v_8917;
assign v_10703 = v_8751 & v_10702;
assign v_10704 = v_8733 & v_8782;
assign v_10706 = v_8606 & v_10705;
assign v_10707 = v_8597 & v_8621;
assign v_10709 = v_8463 & v_10708;
assign v_10710 = v_8451 & v_8488;
assign v_10712 = v_8322 & v_10711;
assign v_10713 = v_8313 & v_8337;
assign v_10715 = v_8176 & v_10714;
assign v_10716 = v_8161 & v_8203;
assign v_10718 = v_8034 & v_10717;
assign v_10719 = v_8025 & v_8049;
assign v_10721 = v_7892 & v_10720;
assign v_10722 = v_7880 & v_7916;
assign v_10724 = v_7752 & v_10723;
assign v_10725 = v_7743 & v_7767;
assign v_10727 = v_7596 & v_10726;
assign v_10728 = v_7575 & v_7631;
assign v_10730 = v_7448 & v_10729;
assign v_10731 = v_7439 & v_7463;
assign v_10733 = v_7304 & v_10732;
assign v_10734 = v_7292 & v_7330;
assign v_10736 = v_7162 & v_10735;
assign v_10737 = v_7153 & v_7177;
assign v_10739 = v_7016 & v_10738;
assign v_10740 = v_7001 & v_7043;
assign v_10742 = v_6874 & v_10741;
assign v_10743 = v_6865 & v_6889;
assign v_10745 = v_6732 & v_10744;
assign v_10746 = v_6720 & v_6756;
assign v_10748 = v_6592 & v_10747;
assign v_10749 = v_6583 & v_6607;
assign v_10751 = v_6441 & v_10750;
assign v_10752 = v_6423 & v_6472;
assign v_10754 = v_6296 & v_10753;
assign v_10755 = v_6287 & v_6311;
assign v_10757 = v_6153 & v_10756;
assign v_10758 = v_6141 & v_6178;
assign v_10760 = v_6012 & v_10759;
assign v_10761 = v_6003 & v_6027;
assign v_10763 = v_5866 & v_10762;
assign v_10764 = v_5851 & v_5893;
assign v_10766 = v_5724 & v_10765;
assign v_10767 = v_5715 & v_5739;
assign v_10769 = v_5582 & v_10768;
assign v_10770 = v_5570 & v_5606;
assign v_10772 = v_5442 & v_10771;
assign v_10773 = v_5433 & v_5457;
assign v_10775 = v_5281 & v_10774;
assign v_10776 = v_5257 & v_5320;
assign v_10778 = v_5130 & v_10777;
assign v_10779 = v_5121 & v_5145;
assign v_10781 = v_4985 & v_10780;
assign v_10782 = v_4973 & v_5012;
assign v_10784 = v_4842 & v_10783;
assign v_10785 = v_4833 & v_4857;
assign v_10787 = v_4696 & v_10786;
assign v_10788 = v_4681 & v_4723;
assign v_10790 = v_4554 & v_10789;
assign v_10791 = v_4545 & v_4569;
assign v_10793 = v_4412 & v_10792;
assign v_10794 = v_4400 & v_4436;
assign v_10796 = v_4272 & v_10795;
assign v_10797 = v_4263 & v_4287;
assign v_10799 = v_4121 & v_10798;
assign v_10800 = v_4103 & v_4152;
assign v_10802 = v_3976 & v_10801;
assign v_10803 = v_3967 & v_3991;
assign v_10805 = v_3833 & v_10804;
assign v_10806 = v_3821 & v_3858;
assign v_10808 = v_3692 & v_10807;
assign v_10809 = v_3683 & v_3707;
assign v_10811 = v_3546 & v_10810;
assign v_10812 = v_3531 & v_3573;
assign v_10814 = v_3404 & v_10813;
assign v_10815 = v_3395 & v_3419;
assign v_10817 = v_3262 & v_10816;
assign v_10818 = v_3250 & v_3286;
assign v_10820 = v_3122 & v_10819;
assign v_10821 = v_3113 & v_3137;
assign v_10823 = v_2966 & v_10822;
assign v_10824 = v_2945 & v_3001;
assign v_10826 = v_2818 & v_10825;
assign v_10827 = v_2809 & v_2833;
assign v_10829 = v_2674 & v_10828;
assign v_10830 = v_2662 & v_2700;
assign v_10832 = v_2532 & v_10831;
assign v_10833 = v_2523 & v_2547;
assign v_10835 = v_2386 & v_10834;
assign v_10836 = v_2371 & v_2413;
assign v_10838 = v_2244 & v_10837;
assign v_10839 = v_2235 & v_2259;
assign v_10841 = v_2102 & v_10840;
assign v_10842 = v_2090 & v_2126;
assign v_10844 = v_1962 & v_10843;
assign v_10845 = v_1953 & v_1977;
assign v_10847 = v_1811 & v_10846;
assign v_10848 = v_1793 & v_1842;
assign v_10850 = v_1666 & v_10849;
assign v_10851 = v_1657 & v_1681;
assign v_10853 = v_1523 & v_10852;
assign v_10854 = v_1511 & v_1548;
assign v_10856 = v_1382 & v_10855;
assign v_10857 = v_1373 & v_1397;
assign v_10859 = v_1236 & v_10858;
assign v_10860 = v_1221 & v_1263;
assign v_10862 = v_1094 & v_10861;
assign v_10863 = v_1085 & v_1109;
assign v_10865 = v_952 & v_10864;
assign v_10866 = v_940 & v_976;
assign v_10868 = v_815 & v_10867;
assign v_10869 = v_804 & v_831;
assign v_10871 = v_453 & v_10870;
assign v_10872 = v_98 & v_687;
assign v_10875 = v_9616 & v_9796;
assign v_10876 = v_9644 & v_9664;
assign v_10878 = v_9472 & v_10877;
assign v_10879 = v_9487 & v_9506;
assign v_10881 = v_9326 & v_10880;
assign v_10882 = v_9353 & v_9374;
assign v_10884 = v_9184 & v_10883;
assign v_10885 = v_9199 & v_9218;
assign v_10887 = v_9042 & v_10886;
assign v_10888 = v_9066 & v_9086;
assign v_10890 = v_8902 & v_10889;
assign v_10891 = v_8917 & v_8936;
assign v_10893 = v_8751 & v_10892;
assign v_10894 = v_8782 & v_8804;
assign v_10896 = v_8606 & v_10895;
assign v_10897 = v_8621 & v_8640;
assign v_10899 = v_8463 & v_10898;
assign v_10900 = v_8488 & v_8508;
assign v_10902 = v_8322 & v_10901;
assign v_10903 = v_8337 & v_8356;
assign v_10905 = v_8176 & v_10904;
assign v_10906 = v_8203 & v_8224;
assign v_10908 = v_8034 & v_10907;
assign v_10909 = v_8049 & v_8068;
assign v_10911 = v_7892 & v_10910;
assign v_10912 = v_7916 & v_7936;
assign v_10914 = v_7752 & v_10913;
assign v_10915 = v_7767 & v_7786;
assign v_10917 = v_7596 & v_10916;
assign v_10918 = v_7631 & v_7654;
assign v_10920 = v_7448 & v_10919;
assign v_10921 = v_7463 & v_7482;
assign v_10923 = v_7304 & v_10922;
assign v_10924 = v_7330 & v_7350;
assign v_10926 = v_7162 & v_10925;
assign v_10927 = v_7177 & v_7196;
assign v_10929 = v_7016 & v_10928;
assign v_10930 = v_7043 & v_7064;
assign v_10932 = v_6874 & v_10931;
assign v_10933 = v_6889 & v_6908;
assign v_10935 = v_6732 & v_10934;
assign v_10936 = v_6756 & v_6776;
assign v_10938 = v_6592 & v_10937;
assign v_10939 = v_6607 & v_6626;
assign v_10941 = v_6441 & v_10940;
assign v_10942 = v_6472 & v_6494;
assign v_10944 = v_6296 & v_10943;
assign v_10945 = v_6311 & v_6330;
assign v_10947 = v_6153 & v_10946;
assign v_10948 = v_6178 & v_6198;
assign v_10950 = v_6012 & v_10949;
assign v_10951 = v_6027 & v_6046;
assign v_10953 = v_5866 & v_10952;
assign v_10954 = v_5893 & v_5914;
assign v_10956 = v_5724 & v_10955;
assign v_10957 = v_5739 & v_5758;
assign v_10959 = v_5582 & v_10958;
assign v_10960 = v_5606 & v_5626;
assign v_10962 = v_5442 & v_10961;
assign v_10963 = v_5457 & v_5476;
assign v_10965 = v_5281 & v_10964;
assign v_10966 = v_5320 & v_5344;
assign v_10968 = v_5130 & v_10967;
assign v_10969 = v_5145 & v_5164;
assign v_10971 = v_4985 & v_10970;
assign v_10972 = v_5012 & v_5032;
assign v_10974 = v_4842 & v_10973;
assign v_10975 = v_4857 & v_4876;
assign v_10977 = v_4696 & v_10976;
assign v_10978 = v_4723 & v_4744;
assign v_10980 = v_4554 & v_10979;
assign v_10981 = v_4569 & v_4588;
assign v_10983 = v_4412 & v_10982;
assign v_10984 = v_4436 & v_4456;
assign v_10986 = v_4272 & v_10985;
assign v_10987 = v_4287 & v_4306;
assign v_10989 = v_4121 & v_10988;
assign v_10990 = v_4152 & v_4174;
assign v_10992 = v_3976 & v_10991;
assign v_10993 = v_3991 & v_4010;
assign v_10995 = v_3833 & v_10994;
assign v_10996 = v_3858 & v_3878;
assign v_10998 = v_3692 & v_10997;
assign v_10999 = v_3707 & v_3726;
assign v_11001 = v_3546 & v_11000;
assign v_11002 = v_3573 & v_3594;
assign v_11004 = v_3404 & v_11003;
assign v_11005 = v_3419 & v_3438;
assign v_11007 = v_3262 & v_11006;
assign v_11008 = v_3286 & v_3306;
assign v_11010 = v_3122 & v_11009;
assign v_11011 = v_3137 & v_3156;
assign v_11013 = v_2966 & v_11012;
assign v_11014 = v_3001 & v_3024;
assign v_11016 = v_2818 & v_11015;
assign v_11017 = v_2833 & v_2852;
assign v_11019 = v_2674 & v_11018;
assign v_11020 = v_2700 & v_2720;
assign v_11022 = v_2532 & v_11021;
assign v_11023 = v_2547 & v_2566;
assign v_11025 = v_2386 & v_11024;
assign v_11026 = v_2413 & v_2434;
assign v_11028 = v_2244 & v_11027;
assign v_11029 = v_2259 & v_2278;
assign v_11031 = v_2102 & v_11030;
assign v_11032 = v_2126 & v_2146;
assign v_11034 = v_1962 & v_11033;
assign v_11035 = v_1977 & v_1996;
assign v_11037 = v_1811 & v_11036;
assign v_11038 = v_1842 & v_1864;
assign v_11040 = v_1666 & v_11039;
assign v_11041 = v_1681 & v_1700;
assign v_11043 = v_1523 & v_11042;
assign v_11044 = v_1548 & v_1568;
assign v_11046 = v_1382 & v_11045;
assign v_11047 = v_1397 & v_1416;
assign v_11049 = v_1236 & v_11048;
assign v_11050 = v_1263 & v_1284;
assign v_11052 = v_1094 & v_11051;
assign v_11053 = v_1109 & v_1128;
assign v_11055 = v_952 & v_11054;
assign v_11056 = v_976 & v_996;
assign v_11058 = v_815 & v_11057;
assign v_11059 = v_831 & v_850;
assign v_11061 = v_453 & v_11060;
assign v_11062 = v_687 & v_731;
assign v_11065 = v_9616 & v_9808;
assign v_11066 = v_9644 & v_9676;
assign v_11068 = v_9472 & v_11067;
assign v_11069 = v_9487 & v_9518;
assign v_11071 = v_9326 & v_11070;
assign v_11072 = v_9353 & v_9386;
assign v_11074 = v_9184 & v_11073;
assign v_11075 = v_9199 & v_9230;
assign v_11077 = v_9042 & v_11076;
assign v_11078 = v_9066 & v_9098;
assign v_11080 = v_8902 & v_11079;
assign v_11081 = v_8917 & v_8948;
assign v_11083 = v_8751 & v_11082;
assign v_11084 = v_8782 & v_8816;
assign v_11086 = v_8606 & v_11085;
assign v_11087 = v_8621 & v_8652;
assign v_11089 = v_8463 & v_11088;
assign v_11090 = v_8488 & v_8520;
assign v_11092 = v_8322 & v_11091;
assign v_11093 = v_8337 & v_8368;
assign v_11095 = v_8176 & v_11094;
assign v_11096 = v_8203 & v_8236;
assign v_11098 = v_8034 & v_11097;
assign v_11099 = v_8049 & v_8080;
assign v_11101 = v_7892 & v_11100;
assign v_11102 = v_7916 & v_7948;
assign v_11104 = v_7752 & v_11103;
assign v_11105 = v_7767 & v_7798;
assign v_11107 = v_7596 & v_11106;
assign v_11108 = v_7631 & v_7666;
assign v_11110 = v_7448 & v_11109;
assign v_11111 = v_7463 & v_7494;
assign v_11113 = v_7304 & v_11112;
assign v_11114 = v_7330 & v_7362;
assign v_11116 = v_7162 & v_11115;
assign v_11117 = v_7177 & v_7208;
assign v_11119 = v_7016 & v_11118;
assign v_11120 = v_7043 & v_7076;
assign v_11122 = v_6874 & v_11121;
assign v_11123 = v_6889 & v_6920;
assign v_11125 = v_6732 & v_11124;
assign v_11126 = v_6756 & v_6788;
assign v_11128 = v_6592 & v_11127;
assign v_11129 = v_6607 & v_6638;
assign v_11131 = v_6441 & v_11130;
assign v_11132 = v_6472 & v_6506;
assign v_11134 = v_6296 & v_11133;
assign v_11135 = v_6311 & v_6342;
assign v_11137 = v_6153 & v_11136;
assign v_11138 = v_6178 & v_6210;
assign v_11140 = v_6012 & v_11139;
assign v_11141 = v_6027 & v_6058;
assign v_11143 = v_5866 & v_11142;
assign v_11144 = v_5893 & v_5926;
assign v_11146 = v_5724 & v_11145;
assign v_11147 = v_5739 & v_5770;
assign v_11149 = v_5582 & v_11148;
assign v_11150 = v_5606 & v_5638;
assign v_11152 = v_5442 & v_11151;
assign v_11153 = v_5457 & v_5488;
assign v_11155 = v_5281 & v_11154;
assign v_11156 = v_5320 & v_5356;
assign v_11158 = v_5130 & v_11157;
assign v_11159 = v_5145 & v_5176;
assign v_11161 = v_4985 & v_11160;
assign v_11162 = v_5012 & v_5044;
assign v_11164 = v_4842 & v_11163;
assign v_11165 = v_4857 & v_4888;
assign v_11167 = v_4696 & v_11166;
assign v_11168 = v_4723 & v_4756;
assign v_11170 = v_4554 & v_11169;
assign v_11171 = v_4569 & v_4600;
assign v_11173 = v_4412 & v_11172;
assign v_11174 = v_4436 & v_4468;
assign v_11176 = v_4272 & v_11175;
assign v_11177 = v_4287 & v_4318;
assign v_11179 = v_4121 & v_11178;
assign v_11180 = v_4152 & v_4186;
assign v_11182 = v_3976 & v_11181;
assign v_11183 = v_3991 & v_4022;
assign v_11185 = v_3833 & v_11184;
assign v_11186 = v_3858 & v_3890;
assign v_11188 = v_3692 & v_11187;
assign v_11189 = v_3707 & v_3738;
assign v_11191 = v_3546 & v_11190;
assign v_11192 = v_3573 & v_3606;
assign v_11194 = v_3404 & v_11193;
assign v_11195 = v_3419 & v_3450;
assign v_11197 = v_3262 & v_11196;
assign v_11198 = v_3286 & v_3318;
assign v_11200 = v_3122 & v_11199;
assign v_11201 = v_3137 & v_3168;
assign v_11203 = v_2966 & v_11202;
assign v_11204 = v_3001 & v_3036;
assign v_11206 = v_2818 & v_11205;
assign v_11207 = v_2833 & v_2864;
assign v_11209 = v_2674 & v_11208;
assign v_11210 = v_2700 & v_2732;
assign v_11212 = v_2532 & v_11211;
assign v_11213 = v_2547 & v_2578;
assign v_11215 = v_2386 & v_11214;
assign v_11216 = v_2413 & v_2446;
assign v_11218 = v_2244 & v_11217;
assign v_11219 = v_2259 & v_2290;
assign v_11221 = v_2102 & v_11220;
assign v_11222 = v_2126 & v_2158;
assign v_11224 = v_1962 & v_11223;
assign v_11225 = v_1977 & v_2008;
assign v_11227 = v_1811 & v_11226;
assign v_11228 = v_1842 & v_1876;
assign v_11230 = v_1666 & v_11229;
assign v_11231 = v_1681 & v_1712;
assign v_11233 = v_1523 & v_11232;
assign v_11234 = v_1548 & v_1580;
assign v_11236 = v_1382 & v_11235;
assign v_11237 = v_1397 & v_1428;
assign v_11239 = v_1236 & v_11238;
assign v_11240 = v_1263 & v_1296;
assign v_11242 = v_1094 & v_11241;
assign v_11243 = v_1109 & v_1140;
assign v_11245 = v_952 & v_11244;
assign v_11246 = v_976 & v_1008;
assign v_11248 = v_815 & v_11247;
assign v_11249 = v_831 & v_862;
assign v_11251 = v_453 & v_11250;
assign v_11252 = v_687 & v_741;
assign v_11255 = v_9616 & v_9820;
assign v_11256 = v_9644 & v_9688;
assign v_11258 = v_9472 & v_11257;
assign v_11259 = v_9487 & v_9530;
assign v_11261 = v_9326 & v_11260;
assign v_11262 = v_9353 & v_9398;
assign v_11264 = v_9184 & v_11263;
assign v_11265 = v_9199 & v_9242;
assign v_11267 = v_9042 & v_11266;
assign v_11268 = v_9066 & v_9110;
assign v_11270 = v_8902 & v_11269;
assign v_11271 = v_8917 & v_8960;
assign v_11273 = v_8751 & v_11272;
assign v_11274 = v_8782 & v_8828;
assign v_11276 = v_8606 & v_11275;
assign v_11277 = v_8621 & v_8664;
assign v_11279 = v_8463 & v_11278;
assign v_11280 = v_8488 & v_8532;
assign v_11282 = v_8322 & v_11281;
assign v_11283 = v_8337 & v_8380;
assign v_11285 = v_8176 & v_11284;
assign v_11286 = v_8203 & v_8248;
assign v_11288 = v_8034 & v_11287;
assign v_11289 = v_8049 & v_8092;
assign v_11291 = v_7892 & v_11290;
assign v_11292 = v_7916 & v_7960;
assign v_11294 = v_7752 & v_11293;
assign v_11295 = v_7767 & v_7810;
assign v_11297 = v_7596 & v_11296;
assign v_11298 = v_7631 & v_7678;
assign v_11300 = v_7448 & v_11299;
assign v_11301 = v_7463 & v_7506;
assign v_11303 = v_7304 & v_11302;
assign v_11304 = v_7330 & v_7374;
assign v_11306 = v_7162 & v_11305;
assign v_11307 = v_7177 & v_7220;
assign v_11309 = v_7016 & v_11308;
assign v_11310 = v_7043 & v_7088;
assign v_11312 = v_6874 & v_11311;
assign v_11313 = v_6889 & v_6932;
assign v_11315 = v_6732 & v_11314;
assign v_11316 = v_6756 & v_6800;
assign v_11318 = v_6592 & v_11317;
assign v_11319 = v_6607 & v_6650;
assign v_11321 = v_6441 & v_11320;
assign v_11322 = v_6472 & v_6518;
assign v_11324 = v_6296 & v_11323;
assign v_11325 = v_6311 & v_6354;
assign v_11327 = v_6153 & v_11326;
assign v_11328 = v_6178 & v_6222;
assign v_11330 = v_6012 & v_11329;
assign v_11331 = v_6027 & v_6070;
assign v_11333 = v_5866 & v_11332;
assign v_11334 = v_5893 & v_5938;
assign v_11336 = v_5724 & v_11335;
assign v_11337 = v_5739 & v_5782;
assign v_11339 = v_5582 & v_11338;
assign v_11340 = v_5606 & v_5650;
assign v_11342 = v_5442 & v_11341;
assign v_11343 = v_5457 & v_5500;
assign v_11345 = v_5281 & v_11344;
assign v_11346 = v_5320 & v_5368;
assign v_11348 = v_5130 & v_11347;
assign v_11349 = v_5145 & v_5188;
assign v_11351 = v_4985 & v_11350;
assign v_11352 = v_5012 & v_5056;
assign v_11354 = v_4842 & v_11353;
assign v_11355 = v_4857 & v_4900;
assign v_11357 = v_4696 & v_11356;
assign v_11358 = v_4723 & v_4768;
assign v_11360 = v_4554 & v_11359;
assign v_11361 = v_4569 & v_4612;
assign v_11363 = v_4412 & v_11362;
assign v_11364 = v_4436 & v_4480;
assign v_11366 = v_4272 & v_11365;
assign v_11367 = v_4287 & v_4330;
assign v_11369 = v_4121 & v_11368;
assign v_11370 = v_4152 & v_4198;
assign v_11372 = v_3976 & v_11371;
assign v_11373 = v_3991 & v_4034;
assign v_11375 = v_3833 & v_11374;
assign v_11376 = v_3858 & v_3902;
assign v_11378 = v_3692 & v_11377;
assign v_11379 = v_3707 & v_3750;
assign v_11381 = v_3546 & v_11380;
assign v_11382 = v_3573 & v_3618;
assign v_11384 = v_3404 & v_11383;
assign v_11385 = v_3419 & v_3462;
assign v_11387 = v_3262 & v_11386;
assign v_11388 = v_3286 & v_3330;
assign v_11390 = v_3122 & v_11389;
assign v_11391 = v_3137 & v_3180;
assign v_11393 = v_2966 & v_11392;
assign v_11394 = v_3001 & v_3048;
assign v_11396 = v_2818 & v_11395;
assign v_11397 = v_2833 & v_2876;
assign v_11399 = v_2674 & v_11398;
assign v_11400 = v_2700 & v_2744;
assign v_11402 = v_2532 & v_11401;
assign v_11403 = v_2547 & v_2590;
assign v_11405 = v_2386 & v_11404;
assign v_11406 = v_2413 & v_2458;
assign v_11408 = v_2244 & v_11407;
assign v_11409 = v_2259 & v_2302;
assign v_11411 = v_2102 & v_11410;
assign v_11412 = v_2126 & v_2170;
assign v_11414 = v_1962 & v_11413;
assign v_11415 = v_1977 & v_2020;
assign v_11417 = v_1811 & v_11416;
assign v_11418 = v_1842 & v_1888;
assign v_11420 = v_1666 & v_11419;
assign v_11421 = v_1681 & v_1724;
assign v_11423 = v_1523 & v_11422;
assign v_11424 = v_1548 & v_1592;
assign v_11426 = v_1382 & v_11425;
assign v_11427 = v_1397 & v_1440;
assign v_11429 = v_1236 & v_11428;
assign v_11430 = v_1263 & v_1308;
assign v_11432 = v_1094 & v_11431;
assign v_11433 = v_1109 & v_1152;
assign v_11435 = v_952 & v_11434;
assign v_11436 = v_976 & v_1020;
assign v_11438 = v_815 & v_11437;
assign v_11439 = v_831 & v_874;
assign v_11441 = v_453 & v_11440;
assign v_11442 = v_687 & v_751;
assign v_11445 = v_9616 & v_9832;
assign v_11446 = v_9644 & v_9700;
assign v_11448 = v_9472 & v_11447;
assign v_11449 = v_9487 & v_9542;
assign v_11451 = v_9326 & v_11450;
assign v_11452 = v_9353 & v_9410;
assign v_11454 = v_9184 & v_11453;
assign v_11455 = v_9199 & v_9254;
assign v_11457 = v_9042 & v_11456;
assign v_11458 = v_9066 & v_9122;
assign v_11460 = v_8902 & v_11459;
assign v_11461 = v_8917 & v_8972;
assign v_11463 = v_8751 & v_11462;
assign v_11464 = v_8782 & v_8840;
assign v_11466 = v_8606 & v_11465;
assign v_11467 = v_8621 & v_8676;
assign v_11469 = v_8463 & v_11468;
assign v_11470 = v_8488 & v_8544;
assign v_11472 = v_8322 & v_11471;
assign v_11473 = v_8337 & v_8392;
assign v_11475 = v_8176 & v_11474;
assign v_11476 = v_8203 & v_8260;
assign v_11478 = v_8034 & v_11477;
assign v_11479 = v_8049 & v_8104;
assign v_11481 = v_7892 & v_11480;
assign v_11482 = v_7916 & v_7972;
assign v_11484 = v_7752 & v_11483;
assign v_11485 = v_7767 & v_7822;
assign v_11487 = v_7596 & v_11486;
assign v_11488 = v_7631 & v_7690;
assign v_11490 = v_7448 & v_11489;
assign v_11491 = v_7463 & v_7518;
assign v_11493 = v_7304 & v_11492;
assign v_11494 = v_7330 & v_7386;
assign v_11496 = v_7162 & v_11495;
assign v_11497 = v_7177 & v_7232;
assign v_11499 = v_7016 & v_11498;
assign v_11500 = v_7043 & v_7100;
assign v_11502 = v_6874 & v_11501;
assign v_11503 = v_6889 & v_6944;
assign v_11505 = v_6732 & v_11504;
assign v_11506 = v_6756 & v_6812;
assign v_11508 = v_6592 & v_11507;
assign v_11509 = v_6607 & v_6662;
assign v_11511 = v_6441 & v_11510;
assign v_11512 = v_6472 & v_6530;
assign v_11514 = v_6296 & v_11513;
assign v_11515 = v_6311 & v_6366;
assign v_11517 = v_6153 & v_11516;
assign v_11518 = v_6178 & v_6234;
assign v_11520 = v_6012 & v_11519;
assign v_11521 = v_6027 & v_6082;
assign v_11523 = v_5866 & v_11522;
assign v_11524 = v_5893 & v_5950;
assign v_11526 = v_5724 & v_11525;
assign v_11527 = v_5739 & v_5794;
assign v_11529 = v_5582 & v_11528;
assign v_11530 = v_5606 & v_5662;
assign v_11532 = v_5442 & v_11531;
assign v_11533 = v_5457 & v_5512;
assign v_11535 = v_5281 & v_11534;
assign v_11536 = v_5320 & v_5380;
assign v_11538 = v_5130 & v_11537;
assign v_11539 = v_5145 & v_5200;
assign v_11541 = v_4985 & v_11540;
assign v_11542 = v_5012 & v_5068;
assign v_11544 = v_4842 & v_11543;
assign v_11545 = v_4857 & v_4912;
assign v_11547 = v_4696 & v_11546;
assign v_11548 = v_4723 & v_4780;
assign v_11550 = v_4554 & v_11549;
assign v_11551 = v_4569 & v_4624;
assign v_11553 = v_4412 & v_11552;
assign v_11554 = v_4436 & v_4492;
assign v_11556 = v_4272 & v_11555;
assign v_11557 = v_4287 & v_4342;
assign v_11559 = v_4121 & v_11558;
assign v_11560 = v_4152 & v_4210;
assign v_11562 = v_3976 & v_11561;
assign v_11563 = v_3991 & v_4046;
assign v_11565 = v_3833 & v_11564;
assign v_11566 = v_3858 & v_3914;
assign v_11568 = v_3692 & v_11567;
assign v_11569 = v_3707 & v_3762;
assign v_11571 = v_3546 & v_11570;
assign v_11572 = v_3573 & v_3630;
assign v_11574 = v_3404 & v_11573;
assign v_11575 = v_3419 & v_3474;
assign v_11577 = v_3262 & v_11576;
assign v_11578 = v_3286 & v_3342;
assign v_11580 = v_3122 & v_11579;
assign v_11581 = v_3137 & v_3192;
assign v_11583 = v_2966 & v_11582;
assign v_11584 = v_3001 & v_3060;
assign v_11586 = v_2818 & v_11585;
assign v_11587 = v_2833 & v_2888;
assign v_11589 = v_2674 & v_11588;
assign v_11590 = v_2700 & v_2756;
assign v_11592 = v_2532 & v_11591;
assign v_11593 = v_2547 & v_2602;
assign v_11595 = v_2386 & v_11594;
assign v_11596 = v_2413 & v_2470;
assign v_11598 = v_2244 & v_11597;
assign v_11599 = v_2259 & v_2314;
assign v_11601 = v_2102 & v_11600;
assign v_11602 = v_2126 & v_2182;
assign v_11604 = v_1962 & v_11603;
assign v_11605 = v_1977 & v_2032;
assign v_11607 = v_1811 & v_11606;
assign v_11608 = v_1842 & v_1900;
assign v_11610 = v_1666 & v_11609;
assign v_11611 = v_1681 & v_1736;
assign v_11613 = v_1523 & v_11612;
assign v_11614 = v_1548 & v_1604;
assign v_11616 = v_1382 & v_11615;
assign v_11617 = v_1397 & v_1452;
assign v_11619 = v_1236 & v_11618;
assign v_11620 = v_1263 & v_1320;
assign v_11622 = v_1094 & v_11621;
assign v_11623 = v_1109 & v_1164;
assign v_11625 = v_952 & v_11624;
assign v_11626 = v_976 & v_1032;
assign v_11628 = v_815 & v_11627;
assign v_11629 = v_831 & v_886;
assign v_11631 = v_453 & v_11630;
assign v_11632 = v_687 & v_761;
assign v_11635 = v_9616 & v_9844;
assign v_11636 = v_9644 & v_9712;
assign v_11638 = v_9472 & v_11637;
assign v_11639 = v_9487 & v_9554;
assign v_11641 = v_9326 & v_11640;
assign v_11642 = v_9353 & v_9422;
assign v_11644 = v_9184 & v_11643;
assign v_11645 = v_9199 & v_9266;
assign v_11647 = v_9042 & v_11646;
assign v_11648 = v_9066 & v_9134;
assign v_11650 = v_8902 & v_11649;
assign v_11651 = v_8917 & v_8984;
assign v_11653 = v_8751 & v_11652;
assign v_11654 = v_8782 & v_8852;
assign v_11656 = v_8606 & v_11655;
assign v_11657 = v_8621 & v_8688;
assign v_11659 = v_8463 & v_11658;
assign v_11660 = v_8488 & v_8556;
assign v_11662 = v_8322 & v_11661;
assign v_11663 = v_8337 & v_8404;
assign v_11665 = v_8176 & v_11664;
assign v_11666 = v_8203 & v_8272;
assign v_11668 = v_8034 & v_11667;
assign v_11669 = v_8049 & v_8116;
assign v_11671 = v_7892 & v_11670;
assign v_11672 = v_7916 & v_7984;
assign v_11674 = v_7752 & v_11673;
assign v_11675 = v_7767 & v_7834;
assign v_11677 = v_7596 & v_11676;
assign v_11678 = v_7631 & v_7702;
assign v_11680 = v_7448 & v_11679;
assign v_11681 = v_7463 & v_7530;
assign v_11683 = v_7304 & v_11682;
assign v_11684 = v_7330 & v_7398;
assign v_11686 = v_7162 & v_11685;
assign v_11687 = v_7177 & v_7244;
assign v_11689 = v_7016 & v_11688;
assign v_11690 = v_7043 & v_7112;
assign v_11692 = v_6874 & v_11691;
assign v_11693 = v_6889 & v_6956;
assign v_11695 = v_6732 & v_11694;
assign v_11696 = v_6756 & ~v_6824;
assign v_11698 = v_6592 & v_11697;
assign v_11699 = v_6607 & v_6674;
assign v_11701 = v_6441 & v_11700;
assign v_11702 = v_6472 & v_6542;
assign v_11704 = v_6296 & v_11703;
assign v_11705 = v_6311 & v_6378;
assign v_11707 = v_6153 & v_11706;
assign v_11708 = v_6178 & v_6246;
assign v_11710 = v_6012 & v_11709;
assign v_11711 = v_6027 & ~v_6094;
assign v_11713 = v_5866 & v_11712;
assign v_11714 = v_5893 & v_5962;
assign v_11716 = v_5724 & v_11715;
assign v_11717 = v_5739 & ~v_5806;
assign v_11719 = v_5582 & v_11718;
assign v_11720 = v_5606 & v_5674;
assign v_11722 = v_5442 & v_11721;
assign v_11723 = v_5457 & v_5524;
assign v_11725 = v_5281 & v_11724;
assign v_11726 = v_5320 & v_5392;
assign v_11728 = v_5130 & v_11727;
assign v_11729 = v_5145 & v_5212;
assign v_11731 = v_4985 & v_11730;
assign v_11732 = v_5012 & v_5080;
assign v_11734 = v_4842 & v_11733;
assign v_11735 = v_4857 & v_4924;
assign v_11737 = v_4696 & v_11736;
assign v_11738 = v_4723 & v_4792;
assign v_11740 = v_4554 & v_11739;
assign v_11741 = v_4569 & v_4636;
assign v_11743 = v_4412 & v_11742;
assign v_11744 = v_4436 & v_4504;
assign v_11746 = v_4272 & v_11745;
assign v_11747 = v_4287 & v_4354;
assign v_11749 = v_4121 & v_11748;
assign v_11750 = v_4152 & v_4222;
assign v_11752 = v_3976 & v_11751;
assign v_11753 = v_3991 & v_4058;
assign v_11755 = v_3833 & v_11754;
assign v_11756 = v_3858 & v_3926;
assign v_11758 = v_3692 & v_11757;
assign v_11759 = v_3707 & v_3774;
assign v_11761 = v_3546 & v_11760;
assign v_11762 = v_3573 & v_3642;
assign v_11764 = v_3404 & v_11763;
assign v_11765 = v_3419 & v_3486;
assign v_11767 = v_3262 & v_11766;
assign v_11768 = v_3286 & v_3354;
assign v_11770 = v_3122 & v_11769;
assign v_11771 = v_3137 & ~v_3204;
assign v_11773 = v_2966 & v_11772;
assign v_11774 = v_3001 & v_3072;
assign v_11776 = v_2818 & v_11775;
assign v_11777 = v_2833 & v_2900;
assign v_11779 = v_2674 & v_11778;
assign v_11780 = v_2700 & v_2768;
assign v_11782 = v_2532 & v_11781;
assign v_11783 = v_2547 & v_2614;
assign v_11785 = v_2386 & v_11784;
assign v_11786 = v_2413 & v_2482;
assign v_11788 = v_2244 & v_11787;
assign v_11789 = v_2259 & v_2326;
assign v_11791 = v_2102 & v_11790;
assign v_11792 = v_2126 & v_2194;
assign v_11794 = v_1962 & v_11793;
assign v_11795 = v_1977 & v_2044;
assign v_11797 = v_1811 & v_11796;
assign v_11798 = v_1842 & v_1912;
assign v_11800 = v_1666 & v_11799;
assign v_11801 = v_1681 & v_1748;
assign v_11803 = v_1523 & v_11802;
assign v_11804 = v_1548 & v_1616;
assign v_11806 = v_1382 & v_11805;
assign v_11807 = v_1397 & v_1464;
assign v_11809 = v_1236 & v_11808;
assign v_11810 = v_1263 & v_1332;
assign v_11812 = v_1094 & v_11811;
assign v_11813 = v_1109 & v_1176;
assign v_11815 = v_952 & v_11814;
assign v_11816 = v_976 & v_1044;
assign v_11818 = v_815 & v_11817;
assign v_11819 = v_831 & v_898;
assign v_11821 = v_453 & v_11820;
assign v_11822 = v_687 & v_771;
assign v_11825 = v_9616 & ~v_9872;
assign v_11826 = v_9644 & ~v_9740;
assign v_11828 = v_9472 & v_11827;
assign v_11829 = v_9487 & ~v_9582;
assign v_11831 = v_9326 & v_11830;
assign v_11832 = v_9353 & ~v_9450;
assign v_11834 = v_9184 & v_11833;
assign v_11835 = v_9199 & ~v_9294;
assign v_11837 = v_9042 & v_11836;
assign v_11838 = v_9066 & ~v_9162;
assign v_11840 = v_8902 & v_11839;
assign v_11841 = v_8917 & ~v_9012;
assign v_11843 = v_8751 & v_11842;
assign v_11844 = v_8782 & ~v_8880;
assign v_11846 = v_8606 & v_11845;
assign v_11847 = v_8621 & ~v_8716;
assign v_11849 = v_8463 & v_11848;
assign v_11850 = v_8488 & ~v_8584;
assign v_11852 = v_8322 & v_11851;
assign v_11853 = v_8337 & v_8432;
assign v_11855 = v_8176 & v_11854;
assign v_11856 = v_8203 & v_8300;
assign v_11858 = v_8034 & v_11857;
assign v_11859 = v_8049 & v_8144;
assign v_11861 = v_7892 & v_11860;
assign v_11862 = v_7916 & ~v_8012;
assign v_11864 = v_7752 & v_11863;
assign v_11865 = v_7767 & ~v_7862;
assign v_11867 = v_7596 & v_11866;
assign v_11868 = v_7631 & ~v_7730;
assign v_11870 = v_7448 & v_11869;
assign v_11871 = v_7463 & ~v_7558;
assign v_11873 = v_7304 & v_11872;
assign v_11874 = v_7330 & ~v_7426;
assign v_11876 = v_7162 & v_11875;
assign v_11877 = v_7177 & v_7272;
assign v_11879 = v_7016 & v_11878;
assign v_11880 = v_7043 & ~v_7140;
assign v_11882 = v_6874 & v_11881;
assign v_11883 = v_6889 & v_6984;
assign v_11885 = v_6732 & v_11884;
assign v_11886 = v_6756 & v_6852;
assign v_11888 = v_6592 & v_11887;
assign v_11889 = v_6607 & v_6702;
assign v_11891 = v_6441 & v_11890;
assign v_11892 = v_6472 & ~v_6570;
assign v_11894 = v_6296 & v_11893;
assign v_11895 = v_6311 & ~v_6406;
assign v_11897 = v_6153 & v_11896;
assign v_11898 = v_6178 & v_6274;
assign v_11900 = v_6012 & v_11899;
assign v_11901 = v_6027 & v_6122;
assign v_11903 = v_5866 & v_11902;
assign v_11904 = v_5893 & v_5990;
assign v_11906 = v_5724 & v_11905;
assign v_11907 = v_5739 & v_5834;
assign v_11909 = v_5582 & v_11908;
assign v_11910 = v_5606 & v_5702;
assign v_11912 = v_5442 & v_11911;
assign v_11913 = v_5457 & v_5552;
assign v_11915 = v_5281 & v_11914;
assign v_11916 = v_5320 & ~v_5420;
assign v_11918 = v_5130 & v_11917;
assign v_11919 = v_5145 & ~v_5240;
assign v_11921 = v_4985 & v_11920;
assign v_11922 = v_5012 & v_5108;
assign v_11924 = v_4842 & v_11923;
assign v_11925 = v_4857 & v_4952;
assign v_11927 = v_4696 & v_11926;
assign v_11928 = v_4723 & v_4820;
assign v_11930 = v_4554 & v_11929;
assign v_11931 = v_4569 & v_4664;
assign v_11933 = v_4412 & v_11932;
assign v_11934 = v_4436 & v_4532;
assign v_11936 = v_4272 & v_11935;
assign v_11937 = v_4287 & v_4382;
assign v_11939 = v_4121 & v_11938;
assign v_11940 = v_4152 & ~v_4250;
assign v_11942 = v_3976 & v_11941;
assign v_11943 = v_3991 & ~v_4086;
assign v_11945 = v_3833 & v_11944;
assign v_11946 = v_3858 & ~v_3954;
assign v_11948 = v_3692 & v_11947;
assign v_11949 = v_3707 & ~v_3802;
assign v_11951 = v_3546 & v_11950;
assign v_11952 = v_3573 & ~v_3670;
assign v_11954 = v_3404 & v_11953;
assign v_11955 = v_3419 & v_3514;
assign v_11957 = v_3262 & v_11956;
assign v_11958 = v_3286 & ~v_3382;
assign v_11960 = v_3122 & v_11959;
assign v_11961 = v_3137 & v_3232;
assign v_11963 = v_2966 & v_11962;
assign v_11964 = v_3001 & ~v_3100;
assign v_11966 = v_2818 & v_11965;
assign v_11967 = v_2833 & ~v_2928;
assign v_11969 = v_2674 & v_11968;
assign v_11970 = v_2700 & ~v_2796;
assign v_11972 = v_2532 & v_11971;
assign v_11973 = v_2547 & ~v_2642;
assign v_11975 = v_2386 & v_11974;
assign v_11976 = v_2413 & ~v_2510;
assign v_11978 = v_2244 & v_11977;
assign v_11979 = v_2259 & v_2354;
assign v_11981 = v_2102 & v_11980;
assign v_11982 = v_2126 & v_2222;
assign v_11984 = v_1962 & v_11983;
assign v_11985 = v_1977 & v_2072;
assign v_11987 = v_1811 & v_11986;
assign v_11988 = v_1842 & ~v_1940;
assign v_11990 = v_1666 & v_11989;
assign v_11991 = v_1681 & ~v_1776;
assign v_11993 = v_1523 & v_11992;
assign v_11994 = v_1548 & ~v_1644;
assign v_11996 = v_1382 & v_11995;
assign v_11997 = v_1397 & ~v_1492;
assign v_11999 = v_1236 & v_11998;
assign v_12000 = v_1263 & ~v_1360;
assign v_12002 = v_1094 & v_12001;
assign v_12003 = v_1109 & ~v_1204;
assign v_12005 = v_952 & v_12004;
assign v_12006 = v_976 & ~v_1072;
assign v_12008 = v_815 & v_12007;
assign v_12009 = v_831 & ~v_922;
assign v_12011 = v_453 & v_12010;
assign v_12012 = v_687 & ~v_793;
assign v_12015 = v_9618 & v_9784;
assign v_12016 = v_9646 & v_9652;
assign v_12018 = v_9473 & v_12017;
assign v_12019 = v_9488 & v_9494;
assign v_12021 = v_9329 & v_12020;
assign v_12022 = v_9356 & v_9362;
assign v_12024 = v_9185 & v_12023;
assign v_12025 = v_9200 & v_9206;
assign v_12027 = v_9044 & v_12026;
assign v_12028 = v_9068 & v_9074;
assign v_12030 = v_8903 & v_12029;
assign v_12031 = v_8918 & v_8924;
assign v_12033 = v_8755 & v_12032;
assign v_12034 = v_8786 & v_8792;
assign v_12036 = v_8607 & v_12035;
assign v_12037 = v_8622 & v_8628;
assign v_12039 = v_8465 & v_12038;
assign v_12040 = v_8490 & v_8496;
assign v_12042 = v_8323 & v_12041;
assign v_12043 = v_8338 & v_8344;
assign v_12045 = v_8179 & v_12044;
assign v_12046 = v_8206 & v_8212;
assign v_12048 = v_8035 & v_12047;
assign v_12049 = v_8050 & v_8056;
assign v_12051 = v_7894 & v_12050;
assign v_12052 = v_7918 & v_7924;
assign v_12054 = v_7753 & v_12053;
assign v_12055 = v_7768 & v_7774;
assign v_12057 = v_7601 & v_12056;
assign v_12058 = v_7636 & v_7642;
assign v_12060 = v_7449 & v_12059;
assign v_12061 = v_7464 & v_7470;
assign v_12063 = v_7306 & v_12062;
assign v_12064 = v_7332 & v_7338;
assign v_12066 = v_7163 & v_12065;
assign v_12067 = v_7178 & v_7184;
assign v_12069 = v_7019 & v_12068;
assign v_12070 = v_7046 & v_7052;
assign v_12072 = v_6875 & v_12071;
assign v_12073 = v_6890 & v_6896;
assign v_12075 = v_6734 & v_12074;
assign v_12076 = v_6758 & v_6764;
assign v_12078 = v_6593 & v_12077;
assign v_12079 = v_6608 & v_6614;
assign v_12081 = v_6445 & v_12080;
assign v_12082 = v_6476 & v_6482;
assign v_12084 = v_6297 & v_12083;
assign v_12085 = v_6312 & v_6318;
assign v_12087 = v_6155 & v_12086;
assign v_12088 = v_6180 & v_6186;
assign v_12090 = v_6013 & v_12089;
assign v_12091 = v_6028 & v_6034;
assign v_12093 = v_5869 & v_12092;
assign v_12094 = v_5896 & v_5902;
assign v_12096 = v_5725 & v_12095;
assign v_12097 = v_5740 & v_5746;
assign v_12099 = v_5584 & v_12098;
assign v_12100 = v_5608 & v_5614;
assign v_12102 = v_5443 & v_12101;
assign v_12103 = v_5458 & v_5464;
assign v_12105 = v_5287 & v_12104;
assign v_12106 = v_5326 & v_5332;
assign v_12108 = v_5131 & v_12107;
assign v_12109 = v_5146 & v_5152;
assign v_12111 = v_4987 & v_12110;
assign v_12112 = v_5014 & v_5020;
assign v_12114 = v_4843 & v_12113;
assign v_12115 = v_4858 & v_4864;
assign v_12117 = v_4699 & v_12116;
assign v_12118 = v_4726 & v_4732;
assign v_12120 = v_4555 & v_12119;
assign v_12121 = v_4570 & v_4576;
assign v_12123 = v_4414 & v_12122;
assign v_12124 = v_4438 & v_4444;
assign v_12126 = v_4273 & v_12125;
assign v_12127 = v_4288 & v_4294;
assign v_12129 = v_4125 & v_12128;
assign v_12130 = v_4156 & v_4162;
assign v_12132 = v_3977 & v_12131;
assign v_12133 = v_3992 & v_3998;
assign v_12135 = v_3835 & v_12134;
assign v_12136 = v_3860 & v_3866;
assign v_12138 = v_3693 & v_12137;
assign v_12139 = v_3708 & v_3714;
assign v_12141 = v_3549 & v_12140;
assign v_12142 = v_3576 & v_3582;
assign v_12144 = v_3405 & v_12143;
assign v_12145 = v_3420 & v_3426;
assign v_12147 = v_3264 & v_12146;
assign v_12148 = v_3288 & v_3294;
assign v_12150 = v_3123 & v_12149;
assign v_12151 = v_3138 & v_3144;
assign v_12153 = v_2971 & v_12152;
assign v_12154 = v_3006 & v_3012;
assign v_12156 = v_2819 & v_12155;
assign v_12157 = v_2834 & v_2840;
assign v_12159 = v_2676 & v_12158;
assign v_12160 = v_2702 & v_2708;
assign v_12162 = v_2533 & v_12161;
assign v_12163 = v_2548 & v_2554;
assign v_12165 = v_2389 & v_12164;
assign v_12166 = v_2416 & v_2422;
assign v_12168 = v_2245 & v_12167;
assign v_12169 = v_2260 & v_2266;
assign v_12171 = v_2104 & v_12170;
assign v_12172 = v_2128 & v_2134;
assign v_12174 = v_1963 & v_12173;
assign v_12175 = v_1978 & v_1984;
assign v_12177 = v_1815 & v_12176;
assign v_12178 = v_1846 & v_1852;
assign v_12180 = v_1667 & v_12179;
assign v_12181 = v_1682 & v_1688;
assign v_12183 = v_1525 & v_12182;
assign v_12184 = v_1550 & v_1556;
assign v_12186 = v_1383 & v_12185;
assign v_12187 = v_1398 & v_1404;
assign v_12189 = v_1239 & v_12188;
assign v_12190 = v_1266 & v_1272;
assign v_12192 = v_1095 & v_12191;
assign v_12193 = v_1110 & v_1116;
assign v_12195 = v_954 & v_12194;
assign v_12196 = v_978 & v_984;
assign v_12198 = v_816 & v_12197;
assign v_12199 = v_832 & v_838;
assign v_12201 = v_561 & v_12200;
assign v_12202 = v_715 & v_721;
assign v_12204 = v_9618 & v_9753;
assign v_12205 = v_9604 & v_9646;
assign v_12207 = v_9473 & v_12206;
assign v_12208 = v_9463 & v_9488;
assign v_12210 = v_9329 & v_12209;
assign v_12211 = v_9311 & v_9356;
assign v_12213 = v_9185 & v_12212;
assign v_12214 = v_9175 & v_9200;
assign v_12216 = v_9044 & v_12215;
assign v_12217 = v_9030 & v_9068;
assign v_12219 = v_8903 & v_12218;
assign v_12220 = v_8893 & v_8918;
assign v_12222 = v_8755 & v_12221;
assign v_12223 = v_8733 & v_8786;
assign v_12225 = v_8607 & v_12224;
assign v_12226 = v_8597 & v_8622;
assign v_12228 = v_8465 & v_12227;
assign v_12229 = v_8451 & v_8490;
assign v_12231 = v_8323 & v_12230;
assign v_12232 = v_8313 & v_8338;
assign v_12234 = v_8179 & v_12233;
assign v_12235 = v_8161 & v_8206;
assign v_12237 = v_8035 & v_12236;
assign v_12238 = v_8025 & v_8050;
assign v_12240 = v_7894 & v_12239;
assign v_12241 = v_7880 & v_7918;
assign v_12243 = v_7753 & v_12242;
assign v_12244 = v_7743 & v_7768;
assign v_12246 = v_7601 & v_12245;
assign v_12247 = v_7575 & v_7636;
assign v_12249 = v_7449 & v_12248;
assign v_12250 = v_7439 & v_7464;
assign v_12252 = v_7306 & v_12251;
assign v_12253 = v_7292 & v_7332;
assign v_12255 = v_7163 & v_12254;
assign v_12256 = v_7153 & v_7178;
assign v_12258 = v_7019 & v_12257;
assign v_12259 = v_7001 & v_7046;
assign v_12261 = v_6875 & v_12260;
assign v_12262 = v_6865 & v_6890;
assign v_12264 = v_6734 & v_12263;
assign v_12265 = v_6720 & v_6758;
assign v_12267 = v_6593 & v_12266;
assign v_12268 = v_6583 & v_6608;
assign v_12270 = v_6445 & v_12269;
assign v_12271 = v_6423 & v_6476;
assign v_12273 = v_6297 & v_12272;
assign v_12274 = v_6287 & v_6312;
assign v_12276 = v_6155 & v_12275;
assign v_12277 = v_6141 & v_6180;
assign v_12279 = v_6013 & v_12278;
assign v_12280 = v_6003 & v_6028;
assign v_12282 = v_5869 & v_12281;
assign v_12283 = v_5851 & v_5896;
assign v_12285 = v_5725 & v_12284;
assign v_12286 = v_5715 & v_5740;
assign v_12288 = v_5584 & v_12287;
assign v_12289 = v_5570 & v_5608;
assign v_12291 = v_5443 & v_12290;
assign v_12292 = v_5433 & v_5458;
assign v_12294 = v_5287 & v_12293;
assign v_12295 = v_5257 & v_5326;
assign v_12297 = v_5131 & v_12296;
assign v_12298 = v_5121 & v_5146;
assign v_12300 = v_4987 & v_12299;
assign v_12301 = v_4973 & v_5014;
assign v_12303 = v_4843 & v_12302;
assign v_12304 = v_4833 & v_4858;
assign v_12306 = v_4699 & v_12305;
assign v_12307 = v_4681 & v_4726;
assign v_12309 = v_4555 & v_12308;
assign v_12310 = v_4545 & v_4570;
assign v_12312 = v_4414 & v_12311;
assign v_12313 = v_4400 & v_4438;
assign v_12315 = v_4273 & v_12314;
assign v_12316 = v_4263 & v_4288;
assign v_12318 = v_4125 & v_12317;
assign v_12319 = v_4103 & v_4156;
assign v_12321 = v_3977 & v_12320;
assign v_12322 = v_3967 & v_3992;
assign v_12324 = v_3835 & v_12323;
assign v_12325 = v_3821 & v_3860;
assign v_12327 = v_3693 & v_12326;
assign v_12328 = v_3683 & v_3708;
assign v_12330 = v_3549 & v_12329;
assign v_12331 = v_3531 & v_3576;
assign v_12333 = v_3405 & v_12332;
assign v_12334 = v_3395 & v_3420;
assign v_12336 = v_3264 & v_12335;
assign v_12337 = v_3250 & v_3288;
assign v_12339 = v_3123 & v_12338;
assign v_12340 = v_3113 & v_3138;
assign v_12342 = v_2971 & v_12341;
assign v_12343 = v_2945 & v_3006;
assign v_12345 = v_2819 & v_12344;
assign v_12346 = v_2809 & v_2834;
assign v_12348 = v_2676 & v_12347;
assign v_12349 = v_2662 & v_2702;
assign v_12351 = v_2533 & v_12350;
assign v_12352 = v_2523 & v_2548;
assign v_12354 = v_2389 & v_12353;
assign v_12355 = v_2371 & v_2416;
assign v_12357 = v_2245 & v_12356;
assign v_12358 = v_2235 & v_2260;
assign v_12360 = v_2104 & v_12359;
assign v_12361 = v_2090 & v_2128;
assign v_12363 = v_1963 & v_12362;
assign v_12364 = v_1953 & v_1978;
assign v_12366 = v_1815 & v_12365;
assign v_12367 = v_1793 & v_1846;
assign v_12369 = v_1667 & v_12368;
assign v_12370 = v_1657 & v_1682;
assign v_12372 = v_1525 & v_12371;
assign v_12373 = v_1511 & v_1550;
assign v_12375 = v_1383 & v_12374;
assign v_12376 = v_1373 & v_1398;
assign v_12378 = v_1239 & v_12377;
assign v_12379 = v_1221 & v_1266;
assign v_12381 = v_1095 & v_12380;
assign v_12382 = v_1085 & v_1110;
assign v_12384 = v_954 & v_12383;
assign v_12385 = v_940 & v_978;
assign v_12387 = v_816 & v_12386;
assign v_12388 = v_804 & v_832;
assign v_12390 = v_561 & v_12389;
assign v_12391 = v_98 & v_715;
assign v_12394 = v_9618 & v_9796;
assign v_12395 = v_9646 & v_9664;
assign v_12397 = v_9473 & v_12396;
assign v_12398 = v_9488 & v_9506;
assign v_12400 = v_9329 & v_12399;
assign v_12401 = v_9356 & v_9374;
assign v_12403 = v_9185 & v_12402;
assign v_12404 = v_9200 & v_9218;
assign v_12406 = v_9044 & v_12405;
assign v_12407 = v_9068 & v_9086;
assign v_12409 = v_8903 & v_12408;
assign v_12410 = v_8918 & v_8936;
assign v_12412 = v_8755 & v_12411;
assign v_12413 = v_8786 & v_8804;
assign v_12415 = v_8607 & v_12414;
assign v_12416 = v_8622 & v_8640;
assign v_12418 = v_8465 & v_12417;
assign v_12419 = v_8490 & v_8508;
assign v_12421 = v_8323 & v_12420;
assign v_12422 = v_8338 & v_8356;
assign v_12424 = v_8179 & v_12423;
assign v_12425 = v_8206 & v_8224;
assign v_12427 = v_8035 & v_12426;
assign v_12428 = v_8050 & v_8068;
assign v_12430 = v_7894 & v_12429;
assign v_12431 = v_7918 & v_7936;
assign v_12433 = v_7753 & v_12432;
assign v_12434 = v_7768 & v_7786;
assign v_12436 = v_7601 & v_12435;
assign v_12437 = v_7636 & v_7654;
assign v_12439 = v_7449 & v_12438;
assign v_12440 = v_7464 & v_7482;
assign v_12442 = v_7306 & v_12441;
assign v_12443 = v_7332 & v_7350;
assign v_12445 = v_7163 & v_12444;
assign v_12446 = v_7178 & v_7196;
assign v_12448 = v_7019 & v_12447;
assign v_12449 = v_7046 & v_7064;
assign v_12451 = v_6875 & v_12450;
assign v_12452 = v_6890 & v_6908;
assign v_12454 = v_6734 & v_12453;
assign v_12455 = v_6758 & v_6776;
assign v_12457 = v_6593 & v_12456;
assign v_12458 = v_6608 & v_6626;
assign v_12460 = v_6445 & v_12459;
assign v_12461 = v_6476 & v_6494;
assign v_12463 = v_6297 & v_12462;
assign v_12464 = v_6312 & v_6330;
assign v_12466 = v_6155 & v_12465;
assign v_12467 = v_6180 & v_6198;
assign v_12469 = v_6013 & v_12468;
assign v_12470 = v_6028 & v_6046;
assign v_12472 = v_5869 & v_12471;
assign v_12473 = v_5896 & v_5914;
assign v_12475 = v_5725 & v_12474;
assign v_12476 = v_5740 & v_5758;
assign v_12478 = v_5584 & v_12477;
assign v_12479 = v_5608 & v_5626;
assign v_12481 = v_5443 & v_12480;
assign v_12482 = v_5458 & v_5476;
assign v_12484 = v_5287 & v_12483;
assign v_12485 = v_5326 & v_5344;
assign v_12487 = v_5131 & v_12486;
assign v_12488 = v_5146 & v_5164;
assign v_12490 = v_4987 & v_12489;
assign v_12491 = v_5014 & v_5032;
assign v_12493 = v_4843 & v_12492;
assign v_12494 = v_4858 & v_4876;
assign v_12496 = v_4699 & v_12495;
assign v_12497 = v_4726 & v_4744;
assign v_12499 = v_4555 & v_12498;
assign v_12500 = v_4570 & v_4588;
assign v_12502 = v_4414 & v_12501;
assign v_12503 = v_4438 & v_4456;
assign v_12505 = v_4273 & v_12504;
assign v_12506 = v_4288 & v_4306;
assign v_12508 = v_4125 & v_12507;
assign v_12509 = v_4156 & v_4174;
assign v_12511 = v_3977 & v_12510;
assign v_12512 = v_3992 & v_4010;
assign v_12514 = v_3835 & v_12513;
assign v_12515 = v_3860 & v_3878;
assign v_12517 = v_3693 & v_12516;
assign v_12518 = v_3708 & v_3726;
assign v_12520 = v_3549 & v_12519;
assign v_12521 = v_3576 & v_3594;
assign v_12523 = v_3405 & v_12522;
assign v_12524 = v_3420 & v_3438;
assign v_12526 = v_3264 & v_12525;
assign v_12527 = v_3288 & v_3306;
assign v_12529 = v_3123 & v_12528;
assign v_12530 = v_3138 & v_3156;
assign v_12532 = v_2971 & v_12531;
assign v_12533 = v_3006 & v_3024;
assign v_12535 = v_2819 & v_12534;
assign v_12536 = v_2834 & v_2852;
assign v_12538 = v_2676 & v_12537;
assign v_12539 = v_2702 & v_2720;
assign v_12541 = v_2533 & v_12540;
assign v_12542 = v_2548 & v_2566;
assign v_12544 = v_2389 & v_12543;
assign v_12545 = v_2416 & v_2434;
assign v_12547 = v_2245 & v_12546;
assign v_12548 = v_2260 & v_2278;
assign v_12550 = v_2104 & v_12549;
assign v_12551 = v_2128 & v_2146;
assign v_12553 = v_1963 & v_12552;
assign v_12554 = v_1978 & v_1996;
assign v_12556 = v_1815 & v_12555;
assign v_12557 = v_1846 & v_1864;
assign v_12559 = v_1667 & v_12558;
assign v_12560 = v_1682 & v_1700;
assign v_12562 = v_1525 & v_12561;
assign v_12563 = v_1550 & v_1568;
assign v_12565 = v_1383 & v_12564;
assign v_12566 = v_1398 & v_1416;
assign v_12568 = v_1239 & v_12567;
assign v_12569 = v_1266 & v_1284;
assign v_12571 = v_1095 & v_12570;
assign v_12572 = v_1110 & v_1128;
assign v_12574 = v_954 & v_12573;
assign v_12575 = v_978 & v_996;
assign v_12577 = v_816 & v_12576;
assign v_12578 = v_832 & v_850;
assign v_12580 = v_561 & v_12579;
assign v_12581 = v_715 & v_731;
assign v_12584 = v_9618 & v_9808;
assign v_12585 = v_9646 & v_9676;
assign v_12587 = v_9473 & v_12586;
assign v_12588 = v_9488 & v_9518;
assign v_12590 = v_9329 & v_12589;
assign v_12591 = v_9356 & v_9386;
assign v_12593 = v_9185 & v_12592;
assign v_12594 = v_9200 & v_9230;
assign v_12596 = v_9044 & v_12595;
assign v_12597 = v_9068 & v_9098;
assign v_12599 = v_8903 & v_12598;
assign v_12600 = v_8918 & v_8948;
assign v_12602 = v_8755 & v_12601;
assign v_12603 = v_8786 & v_8816;
assign v_12605 = v_8607 & v_12604;
assign v_12606 = v_8622 & v_8652;
assign v_12608 = v_8465 & v_12607;
assign v_12609 = v_8490 & v_8520;
assign v_12611 = v_8323 & v_12610;
assign v_12612 = v_8338 & v_8368;
assign v_12614 = v_8179 & v_12613;
assign v_12615 = v_8206 & v_8236;
assign v_12617 = v_8035 & v_12616;
assign v_12618 = v_8050 & v_8080;
assign v_12620 = v_7894 & v_12619;
assign v_12621 = v_7918 & v_7948;
assign v_12623 = v_7753 & v_12622;
assign v_12624 = v_7768 & v_7798;
assign v_12626 = v_7601 & v_12625;
assign v_12627 = v_7636 & v_7666;
assign v_12629 = v_7449 & v_12628;
assign v_12630 = v_7464 & v_7494;
assign v_12632 = v_7306 & v_12631;
assign v_12633 = v_7332 & v_7362;
assign v_12635 = v_7163 & v_12634;
assign v_12636 = v_7178 & v_7208;
assign v_12638 = v_7019 & v_12637;
assign v_12639 = v_7046 & v_7076;
assign v_12641 = v_6875 & v_12640;
assign v_12642 = v_6890 & v_6920;
assign v_12644 = v_6734 & v_12643;
assign v_12645 = v_6758 & v_6788;
assign v_12647 = v_6593 & v_12646;
assign v_12648 = v_6608 & v_6638;
assign v_12650 = v_6445 & v_12649;
assign v_12651 = v_6476 & v_6506;
assign v_12653 = v_6297 & v_12652;
assign v_12654 = v_6312 & v_6342;
assign v_12656 = v_6155 & v_12655;
assign v_12657 = v_6180 & v_6210;
assign v_12659 = v_6013 & v_12658;
assign v_12660 = v_6028 & v_6058;
assign v_12662 = v_5869 & v_12661;
assign v_12663 = v_5896 & v_5926;
assign v_12665 = v_5725 & v_12664;
assign v_12666 = v_5740 & v_5770;
assign v_12668 = v_5584 & v_12667;
assign v_12669 = v_5608 & v_5638;
assign v_12671 = v_5443 & v_12670;
assign v_12672 = v_5458 & v_5488;
assign v_12674 = v_5287 & v_12673;
assign v_12675 = v_5326 & v_5356;
assign v_12677 = v_5131 & v_12676;
assign v_12678 = v_5146 & v_5176;
assign v_12680 = v_4987 & v_12679;
assign v_12681 = v_5014 & v_5044;
assign v_12683 = v_4843 & v_12682;
assign v_12684 = v_4858 & v_4888;
assign v_12686 = v_4699 & v_12685;
assign v_12687 = v_4726 & v_4756;
assign v_12689 = v_4555 & v_12688;
assign v_12690 = v_4570 & v_4600;
assign v_12692 = v_4414 & v_12691;
assign v_12693 = v_4438 & v_4468;
assign v_12695 = v_4273 & v_12694;
assign v_12696 = v_4288 & v_4318;
assign v_12698 = v_4125 & v_12697;
assign v_12699 = v_4156 & v_4186;
assign v_12701 = v_3977 & v_12700;
assign v_12702 = v_3992 & v_4022;
assign v_12704 = v_3835 & v_12703;
assign v_12705 = v_3860 & v_3890;
assign v_12707 = v_3693 & v_12706;
assign v_12708 = v_3708 & v_3738;
assign v_12710 = v_3549 & v_12709;
assign v_12711 = v_3576 & v_3606;
assign v_12713 = v_3405 & v_12712;
assign v_12714 = v_3420 & v_3450;
assign v_12716 = v_3264 & v_12715;
assign v_12717 = v_3288 & v_3318;
assign v_12719 = v_3123 & v_12718;
assign v_12720 = v_3138 & v_3168;
assign v_12722 = v_2971 & v_12721;
assign v_12723 = v_3006 & v_3036;
assign v_12725 = v_2819 & v_12724;
assign v_12726 = v_2834 & v_2864;
assign v_12728 = v_2676 & v_12727;
assign v_12729 = v_2702 & v_2732;
assign v_12731 = v_2533 & v_12730;
assign v_12732 = v_2548 & v_2578;
assign v_12734 = v_2389 & v_12733;
assign v_12735 = v_2416 & v_2446;
assign v_12737 = v_2245 & v_12736;
assign v_12738 = v_2260 & v_2290;
assign v_12740 = v_2104 & v_12739;
assign v_12741 = v_2128 & v_2158;
assign v_12743 = v_1963 & v_12742;
assign v_12744 = v_1978 & v_2008;
assign v_12746 = v_1815 & v_12745;
assign v_12747 = v_1846 & v_1876;
assign v_12749 = v_1667 & v_12748;
assign v_12750 = v_1682 & v_1712;
assign v_12752 = v_1525 & v_12751;
assign v_12753 = v_1550 & v_1580;
assign v_12755 = v_1383 & v_12754;
assign v_12756 = v_1398 & v_1428;
assign v_12758 = v_1239 & v_12757;
assign v_12759 = v_1266 & v_1296;
assign v_12761 = v_1095 & v_12760;
assign v_12762 = v_1110 & v_1140;
assign v_12764 = v_954 & v_12763;
assign v_12765 = v_978 & v_1008;
assign v_12767 = v_816 & v_12766;
assign v_12768 = v_832 & v_862;
assign v_12770 = v_561 & v_12769;
assign v_12771 = v_715 & v_741;
assign v_12774 = v_9618 & v_9820;
assign v_12775 = v_9646 & v_9688;
assign v_12777 = v_9473 & v_12776;
assign v_12778 = v_9488 & v_9530;
assign v_12780 = v_9329 & v_12779;
assign v_12781 = v_9356 & v_9398;
assign v_12783 = v_9185 & v_12782;
assign v_12784 = v_9200 & v_9242;
assign v_12786 = v_9044 & v_12785;
assign v_12787 = v_9068 & v_9110;
assign v_12789 = v_8903 & v_12788;
assign v_12790 = v_8918 & v_8960;
assign v_12792 = v_8755 & v_12791;
assign v_12793 = v_8786 & v_8828;
assign v_12795 = v_8607 & v_12794;
assign v_12796 = v_8622 & v_8664;
assign v_12798 = v_8465 & v_12797;
assign v_12799 = v_8490 & v_8532;
assign v_12801 = v_8323 & v_12800;
assign v_12802 = v_8338 & v_8380;
assign v_12804 = v_8179 & v_12803;
assign v_12805 = v_8206 & v_8248;
assign v_12807 = v_8035 & v_12806;
assign v_12808 = v_8050 & v_8092;
assign v_12810 = v_7894 & v_12809;
assign v_12811 = v_7918 & v_7960;
assign v_12813 = v_7753 & v_12812;
assign v_12814 = v_7768 & v_7810;
assign v_12816 = v_7601 & v_12815;
assign v_12817 = v_7636 & v_7678;
assign v_12819 = v_7449 & v_12818;
assign v_12820 = v_7464 & v_7506;
assign v_12822 = v_7306 & v_12821;
assign v_12823 = v_7332 & v_7374;
assign v_12825 = v_7163 & v_12824;
assign v_12826 = v_7178 & v_7220;
assign v_12828 = v_7019 & v_12827;
assign v_12829 = v_7046 & v_7088;
assign v_12831 = v_6875 & v_12830;
assign v_12832 = v_6890 & v_6932;
assign v_12834 = v_6734 & v_12833;
assign v_12835 = v_6758 & v_6800;
assign v_12837 = v_6593 & v_12836;
assign v_12838 = v_6608 & v_6650;
assign v_12840 = v_6445 & v_12839;
assign v_12841 = v_6476 & v_6518;
assign v_12843 = v_6297 & v_12842;
assign v_12844 = v_6312 & v_6354;
assign v_12846 = v_6155 & v_12845;
assign v_12847 = v_6180 & v_6222;
assign v_12849 = v_6013 & v_12848;
assign v_12850 = v_6028 & v_6070;
assign v_12852 = v_5869 & v_12851;
assign v_12853 = v_5896 & v_5938;
assign v_12855 = v_5725 & v_12854;
assign v_12856 = v_5740 & v_5782;
assign v_12858 = v_5584 & v_12857;
assign v_12859 = v_5608 & v_5650;
assign v_12861 = v_5443 & v_12860;
assign v_12862 = v_5458 & v_5500;
assign v_12864 = v_5287 & v_12863;
assign v_12865 = v_5326 & v_5368;
assign v_12867 = v_5131 & v_12866;
assign v_12868 = v_5146 & v_5188;
assign v_12870 = v_4987 & v_12869;
assign v_12871 = v_5014 & v_5056;
assign v_12873 = v_4843 & v_12872;
assign v_12874 = v_4858 & v_4900;
assign v_12876 = v_4699 & v_12875;
assign v_12877 = v_4726 & v_4768;
assign v_12879 = v_4555 & v_12878;
assign v_12880 = v_4570 & v_4612;
assign v_12882 = v_4414 & v_12881;
assign v_12883 = v_4438 & v_4480;
assign v_12885 = v_4273 & v_12884;
assign v_12886 = v_4288 & v_4330;
assign v_12888 = v_4125 & v_12887;
assign v_12889 = v_4156 & v_4198;
assign v_12891 = v_3977 & v_12890;
assign v_12892 = v_3992 & v_4034;
assign v_12894 = v_3835 & v_12893;
assign v_12895 = v_3860 & v_3902;
assign v_12897 = v_3693 & v_12896;
assign v_12898 = v_3708 & v_3750;
assign v_12900 = v_3549 & v_12899;
assign v_12901 = v_3576 & v_3618;
assign v_12903 = v_3405 & v_12902;
assign v_12904 = v_3420 & v_3462;
assign v_12906 = v_3264 & v_12905;
assign v_12907 = v_3288 & v_3330;
assign v_12909 = v_3123 & v_12908;
assign v_12910 = v_3138 & v_3180;
assign v_12912 = v_2971 & v_12911;
assign v_12913 = v_3006 & v_3048;
assign v_12915 = v_2819 & v_12914;
assign v_12916 = v_2834 & v_2876;
assign v_12918 = v_2676 & v_12917;
assign v_12919 = v_2702 & v_2744;
assign v_12921 = v_2533 & v_12920;
assign v_12922 = v_2548 & v_2590;
assign v_12924 = v_2389 & v_12923;
assign v_12925 = v_2416 & v_2458;
assign v_12927 = v_2245 & v_12926;
assign v_12928 = v_2260 & v_2302;
assign v_12930 = v_2104 & v_12929;
assign v_12931 = v_2128 & v_2170;
assign v_12933 = v_1963 & v_12932;
assign v_12934 = v_1978 & v_2020;
assign v_12936 = v_1815 & v_12935;
assign v_12937 = v_1846 & v_1888;
assign v_12939 = v_1667 & v_12938;
assign v_12940 = v_1682 & v_1724;
assign v_12942 = v_1525 & v_12941;
assign v_12943 = v_1550 & v_1592;
assign v_12945 = v_1383 & v_12944;
assign v_12946 = v_1398 & v_1440;
assign v_12948 = v_1239 & v_12947;
assign v_12949 = v_1266 & v_1308;
assign v_12951 = v_1095 & v_12950;
assign v_12952 = v_1110 & v_1152;
assign v_12954 = v_954 & v_12953;
assign v_12955 = v_978 & v_1020;
assign v_12957 = v_816 & v_12956;
assign v_12958 = v_832 & v_874;
assign v_12960 = v_561 & v_12959;
assign v_12961 = v_715 & v_751;
assign v_12964 = v_9618 & v_9832;
assign v_12965 = v_9646 & v_9700;
assign v_12967 = v_9473 & v_12966;
assign v_12968 = v_9488 & v_9542;
assign v_12970 = v_9329 & v_12969;
assign v_12971 = v_9356 & v_9410;
assign v_12973 = v_9185 & v_12972;
assign v_12974 = v_9200 & v_9254;
assign v_12976 = v_9044 & v_12975;
assign v_12977 = v_9068 & v_9122;
assign v_12979 = v_8903 & v_12978;
assign v_12980 = v_8918 & v_8972;
assign v_12982 = v_8755 & v_12981;
assign v_12983 = v_8786 & v_8840;
assign v_12985 = v_8607 & v_12984;
assign v_12986 = v_8622 & v_8676;
assign v_12988 = v_8465 & v_12987;
assign v_12989 = v_8490 & v_8544;
assign v_12991 = v_8323 & v_12990;
assign v_12992 = v_8338 & v_8392;
assign v_12994 = v_8179 & v_12993;
assign v_12995 = v_8206 & v_8260;
assign v_12997 = v_8035 & v_12996;
assign v_12998 = v_8050 & v_8104;
assign v_13000 = v_7894 & v_12999;
assign v_13001 = v_7918 & v_7972;
assign v_13003 = v_7753 & v_13002;
assign v_13004 = v_7768 & v_7822;
assign v_13006 = v_7601 & v_13005;
assign v_13007 = v_7636 & v_7690;
assign v_13009 = v_7449 & v_13008;
assign v_13010 = v_7464 & v_7518;
assign v_13012 = v_7306 & v_13011;
assign v_13013 = v_7332 & v_7386;
assign v_13015 = v_7163 & v_13014;
assign v_13016 = v_7178 & v_7232;
assign v_13018 = v_7019 & v_13017;
assign v_13019 = v_7046 & v_7100;
assign v_13021 = v_6875 & v_13020;
assign v_13022 = v_6890 & v_6944;
assign v_13024 = v_6734 & v_13023;
assign v_13025 = v_6758 & v_6812;
assign v_13027 = v_6593 & v_13026;
assign v_13028 = v_6608 & v_6662;
assign v_13030 = v_6445 & v_13029;
assign v_13031 = v_6476 & v_6530;
assign v_13033 = v_6297 & v_13032;
assign v_13034 = v_6312 & v_6366;
assign v_13036 = v_6155 & v_13035;
assign v_13037 = v_6180 & v_6234;
assign v_13039 = v_6013 & v_13038;
assign v_13040 = v_6028 & v_6082;
assign v_13042 = v_5869 & v_13041;
assign v_13043 = v_5896 & v_5950;
assign v_13045 = v_5725 & v_13044;
assign v_13046 = v_5740 & v_5794;
assign v_13048 = v_5584 & v_13047;
assign v_13049 = v_5608 & v_5662;
assign v_13051 = v_5443 & v_13050;
assign v_13052 = v_5458 & v_5512;
assign v_13054 = v_5287 & v_13053;
assign v_13055 = v_5326 & v_5380;
assign v_13057 = v_5131 & v_13056;
assign v_13058 = v_5146 & v_5200;
assign v_13060 = v_4987 & v_13059;
assign v_13061 = v_5014 & v_5068;
assign v_13063 = v_4843 & v_13062;
assign v_13064 = v_4858 & v_4912;
assign v_13066 = v_4699 & v_13065;
assign v_13067 = v_4726 & v_4780;
assign v_13069 = v_4555 & v_13068;
assign v_13070 = v_4570 & v_4624;
assign v_13072 = v_4414 & v_13071;
assign v_13073 = v_4438 & v_4492;
assign v_13075 = v_4273 & v_13074;
assign v_13076 = v_4288 & v_4342;
assign v_13078 = v_4125 & v_13077;
assign v_13079 = v_4156 & v_4210;
assign v_13081 = v_3977 & v_13080;
assign v_13082 = v_3992 & v_4046;
assign v_13084 = v_3835 & v_13083;
assign v_13085 = v_3860 & v_3914;
assign v_13087 = v_3693 & v_13086;
assign v_13088 = v_3708 & v_3762;
assign v_13090 = v_3549 & v_13089;
assign v_13091 = v_3576 & v_3630;
assign v_13093 = v_3405 & v_13092;
assign v_13094 = v_3420 & v_3474;
assign v_13096 = v_3264 & v_13095;
assign v_13097 = v_3288 & v_3342;
assign v_13099 = v_3123 & v_13098;
assign v_13100 = v_3138 & v_3192;
assign v_13102 = v_2971 & v_13101;
assign v_13103 = v_3006 & v_3060;
assign v_13105 = v_2819 & v_13104;
assign v_13106 = v_2834 & v_2888;
assign v_13108 = v_2676 & v_13107;
assign v_13109 = v_2702 & v_2756;
assign v_13111 = v_2533 & v_13110;
assign v_13112 = v_2548 & v_2602;
assign v_13114 = v_2389 & v_13113;
assign v_13115 = v_2416 & v_2470;
assign v_13117 = v_2245 & v_13116;
assign v_13118 = v_2260 & v_2314;
assign v_13120 = v_2104 & v_13119;
assign v_13121 = v_2128 & v_2182;
assign v_13123 = v_1963 & v_13122;
assign v_13124 = v_1978 & v_2032;
assign v_13126 = v_1815 & v_13125;
assign v_13127 = v_1846 & v_1900;
assign v_13129 = v_1667 & v_13128;
assign v_13130 = v_1682 & v_1736;
assign v_13132 = v_1525 & v_13131;
assign v_13133 = v_1550 & v_1604;
assign v_13135 = v_1383 & v_13134;
assign v_13136 = v_1398 & v_1452;
assign v_13138 = v_1239 & v_13137;
assign v_13139 = v_1266 & v_1320;
assign v_13141 = v_1095 & v_13140;
assign v_13142 = v_1110 & v_1164;
assign v_13144 = v_954 & v_13143;
assign v_13145 = v_978 & v_1032;
assign v_13147 = v_816 & v_13146;
assign v_13148 = v_832 & v_886;
assign v_13150 = v_561 & v_13149;
assign v_13151 = v_715 & v_761;
assign v_13156 = v_13154 & v_13155;
assign v_13159 = v_13157 & v_13158;
assign v_13162 = v_13160 & v_13161;
assign v_13165 = v_13163 & v_13164;
assign v_13168 = v_13166 & v_13167;
assign v_13171 = v_13169 & v_13170;
assign v_13174 = v_13172 & v_13173;
assign v_13177 = v_13175 & v_13176;
assign v_13180 = v_13178 & v_13179;
assign v_13183 = v_13181 & v_13182;
assign v_13186 = v_13184 & v_13185;
assign v_13189 = v_13187 & v_13188;
assign v_13192 = v_13190 & v_13191;
assign v_13195 = v_13193 & v_13194;
assign v_13198 = v_13196 & v_13197;
assign v_13201 = v_13199 & v_13200;
assign v_13204 = v_13202 & v_13203;
assign v_13207 = v_13205 & v_13206;
assign v_13210 = v_13208 & v_13209;
assign v_13213 = v_13211 & v_13212;
assign v_13216 = v_13214 & v_13215;
assign v_13219 = v_13217 & v_13218;
assign v_13222 = v_13220 & v_13221;
assign v_13225 = v_13223 & v_13224;
assign v_13228 = v_13226 & v_13227;
assign v_13231 = v_13229 & v_13230;
assign v_13234 = v_13232 & v_13233;
assign v_13237 = v_13235 & v_13236;
assign v_13240 = v_13238 & v_13239;
assign v_13243 = v_13241 & v_13242;
assign v_13246 = v_13244 & v_13245;
assign v_13249 = v_13247 & v_13248;
assign v_13252 = v_13250 & v_13251;
assign v_13255 = v_13253 & v_13254;
assign v_13258 = v_13256 & v_13257;
assign v_13261 = v_13259 & v_13260;
assign v_13264 = v_13262 & v_13263;
assign v_13267 = v_13265 & v_13266;
assign v_13270 = v_13268 & v_13269;
assign v_13273 = v_13271 & v_13272;
assign v_13276 = v_13274 & v_13275;
assign v_13279 = v_13277 & v_13278;
assign v_13282 = v_13280 & v_13281;
assign v_13285 = v_13283 & v_13284;
assign v_13288 = v_13286 & v_13287;
assign v_13291 = v_13289 & v_13290;
assign v_13294 = v_13292 & v_13293;
assign v_13297 = v_13295 & v_13296;
assign v_13300 = v_13298 & v_13299;
assign v_13303 = v_13301 & v_13302;
assign v_13306 = v_13304 & v_13305;
assign v_13309 = v_13307 & v_13308;
assign v_13312 = v_13310 & v_13311;
assign v_13315 = v_13313 & v_13314;
assign v_13318 = v_13316 & v_13317;
assign v_13321 = v_13319 & v_13320;
assign v_13324 = v_13322 & v_13323;
assign v_13327 = v_13325 & v_13326;
assign v_13330 = v_13328 & v_13329;
assign v_13333 = v_13331 & v_13332;
assign v_13336 = v_13334 & v_13335;
assign v_13339 = v_13337 & v_13338;
assign v_13342 = v_13340 & v_13341;
assign v_13344 = v_9618 & ~v_9872;
assign v_13345 = v_9646 & ~v_9740;
assign v_13347 = v_9473 & v_13346;
assign v_13348 = v_9488 & ~v_9582;
assign v_13350 = v_9329 & v_13349;
assign v_13351 = v_9356 & ~v_9450;
assign v_13353 = v_9185 & v_13352;
assign v_13354 = v_9200 & ~v_9294;
assign v_13356 = v_9044 & v_13355;
assign v_13357 = v_9068 & ~v_9162;
assign v_13359 = v_8903 & v_13358;
assign v_13360 = v_8918 & ~v_9012;
assign v_13362 = v_8755 & v_13361;
assign v_13363 = v_8786 & ~v_8880;
assign v_13365 = v_8607 & v_13364;
assign v_13366 = v_8622 & ~v_8716;
assign v_13368 = v_8465 & v_13367;
assign v_13369 = v_8490 & ~v_8584;
assign v_13371 = v_8323 & v_13370;
assign v_13372 = v_8338 & v_8432;
assign v_13374 = v_8179 & v_13373;
assign v_13375 = v_8206 & v_8300;
assign v_13377 = v_8035 & v_13376;
assign v_13378 = v_8050 & v_8144;
assign v_13380 = v_7894 & v_13379;
assign v_13381 = v_7918 & ~v_8012;
assign v_13383 = v_7753 & v_13382;
assign v_13384 = v_7768 & ~v_7862;
assign v_13386 = v_7601 & v_13385;
assign v_13387 = v_7636 & ~v_7730;
assign v_13389 = v_7449 & v_13388;
assign v_13390 = v_7464 & ~v_7558;
assign v_13392 = v_7306 & v_13391;
assign v_13393 = v_7332 & ~v_7426;
assign v_13395 = v_7163 & v_13394;
assign v_13396 = v_7178 & v_7272;
assign v_13398 = v_7019 & v_13397;
assign v_13399 = v_7046 & ~v_7140;
assign v_13401 = v_6875 & v_13400;
assign v_13402 = v_6890 & v_6984;
assign v_13404 = v_6734 & v_13403;
assign v_13405 = v_6758 & v_6852;
assign v_13407 = v_6593 & v_13406;
assign v_13408 = v_6608 & v_6702;
assign v_13410 = v_6445 & v_13409;
assign v_13411 = v_6476 & ~v_6570;
assign v_13413 = v_6297 & v_13412;
assign v_13414 = v_6312 & ~v_6406;
assign v_13416 = v_6155 & v_13415;
assign v_13417 = v_6180 & v_6274;
assign v_13419 = v_6013 & v_13418;
assign v_13420 = v_6028 & v_6122;
assign v_13422 = v_5869 & v_13421;
assign v_13423 = v_5896 & v_5990;
assign v_13425 = v_5725 & v_13424;
assign v_13426 = v_5740 & v_5834;
assign v_13428 = v_5584 & v_13427;
assign v_13429 = v_5608 & v_5702;
assign v_13431 = v_5443 & v_13430;
assign v_13432 = v_5458 & v_5552;
assign v_13434 = v_5287 & v_13433;
assign v_13435 = v_5326 & ~v_5420;
assign v_13437 = v_5131 & v_13436;
assign v_13438 = v_5146 & ~v_5240;
assign v_13440 = v_4987 & v_13439;
assign v_13441 = v_5014 & v_5108;
assign v_13443 = v_4843 & v_13442;
assign v_13444 = v_4858 & v_4952;
assign v_13446 = v_4699 & v_13445;
assign v_13447 = v_4726 & v_4820;
assign v_13449 = v_4555 & v_13448;
assign v_13450 = v_4570 & v_4664;
assign v_13452 = v_4414 & v_13451;
assign v_13453 = v_4438 & v_4532;
assign v_13455 = v_4273 & v_13454;
assign v_13456 = v_4288 & v_4382;
assign v_13458 = v_4125 & v_13457;
assign v_13459 = v_4156 & ~v_4250;
assign v_13461 = v_3977 & v_13460;
assign v_13462 = v_3992 & ~v_4086;
assign v_13464 = v_3835 & v_13463;
assign v_13465 = v_3860 & ~v_3954;
assign v_13467 = v_3693 & v_13466;
assign v_13468 = v_3708 & ~v_3802;
assign v_13470 = v_3549 & v_13469;
assign v_13471 = v_3576 & ~v_3670;
assign v_13473 = v_3405 & v_13472;
assign v_13474 = v_3420 & v_3514;
assign v_13476 = v_3264 & v_13475;
assign v_13477 = v_3288 & ~v_3382;
assign v_13479 = v_3123 & v_13478;
assign v_13480 = v_3138 & v_3232;
assign v_13482 = v_2971 & v_13481;
assign v_13483 = v_3006 & ~v_3100;
assign v_13485 = v_2819 & v_13484;
assign v_13486 = v_2834 & ~v_2928;
assign v_13488 = v_2676 & v_13487;
assign v_13489 = v_2702 & ~v_2796;
assign v_13491 = v_2533 & v_13490;
assign v_13492 = v_2548 & ~v_2642;
assign v_13494 = v_2389 & v_13493;
assign v_13495 = v_2416 & ~v_2510;
assign v_13497 = v_2245 & v_13496;
assign v_13498 = v_2260 & v_2354;
assign v_13500 = v_2104 & v_13499;
assign v_13501 = v_2128 & v_2222;
assign v_13503 = v_1963 & v_13502;
assign v_13504 = v_1978 & v_2072;
assign v_13506 = v_1815 & v_13505;
assign v_13507 = v_1846 & ~v_1940;
assign v_13509 = v_1667 & v_13508;
assign v_13510 = v_1682 & ~v_1776;
assign v_13512 = v_1525 & v_13511;
assign v_13513 = v_1550 & ~v_1644;
assign v_13515 = v_1383 & v_13514;
assign v_13516 = v_1398 & ~v_1492;
assign v_13518 = v_1239 & v_13517;
assign v_13519 = v_1266 & ~v_1360;
assign v_13521 = v_1095 & v_13520;
assign v_13522 = v_1110 & ~v_1204;
assign v_13524 = v_954 & v_13523;
assign v_13525 = v_978 & ~v_1072;
assign v_13527 = v_816 & v_13526;
assign v_13528 = v_832 & ~v_922;
assign v_13530 = v_561 & v_13529;
assign v_13531 = v_715 & ~v_793;
assign v_13544 = v_563 & v_13543;
assign v_13545 = v_9609 & v_9784;
assign v_13546 = v_9637 & v_9652;
assign v_13548 = v_9467 & v_13547;
assign v_13549 = v_9482 & v_9494;
assign v_13551 = v_9317 & v_13550;
assign v_13552 = v_9344 & v_9362;
assign v_13554 = v_9179 & v_13553;
assign v_13555 = v_9194 & v_9206;
assign v_13557 = v_9035 & v_13556;
assign v_13558 = v_9059 & v_9074;
assign v_13560 = v_8897 & v_13559;
assign v_13561 = v_8912 & v_8924;
assign v_13563 = v_8740 & v_13562;
assign v_13564 = v_8771 & v_8792;
assign v_13566 = v_8601 & v_13565;
assign v_13567 = v_8616 & v_8628;
assign v_13569 = v_8456 & v_13568;
assign v_13570 = v_8481 & v_8496;
assign v_13572 = v_8317 & v_13571;
assign v_13573 = v_8332 & v_8344;
assign v_13575 = v_8167 & v_13574;
assign v_13576 = v_8194 & v_8212;
assign v_13578 = v_8029 & v_13577;
assign v_13579 = v_8044 & v_8056;
assign v_13581 = v_7885 & v_13580;
assign v_13582 = v_7909 & v_7924;
assign v_13584 = v_7747 & v_13583;
assign v_13585 = v_7762 & v_7774;
assign v_13587 = v_7583 & v_13586;
assign v_13588 = v_7618 & v_7642;
assign v_13590 = v_7443 & v_13589;
assign v_13591 = v_7458 & v_7470;
assign v_13593 = v_7297 & v_13592;
assign v_13594 = v_7323 & v_7338;
assign v_13596 = v_7157 & v_13595;
assign v_13597 = v_7172 & v_7184;
assign v_13599 = v_7007 & v_13598;
assign v_13600 = v_7034 & v_7052;
assign v_13602 = v_6869 & v_13601;
assign v_13603 = v_6884 & v_6896;
assign v_13605 = v_6725 & v_13604;
assign v_13606 = v_6749 & v_6764;
assign v_13608 = v_6587 & v_13607;
assign v_13609 = v_6602 & v_6614;
assign v_13611 = v_6430 & v_13610;
assign v_13612 = v_6461 & v_6482;
assign v_13614 = v_6291 & v_13613;
assign v_13615 = v_6306 & v_6318;
assign v_13617 = v_6146 & v_13616;
assign v_13618 = v_6171 & v_6186;
assign v_13620 = v_6007 & v_13619;
assign v_13621 = v_6022 & v_6034;
assign v_13623 = v_5857 & v_13622;
assign v_13624 = v_5884 & v_5902;
assign v_13626 = v_5719 & v_13625;
assign v_13627 = v_5734 & v_5746;
assign v_13629 = v_5575 & v_13628;
assign v_13630 = v_5599 & v_5614;
assign v_13632 = v_5437 & v_13631;
assign v_13633 = v_5452 & v_5464;
assign v_13635 = v_5266 & v_13634;
assign v_13636 = v_5305 & v_5332;
assign v_13638 = v_5125 & v_13637;
assign v_13639 = v_5140 & v_5152;
assign v_13641 = v_4978 & v_13640;
assign v_13642 = v_5005 & v_5020;
assign v_13644 = v_4837 & v_13643;
assign v_13645 = v_4852 & v_4864;
assign v_13647 = v_4687 & v_13646;
assign v_13648 = v_4714 & v_4732;
assign v_13650 = v_4549 & v_13649;
assign v_13651 = v_4564 & v_4576;
assign v_13653 = v_4405 & v_13652;
assign v_13654 = v_4429 & v_4444;
assign v_13656 = v_4267 & v_13655;
assign v_13657 = v_4282 & v_4294;
assign v_13659 = v_4110 & v_13658;
assign v_13660 = v_4141 & v_4162;
assign v_13662 = v_3971 & v_13661;
assign v_13663 = v_3986 & v_3998;
assign v_13665 = v_3826 & v_13664;
assign v_13666 = v_3851 & v_3866;
assign v_13668 = v_3687 & v_13667;
assign v_13669 = v_3702 & v_3714;
assign v_13671 = v_3537 & v_13670;
assign v_13672 = v_3564 & v_3582;
assign v_13674 = v_3399 & v_13673;
assign v_13675 = v_3414 & v_3426;
assign v_13677 = v_3255 & v_13676;
assign v_13678 = v_3279 & v_3294;
assign v_13680 = v_3117 & v_13679;
assign v_13681 = v_3132 & v_3144;
assign v_13683 = v_2953 & v_13682;
assign v_13684 = v_2988 & v_3012;
assign v_13686 = v_2813 & v_13685;
assign v_13687 = v_2828 & v_2840;
assign v_13689 = v_2667 & v_13688;
assign v_13690 = v_2693 & v_2708;
assign v_13692 = v_2527 & v_13691;
assign v_13693 = v_2542 & v_2554;
assign v_13695 = v_2377 & v_13694;
assign v_13696 = v_2404 & v_2422;
assign v_13698 = v_2239 & v_13697;
assign v_13699 = v_2254 & v_2266;
assign v_13701 = v_2095 & v_13700;
assign v_13702 = v_2119 & v_2134;
assign v_13704 = v_1957 & v_13703;
assign v_13705 = v_1972 & v_1984;
assign v_13707 = v_1800 & v_13706;
assign v_13708 = v_1831 & v_1852;
assign v_13710 = v_1661 & v_13709;
assign v_13711 = v_1676 & v_1688;
assign v_13713 = v_1516 & v_13712;
assign v_13714 = v_1541 & v_1556;
assign v_13716 = v_1377 & v_13715;
assign v_13717 = v_1392 & v_1404;
assign v_13719 = v_1227 & v_13718;
assign v_13720 = v_1254 & v_1272;
assign v_13722 = v_1089 & v_13721;
assign v_13723 = v_1104 & v_1116;
assign v_13725 = v_945 & v_13724;
assign v_13726 = v_969 & v_984;
assign v_13728 = v_810 & v_13727;
assign v_13729 = v_826 & v_838;
assign v_13731 = v_223 & v_13730;
assign v_13732 = v_626 & v_721;
assign v_13734 = v_9609 & v_9753;
assign v_13735 = v_9604 & v_9637;
assign v_13737 = v_9467 & v_13736;
assign v_13738 = v_9463 & v_9482;
assign v_13740 = v_9317 & v_13739;
assign v_13741 = v_9311 & v_9344;
assign v_13743 = v_9179 & v_13742;
assign v_13744 = v_9175 & v_9194;
assign v_13746 = v_9035 & v_13745;
assign v_13747 = v_9030 & v_9059;
assign v_13749 = v_8897 & v_13748;
assign v_13750 = v_8893 & v_8912;
assign v_13752 = v_8740 & v_13751;
assign v_13753 = v_8733 & v_8771;
assign v_13755 = v_8601 & v_13754;
assign v_13756 = v_8597 & v_8616;
assign v_13758 = v_8456 & v_13757;
assign v_13759 = v_8451 & v_8481;
assign v_13761 = v_8317 & v_13760;
assign v_13762 = v_8313 & v_8332;
assign v_13764 = v_8167 & v_13763;
assign v_13765 = v_8161 & v_8194;
assign v_13767 = v_8029 & v_13766;
assign v_13768 = v_8025 & v_8044;
assign v_13770 = v_7885 & v_13769;
assign v_13771 = v_7880 & v_7909;
assign v_13773 = v_7747 & v_13772;
assign v_13774 = v_7743 & v_7762;
assign v_13776 = v_7583 & v_13775;
assign v_13777 = v_7575 & v_7618;
assign v_13779 = v_7443 & v_13778;
assign v_13780 = v_7439 & v_7458;
assign v_13782 = v_7297 & v_13781;
assign v_13783 = v_7292 & v_7323;
assign v_13785 = v_7157 & v_13784;
assign v_13786 = v_7153 & v_7172;
assign v_13788 = v_7007 & v_13787;
assign v_13789 = v_7001 & v_7034;
assign v_13791 = v_6869 & v_13790;
assign v_13792 = v_6865 & v_6884;
assign v_13794 = v_6725 & v_13793;
assign v_13795 = v_6720 & v_6749;
assign v_13797 = v_6587 & v_13796;
assign v_13798 = v_6583 & v_6602;
assign v_13800 = v_6430 & v_13799;
assign v_13801 = v_6423 & v_6461;
assign v_13803 = v_6291 & v_13802;
assign v_13804 = v_6287 & v_6306;
assign v_13806 = v_6146 & v_13805;
assign v_13807 = v_6141 & v_6171;
assign v_13809 = v_6007 & v_13808;
assign v_13810 = v_6003 & v_6022;
assign v_13812 = v_5857 & v_13811;
assign v_13813 = v_5851 & v_5884;
assign v_13815 = v_5719 & v_13814;
assign v_13816 = v_5715 & v_5734;
assign v_13818 = v_5575 & v_13817;
assign v_13819 = v_5570 & v_5599;
assign v_13821 = v_5437 & v_13820;
assign v_13822 = v_5433 & v_5452;
assign v_13824 = v_5266 & v_13823;
assign v_13825 = v_5257 & v_5305;
assign v_13827 = v_5125 & v_13826;
assign v_13828 = v_5121 & v_5140;
assign v_13830 = v_4978 & v_13829;
assign v_13831 = v_4973 & v_5005;
assign v_13833 = v_4837 & v_13832;
assign v_13834 = v_4833 & v_4852;
assign v_13836 = v_4687 & v_13835;
assign v_13837 = v_4681 & v_4714;
assign v_13839 = v_4549 & v_13838;
assign v_13840 = v_4545 & v_4564;
assign v_13842 = v_4405 & v_13841;
assign v_13843 = v_4400 & v_4429;
assign v_13845 = v_4267 & v_13844;
assign v_13846 = v_4263 & v_4282;
assign v_13848 = v_4110 & v_13847;
assign v_13849 = v_4103 & v_4141;
assign v_13851 = v_3971 & v_13850;
assign v_13852 = v_3967 & v_3986;
assign v_13854 = v_3826 & v_13853;
assign v_13855 = v_3821 & v_3851;
assign v_13857 = v_3687 & v_13856;
assign v_13858 = v_3683 & v_3702;
assign v_13860 = v_3537 & v_13859;
assign v_13861 = v_3531 & v_3564;
assign v_13863 = v_3399 & v_13862;
assign v_13864 = v_3395 & v_3414;
assign v_13866 = v_3255 & v_13865;
assign v_13867 = v_3250 & v_3279;
assign v_13869 = v_3117 & v_13868;
assign v_13870 = v_3113 & v_3132;
assign v_13872 = v_2953 & v_13871;
assign v_13873 = v_2945 & v_2988;
assign v_13875 = v_2813 & v_13874;
assign v_13876 = v_2809 & v_2828;
assign v_13878 = v_2667 & v_13877;
assign v_13879 = v_2662 & v_2693;
assign v_13881 = v_2527 & v_13880;
assign v_13882 = v_2523 & v_2542;
assign v_13884 = v_2377 & v_13883;
assign v_13885 = v_2371 & v_2404;
assign v_13887 = v_2239 & v_13886;
assign v_13888 = v_2235 & v_2254;
assign v_13890 = v_2095 & v_13889;
assign v_13891 = v_2090 & v_2119;
assign v_13893 = v_1957 & v_13892;
assign v_13894 = v_1953 & v_1972;
assign v_13896 = v_1800 & v_13895;
assign v_13897 = v_1793 & v_1831;
assign v_13899 = v_1661 & v_13898;
assign v_13900 = v_1657 & v_1676;
assign v_13902 = v_1516 & v_13901;
assign v_13903 = v_1511 & v_1541;
assign v_13905 = v_1377 & v_13904;
assign v_13906 = v_1373 & v_1392;
assign v_13908 = v_1227 & v_13907;
assign v_13909 = v_1221 & v_1254;
assign v_13911 = v_1089 & v_13910;
assign v_13912 = v_1085 & v_1104;
assign v_13914 = v_945 & v_13913;
assign v_13915 = v_940 & v_969;
assign v_13917 = v_810 & v_13916;
assign v_13918 = v_804 & v_826;
assign v_13920 = v_223 & v_13919;
assign v_13921 = v_98 & v_626;
assign v_13924 = v_9609 & v_9796;
assign v_13925 = v_9637 & v_9664;
assign v_13927 = v_9467 & v_13926;
assign v_13928 = v_9482 & v_9506;
assign v_13930 = v_9317 & v_13929;
assign v_13931 = v_9344 & v_9374;
assign v_13933 = v_9179 & v_13932;
assign v_13934 = v_9194 & v_9218;
assign v_13936 = v_9035 & v_13935;
assign v_13937 = v_9059 & v_9086;
assign v_13939 = v_8897 & v_13938;
assign v_13940 = v_8912 & v_8936;
assign v_13942 = v_8740 & v_13941;
assign v_13943 = v_8771 & v_8804;
assign v_13945 = v_8601 & v_13944;
assign v_13946 = v_8616 & v_8640;
assign v_13948 = v_8456 & v_13947;
assign v_13949 = v_8481 & v_8508;
assign v_13951 = v_8317 & v_13950;
assign v_13952 = v_8332 & v_8356;
assign v_13954 = v_8167 & v_13953;
assign v_13955 = v_8194 & v_8224;
assign v_13957 = v_8029 & v_13956;
assign v_13958 = v_8044 & v_8068;
assign v_13960 = v_7885 & v_13959;
assign v_13961 = v_7909 & v_7936;
assign v_13963 = v_7747 & v_13962;
assign v_13964 = v_7762 & v_7786;
assign v_13966 = v_7583 & v_13965;
assign v_13967 = v_7618 & v_7654;
assign v_13969 = v_7443 & v_13968;
assign v_13970 = v_7458 & v_7482;
assign v_13972 = v_7297 & v_13971;
assign v_13973 = v_7323 & v_7350;
assign v_13975 = v_7157 & v_13974;
assign v_13976 = v_7172 & v_7196;
assign v_13978 = v_7007 & v_13977;
assign v_13979 = v_7034 & v_7064;
assign v_13981 = v_6869 & v_13980;
assign v_13982 = v_6884 & v_6908;
assign v_13984 = v_6725 & v_13983;
assign v_13985 = v_6749 & v_6776;
assign v_13987 = v_6587 & v_13986;
assign v_13988 = v_6602 & v_6626;
assign v_13990 = v_6430 & v_13989;
assign v_13991 = v_6461 & v_6494;
assign v_13993 = v_6291 & v_13992;
assign v_13994 = v_6306 & v_6330;
assign v_13996 = v_6146 & v_13995;
assign v_13997 = v_6171 & v_6198;
assign v_13999 = v_6007 & v_13998;
assign v_14000 = v_6022 & v_6046;
assign v_14002 = v_5857 & v_14001;
assign v_14003 = v_5884 & v_5914;
assign v_14005 = v_5719 & v_14004;
assign v_14006 = v_5734 & v_5758;
assign v_14008 = v_5575 & v_14007;
assign v_14009 = v_5599 & v_5626;
assign v_14011 = v_5437 & v_14010;
assign v_14012 = v_5452 & v_5476;
assign v_14014 = v_5266 & v_14013;
assign v_14015 = v_5305 & v_5344;
assign v_14017 = v_5125 & v_14016;
assign v_14018 = v_5140 & v_5164;
assign v_14020 = v_4978 & v_14019;
assign v_14021 = v_5005 & v_5032;
assign v_14023 = v_4837 & v_14022;
assign v_14024 = v_4852 & v_4876;
assign v_14026 = v_4687 & v_14025;
assign v_14027 = v_4714 & v_4744;
assign v_14029 = v_4549 & v_14028;
assign v_14030 = v_4564 & v_4588;
assign v_14032 = v_4405 & v_14031;
assign v_14033 = v_4429 & v_4456;
assign v_14035 = v_4267 & v_14034;
assign v_14036 = v_4282 & v_4306;
assign v_14038 = v_4110 & v_14037;
assign v_14039 = v_4141 & v_4174;
assign v_14041 = v_3971 & v_14040;
assign v_14042 = v_3986 & v_4010;
assign v_14044 = v_3826 & v_14043;
assign v_14045 = v_3851 & v_3878;
assign v_14047 = v_3687 & v_14046;
assign v_14048 = v_3702 & v_3726;
assign v_14050 = v_3537 & v_14049;
assign v_14051 = v_3564 & v_3594;
assign v_14053 = v_3399 & v_14052;
assign v_14054 = v_3414 & v_3438;
assign v_14056 = v_3255 & v_14055;
assign v_14057 = v_3279 & v_3306;
assign v_14059 = v_3117 & v_14058;
assign v_14060 = v_3132 & v_3156;
assign v_14062 = v_2953 & v_14061;
assign v_14063 = v_2988 & v_3024;
assign v_14065 = v_2813 & v_14064;
assign v_14066 = v_2828 & v_2852;
assign v_14068 = v_2667 & v_14067;
assign v_14069 = v_2693 & v_2720;
assign v_14071 = v_2527 & v_14070;
assign v_14072 = v_2542 & v_2566;
assign v_14074 = v_2377 & v_14073;
assign v_14075 = v_2404 & v_2434;
assign v_14077 = v_2239 & v_14076;
assign v_14078 = v_2254 & v_2278;
assign v_14080 = v_2095 & v_14079;
assign v_14081 = v_2119 & v_2146;
assign v_14083 = v_1957 & v_14082;
assign v_14084 = v_1972 & v_1996;
assign v_14086 = v_1800 & v_14085;
assign v_14087 = v_1831 & v_1864;
assign v_14089 = v_1661 & v_14088;
assign v_14090 = v_1676 & v_1700;
assign v_14092 = v_1516 & v_14091;
assign v_14093 = v_1541 & v_1568;
assign v_14095 = v_1377 & v_14094;
assign v_14096 = v_1392 & v_1416;
assign v_14098 = v_1227 & v_14097;
assign v_14099 = v_1254 & v_1284;
assign v_14101 = v_1089 & v_14100;
assign v_14102 = v_1104 & v_1128;
assign v_14104 = v_945 & v_14103;
assign v_14105 = v_969 & v_996;
assign v_14107 = v_810 & v_14106;
assign v_14108 = v_826 & v_850;
assign v_14110 = v_223 & v_14109;
assign v_14111 = v_626 & v_731;
assign v_14114 = v_9609 & v_9808;
assign v_14115 = v_9637 & v_9676;
assign v_14117 = v_9467 & v_14116;
assign v_14118 = v_9482 & v_9518;
assign v_14120 = v_9317 & v_14119;
assign v_14121 = v_9344 & v_9386;
assign v_14123 = v_9179 & v_14122;
assign v_14124 = v_9194 & v_9230;
assign v_14126 = v_9035 & v_14125;
assign v_14127 = v_9059 & v_9098;
assign v_14129 = v_8897 & v_14128;
assign v_14130 = v_8912 & v_8948;
assign v_14132 = v_8740 & v_14131;
assign v_14133 = v_8771 & v_8816;
assign v_14135 = v_8601 & v_14134;
assign v_14136 = v_8616 & v_8652;
assign v_14138 = v_8456 & v_14137;
assign v_14139 = v_8481 & v_8520;
assign v_14141 = v_8317 & v_14140;
assign v_14142 = v_8332 & v_8368;
assign v_14144 = v_8167 & v_14143;
assign v_14145 = v_8194 & v_8236;
assign v_14147 = v_8029 & v_14146;
assign v_14148 = v_8044 & v_8080;
assign v_14150 = v_7885 & v_14149;
assign v_14151 = v_7909 & v_7948;
assign v_14153 = v_7747 & v_14152;
assign v_14154 = v_7762 & v_7798;
assign v_14156 = v_7583 & v_14155;
assign v_14157 = v_7618 & v_7666;
assign v_14159 = v_7443 & v_14158;
assign v_14160 = v_7458 & v_7494;
assign v_14162 = v_7297 & v_14161;
assign v_14163 = v_7323 & v_7362;
assign v_14165 = v_7157 & v_14164;
assign v_14166 = v_7172 & v_7208;
assign v_14168 = v_7007 & v_14167;
assign v_14169 = v_7034 & v_7076;
assign v_14171 = v_6869 & v_14170;
assign v_14172 = v_6884 & v_6920;
assign v_14174 = v_6725 & v_14173;
assign v_14175 = v_6749 & v_6788;
assign v_14177 = v_6587 & v_14176;
assign v_14178 = v_6602 & v_6638;
assign v_14180 = v_6430 & v_14179;
assign v_14181 = v_6461 & v_6506;
assign v_14183 = v_6291 & v_14182;
assign v_14184 = v_6306 & v_6342;
assign v_14186 = v_6146 & v_14185;
assign v_14187 = v_6171 & v_6210;
assign v_14189 = v_6007 & v_14188;
assign v_14190 = v_6022 & v_6058;
assign v_14192 = v_5857 & v_14191;
assign v_14193 = v_5884 & v_5926;
assign v_14195 = v_5719 & v_14194;
assign v_14196 = v_5734 & v_5770;
assign v_14198 = v_5575 & v_14197;
assign v_14199 = v_5599 & v_5638;
assign v_14201 = v_5437 & v_14200;
assign v_14202 = v_5452 & v_5488;
assign v_14204 = v_5266 & v_14203;
assign v_14205 = v_5305 & v_5356;
assign v_14207 = v_5125 & v_14206;
assign v_14208 = v_5140 & v_5176;
assign v_14210 = v_4978 & v_14209;
assign v_14211 = v_5005 & v_5044;
assign v_14213 = v_4837 & v_14212;
assign v_14214 = v_4852 & v_4888;
assign v_14216 = v_4687 & v_14215;
assign v_14217 = v_4714 & v_4756;
assign v_14219 = v_4549 & v_14218;
assign v_14220 = v_4564 & v_4600;
assign v_14222 = v_4405 & v_14221;
assign v_14223 = v_4429 & v_4468;
assign v_14225 = v_4267 & v_14224;
assign v_14226 = v_4282 & v_4318;
assign v_14228 = v_4110 & v_14227;
assign v_14229 = v_4141 & v_4186;
assign v_14231 = v_3971 & v_14230;
assign v_14232 = v_3986 & v_4022;
assign v_14234 = v_3826 & v_14233;
assign v_14235 = v_3851 & v_3890;
assign v_14237 = v_3687 & v_14236;
assign v_14238 = v_3702 & v_3738;
assign v_14240 = v_3537 & v_14239;
assign v_14241 = v_3564 & v_3606;
assign v_14243 = v_3399 & v_14242;
assign v_14244 = v_3414 & v_3450;
assign v_14246 = v_3255 & v_14245;
assign v_14247 = v_3279 & v_3318;
assign v_14249 = v_3117 & v_14248;
assign v_14250 = v_3132 & v_3168;
assign v_14252 = v_2953 & v_14251;
assign v_14253 = v_2988 & v_3036;
assign v_14255 = v_2813 & v_14254;
assign v_14256 = v_2828 & v_2864;
assign v_14258 = v_2667 & v_14257;
assign v_14259 = v_2693 & v_2732;
assign v_14261 = v_2527 & v_14260;
assign v_14262 = v_2542 & v_2578;
assign v_14264 = v_2377 & v_14263;
assign v_14265 = v_2404 & v_2446;
assign v_14267 = v_2239 & v_14266;
assign v_14268 = v_2254 & v_2290;
assign v_14270 = v_2095 & v_14269;
assign v_14271 = v_2119 & v_2158;
assign v_14273 = v_1957 & v_14272;
assign v_14274 = v_1972 & v_2008;
assign v_14276 = v_1800 & v_14275;
assign v_14277 = v_1831 & v_1876;
assign v_14279 = v_1661 & v_14278;
assign v_14280 = v_1676 & v_1712;
assign v_14282 = v_1516 & v_14281;
assign v_14283 = v_1541 & v_1580;
assign v_14285 = v_1377 & v_14284;
assign v_14286 = v_1392 & v_1428;
assign v_14288 = v_1227 & v_14287;
assign v_14289 = v_1254 & v_1296;
assign v_14291 = v_1089 & v_14290;
assign v_14292 = v_1104 & v_1140;
assign v_14294 = v_945 & v_14293;
assign v_14295 = v_969 & v_1008;
assign v_14297 = v_810 & v_14296;
assign v_14298 = v_826 & v_862;
assign v_14300 = v_223 & v_14299;
assign v_14301 = v_626 & v_741;
assign v_14304 = v_9609 & v_9820;
assign v_14305 = v_9637 & v_9688;
assign v_14307 = v_9467 & v_14306;
assign v_14308 = v_9482 & v_9530;
assign v_14310 = v_9317 & v_14309;
assign v_14311 = v_9344 & v_9398;
assign v_14313 = v_9179 & v_14312;
assign v_14314 = v_9194 & v_9242;
assign v_14316 = v_9035 & v_14315;
assign v_14317 = v_9059 & v_9110;
assign v_14319 = v_8897 & v_14318;
assign v_14320 = v_8912 & v_8960;
assign v_14322 = v_8740 & v_14321;
assign v_14323 = v_8771 & v_8828;
assign v_14325 = v_8601 & v_14324;
assign v_14326 = v_8616 & v_8664;
assign v_14328 = v_8456 & v_14327;
assign v_14329 = v_8481 & v_8532;
assign v_14331 = v_8317 & v_14330;
assign v_14332 = v_8332 & v_8380;
assign v_14334 = v_8167 & v_14333;
assign v_14335 = v_8194 & v_8248;
assign v_14337 = v_8029 & v_14336;
assign v_14338 = v_8044 & v_8092;
assign v_14340 = v_7885 & v_14339;
assign v_14341 = v_7909 & v_7960;
assign v_14343 = v_7747 & v_14342;
assign v_14344 = v_7762 & v_7810;
assign v_14346 = v_7583 & v_14345;
assign v_14347 = v_7618 & v_7678;
assign v_14349 = v_7443 & v_14348;
assign v_14350 = v_7458 & v_7506;
assign v_14352 = v_7297 & v_14351;
assign v_14353 = v_7323 & v_7374;
assign v_14355 = v_7157 & v_14354;
assign v_14356 = v_7172 & v_7220;
assign v_14358 = v_7007 & v_14357;
assign v_14359 = v_7034 & v_7088;
assign v_14361 = v_6869 & v_14360;
assign v_14362 = v_6884 & v_6932;
assign v_14364 = v_6725 & v_14363;
assign v_14365 = v_6749 & v_6800;
assign v_14367 = v_6587 & v_14366;
assign v_14368 = v_6602 & v_6650;
assign v_14370 = v_6430 & v_14369;
assign v_14371 = v_6461 & v_6518;
assign v_14373 = v_6291 & v_14372;
assign v_14374 = v_6306 & v_6354;
assign v_14376 = v_6146 & v_14375;
assign v_14377 = v_6171 & v_6222;
assign v_14379 = v_6007 & v_14378;
assign v_14380 = v_6022 & v_6070;
assign v_14382 = v_5857 & v_14381;
assign v_14383 = v_5884 & v_5938;
assign v_14385 = v_5719 & v_14384;
assign v_14386 = v_5734 & v_5782;
assign v_14388 = v_5575 & v_14387;
assign v_14389 = v_5599 & v_5650;
assign v_14391 = v_5437 & v_14390;
assign v_14392 = v_5452 & v_5500;
assign v_14394 = v_5266 & v_14393;
assign v_14395 = v_5305 & v_5368;
assign v_14397 = v_5125 & v_14396;
assign v_14398 = v_5140 & v_5188;
assign v_14400 = v_4978 & v_14399;
assign v_14401 = v_5005 & v_5056;
assign v_14403 = v_4837 & v_14402;
assign v_14404 = v_4852 & v_4900;
assign v_14406 = v_4687 & v_14405;
assign v_14407 = v_4714 & v_4768;
assign v_14409 = v_4549 & v_14408;
assign v_14410 = v_4564 & v_4612;
assign v_14412 = v_4405 & v_14411;
assign v_14413 = v_4429 & v_4480;
assign v_14415 = v_4267 & v_14414;
assign v_14416 = v_4282 & v_4330;
assign v_14418 = v_4110 & v_14417;
assign v_14419 = v_4141 & v_4198;
assign v_14421 = v_3971 & v_14420;
assign v_14422 = v_3986 & v_4034;
assign v_14424 = v_3826 & v_14423;
assign v_14425 = v_3851 & v_3902;
assign v_14427 = v_3687 & v_14426;
assign v_14428 = v_3702 & v_3750;
assign v_14430 = v_3537 & v_14429;
assign v_14431 = v_3564 & v_3618;
assign v_14433 = v_3399 & v_14432;
assign v_14434 = v_3414 & v_3462;
assign v_14436 = v_3255 & v_14435;
assign v_14437 = v_3279 & v_3330;
assign v_14439 = v_3117 & v_14438;
assign v_14440 = v_3132 & v_3180;
assign v_14442 = v_2953 & v_14441;
assign v_14443 = v_2988 & v_3048;
assign v_14445 = v_2813 & v_14444;
assign v_14446 = v_2828 & v_2876;
assign v_14448 = v_2667 & v_14447;
assign v_14449 = v_2693 & v_2744;
assign v_14451 = v_2527 & v_14450;
assign v_14452 = v_2542 & v_2590;
assign v_14454 = v_2377 & v_14453;
assign v_14455 = v_2404 & v_2458;
assign v_14457 = v_2239 & v_14456;
assign v_14458 = v_2254 & v_2302;
assign v_14460 = v_2095 & v_14459;
assign v_14461 = v_2119 & v_2170;
assign v_14463 = v_1957 & v_14462;
assign v_14464 = v_1972 & v_2020;
assign v_14466 = v_1800 & v_14465;
assign v_14467 = v_1831 & v_1888;
assign v_14469 = v_1661 & v_14468;
assign v_14470 = v_1676 & v_1724;
assign v_14472 = v_1516 & v_14471;
assign v_14473 = v_1541 & v_1592;
assign v_14475 = v_1377 & v_14474;
assign v_14476 = v_1392 & v_1440;
assign v_14478 = v_1227 & v_14477;
assign v_14479 = v_1254 & v_1308;
assign v_14481 = v_1089 & v_14480;
assign v_14482 = v_1104 & v_1152;
assign v_14484 = v_945 & v_14483;
assign v_14485 = v_969 & v_1020;
assign v_14487 = v_810 & v_14486;
assign v_14488 = v_826 & v_874;
assign v_14490 = v_223 & v_14489;
assign v_14491 = v_626 & v_751;
assign v_14494 = v_9609 & v_9832;
assign v_14495 = v_9637 & v_9700;
assign v_14497 = v_9467 & v_14496;
assign v_14498 = v_9482 & v_9542;
assign v_14500 = v_9317 & v_14499;
assign v_14501 = v_9344 & v_9410;
assign v_14503 = v_9179 & v_14502;
assign v_14504 = v_9194 & v_9254;
assign v_14506 = v_9035 & v_14505;
assign v_14507 = v_9059 & v_9122;
assign v_14509 = v_8897 & v_14508;
assign v_14510 = v_8912 & v_8972;
assign v_14512 = v_8740 & v_14511;
assign v_14513 = v_8771 & v_8840;
assign v_14515 = v_8601 & v_14514;
assign v_14516 = v_8616 & v_8676;
assign v_14518 = v_8456 & v_14517;
assign v_14519 = v_8481 & v_8544;
assign v_14521 = v_8317 & v_14520;
assign v_14522 = v_8332 & v_8392;
assign v_14524 = v_8167 & v_14523;
assign v_14525 = v_8194 & v_8260;
assign v_14527 = v_8029 & v_14526;
assign v_14528 = v_8044 & v_8104;
assign v_14530 = v_7885 & v_14529;
assign v_14531 = v_7909 & v_7972;
assign v_14533 = v_7747 & v_14532;
assign v_14534 = v_7762 & v_7822;
assign v_14536 = v_7583 & v_14535;
assign v_14537 = v_7618 & v_7690;
assign v_14539 = v_7443 & v_14538;
assign v_14540 = v_7458 & v_7518;
assign v_14542 = v_7297 & v_14541;
assign v_14543 = v_7323 & v_7386;
assign v_14545 = v_7157 & v_14544;
assign v_14546 = v_7172 & v_7232;
assign v_14548 = v_7007 & v_14547;
assign v_14549 = v_7034 & v_7100;
assign v_14551 = v_6869 & v_14550;
assign v_14552 = v_6884 & v_6944;
assign v_14554 = v_6725 & v_14553;
assign v_14555 = v_6749 & v_6812;
assign v_14557 = v_6587 & v_14556;
assign v_14558 = v_6602 & v_6662;
assign v_14560 = v_6430 & v_14559;
assign v_14561 = v_6461 & v_6530;
assign v_14563 = v_6291 & v_14562;
assign v_14564 = v_6306 & v_6366;
assign v_14566 = v_6146 & v_14565;
assign v_14567 = v_6171 & v_6234;
assign v_14569 = v_6007 & v_14568;
assign v_14570 = v_6022 & v_6082;
assign v_14572 = v_5857 & v_14571;
assign v_14573 = v_5884 & v_5950;
assign v_14575 = v_5719 & v_14574;
assign v_14576 = v_5734 & v_5794;
assign v_14578 = v_5575 & v_14577;
assign v_14579 = v_5599 & v_5662;
assign v_14581 = v_5437 & v_14580;
assign v_14582 = v_5452 & v_5512;
assign v_14584 = v_5266 & v_14583;
assign v_14585 = v_5305 & v_5380;
assign v_14587 = v_5125 & v_14586;
assign v_14588 = v_5140 & v_5200;
assign v_14590 = v_4978 & v_14589;
assign v_14591 = v_5005 & v_5068;
assign v_14593 = v_4837 & v_14592;
assign v_14594 = v_4852 & v_4912;
assign v_14596 = v_4687 & v_14595;
assign v_14597 = v_4714 & v_4780;
assign v_14599 = v_4549 & v_14598;
assign v_14600 = v_4564 & v_4624;
assign v_14602 = v_4405 & v_14601;
assign v_14603 = v_4429 & v_4492;
assign v_14605 = v_4267 & v_14604;
assign v_14606 = v_4282 & v_4342;
assign v_14608 = v_4110 & v_14607;
assign v_14609 = v_4141 & v_4210;
assign v_14611 = v_3971 & v_14610;
assign v_14612 = v_3986 & v_4046;
assign v_14614 = v_3826 & v_14613;
assign v_14615 = v_3851 & v_3914;
assign v_14617 = v_3687 & v_14616;
assign v_14618 = v_3702 & v_3762;
assign v_14620 = v_3537 & v_14619;
assign v_14621 = v_3564 & v_3630;
assign v_14623 = v_3399 & v_14622;
assign v_14624 = v_3414 & v_3474;
assign v_14626 = v_3255 & v_14625;
assign v_14627 = v_3279 & v_3342;
assign v_14629 = v_3117 & v_14628;
assign v_14630 = v_3132 & v_3192;
assign v_14632 = v_2953 & v_14631;
assign v_14633 = v_2988 & v_3060;
assign v_14635 = v_2813 & v_14634;
assign v_14636 = v_2828 & v_2888;
assign v_14638 = v_2667 & v_14637;
assign v_14639 = v_2693 & v_2756;
assign v_14641 = v_2527 & v_14640;
assign v_14642 = v_2542 & v_2602;
assign v_14644 = v_2377 & v_14643;
assign v_14645 = v_2404 & v_2470;
assign v_14647 = v_2239 & v_14646;
assign v_14648 = v_2254 & v_2314;
assign v_14650 = v_2095 & v_14649;
assign v_14651 = v_2119 & v_2182;
assign v_14653 = v_1957 & v_14652;
assign v_14654 = v_1972 & v_2032;
assign v_14656 = v_1800 & v_14655;
assign v_14657 = v_1831 & v_1900;
assign v_14659 = v_1661 & v_14658;
assign v_14660 = v_1676 & v_1736;
assign v_14662 = v_1516 & v_14661;
assign v_14663 = v_1541 & v_1604;
assign v_14665 = v_1377 & v_14664;
assign v_14666 = v_1392 & v_1452;
assign v_14668 = v_1227 & v_14667;
assign v_14669 = v_1254 & v_1320;
assign v_14671 = v_1089 & v_14670;
assign v_14672 = v_1104 & v_1164;
assign v_14674 = v_945 & v_14673;
assign v_14675 = v_969 & v_1032;
assign v_14677 = v_810 & v_14676;
assign v_14678 = v_826 & v_886;
assign v_14680 = v_223 & v_14679;
assign v_14681 = v_626 & v_761;
assign v_14684 = v_9609 & v_9844;
assign v_14685 = v_9637 & v_9712;
assign v_14687 = v_9467 & v_14686;
assign v_14688 = v_9482 & v_9554;
assign v_14690 = v_9317 & v_14689;
assign v_14691 = v_9344 & v_9422;
assign v_14693 = v_9179 & v_14692;
assign v_14694 = v_9194 & v_9266;
assign v_14696 = v_9035 & v_14695;
assign v_14697 = v_9059 & v_9134;
assign v_14699 = v_8897 & v_14698;
assign v_14700 = v_8912 & v_8984;
assign v_14702 = v_8740 & v_14701;
assign v_14703 = v_8771 & v_8852;
assign v_14705 = v_8601 & v_14704;
assign v_14706 = v_8616 & v_8688;
assign v_14708 = v_8456 & v_14707;
assign v_14709 = v_8481 & v_8556;
assign v_14711 = v_8317 & v_14710;
assign v_14712 = v_8332 & v_8404;
assign v_14714 = v_8167 & v_14713;
assign v_14715 = v_8194 & v_8272;
assign v_14717 = v_8029 & v_14716;
assign v_14718 = v_8044 & v_8116;
assign v_14720 = v_7885 & v_14719;
assign v_14721 = v_7909 & v_7984;
assign v_14723 = v_7747 & v_14722;
assign v_14724 = v_7762 & v_7834;
assign v_14726 = v_7583 & v_14725;
assign v_14727 = v_7618 & v_7702;
assign v_14729 = v_7443 & v_14728;
assign v_14730 = v_7458 & v_7530;
assign v_14732 = v_7297 & v_14731;
assign v_14733 = v_7323 & v_7398;
assign v_14735 = v_7157 & v_14734;
assign v_14736 = v_7172 & v_7244;
assign v_14738 = v_7007 & v_14737;
assign v_14739 = v_7034 & v_7112;
assign v_14741 = v_6869 & v_14740;
assign v_14742 = v_6884 & v_6956;
assign v_14744 = v_6725 & v_14743;
assign v_14745 = v_6749 & ~v_6824;
assign v_14747 = v_6587 & v_14746;
assign v_14748 = v_6602 & v_6674;
assign v_14750 = v_6430 & v_14749;
assign v_14751 = v_6461 & v_6542;
assign v_14753 = v_6291 & v_14752;
assign v_14754 = v_6306 & v_6378;
assign v_14756 = v_6146 & v_14755;
assign v_14757 = v_6171 & v_6246;
assign v_14759 = v_6007 & v_14758;
assign v_14760 = v_6022 & ~v_6094;
assign v_14762 = v_5857 & v_14761;
assign v_14763 = v_5884 & v_5962;
assign v_14765 = v_5719 & v_14764;
assign v_14766 = v_5734 & ~v_5806;
assign v_14768 = v_5575 & v_14767;
assign v_14769 = v_5599 & v_5674;
assign v_14771 = v_5437 & v_14770;
assign v_14772 = v_5452 & v_5524;
assign v_14774 = v_5266 & v_14773;
assign v_14775 = v_5305 & v_5392;
assign v_14777 = v_5125 & v_14776;
assign v_14778 = v_5140 & v_5212;
assign v_14780 = v_4978 & v_14779;
assign v_14781 = v_5005 & v_5080;
assign v_14783 = v_4837 & v_14782;
assign v_14784 = v_4852 & v_4924;
assign v_14786 = v_4687 & v_14785;
assign v_14787 = v_4714 & v_4792;
assign v_14789 = v_4549 & v_14788;
assign v_14790 = v_4564 & v_4636;
assign v_14792 = v_4405 & v_14791;
assign v_14793 = v_4429 & v_4504;
assign v_14795 = v_4267 & v_14794;
assign v_14796 = v_4282 & v_4354;
assign v_14798 = v_4110 & v_14797;
assign v_14799 = v_4141 & v_4222;
assign v_14801 = v_3971 & v_14800;
assign v_14802 = v_3986 & v_4058;
assign v_14804 = v_3826 & v_14803;
assign v_14805 = v_3851 & v_3926;
assign v_14807 = v_3687 & v_14806;
assign v_14808 = v_3702 & v_3774;
assign v_14810 = v_3537 & v_14809;
assign v_14811 = v_3564 & v_3642;
assign v_14813 = v_3399 & v_14812;
assign v_14814 = v_3414 & v_3486;
assign v_14816 = v_3255 & v_14815;
assign v_14817 = v_3279 & v_3354;
assign v_14819 = v_3117 & v_14818;
assign v_14820 = v_3132 & ~v_3204;
assign v_14822 = v_2953 & v_14821;
assign v_14823 = v_2988 & v_3072;
assign v_14825 = v_2813 & v_14824;
assign v_14826 = v_2828 & v_2900;
assign v_14828 = v_2667 & v_14827;
assign v_14829 = v_2693 & v_2768;
assign v_14831 = v_2527 & v_14830;
assign v_14832 = v_2542 & v_2614;
assign v_14834 = v_2377 & v_14833;
assign v_14835 = v_2404 & v_2482;
assign v_14837 = v_2239 & v_14836;
assign v_14838 = v_2254 & v_2326;
assign v_14840 = v_2095 & v_14839;
assign v_14841 = v_2119 & v_2194;
assign v_14843 = v_1957 & v_14842;
assign v_14844 = v_1972 & v_2044;
assign v_14846 = v_1800 & v_14845;
assign v_14847 = v_1831 & v_1912;
assign v_14849 = v_1661 & v_14848;
assign v_14850 = v_1676 & v_1748;
assign v_14852 = v_1516 & v_14851;
assign v_14853 = v_1541 & v_1616;
assign v_14855 = v_1377 & v_14854;
assign v_14856 = v_1392 & v_1464;
assign v_14858 = v_1227 & v_14857;
assign v_14859 = v_1254 & v_1332;
assign v_14861 = v_1089 & v_14860;
assign v_14862 = v_1104 & v_1176;
assign v_14864 = v_945 & v_14863;
assign v_14865 = v_969 & v_1044;
assign v_14867 = v_810 & v_14866;
assign v_14868 = v_826 & v_898;
assign v_14870 = v_223 & v_14869;
assign v_14871 = v_626 & v_771;
assign v_14874 = v_9609 & ~v_9872;
assign v_14875 = v_9637 & ~v_9740;
assign v_14877 = v_9467 & v_14876;
assign v_14878 = v_9482 & ~v_9582;
assign v_14880 = v_9317 & v_14879;
assign v_14881 = v_9344 & ~v_9450;
assign v_14883 = v_9179 & v_14882;
assign v_14884 = v_9194 & ~v_9294;
assign v_14886 = v_9035 & v_14885;
assign v_14887 = v_9059 & ~v_9162;
assign v_14889 = v_8897 & v_14888;
assign v_14890 = v_8912 & ~v_9012;
assign v_14892 = v_8740 & v_14891;
assign v_14893 = v_8771 & ~v_8880;
assign v_14895 = v_8601 & v_14894;
assign v_14896 = v_8616 & ~v_8716;
assign v_14898 = v_8456 & v_14897;
assign v_14899 = v_8481 & ~v_8584;
assign v_14901 = v_8317 & v_14900;
assign v_14902 = v_8332 & v_8432;
assign v_14904 = v_8167 & v_14903;
assign v_14905 = v_8194 & v_8300;
assign v_14907 = v_8029 & v_14906;
assign v_14908 = v_8044 & v_8144;
assign v_14910 = v_7885 & v_14909;
assign v_14911 = v_7909 & ~v_8012;
assign v_14913 = v_7747 & v_14912;
assign v_14914 = v_7762 & ~v_7862;
assign v_14916 = v_7583 & v_14915;
assign v_14917 = v_7618 & ~v_7730;
assign v_14919 = v_7443 & v_14918;
assign v_14920 = v_7458 & ~v_7558;
assign v_14922 = v_7297 & v_14921;
assign v_14923 = v_7323 & ~v_7426;
assign v_14925 = v_7157 & v_14924;
assign v_14926 = v_7172 & v_7272;
assign v_14928 = v_7007 & v_14927;
assign v_14929 = v_7034 & ~v_7140;
assign v_14931 = v_6869 & v_14930;
assign v_14932 = v_6884 & v_6984;
assign v_14934 = v_6725 & v_14933;
assign v_14935 = v_6749 & v_6852;
assign v_14937 = v_6587 & v_14936;
assign v_14938 = v_6602 & v_6702;
assign v_14940 = v_6430 & v_14939;
assign v_14941 = v_6461 & ~v_6570;
assign v_14943 = v_6291 & v_14942;
assign v_14944 = v_6306 & ~v_6406;
assign v_14946 = v_6146 & v_14945;
assign v_14947 = v_6171 & v_6274;
assign v_14949 = v_6007 & v_14948;
assign v_14950 = v_6022 & v_6122;
assign v_14952 = v_5857 & v_14951;
assign v_14953 = v_5884 & v_5990;
assign v_14955 = v_5719 & v_14954;
assign v_14956 = v_5734 & v_5834;
assign v_14958 = v_5575 & v_14957;
assign v_14959 = v_5599 & v_5702;
assign v_14961 = v_5437 & v_14960;
assign v_14962 = v_5452 & v_5552;
assign v_14964 = v_5266 & v_14963;
assign v_14965 = v_5305 & ~v_5420;
assign v_14967 = v_5125 & v_14966;
assign v_14968 = v_5140 & ~v_5240;
assign v_14970 = v_4978 & v_14969;
assign v_14971 = v_5005 & v_5108;
assign v_14973 = v_4837 & v_14972;
assign v_14974 = v_4852 & v_4952;
assign v_14976 = v_4687 & v_14975;
assign v_14977 = v_4714 & v_4820;
assign v_14979 = v_4549 & v_14978;
assign v_14980 = v_4564 & v_4664;
assign v_14982 = v_4405 & v_14981;
assign v_14983 = v_4429 & v_4532;
assign v_14985 = v_4267 & v_14984;
assign v_14986 = v_4282 & v_4382;
assign v_14988 = v_4110 & v_14987;
assign v_14989 = v_4141 & ~v_4250;
assign v_14991 = v_3971 & v_14990;
assign v_14992 = v_3986 & ~v_4086;
assign v_14994 = v_3826 & v_14993;
assign v_14995 = v_3851 & ~v_3954;
assign v_14997 = v_3687 & v_14996;
assign v_14998 = v_3702 & ~v_3802;
assign v_15000 = v_3537 & v_14999;
assign v_15001 = v_3564 & ~v_3670;
assign v_15003 = v_3399 & v_15002;
assign v_15004 = v_3414 & v_3514;
assign v_15006 = v_3255 & v_15005;
assign v_15007 = v_3279 & ~v_3382;
assign v_15009 = v_3117 & v_15008;
assign v_15010 = v_3132 & v_3232;
assign v_15012 = v_2953 & v_15011;
assign v_15013 = v_2988 & ~v_3100;
assign v_15015 = v_2813 & v_15014;
assign v_15016 = v_2828 & ~v_2928;
assign v_15018 = v_2667 & v_15017;
assign v_15019 = v_2693 & ~v_2796;
assign v_15021 = v_2527 & v_15020;
assign v_15022 = v_2542 & ~v_2642;
assign v_15024 = v_2377 & v_15023;
assign v_15025 = v_2404 & ~v_2510;
assign v_15027 = v_2239 & v_15026;
assign v_15028 = v_2254 & v_2354;
assign v_15030 = v_2095 & v_15029;
assign v_15031 = v_2119 & v_2222;
assign v_15033 = v_1957 & v_15032;
assign v_15034 = v_1972 & v_2072;
assign v_15036 = v_1800 & v_15035;
assign v_15037 = v_1831 & ~v_1940;
assign v_15039 = v_1661 & v_15038;
assign v_15040 = v_1676 & ~v_1776;
assign v_15042 = v_1516 & v_15041;
assign v_15043 = v_1541 & ~v_1644;
assign v_15045 = v_1377 & v_15044;
assign v_15046 = v_1392 & ~v_1492;
assign v_15048 = v_1227 & v_15047;
assign v_15049 = v_1254 & ~v_1360;
assign v_15051 = v_1089 & v_15050;
assign v_15052 = v_1104 & ~v_1204;
assign v_15054 = v_945 & v_15053;
assign v_15055 = v_969 & ~v_1072;
assign v_15057 = v_810 & v_15056;
assign v_15058 = v_826 & ~v_922;
assign v_15060 = v_223 & v_15059;
assign v_15061 = v_626 & ~v_793;
assign v_15064 = v_9611 & v_9784;
assign v_15065 = v_9639 & v_9652;
assign v_15067 = v_9468 & v_15066;
assign v_15068 = v_9483 & v_9494;
assign v_15070 = v_9320 & v_15069;
assign v_15071 = v_9347 & v_9362;
assign v_15073 = v_9180 & v_15072;
assign v_15074 = v_9195 & v_9206;
assign v_15076 = v_9037 & v_15075;
assign v_15077 = v_9061 & v_9074;
assign v_15079 = v_8898 & v_15078;
assign v_15080 = v_8913 & v_8924;
assign v_15082 = v_8744 & v_15081;
assign v_15083 = v_8775 & v_8792;
assign v_15085 = v_8602 & v_15084;
assign v_15086 = v_8617 & v_8628;
assign v_15088 = v_8458 & v_15087;
assign v_15089 = v_8483 & v_8496;
assign v_15091 = v_8318 & v_15090;
assign v_15092 = v_8333 & v_8344;
assign v_15094 = v_8170 & v_15093;
assign v_15095 = v_8197 & v_8212;
assign v_15097 = v_8030 & v_15096;
assign v_15098 = v_8045 & v_8056;
assign v_15100 = v_7887 & v_15099;
assign v_15101 = v_7911 & v_7924;
assign v_15103 = v_7748 & v_15102;
assign v_15104 = v_7763 & v_7774;
assign v_15106 = v_7588 & v_15105;
assign v_15107 = v_7623 & v_7642;
assign v_15109 = v_7444 & v_15108;
assign v_15110 = v_7459 & v_7470;
assign v_15112 = v_7299 & v_15111;
assign v_15113 = v_7325 & v_7338;
assign v_15115 = v_7158 & v_15114;
assign v_15116 = v_7173 & v_7184;
assign v_15118 = v_7010 & v_15117;
assign v_15119 = v_7037 & v_7052;
assign v_15121 = v_6870 & v_15120;
assign v_15122 = v_6885 & v_6896;
assign v_15124 = v_6727 & v_15123;
assign v_15125 = v_6751 & v_6764;
assign v_15127 = v_6588 & v_15126;
assign v_15128 = v_6603 & v_6614;
assign v_15130 = v_6434 & v_15129;
assign v_15131 = v_6465 & v_6482;
assign v_15133 = v_6292 & v_15132;
assign v_15134 = v_6307 & v_6318;
assign v_15136 = v_6148 & v_15135;
assign v_15137 = v_6173 & v_6186;
assign v_15139 = v_6008 & v_15138;
assign v_15140 = v_6023 & v_6034;
assign v_15142 = v_5860 & v_15141;
assign v_15143 = v_5887 & v_5902;
assign v_15145 = v_5720 & v_15144;
assign v_15146 = v_5735 & v_5746;
assign v_15148 = v_5577 & v_15147;
assign v_15149 = v_5601 & v_5614;
assign v_15151 = v_5438 & v_15150;
assign v_15152 = v_5453 & v_5464;
assign v_15154 = v_5272 & v_15153;
assign v_15155 = v_5311 & v_5332;
assign v_15157 = v_5126 & v_15156;
assign v_15158 = v_5141 & v_5152;
assign v_15160 = v_4980 & v_15159;
assign v_15161 = v_5007 & v_5020;
assign v_15163 = v_4838 & v_15162;
assign v_15164 = v_4853 & v_4864;
assign v_15166 = v_4690 & v_15165;
assign v_15167 = v_4717 & v_4732;
assign v_15169 = v_4550 & v_15168;
assign v_15170 = v_4565 & v_4576;
assign v_15172 = v_4407 & v_15171;
assign v_15173 = v_4431 & v_4444;
assign v_15175 = v_4268 & v_15174;
assign v_15176 = v_4283 & v_4294;
assign v_15178 = v_4114 & v_15177;
assign v_15179 = v_4145 & v_4162;
assign v_15181 = v_3972 & v_15180;
assign v_15182 = v_3987 & v_3998;
assign v_15184 = v_3828 & v_15183;
assign v_15185 = v_3853 & v_3866;
assign v_15187 = v_3688 & v_15186;
assign v_15188 = v_3703 & v_3714;
assign v_15190 = v_3540 & v_15189;
assign v_15191 = v_3567 & v_3582;
assign v_15193 = v_3400 & v_15192;
assign v_15194 = v_3415 & v_3426;
assign v_15196 = v_3257 & v_15195;
assign v_15197 = v_3281 & v_3294;
assign v_15199 = v_3118 & v_15198;
assign v_15200 = v_3133 & v_3144;
assign v_15202 = v_2958 & v_15201;
assign v_15203 = v_2993 & v_3012;
assign v_15205 = v_2814 & v_15204;
assign v_15206 = v_2829 & v_2840;
assign v_15208 = v_2669 & v_15207;
assign v_15209 = v_2695 & v_2708;
assign v_15211 = v_2528 & v_15210;
assign v_15212 = v_2543 & v_2554;
assign v_15214 = v_2380 & v_15213;
assign v_15215 = v_2407 & v_2422;
assign v_15217 = v_2240 & v_15216;
assign v_15218 = v_2255 & v_2266;
assign v_15220 = v_2097 & v_15219;
assign v_15221 = v_2121 & v_2134;
assign v_15223 = v_1958 & v_15222;
assign v_15224 = v_1973 & v_1984;
assign v_15226 = v_1804 & v_15225;
assign v_15227 = v_1835 & v_1852;
assign v_15229 = v_1662 & v_15228;
assign v_15230 = v_1677 & v_1688;
assign v_15232 = v_1518 & v_15231;
assign v_15233 = v_1543 & v_1556;
assign v_15235 = v_1378 & v_15234;
assign v_15236 = v_1393 & v_1404;
assign v_15238 = v_1230 & v_15237;
assign v_15239 = v_1257 & v_1272;
assign v_15241 = v_1090 & v_15240;
assign v_15242 = v_1105 & v_1116;
assign v_15244 = v_947 & v_15243;
assign v_15245 = v_971 & v_984;
assign v_15247 = v_811 & v_15246;
assign v_15248 = v_827 & v_838;
assign v_15250 = v_359 & v_15249;
assign v_15251 = v_658 & v_721;
assign v_15253 = v_9611 & v_9753;
assign v_15254 = v_9604 & v_9639;
assign v_15256 = v_9468 & v_15255;
assign v_15257 = v_9463 & v_9483;
assign v_15259 = v_9320 & v_15258;
assign v_15260 = v_9311 & v_9347;
assign v_15262 = v_9180 & v_15261;
assign v_15263 = v_9175 & v_9195;
assign v_15265 = v_9037 & v_15264;
assign v_15266 = v_9030 & v_9061;
assign v_15268 = v_8898 & v_15267;
assign v_15269 = v_8893 & v_8913;
assign v_15271 = v_8744 & v_15270;
assign v_15272 = v_8733 & v_8775;
assign v_15274 = v_8602 & v_15273;
assign v_15275 = v_8597 & v_8617;
assign v_15277 = v_8458 & v_15276;
assign v_15278 = v_8451 & v_8483;
assign v_15280 = v_8318 & v_15279;
assign v_15281 = v_8313 & v_8333;
assign v_15283 = v_8170 & v_15282;
assign v_15284 = v_8161 & v_8197;
assign v_15286 = v_8030 & v_15285;
assign v_15287 = v_8025 & v_8045;
assign v_15289 = v_7887 & v_15288;
assign v_15290 = v_7880 & v_7911;
assign v_15292 = v_7748 & v_15291;
assign v_15293 = v_7743 & v_7763;
assign v_15295 = v_7588 & v_15294;
assign v_15296 = v_7575 & v_7623;
assign v_15298 = v_7444 & v_15297;
assign v_15299 = v_7439 & v_7459;
assign v_15301 = v_7299 & v_15300;
assign v_15302 = v_7292 & v_7325;
assign v_15304 = v_7158 & v_15303;
assign v_15305 = v_7153 & v_7173;
assign v_15307 = v_7010 & v_15306;
assign v_15308 = v_7001 & v_7037;
assign v_15310 = v_6870 & v_15309;
assign v_15311 = v_6865 & v_6885;
assign v_15313 = v_6727 & v_15312;
assign v_15314 = v_6720 & v_6751;
assign v_15316 = v_6588 & v_15315;
assign v_15317 = v_6583 & v_6603;
assign v_15319 = v_6434 & v_15318;
assign v_15320 = v_6423 & v_6465;
assign v_15322 = v_6292 & v_15321;
assign v_15323 = v_6287 & v_6307;
assign v_15325 = v_6148 & v_15324;
assign v_15326 = v_6141 & v_6173;
assign v_15328 = v_6008 & v_15327;
assign v_15329 = v_6003 & v_6023;
assign v_15331 = v_5860 & v_15330;
assign v_15332 = v_5851 & v_5887;
assign v_15334 = v_5720 & v_15333;
assign v_15335 = v_5715 & v_5735;
assign v_15337 = v_5577 & v_15336;
assign v_15338 = v_5570 & v_5601;
assign v_15340 = v_5438 & v_15339;
assign v_15341 = v_5433 & v_5453;
assign v_15343 = v_5272 & v_15342;
assign v_15344 = v_5257 & v_5311;
assign v_15346 = v_5126 & v_15345;
assign v_15347 = v_5121 & v_5141;
assign v_15349 = v_4980 & v_15348;
assign v_15350 = v_4973 & v_5007;
assign v_15352 = v_4838 & v_15351;
assign v_15353 = v_4833 & v_4853;
assign v_15355 = v_4690 & v_15354;
assign v_15356 = v_4681 & v_4717;
assign v_15358 = v_4550 & v_15357;
assign v_15359 = v_4545 & v_4565;
assign v_15361 = v_4407 & v_15360;
assign v_15362 = v_4400 & v_4431;
assign v_15364 = v_4268 & v_15363;
assign v_15365 = v_4263 & v_4283;
assign v_15367 = v_4114 & v_15366;
assign v_15368 = v_4103 & v_4145;
assign v_15370 = v_3972 & v_15369;
assign v_15371 = v_3967 & v_3987;
assign v_15373 = v_3828 & v_15372;
assign v_15374 = v_3821 & v_3853;
assign v_15376 = v_3688 & v_15375;
assign v_15377 = v_3683 & v_3703;
assign v_15379 = v_3540 & v_15378;
assign v_15380 = v_3531 & v_3567;
assign v_15382 = v_3400 & v_15381;
assign v_15383 = v_3395 & v_3415;
assign v_15385 = v_3257 & v_15384;
assign v_15386 = v_3250 & v_3281;
assign v_15388 = v_3118 & v_15387;
assign v_15389 = v_3113 & v_3133;
assign v_15391 = v_2958 & v_15390;
assign v_15392 = v_2945 & v_2993;
assign v_15394 = v_2814 & v_15393;
assign v_15395 = v_2809 & v_2829;
assign v_15397 = v_2669 & v_15396;
assign v_15398 = v_2662 & v_2695;
assign v_15400 = v_2528 & v_15399;
assign v_15401 = v_2523 & v_2543;
assign v_15403 = v_2380 & v_15402;
assign v_15404 = v_2371 & v_2407;
assign v_15406 = v_2240 & v_15405;
assign v_15407 = v_2235 & v_2255;
assign v_15409 = v_2097 & v_15408;
assign v_15410 = v_2090 & v_2121;
assign v_15412 = v_1958 & v_15411;
assign v_15413 = v_1953 & v_1973;
assign v_15415 = v_1804 & v_15414;
assign v_15416 = v_1793 & v_1835;
assign v_15418 = v_1662 & v_15417;
assign v_15419 = v_1657 & v_1677;
assign v_15421 = v_1518 & v_15420;
assign v_15422 = v_1511 & v_1543;
assign v_15424 = v_1378 & v_15423;
assign v_15425 = v_1373 & v_1393;
assign v_15427 = v_1230 & v_15426;
assign v_15428 = v_1221 & v_1257;
assign v_15430 = v_1090 & v_15429;
assign v_15431 = v_1085 & v_1105;
assign v_15433 = v_947 & v_15432;
assign v_15434 = v_940 & v_971;
assign v_15436 = v_811 & v_15435;
assign v_15437 = v_804 & v_827;
assign v_15439 = v_359 & v_15438;
assign v_15440 = v_98 & v_658;
assign v_15443 = v_9611 & v_9796;
assign v_15444 = v_9639 & v_9664;
assign v_15446 = v_9468 & v_15445;
assign v_15447 = v_9483 & v_9506;
assign v_15449 = v_9320 & v_15448;
assign v_15450 = v_9347 & v_9374;
assign v_15452 = v_9180 & v_15451;
assign v_15453 = v_9195 & v_9218;
assign v_15455 = v_9037 & v_15454;
assign v_15456 = v_9061 & v_9086;
assign v_15458 = v_8898 & v_15457;
assign v_15459 = v_8913 & v_8936;
assign v_15461 = v_8744 & v_15460;
assign v_15462 = v_8775 & v_8804;
assign v_15464 = v_8602 & v_15463;
assign v_15465 = v_8617 & v_8640;
assign v_15467 = v_8458 & v_15466;
assign v_15468 = v_8483 & v_8508;
assign v_15470 = v_8318 & v_15469;
assign v_15471 = v_8333 & v_8356;
assign v_15473 = v_8170 & v_15472;
assign v_15474 = v_8197 & v_8224;
assign v_15476 = v_8030 & v_15475;
assign v_15477 = v_8045 & v_8068;
assign v_15479 = v_7887 & v_15478;
assign v_15480 = v_7911 & v_7936;
assign v_15482 = v_7748 & v_15481;
assign v_15483 = v_7763 & v_7786;
assign v_15485 = v_7588 & v_15484;
assign v_15486 = v_7623 & v_7654;
assign v_15488 = v_7444 & v_15487;
assign v_15489 = v_7459 & v_7482;
assign v_15491 = v_7299 & v_15490;
assign v_15492 = v_7325 & v_7350;
assign v_15494 = v_7158 & v_15493;
assign v_15495 = v_7173 & v_7196;
assign v_15497 = v_7010 & v_15496;
assign v_15498 = v_7037 & v_7064;
assign v_15500 = v_6870 & v_15499;
assign v_15501 = v_6885 & v_6908;
assign v_15503 = v_6727 & v_15502;
assign v_15504 = v_6751 & v_6776;
assign v_15506 = v_6588 & v_15505;
assign v_15507 = v_6603 & v_6626;
assign v_15509 = v_6434 & v_15508;
assign v_15510 = v_6465 & v_6494;
assign v_15512 = v_6292 & v_15511;
assign v_15513 = v_6307 & v_6330;
assign v_15515 = v_6148 & v_15514;
assign v_15516 = v_6173 & v_6198;
assign v_15518 = v_6008 & v_15517;
assign v_15519 = v_6023 & v_6046;
assign v_15521 = v_5860 & v_15520;
assign v_15522 = v_5887 & v_5914;
assign v_15524 = v_5720 & v_15523;
assign v_15525 = v_5735 & v_5758;
assign v_15527 = v_5577 & v_15526;
assign v_15528 = v_5601 & v_5626;
assign v_15530 = v_5438 & v_15529;
assign v_15531 = v_5453 & v_5476;
assign v_15533 = v_5272 & v_15532;
assign v_15534 = v_5311 & v_5344;
assign v_15536 = v_5126 & v_15535;
assign v_15537 = v_5141 & v_5164;
assign v_15539 = v_4980 & v_15538;
assign v_15540 = v_5007 & v_5032;
assign v_15542 = v_4838 & v_15541;
assign v_15543 = v_4853 & v_4876;
assign v_15545 = v_4690 & v_15544;
assign v_15546 = v_4717 & v_4744;
assign v_15548 = v_4550 & v_15547;
assign v_15549 = v_4565 & v_4588;
assign v_15551 = v_4407 & v_15550;
assign v_15552 = v_4431 & v_4456;
assign v_15554 = v_4268 & v_15553;
assign v_15555 = v_4283 & v_4306;
assign v_15557 = v_4114 & v_15556;
assign v_15558 = v_4145 & v_4174;
assign v_15560 = v_3972 & v_15559;
assign v_15561 = v_3987 & v_4010;
assign v_15563 = v_3828 & v_15562;
assign v_15564 = v_3853 & v_3878;
assign v_15566 = v_3688 & v_15565;
assign v_15567 = v_3703 & v_3726;
assign v_15569 = v_3540 & v_15568;
assign v_15570 = v_3567 & v_3594;
assign v_15572 = v_3400 & v_15571;
assign v_15573 = v_3415 & v_3438;
assign v_15575 = v_3257 & v_15574;
assign v_15576 = v_3281 & v_3306;
assign v_15578 = v_3118 & v_15577;
assign v_15579 = v_3133 & v_3156;
assign v_15581 = v_2958 & v_15580;
assign v_15582 = v_2993 & v_3024;
assign v_15584 = v_2814 & v_15583;
assign v_15585 = v_2829 & v_2852;
assign v_15587 = v_2669 & v_15586;
assign v_15588 = v_2695 & v_2720;
assign v_15590 = v_2528 & v_15589;
assign v_15591 = v_2543 & v_2566;
assign v_15593 = v_2380 & v_15592;
assign v_15594 = v_2407 & v_2434;
assign v_15596 = v_2240 & v_15595;
assign v_15597 = v_2255 & v_2278;
assign v_15599 = v_2097 & v_15598;
assign v_15600 = v_2121 & v_2146;
assign v_15602 = v_1958 & v_15601;
assign v_15603 = v_1973 & v_1996;
assign v_15605 = v_1804 & v_15604;
assign v_15606 = v_1835 & v_1864;
assign v_15608 = v_1662 & v_15607;
assign v_15609 = v_1677 & v_1700;
assign v_15611 = v_1518 & v_15610;
assign v_15612 = v_1543 & v_1568;
assign v_15614 = v_1378 & v_15613;
assign v_15615 = v_1393 & v_1416;
assign v_15617 = v_1230 & v_15616;
assign v_15618 = v_1257 & v_1284;
assign v_15620 = v_1090 & v_15619;
assign v_15621 = v_1105 & v_1128;
assign v_15623 = v_947 & v_15622;
assign v_15624 = v_971 & v_996;
assign v_15626 = v_811 & v_15625;
assign v_15627 = v_827 & v_850;
assign v_15629 = v_359 & v_15628;
assign v_15630 = v_658 & v_731;
assign v_15633 = v_9611 & v_9808;
assign v_15634 = v_9639 & v_9676;
assign v_15636 = v_9468 & v_15635;
assign v_15637 = v_9483 & v_9518;
assign v_15639 = v_9320 & v_15638;
assign v_15640 = v_9347 & v_9386;
assign v_15642 = v_9180 & v_15641;
assign v_15643 = v_9195 & v_9230;
assign v_15645 = v_9037 & v_15644;
assign v_15646 = v_9061 & v_9098;
assign v_15648 = v_8898 & v_15647;
assign v_15649 = v_8913 & v_8948;
assign v_15651 = v_8744 & v_15650;
assign v_15652 = v_8775 & v_8816;
assign v_15654 = v_8602 & v_15653;
assign v_15655 = v_8617 & v_8652;
assign v_15657 = v_8458 & v_15656;
assign v_15658 = v_8483 & v_8520;
assign v_15660 = v_8318 & v_15659;
assign v_15661 = v_8333 & v_8368;
assign v_15663 = v_8170 & v_15662;
assign v_15664 = v_8197 & v_8236;
assign v_15666 = v_8030 & v_15665;
assign v_15667 = v_8045 & v_8080;
assign v_15669 = v_7887 & v_15668;
assign v_15670 = v_7911 & v_7948;
assign v_15672 = v_7748 & v_15671;
assign v_15673 = v_7763 & v_7798;
assign v_15675 = v_7588 & v_15674;
assign v_15676 = v_7623 & v_7666;
assign v_15678 = v_7444 & v_15677;
assign v_15679 = v_7459 & v_7494;
assign v_15681 = v_7299 & v_15680;
assign v_15682 = v_7325 & v_7362;
assign v_15684 = v_7158 & v_15683;
assign v_15685 = v_7173 & v_7208;
assign v_15687 = v_7010 & v_15686;
assign v_15688 = v_7037 & v_7076;
assign v_15690 = v_6870 & v_15689;
assign v_15691 = v_6885 & v_6920;
assign v_15693 = v_6727 & v_15692;
assign v_15694 = v_6751 & v_6788;
assign v_15696 = v_6588 & v_15695;
assign v_15697 = v_6603 & v_6638;
assign v_15699 = v_6434 & v_15698;
assign v_15700 = v_6465 & v_6506;
assign v_15702 = v_6292 & v_15701;
assign v_15703 = v_6307 & v_6342;
assign v_15705 = v_6148 & v_15704;
assign v_15706 = v_6173 & v_6210;
assign v_15708 = v_6008 & v_15707;
assign v_15709 = v_6023 & v_6058;
assign v_15711 = v_5860 & v_15710;
assign v_15712 = v_5887 & v_5926;
assign v_15714 = v_5720 & v_15713;
assign v_15715 = v_5735 & v_5770;
assign v_15717 = v_5577 & v_15716;
assign v_15718 = v_5601 & v_5638;
assign v_15720 = v_5438 & v_15719;
assign v_15721 = v_5453 & v_5488;
assign v_15723 = v_5272 & v_15722;
assign v_15724 = v_5311 & v_5356;
assign v_15726 = v_5126 & v_15725;
assign v_15727 = v_5141 & v_5176;
assign v_15729 = v_4980 & v_15728;
assign v_15730 = v_5007 & v_5044;
assign v_15732 = v_4838 & v_15731;
assign v_15733 = v_4853 & v_4888;
assign v_15735 = v_4690 & v_15734;
assign v_15736 = v_4717 & v_4756;
assign v_15738 = v_4550 & v_15737;
assign v_15739 = v_4565 & v_4600;
assign v_15741 = v_4407 & v_15740;
assign v_15742 = v_4431 & v_4468;
assign v_15744 = v_4268 & v_15743;
assign v_15745 = v_4283 & v_4318;
assign v_15747 = v_4114 & v_15746;
assign v_15748 = v_4145 & v_4186;
assign v_15750 = v_3972 & v_15749;
assign v_15751 = v_3987 & v_4022;
assign v_15753 = v_3828 & v_15752;
assign v_15754 = v_3853 & v_3890;
assign v_15756 = v_3688 & v_15755;
assign v_15757 = v_3703 & v_3738;
assign v_15759 = v_3540 & v_15758;
assign v_15760 = v_3567 & v_3606;
assign v_15762 = v_3400 & v_15761;
assign v_15763 = v_3415 & v_3450;
assign v_15765 = v_3257 & v_15764;
assign v_15766 = v_3281 & v_3318;
assign v_15768 = v_3118 & v_15767;
assign v_15769 = v_3133 & v_3168;
assign v_15771 = v_2958 & v_15770;
assign v_15772 = v_2993 & v_3036;
assign v_15774 = v_2814 & v_15773;
assign v_15775 = v_2829 & v_2864;
assign v_15777 = v_2669 & v_15776;
assign v_15778 = v_2695 & v_2732;
assign v_15780 = v_2528 & v_15779;
assign v_15781 = v_2543 & v_2578;
assign v_15783 = v_2380 & v_15782;
assign v_15784 = v_2407 & v_2446;
assign v_15786 = v_2240 & v_15785;
assign v_15787 = v_2255 & v_2290;
assign v_15789 = v_2097 & v_15788;
assign v_15790 = v_2121 & v_2158;
assign v_15792 = v_1958 & v_15791;
assign v_15793 = v_1973 & v_2008;
assign v_15795 = v_1804 & v_15794;
assign v_15796 = v_1835 & v_1876;
assign v_15798 = v_1662 & v_15797;
assign v_15799 = v_1677 & v_1712;
assign v_15801 = v_1518 & v_15800;
assign v_15802 = v_1543 & v_1580;
assign v_15804 = v_1378 & v_15803;
assign v_15805 = v_1393 & v_1428;
assign v_15807 = v_1230 & v_15806;
assign v_15808 = v_1257 & v_1296;
assign v_15810 = v_1090 & v_15809;
assign v_15811 = v_1105 & v_1140;
assign v_15813 = v_947 & v_15812;
assign v_15814 = v_971 & v_1008;
assign v_15816 = v_811 & v_15815;
assign v_15817 = v_827 & v_862;
assign v_15819 = v_359 & v_15818;
assign v_15820 = v_658 & v_741;
assign v_15823 = v_9611 & v_9820;
assign v_15824 = v_9639 & v_9688;
assign v_15826 = v_9468 & v_15825;
assign v_15827 = v_9483 & v_9530;
assign v_15829 = v_9320 & v_15828;
assign v_15830 = v_9347 & v_9398;
assign v_15832 = v_9180 & v_15831;
assign v_15833 = v_9195 & v_9242;
assign v_15835 = v_9037 & v_15834;
assign v_15836 = v_9061 & v_9110;
assign v_15838 = v_8898 & v_15837;
assign v_15839 = v_8913 & v_8960;
assign v_15841 = v_8744 & v_15840;
assign v_15842 = v_8775 & v_8828;
assign v_15844 = v_8602 & v_15843;
assign v_15845 = v_8617 & v_8664;
assign v_15847 = v_8458 & v_15846;
assign v_15848 = v_8483 & v_8532;
assign v_15850 = v_8318 & v_15849;
assign v_15851 = v_8333 & v_8380;
assign v_15853 = v_8170 & v_15852;
assign v_15854 = v_8197 & v_8248;
assign v_15856 = v_8030 & v_15855;
assign v_15857 = v_8045 & v_8092;
assign v_15859 = v_7887 & v_15858;
assign v_15860 = v_7911 & v_7960;
assign v_15862 = v_7748 & v_15861;
assign v_15863 = v_7763 & v_7810;
assign v_15865 = v_7588 & v_15864;
assign v_15866 = v_7623 & v_7678;
assign v_15868 = v_7444 & v_15867;
assign v_15869 = v_7459 & v_7506;
assign v_15871 = v_7299 & v_15870;
assign v_15872 = v_7325 & v_7374;
assign v_15874 = v_7158 & v_15873;
assign v_15875 = v_7173 & v_7220;
assign v_15877 = v_7010 & v_15876;
assign v_15878 = v_7037 & v_7088;
assign v_15880 = v_6870 & v_15879;
assign v_15881 = v_6885 & v_6932;
assign v_15883 = v_6727 & v_15882;
assign v_15884 = v_6751 & v_6800;
assign v_15886 = v_6588 & v_15885;
assign v_15887 = v_6603 & v_6650;
assign v_15889 = v_6434 & v_15888;
assign v_15890 = v_6465 & v_6518;
assign v_15892 = v_6292 & v_15891;
assign v_15893 = v_6307 & v_6354;
assign v_15895 = v_6148 & v_15894;
assign v_15896 = v_6173 & v_6222;
assign v_15898 = v_6008 & v_15897;
assign v_15899 = v_6023 & v_6070;
assign v_15901 = v_5860 & v_15900;
assign v_15902 = v_5887 & v_5938;
assign v_15904 = v_5720 & v_15903;
assign v_15905 = v_5735 & v_5782;
assign v_15907 = v_5577 & v_15906;
assign v_15908 = v_5601 & v_5650;
assign v_15910 = v_5438 & v_15909;
assign v_15911 = v_5453 & v_5500;
assign v_15913 = v_5272 & v_15912;
assign v_15914 = v_5311 & v_5368;
assign v_15916 = v_5126 & v_15915;
assign v_15917 = v_5141 & v_5188;
assign v_15919 = v_4980 & v_15918;
assign v_15920 = v_5007 & v_5056;
assign v_15922 = v_4838 & v_15921;
assign v_15923 = v_4853 & v_4900;
assign v_15925 = v_4690 & v_15924;
assign v_15926 = v_4717 & v_4768;
assign v_15928 = v_4550 & v_15927;
assign v_15929 = v_4565 & v_4612;
assign v_15931 = v_4407 & v_15930;
assign v_15932 = v_4431 & v_4480;
assign v_15934 = v_4268 & v_15933;
assign v_15935 = v_4283 & v_4330;
assign v_15937 = v_4114 & v_15936;
assign v_15938 = v_4145 & v_4198;
assign v_15940 = v_3972 & v_15939;
assign v_15941 = v_3987 & v_4034;
assign v_15943 = v_3828 & v_15942;
assign v_15944 = v_3853 & v_3902;
assign v_15946 = v_3688 & v_15945;
assign v_15947 = v_3703 & v_3750;
assign v_15949 = v_3540 & v_15948;
assign v_15950 = v_3567 & v_3618;
assign v_15952 = v_3400 & v_15951;
assign v_15953 = v_3415 & v_3462;
assign v_15955 = v_3257 & v_15954;
assign v_15956 = v_3281 & v_3330;
assign v_15958 = v_3118 & v_15957;
assign v_15959 = v_3133 & v_3180;
assign v_15961 = v_2958 & v_15960;
assign v_15962 = v_2993 & v_3048;
assign v_15964 = v_2814 & v_15963;
assign v_15965 = v_2829 & v_2876;
assign v_15967 = v_2669 & v_15966;
assign v_15968 = v_2695 & v_2744;
assign v_15970 = v_2528 & v_15969;
assign v_15971 = v_2543 & v_2590;
assign v_15973 = v_2380 & v_15972;
assign v_15974 = v_2407 & v_2458;
assign v_15976 = v_2240 & v_15975;
assign v_15977 = v_2255 & v_2302;
assign v_15979 = v_2097 & v_15978;
assign v_15980 = v_2121 & v_2170;
assign v_15982 = v_1958 & v_15981;
assign v_15983 = v_1973 & v_2020;
assign v_15985 = v_1804 & v_15984;
assign v_15986 = v_1835 & v_1888;
assign v_15988 = v_1662 & v_15987;
assign v_15989 = v_1677 & v_1724;
assign v_15991 = v_1518 & v_15990;
assign v_15992 = v_1543 & v_1592;
assign v_15994 = v_1378 & v_15993;
assign v_15995 = v_1393 & v_1440;
assign v_15997 = v_1230 & v_15996;
assign v_15998 = v_1257 & v_1308;
assign v_16000 = v_1090 & v_15999;
assign v_16001 = v_1105 & v_1152;
assign v_16003 = v_947 & v_16002;
assign v_16004 = v_971 & v_1020;
assign v_16006 = v_811 & v_16005;
assign v_16007 = v_827 & v_874;
assign v_16009 = v_359 & v_16008;
assign v_16010 = v_658 & v_751;
assign v_16013 = v_9611 & v_9832;
assign v_16014 = v_9639 & v_9700;
assign v_16016 = v_9468 & v_16015;
assign v_16017 = v_9483 & v_9542;
assign v_16019 = v_9320 & v_16018;
assign v_16020 = v_9347 & v_9410;
assign v_16022 = v_9180 & v_16021;
assign v_16023 = v_9195 & v_9254;
assign v_16025 = v_9037 & v_16024;
assign v_16026 = v_9061 & v_9122;
assign v_16028 = v_8898 & v_16027;
assign v_16029 = v_8913 & v_8972;
assign v_16031 = v_8744 & v_16030;
assign v_16032 = v_8775 & v_8840;
assign v_16034 = v_8602 & v_16033;
assign v_16035 = v_8617 & v_8676;
assign v_16037 = v_8458 & v_16036;
assign v_16038 = v_8483 & v_8544;
assign v_16040 = v_8318 & v_16039;
assign v_16041 = v_8333 & v_8392;
assign v_16043 = v_8170 & v_16042;
assign v_16044 = v_8197 & v_8260;
assign v_16046 = v_8030 & v_16045;
assign v_16047 = v_8045 & v_8104;
assign v_16049 = v_7887 & v_16048;
assign v_16050 = v_7911 & v_7972;
assign v_16052 = v_7748 & v_16051;
assign v_16053 = v_7763 & v_7822;
assign v_16055 = v_7588 & v_16054;
assign v_16056 = v_7623 & v_7690;
assign v_16058 = v_7444 & v_16057;
assign v_16059 = v_7459 & v_7518;
assign v_16061 = v_7299 & v_16060;
assign v_16062 = v_7325 & v_7386;
assign v_16064 = v_7158 & v_16063;
assign v_16065 = v_7173 & v_7232;
assign v_16067 = v_7010 & v_16066;
assign v_16068 = v_7037 & v_7100;
assign v_16070 = v_6870 & v_16069;
assign v_16071 = v_6885 & v_6944;
assign v_16073 = v_6727 & v_16072;
assign v_16074 = v_6751 & v_6812;
assign v_16076 = v_6588 & v_16075;
assign v_16077 = v_6603 & v_6662;
assign v_16079 = v_6434 & v_16078;
assign v_16080 = v_6465 & v_6530;
assign v_16082 = v_6292 & v_16081;
assign v_16083 = v_6307 & v_6366;
assign v_16085 = v_6148 & v_16084;
assign v_16086 = v_6173 & v_6234;
assign v_16088 = v_6008 & v_16087;
assign v_16089 = v_6023 & v_6082;
assign v_16091 = v_5860 & v_16090;
assign v_16092 = v_5887 & v_5950;
assign v_16094 = v_5720 & v_16093;
assign v_16095 = v_5735 & v_5794;
assign v_16097 = v_5577 & v_16096;
assign v_16098 = v_5601 & v_5662;
assign v_16100 = v_5438 & v_16099;
assign v_16101 = v_5453 & v_5512;
assign v_16103 = v_5272 & v_16102;
assign v_16104 = v_5311 & v_5380;
assign v_16106 = v_5126 & v_16105;
assign v_16107 = v_5141 & v_5200;
assign v_16109 = v_4980 & v_16108;
assign v_16110 = v_5007 & v_5068;
assign v_16112 = v_4838 & v_16111;
assign v_16113 = v_4853 & v_4912;
assign v_16115 = v_4690 & v_16114;
assign v_16116 = v_4717 & v_4780;
assign v_16118 = v_4550 & v_16117;
assign v_16119 = v_4565 & v_4624;
assign v_16121 = v_4407 & v_16120;
assign v_16122 = v_4431 & v_4492;
assign v_16124 = v_4268 & v_16123;
assign v_16125 = v_4283 & v_4342;
assign v_16127 = v_4114 & v_16126;
assign v_16128 = v_4145 & v_4210;
assign v_16130 = v_3972 & v_16129;
assign v_16131 = v_3987 & v_4046;
assign v_16133 = v_3828 & v_16132;
assign v_16134 = v_3853 & v_3914;
assign v_16136 = v_3688 & v_16135;
assign v_16137 = v_3703 & v_3762;
assign v_16139 = v_3540 & v_16138;
assign v_16140 = v_3567 & v_3630;
assign v_16142 = v_3400 & v_16141;
assign v_16143 = v_3415 & v_3474;
assign v_16145 = v_3257 & v_16144;
assign v_16146 = v_3281 & v_3342;
assign v_16148 = v_3118 & v_16147;
assign v_16149 = v_3133 & v_3192;
assign v_16151 = v_2958 & v_16150;
assign v_16152 = v_2993 & v_3060;
assign v_16154 = v_2814 & v_16153;
assign v_16155 = v_2829 & v_2888;
assign v_16157 = v_2669 & v_16156;
assign v_16158 = v_2695 & v_2756;
assign v_16160 = v_2528 & v_16159;
assign v_16161 = v_2543 & v_2602;
assign v_16163 = v_2380 & v_16162;
assign v_16164 = v_2407 & v_2470;
assign v_16166 = v_2240 & v_16165;
assign v_16167 = v_2255 & v_2314;
assign v_16169 = v_2097 & v_16168;
assign v_16170 = v_2121 & v_2182;
assign v_16172 = v_1958 & v_16171;
assign v_16173 = v_1973 & v_2032;
assign v_16175 = v_1804 & v_16174;
assign v_16176 = v_1835 & v_1900;
assign v_16178 = v_1662 & v_16177;
assign v_16179 = v_1677 & v_1736;
assign v_16181 = v_1518 & v_16180;
assign v_16182 = v_1543 & v_1604;
assign v_16184 = v_1378 & v_16183;
assign v_16185 = v_1393 & v_1452;
assign v_16187 = v_1230 & v_16186;
assign v_16188 = v_1257 & v_1320;
assign v_16190 = v_1090 & v_16189;
assign v_16191 = v_1105 & v_1164;
assign v_16193 = v_947 & v_16192;
assign v_16194 = v_971 & v_1032;
assign v_16196 = v_811 & v_16195;
assign v_16197 = v_827 & v_886;
assign v_16199 = v_359 & v_16198;
assign v_16200 = v_658 & v_761;
assign v_16205 = v_16203 & v_16204;
assign v_16208 = v_16206 & v_16207;
assign v_16211 = v_16209 & v_16210;
assign v_16214 = v_16212 & v_16213;
assign v_16217 = v_16215 & v_16216;
assign v_16220 = v_16218 & v_16219;
assign v_16223 = v_16221 & v_16222;
assign v_16226 = v_16224 & v_16225;
assign v_16229 = v_16227 & v_16228;
assign v_16232 = v_16230 & v_16231;
assign v_16235 = v_16233 & v_16234;
assign v_16238 = v_16236 & v_16237;
assign v_16241 = v_16239 & v_16240;
assign v_16244 = v_16242 & v_16243;
assign v_16247 = v_16245 & v_16246;
assign v_16250 = v_16248 & v_16249;
assign v_16253 = v_16251 & v_16252;
assign v_16256 = v_16254 & v_16255;
assign v_16259 = v_16257 & v_16258;
assign v_16262 = v_16260 & v_16261;
assign v_16265 = v_16263 & v_16264;
assign v_16268 = v_16266 & v_16267;
assign v_16271 = v_16269 & v_16270;
assign v_16274 = v_16272 & v_16273;
assign v_16277 = v_16275 & v_16276;
assign v_16280 = v_16278 & v_16279;
assign v_16283 = v_16281 & v_16282;
assign v_16286 = v_16284 & v_16285;
assign v_16289 = v_16287 & v_16288;
assign v_16292 = v_16290 & v_16291;
assign v_16295 = v_16293 & v_16294;
assign v_16298 = v_16296 & v_16297;
assign v_16301 = v_16299 & v_16300;
assign v_16304 = v_16302 & v_16303;
assign v_16307 = v_16305 & v_16306;
assign v_16310 = v_16308 & v_16309;
assign v_16313 = v_16311 & v_16312;
assign v_16316 = v_16314 & v_16315;
assign v_16319 = v_16317 & v_16318;
assign v_16322 = v_16320 & v_16321;
assign v_16325 = v_16323 & v_16324;
assign v_16328 = v_16326 & v_16327;
assign v_16331 = v_16329 & v_16330;
assign v_16334 = v_16332 & v_16333;
assign v_16337 = v_16335 & v_16336;
assign v_16340 = v_16338 & v_16339;
assign v_16343 = v_16341 & v_16342;
assign v_16346 = v_16344 & v_16345;
assign v_16349 = v_16347 & v_16348;
assign v_16352 = v_16350 & v_16351;
assign v_16355 = v_16353 & v_16354;
assign v_16358 = v_16356 & v_16357;
assign v_16361 = v_16359 & v_16360;
assign v_16364 = v_16362 & v_16363;
assign v_16367 = v_16365 & v_16366;
assign v_16370 = v_16368 & v_16369;
assign v_16373 = v_16371 & v_16372;
assign v_16376 = v_16374 & v_16375;
assign v_16379 = v_16377 & v_16378;
assign v_16382 = v_16380 & v_16381;
assign v_16385 = v_16383 & v_16384;
assign v_16388 = v_16386 & v_16387;
assign v_16391 = v_16389 & v_16390;
assign v_16393 = v_9611 & ~v_9872;
assign v_16394 = v_9639 & ~v_9740;
assign v_16396 = v_9468 & v_16395;
assign v_16397 = v_9483 & ~v_9582;
assign v_16399 = v_9320 & v_16398;
assign v_16400 = v_9347 & ~v_9450;
assign v_16402 = v_9180 & v_16401;
assign v_16403 = v_9195 & ~v_9294;
assign v_16405 = v_9037 & v_16404;
assign v_16406 = v_9061 & ~v_9162;
assign v_16408 = v_8898 & v_16407;
assign v_16409 = v_8913 & ~v_9012;
assign v_16411 = v_8744 & v_16410;
assign v_16412 = v_8775 & ~v_8880;
assign v_16414 = v_8602 & v_16413;
assign v_16415 = v_8617 & ~v_8716;
assign v_16417 = v_8458 & v_16416;
assign v_16418 = v_8483 & ~v_8584;
assign v_16420 = v_8318 & v_16419;
assign v_16421 = v_8333 & v_8432;
assign v_16423 = v_8170 & v_16422;
assign v_16424 = v_8197 & v_8300;
assign v_16426 = v_8030 & v_16425;
assign v_16427 = v_8045 & v_8144;
assign v_16429 = v_7887 & v_16428;
assign v_16430 = v_7911 & ~v_8012;
assign v_16432 = v_7748 & v_16431;
assign v_16433 = v_7763 & ~v_7862;
assign v_16435 = v_7588 & v_16434;
assign v_16436 = v_7623 & ~v_7730;
assign v_16438 = v_7444 & v_16437;
assign v_16439 = v_7459 & ~v_7558;
assign v_16441 = v_7299 & v_16440;
assign v_16442 = v_7325 & ~v_7426;
assign v_16444 = v_7158 & v_16443;
assign v_16445 = v_7173 & v_7272;
assign v_16447 = v_7010 & v_16446;
assign v_16448 = v_7037 & ~v_7140;
assign v_16450 = v_6870 & v_16449;
assign v_16451 = v_6885 & v_6984;
assign v_16453 = v_6727 & v_16452;
assign v_16454 = v_6751 & v_6852;
assign v_16456 = v_6588 & v_16455;
assign v_16457 = v_6603 & v_6702;
assign v_16459 = v_6434 & v_16458;
assign v_16460 = v_6465 & ~v_6570;
assign v_16462 = v_6292 & v_16461;
assign v_16463 = v_6307 & ~v_6406;
assign v_16465 = v_6148 & v_16464;
assign v_16466 = v_6173 & v_6274;
assign v_16468 = v_6008 & v_16467;
assign v_16469 = v_6023 & v_6122;
assign v_16471 = v_5860 & v_16470;
assign v_16472 = v_5887 & v_5990;
assign v_16474 = v_5720 & v_16473;
assign v_16475 = v_5735 & v_5834;
assign v_16477 = v_5577 & v_16476;
assign v_16478 = v_5601 & v_5702;
assign v_16480 = v_5438 & v_16479;
assign v_16481 = v_5453 & v_5552;
assign v_16483 = v_5272 & v_16482;
assign v_16484 = v_5311 & ~v_5420;
assign v_16486 = v_5126 & v_16485;
assign v_16487 = v_5141 & ~v_5240;
assign v_16489 = v_4980 & v_16488;
assign v_16490 = v_5007 & v_5108;
assign v_16492 = v_4838 & v_16491;
assign v_16493 = v_4853 & v_4952;
assign v_16495 = v_4690 & v_16494;
assign v_16496 = v_4717 & v_4820;
assign v_16498 = v_4550 & v_16497;
assign v_16499 = v_4565 & v_4664;
assign v_16501 = v_4407 & v_16500;
assign v_16502 = v_4431 & v_4532;
assign v_16504 = v_4268 & v_16503;
assign v_16505 = v_4283 & v_4382;
assign v_16507 = v_4114 & v_16506;
assign v_16508 = v_4145 & ~v_4250;
assign v_16510 = v_3972 & v_16509;
assign v_16511 = v_3987 & ~v_4086;
assign v_16513 = v_3828 & v_16512;
assign v_16514 = v_3853 & ~v_3954;
assign v_16516 = v_3688 & v_16515;
assign v_16517 = v_3703 & ~v_3802;
assign v_16519 = v_3540 & v_16518;
assign v_16520 = v_3567 & ~v_3670;
assign v_16522 = v_3400 & v_16521;
assign v_16523 = v_3415 & v_3514;
assign v_16525 = v_3257 & v_16524;
assign v_16526 = v_3281 & ~v_3382;
assign v_16528 = v_3118 & v_16527;
assign v_16529 = v_3133 & v_3232;
assign v_16531 = v_2958 & v_16530;
assign v_16532 = v_2993 & ~v_3100;
assign v_16534 = v_2814 & v_16533;
assign v_16535 = v_2829 & ~v_2928;
assign v_16537 = v_2669 & v_16536;
assign v_16538 = v_2695 & ~v_2796;
assign v_16540 = v_2528 & v_16539;
assign v_16541 = v_2543 & ~v_2642;
assign v_16543 = v_2380 & v_16542;
assign v_16544 = v_2407 & ~v_2510;
assign v_16546 = v_2240 & v_16545;
assign v_16547 = v_2255 & v_2354;
assign v_16549 = v_2097 & v_16548;
assign v_16550 = v_2121 & v_2222;
assign v_16552 = v_1958 & v_16551;
assign v_16553 = v_1973 & v_2072;
assign v_16555 = v_1804 & v_16554;
assign v_16556 = v_1835 & ~v_1940;
assign v_16558 = v_1662 & v_16557;
assign v_16559 = v_1677 & ~v_1776;
assign v_16561 = v_1518 & v_16560;
assign v_16562 = v_1543 & ~v_1644;
assign v_16564 = v_1378 & v_16563;
assign v_16565 = v_1393 & ~v_1492;
assign v_16567 = v_1230 & v_16566;
assign v_16568 = v_1257 & ~v_1360;
assign v_16570 = v_1090 & v_16569;
assign v_16571 = v_1105 & ~v_1204;
assign v_16573 = v_947 & v_16572;
assign v_16574 = v_971 & ~v_1072;
assign v_16576 = v_811 & v_16575;
assign v_16577 = v_827 & ~v_922;
assign v_16579 = v_359 & v_16578;
assign v_16580 = v_658 & ~v_793;
assign v_16586 = v_361 & v_16585;
assign v_16587 = v_9026 & v_9784;
assign v_16588 = v_9051 & v_9652;
assign v_16590 = v_9027 & v_16589;
assign v_16591 = v_9052 & v_9494;
assign v_16593 = v_8729 & v_16592;
assign v_16594 = v_8761 & v_9362;
assign v_16596 = v_8730 & v_16595;
assign v_16597 = v_8762 & v_9206;
assign v_16599 = v_8447 & v_16598;
assign v_16600 = v_8473 & v_9074;
assign v_16602 = v_8448 & v_16601;
assign v_16603 = v_8474 & v_8924;
assign v_16605 = v_8157 & v_16604;
assign v_16606 = v_8185 & v_8792;
assign v_16608 = v_8158 & v_16607;
assign v_16609 = v_8186 & v_8628;
assign v_16611 = v_7876 & v_16610;
assign v_16612 = v_7901 & v_8496;
assign v_16614 = v_7877 & v_16613;
assign v_16615 = v_7902 & v_8344;
assign v_16617 = v_7571 & v_16616;
assign v_16618 = v_7607 & v_8212;
assign v_16620 = v_7572 & v_16619;
assign v_16621 = v_7608 & v_8056;
assign v_16623 = v_7288 & v_16622;
assign v_16624 = v_7315 & v_7924;
assign v_16626 = v_7289 & v_16625;
assign v_16627 = v_7316 & v_7774;
assign v_16629 = v_6997 & v_16628;
assign v_16630 = v_7025 & v_7642;
assign v_16632 = v_6998 & v_16631;
assign v_16633 = v_7026 & v_7470;
assign v_16635 = v_6716 & v_16634;
assign v_16636 = v_6741 & v_7338;
assign v_16638 = v_6717 & v_16637;
assign v_16639 = v_6742 & v_7184;
assign v_16641 = v_6419 & v_16640;
assign v_16642 = v_6451 & v_7052;
assign v_16644 = v_6420 & v_16643;
assign v_16645 = v_6452 & v_6896;
assign v_16647 = v_6137 & v_16646;
assign v_16648 = v_6163 & v_6764;
assign v_16650 = v_6138 & v_16649;
assign v_16651 = v_6164 & v_6614;
assign v_16653 = v_5847 & v_16652;
assign v_16654 = v_5875 & v_6482;
assign v_16656 = v_5848 & v_16655;
assign v_16657 = v_5876 & v_6318;
assign v_16659 = v_5566 & v_16658;
assign v_16660 = v_5591 & v_6186;
assign v_16662 = v_5567 & v_16661;
assign v_16663 = v_5592 & v_6034;
assign v_16665 = v_5253 & v_16664;
assign v_16666 = v_5293 & v_5902;
assign v_16668 = v_5254 & v_16667;
assign v_16669 = v_5294 & v_5746;
assign v_16671 = v_4969 & v_16670;
assign v_16672 = v_4997 & v_5614;
assign v_16674 = v_4970 & v_16673;
assign v_16675 = v_4998 & v_5464;
assign v_16677 = v_4677 & v_16676;
assign v_16678 = v_4705 & v_5332;
assign v_16680 = v_4678 & v_16679;
assign v_16681 = v_4706 & v_5152;
assign v_16683 = v_4396 & v_16682;
assign v_16684 = v_4421 & v_5020;
assign v_16686 = v_4397 & v_16685;
assign v_16687 = v_4422 & v_4864;
assign v_16689 = v_4099 & v_16688;
assign v_16690 = v_4131 & v_4732;
assign v_16692 = v_4100 & v_16691;
assign v_16693 = v_4132 & v_4576;
assign v_16695 = v_3817 & v_16694;
assign v_16696 = v_3843 & v_4444;
assign v_16698 = v_3818 & v_16697;
assign v_16699 = v_3844 & v_4294;
assign v_16701 = v_3527 & v_16700;
assign v_16702 = v_3555 & v_4162;
assign v_16704 = v_3528 & v_16703;
assign v_16705 = v_3556 & v_3998;
assign v_16707 = v_3246 & v_16706;
assign v_16708 = v_3271 & v_3866;
assign v_16710 = v_3247 & v_16709;
assign v_16711 = v_3272 & v_3714;
assign v_16713 = v_2941 & v_16712;
assign v_16714 = v_2977 & v_3582;
assign v_16716 = v_2942 & v_16715;
assign v_16717 = v_2978 & v_3426;
assign v_16719 = v_2658 & v_16718;
assign v_16720 = v_2685 & v_3294;
assign v_16722 = v_2659 & v_16721;
assign v_16723 = v_2686 & v_3144;
assign v_16725 = v_2367 & v_16724;
assign v_16726 = v_2395 & v_3012;
assign v_16728 = v_2368 & v_16727;
assign v_16729 = v_2396 & v_2840;
assign v_16731 = v_2086 & v_16730;
assign v_16732 = v_2111 & v_2708;
assign v_16734 = v_2087 & v_16733;
assign v_16735 = v_2112 & v_2554;
assign v_16737 = v_1789 & v_16736;
assign v_16738 = v_1821 & v_2422;
assign v_16740 = v_1790 & v_16739;
assign v_16741 = v_1822 & v_2266;
assign v_16743 = v_1507 & v_16742;
assign v_16744 = v_1533 & v_2134;
assign v_16746 = v_1508 & v_16745;
assign v_16747 = v_1534 & v_1984;
assign v_16749 = v_1217 & v_16748;
assign v_16750 = v_1245 & v_1852;
assign v_16752 = v_1218 & v_16751;
assign v_16753 = v_1246 & v_1688;
assign v_16755 = v_936 & v_16754;
assign v_16756 = v_961 & v_1556;
assign v_16758 = v_937 & v_16757;
assign v_16759 = v_962 & v_1404;
assign v_16761 = v_92 & v_16760;
assign v_16762 = v_591 & v_1272;
assign v_16764 = v_94 & v_16763;
assign v_16765 = v_593 & v_1116;
assign v_16767 = v_806 & v_16766;
assign v_16768 = v_823 & v_984;
assign v_16770 = v_9026 & v_9753;
assign v_16771 = v_9051 & v_9604;
assign v_16773 = v_9027 & v_16772;
assign v_16774 = v_9052 & v_9463;
assign v_16776 = v_8729 & v_16775;
assign v_16777 = v_8761 & v_9311;
assign v_16779 = v_8730 & v_16778;
assign v_16780 = v_8762 & v_9175;
assign v_16782 = v_8447 & v_16781;
assign v_16783 = v_8473 & v_9030;
assign v_16785 = v_8448 & v_16784;
assign v_16786 = v_8474 & v_8893;
assign v_16788 = v_8157 & v_16787;
assign v_16789 = v_8185 & v_8733;
assign v_16791 = v_8158 & v_16790;
assign v_16792 = v_8186 & v_8597;
assign v_16794 = v_7876 & v_16793;
assign v_16795 = v_7901 & v_8451;
assign v_16797 = v_7877 & v_16796;
assign v_16798 = v_7902 & v_8313;
assign v_16800 = v_7571 & v_16799;
assign v_16801 = v_7607 & v_8161;
assign v_16803 = v_7572 & v_16802;
assign v_16804 = v_7608 & v_8025;
assign v_16806 = v_7288 & v_16805;
assign v_16807 = v_7315 & v_7880;
assign v_16809 = v_7289 & v_16808;
assign v_16810 = v_7316 & v_7743;
assign v_16812 = v_6997 & v_16811;
assign v_16813 = v_7025 & v_7575;
assign v_16815 = v_6998 & v_16814;
assign v_16816 = v_7026 & v_7439;
assign v_16818 = v_6716 & v_16817;
assign v_16819 = v_6741 & v_7292;
assign v_16821 = v_6717 & v_16820;
assign v_16822 = v_6742 & v_7153;
assign v_16824 = v_6419 & v_16823;
assign v_16825 = v_6451 & v_7001;
assign v_16827 = v_6420 & v_16826;
assign v_16828 = v_6452 & v_6865;
assign v_16830 = v_6137 & v_16829;
assign v_16831 = v_6163 & v_6720;
assign v_16833 = v_6138 & v_16832;
assign v_16834 = v_6164 & v_6583;
assign v_16836 = v_5847 & v_16835;
assign v_16837 = v_5875 & v_6423;
assign v_16839 = v_5848 & v_16838;
assign v_16840 = v_5876 & v_6287;
assign v_16842 = v_5566 & v_16841;
assign v_16843 = v_5591 & v_6141;
assign v_16845 = v_5567 & v_16844;
assign v_16846 = v_5592 & v_6003;
assign v_16848 = v_5253 & v_16847;
assign v_16849 = v_5293 & v_5851;
assign v_16851 = v_5254 & v_16850;
assign v_16852 = v_5294 & v_5715;
assign v_16854 = v_4969 & v_16853;
assign v_16855 = v_4997 & v_5570;
assign v_16857 = v_4970 & v_16856;
assign v_16858 = v_4998 & v_5433;
assign v_16860 = v_4677 & v_16859;
assign v_16861 = v_4705 & v_5257;
assign v_16863 = v_4678 & v_16862;
assign v_16864 = v_4706 & v_5121;
assign v_16866 = v_4396 & v_16865;
assign v_16867 = v_4421 & v_4973;
assign v_16869 = v_4397 & v_16868;
assign v_16870 = v_4422 & v_4833;
assign v_16872 = v_4099 & v_16871;
assign v_16873 = v_4131 & v_4681;
assign v_16875 = v_4100 & v_16874;
assign v_16876 = v_4132 & v_4545;
assign v_16878 = v_3817 & v_16877;
assign v_16879 = v_3843 & v_4400;
assign v_16881 = v_3818 & v_16880;
assign v_16882 = v_3844 & v_4263;
assign v_16884 = v_3527 & v_16883;
assign v_16885 = v_3555 & v_4103;
assign v_16887 = v_3528 & v_16886;
assign v_16888 = v_3556 & v_3967;
assign v_16890 = v_3246 & v_16889;
assign v_16891 = v_3271 & v_3821;
assign v_16893 = v_3247 & v_16892;
assign v_16894 = v_3272 & v_3683;
assign v_16896 = v_2941 & v_16895;
assign v_16897 = v_2977 & v_3531;
assign v_16899 = v_2942 & v_16898;
assign v_16900 = v_2978 & v_3395;
assign v_16902 = v_2658 & v_16901;
assign v_16903 = v_2685 & v_3250;
assign v_16905 = v_2659 & v_16904;
assign v_16906 = v_2686 & v_3113;
assign v_16908 = v_2367 & v_16907;
assign v_16909 = v_2395 & v_2945;
assign v_16911 = v_2368 & v_16910;
assign v_16912 = v_2396 & v_2809;
assign v_16914 = v_2086 & v_16913;
assign v_16915 = v_2111 & v_2662;
assign v_16917 = v_2087 & v_16916;
assign v_16918 = v_2112 & v_2523;
assign v_16920 = v_1789 & v_16919;
assign v_16921 = v_1821 & v_2371;
assign v_16923 = v_1790 & v_16922;
assign v_16924 = v_1822 & v_2235;
assign v_16926 = v_1507 & v_16925;
assign v_16927 = v_1533 & v_2090;
assign v_16929 = v_1508 & v_16928;
assign v_16930 = v_1534 & v_1953;
assign v_16932 = v_1217 & v_16931;
assign v_16933 = v_1245 & v_1793;
assign v_16935 = v_1218 & v_16934;
assign v_16936 = v_1246 & v_1657;
assign v_16938 = v_936 & v_16937;
assign v_16939 = v_961 & v_1511;
assign v_16941 = v_937 & v_16940;
assign v_16942 = v_962 & v_1373;
assign v_16944 = v_92 & v_16943;
assign v_16945 = v_591 & v_1221;
assign v_16947 = v_94 & v_16946;
assign v_16948 = v_593 & v_1085;
assign v_16950 = v_806 & v_16949;
assign v_16951 = v_823 & v_940;
assign v_16954 = v_9026 & v_9796;
assign v_16955 = v_9051 & v_9664;
assign v_16957 = v_9027 & v_16956;
assign v_16958 = v_9052 & v_9506;
assign v_16960 = v_8729 & v_16959;
assign v_16961 = v_8761 & v_9374;
assign v_16963 = v_8730 & v_16962;
assign v_16964 = v_8762 & v_9218;
assign v_16966 = v_8447 & v_16965;
assign v_16967 = v_8473 & v_9086;
assign v_16969 = v_8448 & v_16968;
assign v_16970 = v_8474 & v_8936;
assign v_16972 = v_8157 & v_16971;
assign v_16973 = v_8185 & v_8804;
assign v_16975 = v_8158 & v_16974;
assign v_16976 = v_8186 & v_8640;
assign v_16978 = v_7876 & v_16977;
assign v_16979 = v_7901 & v_8508;
assign v_16981 = v_7877 & v_16980;
assign v_16982 = v_7902 & v_8356;
assign v_16984 = v_7571 & v_16983;
assign v_16985 = v_7607 & v_8224;
assign v_16987 = v_7572 & v_16986;
assign v_16988 = v_7608 & v_8068;
assign v_16990 = v_7288 & v_16989;
assign v_16991 = v_7315 & v_7936;
assign v_16993 = v_7289 & v_16992;
assign v_16994 = v_7316 & v_7786;
assign v_16996 = v_6997 & v_16995;
assign v_16997 = v_7025 & v_7654;
assign v_16999 = v_6998 & v_16998;
assign v_17000 = v_7026 & v_7482;
assign v_17002 = v_6716 & v_17001;
assign v_17003 = v_6741 & v_7350;
assign v_17005 = v_6717 & v_17004;
assign v_17006 = v_6742 & v_7196;
assign v_17008 = v_6419 & v_17007;
assign v_17009 = v_6451 & v_7064;
assign v_17011 = v_6420 & v_17010;
assign v_17012 = v_6452 & v_6908;
assign v_17014 = v_6137 & v_17013;
assign v_17015 = v_6163 & v_6776;
assign v_17017 = v_6138 & v_17016;
assign v_17018 = v_6164 & v_6626;
assign v_17020 = v_5847 & v_17019;
assign v_17021 = v_5875 & v_6494;
assign v_17023 = v_5848 & v_17022;
assign v_17024 = v_5876 & v_6330;
assign v_17026 = v_5566 & v_17025;
assign v_17027 = v_5591 & v_6198;
assign v_17029 = v_5567 & v_17028;
assign v_17030 = v_5592 & v_6046;
assign v_17032 = v_5253 & v_17031;
assign v_17033 = v_5293 & v_5914;
assign v_17035 = v_5254 & v_17034;
assign v_17036 = v_5294 & v_5758;
assign v_17038 = v_4969 & v_17037;
assign v_17039 = v_4997 & v_5626;
assign v_17041 = v_4970 & v_17040;
assign v_17042 = v_4998 & v_5476;
assign v_17044 = v_4677 & v_17043;
assign v_17045 = v_4705 & v_5344;
assign v_17047 = v_4678 & v_17046;
assign v_17048 = v_4706 & v_5164;
assign v_17050 = v_4396 & v_17049;
assign v_17051 = v_4421 & v_5032;
assign v_17053 = v_4397 & v_17052;
assign v_17054 = v_4422 & v_4876;
assign v_17056 = v_4099 & v_17055;
assign v_17057 = v_4131 & v_4744;
assign v_17059 = v_4100 & v_17058;
assign v_17060 = v_4132 & v_4588;
assign v_17062 = v_3817 & v_17061;
assign v_17063 = v_3843 & v_4456;
assign v_17065 = v_3818 & v_17064;
assign v_17066 = v_3844 & v_4306;
assign v_17068 = v_3527 & v_17067;
assign v_17069 = v_3555 & v_4174;
assign v_17071 = v_3528 & v_17070;
assign v_17072 = v_3556 & v_4010;
assign v_17074 = v_3246 & v_17073;
assign v_17075 = v_3271 & v_3878;
assign v_17077 = v_3247 & v_17076;
assign v_17078 = v_3272 & v_3726;
assign v_17080 = v_2941 & v_17079;
assign v_17081 = v_2977 & v_3594;
assign v_17083 = v_2942 & v_17082;
assign v_17084 = v_2978 & v_3438;
assign v_17086 = v_2658 & v_17085;
assign v_17087 = v_2685 & v_3306;
assign v_17089 = v_2659 & v_17088;
assign v_17090 = v_2686 & v_3156;
assign v_17092 = v_2367 & v_17091;
assign v_17093 = v_2395 & v_3024;
assign v_17095 = v_2368 & v_17094;
assign v_17096 = v_2396 & v_2852;
assign v_17098 = v_2086 & v_17097;
assign v_17099 = v_2111 & v_2720;
assign v_17101 = v_2087 & v_17100;
assign v_17102 = v_2112 & v_2566;
assign v_17104 = v_1789 & v_17103;
assign v_17105 = v_1821 & v_2434;
assign v_17107 = v_1790 & v_17106;
assign v_17108 = v_1822 & v_2278;
assign v_17110 = v_1507 & v_17109;
assign v_17111 = v_1533 & v_2146;
assign v_17113 = v_1508 & v_17112;
assign v_17114 = v_1534 & v_1996;
assign v_17116 = v_1217 & v_17115;
assign v_17117 = v_1245 & v_1864;
assign v_17119 = v_1218 & v_17118;
assign v_17120 = v_1246 & v_1700;
assign v_17122 = v_936 & v_17121;
assign v_17123 = v_961 & v_1568;
assign v_17125 = v_937 & v_17124;
assign v_17126 = v_962 & v_1416;
assign v_17128 = v_92 & v_17127;
assign v_17129 = v_591 & v_1284;
assign v_17131 = v_94 & v_17130;
assign v_17132 = v_593 & v_1128;
assign v_17134 = v_806 & v_17133;
assign v_17135 = v_823 & v_996;
assign v_17138 = v_9026 & v_9808;
assign v_17139 = v_9051 & v_9676;
assign v_17141 = v_9027 & v_17140;
assign v_17142 = v_9052 & v_9518;
assign v_17144 = v_8729 & v_17143;
assign v_17145 = v_8761 & v_9386;
assign v_17147 = v_8730 & v_17146;
assign v_17148 = v_8762 & v_9230;
assign v_17150 = v_8447 & v_17149;
assign v_17151 = v_8473 & v_9098;
assign v_17153 = v_8448 & v_17152;
assign v_17154 = v_8474 & v_8948;
assign v_17156 = v_8157 & v_17155;
assign v_17157 = v_8185 & v_8816;
assign v_17159 = v_8158 & v_17158;
assign v_17160 = v_8186 & v_8652;
assign v_17162 = v_7876 & v_17161;
assign v_17163 = v_7901 & v_8520;
assign v_17165 = v_7877 & v_17164;
assign v_17166 = v_7902 & v_8368;
assign v_17168 = v_7571 & v_17167;
assign v_17169 = v_7607 & v_8236;
assign v_17171 = v_7572 & v_17170;
assign v_17172 = v_7608 & v_8080;
assign v_17174 = v_7288 & v_17173;
assign v_17175 = v_7315 & v_7948;
assign v_17177 = v_7289 & v_17176;
assign v_17178 = v_7316 & v_7798;
assign v_17180 = v_6997 & v_17179;
assign v_17181 = v_7025 & v_7666;
assign v_17183 = v_6998 & v_17182;
assign v_17184 = v_7026 & v_7494;
assign v_17186 = v_6716 & v_17185;
assign v_17187 = v_6741 & v_7362;
assign v_17189 = v_6717 & v_17188;
assign v_17190 = v_6742 & v_7208;
assign v_17192 = v_6419 & v_17191;
assign v_17193 = v_6451 & v_7076;
assign v_17195 = v_6420 & v_17194;
assign v_17196 = v_6452 & v_6920;
assign v_17198 = v_6137 & v_17197;
assign v_17199 = v_6163 & v_6788;
assign v_17201 = v_6138 & v_17200;
assign v_17202 = v_6164 & v_6638;
assign v_17204 = v_5847 & v_17203;
assign v_17205 = v_5875 & v_6506;
assign v_17207 = v_5848 & v_17206;
assign v_17208 = v_5876 & v_6342;
assign v_17210 = v_5566 & v_17209;
assign v_17211 = v_5591 & v_6210;
assign v_17213 = v_5567 & v_17212;
assign v_17214 = v_5592 & v_6058;
assign v_17216 = v_5253 & v_17215;
assign v_17217 = v_5293 & v_5926;
assign v_17219 = v_5254 & v_17218;
assign v_17220 = v_5294 & v_5770;
assign v_17222 = v_4969 & v_17221;
assign v_17223 = v_4997 & v_5638;
assign v_17225 = v_4970 & v_17224;
assign v_17226 = v_4998 & v_5488;
assign v_17228 = v_4677 & v_17227;
assign v_17229 = v_4705 & v_5356;
assign v_17231 = v_4678 & v_17230;
assign v_17232 = v_4706 & v_5176;
assign v_17234 = v_4396 & v_17233;
assign v_17235 = v_4421 & v_5044;
assign v_17237 = v_4397 & v_17236;
assign v_17238 = v_4422 & v_4888;
assign v_17240 = v_4099 & v_17239;
assign v_17241 = v_4131 & v_4756;
assign v_17243 = v_4100 & v_17242;
assign v_17244 = v_4132 & v_4600;
assign v_17246 = v_3817 & v_17245;
assign v_17247 = v_3843 & v_4468;
assign v_17249 = v_3818 & v_17248;
assign v_17250 = v_3844 & v_4318;
assign v_17252 = v_3527 & v_17251;
assign v_17253 = v_3555 & v_4186;
assign v_17255 = v_3528 & v_17254;
assign v_17256 = v_3556 & v_4022;
assign v_17258 = v_3246 & v_17257;
assign v_17259 = v_3271 & v_3890;
assign v_17261 = v_3247 & v_17260;
assign v_17262 = v_3272 & v_3738;
assign v_17264 = v_2941 & v_17263;
assign v_17265 = v_2977 & v_3606;
assign v_17267 = v_2942 & v_17266;
assign v_17268 = v_2978 & v_3450;
assign v_17270 = v_2658 & v_17269;
assign v_17271 = v_2685 & v_3318;
assign v_17273 = v_2659 & v_17272;
assign v_17274 = v_2686 & v_3168;
assign v_17276 = v_2367 & v_17275;
assign v_17277 = v_2395 & v_3036;
assign v_17279 = v_2368 & v_17278;
assign v_17280 = v_2396 & v_2864;
assign v_17282 = v_2086 & v_17281;
assign v_17283 = v_2111 & v_2732;
assign v_17285 = v_2087 & v_17284;
assign v_17286 = v_2112 & v_2578;
assign v_17288 = v_1789 & v_17287;
assign v_17289 = v_1821 & v_2446;
assign v_17291 = v_1790 & v_17290;
assign v_17292 = v_1822 & v_2290;
assign v_17294 = v_1507 & v_17293;
assign v_17295 = v_1533 & v_2158;
assign v_17297 = v_1508 & v_17296;
assign v_17298 = v_1534 & v_2008;
assign v_17300 = v_1217 & v_17299;
assign v_17301 = v_1245 & v_1876;
assign v_17303 = v_1218 & v_17302;
assign v_17304 = v_1246 & v_1712;
assign v_17306 = v_936 & v_17305;
assign v_17307 = v_961 & v_1580;
assign v_17309 = v_937 & v_17308;
assign v_17310 = v_962 & v_1428;
assign v_17312 = v_92 & v_17311;
assign v_17313 = v_591 & v_1296;
assign v_17315 = v_94 & v_17314;
assign v_17316 = v_593 & v_1140;
assign v_17318 = v_806 & v_17317;
assign v_17319 = v_823 & v_1008;
assign v_17322 = v_9026 & v_9820;
assign v_17323 = v_9051 & v_9688;
assign v_17325 = v_9027 & v_17324;
assign v_17326 = v_9052 & v_9530;
assign v_17328 = v_8729 & v_17327;
assign v_17329 = v_8761 & v_9398;
assign v_17331 = v_8730 & v_17330;
assign v_17332 = v_8762 & v_9242;
assign v_17334 = v_8447 & v_17333;
assign v_17335 = v_8473 & v_9110;
assign v_17337 = v_8448 & v_17336;
assign v_17338 = v_8474 & v_8960;
assign v_17340 = v_8157 & v_17339;
assign v_17341 = v_8185 & v_8828;
assign v_17343 = v_8158 & v_17342;
assign v_17344 = v_8186 & v_8664;
assign v_17346 = v_7876 & v_17345;
assign v_17347 = v_7901 & v_8532;
assign v_17349 = v_7877 & v_17348;
assign v_17350 = v_7902 & v_8380;
assign v_17352 = v_7571 & v_17351;
assign v_17353 = v_7607 & v_8248;
assign v_17355 = v_7572 & v_17354;
assign v_17356 = v_7608 & v_8092;
assign v_17358 = v_7288 & v_17357;
assign v_17359 = v_7315 & v_7960;
assign v_17361 = v_7289 & v_17360;
assign v_17362 = v_7316 & v_7810;
assign v_17364 = v_6997 & v_17363;
assign v_17365 = v_7025 & v_7678;
assign v_17367 = v_6998 & v_17366;
assign v_17368 = v_7026 & v_7506;
assign v_17370 = v_6716 & v_17369;
assign v_17371 = v_6741 & v_7374;
assign v_17373 = v_6717 & v_17372;
assign v_17374 = v_6742 & v_7220;
assign v_17376 = v_6419 & v_17375;
assign v_17377 = v_6451 & v_7088;
assign v_17379 = v_6420 & v_17378;
assign v_17380 = v_6452 & v_6932;
assign v_17382 = v_6137 & v_17381;
assign v_17383 = v_6163 & v_6800;
assign v_17385 = v_6138 & v_17384;
assign v_17386 = v_6164 & v_6650;
assign v_17388 = v_5847 & v_17387;
assign v_17389 = v_5875 & v_6518;
assign v_17391 = v_5848 & v_17390;
assign v_17392 = v_5876 & v_6354;
assign v_17394 = v_5566 & v_17393;
assign v_17395 = v_5591 & v_6222;
assign v_17397 = v_5567 & v_17396;
assign v_17398 = v_5592 & v_6070;
assign v_17400 = v_5253 & v_17399;
assign v_17401 = v_5293 & v_5938;
assign v_17403 = v_5254 & v_17402;
assign v_17404 = v_5294 & v_5782;
assign v_17406 = v_4969 & v_17405;
assign v_17407 = v_4997 & v_5650;
assign v_17409 = v_4970 & v_17408;
assign v_17410 = v_4998 & v_5500;
assign v_17412 = v_4677 & v_17411;
assign v_17413 = v_4705 & v_5368;
assign v_17415 = v_4678 & v_17414;
assign v_17416 = v_4706 & v_5188;
assign v_17418 = v_4396 & v_17417;
assign v_17419 = v_4421 & v_5056;
assign v_17421 = v_4397 & v_17420;
assign v_17422 = v_4422 & v_4900;
assign v_17424 = v_4099 & v_17423;
assign v_17425 = v_4131 & v_4768;
assign v_17427 = v_4100 & v_17426;
assign v_17428 = v_4132 & v_4612;
assign v_17430 = v_3817 & v_17429;
assign v_17431 = v_3843 & v_4480;
assign v_17433 = v_3818 & v_17432;
assign v_17434 = v_3844 & v_4330;
assign v_17436 = v_3527 & v_17435;
assign v_17437 = v_3555 & v_4198;
assign v_17439 = v_3528 & v_17438;
assign v_17440 = v_3556 & v_4034;
assign v_17442 = v_3246 & v_17441;
assign v_17443 = v_3271 & v_3902;
assign v_17445 = v_3247 & v_17444;
assign v_17446 = v_3272 & v_3750;
assign v_17448 = v_2941 & v_17447;
assign v_17449 = v_2977 & v_3618;
assign v_17451 = v_2942 & v_17450;
assign v_17452 = v_2978 & v_3462;
assign v_17454 = v_2658 & v_17453;
assign v_17455 = v_2685 & v_3330;
assign v_17457 = v_2659 & v_17456;
assign v_17458 = v_2686 & v_3180;
assign v_17460 = v_2367 & v_17459;
assign v_17461 = v_2395 & v_3048;
assign v_17463 = v_2368 & v_17462;
assign v_17464 = v_2396 & v_2876;
assign v_17466 = v_2086 & v_17465;
assign v_17467 = v_2111 & v_2744;
assign v_17469 = v_2087 & v_17468;
assign v_17470 = v_2112 & v_2590;
assign v_17472 = v_1789 & v_17471;
assign v_17473 = v_1821 & v_2458;
assign v_17475 = v_1790 & v_17474;
assign v_17476 = v_1822 & v_2302;
assign v_17478 = v_1507 & v_17477;
assign v_17479 = v_1533 & v_2170;
assign v_17481 = v_1508 & v_17480;
assign v_17482 = v_1534 & v_2020;
assign v_17484 = v_1217 & v_17483;
assign v_17485 = v_1245 & v_1888;
assign v_17487 = v_1218 & v_17486;
assign v_17488 = v_1246 & v_1724;
assign v_17490 = v_936 & v_17489;
assign v_17491 = v_961 & v_1592;
assign v_17493 = v_937 & v_17492;
assign v_17494 = v_962 & v_1440;
assign v_17496 = v_92 & v_17495;
assign v_17497 = v_591 & v_1308;
assign v_17499 = v_94 & v_17498;
assign v_17500 = v_593 & v_1152;
assign v_17502 = v_806 & v_17501;
assign v_17503 = v_823 & v_1020;
assign v_17506 = v_9026 & v_9832;
assign v_17507 = v_9051 & v_9700;
assign v_17509 = v_9027 & v_17508;
assign v_17510 = v_9052 & v_9542;
assign v_17512 = v_8729 & v_17511;
assign v_17513 = v_8761 & v_9410;
assign v_17515 = v_8730 & v_17514;
assign v_17516 = v_8762 & v_9254;
assign v_17518 = v_8447 & v_17517;
assign v_17519 = v_8473 & v_9122;
assign v_17521 = v_8448 & v_17520;
assign v_17522 = v_8474 & v_8972;
assign v_17524 = v_8157 & v_17523;
assign v_17525 = v_8185 & v_8840;
assign v_17527 = v_8158 & v_17526;
assign v_17528 = v_8186 & v_8676;
assign v_17530 = v_7876 & v_17529;
assign v_17531 = v_7901 & v_8544;
assign v_17533 = v_7877 & v_17532;
assign v_17534 = v_7902 & v_8392;
assign v_17536 = v_7571 & v_17535;
assign v_17537 = v_7607 & v_8260;
assign v_17539 = v_7572 & v_17538;
assign v_17540 = v_7608 & v_8104;
assign v_17542 = v_7288 & v_17541;
assign v_17543 = v_7315 & v_7972;
assign v_17545 = v_7289 & v_17544;
assign v_17546 = v_7316 & v_7822;
assign v_17548 = v_6997 & v_17547;
assign v_17549 = v_7025 & v_7690;
assign v_17551 = v_6998 & v_17550;
assign v_17552 = v_7026 & v_7518;
assign v_17554 = v_6716 & v_17553;
assign v_17555 = v_6741 & v_7386;
assign v_17557 = v_6717 & v_17556;
assign v_17558 = v_6742 & v_7232;
assign v_17560 = v_6419 & v_17559;
assign v_17561 = v_6451 & v_7100;
assign v_17563 = v_6420 & v_17562;
assign v_17564 = v_6452 & v_6944;
assign v_17566 = v_6137 & v_17565;
assign v_17567 = v_6163 & v_6812;
assign v_17569 = v_6138 & v_17568;
assign v_17570 = v_6164 & v_6662;
assign v_17572 = v_5847 & v_17571;
assign v_17573 = v_5875 & v_6530;
assign v_17575 = v_5848 & v_17574;
assign v_17576 = v_5876 & v_6366;
assign v_17578 = v_5566 & v_17577;
assign v_17579 = v_5591 & v_6234;
assign v_17581 = v_5567 & v_17580;
assign v_17582 = v_5592 & v_6082;
assign v_17584 = v_5253 & v_17583;
assign v_17585 = v_5293 & v_5950;
assign v_17587 = v_5254 & v_17586;
assign v_17588 = v_5294 & v_5794;
assign v_17590 = v_4969 & v_17589;
assign v_17591 = v_4997 & v_5662;
assign v_17593 = v_4970 & v_17592;
assign v_17594 = v_4998 & v_5512;
assign v_17596 = v_4677 & v_17595;
assign v_17597 = v_4705 & v_5380;
assign v_17599 = v_4678 & v_17598;
assign v_17600 = v_4706 & v_5200;
assign v_17602 = v_4396 & v_17601;
assign v_17603 = v_4421 & v_5068;
assign v_17605 = v_4397 & v_17604;
assign v_17606 = v_4422 & v_4912;
assign v_17608 = v_4099 & v_17607;
assign v_17609 = v_4131 & v_4780;
assign v_17611 = v_4100 & v_17610;
assign v_17612 = v_4132 & v_4624;
assign v_17614 = v_3817 & v_17613;
assign v_17615 = v_3843 & v_4492;
assign v_17617 = v_3818 & v_17616;
assign v_17618 = v_3844 & v_4342;
assign v_17620 = v_3527 & v_17619;
assign v_17621 = v_3555 & v_4210;
assign v_17623 = v_3528 & v_17622;
assign v_17624 = v_3556 & v_4046;
assign v_17626 = v_3246 & v_17625;
assign v_17627 = v_3271 & v_3914;
assign v_17629 = v_3247 & v_17628;
assign v_17630 = v_3272 & v_3762;
assign v_17632 = v_2941 & v_17631;
assign v_17633 = v_2977 & v_3630;
assign v_17635 = v_2942 & v_17634;
assign v_17636 = v_2978 & v_3474;
assign v_17638 = v_2658 & v_17637;
assign v_17639 = v_2685 & v_3342;
assign v_17641 = v_2659 & v_17640;
assign v_17642 = v_2686 & v_3192;
assign v_17644 = v_2367 & v_17643;
assign v_17645 = v_2395 & v_3060;
assign v_17647 = v_2368 & v_17646;
assign v_17648 = v_2396 & v_2888;
assign v_17650 = v_2086 & v_17649;
assign v_17651 = v_2111 & v_2756;
assign v_17653 = v_2087 & v_17652;
assign v_17654 = v_2112 & v_2602;
assign v_17656 = v_1789 & v_17655;
assign v_17657 = v_1821 & v_2470;
assign v_17659 = v_1790 & v_17658;
assign v_17660 = v_1822 & v_2314;
assign v_17662 = v_1507 & v_17661;
assign v_17663 = v_1533 & v_2182;
assign v_17665 = v_1508 & v_17664;
assign v_17666 = v_1534 & v_2032;
assign v_17668 = v_1217 & v_17667;
assign v_17669 = v_1245 & v_1900;
assign v_17671 = v_1218 & v_17670;
assign v_17672 = v_1246 & v_1736;
assign v_17674 = v_936 & v_17673;
assign v_17675 = v_961 & v_1604;
assign v_17677 = v_937 & v_17676;
assign v_17678 = v_962 & v_1452;
assign v_17680 = v_92 & v_17679;
assign v_17681 = v_591 & v_1320;
assign v_17683 = v_94 & v_17682;
assign v_17684 = v_593 & v_1164;
assign v_17686 = v_806 & v_17685;
assign v_17687 = v_823 & v_1032;
assign v_17690 = v_9026 & v_9844;
assign v_17691 = v_9051 & v_9712;
assign v_17693 = v_9027 & v_17692;
assign v_17694 = v_9052 & v_9554;
assign v_17696 = v_8729 & v_17695;
assign v_17697 = v_8761 & v_9422;
assign v_17699 = v_8730 & v_17698;
assign v_17700 = v_8762 & v_9266;
assign v_17702 = v_8447 & v_17701;
assign v_17703 = v_8473 & v_9134;
assign v_17705 = v_8448 & v_17704;
assign v_17706 = v_8474 & v_8984;
assign v_17708 = v_8157 & v_17707;
assign v_17709 = v_8185 & v_8852;
assign v_17711 = v_8158 & v_17710;
assign v_17712 = v_8186 & v_8688;
assign v_17714 = v_7876 & v_17713;
assign v_17715 = v_7901 & v_8556;
assign v_17717 = v_7877 & v_17716;
assign v_17718 = v_7902 & v_8404;
assign v_17720 = v_7571 & v_17719;
assign v_17721 = v_7607 & v_8272;
assign v_17723 = v_7572 & v_17722;
assign v_17724 = v_7608 & v_8116;
assign v_17726 = v_7288 & v_17725;
assign v_17727 = v_7315 & v_7984;
assign v_17729 = v_7289 & v_17728;
assign v_17730 = v_7316 & v_7834;
assign v_17732 = v_6997 & v_17731;
assign v_17733 = v_7025 & v_7702;
assign v_17735 = v_6998 & v_17734;
assign v_17736 = v_7026 & v_7530;
assign v_17738 = v_6716 & v_17737;
assign v_17739 = v_6741 & v_7398;
assign v_17741 = v_6717 & v_17740;
assign v_17742 = v_6742 & v_7244;
assign v_17744 = v_6419 & v_17743;
assign v_17745 = v_6451 & v_7112;
assign v_17747 = v_6420 & v_17746;
assign v_17748 = v_6452 & v_6956;
assign v_17750 = v_6137 & v_17749;
assign v_17751 = v_6163 & ~v_6824;
assign v_17753 = v_6138 & v_17752;
assign v_17754 = v_6164 & v_6674;
assign v_17756 = v_5847 & v_17755;
assign v_17757 = v_5875 & v_6542;
assign v_17759 = v_5848 & v_17758;
assign v_17760 = v_5876 & v_6378;
assign v_17762 = v_5566 & v_17761;
assign v_17763 = v_5591 & v_6246;
assign v_17765 = v_5567 & v_17764;
assign v_17766 = v_5592 & ~v_6094;
assign v_17768 = v_5253 & v_17767;
assign v_17769 = v_5293 & v_5962;
assign v_17771 = v_5254 & v_17770;
assign v_17772 = v_5294 & ~v_5806;
assign v_17774 = v_4969 & v_17773;
assign v_17775 = v_4997 & v_5674;
assign v_17777 = v_4970 & v_17776;
assign v_17778 = v_4998 & v_5524;
assign v_17780 = v_4677 & v_17779;
assign v_17781 = v_4705 & v_5392;
assign v_17783 = v_4678 & v_17782;
assign v_17784 = v_4706 & v_5212;
assign v_17786 = v_4396 & v_17785;
assign v_17787 = v_4421 & v_5080;
assign v_17789 = v_4397 & v_17788;
assign v_17790 = v_4422 & v_4924;
assign v_17792 = v_4099 & v_17791;
assign v_17793 = v_4131 & v_4792;
assign v_17795 = v_4100 & v_17794;
assign v_17796 = v_4132 & v_4636;
assign v_17798 = v_3817 & v_17797;
assign v_17799 = v_3843 & v_4504;
assign v_17801 = v_3818 & v_17800;
assign v_17802 = v_3844 & v_4354;
assign v_17804 = v_3527 & v_17803;
assign v_17805 = v_3555 & v_4222;
assign v_17807 = v_3528 & v_17806;
assign v_17808 = v_3556 & v_4058;
assign v_17810 = v_3246 & v_17809;
assign v_17811 = v_3271 & v_3926;
assign v_17813 = v_3247 & v_17812;
assign v_17814 = v_3272 & v_3774;
assign v_17816 = v_2941 & v_17815;
assign v_17817 = v_2977 & v_3642;
assign v_17819 = v_2942 & v_17818;
assign v_17820 = v_2978 & v_3486;
assign v_17822 = v_2658 & v_17821;
assign v_17823 = v_2685 & v_3354;
assign v_17825 = v_2659 & v_17824;
assign v_17826 = v_2686 & ~v_3204;
assign v_17828 = v_2367 & v_17827;
assign v_17829 = v_2395 & v_3072;
assign v_17831 = v_2368 & v_17830;
assign v_17832 = v_2396 & v_2900;
assign v_17834 = v_2086 & v_17833;
assign v_17835 = v_2111 & v_2768;
assign v_17837 = v_2087 & v_17836;
assign v_17838 = v_2112 & v_2614;
assign v_17840 = v_1789 & v_17839;
assign v_17841 = v_1821 & v_2482;
assign v_17843 = v_1790 & v_17842;
assign v_17844 = v_1822 & v_2326;
assign v_17846 = v_1507 & v_17845;
assign v_17847 = v_1533 & v_2194;
assign v_17849 = v_1508 & v_17848;
assign v_17850 = v_1534 & v_2044;
assign v_17852 = v_1217 & v_17851;
assign v_17853 = v_1245 & v_1912;
assign v_17855 = v_1218 & v_17854;
assign v_17856 = v_1246 & v_1748;
assign v_17858 = v_936 & v_17857;
assign v_17859 = v_961 & v_1616;
assign v_17861 = v_937 & v_17860;
assign v_17862 = v_962 & v_1464;
assign v_17864 = v_92 & v_17863;
assign v_17865 = v_591 & v_1332;
assign v_17867 = v_94 & v_17866;
assign v_17868 = v_593 & v_1176;
assign v_17870 = v_806 & v_17869;
assign v_17871 = v_823 & v_1044;
assign v_17874 = v_9026 & ~v_9872;
assign v_17875 = v_9051 & ~v_9740;
assign v_17877 = v_9027 & v_17876;
assign v_17878 = v_9052 & ~v_9582;
assign v_17880 = v_8729 & v_17879;
assign v_17881 = v_8761 & ~v_9450;
assign v_17883 = v_8730 & v_17882;
assign v_17884 = v_8762 & ~v_9294;
assign v_17886 = v_8447 & v_17885;
assign v_17887 = v_8473 & ~v_9162;
assign v_17889 = v_8448 & v_17888;
assign v_17890 = v_8474 & ~v_9012;
assign v_17892 = v_8157 & v_17891;
assign v_17893 = v_8185 & ~v_8880;
assign v_17895 = v_8158 & v_17894;
assign v_17896 = v_8186 & ~v_8716;
assign v_17898 = v_7876 & v_17897;
assign v_17899 = v_7901 & ~v_8584;
assign v_17901 = v_7877 & v_17900;
assign v_17902 = v_7902 & v_8432;
assign v_17904 = v_7571 & v_17903;
assign v_17905 = v_7607 & v_8300;
assign v_17907 = v_7572 & v_17906;
assign v_17908 = v_7608 & v_8144;
assign v_17910 = v_7288 & v_17909;
assign v_17911 = v_7315 & ~v_8012;
assign v_17913 = v_7289 & v_17912;
assign v_17914 = v_7316 & ~v_7862;
assign v_17916 = v_6997 & v_17915;
assign v_17917 = v_7025 & ~v_7730;
assign v_17919 = v_6998 & v_17918;
assign v_17920 = v_7026 & ~v_7558;
assign v_17922 = v_6716 & v_17921;
assign v_17923 = v_6741 & ~v_7426;
assign v_17925 = v_6717 & v_17924;
assign v_17926 = v_6742 & v_7272;
assign v_17928 = v_6419 & v_17927;
assign v_17929 = v_6451 & ~v_7140;
assign v_17931 = v_6420 & v_17930;
assign v_17932 = v_6452 & v_6984;
assign v_17934 = v_6137 & v_17933;
assign v_17935 = v_6163 & v_6852;
assign v_17937 = v_6138 & v_17936;
assign v_17938 = v_6164 & v_6702;
assign v_17940 = v_5847 & v_17939;
assign v_17941 = v_5875 & ~v_6570;
assign v_17943 = v_5848 & v_17942;
assign v_17944 = v_5876 & ~v_6406;
assign v_17946 = v_5566 & v_17945;
assign v_17947 = v_5591 & v_6274;
assign v_17949 = v_5567 & v_17948;
assign v_17950 = v_5592 & v_6122;
assign v_17952 = v_5253 & v_17951;
assign v_17953 = v_5293 & v_5990;
assign v_17955 = v_5254 & v_17954;
assign v_17956 = v_5294 & v_5834;
assign v_17958 = v_4969 & v_17957;
assign v_17959 = v_4997 & v_5702;
assign v_17961 = v_4970 & v_17960;
assign v_17962 = v_4998 & v_5552;
assign v_17964 = v_4677 & v_17963;
assign v_17965 = v_4705 & ~v_5420;
assign v_17967 = v_4678 & v_17966;
assign v_17968 = v_4706 & ~v_5240;
assign v_17970 = v_4396 & v_17969;
assign v_17971 = v_4421 & v_5108;
assign v_17973 = v_4397 & v_17972;
assign v_17974 = v_4422 & v_4952;
assign v_17976 = v_4099 & v_17975;
assign v_17977 = v_4131 & v_4820;
assign v_17979 = v_4100 & v_17978;
assign v_17980 = v_4132 & v_4664;
assign v_17982 = v_3817 & v_17981;
assign v_17983 = v_3843 & v_4532;
assign v_17985 = v_3818 & v_17984;
assign v_17986 = v_3844 & v_4382;
assign v_17988 = v_3527 & v_17987;
assign v_17989 = v_3555 & ~v_4250;
assign v_17991 = v_3528 & v_17990;
assign v_17992 = v_3556 & ~v_4086;
assign v_17994 = v_3246 & v_17993;
assign v_17995 = v_3271 & ~v_3954;
assign v_17997 = v_3247 & v_17996;
assign v_17998 = v_3272 & ~v_3802;
assign v_18000 = v_2941 & v_17999;
assign v_18001 = v_2977 & ~v_3670;
assign v_18003 = v_2942 & v_18002;
assign v_18004 = v_2978 & v_3514;
assign v_18006 = v_2658 & v_18005;
assign v_18007 = v_2685 & ~v_3382;
assign v_18009 = v_2659 & v_18008;
assign v_18010 = v_2686 & v_3232;
assign v_18012 = v_2367 & v_18011;
assign v_18013 = v_2395 & ~v_3100;
assign v_18015 = v_2368 & v_18014;
assign v_18016 = v_2396 & ~v_2928;
assign v_18018 = v_2086 & v_18017;
assign v_18019 = v_2111 & ~v_2796;
assign v_18021 = v_2087 & v_18020;
assign v_18022 = v_2112 & ~v_2642;
assign v_18024 = v_1789 & v_18023;
assign v_18025 = v_1821 & ~v_2510;
assign v_18027 = v_1790 & v_18026;
assign v_18028 = v_1822 & v_2354;
assign v_18030 = v_1507 & v_18029;
assign v_18031 = v_1533 & v_2222;
assign v_18033 = v_1508 & v_18032;
assign v_18034 = v_1534 & v_2072;
assign v_18036 = v_1217 & v_18035;
assign v_18037 = v_1245 & ~v_1940;
assign v_18039 = v_1218 & v_18038;
assign v_18040 = v_1246 & ~v_1776;
assign v_18042 = v_936 & v_18041;
assign v_18043 = v_961 & ~v_1644;
assign v_18045 = v_937 & v_18044;
assign v_18046 = v_962 & ~v_1492;
assign v_18048 = v_92 & v_18047;
assign v_18049 = v_591 & ~v_1360;
assign v_18051 = v_94 & v_18050;
assign v_18052 = v_593 & ~v_1204;
assign v_18054 = v_806 & v_18053;
assign v_18055 = v_823 & ~v_1072;
assign v_18058 = v_9308 & v_9784;
assign v_18059 = v_9336 & v_9652;
assign v_18061 = v_9026 & v_18060;
assign v_18062 = v_9051 & v_9494;
assign v_18064 = v_9027 & v_18063;
assign v_18065 = v_9052 & v_9362;
assign v_18067 = v_8729 & v_18066;
assign v_18068 = v_8761 & v_9206;
assign v_18070 = v_8730 & v_18069;
assign v_18071 = v_8762 & v_9074;
assign v_18073 = v_8447 & v_18072;
assign v_18074 = v_8473 & v_8924;
assign v_18076 = v_8448 & v_18075;
assign v_18077 = v_8474 & v_8792;
assign v_18079 = v_8157 & v_18078;
assign v_18080 = v_8185 & v_8628;
assign v_18082 = v_8158 & v_18081;
assign v_18083 = v_8186 & v_8496;
assign v_18085 = v_7876 & v_18084;
assign v_18086 = v_7901 & v_8344;
assign v_18088 = v_7877 & v_18087;
assign v_18089 = v_7902 & v_8212;
assign v_18091 = v_7571 & v_18090;
assign v_18092 = v_7607 & v_8056;
assign v_18094 = v_7572 & v_18093;
assign v_18095 = v_7608 & v_7924;
assign v_18097 = v_7288 & v_18096;
assign v_18098 = v_7315 & v_7774;
assign v_18100 = v_7289 & v_18099;
assign v_18101 = v_7316 & v_7642;
assign v_18103 = v_6997 & v_18102;
assign v_18104 = v_7025 & v_7470;
assign v_18106 = v_6998 & v_18105;
assign v_18107 = v_7026 & v_7338;
assign v_18109 = v_6716 & v_18108;
assign v_18110 = v_6741 & v_7184;
assign v_18112 = v_6717 & v_18111;
assign v_18113 = v_6742 & v_7052;
assign v_18115 = v_6419 & v_18114;
assign v_18116 = v_6451 & v_6896;
assign v_18118 = v_6420 & v_18117;
assign v_18119 = v_6452 & v_6764;
assign v_18121 = v_6137 & v_18120;
assign v_18122 = v_6163 & v_6614;
assign v_18124 = v_6138 & v_18123;
assign v_18125 = v_6164 & v_6482;
assign v_18127 = v_5847 & v_18126;
assign v_18128 = v_5875 & v_6318;
assign v_18130 = v_5848 & v_18129;
assign v_18131 = v_5876 & v_6186;
assign v_18133 = v_5566 & v_18132;
assign v_18134 = v_5591 & v_6034;
assign v_18136 = v_5567 & v_18135;
assign v_18137 = v_5592 & v_5902;
assign v_18139 = v_5253 & v_18138;
assign v_18140 = v_5293 & v_5746;
assign v_18142 = v_5254 & v_18141;
assign v_18143 = v_5294 & v_5614;
assign v_18145 = v_4969 & v_18144;
assign v_18146 = v_4997 & v_5464;
assign v_18148 = v_4970 & v_18147;
assign v_18149 = v_4998 & v_5332;
assign v_18151 = v_4677 & v_18150;
assign v_18152 = v_4705 & v_5152;
assign v_18154 = v_4678 & v_18153;
assign v_18155 = v_4706 & v_5020;
assign v_18157 = v_4396 & v_18156;
assign v_18158 = v_4421 & v_4864;
assign v_18160 = v_4397 & v_18159;
assign v_18161 = v_4422 & v_4732;
assign v_18163 = v_4099 & v_18162;
assign v_18164 = v_4131 & v_4576;
assign v_18166 = v_4100 & v_18165;
assign v_18167 = v_4132 & v_4444;
assign v_18169 = v_3817 & v_18168;
assign v_18170 = v_3843 & v_4294;
assign v_18172 = v_3818 & v_18171;
assign v_18173 = v_3844 & v_4162;
assign v_18175 = v_3527 & v_18174;
assign v_18176 = v_3555 & v_3998;
assign v_18178 = v_3528 & v_18177;
assign v_18179 = v_3556 & v_3866;
assign v_18181 = v_3246 & v_18180;
assign v_18182 = v_3271 & v_3714;
assign v_18184 = v_3247 & v_18183;
assign v_18185 = v_3272 & v_3582;
assign v_18187 = v_2941 & v_18186;
assign v_18188 = v_2977 & v_3426;
assign v_18190 = v_2942 & v_18189;
assign v_18191 = v_2978 & v_3294;
assign v_18193 = v_2658 & v_18192;
assign v_18194 = v_2685 & v_3144;
assign v_18196 = v_2659 & v_18195;
assign v_18197 = v_2686 & v_3012;
assign v_18199 = v_2367 & v_18198;
assign v_18200 = v_2395 & v_2840;
assign v_18202 = v_2368 & v_18201;
assign v_18203 = v_2396 & v_2708;
assign v_18205 = v_2086 & v_18204;
assign v_18206 = v_2111 & v_2554;
assign v_18208 = v_2087 & v_18207;
assign v_18209 = v_2112 & v_2422;
assign v_18211 = v_1789 & v_18210;
assign v_18212 = v_1821 & v_2266;
assign v_18214 = v_1790 & v_18213;
assign v_18215 = v_1822 & v_2134;
assign v_18217 = v_1507 & v_18216;
assign v_18218 = v_1533 & v_1984;
assign v_18220 = v_1508 & v_18219;
assign v_18221 = v_1534 & v_1852;
assign v_18223 = v_1217 & v_18222;
assign v_18224 = v_1245 & v_1688;
assign v_18226 = v_1218 & v_18225;
assign v_18227 = v_1246 & v_1556;
assign v_18229 = v_936 & v_18228;
assign v_18230 = v_961 & v_1404;
assign v_18232 = v_937 & v_18231;
assign v_18233 = v_962 & v_1272;
assign v_18235 = v_92 & v_18234;
assign v_18236 = v_591 & v_1116;
assign v_18238 = v_94 & v_18237;
assign v_18239 = v_593 & v_984;
assign v_18241 = v_806 & v_18240;
assign v_18242 = v_823 & v_838;
assign v_18244 = v_9308 & v_9753;
assign v_18245 = v_9336 & v_9604;
assign v_18247 = v_9026 & v_18246;
assign v_18248 = v_9051 & v_9463;
assign v_18250 = v_9027 & v_18249;
assign v_18251 = v_9052 & v_9311;
assign v_18253 = v_8729 & v_18252;
assign v_18254 = v_8761 & v_9175;
assign v_18256 = v_8730 & v_18255;
assign v_18257 = v_8762 & v_9030;
assign v_18259 = v_8447 & v_18258;
assign v_18260 = v_8473 & v_8893;
assign v_18262 = v_8448 & v_18261;
assign v_18263 = v_8474 & v_8733;
assign v_18265 = v_8157 & v_18264;
assign v_18266 = v_8185 & v_8597;
assign v_18268 = v_8158 & v_18267;
assign v_18269 = v_8186 & v_8451;
assign v_18271 = v_7876 & v_18270;
assign v_18272 = v_7901 & v_8313;
assign v_18274 = v_7877 & v_18273;
assign v_18275 = v_7902 & v_8161;
assign v_18277 = v_7571 & v_18276;
assign v_18278 = v_7607 & v_8025;
assign v_18280 = v_7572 & v_18279;
assign v_18281 = v_7608 & v_7880;
assign v_18283 = v_7288 & v_18282;
assign v_18284 = v_7315 & v_7743;
assign v_18286 = v_7289 & v_18285;
assign v_18287 = v_7316 & v_7575;
assign v_18289 = v_6997 & v_18288;
assign v_18290 = v_7025 & v_7439;
assign v_18292 = v_6998 & v_18291;
assign v_18293 = v_7026 & v_7292;
assign v_18295 = v_6716 & v_18294;
assign v_18296 = v_6741 & v_7153;
assign v_18298 = v_6717 & v_18297;
assign v_18299 = v_6742 & v_7001;
assign v_18301 = v_6419 & v_18300;
assign v_18302 = v_6451 & v_6865;
assign v_18304 = v_6420 & v_18303;
assign v_18305 = v_6452 & v_6720;
assign v_18307 = v_6137 & v_18306;
assign v_18308 = v_6163 & v_6583;
assign v_18310 = v_6138 & v_18309;
assign v_18311 = v_6164 & v_6423;
assign v_18313 = v_5847 & v_18312;
assign v_18314 = v_5875 & v_6287;
assign v_18316 = v_5848 & v_18315;
assign v_18317 = v_5876 & v_6141;
assign v_18319 = v_5566 & v_18318;
assign v_18320 = v_5591 & v_6003;
assign v_18322 = v_5567 & v_18321;
assign v_18323 = v_5592 & v_5851;
assign v_18325 = v_5253 & v_18324;
assign v_18326 = v_5293 & v_5715;
assign v_18328 = v_5254 & v_18327;
assign v_18329 = v_5294 & v_5570;
assign v_18331 = v_4969 & v_18330;
assign v_18332 = v_4997 & v_5433;
assign v_18334 = v_4970 & v_18333;
assign v_18335 = v_4998 & v_5257;
assign v_18337 = v_4677 & v_18336;
assign v_18338 = v_4705 & v_5121;
assign v_18340 = v_4678 & v_18339;
assign v_18341 = v_4706 & v_4973;
assign v_18343 = v_4396 & v_18342;
assign v_18344 = v_4421 & v_4833;
assign v_18346 = v_4397 & v_18345;
assign v_18347 = v_4422 & v_4681;
assign v_18349 = v_4099 & v_18348;
assign v_18350 = v_4131 & v_4545;
assign v_18352 = v_4100 & v_18351;
assign v_18353 = v_4132 & v_4400;
assign v_18355 = v_3817 & v_18354;
assign v_18356 = v_3843 & v_4263;
assign v_18358 = v_3818 & v_18357;
assign v_18359 = v_3844 & v_4103;
assign v_18361 = v_3527 & v_18360;
assign v_18362 = v_3555 & v_3967;
assign v_18364 = v_3528 & v_18363;
assign v_18365 = v_3556 & v_3821;
assign v_18367 = v_3246 & v_18366;
assign v_18368 = v_3271 & v_3683;
assign v_18370 = v_3247 & v_18369;
assign v_18371 = v_3272 & v_3531;
assign v_18373 = v_2941 & v_18372;
assign v_18374 = v_2977 & v_3395;
assign v_18376 = v_2942 & v_18375;
assign v_18377 = v_2978 & v_3250;
assign v_18379 = v_2658 & v_18378;
assign v_18380 = v_2685 & v_3113;
assign v_18382 = v_2659 & v_18381;
assign v_18383 = v_2686 & v_2945;
assign v_18385 = v_2367 & v_18384;
assign v_18386 = v_2395 & v_2809;
assign v_18388 = v_2368 & v_18387;
assign v_18389 = v_2396 & v_2662;
assign v_18391 = v_2086 & v_18390;
assign v_18392 = v_2111 & v_2523;
assign v_18394 = v_2087 & v_18393;
assign v_18395 = v_2112 & v_2371;
assign v_18397 = v_1789 & v_18396;
assign v_18398 = v_1821 & v_2235;
assign v_18400 = v_1790 & v_18399;
assign v_18401 = v_1822 & v_2090;
assign v_18403 = v_1507 & v_18402;
assign v_18404 = v_1533 & v_1953;
assign v_18406 = v_1508 & v_18405;
assign v_18407 = v_1534 & v_1793;
assign v_18409 = v_1217 & v_18408;
assign v_18410 = v_1245 & v_1657;
assign v_18412 = v_1218 & v_18411;
assign v_18413 = v_1246 & v_1511;
assign v_18415 = v_936 & v_18414;
assign v_18416 = v_961 & v_1373;
assign v_18418 = v_937 & v_18417;
assign v_18419 = v_962 & v_1221;
assign v_18421 = v_92 & v_18420;
assign v_18422 = v_591 & v_1085;
assign v_18424 = v_94 & v_18423;
assign v_18425 = v_593 & v_940;
assign v_18427 = v_806 & v_18426;
assign v_18428 = v_804 & v_823;
assign v_18431 = v_9308 & v_9796;
assign v_18432 = v_9336 & v_9664;
assign v_18434 = v_9026 & v_18433;
assign v_18435 = v_9051 & v_9506;
assign v_18437 = v_9027 & v_18436;
assign v_18438 = v_9052 & v_9374;
assign v_18440 = v_8729 & v_18439;
assign v_18441 = v_8761 & v_9218;
assign v_18443 = v_8730 & v_18442;
assign v_18444 = v_8762 & v_9086;
assign v_18446 = v_8447 & v_18445;
assign v_18447 = v_8473 & v_8936;
assign v_18449 = v_8448 & v_18448;
assign v_18450 = v_8474 & v_8804;
assign v_18452 = v_8157 & v_18451;
assign v_18453 = v_8185 & v_8640;
assign v_18455 = v_8158 & v_18454;
assign v_18456 = v_8186 & v_8508;
assign v_18458 = v_7876 & v_18457;
assign v_18459 = v_7901 & v_8356;
assign v_18461 = v_7877 & v_18460;
assign v_18462 = v_7902 & v_8224;
assign v_18464 = v_7571 & v_18463;
assign v_18465 = v_7607 & v_8068;
assign v_18467 = v_7572 & v_18466;
assign v_18468 = v_7608 & v_7936;
assign v_18470 = v_7288 & v_18469;
assign v_18471 = v_7315 & v_7786;
assign v_18473 = v_7289 & v_18472;
assign v_18474 = v_7316 & v_7654;
assign v_18476 = v_6997 & v_18475;
assign v_18477 = v_7025 & v_7482;
assign v_18479 = v_6998 & v_18478;
assign v_18480 = v_7026 & v_7350;
assign v_18482 = v_6716 & v_18481;
assign v_18483 = v_6741 & v_7196;
assign v_18485 = v_6717 & v_18484;
assign v_18486 = v_6742 & v_7064;
assign v_18488 = v_6419 & v_18487;
assign v_18489 = v_6451 & v_6908;
assign v_18491 = v_6420 & v_18490;
assign v_18492 = v_6452 & v_6776;
assign v_18494 = v_6137 & v_18493;
assign v_18495 = v_6163 & v_6626;
assign v_18497 = v_6138 & v_18496;
assign v_18498 = v_6164 & v_6494;
assign v_18500 = v_5847 & v_18499;
assign v_18501 = v_5875 & v_6330;
assign v_18503 = v_5848 & v_18502;
assign v_18504 = v_5876 & v_6198;
assign v_18506 = v_5566 & v_18505;
assign v_18507 = v_5591 & v_6046;
assign v_18509 = v_5567 & v_18508;
assign v_18510 = v_5592 & v_5914;
assign v_18512 = v_5253 & v_18511;
assign v_18513 = v_5293 & v_5758;
assign v_18515 = v_5254 & v_18514;
assign v_18516 = v_5294 & v_5626;
assign v_18518 = v_4969 & v_18517;
assign v_18519 = v_4997 & v_5476;
assign v_18521 = v_4970 & v_18520;
assign v_18522 = v_4998 & v_5344;
assign v_18524 = v_4677 & v_18523;
assign v_18525 = v_4705 & v_5164;
assign v_18527 = v_4678 & v_18526;
assign v_18528 = v_4706 & v_5032;
assign v_18530 = v_4396 & v_18529;
assign v_18531 = v_4421 & v_4876;
assign v_18533 = v_4397 & v_18532;
assign v_18534 = v_4422 & v_4744;
assign v_18536 = v_4099 & v_18535;
assign v_18537 = v_4131 & v_4588;
assign v_18539 = v_4100 & v_18538;
assign v_18540 = v_4132 & v_4456;
assign v_18542 = v_3817 & v_18541;
assign v_18543 = v_3843 & v_4306;
assign v_18545 = v_3818 & v_18544;
assign v_18546 = v_3844 & v_4174;
assign v_18548 = v_3527 & v_18547;
assign v_18549 = v_3555 & v_4010;
assign v_18551 = v_3528 & v_18550;
assign v_18552 = v_3556 & v_3878;
assign v_18554 = v_3246 & v_18553;
assign v_18555 = v_3271 & v_3726;
assign v_18557 = v_3247 & v_18556;
assign v_18558 = v_3272 & v_3594;
assign v_18560 = v_2941 & v_18559;
assign v_18561 = v_2977 & v_3438;
assign v_18563 = v_2942 & v_18562;
assign v_18564 = v_2978 & v_3306;
assign v_18566 = v_2658 & v_18565;
assign v_18567 = v_2685 & v_3156;
assign v_18569 = v_2659 & v_18568;
assign v_18570 = v_2686 & v_3024;
assign v_18572 = v_2367 & v_18571;
assign v_18573 = v_2395 & v_2852;
assign v_18575 = v_2368 & v_18574;
assign v_18576 = v_2396 & v_2720;
assign v_18578 = v_2086 & v_18577;
assign v_18579 = v_2111 & v_2566;
assign v_18581 = v_2087 & v_18580;
assign v_18582 = v_2112 & v_2434;
assign v_18584 = v_1789 & v_18583;
assign v_18585 = v_1821 & v_2278;
assign v_18587 = v_1790 & v_18586;
assign v_18588 = v_1822 & v_2146;
assign v_18590 = v_1507 & v_18589;
assign v_18591 = v_1533 & v_1996;
assign v_18593 = v_1508 & v_18592;
assign v_18594 = v_1534 & v_1864;
assign v_18596 = v_1217 & v_18595;
assign v_18597 = v_1245 & v_1700;
assign v_18599 = v_1218 & v_18598;
assign v_18600 = v_1246 & v_1568;
assign v_18602 = v_936 & v_18601;
assign v_18603 = v_961 & v_1416;
assign v_18605 = v_937 & v_18604;
assign v_18606 = v_962 & v_1284;
assign v_18608 = v_92 & v_18607;
assign v_18609 = v_591 & v_1128;
assign v_18611 = v_94 & v_18610;
assign v_18612 = v_593 & v_996;
assign v_18614 = v_806 & v_18613;
assign v_18615 = v_823 & v_850;
assign v_18618 = v_9308 & v_9808;
assign v_18619 = v_9336 & v_9676;
assign v_18621 = v_9026 & v_18620;
assign v_18622 = v_9051 & v_9518;
assign v_18624 = v_9027 & v_18623;
assign v_18625 = v_9052 & v_9386;
assign v_18627 = v_8729 & v_18626;
assign v_18628 = v_8761 & v_9230;
assign v_18630 = v_8730 & v_18629;
assign v_18631 = v_8762 & v_9098;
assign v_18633 = v_8447 & v_18632;
assign v_18634 = v_8473 & v_8948;
assign v_18636 = v_8448 & v_18635;
assign v_18637 = v_8474 & v_8816;
assign v_18639 = v_8157 & v_18638;
assign v_18640 = v_8185 & v_8652;
assign v_18642 = v_8158 & v_18641;
assign v_18643 = v_8186 & v_8520;
assign v_18645 = v_7876 & v_18644;
assign v_18646 = v_7901 & v_8368;
assign v_18648 = v_7877 & v_18647;
assign v_18649 = v_7902 & v_8236;
assign v_18651 = v_7571 & v_18650;
assign v_18652 = v_7607 & v_8080;
assign v_18654 = v_7572 & v_18653;
assign v_18655 = v_7608 & v_7948;
assign v_18657 = v_7288 & v_18656;
assign v_18658 = v_7315 & v_7798;
assign v_18660 = v_7289 & v_18659;
assign v_18661 = v_7316 & v_7666;
assign v_18663 = v_6997 & v_18662;
assign v_18664 = v_7025 & v_7494;
assign v_18666 = v_6998 & v_18665;
assign v_18667 = v_7026 & v_7362;
assign v_18669 = v_6716 & v_18668;
assign v_18670 = v_6741 & v_7208;
assign v_18672 = v_6717 & v_18671;
assign v_18673 = v_6742 & v_7076;
assign v_18675 = v_6419 & v_18674;
assign v_18676 = v_6451 & v_6920;
assign v_18678 = v_6420 & v_18677;
assign v_18679 = v_6452 & v_6788;
assign v_18681 = v_6137 & v_18680;
assign v_18682 = v_6163 & v_6638;
assign v_18684 = v_6138 & v_18683;
assign v_18685 = v_6164 & v_6506;
assign v_18687 = v_5847 & v_18686;
assign v_18688 = v_5875 & v_6342;
assign v_18690 = v_5848 & v_18689;
assign v_18691 = v_5876 & v_6210;
assign v_18693 = v_5566 & v_18692;
assign v_18694 = v_5591 & v_6058;
assign v_18696 = v_5567 & v_18695;
assign v_18697 = v_5592 & v_5926;
assign v_18699 = v_5253 & v_18698;
assign v_18700 = v_5293 & v_5770;
assign v_18702 = v_5254 & v_18701;
assign v_18703 = v_5294 & v_5638;
assign v_18705 = v_4969 & v_18704;
assign v_18706 = v_4997 & v_5488;
assign v_18708 = v_4970 & v_18707;
assign v_18709 = v_4998 & v_5356;
assign v_18711 = v_4677 & v_18710;
assign v_18712 = v_4705 & v_5176;
assign v_18714 = v_4678 & v_18713;
assign v_18715 = v_4706 & v_5044;
assign v_18717 = v_4396 & v_18716;
assign v_18718 = v_4421 & v_4888;
assign v_18720 = v_4397 & v_18719;
assign v_18721 = v_4422 & v_4756;
assign v_18723 = v_4099 & v_18722;
assign v_18724 = v_4131 & v_4600;
assign v_18726 = v_4100 & v_18725;
assign v_18727 = v_4132 & v_4468;
assign v_18729 = v_3817 & v_18728;
assign v_18730 = v_3843 & v_4318;
assign v_18732 = v_3818 & v_18731;
assign v_18733 = v_3844 & v_4186;
assign v_18735 = v_3527 & v_18734;
assign v_18736 = v_3555 & v_4022;
assign v_18738 = v_3528 & v_18737;
assign v_18739 = v_3556 & v_3890;
assign v_18741 = v_3246 & v_18740;
assign v_18742 = v_3271 & v_3738;
assign v_18744 = v_3247 & v_18743;
assign v_18745 = v_3272 & v_3606;
assign v_18747 = v_2941 & v_18746;
assign v_18748 = v_2977 & v_3450;
assign v_18750 = v_2942 & v_18749;
assign v_18751 = v_2978 & v_3318;
assign v_18753 = v_2658 & v_18752;
assign v_18754 = v_2685 & v_3168;
assign v_18756 = v_2659 & v_18755;
assign v_18757 = v_2686 & v_3036;
assign v_18759 = v_2367 & v_18758;
assign v_18760 = v_2395 & v_2864;
assign v_18762 = v_2368 & v_18761;
assign v_18763 = v_2396 & v_2732;
assign v_18765 = v_2086 & v_18764;
assign v_18766 = v_2111 & v_2578;
assign v_18768 = v_2087 & v_18767;
assign v_18769 = v_2112 & v_2446;
assign v_18771 = v_1789 & v_18770;
assign v_18772 = v_1821 & v_2290;
assign v_18774 = v_1790 & v_18773;
assign v_18775 = v_1822 & v_2158;
assign v_18777 = v_1507 & v_18776;
assign v_18778 = v_1533 & v_2008;
assign v_18780 = v_1508 & v_18779;
assign v_18781 = v_1534 & v_1876;
assign v_18783 = v_1217 & v_18782;
assign v_18784 = v_1245 & v_1712;
assign v_18786 = v_1218 & v_18785;
assign v_18787 = v_1246 & v_1580;
assign v_18789 = v_936 & v_18788;
assign v_18790 = v_961 & v_1428;
assign v_18792 = v_937 & v_18791;
assign v_18793 = v_962 & v_1296;
assign v_18795 = v_92 & v_18794;
assign v_18796 = v_591 & v_1140;
assign v_18798 = v_94 & v_18797;
assign v_18799 = v_593 & v_1008;
assign v_18801 = v_806 & v_18800;
assign v_18802 = v_823 & v_862;
assign v_18805 = v_9308 & v_9820;
assign v_18806 = v_9336 & v_9688;
assign v_18808 = v_9026 & v_18807;
assign v_18809 = v_9051 & v_9530;
assign v_18811 = v_9027 & v_18810;
assign v_18812 = v_9052 & v_9398;
assign v_18814 = v_8729 & v_18813;
assign v_18815 = v_8761 & v_9242;
assign v_18817 = v_8730 & v_18816;
assign v_18818 = v_8762 & v_9110;
assign v_18820 = v_8447 & v_18819;
assign v_18821 = v_8473 & v_8960;
assign v_18823 = v_8448 & v_18822;
assign v_18824 = v_8474 & v_8828;
assign v_18826 = v_8157 & v_18825;
assign v_18827 = v_8185 & v_8664;
assign v_18829 = v_8158 & v_18828;
assign v_18830 = v_8186 & v_8532;
assign v_18832 = v_7876 & v_18831;
assign v_18833 = v_7901 & v_8380;
assign v_18835 = v_7877 & v_18834;
assign v_18836 = v_7902 & v_8248;
assign v_18838 = v_7571 & v_18837;
assign v_18839 = v_7607 & v_8092;
assign v_18841 = v_7572 & v_18840;
assign v_18842 = v_7608 & v_7960;
assign v_18844 = v_7288 & v_18843;
assign v_18845 = v_7315 & v_7810;
assign v_18847 = v_7289 & v_18846;
assign v_18848 = v_7316 & v_7678;
assign v_18850 = v_6997 & v_18849;
assign v_18851 = v_7025 & v_7506;
assign v_18853 = v_6998 & v_18852;
assign v_18854 = v_7026 & v_7374;
assign v_18856 = v_6716 & v_18855;
assign v_18857 = v_6741 & v_7220;
assign v_18859 = v_6717 & v_18858;
assign v_18860 = v_6742 & v_7088;
assign v_18862 = v_6419 & v_18861;
assign v_18863 = v_6451 & v_6932;
assign v_18865 = v_6420 & v_18864;
assign v_18866 = v_6452 & v_6800;
assign v_18868 = v_6137 & v_18867;
assign v_18869 = v_6163 & v_6650;
assign v_18871 = v_6138 & v_18870;
assign v_18872 = v_6164 & v_6518;
assign v_18874 = v_5847 & v_18873;
assign v_18875 = v_5875 & v_6354;
assign v_18877 = v_5848 & v_18876;
assign v_18878 = v_5876 & v_6222;
assign v_18880 = v_5566 & v_18879;
assign v_18881 = v_5591 & v_6070;
assign v_18883 = v_5567 & v_18882;
assign v_18884 = v_5592 & v_5938;
assign v_18886 = v_5253 & v_18885;
assign v_18887 = v_5293 & v_5782;
assign v_18889 = v_5254 & v_18888;
assign v_18890 = v_5294 & v_5650;
assign v_18892 = v_4969 & v_18891;
assign v_18893 = v_4997 & v_5500;
assign v_18895 = v_4970 & v_18894;
assign v_18896 = v_4998 & v_5368;
assign v_18898 = v_4677 & v_18897;
assign v_18899 = v_4705 & v_5188;
assign v_18901 = v_4678 & v_18900;
assign v_18902 = v_4706 & v_5056;
assign v_18904 = v_4396 & v_18903;
assign v_18905 = v_4421 & v_4900;
assign v_18907 = v_4397 & v_18906;
assign v_18908 = v_4422 & v_4768;
assign v_18910 = v_4099 & v_18909;
assign v_18911 = v_4131 & v_4612;
assign v_18913 = v_4100 & v_18912;
assign v_18914 = v_4132 & v_4480;
assign v_18916 = v_3817 & v_18915;
assign v_18917 = v_3843 & v_4330;
assign v_18919 = v_3818 & v_18918;
assign v_18920 = v_3844 & v_4198;
assign v_18922 = v_3527 & v_18921;
assign v_18923 = v_3555 & v_4034;
assign v_18925 = v_3528 & v_18924;
assign v_18926 = v_3556 & v_3902;
assign v_18928 = v_3246 & v_18927;
assign v_18929 = v_3271 & v_3750;
assign v_18931 = v_3247 & v_18930;
assign v_18932 = v_3272 & v_3618;
assign v_18934 = v_2941 & v_18933;
assign v_18935 = v_2977 & v_3462;
assign v_18937 = v_2942 & v_18936;
assign v_18938 = v_2978 & v_3330;
assign v_18940 = v_2658 & v_18939;
assign v_18941 = v_2685 & v_3180;
assign v_18943 = v_2659 & v_18942;
assign v_18944 = v_2686 & v_3048;
assign v_18946 = v_2367 & v_18945;
assign v_18947 = v_2395 & v_2876;
assign v_18949 = v_2368 & v_18948;
assign v_18950 = v_2396 & v_2744;
assign v_18952 = v_2086 & v_18951;
assign v_18953 = v_2111 & v_2590;
assign v_18955 = v_2087 & v_18954;
assign v_18956 = v_2112 & v_2458;
assign v_18958 = v_1789 & v_18957;
assign v_18959 = v_1821 & v_2302;
assign v_18961 = v_1790 & v_18960;
assign v_18962 = v_1822 & v_2170;
assign v_18964 = v_1507 & v_18963;
assign v_18965 = v_1533 & v_2020;
assign v_18967 = v_1508 & v_18966;
assign v_18968 = v_1534 & v_1888;
assign v_18970 = v_1217 & v_18969;
assign v_18971 = v_1245 & v_1724;
assign v_18973 = v_1218 & v_18972;
assign v_18974 = v_1246 & v_1592;
assign v_18976 = v_936 & v_18975;
assign v_18977 = v_961 & v_1440;
assign v_18979 = v_937 & v_18978;
assign v_18980 = v_962 & v_1308;
assign v_18982 = v_92 & v_18981;
assign v_18983 = v_591 & v_1152;
assign v_18985 = v_94 & v_18984;
assign v_18986 = v_593 & v_1020;
assign v_18988 = v_806 & v_18987;
assign v_18989 = v_823 & v_874;
assign v_18992 = v_9308 & v_9832;
assign v_18993 = v_9336 & v_9700;
assign v_18995 = v_9026 & v_18994;
assign v_18996 = v_9051 & v_9542;
assign v_18998 = v_9027 & v_18997;
assign v_18999 = v_9052 & v_9410;
assign v_19001 = v_8729 & v_19000;
assign v_19002 = v_8761 & v_9254;
assign v_19004 = v_8730 & v_19003;
assign v_19005 = v_8762 & v_9122;
assign v_19007 = v_8447 & v_19006;
assign v_19008 = v_8473 & v_8972;
assign v_19010 = v_8448 & v_19009;
assign v_19011 = v_8474 & v_8840;
assign v_19013 = v_8157 & v_19012;
assign v_19014 = v_8185 & v_8676;
assign v_19016 = v_8158 & v_19015;
assign v_19017 = v_8186 & v_8544;
assign v_19019 = v_7876 & v_19018;
assign v_19020 = v_7901 & v_8392;
assign v_19022 = v_7877 & v_19021;
assign v_19023 = v_7902 & v_8260;
assign v_19025 = v_7571 & v_19024;
assign v_19026 = v_7607 & v_8104;
assign v_19028 = v_7572 & v_19027;
assign v_19029 = v_7608 & v_7972;
assign v_19031 = v_7288 & v_19030;
assign v_19032 = v_7315 & v_7822;
assign v_19034 = v_7289 & v_19033;
assign v_19035 = v_7316 & v_7690;
assign v_19037 = v_6997 & v_19036;
assign v_19038 = v_7025 & v_7518;
assign v_19040 = v_6998 & v_19039;
assign v_19041 = v_7026 & v_7386;
assign v_19043 = v_6716 & v_19042;
assign v_19044 = v_6741 & v_7232;
assign v_19046 = v_6717 & v_19045;
assign v_19047 = v_6742 & v_7100;
assign v_19049 = v_6419 & v_19048;
assign v_19050 = v_6451 & v_6944;
assign v_19052 = v_6420 & v_19051;
assign v_19053 = v_6452 & v_6812;
assign v_19055 = v_6137 & v_19054;
assign v_19056 = v_6163 & v_6662;
assign v_19058 = v_6138 & v_19057;
assign v_19059 = v_6164 & v_6530;
assign v_19061 = v_5847 & v_19060;
assign v_19062 = v_5875 & v_6366;
assign v_19064 = v_5848 & v_19063;
assign v_19065 = v_5876 & v_6234;
assign v_19067 = v_5566 & v_19066;
assign v_19068 = v_5591 & v_6082;
assign v_19070 = v_5567 & v_19069;
assign v_19071 = v_5592 & v_5950;
assign v_19073 = v_5253 & v_19072;
assign v_19074 = v_5293 & v_5794;
assign v_19076 = v_5254 & v_19075;
assign v_19077 = v_5294 & v_5662;
assign v_19079 = v_4969 & v_19078;
assign v_19080 = v_4997 & v_5512;
assign v_19082 = v_4970 & v_19081;
assign v_19083 = v_4998 & v_5380;
assign v_19085 = v_4677 & v_19084;
assign v_19086 = v_4705 & v_5200;
assign v_19088 = v_4678 & v_19087;
assign v_19089 = v_4706 & v_5068;
assign v_19091 = v_4396 & v_19090;
assign v_19092 = v_4421 & v_4912;
assign v_19094 = v_4397 & v_19093;
assign v_19095 = v_4422 & v_4780;
assign v_19097 = v_4099 & v_19096;
assign v_19098 = v_4131 & v_4624;
assign v_19100 = v_4100 & v_19099;
assign v_19101 = v_4132 & v_4492;
assign v_19103 = v_3817 & v_19102;
assign v_19104 = v_3843 & v_4342;
assign v_19106 = v_3818 & v_19105;
assign v_19107 = v_3844 & v_4210;
assign v_19109 = v_3527 & v_19108;
assign v_19110 = v_3555 & v_4046;
assign v_19112 = v_3528 & v_19111;
assign v_19113 = v_3556 & v_3914;
assign v_19115 = v_3246 & v_19114;
assign v_19116 = v_3271 & v_3762;
assign v_19118 = v_3247 & v_19117;
assign v_19119 = v_3272 & v_3630;
assign v_19121 = v_2941 & v_19120;
assign v_19122 = v_2977 & v_3474;
assign v_19124 = v_2942 & v_19123;
assign v_19125 = v_2978 & v_3342;
assign v_19127 = v_2658 & v_19126;
assign v_19128 = v_2685 & v_3192;
assign v_19130 = v_2659 & v_19129;
assign v_19131 = v_2686 & v_3060;
assign v_19133 = v_2367 & v_19132;
assign v_19134 = v_2395 & v_2888;
assign v_19136 = v_2368 & v_19135;
assign v_19137 = v_2396 & v_2756;
assign v_19139 = v_2086 & v_19138;
assign v_19140 = v_2111 & v_2602;
assign v_19142 = v_2087 & v_19141;
assign v_19143 = v_2112 & v_2470;
assign v_19145 = v_1789 & v_19144;
assign v_19146 = v_1821 & v_2314;
assign v_19148 = v_1790 & v_19147;
assign v_19149 = v_1822 & v_2182;
assign v_19151 = v_1507 & v_19150;
assign v_19152 = v_1533 & v_2032;
assign v_19154 = v_1508 & v_19153;
assign v_19155 = v_1534 & v_1900;
assign v_19157 = v_1217 & v_19156;
assign v_19158 = v_1245 & v_1736;
assign v_19160 = v_1218 & v_19159;
assign v_19161 = v_1246 & v_1604;
assign v_19163 = v_936 & v_19162;
assign v_19164 = v_961 & v_1452;
assign v_19166 = v_937 & v_19165;
assign v_19167 = v_962 & v_1320;
assign v_19169 = v_92 & v_19168;
assign v_19170 = v_591 & v_1164;
assign v_19172 = v_94 & v_19171;
assign v_19173 = v_593 & v_1032;
assign v_19175 = v_806 & v_19174;
assign v_19176 = v_823 & v_886;
assign v_19181 = v_19179 & v_19180;
assign v_19184 = v_19182 & v_19183;
assign v_19187 = v_19185 & v_19186;
assign v_19190 = v_19188 & v_19189;
assign v_19193 = v_19191 & v_19192;
assign v_19196 = v_19194 & v_19195;
assign v_19199 = v_19197 & v_19198;
assign v_19202 = v_19200 & v_19201;
assign v_19205 = v_19203 & v_19204;
assign v_19208 = v_19206 & v_19207;
assign v_19211 = v_19209 & v_19210;
assign v_19214 = v_19212 & v_19213;
assign v_19217 = v_19215 & v_19216;
assign v_19220 = v_19218 & v_19219;
assign v_19223 = v_19221 & v_19222;
assign v_19226 = v_19224 & v_19225;
assign v_19229 = v_19227 & v_19228;
assign v_19232 = v_19230 & v_19231;
assign v_19235 = v_19233 & v_19234;
assign v_19238 = v_19236 & v_19237;
assign v_19241 = v_19239 & v_19240;
assign v_19244 = v_19242 & v_19243;
assign v_19247 = v_19245 & v_19246;
assign v_19250 = v_19248 & v_19249;
assign v_19253 = v_19251 & v_19252;
assign v_19256 = v_19254 & v_19255;
assign v_19259 = v_19257 & v_19258;
assign v_19262 = v_19260 & v_19261;
assign v_19265 = v_19263 & v_19264;
assign v_19268 = v_19266 & v_19267;
assign v_19271 = v_19269 & v_19270;
assign v_19274 = v_19272 & v_19273;
assign v_19277 = v_19275 & v_19276;
assign v_19280 = v_19278 & v_19279;
assign v_19283 = v_19281 & v_19282;
assign v_19286 = v_19284 & v_19285;
assign v_19289 = v_19287 & v_19288;
assign v_19292 = v_19290 & v_19291;
assign v_19295 = v_19293 & v_19294;
assign v_19298 = v_19296 & v_19297;
assign v_19301 = v_19299 & v_19300;
assign v_19304 = v_19302 & v_19303;
assign v_19307 = v_19305 & v_19306;
assign v_19310 = v_19308 & v_19309;
assign v_19313 = v_19311 & v_19312;
assign v_19316 = v_19314 & v_19315;
assign v_19319 = v_19317 & v_19318;
assign v_19322 = v_19320 & v_19321;
assign v_19325 = v_19323 & v_19324;
assign v_19328 = v_19326 & v_19327;
assign v_19331 = v_19329 & v_19330;
assign v_19334 = v_19332 & v_19333;
assign v_19337 = v_19335 & v_19336;
assign v_19340 = v_19338 & v_19339;
assign v_19343 = v_19341 & v_19342;
assign v_19346 = v_19344 & v_19345;
assign v_19349 = v_19347 & v_19348;
assign v_19352 = v_19350 & v_19351;
assign v_19355 = v_19353 & v_19354;
assign v_19358 = v_19356 & v_19357;
assign v_19361 = v_19359 & v_19360;
assign v_19364 = v_19362 & v_19363;
assign v_19366 = v_9308 & ~v_9872;
assign v_19367 = v_9336 & ~v_9740;
assign v_19369 = v_9026 & v_19368;
assign v_19370 = v_9051 & ~v_9582;
assign v_19372 = v_9027 & v_19371;
assign v_19373 = v_9052 & ~v_9450;
assign v_19375 = v_8729 & v_19374;
assign v_19376 = v_8761 & ~v_9294;
assign v_19378 = v_8730 & v_19377;
assign v_19379 = v_8762 & ~v_9162;
assign v_19381 = v_8447 & v_19380;
assign v_19382 = v_8473 & ~v_9012;
assign v_19384 = v_8448 & v_19383;
assign v_19385 = v_8474 & ~v_8880;
assign v_19387 = v_8157 & v_19386;
assign v_19388 = v_8185 & ~v_8716;
assign v_19390 = v_8158 & v_19389;
assign v_19391 = v_8186 & ~v_8584;
assign v_19393 = v_7876 & v_19392;
assign v_19394 = v_7901 & v_8432;
assign v_19396 = v_7877 & v_19395;
assign v_19397 = v_7902 & v_8300;
assign v_19399 = v_7571 & v_19398;
assign v_19400 = v_7607 & v_8144;
assign v_19402 = v_7572 & v_19401;
assign v_19403 = v_7608 & ~v_8012;
assign v_19405 = v_7288 & v_19404;
assign v_19406 = v_7315 & ~v_7862;
assign v_19408 = v_7289 & v_19407;
assign v_19409 = v_7316 & ~v_7730;
assign v_19411 = v_6997 & v_19410;
assign v_19412 = v_7025 & ~v_7558;
assign v_19414 = v_6998 & v_19413;
assign v_19415 = v_7026 & ~v_7426;
assign v_19417 = v_6716 & v_19416;
assign v_19418 = v_6741 & v_7272;
assign v_19420 = v_6717 & v_19419;
assign v_19421 = v_6742 & ~v_7140;
assign v_19423 = v_6419 & v_19422;
assign v_19424 = v_6451 & v_6984;
assign v_19426 = v_6420 & v_19425;
assign v_19427 = v_6452 & v_6852;
assign v_19429 = v_6137 & v_19428;
assign v_19430 = v_6163 & v_6702;
assign v_19432 = v_6138 & v_19431;
assign v_19433 = v_6164 & ~v_6570;
assign v_19435 = v_5847 & v_19434;
assign v_19436 = v_5875 & ~v_6406;
assign v_19438 = v_5848 & v_19437;
assign v_19439 = v_5876 & v_6274;
assign v_19441 = v_5566 & v_19440;
assign v_19442 = v_5591 & v_6122;
assign v_19444 = v_5567 & v_19443;
assign v_19445 = v_5592 & v_5990;
assign v_19447 = v_5253 & v_19446;
assign v_19448 = v_5293 & v_5834;
assign v_19450 = v_5254 & v_19449;
assign v_19451 = v_5294 & v_5702;
assign v_19453 = v_4969 & v_19452;
assign v_19454 = v_4997 & v_5552;
assign v_19456 = v_4970 & v_19455;
assign v_19457 = v_4998 & ~v_5420;
assign v_19459 = v_4677 & v_19458;
assign v_19460 = v_4705 & ~v_5240;
assign v_19462 = v_4678 & v_19461;
assign v_19463 = v_4706 & v_5108;
assign v_19465 = v_4396 & v_19464;
assign v_19466 = v_4421 & v_4952;
assign v_19468 = v_4397 & v_19467;
assign v_19469 = v_4422 & v_4820;
assign v_19471 = v_4099 & v_19470;
assign v_19472 = v_4131 & v_4664;
assign v_19474 = v_4100 & v_19473;
assign v_19475 = v_4132 & v_4532;
assign v_19477 = v_3817 & v_19476;
assign v_19478 = v_3843 & v_4382;
assign v_19480 = v_3818 & v_19479;
assign v_19481 = v_3844 & ~v_4250;
assign v_19483 = v_3527 & v_19482;
assign v_19484 = v_3555 & ~v_4086;
assign v_19486 = v_3528 & v_19485;
assign v_19487 = v_3556 & ~v_3954;
assign v_19489 = v_3246 & v_19488;
assign v_19490 = v_3271 & ~v_3802;
assign v_19492 = v_3247 & v_19491;
assign v_19493 = v_3272 & ~v_3670;
assign v_19495 = v_2941 & v_19494;
assign v_19496 = v_2977 & v_3514;
assign v_19498 = v_2942 & v_19497;
assign v_19499 = v_2978 & ~v_3382;
assign v_19501 = v_2658 & v_19500;
assign v_19502 = v_2685 & v_3232;
assign v_19504 = v_2659 & v_19503;
assign v_19505 = v_2686 & ~v_3100;
assign v_19507 = v_2367 & v_19506;
assign v_19508 = v_2395 & ~v_2928;
assign v_19510 = v_2368 & v_19509;
assign v_19511 = v_2396 & ~v_2796;
assign v_19513 = v_2086 & v_19512;
assign v_19514 = v_2111 & ~v_2642;
assign v_19516 = v_2087 & v_19515;
assign v_19517 = v_2112 & ~v_2510;
assign v_19519 = v_1789 & v_19518;
assign v_19520 = v_1821 & v_2354;
assign v_19522 = v_1790 & v_19521;
assign v_19523 = v_1822 & v_2222;
assign v_19525 = v_1507 & v_19524;
assign v_19526 = v_1533 & v_2072;
assign v_19528 = v_1508 & v_19527;
assign v_19529 = v_1534 & ~v_1940;
assign v_19531 = v_1217 & v_19530;
assign v_19532 = v_1245 & ~v_1776;
assign v_19534 = v_1218 & v_19533;
assign v_19535 = v_1246 & ~v_1644;
assign v_19537 = v_936 & v_19536;
assign v_19538 = v_961 & ~v_1492;
assign v_19540 = v_937 & v_19539;
assign v_19541 = v_962 & ~v_1360;
assign v_19543 = v_92 & v_19542;
assign v_19544 = v_591 & ~v_1204;
assign v_19546 = v_94 & v_19545;
assign v_19547 = v_593 & ~v_1072;
assign v_19549 = v_806 & v_19548;
assign v_19550 = v_823 & ~v_922;
assign v_19556 = v_807 & v_19555;
assign v_19557 = v_9600 & v_9784;
assign v_19558 = v_9629 & v_9652;
assign v_19560 = v_9601 & v_19559;
assign v_19561 = v_9494 & v_9630;
assign v_19563 = v_9307 & v_19562;
assign v_19564 = v_9335 & v_9362;
assign v_19566 = v_9308 & v_19565;
assign v_19567 = v_9206 & v_9336;
assign v_19569 = v_9026 & v_19568;
assign v_19570 = v_9051 & v_9074;
assign v_19572 = v_9027 & v_19571;
assign v_19573 = v_8924 & v_9052;
assign v_19575 = v_8729 & v_19574;
assign v_19576 = v_8761 & v_8792;
assign v_19578 = v_8730 & v_19577;
assign v_19579 = v_8628 & v_8762;
assign v_19581 = v_8447 & v_19580;
assign v_19582 = v_8473 & v_8496;
assign v_19584 = v_8448 & v_19583;
assign v_19585 = v_8344 & v_8474;
assign v_19587 = v_8157 & v_19586;
assign v_19588 = v_8185 & v_8212;
assign v_19590 = v_8158 & v_19589;
assign v_19591 = v_8056 & v_8186;
assign v_19593 = v_7876 & v_19592;
assign v_19594 = v_7901 & v_7924;
assign v_19596 = v_7877 & v_19595;
assign v_19597 = v_7774 & v_7902;
assign v_19599 = v_7571 & v_19598;
assign v_19600 = v_7607 & v_7642;
assign v_19602 = v_7572 & v_19601;
assign v_19603 = v_7470 & v_7608;
assign v_19605 = v_7288 & v_19604;
assign v_19606 = v_7315 & v_7338;
assign v_19608 = v_7289 & v_19607;
assign v_19609 = v_7184 & v_7316;
assign v_19611 = v_6997 & v_19610;
assign v_19612 = v_7025 & v_7052;
assign v_19614 = v_6998 & v_19613;
assign v_19615 = v_6896 & v_7026;
assign v_19617 = v_6716 & v_19616;
assign v_19618 = v_6741 & v_6764;
assign v_19620 = v_6717 & v_19619;
assign v_19621 = v_6614 & v_6742;
assign v_19623 = v_6419 & v_19622;
assign v_19624 = v_6451 & v_6482;
assign v_19626 = v_6420 & v_19625;
assign v_19627 = v_6318 & v_6452;
assign v_19629 = v_6137 & v_19628;
assign v_19630 = v_6163 & v_6186;
assign v_19632 = v_6138 & v_19631;
assign v_19633 = v_6034 & v_6164;
assign v_19635 = v_5847 & v_19634;
assign v_19636 = v_5875 & v_5902;
assign v_19638 = v_5848 & v_19637;
assign v_19639 = v_5746 & v_5876;
assign v_19641 = v_5566 & v_19640;
assign v_19642 = v_5591 & v_5614;
assign v_19644 = v_5567 & v_19643;
assign v_19645 = v_5464 & v_5592;
assign v_19647 = v_5253 & v_19646;
assign v_19648 = v_5293 & v_5332;
assign v_19650 = v_5254 & v_19649;
assign v_19651 = v_5152 & v_5294;
assign v_19653 = v_4969 & v_19652;
assign v_19654 = v_4997 & v_5020;
assign v_19656 = v_4970 & v_19655;
assign v_19657 = v_4864 & v_4998;
assign v_19659 = v_4677 & v_19658;
assign v_19660 = v_4705 & v_4732;
assign v_19662 = v_4678 & v_19661;
assign v_19663 = v_4576 & v_4706;
assign v_19665 = v_4396 & v_19664;
assign v_19666 = v_4421 & v_4444;
assign v_19668 = v_4397 & v_19667;
assign v_19669 = v_4294 & v_4422;
assign v_19671 = v_4099 & v_19670;
assign v_19672 = v_4131 & v_4162;
assign v_19674 = v_4100 & v_19673;
assign v_19675 = v_3998 & v_4132;
assign v_19677 = v_3817 & v_19676;
assign v_19678 = v_3843 & v_3866;
assign v_19680 = v_3818 & v_19679;
assign v_19681 = v_3714 & v_3844;
assign v_19683 = v_3527 & v_19682;
assign v_19684 = v_3555 & v_3582;
assign v_19686 = v_3528 & v_19685;
assign v_19687 = v_3426 & v_3556;
assign v_19689 = v_3246 & v_19688;
assign v_19690 = v_3271 & v_3294;
assign v_19692 = v_3247 & v_19691;
assign v_19693 = v_3144 & v_3272;
assign v_19695 = v_2941 & v_19694;
assign v_19696 = v_2977 & v_3012;
assign v_19698 = v_2942 & v_19697;
assign v_19699 = v_2840 & v_2978;
assign v_19701 = v_2658 & v_19700;
assign v_19702 = v_2685 & v_2708;
assign v_19704 = v_2659 & v_19703;
assign v_19705 = v_2554 & v_2686;
assign v_19707 = v_2367 & v_19706;
assign v_19708 = v_2395 & v_2422;
assign v_19710 = v_2368 & v_19709;
assign v_19711 = v_2266 & v_2396;
assign v_19713 = v_2086 & v_19712;
assign v_19714 = v_2111 & v_2134;
assign v_19716 = v_2087 & v_19715;
assign v_19717 = v_1984 & v_2112;
assign v_19719 = v_1789 & v_19718;
assign v_19720 = v_1821 & v_1852;
assign v_19722 = v_1790 & v_19721;
assign v_19723 = v_1688 & v_1822;
assign v_19725 = v_1507 & v_19724;
assign v_19726 = v_1533 & v_1556;
assign v_19728 = v_1508 & v_19727;
assign v_19729 = v_1404 & v_1534;
assign v_19731 = v_1217 & v_19730;
assign v_19732 = v_1245 & v_1272;
assign v_19734 = v_1218 & v_19733;
assign v_19735 = v_1116 & v_1246;
assign v_19737 = v_936 & v_19736;
assign v_19738 = v_961 & v_984;
assign v_19740 = v_937 & v_19739;
assign v_19741 = v_838 & v_962;
assign v_19743 = v_92 & v_19742;
assign v_19744 = v_591 & v_721;
assign v_19746 = v_9600 & v_9753;
assign v_19747 = v_9604 & v_9629;
assign v_19749 = v_9601 & v_19748;
assign v_19750 = v_9463 & v_9630;
assign v_19752 = v_9307 & v_19751;
assign v_19753 = v_9311 & v_9335;
assign v_19755 = v_9308 & v_19754;
assign v_19756 = v_9175 & v_9336;
assign v_19758 = v_9026 & v_19757;
assign v_19759 = v_9030 & v_9051;
assign v_19761 = v_9027 & v_19760;
assign v_19762 = v_8893 & v_9052;
assign v_19764 = v_8729 & v_19763;
assign v_19765 = v_8733 & v_8761;
assign v_19767 = v_8730 & v_19766;
assign v_19768 = v_8597 & v_8762;
assign v_19770 = v_8447 & v_19769;
assign v_19771 = v_8451 & v_8473;
assign v_19773 = v_8448 & v_19772;
assign v_19774 = v_8313 & v_8474;
assign v_19776 = v_8157 & v_19775;
assign v_19777 = v_8161 & v_8185;
assign v_19779 = v_8158 & v_19778;
assign v_19780 = v_8025 & v_8186;
assign v_19782 = v_7876 & v_19781;
assign v_19783 = v_7880 & v_7901;
assign v_19785 = v_7877 & v_19784;
assign v_19786 = v_7743 & v_7902;
assign v_19788 = v_7571 & v_19787;
assign v_19789 = v_7575 & v_7607;
assign v_19791 = v_7572 & v_19790;
assign v_19792 = v_7439 & v_7608;
assign v_19794 = v_7288 & v_19793;
assign v_19795 = v_7292 & v_7315;
assign v_19797 = v_7289 & v_19796;
assign v_19798 = v_7153 & v_7316;
assign v_19800 = v_6997 & v_19799;
assign v_19801 = v_7001 & v_7025;
assign v_19803 = v_6998 & v_19802;
assign v_19804 = v_6865 & v_7026;
assign v_19806 = v_6716 & v_19805;
assign v_19807 = v_6720 & v_6741;
assign v_19809 = v_6717 & v_19808;
assign v_19810 = v_6583 & v_6742;
assign v_19812 = v_6419 & v_19811;
assign v_19813 = v_6423 & v_6451;
assign v_19815 = v_6420 & v_19814;
assign v_19816 = v_6287 & v_6452;
assign v_19818 = v_6137 & v_19817;
assign v_19819 = v_6141 & v_6163;
assign v_19821 = v_6138 & v_19820;
assign v_19822 = v_6003 & v_6164;
assign v_19824 = v_5847 & v_19823;
assign v_19825 = v_5851 & v_5875;
assign v_19827 = v_5848 & v_19826;
assign v_19828 = v_5715 & v_5876;
assign v_19830 = v_5566 & v_19829;
assign v_19831 = v_5570 & v_5591;
assign v_19833 = v_5567 & v_19832;
assign v_19834 = v_5433 & v_5592;
assign v_19836 = v_5253 & v_19835;
assign v_19837 = v_5257 & v_5293;
assign v_19839 = v_5254 & v_19838;
assign v_19840 = v_5121 & v_5294;
assign v_19842 = v_4969 & v_19841;
assign v_19843 = v_4973 & v_4997;
assign v_19845 = v_4970 & v_19844;
assign v_19846 = v_4833 & v_4998;
assign v_19848 = v_4677 & v_19847;
assign v_19849 = v_4681 & v_4705;
assign v_19851 = v_4678 & v_19850;
assign v_19852 = v_4545 & v_4706;
assign v_19854 = v_4396 & v_19853;
assign v_19855 = v_4400 & v_4421;
assign v_19857 = v_4397 & v_19856;
assign v_19858 = v_4263 & v_4422;
assign v_19860 = v_4099 & v_19859;
assign v_19861 = v_4103 & v_4131;
assign v_19863 = v_4100 & v_19862;
assign v_19864 = v_3967 & v_4132;
assign v_19866 = v_3817 & v_19865;
assign v_19867 = v_3821 & v_3843;
assign v_19869 = v_3818 & v_19868;
assign v_19870 = v_3683 & v_3844;
assign v_19872 = v_3527 & v_19871;
assign v_19873 = v_3531 & v_3555;
assign v_19875 = v_3528 & v_19874;
assign v_19876 = v_3395 & v_3556;
assign v_19878 = v_3246 & v_19877;
assign v_19879 = v_3250 & v_3271;
assign v_19881 = v_3247 & v_19880;
assign v_19882 = v_3113 & v_3272;
assign v_19884 = v_2941 & v_19883;
assign v_19885 = v_2945 & v_2977;
assign v_19887 = v_2942 & v_19886;
assign v_19888 = v_2809 & v_2978;
assign v_19890 = v_2658 & v_19889;
assign v_19891 = v_2662 & v_2685;
assign v_19893 = v_2659 & v_19892;
assign v_19894 = v_2523 & v_2686;
assign v_19896 = v_2367 & v_19895;
assign v_19897 = v_2371 & v_2395;
assign v_19899 = v_2368 & v_19898;
assign v_19900 = v_2235 & v_2396;
assign v_19902 = v_2086 & v_19901;
assign v_19903 = v_2090 & v_2111;
assign v_19905 = v_2087 & v_19904;
assign v_19906 = v_1953 & v_2112;
assign v_19908 = v_1789 & v_19907;
assign v_19909 = v_1793 & v_1821;
assign v_19911 = v_1790 & v_19910;
assign v_19912 = v_1657 & v_1822;
assign v_19914 = v_1507 & v_19913;
assign v_19915 = v_1511 & v_1533;
assign v_19917 = v_1508 & v_19916;
assign v_19918 = v_1373 & v_1534;
assign v_19920 = v_1217 & v_19919;
assign v_19921 = v_1221 & v_1245;
assign v_19923 = v_1218 & v_19922;
assign v_19924 = v_1085 & v_1246;
assign v_19926 = v_936 & v_19925;
assign v_19927 = v_940 & v_961;
assign v_19929 = v_937 & v_19928;
assign v_19930 = v_804 & v_962;
assign v_19932 = v_92 & v_19931;
assign v_19933 = v_98 & v_591;
assign v_19936 = v_9600 & v_9796;
assign v_19937 = v_9629 & v_9664;
assign v_19939 = v_9601 & v_19938;
assign v_19940 = v_9506 & v_9630;
assign v_19942 = v_9307 & v_19941;
assign v_19943 = v_9335 & v_9374;
assign v_19945 = v_9308 & v_19944;
assign v_19946 = v_9218 & v_9336;
assign v_19948 = v_9026 & v_19947;
assign v_19949 = v_9051 & v_9086;
assign v_19951 = v_9027 & v_19950;
assign v_19952 = v_8936 & v_9052;
assign v_19954 = v_8729 & v_19953;
assign v_19955 = v_8761 & v_8804;
assign v_19957 = v_8730 & v_19956;
assign v_19958 = v_8640 & v_8762;
assign v_19960 = v_8447 & v_19959;
assign v_19961 = v_8473 & v_8508;
assign v_19963 = v_8448 & v_19962;
assign v_19964 = v_8356 & v_8474;
assign v_19966 = v_8157 & v_19965;
assign v_19967 = v_8185 & v_8224;
assign v_19969 = v_8158 & v_19968;
assign v_19970 = v_8068 & v_8186;
assign v_19972 = v_7876 & v_19971;
assign v_19973 = v_7901 & v_7936;
assign v_19975 = v_7877 & v_19974;
assign v_19976 = v_7786 & v_7902;
assign v_19978 = v_7571 & v_19977;
assign v_19979 = v_7607 & v_7654;
assign v_19981 = v_7572 & v_19980;
assign v_19982 = v_7482 & v_7608;
assign v_19984 = v_7288 & v_19983;
assign v_19985 = v_7315 & v_7350;
assign v_19987 = v_7289 & v_19986;
assign v_19988 = v_7196 & v_7316;
assign v_19990 = v_6997 & v_19989;
assign v_19991 = v_7025 & v_7064;
assign v_19993 = v_6998 & v_19992;
assign v_19994 = v_6908 & v_7026;
assign v_19996 = v_6716 & v_19995;
assign v_19997 = v_6741 & v_6776;
assign v_19999 = v_6717 & v_19998;
assign v_20000 = v_6626 & v_6742;
assign v_20002 = v_6419 & v_20001;
assign v_20003 = v_6451 & v_6494;
assign v_20005 = v_6420 & v_20004;
assign v_20006 = v_6330 & v_6452;
assign v_20008 = v_6137 & v_20007;
assign v_20009 = v_6163 & v_6198;
assign v_20011 = v_6138 & v_20010;
assign v_20012 = v_6046 & v_6164;
assign v_20014 = v_5847 & v_20013;
assign v_20015 = v_5875 & v_5914;
assign v_20017 = v_5848 & v_20016;
assign v_20018 = v_5758 & v_5876;
assign v_20020 = v_5566 & v_20019;
assign v_20021 = v_5591 & v_5626;
assign v_20023 = v_5567 & v_20022;
assign v_20024 = v_5476 & v_5592;
assign v_20026 = v_5253 & v_20025;
assign v_20027 = v_5293 & v_5344;
assign v_20029 = v_5254 & v_20028;
assign v_20030 = v_5164 & v_5294;
assign v_20032 = v_4969 & v_20031;
assign v_20033 = v_4997 & v_5032;
assign v_20035 = v_4970 & v_20034;
assign v_20036 = v_4876 & v_4998;
assign v_20038 = v_4677 & v_20037;
assign v_20039 = v_4705 & v_4744;
assign v_20041 = v_4678 & v_20040;
assign v_20042 = v_4588 & v_4706;
assign v_20044 = v_4396 & v_20043;
assign v_20045 = v_4421 & v_4456;
assign v_20047 = v_4397 & v_20046;
assign v_20048 = v_4306 & v_4422;
assign v_20050 = v_4099 & v_20049;
assign v_20051 = v_4131 & v_4174;
assign v_20053 = v_4100 & v_20052;
assign v_20054 = v_4010 & v_4132;
assign v_20056 = v_3817 & v_20055;
assign v_20057 = v_3843 & v_3878;
assign v_20059 = v_3818 & v_20058;
assign v_20060 = v_3726 & v_3844;
assign v_20062 = v_3527 & v_20061;
assign v_20063 = v_3555 & v_3594;
assign v_20065 = v_3528 & v_20064;
assign v_20066 = v_3438 & v_3556;
assign v_20068 = v_3246 & v_20067;
assign v_20069 = v_3271 & v_3306;
assign v_20071 = v_3247 & v_20070;
assign v_20072 = v_3156 & v_3272;
assign v_20074 = v_2941 & v_20073;
assign v_20075 = v_2977 & v_3024;
assign v_20077 = v_2942 & v_20076;
assign v_20078 = v_2852 & v_2978;
assign v_20080 = v_2658 & v_20079;
assign v_20081 = v_2685 & v_2720;
assign v_20083 = v_2659 & v_20082;
assign v_20084 = v_2566 & v_2686;
assign v_20086 = v_2367 & v_20085;
assign v_20087 = v_2395 & v_2434;
assign v_20089 = v_2368 & v_20088;
assign v_20090 = v_2278 & v_2396;
assign v_20092 = v_2086 & v_20091;
assign v_20093 = v_2111 & v_2146;
assign v_20095 = v_2087 & v_20094;
assign v_20096 = v_1996 & v_2112;
assign v_20098 = v_1789 & v_20097;
assign v_20099 = v_1821 & v_1864;
assign v_20101 = v_1790 & v_20100;
assign v_20102 = v_1700 & v_1822;
assign v_20104 = v_1507 & v_20103;
assign v_20105 = v_1533 & v_1568;
assign v_20107 = v_1508 & v_20106;
assign v_20108 = v_1416 & v_1534;
assign v_20110 = v_1217 & v_20109;
assign v_20111 = v_1245 & v_1284;
assign v_20113 = v_1218 & v_20112;
assign v_20114 = v_1128 & v_1246;
assign v_20116 = v_936 & v_20115;
assign v_20117 = v_961 & v_996;
assign v_20119 = v_937 & v_20118;
assign v_20120 = v_850 & v_962;
assign v_20122 = v_92 & v_20121;
assign v_20123 = v_591 & v_731;
assign v_20126 = v_9600 & v_9808;
assign v_20127 = v_9629 & v_9676;
assign v_20129 = v_9601 & v_20128;
assign v_20130 = v_9518 & v_9630;
assign v_20132 = v_9307 & v_20131;
assign v_20133 = v_9335 & v_9386;
assign v_20135 = v_9308 & v_20134;
assign v_20136 = v_9230 & v_9336;
assign v_20138 = v_9026 & v_20137;
assign v_20139 = v_9051 & v_9098;
assign v_20141 = v_9027 & v_20140;
assign v_20142 = v_8948 & v_9052;
assign v_20144 = v_8729 & v_20143;
assign v_20145 = v_8761 & v_8816;
assign v_20147 = v_8730 & v_20146;
assign v_20148 = v_8652 & v_8762;
assign v_20150 = v_8447 & v_20149;
assign v_20151 = v_8473 & v_8520;
assign v_20153 = v_8448 & v_20152;
assign v_20154 = v_8368 & v_8474;
assign v_20156 = v_8157 & v_20155;
assign v_20157 = v_8185 & v_8236;
assign v_20159 = v_8158 & v_20158;
assign v_20160 = v_8080 & v_8186;
assign v_20162 = v_7876 & v_20161;
assign v_20163 = v_7901 & v_7948;
assign v_20165 = v_7877 & v_20164;
assign v_20166 = v_7798 & v_7902;
assign v_20168 = v_7571 & v_20167;
assign v_20169 = v_7607 & v_7666;
assign v_20171 = v_7572 & v_20170;
assign v_20172 = v_7494 & v_7608;
assign v_20174 = v_7288 & v_20173;
assign v_20175 = v_7315 & v_7362;
assign v_20177 = v_7289 & v_20176;
assign v_20178 = v_7208 & v_7316;
assign v_20180 = v_6997 & v_20179;
assign v_20181 = v_7025 & v_7076;
assign v_20183 = v_6998 & v_20182;
assign v_20184 = v_6920 & v_7026;
assign v_20186 = v_6716 & v_20185;
assign v_20187 = v_6741 & v_6788;
assign v_20189 = v_6717 & v_20188;
assign v_20190 = v_6638 & v_6742;
assign v_20192 = v_6419 & v_20191;
assign v_20193 = v_6451 & v_6506;
assign v_20195 = v_6420 & v_20194;
assign v_20196 = v_6342 & v_6452;
assign v_20198 = v_6137 & v_20197;
assign v_20199 = v_6163 & v_6210;
assign v_20201 = v_6138 & v_20200;
assign v_20202 = v_6058 & v_6164;
assign v_20204 = v_5847 & v_20203;
assign v_20205 = v_5875 & v_5926;
assign v_20207 = v_5848 & v_20206;
assign v_20208 = v_5770 & v_5876;
assign v_20210 = v_5566 & v_20209;
assign v_20211 = v_5591 & v_5638;
assign v_20213 = v_5567 & v_20212;
assign v_20214 = v_5488 & v_5592;
assign v_20216 = v_5253 & v_20215;
assign v_20217 = v_5293 & v_5356;
assign v_20219 = v_5254 & v_20218;
assign v_20220 = v_5176 & v_5294;
assign v_20222 = v_4969 & v_20221;
assign v_20223 = v_4997 & v_5044;
assign v_20225 = v_4970 & v_20224;
assign v_20226 = v_4888 & v_4998;
assign v_20228 = v_4677 & v_20227;
assign v_20229 = v_4705 & v_4756;
assign v_20231 = v_4678 & v_20230;
assign v_20232 = v_4600 & v_4706;
assign v_20234 = v_4396 & v_20233;
assign v_20235 = v_4421 & v_4468;
assign v_20237 = v_4397 & v_20236;
assign v_20238 = v_4318 & v_4422;
assign v_20240 = v_4099 & v_20239;
assign v_20241 = v_4131 & v_4186;
assign v_20243 = v_4100 & v_20242;
assign v_20244 = v_4022 & v_4132;
assign v_20246 = v_3817 & v_20245;
assign v_20247 = v_3843 & v_3890;
assign v_20249 = v_3818 & v_20248;
assign v_20250 = v_3738 & v_3844;
assign v_20252 = v_3527 & v_20251;
assign v_20253 = v_3555 & v_3606;
assign v_20255 = v_3528 & v_20254;
assign v_20256 = v_3450 & v_3556;
assign v_20258 = v_3246 & v_20257;
assign v_20259 = v_3271 & v_3318;
assign v_20261 = v_3247 & v_20260;
assign v_20262 = v_3168 & v_3272;
assign v_20264 = v_2941 & v_20263;
assign v_20265 = v_2977 & v_3036;
assign v_20267 = v_2942 & v_20266;
assign v_20268 = v_2864 & v_2978;
assign v_20270 = v_2658 & v_20269;
assign v_20271 = v_2685 & v_2732;
assign v_20273 = v_2659 & v_20272;
assign v_20274 = v_2578 & v_2686;
assign v_20276 = v_2367 & v_20275;
assign v_20277 = v_2395 & v_2446;
assign v_20279 = v_2368 & v_20278;
assign v_20280 = v_2290 & v_2396;
assign v_20282 = v_2086 & v_20281;
assign v_20283 = v_2111 & v_2158;
assign v_20285 = v_2087 & v_20284;
assign v_20286 = v_2008 & v_2112;
assign v_20288 = v_1789 & v_20287;
assign v_20289 = v_1821 & v_1876;
assign v_20291 = v_1790 & v_20290;
assign v_20292 = v_1712 & v_1822;
assign v_20294 = v_1507 & v_20293;
assign v_20295 = v_1533 & v_1580;
assign v_20297 = v_1508 & v_20296;
assign v_20298 = v_1428 & v_1534;
assign v_20300 = v_1217 & v_20299;
assign v_20301 = v_1245 & v_1296;
assign v_20303 = v_1218 & v_20302;
assign v_20304 = v_1140 & v_1246;
assign v_20306 = v_936 & v_20305;
assign v_20307 = v_961 & v_1008;
assign v_20309 = v_937 & v_20308;
assign v_20310 = v_862 & v_962;
assign v_20312 = v_92 & v_20311;
assign v_20313 = v_591 & v_741;
assign v_20316 = v_9600 & v_9820;
assign v_20317 = v_9629 & v_9688;
assign v_20319 = v_9601 & v_20318;
assign v_20320 = v_9530 & v_9630;
assign v_20322 = v_9307 & v_20321;
assign v_20323 = v_9335 & v_9398;
assign v_20325 = v_9308 & v_20324;
assign v_20326 = v_9242 & v_9336;
assign v_20328 = v_9026 & v_20327;
assign v_20329 = v_9051 & v_9110;
assign v_20331 = v_9027 & v_20330;
assign v_20332 = v_8960 & v_9052;
assign v_20334 = v_8729 & v_20333;
assign v_20335 = v_8761 & v_8828;
assign v_20337 = v_8730 & v_20336;
assign v_20338 = v_8664 & v_8762;
assign v_20340 = v_8447 & v_20339;
assign v_20341 = v_8473 & v_8532;
assign v_20343 = v_8448 & v_20342;
assign v_20344 = v_8380 & v_8474;
assign v_20346 = v_8157 & v_20345;
assign v_20347 = v_8185 & v_8248;
assign v_20349 = v_8158 & v_20348;
assign v_20350 = v_8092 & v_8186;
assign v_20352 = v_7876 & v_20351;
assign v_20353 = v_7901 & v_7960;
assign v_20355 = v_7877 & v_20354;
assign v_20356 = v_7810 & v_7902;
assign v_20358 = v_7571 & v_20357;
assign v_20359 = v_7607 & v_7678;
assign v_20361 = v_7572 & v_20360;
assign v_20362 = v_7506 & v_7608;
assign v_20364 = v_7288 & v_20363;
assign v_20365 = v_7315 & v_7374;
assign v_20367 = v_7289 & v_20366;
assign v_20368 = v_7220 & v_7316;
assign v_20370 = v_6997 & v_20369;
assign v_20371 = v_7025 & v_7088;
assign v_20373 = v_6998 & v_20372;
assign v_20374 = v_6932 & v_7026;
assign v_20376 = v_6716 & v_20375;
assign v_20377 = v_6741 & v_6800;
assign v_20379 = v_6717 & v_20378;
assign v_20380 = v_6650 & v_6742;
assign v_20382 = v_6419 & v_20381;
assign v_20383 = v_6451 & v_6518;
assign v_20385 = v_6420 & v_20384;
assign v_20386 = v_6354 & v_6452;
assign v_20388 = v_6137 & v_20387;
assign v_20389 = v_6163 & v_6222;
assign v_20391 = v_6138 & v_20390;
assign v_20392 = v_6070 & v_6164;
assign v_20394 = v_5847 & v_20393;
assign v_20395 = v_5875 & v_5938;
assign v_20397 = v_5848 & v_20396;
assign v_20398 = v_5782 & v_5876;
assign v_20400 = v_5566 & v_20399;
assign v_20401 = v_5591 & v_5650;
assign v_20403 = v_5567 & v_20402;
assign v_20404 = v_5500 & v_5592;
assign v_20406 = v_5253 & v_20405;
assign v_20407 = v_5293 & v_5368;
assign v_20409 = v_5254 & v_20408;
assign v_20410 = v_5188 & v_5294;
assign v_20412 = v_4969 & v_20411;
assign v_20413 = v_4997 & v_5056;
assign v_20415 = v_4970 & v_20414;
assign v_20416 = v_4900 & v_4998;
assign v_20418 = v_4677 & v_20417;
assign v_20419 = v_4705 & v_4768;
assign v_20421 = v_4678 & v_20420;
assign v_20422 = v_4612 & v_4706;
assign v_20424 = v_4396 & v_20423;
assign v_20425 = v_4421 & v_4480;
assign v_20427 = v_4397 & v_20426;
assign v_20428 = v_4330 & v_4422;
assign v_20430 = v_4099 & v_20429;
assign v_20431 = v_4131 & v_4198;
assign v_20433 = v_4100 & v_20432;
assign v_20434 = v_4034 & v_4132;
assign v_20436 = v_3817 & v_20435;
assign v_20437 = v_3843 & v_3902;
assign v_20439 = v_3818 & v_20438;
assign v_20440 = v_3750 & v_3844;
assign v_20442 = v_3527 & v_20441;
assign v_20443 = v_3555 & v_3618;
assign v_20445 = v_3528 & v_20444;
assign v_20446 = v_3462 & v_3556;
assign v_20448 = v_3246 & v_20447;
assign v_20449 = v_3271 & v_3330;
assign v_20451 = v_3247 & v_20450;
assign v_20452 = v_3180 & v_3272;
assign v_20454 = v_2941 & v_20453;
assign v_20455 = v_2977 & v_3048;
assign v_20457 = v_2942 & v_20456;
assign v_20458 = v_2876 & v_2978;
assign v_20460 = v_2658 & v_20459;
assign v_20461 = v_2685 & v_2744;
assign v_20463 = v_2659 & v_20462;
assign v_20464 = v_2590 & v_2686;
assign v_20466 = v_2367 & v_20465;
assign v_20467 = v_2395 & v_2458;
assign v_20469 = v_2368 & v_20468;
assign v_20470 = v_2302 & v_2396;
assign v_20472 = v_2086 & v_20471;
assign v_20473 = v_2111 & v_2170;
assign v_20475 = v_2087 & v_20474;
assign v_20476 = v_2020 & v_2112;
assign v_20478 = v_1789 & v_20477;
assign v_20479 = v_1821 & v_1888;
assign v_20481 = v_1790 & v_20480;
assign v_20482 = v_1724 & v_1822;
assign v_20484 = v_1507 & v_20483;
assign v_20485 = v_1533 & v_1592;
assign v_20487 = v_1508 & v_20486;
assign v_20488 = v_1440 & v_1534;
assign v_20490 = v_1217 & v_20489;
assign v_20491 = v_1245 & v_1308;
assign v_20493 = v_1218 & v_20492;
assign v_20494 = v_1152 & v_1246;
assign v_20496 = v_936 & v_20495;
assign v_20497 = v_961 & v_1020;
assign v_20499 = v_937 & v_20498;
assign v_20500 = v_874 & v_962;
assign v_20502 = v_92 & v_20501;
assign v_20503 = v_591 & v_751;
assign v_20506 = v_9600 & v_9832;
assign v_20507 = v_9629 & v_9700;
assign v_20509 = v_9601 & v_20508;
assign v_20510 = v_9542 & v_9630;
assign v_20512 = v_9307 & v_20511;
assign v_20513 = v_9335 & v_9410;
assign v_20515 = v_9308 & v_20514;
assign v_20516 = v_9254 & v_9336;
assign v_20518 = v_9026 & v_20517;
assign v_20519 = v_9051 & v_9122;
assign v_20521 = v_9027 & v_20520;
assign v_20522 = v_8972 & v_9052;
assign v_20524 = v_8729 & v_20523;
assign v_20525 = v_8761 & v_8840;
assign v_20527 = v_8730 & v_20526;
assign v_20528 = v_8676 & v_8762;
assign v_20530 = v_8447 & v_20529;
assign v_20531 = v_8473 & v_8544;
assign v_20533 = v_8448 & v_20532;
assign v_20534 = v_8392 & v_8474;
assign v_20536 = v_8157 & v_20535;
assign v_20537 = v_8185 & v_8260;
assign v_20539 = v_8158 & v_20538;
assign v_20540 = v_8104 & v_8186;
assign v_20542 = v_7876 & v_20541;
assign v_20543 = v_7901 & v_7972;
assign v_20545 = v_7877 & v_20544;
assign v_20546 = v_7822 & v_7902;
assign v_20548 = v_7571 & v_20547;
assign v_20549 = v_7607 & v_7690;
assign v_20551 = v_7572 & v_20550;
assign v_20552 = v_7518 & v_7608;
assign v_20554 = v_7288 & v_20553;
assign v_20555 = v_7315 & v_7386;
assign v_20557 = v_7289 & v_20556;
assign v_20558 = v_7232 & v_7316;
assign v_20560 = v_6997 & v_20559;
assign v_20561 = v_7025 & v_7100;
assign v_20563 = v_6998 & v_20562;
assign v_20564 = v_6944 & v_7026;
assign v_20566 = v_6716 & v_20565;
assign v_20567 = v_6741 & v_6812;
assign v_20569 = v_6717 & v_20568;
assign v_20570 = v_6662 & v_6742;
assign v_20572 = v_6419 & v_20571;
assign v_20573 = v_6451 & v_6530;
assign v_20575 = v_6420 & v_20574;
assign v_20576 = v_6366 & v_6452;
assign v_20578 = v_6137 & v_20577;
assign v_20579 = v_6163 & v_6234;
assign v_20581 = v_6138 & v_20580;
assign v_20582 = v_6082 & v_6164;
assign v_20584 = v_5847 & v_20583;
assign v_20585 = v_5875 & v_5950;
assign v_20587 = v_5848 & v_20586;
assign v_20588 = v_5794 & v_5876;
assign v_20590 = v_5566 & v_20589;
assign v_20591 = v_5591 & v_5662;
assign v_20593 = v_5567 & v_20592;
assign v_20594 = v_5512 & v_5592;
assign v_20596 = v_5253 & v_20595;
assign v_20597 = v_5293 & v_5380;
assign v_20599 = v_5254 & v_20598;
assign v_20600 = v_5200 & v_5294;
assign v_20602 = v_4969 & v_20601;
assign v_20603 = v_4997 & v_5068;
assign v_20605 = v_4970 & v_20604;
assign v_20606 = v_4912 & v_4998;
assign v_20608 = v_4677 & v_20607;
assign v_20609 = v_4705 & v_4780;
assign v_20611 = v_4678 & v_20610;
assign v_20612 = v_4624 & v_4706;
assign v_20614 = v_4396 & v_20613;
assign v_20615 = v_4421 & v_4492;
assign v_20617 = v_4397 & v_20616;
assign v_20618 = v_4342 & v_4422;
assign v_20620 = v_4099 & v_20619;
assign v_20621 = v_4131 & v_4210;
assign v_20623 = v_4100 & v_20622;
assign v_20624 = v_4046 & v_4132;
assign v_20626 = v_3817 & v_20625;
assign v_20627 = v_3843 & v_3914;
assign v_20629 = v_3818 & v_20628;
assign v_20630 = v_3762 & v_3844;
assign v_20632 = v_3527 & v_20631;
assign v_20633 = v_3555 & v_3630;
assign v_20635 = v_3528 & v_20634;
assign v_20636 = v_3474 & v_3556;
assign v_20638 = v_3246 & v_20637;
assign v_20639 = v_3271 & v_3342;
assign v_20641 = v_3247 & v_20640;
assign v_20642 = v_3192 & v_3272;
assign v_20644 = v_2941 & v_20643;
assign v_20645 = v_2977 & v_3060;
assign v_20647 = v_2942 & v_20646;
assign v_20648 = v_2888 & v_2978;
assign v_20650 = v_2658 & v_20649;
assign v_20651 = v_2685 & v_2756;
assign v_20653 = v_2659 & v_20652;
assign v_20654 = v_2602 & v_2686;
assign v_20656 = v_2367 & v_20655;
assign v_20657 = v_2395 & v_2470;
assign v_20659 = v_2368 & v_20658;
assign v_20660 = v_2314 & v_2396;
assign v_20662 = v_2086 & v_20661;
assign v_20663 = v_2111 & v_2182;
assign v_20665 = v_2087 & v_20664;
assign v_20666 = v_2032 & v_2112;
assign v_20668 = v_1789 & v_20667;
assign v_20669 = v_1821 & v_1900;
assign v_20671 = v_1790 & v_20670;
assign v_20672 = v_1736 & v_1822;
assign v_20674 = v_1507 & v_20673;
assign v_20675 = v_1533 & v_1604;
assign v_20677 = v_1508 & v_20676;
assign v_20678 = v_1452 & v_1534;
assign v_20680 = v_1217 & v_20679;
assign v_20681 = v_1245 & v_1320;
assign v_20683 = v_1218 & v_20682;
assign v_20684 = v_1164 & v_1246;
assign v_20686 = v_936 & v_20685;
assign v_20687 = v_961 & v_1032;
assign v_20689 = v_937 & v_20688;
assign v_20690 = v_886 & v_962;
assign v_20692 = v_92 & v_20691;
assign v_20693 = v_591 & v_761;
assign v_20696 = v_9600 & v_9844;
assign v_20697 = v_9629 & v_9712;
assign v_20699 = v_9601 & v_20698;
assign v_20700 = v_9554 & v_9630;
assign v_20702 = v_9307 & v_20701;
assign v_20703 = v_9335 & v_9422;
assign v_20705 = v_9308 & v_20704;
assign v_20706 = v_9266 & v_9336;
assign v_20708 = v_9026 & v_20707;
assign v_20709 = v_9051 & v_9134;
assign v_20711 = v_9027 & v_20710;
assign v_20712 = v_8984 & v_9052;
assign v_20714 = v_8729 & v_20713;
assign v_20715 = v_8761 & v_8852;
assign v_20717 = v_8730 & v_20716;
assign v_20718 = v_8688 & v_8762;
assign v_20720 = v_8447 & v_20719;
assign v_20721 = v_8473 & v_8556;
assign v_20723 = v_8448 & v_20722;
assign v_20724 = v_8404 & v_8474;
assign v_20726 = v_8157 & v_20725;
assign v_20727 = v_8185 & v_8272;
assign v_20729 = v_8158 & v_20728;
assign v_20730 = v_8116 & v_8186;
assign v_20732 = v_7876 & v_20731;
assign v_20733 = v_7901 & v_7984;
assign v_20735 = v_7877 & v_20734;
assign v_20736 = v_7834 & v_7902;
assign v_20738 = v_7571 & v_20737;
assign v_20739 = v_7607 & v_7702;
assign v_20741 = v_7572 & v_20740;
assign v_20742 = v_7530 & v_7608;
assign v_20744 = v_7288 & v_20743;
assign v_20745 = v_7315 & v_7398;
assign v_20747 = v_7289 & v_20746;
assign v_20748 = v_7244 & v_7316;
assign v_20750 = v_6997 & v_20749;
assign v_20751 = v_7025 & v_7112;
assign v_20753 = v_6998 & v_20752;
assign v_20754 = v_6956 & v_7026;
assign v_20756 = v_6716 & v_20755;
assign v_20757 = v_6741 & ~v_6824;
assign v_20759 = v_6717 & v_20758;
assign v_20760 = v_6674 & v_6742;
assign v_20762 = v_6419 & v_20761;
assign v_20763 = v_6451 & v_6542;
assign v_20765 = v_6420 & v_20764;
assign v_20766 = v_6378 & v_6452;
assign v_20768 = v_6137 & v_20767;
assign v_20769 = v_6163 & v_6246;
assign v_20771 = v_6138 & v_20770;
assign v_20772 = ~v_6094 & v_6164;
assign v_20774 = v_5847 & v_20773;
assign v_20775 = v_5875 & v_5962;
assign v_20777 = v_5848 & v_20776;
assign v_20778 = ~v_5806 & v_5876;
assign v_20780 = v_5566 & v_20779;
assign v_20781 = v_5591 & v_5674;
assign v_20783 = v_5567 & v_20782;
assign v_20784 = v_5524 & v_5592;
assign v_20786 = v_5253 & v_20785;
assign v_20787 = v_5293 & v_5392;
assign v_20789 = v_5254 & v_20788;
assign v_20790 = v_5212 & v_5294;
assign v_20792 = v_4969 & v_20791;
assign v_20793 = v_4997 & v_5080;
assign v_20795 = v_4970 & v_20794;
assign v_20796 = v_4924 & v_4998;
assign v_20798 = v_4677 & v_20797;
assign v_20799 = v_4705 & v_4792;
assign v_20801 = v_4678 & v_20800;
assign v_20802 = v_4636 & v_4706;
assign v_20804 = v_4396 & v_20803;
assign v_20805 = v_4421 & v_4504;
assign v_20807 = v_4397 & v_20806;
assign v_20808 = v_4354 & v_4422;
assign v_20810 = v_4099 & v_20809;
assign v_20811 = v_4131 & v_4222;
assign v_20813 = v_4100 & v_20812;
assign v_20814 = v_4058 & v_4132;
assign v_20816 = v_3817 & v_20815;
assign v_20817 = v_3843 & v_3926;
assign v_20819 = v_3818 & v_20818;
assign v_20820 = v_3774 & v_3844;
assign v_20822 = v_3527 & v_20821;
assign v_20823 = v_3555 & v_3642;
assign v_20825 = v_3528 & v_20824;
assign v_20826 = v_3486 & v_3556;
assign v_20828 = v_3246 & v_20827;
assign v_20829 = v_3271 & v_3354;
assign v_20831 = v_3247 & v_20830;
assign v_20832 = ~v_3204 & v_3272;
assign v_20834 = v_2941 & v_20833;
assign v_20835 = v_2977 & v_3072;
assign v_20837 = v_2942 & v_20836;
assign v_20838 = v_2900 & v_2978;
assign v_20840 = v_2658 & v_20839;
assign v_20841 = v_2685 & v_2768;
assign v_20843 = v_2659 & v_20842;
assign v_20844 = v_2614 & v_2686;
assign v_20846 = v_2367 & v_20845;
assign v_20847 = v_2395 & v_2482;
assign v_20849 = v_2368 & v_20848;
assign v_20850 = v_2326 & v_2396;
assign v_20852 = v_2086 & v_20851;
assign v_20853 = v_2111 & v_2194;
assign v_20855 = v_2087 & v_20854;
assign v_20856 = v_2044 & v_2112;
assign v_20858 = v_1789 & v_20857;
assign v_20859 = v_1821 & v_1912;
assign v_20861 = v_1790 & v_20860;
assign v_20862 = v_1748 & v_1822;
assign v_20864 = v_1507 & v_20863;
assign v_20865 = v_1533 & v_1616;
assign v_20867 = v_1508 & v_20866;
assign v_20868 = v_1464 & v_1534;
assign v_20870 = v_1217 & v_20869;
assign v_20871 = v_1245 & v_1332;
assign v_20873 = v_1218 & v_20872;
assign v_20874 = v_1176 & v_1246;
assign v_20876 = v_936 & v_20875;
assign v_20877 = v_961 & v_1044;
assign v_20879 = v_937 & v_20878;
assign v_20880 = v_898 & v_962;
assign v_20882 = v_92 & v_20881;
assign v_20883 = v_591 & v_771;
assign v_20886 = v_9600 & ~v_9872;
assign v_20887 = v_9629 & ~v_9740;
assign v_20889 = v_9601 & v_20888;
assign v_20890 = ~v_9582 & v_9630;
assign v_20892 = v_9307 & v_20891;
assign v_20893 = v_9335 & ~v_9450;
assign v_20895 = v_9308 & v_20894;
assign v_20896 = ~v_9294 & v_9336;
assign v_20898 = v_9026 & v_20897;
assign v_20899 = v_9051 & ~v_9162;
assign v_20901 = v_9027 & v_20900;
assign v_20902 = ~v_9012 & v_9052;
assign v_20904 = v_8729 & v_20903;
assign v_20905 = v_8761 & ~v_8880;
assign v_20907 = v_8730 & v_20906;
assign v_20908 = ~v_8716 & v_8762;
assign v_20910 = v_8447 & v_20909;
assign v_20911 = v_8473 & ~v_8584;
assign v_20913 = v_8448 & v_20912;
assign v_20914 = v_8432 & v_8474;
assign v_20916 = v_8157 & v_20915;
assign v_20917 = v_8185 & v_8300;
assign v_20919 = v_8158 & v_20918;
assign v_20920 = v_8144 & v_8186;
assign v_20922 = v_7876 & v_20921;
assign v_20923 = v_7901 & ~v_8012;
assign v_20925 = v_7877 & v_20924;
assign v_20926 = ~v_7862 & v_7902;
assign v_20928 = v_7571 & v_20927;
assign v_20929 = v_7607 & ~v_7730;
assign v_20931 = v_7572 & v_20930;
assign v_20932 = ~v_7558 & v_7608;
assign v_20934 = v_7288 & v_20933;
assign v_20935 = v_7315 & ~v_7426;
assign v_20937 = v_7289 & v_20936;
assign v_20938 = v_7272 & v_7316;
assign v_20940 = v_6997 & v_20939;
assign v_20941 = v_7025 & ~v_7140;
assign v_20943 = v_6998 & v_20942;
assign v_20944 = v_6984 & v_7026;
assign v_20946 = v_6716 & v_20945;
assign v_20947 = v_6741 & v_6852;
assign v_20949 = v_6717 & v_20948;
assign v_20950 = v_6702 & v_6742;
assign v_20952 = v_6419 & v_20951;
assign v_20953 = v_6451 & ~v_6570;
assign v_20955 = v_6420 & v_20954;
assign v_20956 = ~v_6406 & v_6452;
assign v_20958 = v_6137 & v_20957;
assign v_20959 = v_6163 & v_6274;
assign v_20961 = v_6138 & v_20960;
assign v_20962 = v_6122 & v_6164;
assign v_20964 = v_5847 & v_20963;
assign v_20965 = v_5875 & v_5990;
assign v_20967 = v_5848 & v_20966;
assign v_20968 = v_5834 & v_5876;
assign v_20970 = v_5566 & v_20969;
assign v_20971 = v_5591 & v_5702;
assign v_20973 = v_5567 & v_20972;
assign v_20974 = v_5552 & v_5592;
assign v_20976 = v_5253 & v_20975;
assign v_20977 = v_5293 & ~v_5420;
assign v_20979 = v_5254 & v_20978;
assign v_20980 = ~v_5240 & v_5294;
assign v_20982 = v_4969 & v_20981;
assign v_20983 = v_4997 & v_5108;
assign v_20985 = v_4970 & v_20984;
assign v_20986 = v_4952 & v_4998;
assign v_20988 = v_4677 & v_20987;
assign v_20989 = v_4705 & v_4820;
assign v_20991 = v_4678 & v_20990;
assign v_20992 = v_4664 & v_4706;
assign v_20994 = v_4396 & v_20993;
assign v_20995 = v_4421 & v_4532;
assign v_20997 = v_4397 & v_20996;
assign v_20998 = v_4382 & v_4422;
assign v_21000 = v_4099 & v_20999;
assign v_21001 = v_4131 & ~v_4250;
assign v_21003 = v_4100 & v_21002;
assign v_21004 = ~v_4086 & v_4132;
assign v_21006 = v_3817 & v_21005;
assign v_21007 = v_3843 & ~v_3954;
assign v_21009 = v_3818 & v_21008;
assign v_21010 = ~v_3802 & v_3844;
assign v_21012 = v_3527 & v_21011;
assign v_21013 = v_3555 & ~v_3670;
assign v_21015 = v_3528 & v_21014;
assign v_21016 = v_3514 & v_3556;
assign v_21018 = v_3246 & v_21017;
assign v_21019 = v_3271 & ~v_3382;
assign v_21021 = v_3247 & v_21020;
assign v_21022 = v_3232 & v_3272;
assign v_21024 = v_2941 & v_21023;
assign v_21025 = v_2977 & ~v_3100;
assign v_21027 = v_2942 & v_21026;
assign v_21028 = ~v_2928 & v_2978;
assign v_21030 = v_2658 & v_21029;
assign v_21031 = v_2685 & ~v_2796;
assign v_21033 = v_2659 & v_21032;
assign v_21034 = ~v_2642 & v_2686;
assign v_21036 = v_2367 & v_21035;
assign v_21037 = v_2395 & ~v_2510;
assign v_21039 = v_2368 & v_21038;
assign v_21040 = v_2354 & v_2396;
assign v_21042 = v_2086 & v_21041;
assign v_21043 = v_2111 & v_2222;
assign v_21045 = v_2087 & v_21044;
assign v_21046 = v_2072 & v_2112;
assign v_21048 = v_1789 & v_21047;
assign v_21049 = v_1821 & ~v_1940;
assign v_21051 = v_1790 & v_21050;
assign v_21052 = ~v_1776 & v_1822;
assign v_21054 = v_1507 & v_21053;
assign v_21055 = v_1533 & ~v_1644;
assign v_21057 = v_1508 & v_21056;
assign v_21058 = ~v_1492 & v_1534;
assign v_21060 = v_1217 & v_21059;
assign v_21061 = v_1245 & ~v_1360;
assign v_21063 = v_1218 & v_21062;
assign v_21064 = ~v_1204 & v_1246;
assign v_21066 = v_936 & v_21065;
assign v_21067 = v_961 & ~v_1072;
assign v_21069 = v_937 & v_21068;
assign v_21070 = ~v_922 & v_962;
assign v_21072 = v_92 & v_21071;
assign v_21073 = v_591 & ~v_793;
assign v_21076 = v_9601 & v_9784;
assign v_21077 = v_9630 & v_9652;
assign v_21079 = v_9307 & v_21078;
assign v_21080 = v_9335 & v_9494;
assign v_21082 = v_9308 & v_21081;
assign v_21083 = v_9336 & v_9362;
assign v_21085 = v_9026 & v_21084;
assign v_21086 = v_9051 & v_9206;
assign v_21088 = v_9027 & v_21087;
assign v_21089 = v_9052 & v_9074;
assign v_21091 = v_8729 & v_21090;
assign v_21092 = v_8761 & v_8924;
assign v_21094 = v_8730 & v_21093;
assign v_21095 = v_8762 & v_8792;
assign v_21097 = v_8447 & v_21096;
assign v_21098 = v_8473 & v_8628;
assign v_21100 = v_8448 & v_21099;
assign v_21101 = v_8474 & v_8496;
assign v_21103 = v_8157 & v_21102;
assign v_21104 = v_8185 & v_8344;
assign v_21106 = v_8158 & v_21105;
assign v_21107 = v_8186 & v_8212;
assign v_21109 = v_7876 & v_21108;
assign v_21110 = v_7901 & v_8056;
assign v_21112 = v_7877 & v_21111;
assign v_21113 = v_7902 & v_7924;
assign v_21115 = v_7571 & v_21114;
assign v_21116 = v_7607 & v_7774;
assign v_21118 = v_7572 & v_21117;
assign v_21119 = v_7608 & v_7642;
assign v_21121 = v_7288 & v_21120;
assign v_21122 = v_7315 & v_7470;
assign v_21124 = v_7289 & v_21123;
assign v_21125 = v_7316 & v_7338;
assign v_21127 = v_6997 & v_21126;
assign v_21128 = v_7025 & v_7184;
assign v_21130 = v_6998 & v_21129;
assign v_21131 = v_7026 & v_7052;
assign v_21133 = v_6716 & v_21132;
assign v_21134 = v_6741 & v_6896;
assign v_21136 = v_6717 & v_21135;
assign v_21137 = v_6742 & v_6764;
assign v_21139 = v_6419 & v_21138;
assign v_21140 = v_6451 & v_6614;
assign v_21142 = v_6420 & v_21141;
assign v_21143 = v_6452 & v_6482;
assign v_21145 = v_6137 & v_21144;
assign v_21146 = v_6163 & v_6318;
assign v_21148 = v_6138 & v_21147;
assign v_21149 = v_6164 & v_6186;
assign v_21151 = v_5847 & v_21150;
assign v_21152 = v_5875 & v_6034;
assign v_21154 = v_5848 & v_21153;
assign v_21155 = v_5876 & v_5902;
assign v_21157 = v_5566 & v_21156;
assign v_21158 = v_5591 & v_5746;
assign v_21160 = v_5567 & v_21159;
assign v_21161 = v_5592 & v_5614;
assign v_21163 = v_5253 & v_21162;
assign v_21164 = v_5293 & v_5464;
assign v_21166 = v_5254 & v_21165;
assign v_21167 = v_5294 & v_5332;
assign v_21169 = v_4969 & v_21168;
assign v_21170 = v_4997 & v_5152;
assign v_21172 = v_4970 & v_21171;
assign v_21173 = v_4998 & v_5020;
assign v_21175 = v_4677 & v_21174;
assign v_21176 = v_4705 & v_4864;
assign v_21178 = v_4678 & v_21177;
assign v_21179 = v_4706 & v_4732;
assign v_21181 = v_4396 & v_21180;
assign v_21182 = v_4421 & v_4576;
assign v_21184 = v_4397 & v_21183;
assign v_21185 = v_4422 & v_4444;
assign v_21187 = v_4099 & v_21186;
assign v_21188 = v_4131 & v_4294;
assign v_21190 = v_4100 & v_21189;
assign v_21191 = v_4132 & v_4162;
assign v_21193 = v_3817 & v_21192;
assign v_21194 = v_3843 & v_3998;
assign v_21196 = v_3818 & v_21195;
assign v_21197 = v_3844 & v_3866;
assign v_21199 = v_3527 & v_21198;
assign v_21200 = v_3555 & v_3714;
assign v_21202 = v_3528 & v_21201;
assign v_21203 = v_3556 & v_3582;
assign v_21205 = v_3246 & v_21204;
assign v_21206 = v_3271 & v_3426;
assign v_21208 = v_3247 & v_21207;
assign v_21209 = v_3272 & v_3294;
assign v_21211 = v_2941 & v_21210;
assign v_21212 = v_2977 & v_3144;
assign v_21214 = v_2942 & v_21213;
assign v_21215 = v_2978 & v_3012;
assign v_21217 = v_2658 & v_21216;
assign v_21218 = v_2685 & v_2840;
assign v_21220 = v_2659 & v_21219;
assign v_21221 = v_2686 & v_2708;
assign v_21223 = v_2367 & v_21222;
assign v_21224 = v_2395 & v_2554;
assign v_21226 = v_2368 & v_21225;
assign v_21227 = v_2396 & v_2422;
assign v_21229 = v_2086 & v_21228;
assign v_21230 = v_2111 & v_2266;
assign v_21232 = v_2087 & v_21231;
assign v_21233 = v_2112 & v_2134;
assign v_21235 = v_1789 & v_21234;
assign v_21236 = v_1821 & v_1984;
assign v_21238 = v_1790 & v_21237;
assign v_21239 = v_1822 & v_1852;
assign v_21241 = v_1507 & v_21240;
assign v_21242 = v_1533 & v_1688;
assign v_21244 = v_1508 & v_21243;
assign v_21245 = v_1534 & v_1556;
assign v_21247 = v_1217 & v_21246;
assign v_21248 = v_1245 & v_1404;
assign v_21250 = v_1218 & v_21249;
assign v_21251 = v_1246 & v_1272;
assign v_21253 = v_936 & v_21252;
assign v_21254 = v_961 & v_1116;
assign v_21256 = v_937 & v_21255;
assign v_21257 = v_962 & v_984;
assign v_21259 = v_92 & v_21258;
assign v_21260 = v_591 & v_838;
assign v_21262 = v_94 & v_21261;
assign v_21263 = v_593 & v_721;
assign v_21265 = v_9601 & v_9753;
assign v_21266 = v_9604 & v_9630;
assign v_21268 = v_9307 & v_21267;
assign v_21269 = v_9335 & v_9463;
assign v_21271 = v_9308 & v_21270;
assign v_21272 = v_9311 & v_9336;
assign v_21274 = v_9026 & v_21273;
assign v_21275 = v_9051 & v_9175;
assign v_21277 = v_9027 & v_21276;
assign v_21278 = v_9030 & v_9052;
assign v_21280 = v_8729 & v_21279;
assign v_21281 = v_8761 & v_8893;
assign v_21283 = v_8730 & v_21282;
assign v_21284 = v_8733 & v_8762;
assign v_21286 = v_8447 & v_21285;
assign v_21287 = v_8473 & v_8597;
assign v_21289 = v_8448 & v_21288;
assign v_21290 = v_8451 & v_8474;
assign v_21292 = v_8157 & v_21291;
assign v_21293 = v_8185 & v_8313;
assign v_21295 = v_8158 & v_21294;
assign v_21296 = v_8161 & v_8186;
assign v_21298 = v_7876 & v_21297;
assign v_21299 = v_7901 & v_8025;
assign v_21301 = v_7877 & v_21300;
assign v_21302 = v_7880 & v_7902;
assign v_21304 = v_7571 & v_21303;
assign v_21305 = v_7607 & v_7743;
assign v_21307 = v_7572 & v_21306;
assign v_21308 = v_7575 & v_7608;
assign v_21310 = v_7288 & v_21309;
assign v_21311 = v_7315 & v_7439;
assign v_21313 = v_7289 & v_21312;
assign v_21314 = v_7292 & v_7316;
assign v_21316 = v_6997 & v_21315;
assign v_21317 = v_7025 & v_7153;
assign v_21319 = v_6998 & v_21318;
assign v_21320 = v_7001 & v_7026;
assign v_21322 = v_6716 & v_21321;
assign v_21323 = v_6741 & v_6865;
assign v_21325 = v_6717 & v_21324;
assign v_21326 = v_6720 & v_6742;
assign v_21328 = v_6419 & v_21327;
assign v_21329 = v_6451 & v_6583;
assign v_21331 = v_6420 & v_21330;
assign v_21332 = v_6423 & v_6452;
assign v_21334 = v_6137 & v_21333;
assign v_21335 = v_6163 & v_6287;
assign v_21337 = v_6138 & v_21336;
assign v_21338 = v_6141 & v_6164;
assign v_21340 = v_5847 & v_21339;
assign v_21341 = v_5875 & v_6003;
assign v_21343 = v_5848 & v_21342;
assign v_21344 = v_5851 & v_5876;
assign v_21346 = v_5566 & v_21345;
assign v_21347 = v_5591 & v_5715;
assign v_21349 = v_5567 & v_21348;
assign v_21350 = v_5570 & v_5592;
assign v_21352 = v_5253 & v_21351;
assign v_21353 = v_5293 & v_5433;
assign v_21355 = v_5254 & v_21354;
assign v_21356 = v_5257 & v_5294;
assign v_21358 = v_4969 & v_21357;
assign v_21359 = v_4997 & v_5121;
assign v_21361 = v_4970 & v_21360;
assign v_21362 = v_4973 & v_4998;
assign v_21364 = v_4677 & v_21363;
assign v_21365 = v_4705 & v_4833;
assign v_21367 = v_4678 & v_21366;
assign v_21368 = v_4681 & v_4706;
assign v_21370 = v_4396 & v_21369;
assign v_21371 = v_4421 & v_4545;
assign v_21373 = v_4397 & v_21372;
assign v_21374 = v_4400 & v_4422;
assign v_21376 = v_4099 & v_21375;
assign v_21377 = v_4131 & v_4263;
assign v_21379 = v_4100 & v_21378;
assign v_21380 = v_4103 & v_4132;
assign v_21382 = v_3817 & v_21381;
assign v_21383 = v_3843 & v_3967;
assign v_21385 = v_3818 & v_21384;
assign v_21386 = v_3821 & v_3844;
assign v_21388 = v_3527 & v_21387;
assign v_21389 = v_3555 & v_3683;
assign v_21391 = v_3528 & v_21390;
assign v_21392 = v_3531 & v_3556;
assign v_21394 = v_3246 & v_21393;
assign v_21395 = v_3271 & v_3395;
assign v_21397 = v_3247 & v_21396;
assign v_21398 = v_3250 & v_3272;
assign v_21400 = v_2941 & v_21399;
assign v_21401 = v_2977 & v_3113;
assign v_21403 = v_2942 & v_21402;
assign v_21404 = v_2945 & v_2978;
assign v_21406 = v_2658 & v_21405;
assign v_21407 = v_2685 & v_2809;
assign v_21409 = v_2659 & v_21408;
assign v_21410 = v_2662 & v_2686;
assign v_21412 = v_2367 & v_21411;
assign v_21413 = v_2395 & v_2523;
assign v_21415 = v_2368 & v_21414;
assign v_21416 = v_2371 & v_2396;
assign v_21418 = v_2086 & v_21417;
assign v_21419 = v_2111 & v_2235;
assign v_21421 = v_2087 & v_21420;
assign v_21422 = v_2090 & v_2112;
assign v_21424 = v_1789 & v_21423;
assign v_21425 = v_1821 & v_1953;
assign v_21427 = v_1790 & v_21426;
assign v_21428 = v_1793 & v_1822;
assign v_21430 = v_1507 & v_21429;
assign v_21431 = v_1533 & v_1657;
assign v_21433 = v_1508 & v_21432;
assign v_21434 = v_1511 & v_1534;
assign v_21436 = v_1217 & v_21435;
assign v_21437 = v_1245 & v_1373;
assign v_21439 = v_1218 & v_21438;
assign v_21440 = v_1221 & v_1246;
assign v_21442 = v_936 & v_21441;
assign v_21443 = v_961 & v_1085;
assign v_21445 = v_937 & v_21444;
assign v_21446 = v_940 & v_962;
assign v_21448 = v_92 & v_21447;
assign v_21449 = v_591 & v_804;
assign v_21451 = v_94 & v_21450;
assign v_21452 = v_98 & v_593;
assign v_21455 = v_9601 & v_9796;
assign v_21456 = v_9630 & v_9664;
assign v_21458 = v_9307 & v_21457;
assign v_21459 = v_9335 & v_9506;
assign v_21461 = v_9308 & v_21460;
assign v_21462 = v_9336 & v_9374;
assign v_21464 = v_9026 & v_21463;
assign v_21465 = v_9051 & v_9218;
assign v_21467 = v_9027 & v_21466;
assign v_21468 = v_9052 & v_9086;
assign v_21470 = v_8729 & v_21469;
assign v_21471 = v_8761 & v_8936;
assign v_21473 = v_8730 & v_21472;
assign v_21474 = v_8762 & v_8804;
assign v_21476 = v_8447 & v_21475;
assign v_21477 = v_8473 & v_8640;
assign v_21479 = v_8448 & v_21478;
assign v_21480 = v_8474 & v_8508;
assign v_21482 = v_8157 & v_21481;
assign v_21483 = v_8185 & v_8356;
assign v_21485 = v_8158 & v_21484;
assign v_21486 = v_8186 & v_8224;
assign v_21488 = v_7876 & v_21487;
assign v_21489 = v_7901 & v_8068;
assign v_21491 = v_7877 & v_21490;
assign v_21492 = v_7902 & v_7936;
assign v_21494 = v_7571 & v_21493;
assign v_21495 = v_7607 & v_7786;
assign v_21497 = v_7572 & v_21496;
assign v_21498 = v_7608 & v_7654;
assign v_21500 = v_7288 & v_21499;
assign v_21501 = v_7315 & v_7482;
assign v_21503 = v_7289 & v_21502;
assign v_21504 = v_7316 & v_7350;
assign v_21506 = v_6997 & v_21505;
assign v_21507 = v_7025 & v_7196;
assign v_21509 = v_6998 & v_21508;
assign v_21510 = v_7026 & v_7064;
assign v_21512 = v_6716 & v_21511;
assign v_21513 = v_6741 & v_6908;
assign v_21515 = v_6717 & v_21514;
assign v_21516 = v_6742 & v_6776;
assign v_21518 = v_6419 & v_21517;
assign v_21519 = v_6451 & v_6626;
assign v_21521 = v_6420 & v_21520;
assign v_21522 = v_6452 & v_6494;
assign v_21524 = v_6137 & v_21523;
assign v_21525 = v_6163 & v_6330;
assign v_21527 = v_6138 & v_21526;
assign v_21528 = v_6164 & v_6198;
assign v_21530 = v_5847 & v_21529;
assign v_21531 = v_5875 & v_6046;
assign v_21533 = v_5848 & v_21532;
assign v_21534 = v_5876 & v_5914;
assign v_21536 = v_5566 & v_21535;
assign v_21537 = v_5591 & v_5758;
assign v_21539 = v_5567 & v_21538;
assign v_21540 = v_5592 & v_5626;
assign v_21542 = v_5253 & v_21541;
assign v_21543 = v_5293 & v_5476;
assign v_21545 = v_5254 & v_21544;
assign v_21546 = v_5294 & v_5344;
assign v_21548 = v_4969 & v_21547;
assign v_21549 = v_4997 & v_5164;
assign v_21551 = v_4970 & v_21550;
assign v_21552 = v_4998 & v_5032;
assign v_21554 = v_4677 & v_21553;
assign v_21555 = v_4705 & v_4876;
assign v_21557 = v_4678 & v_21556;
assign v_21558 = v_4706 & v_4744;
assign v_21560 = v_4396 & v_21559;
assign v_21561 = v_4421 & v_4588;
assign v_21563 = v_4397 & v_21562;
assign v_21564 = v_4422 & v_4456;
assign v_21566 = v_4099 & v_21565;
assign v_21567 = v_4131 & v_4306;
assign v_21569 = v_4100 & v_21568;
assign v_21570 = v_4132 & v_4174;
assign v_21572 = v_3817 & v_21571;
assign v_21573 = v_3843 & v_4010;
assign v_21575 = v_3818 & v_21574;
assign v_21576 = v_3844 & v_3878;
assign v_21578 = v_3527 & v_21577;
assign v_21579 = v_3555 & v_3726;
assign v_21581 = v_3528 & v_21580;
assign v_21582 = v_3556 & v_3594;
assign v_21584 = v_3246 & v_21583;
assign v_21585 = v_3271 & v_3438;
assign v_21587 = v_3247 & v_21586;
assign v_21588 = v_3272 & v_3306;
assign v_21590 = v_2941 & v_21589;
assign v_21591 = v_2977 & v_3156;
assign v_21593 = v_2942 & v_21592;
assign v_21594 = v_2978 & v_3024;
assign v_21596 = v_2658 & v_21595;
assign v_21597 = v_2685 & v_2852;
assign v_21599 = v_2659 & v_21598;
assign v_21600 = v_2686 & v_2720;
assign v_21602 = v_2367 & v_21601;
assign v_21603 = v_2395 & v_2566;
assign v_21605 = v_2368 & v_21604;
assign v_21606 = v_2396 & v_2434;
assign v_21608 = v_2086 & v_21607;
assign v_21609 = v_2111 & v_2278;
assign v_21611 = v_2087 & v_21610;
assign v_21612 = v_2112 & v_2146;
assign v_21614 = v_1789 & v_21613;
assign v_21615 = v_1821 & v_1996;
assign v_21617 = v_1790 & v_21616;
assign v_21618 = v_1822 & v_1864;
assign v_21620 = v_1507 & v_21619;
assign v_21621 = v_1533 & v_1700;
assign v_21623 = v_1508 & v_21622;
assign v_21624 = v_1534 & v_1568;
assign v_21626 = v_1217 & v_21625;
assign v_21627 = v_1245 & v_1416;
assign v_21629 = v_1218 & v_21628;
assign v_21630 = v_1246 & v_1284;
assign v_21632 = v_936 & v_21631;
assign v_21633 = v_961 & v_1128;
assign v_21635 = v_937 & v_21634;
assign v_21636 = v_962 & v_996;
assign v_21638 = v_92 & v_21637;
assign v_21639 = v_591 & v_850;
assign v_21641 = v_94 & v_21640;
assign v_21642 = v_593 & v_731;
assign v_21645 = v_9601 & v_9808;
assign v_21646 = v_9630 & v_9676;
assign v_21648 = v_9307 & v_21647;
assign v_21649 = v_9335 & v_9518;
assign v_21651 = v_9308 & v_21650;
assign v_21652 = v_9336 & v_9386;
assign v_21654 = v_9026 & v_21653;
assign v_21655 = v_9051 & v_9230;
assign v_21657 = v_9027 & v_21656;
assign v_21658 = v_9052 & v_9098;
assign v_21660 = v_8729 & v_21659;
assign v_21661 = v_8761 & v_8948;
assign v_21663 = v_8730 & v_21662;
assign v_21664 = v_8762 & v_8816;
assign v_21666 = v_8447 & v_21665;
assign v_21667 = v_8473 & v_8652;
assign v_21669 = v_8448 & v_21668;
assign v_21670 = v_8474 & v_8520;
assign v_21672 = v_8157 & v_21671;
assign v_21673 = v_8185 & v_8368;
assign v_21675 = v_8158 & v_21674;
assign v_21676 = v_8186 & v_8236;
assign v_21678 = v_7876 & v_21677;
assign v_21679 = v_7901 & v_8080;
assign v_21681 = v_7877 & v_21680;
assign v_21682 = v_7902 & v_7948;
assign v_21684 = v_7571 & v_21683;
assign v_21685 = v_7607 & v_7798;
assign v_21687 = v_7572 & v_21686;
assign v_21688 = v_7608 & v_7666;
assign v_21690 = v_7288 & v_21689;
assign v_21691 = v_7315 & v_7494;
assign v_21693 = v_7289 & v_21692;
assign v_21694 = v_7316 & v_7362;
assign v_21696 = v_6997 & v_21695;
assign v_21697 = v_7025 & v_7208;
assign v_21699 = v_6998 & v_21698;
assign v_21700 = v_7026 & v_7076;
assign v_21702 = v_6716 & v_21701;
assign v_21703 = v_6741 & v_6920;
assign v_21705 = v_6717 & v_21704;
assign v_21706 = v_6742 & v_6788;
assign v_21708 = v_6419 & v_21707;
assign v_21709 = v_6451 & v_6638;
assign v_21711 = v_6420 & v_21710;
assign v_21712 = v_6452 & v_6506;
assign v_21714 = v_6137 & v_21713;
assign v_21715 = v_6163 & v_6342;
assign v_21717 = v_6138 & v_21716;
assign v_21718 = v_6164 & v_6210;
assign v_21720 = v_5847 & v_21719;
assign v_21721 = v_5875 & v_6058;
assign v_21723 = v_5848 & v_21722;
assign v_21724 = v_5876 & v_5926;
assign v_21726 = v_5566 & v_21725;
assign v_21727 = v_5591 & v_5770;
assign v_21729 = v_5567 & v_21728;
assign v_21730 = v_5592 & v_5638;
assign v_21732 = v_5253 & v_21731;
assign v_21733 = v_5293 & v_5488;
assign v_21735 = v_5254 & v_21734;
assign v_21736 = v_5294 & v_5356;
assign v_21738 = v_4969 & v_21737;
assign v_21739 = v_4997 & v_5176;
assign v_21741 = v_4970 & v_21740;
assign v_21742 = v_4998 & v_5044;
assign v_21744 = v_4677 & v_21743;
assign v_21745 = v_4705 & v_4888;
assign v_21747 = v_4678 & v_21746;
assign v_21748 = v_4706 & v_4756;
assign v_21750 = v_4396 & v_21749;
assign v_21751 = v_4421 & v_4600;
assign v_21753 = v_4397 & v_21752;
assign v_21754 = v_4422 & v_4468;
assign v_21756 = v_4099 & v_21755;
assign v_21757 = v_4131 & v_4318;
assign v_21759 = v_4100 & v_21758;
assign v_21760 = v_4132 & v_4186;
assign v_21762 = v_3817 & v_21761;
assign v_21763 = v_3843 & v_4022;
assign v_21765 = v_3818 & v_21764;
assign v_21766 = v_3844 & v_3890;
assign v_21768 = v_3527 & v_21767;
assign v_21769 = v_3555 & v_3738;
assign v_21771 = v_3528 & v_21770;
assign v_21772 = v_3556 & v_3606;
assign v_21774 = v_3246 & v_21773;
assign v_21775 = v_3271 & v_3450;
assign v_21777 = v_3247 & v_21776;
assign v_21778 = v_3272 & v_3318;
assign v_21780 = v_2941 & v_21779;
assign v_21781 = v_2977 & v_3168;
assign v_21783 = v_2942 & v_21782;
assign v_21784 = v_2978 & v_3036;
assign v_21786 = v_2658 & v_21785;
assign v_21787 = v_2685 & v_2864;
assign v_21789 = v_2659 & v_21788;
assign v_21790 = v_2686 & v_2732;
assign v_21792 = v_2367 & v_21791;
assign v_21793 = v_2395 & v_2578;
assign v_21795 = v_2368 & v_21794;
assign v_21796 = v_2396 & v_2446;
assign v_21798 = v_2086 & v_21797;
assign v_21799 = v_2111 & v_2290;
assign v_21801 = v_2087 & v_21800;
assign v_21802 = v_2112 & v_2158;
assign v_21804 = v_1789 & v_21803;
assign v_21805 = v_1821 & v_2008;
assign v_21807 = v_1790 & v_21806;
assign v_21808 = v_1822 & v_1876;
assign v_21810 = v_1507 & v_21809;
assign v_21811 = v_1533 & v_1712;
assign v_21813 = v_1508 & v_21812;
assign v_21814 = v_1534 & v_1580;
assign v_21816 = v_1217 & v_21815;
assign v_21817 = v_1245 & v_1428;
assign v_21819 = v_1218 & v_21818;
assign v_21820 = v_1246 & v_1296;
assign v_21822 = v_936 & v_21821;
assign v_21823 = v_961 & v_1140;
assign v_21825 = v_937 & v_21824;
assign v_21826 = v_962 & v_1008;
assign v_21828 = v_92 & v_21827;
assign v_21829 = v_591 & v_862;
assign v_21831 = v_94 & v_21830;
assign v_21832 = v_593 & v_741;
assign v_21835 = v_9601 & v_9820;
assign v_21836 = v_9630 & v_9688;
assign v_21838 = v_9307 & v_21837;
assign v_21839 = v_9335 & v_9530;
assign v_21841 = v_9308 & v_21840;
assign v_21842 = v_9336 & v_9398;
assign v_21844 = v_9026 & v_21843;
assign v_21845 = v_9051 & v_9242;
assign v_21847 = v_9027 & v_21846;
assign v_21848 = v_9052 & v_9110;
assign v_21850 = v_8729 & v_21849;
assign v_21851 = v_8761 & v_8960;
assign v_21853 = v_8730 & v_21852;
assign v_21854 = v_8762 & v_8828;
assign v_21856 = v_8447 & v_21855;
assign v_21857 = v_8473 & v_8664;
assign v_21859 = v_8448 & v_21858;
assign v_21860 = v_8474 & v_8532;
assign v_21862 = v_8157 & v_21861;
assign v_21863 = v_8185 & v_8380;
assign v_21865 = v_8158 & v_21864;
assign v_21866 = v_8186 & v_8248;
assign v_21868 = v_7876 & v_21867;
assign v_21869 = v_7901 & v_8092;
assign v_21871 = v_7877 & v_21870;
assign v_21872 = v_7902 & v_7960;
assign v_21874 = v_7571 & v_21873;
assign v_21875 = v_7607 & v_7810;
assign v_21877 = v_7572 & v_21876;
assign v_21878 = v_7608 & v_7678;
assign v_21880 = v_7288 & v_21879;
assign v_21881 = v_7315 & v_7506;
assign v_21883 = v_7289 & v_21882;
assign v_21884 = v_7316 & v_7374;
assign v_21886 = v_6997 & v_21885;
assign v_21887 = v_7025 & v_7220;
assign v_21889 = v_6998 & v_21888;
assign v_21890 = v_7026 & v_7088;
assign v_21892 = v_6716 & v_21891;
assign v_21893 = v_6741 & v_6932;
assign v_21895 = v_6717 & v_21894;
assign v_21896 = v_6742 & v_6800;
assign v_21898 = v_6419 & v_21897;
assign v_21899 = v_6451 & v_6650;
assign v_21901 = v_6420 & v_21900;
assign v_21902 = v_6452 & v_6518;
assign v_21904 = v_6137 & v_21903;
assign v_21905 = v_6163 & v_6354;
assign v_21907 = v_6138 & v_21906;
assign v_21908 = v_6164 & v_6222;
assign v_21910 = v_5847 & v_21909;
assign v_21911 = v_5875 & v_6070;
assign v_21913 = v_5848 & v_21912;
assign v_21914 = v_5876 & v_5938;
assign v_21916 = v_5566 & v_21915;
assign v_21917 = v_5591 & v_5782;
assign v_21919 = v_5567 & v_21918;
assign v_21920 = v_5592 & v_5650;
assign v_21922 = v_5253 & v_21921;
assign v_21923 = v_5293 & v_5500;
assign v_21925 = v_5254 & v_21924;
assign v_21926 = v_5294 & v_5368;
assign v_21928 = v_4969 & v_21927;
assign v_21929 = v_4997 & v_5188;
assign v_21931 = v_4970 & v_21930;
assign v_21932 = v_4998 & v_5056;
assign v_21934 = v_4677 & v_21933;
assign v_21935 = v_4705 & v_4900;
assign v_21937 = v_4678 & v_21936;
assign v_21938 = v_4706 & v_4768;
assign v_21940 = v_4396 & v_21939;
assign v_21941 = v_4421 & v_4612;
assign v_21943 = v_4397 & v_21942;
assign v_21944 = v_4422 & v_4480;
assign v_21946 = v_4099 & v_21945;
assign v_21947 = v_4131 & v_4330;
assign v_21949 = v_4100 & v_21948;
assign v_21950 = v_4132 & v_4198;
assign v_21952 = v_3817 & v_21951;
assign v_21953 = v_3843 & v_4034;
assign v_21955 = v_3818 & v_21954;
assign v_21956 = v_3844 & v_3902;
assign v_21958 = v_3527 & v_21957;
assign v_21959 = v_3555 & v_3750;
assign v_21961 = v_3528 & v_21960;
assign v_21962 = v_3556 & v_3618;
assign v_21964 = v_3246 & v_21963;
assign v_21965 = v_3271 & v_3462;
assign v_21967 = v_3247 & v_21966;
assign v_21968 = v_3272 & v_3330;
assign v_21970 = v_2941 & v_21969;
assign v_21971 = v_2977 & v_3180;
assign v_21973 = v_2942 & v_21972;
assign v_21974 = v_2978 & v_3048;
assign v_21976 = v_2658 & v_21975;
assign v_21977 = v_2685 & v_2876;
assign v_21979 = v_2659 & v_21978;
assign v_21980 = v_2686 & v_2744;
assign v_21982 = v_2367 & v_21981;
assign v_21983 = v_2395 & v_2590;
assign v_21985 = v_2368 & v_21984;
assign v_21986 = v_2396 & v_2458;
assign v_21988 = v_2086 & v_21987;
assign v_21989 = v_2111 & v_2302;
assign v_21991 = v_2087 & v_21990;
assign v_21992 = v_2112 & v_2170;
assign v_21994 = v_1789 & v_21993;
assign v_21995 = v_1821 & v_2020;
assign v_21997 = v_1790 & v_21996;
assign v_21998 = v_1822 & v_1888;
assign v_22000 = v_1507 & v_21999;
assign v_22001 = v_1533 & v_1724;
assign v_22003 = v_1508 & v_22002;
assign v_22004 = v_1534 & v_1592;
assign v_22006 = v_1217 & v_22005;
assign v_22007 = v_1245 & v_1440;
assign v_22009 = v_1218 & v_22008;
assign v_22010 = v_1246 & v_1308;
assign v_22012 = v_936 & v_22011;
assign v_22013 = v_961 & v_1152;
assign v_22015 = v_937 & v_22014;
assign v_22016 = v_962 & v_1020;
assign v_22018 = v_92 & v_22017;
assign v_22019 = v_591 & v_874;
assign v_22021 = v_94 & v_22020;
assign v_22022 = v_593 & v_751;
assign v_22025 = v_9601 & v_9832;
assign v_22026 = v_9630 & v_9700;
assign v_22028 = v_9307 & v_22027;
assign v_22029 = v_9335 & v_9542;
assign v_22031 = v_9308 & v_22030;
assign v_22032 = v_9336 & v_9410;
assign v_22034 = v_9026 & v_22033;
assign v_22035 = v_9051 & v_9254;
assign v_22037 = v_9027 & v_22036;
assign v_22038 = v_9052 & v_9122;
assign v_22040 = v_8729 & v_22039;
assign v_22041 = v_8761 & v_8972;
assign v_22043 = v_8730 & v_22042;
assign v_22044 = v_8762 & v_8840;
assign v_22046 = v_8447 & v_22045;
assign v_22047 = v_8473 & v_8676;
assign v_22049 = v_8448 & v_22048;
assign v_22050 = v_8474 & v_8544;
assign v_22052 = v_8157 & v_22051;
assign v_22053 = v_8185 & v_8392;
assign v_22055 = v_8158 & v_22054;
assign v_22056 = v_8186 & v_8260;
assign v_22058 = v_7876 & v_22057;
assign v_22059 = v_7901 & v_8104;
assign v_22061 = v_7877 & v_22060;
assign v_22062 = v_7902 & v_7972;
assign v_22064 = v_7571 & v_22063;
assign v_22065 = v_7607 & v_7822;
assign v_22067 = v_7572 & v_22066;
assign v_22068 = v_7608 & v_7690;
assign v_22070 = v_7288 & v_22069;
assign v_22071 = v_7315 & v_7518;
assign v_22073 = v_7289 & v_22072;
assign v_22074 = v_7316 & v_7386;
assign v_22076 = v_6997 & v_22075;
assign v_22077 = v_7025 & v_7232;
assign v_22079 = v_6998 & v_22078;
assign v_22080 = v_7026 & v_7100;
assign v_22082 = v_6716 & v_22081;
assign v_22083 = v_6741 & v_6944;
assign v_22085 = v_6717 & v_22084;
assign v_22086 = v_6742 & v_6812;
assign v_22088 = v_6419 & v_22087;
assign v_22089 = v_6451 & v_6662;
assign v_22091 = v_6420 & v_22090;
assign v_22092 = v_6452 & v_6530;
assign v_22094 = v_6137 & v_22093;
assign v_22095 = v_6163 & v_6366;
assign v_22097 = v_6138 & v_22096;
assign v_22098 = v_6164 & v_6234;
assign v_22100 = v_5847 & v_22099;
assign v_22101 = v_5875 & v_6082;
assign v_22103 = v_5848 & v_22102;
assign v_22104 = v_5876 & v_5950;
assign v_22106 = v_5566 & v_22105;
assign v_22107 = v_5591 & v_5794;
assign v_22109 = v_5567 & v_22108;
assign v_22110 = v_5592 & v_5662;
assign v_22112 = v_5253 & v_22111;
assign v_22113 = v_5293 & v_5512;
assign v_22115 = v_5254 & v_22114;
assign v_22116 = v_5294 & v_5380;
assign v_22118 = v_4969 & v_22117;
assign v_22119 = v_4997 & v_5200;
assign v_22121 = v_4970 & v_22120;
assign v_22122 = v_4998 & v_5068;
assign v_22124 = v_4677 & v_22123;
assign v_22125 = v_4705 & v_4912;
assign v_22127 = v_4678 & v_22126;
assign v_22128 = v_4706 & v_4780;
assign v_22130 = v_4396 & v_22129;
assign v_22131 = v_4421 & v_4624;
assign v_22133 = v_4397 & v_22132;
assign v_22134 = v_4422 & v_4492;
assign v_22136 = v_4099 & v_22135;
assign v_22137 = v_4131 & v_4342;
assign v_22139 = v_4100 & v_22138;
assign v_22140 = v_4132 & v_4210;
assign v_22142 = v_3817 & v_22141;
assign v_22143 = v_3843 & v_4046;
assign v_22145 = v_3818 & v_22144;
assign v_22146 = v_3844 & v_3914;
assign v_22148 = v_3527 & v_22147;
assign v_22149 = v_3555 & v_3762;
assign v_22151 = v_3528 & v_22150;
assign v_22152 = v_3556 & v_3630;
assign v_22154 = v_3246 & v_22153;
assign v_22155 = v_3271 & v_3474;
assign v_22157 = v_3247 & v_22156;
assign v_22158 = v_3272 & v_3342;
assign v_22160 = v_2941 & v_22159;
assign v_22161 = v_2977 & v_3192;
assign v_22163 = v_2942 & v_22162;
assign v_22164 = v_2978 & v_3060;
assign v_22166 = v_2658 & v_22165;
assign v_22167 = v_2685 & v_2888;
assign v_22169 = v_2659 & v_22168;
assign v_22170 = v_2686 & v_2756;
assign v_22172 = v_2367 & v_22171;
assign v_22173 = v_2395 & v_2602;
assign v_22175 = v_2368 & v_22174;
assign v_22176 = v_2396 & v_2470;
assign v_22178 = v_2086 & v_22177;
assign v_22179 = v_2111 & v_2314;
assign v_22181 = v_2087 & v_22180;
assign v_22182 = v_2112 & v_2182;
assign v_22184 = v_1789 & v_22183;
assign v_22185 = v_1821 & v_2032;
assign v_22187 = v_1790 & v_22186;
assign v_22188 = v_1822 & v_1900;
assign v_22190 = v_1507 & v_22189;
assign v_22191 = v_1533 & v_1736;
assign v_22193 = v_1508 & v_22192;
assign v_22194 = v_1534 & v_1604;
assign v_22196 = v_1217 & v_22195;
assign v_22197 = v_1245 & v_1452;
assign v_22199 = v_1218 & v_22198;
assign v_22200 = v_1246 & v_1320;
assign v_22202 = v_936 & v_22201;
assign v_22203 = v_961 & v_1164;
assign v_22205 = v_937 & v_22204;
assign v_22206 = v_962 & v_1032;
assign v_22208 = v_92 & v_22207;
assign v_22209 = v_591 & v_886;
assign v_22211 = v_94 & v_22210;
assign v_22212 = v_593 & v_761;
assign v_22217 = v_22215 & v_22216;
assign v_22220 = v_22218 & v_22219;
assign v_22223 = v_22221 & v_22222;
assign v_22226 = v_22224 & v_22225;
assign v_22229 = v_22227 & v_22228;
assign v_22232 = v_22230 & v_22231;
assign v_22235 = v_22233 & v_22234;
assign v_22238 = v_22236 & v_22237;
assign v_22241 = v_22239 & v_22240;
assign v_22244 = v_22242 & v_22243;
assign v_22247 = v_22245 & v_22246;
assign v_22250 = v_22248 & v_22249;
assign v_22253 = v_22251 & v_22252;
assign v_22256 = v_22254 & v_22255;
assign v_22259 = v_22257 & v_22258;
assign v_22262 = v_22260 & v_22261;
assign v_22265 = v_22263 & v_22264;
assign v_22268 = v_22266 & v_22267;
assign v_22271 = v_22269 & v_22270;
assign v_22274 = v_22272 & v_22273;
assign v_22277 = v_22275 & v_22276;
assign v_22280 = v_22278 & v_22279;
assign v_22283 = v_22281 & v_22282;
assign v_22286 = v_22284 & v_22285;
assign v_22289 = v_22287 & v_22288;
assign v_22292 = v_22290 & v_22291;
assign v_22295 = v_22293 & v_22294;
assign v_22298 = v_22296 & v_22297;
assign v_22301 = v_22299 & v_22300;
assign v_22304 = v_22302 & v_22303;
assign v_22307 = v_22305 & v_22306;
assign v_22310 = v_22308 & v_22309;
assign v_22313 = v_22311 & v_22312;
assign v_22316 = v_22314 & v_22315;
assign v_22319 = v_22317 & v_22318;
assign v_22322 = v_22320 & v_22321;
assign v_22325 = v_22323 & v_22324;
assign v_22328 = v_22326 & v_22327;
assign v_22331 = v_22329 & v_22330;
assign v_22334 = v_22332 & v_22333;
assign v_22337 = v_22335 & v_22336;
assign v_22340 = v_22338 & v_22339;
assign v_22343 = v_22341 & v_22342;
assign v_22346 = v_22344 & v_22345;
assign v_22349 = v_22347 & v_22348;
assign v_22352 = v_22350 & v_22351;
assign v_22355 = v_22353 & v_22354;
assign v_22358 = v_22356 & v_22357;
assign v_22361 = v_22359 & v_22360;
assign v_22364 = v_22362 & v_22363;
assign v_22367 = v_22365 & v_22366;
assign v_22370 = v_22368 & v_22369;
assign v_22373 = v_22371 & v_22372;
assign v_22376 = v_22374 & v_22375;
assign v_22379 = v_22377 & v_22378;
assign v_22382 = v_22380 & v_22381;
assign v_22385 = v_22383 & v_22384;
assign v_22388 = v_22386 & v_22387;
assign v_22391 = v_22389 & v_22390;
assign v_22394 = v_22392 & v_22393;
assign v_22397 = v_22395 & v_22396;
assign v_22400 = v_22398 & v_22399;
assign v_22403 = v_22401 & v_22402;
assign v_22405 = v_9601 & ~v_9872;
assign v_22406 = v_9630 & ~v_9740;
assign v_22408 = v_9307 & v_22407;
assign v_22409 = v_9335 & ~v_9582;
assign v_22411 = v_9308 & v_22410;
assign v_22412 = v_9336 & ~v_9450;
assign v_22414 = v_9026 & v_22413;
assign v_22415 = v_9051 & ~v_9294;
assign v_22417 = v_9027 & v_22416;
assign v_22418 = v_9052 & ~v_9162;
assign v_22420 = v_8729 & v_22419;
assign v_22421 = v_8761 & ~v_9012;
assign v_22423 = v_8730 & v_22422;
assign v_22424 = v_8762 & ~v_8880;
assign v_22426 = v_8447 & v_22425;
assign v_22427 = v_8473 & ~v_8716;
assign v_22429 = v_8448 & v_22428;
assign v_22430 = v_8474 & ~v_8584;
assign v_22432 = v_8157 & v_22431;
assign v_22433 = v_8185 & v_8432;
assign v_22435 = v_8158 & v_22434;
assign v_22436 = v_8186 & v_8300;
assign v_22438 = v_7876 & v_22437;
assign v_22439 = v_7901 & v_8144;
assign v_22441 = v_7877 & v_22440;
assign v_22442 = v_7902 & ~v_8012;
assign v_22444 = v_7571 & v_22443;
assign v_22445 = v_7607 & ~v_7862;
assign v_22447 = v_7572 & v_22446;
assign v_22448 = v_7608 & ~v_7730;
assign v_22450 = v_7288 & v_22449;
assign v_22451 = v_7315 & ~v_7558;
assign v_22453 = v_7289 & v_22452;
assign v_22454 = v_7316 & ~v_7426;
assign v_22456 = v_6997 & v_22455;
assign v_22457 = v_7025 & v_7272;
assign v_22459 = v_6998 & v_22458;
assign v_22460 = v_7026 & ~v_7140;
assign v_22462 = v_6716 & v_22461;
assign v_22463 = v_6741 & v_6984;
assign v_22465 = v_6717 & v_22464;
assign v_22466 = v_6742 & v_6852;
assign v_22468 = v_6419 & v_22467;
assign v_22469 = v_6451 & v_6702;
assign v_22471 = v_6420 & v_22470;
assign v_22472 = v_6452 & ~v_6570;
assign v_22474 = v_6137 & v_22473;
assign v_22475 = v_6163 & ~v_6406;
assign v_22477 = v_6138 & v_22476;
assign v_22478 = v_6164 & v_6274;
assign v_22480 = v_5847 & v_22479;
assign v_22481 = v_5875 & v_6122;
assign v_22483 = v_5848 & v_22482;
assign v_22484 = v_5876 & v_5990;
assign v_22486 = v_5566 & v_22485;
assign v_22487 = v_5591 & v_5834;
assign v_22489 = v_5567 & v_22488;
assign v_22490 = v_5592 & v_5702;
assign v_22492 = v_5253 & v_22491;
assign v_22493 = v_5293 & v_5552;
assign v_22495 = v_5254 & v_22494;
assign v_22496 = v_5294 & ~v_5420;
assign v_22498 = v_4969 & v_22497;
assign v_22499 = v_4997 & ~v_5240;
assign v_22501 = v_4970 & v_22500;
assign v_22502 = v_4998 & v_5108;
assign v_22504 = v_4677 & v_22503;
assign v_22505 = v_4705 & v_4952;
assign v_22507 = v_4678 & v_22506;
assign v_22508 = v_4706 & v_4820;
assign v_22510 = v_4396 & v_22509;
assign v_22511 = v_4421 & v_4664;
assign v_22513 = v_4397 & v_22512;
assign v_22514 = v_4422 & v_4532;
assign v_22516 = v_4099 & v_22515;
assign v_22517 = v_4131 & v_4382;
assign v_22519 = v_4100 & v_22518;
assign v_22520 = v_4132 & ~v_4250;
assign v_22522 = v_3817 & v_22521;
assign v_22523 = v_3843 & ~v_4086;
assign v_22525 = v_3818 & v_22524;
assign v_22526 = v_3844 & ~v_3954;
assign v_22528 = v_3527 & v_22527;
assign v_22529 = v_3555 & ~v_3802;
assign v_22531 = v_3528 & v_22530;
assign v_22532 = v_3556 & ~v_3670;
assign v_22534 = v_3246 & v_22533;
assign v_22535 = v_3271 & v_3514;
assign v_22537 = v_3247 & v_22536;
assign v_22538 = v_3272 & ~v_3382;
assign v_22540 = v_2941 & v_22539;
assign v_22541 = v_2977 & v_3232;
assign v_22543 = v_2942 & v_22542;
assign v_22544 = v_2978 & ~v_3100;
assign v_22546 = v_2658 & v_22545;
assign v_22547 = v_2685 & ~v_2928;
assign v_22549 = v_2659 & v_22548;
assign v_22550 = v_2686 & ~v_2796;
assign v_22552 = v_2367 & v_22551;
assign v_22553 = v_2395 & ~v_2642;
assign v_22555 = v_2368 & v_22554;
assign v_22556 = v_2396 & ~v_2510;
assign v_22558 = v_2086 & v_22557;
assign v_22559 = v_2111 & v_2354;
assign v_22561 = v_2087 & v_22560;
assign v_22562 = v_2112 & v_2222;
assign v_22564 = v_1789 & v_22563;
assign v_22565 = v_1821 & v_2072;
assign v_22567 = v_1790 & v_22566;
assign v_22568 = v_1822 & ~v_1940;
assign v_22570 = v_1507 & v_22569;
assign v_22571 = v_1533 & ~v_1776;
assign v_22573 = v_1508 & v_22572;
assign v_22574 = v_1534 & ~v_1644;
assign v_22576 = v_1217 & v_22575;
assign v_22577 = v_1245 & ~v_1492;
assign v_22579 = v_1218 & v_22578;
assign v_22580 = v_1246 & ~v_1360;
assign v_22582 = v_936 & v_22581;
assign v_22583 = v_961 & ~v_1204;
assign v_22585 = v_937 & v_22584;
assign v_22586 = v_962 & ~v_1072;
assign v_22588 = v_92 & v_22587;
assign v_22589 = v_591 & ~v_922;
assign v_22591 = v_94 & v_22590;
assign v_22592 = v_593 & ~v_793;
assign v_22598 = v_96 & v_22597;
assign v_22599 = v_9618 & v_9844;
assign v_22600 = v_9646 & v_9712;
assign v_22602 = v_9473 & v_22601;
assign v_22603 = v_9488 & v_9554;
assign v_22605 = v_9329 & v_22604;
assign v_22606 = v_9356 & v_9422;
assign v_22608 = v_9185 & v_22607;
assign v_22609 = v_9200 & v_9266;
assign v_22611 = v_9044 & v_22610;
assign v_22612 = v_9068 & v_9134;
assign v_22614 = v_8903 & v_22613;
assign v_22615 = v_8918 & v_8984;
assign v_22617 = v_8755 & v_22616;
assign v_22618 = v_8786 & v_8852;
assign v_22620 = v_8607 & v_22619;
assign v_22621 = v_8622 & v_8688;
assign v_22623 = v_8465 & v_22622;
assign v_22624 = v_8490 & v_8556;
assign v_22626 = v_8323 & v_22625;
assign v_22627 = v_8338 & v_8404;
assign v_22629 = v_8179 & v_22628;
assign v_22630 = v_8206 & v_8272;
assign v_22632 = v_8035 & v_22631;
assign v_22633 = v_8050 & v_8116;
assign v_22635 = v_7894 & v_22634;
assign v_22636 = v_7918 & v_7984;
assign v_22638 = v_7753 & v_22637;
assign v_22639 = v_7768 & v_7834;
assign v_22641 = v_7601 & v_22640;
assign v_22642 = v_7636 & v_7702;
assign v_22644 = v_7449 & v_22643;
assign v_22645 = v_7464 & v_7530;
assign v_22647 = v_7306 & v_22646;
assign v_22648 = v_7332 & v_7398;
assign v_22650 = v_7163 & v_22649;
assign v_22651 = v_7178 & v_7244;
assign v_22653 = v_7019 & v_22652;
assign v_22654 = v_7046 & v_7112;
assign v_22656 = v_6875 & v_22655;
assign v_22657 = v_6890 & v_6956;
assign v_22659 = v_6734 & v_22658;
assign v_22660 = v_6758 & ~v_6824;
assign v_22662 = v_6593 & v_22661;
assign v_22663 = v_6608 & v_6674;
assign v_22665 = v_6445 & v_22664;
assign v_22666 = v_6476 & v_6542;
assign v_22668 = v_6297 & v_22667;
assign v_22669 = v_6312 & v_6378;
assign v_22671 = v_6155 & v_22670;
assign v_22672 = v_6180 & v_6246;
assign v_22674 = v_6013 & v_22673;
assign v_22675 = v_6028 & ~v_6094;
assign v_22677 = v_5869 & v_22676;
assign v_22678 = v_5896 & v_5962;
assign v_22680 = v_5725 & v_22679;
assign v_22681 = v_5740 & ~v_5806;
assign v_22683 = v_5584 & v_22682;
assign v_22684 = v_5608 & v_5674;
assign v_22686 = v_5443 & v_22685;
assign v_22687 = v_5458 & v_5524;
assign v_22689 = v_5287 & v_22688;
assign v_22690 = v_5326 & v_5392;
assign v_22692 = v_5131 & v_22691;
assign v_22693 = v_5146 & v_5212;
assign v_22695 = v_4987 & v_22694;
assign v_22696 = v_5014 & v_5080;
assign v_22698 = v_4843 & v_22697;
assign v_22699 = v_4858 & v_4924;
assign v_22701 = v_4699 & v_22700;
assign v_22702 = v_4726 & v_4792;
assign v_22704 = v_4555 & v_22703;
assign v_22705 = v_4570 & v_4636;
assign v_22707 = v_4414 & v_22706;
assign v_22708 = v_4438 & v_4504;
assign v_22710 = v_4273 & v_22709;
assign v_22711 = v_4288 & v_4354;
assign v_22713 = v_4125 & v_22712;
assign v_22714 = v_4156 & v_4222;
assign v_22716 = v_3977 & v_22715;
assign v_22717 = v_3992 & v_4058;
assign v_22719 = v_3835 & v_22718;
assign v_22720 = v_3860 & v_3926;
assign v_22722 = v_3693 & v_22721;
assign v_22723 = v_3708 & v_3774;
assign v_22725 = v_3549 & v_22724;
assign v_22726 = v_3576 & v_3642;
assign v_22728 = v_3405 & v_22727;
assign v_22729 = v_3420 & v_3486;
assign v_22731 = v_3264 & v_22730;
assign v_22732 = v_3288 & v_3354;
assign v_22734 = v_3123 & v_22733;
assign v_22735 = v_3138 & ~v_3204;
assign v_22737 = v_2971 & v_22736;
assign v_22738 = v_3006 & v_3072;
assign v_22740 = v_2819 & v_22739;
assign v_22741 = v_2834 & v_2900;
assign v_22743 = v_2676 & v_22742;
assign v_22744 = v_2702 & v_2768;
assign v_22746 = v_2533 & v_22745;
assign v_22747 = v_2548 & v_2614;
assign v_22749 = v_2389 & v_22748;
assign v_22750 = v_2416 & v_2482;
assign v_22752 = v_2245 & v_22751;
assign v_22753 = v_2260 & v_2326;
assign v_22755 = v_2104 & v_22754;
assign v_22756 = v_2128 & v_2194;
assign v_22758 = v_1963 & v_22757;
assign v_22759 = v_1978 & v_2044;
assign v_22761 = v_1815 & v_22760;
assign v_22762 = v_1846 & v_1912;
assign v_22764 = v_1667 & v_22763;
assign v_22765 = v_1682 & v_1748;
assign v_22767 = v_1525 & v_22766;
assign v_22768 = v_1550 & v_1616;
assign v_22770 = v_1383 & v_22769;
assign v_22771 = v_1398 & v_1464;
assign v_22773 = v_1239 & v_22772;
assign v_22774 = v_1266 & v_1332;
assign v_22776 = v_1095 & v_22775;
assign v_22777 = v_1110 & v_1176;
assign v_22779 = v_954 & v_22778;
assign v_22780 = v_978 & v_1044;
assign v_22782 = v_816 & v_22781;
assign v_22783 = v_832 & v_898;
assign v_22785 = v_561 & v_22784;
assign v_22786 = v_715 & v_771;
assign v_22792 = v_10200 & v_22791;
assign v_22793 = v_9611 & v_9844;
assign v_22794 = v_9639 & v_9712;
assign v_22796 = v_9468 & v_22795;
assign v_22797 = v_9483 & v_9554;
assign v_22799 = v_9320 & v_22798;
assign v_22800 = v_9347 & v_9422;
assign v_22802 = v_9180 & v_22801;
assign v_22803 = v_9195 & v_9266;
assign v_22805 = v_9037 & v_22804;
assign v_22806 = v_9061 & v_9134;
assign v_22808 = v_8898 & v_22807;
assign v_22809 = v_8913 & v_8984;
assign v_22811 = v_8744 & v_22810;
assign v_22812 = v_8775 & v_8852;
assign v_22814 = v_8602 & v_22813;
assign v_22815 = v_8617 & v_8688;
assign v_22817 = v_8458 & v_22816;
assign v_22818 = v_8483 & v_8556;
assign v_22820 = v_8318 & v_22819;
assign v_22821 = v_8333 & v_8404;
assign v_22823 = v_8170 & v_22822;
assign v_22824 = v_8197 & v_8272;
assign v_22826 = v_8030 & v_22825;
assign v_22827 = v_8045 & v_8116;
assign v_22829 = v_7887 & v_22828;
assign v_22830 = v_7911 & v_7984;
assign v_22832 = v_7748 & v_22831;
assign v_22833 = v_7763 & v_7834;
assign v_22835 = v_7588 & v_22834;
assign v_22836 = v_7623 & v_7702;
assign v_22838 = v_7444 & v_22837;
assign v_22839 = v_7459 & v_7530;
assign v_22841 = v_7299 & v_22840;
assign v_22842 = v_7325 & v_7398;
assign v_22844 = v_7158 & v_22843;
assign v_22845 = v_7173 & v_7244;
assign v_22847 = v_7010 & v_22846;
assign v_22848 = v_7037 & v_7112;
assign v_22850 = v_6870 & v_22849;
assign v_22851 = v_6885 & v_6956;
assign v_22853 = v_6727 & v_22852;
assign v_22854 = v_6751 & ~v_6824;
assign v_22856 = v_6588 & v_22855;
assign v_22857 = v_6603 & v_6674;
assign v_22859 = v_6434 & v_22858;
assign v_22860 = v_6465 & v_6542;
assign v_22862 = v_6292 & v_22861;
assign v_22863 = v_6307 & v_6378;
assign v_22865 = v_6148 & v_22864;
assign v_22866 = v_6173 & v_6246;
assign v_22868 = v_6008 & v_22867;
assign v_22869 = v_6023 & ~v_6094;
assign v_22871 = v_5860 & v_22870;
assign v_22872 = v_5887 & v_5962;
assign v_22874 = v_5720 & v_22873;
assign v_22875 = v_5735 & ~v_5806;
assign v_22877 = v_5577 & v_22876;
assign v_22878 = v_5601 & v_5674;
assign v_22880 = v_5438 & v_22879;
assign v_22881 = v_5453 & v_5524;
assign v_22883 = v_5272 & v_22882;
assign v_22884 = v_5311 & v_5392;
assign v_22886 = v_5126 & v_22885;
assign v_22887 = v_5141 & v_5212;
assign v_22889 = v_4980 & v_22888;
assign v_22890 = v_5007 & v_5080;
assign v_22892 = v_4838 & v_22891;
assign v_22893 = v_4853 & v_4924;
assign v_22895 = v_4690 & v_22894;
assign v_22896 = v_4717 & v_4792;
assign v_22898 = v_4550 & v_22897;
assign v_22899 = v_4565 & v_4636;
assign v_22901 = v_4407 & v_22900;
assign v_22902 = v_4431 & v_4504;
assign v_22904 = v_4268 & v_22903;
assign v_22905 = v_4283 & v_4354;
assign v_22907 = v_4114 & v_22906;
assign v_22908 = v_4145 & v_4222;
assign v_22910 = v_3972 & v_22909;
assign v_22911 = v_3987 & v_4058;
assign v_22913 = v_3828 & v_22912;
assign v_22914 = v_3853 & v_3926;
assign v_22916 = v_3688 & v_22915;
assign v_22917 = v_3703 & v_3774;
assign v_22919 = v_3540 & v_22918;
assign v_22920 = v_3567 & v_3642;
assign v_22922 = v_3400 & v_22921;
assign v_22923 = v_3415 & v_3486;
assign v_22925 = v_3257 & v_22924;
assign v_22926 = v_3281 & v_3354;
assign v_22928 = v_3118 & v_22927;
assign v_22929 = v_3133 & ~v_3204;
assign v_22931 = v_2958 & v_22930;
assign v_22932 = v_2993 & v_3072;
assign v_22934 = v_2814 & v_22933;
assign v_22935 = v_2829 & v_2900;
assign v_22937 = v_2669 & v_22936;
assign v_22938 = v_2695 & v_2768;
assign v_22940 = v_2528 & v_22939;
assign v_22941 = v_2543 & v_2614;
assign v_22943 = v_2380 & v_22942;
assign v_22944 = v_2407 & v_2482;
assign v_22946 = v_2240 & v_22945;
assign v_22947 = v_2255 & v_2326;
assign v_22949 = v_2097 & v_22948;
assign v_22950 = v_2121 & v_2194;
assign v_22952 = v_1958 & v_22951;
assign v_22953 = v_1973 & v_2044;
assign v_22955 = v_1804 & v_22954;
assign v_22956 = v_1835 & v_1912;
assign v_22958 = v_1662 & v_22957;
assign v_22959 = v_1677 & v_1748;
assign v_22961 = v_1518 & v_22960;
assign v_22962 = v_1543 & v_1616;
assign v_22964 = v_1378 & v_22963;
assign v_22965 = v_1393 & v_1464;
assign v_22967 = v_1230 & v_22966;
assign v_22968 = v_1257 & v_1332;
assign v_22970 = v_1090 & v_22969;
assign v_22971 = v_1105 & v_1176;
assign v_22973 = v_947 & v_22972;
assign v_22974 = v_971 & v_1044;
assign v_22976 = v_811 & v_22975;
assign v_22977 = v_827 & v_898;
assign v_22979 = v_359 & v_22978;
assign v_22980 = v_658 & v_771;
assign v_22986 = v_10196 & v_22985;
assign v_22987 = v_9308 & v_9844;
assign v_22988 = v_9336 & v_9712;
assign v_22990 = v_9026 & v_22989;
assign v_22991 = v_9051 & v_9554;
assign v_22993 = v_9027 & v_22992;
assign v_22994 = v_9052 & v_9422;
assign v_22996 = v_8729 & v_22995;
assign v_22997 = v_8761 & v_9266;
assign v_22999 = v_8730 & v_22998;
assign v_23000 = v_8762 & v_9134;
assign v_23002 = v_8447 & v_23001;
assign v_23003 = v_8473 & v_8984;
assign v_23005 = v_8448 & v_23004;
assign v_23006 = v_8474 & v_8852;
assign v_23008 = v_8157 & v_23007;
assign v_23009 = v_8185 & v_8688;
assign v_23011 = v_8158 & v_23010;
assign v_23012 = v_8186 & v_8556;
assign v_23014 = v_7876 & v_23013;
assign v_23015 = v_7901 & v_8404;
assign v_23017 = v_7877 & v_23016;
assign v_23018 = v_7902 & v_8272;
assign v_23020 = v_7571 & v_23019;
assign v_23021 = v_7607 & v_8116;
assign v_23023 = v_7572 & v_23022;
assign v_23024 = v_7608 & v_7984;
assign v_23026 = v_7288 & v_23025;
assign v_23027 = v_7315 & v_7834;
assign v_23029 = v_7289 & v_23028;
assign v_23030 = v_7316 & v_7702;
assign v_23032 = v_6997 & v_23031;
assign v_23033 = v_7025 & v_7530;
assign v_23035 = v_6998 & v_23034;
assign v_23036 = v_7026 & v_7398;
assign v_23038 = v_6716 & v_23037;
assign v_23039 = v_6741 & v_7244;
assign v_23041 = v_6717 & v_23040;
assign v_23042 = v_6742 & v_7112;
assign v_23044 = v_6419 & v_23043;
assign v_23045 = v_6451 & v_6956;
assign v_23047 = v_6420 & v_23046;
assign v_23048 = v_6452 & ~v_6824;
assign v_23050 = v_6137 & v_23049;
assign v_23051 = v_6163 & v_6674;
assign v_23053 = v_6138 & v_23052;
assign v_23054 = v_6164 & v_6542;
assign v_23056 = v_5847 & v_23055;
assign v_23057 = v_5875 & v_6378;
assign v_23059 = v_5848 & v_23058;
assign v_23060 = v_5876 & v_6246;
assign v_23062 = v_5566 & v_23061;
assign v_23063 = v_5591 & ~v_6094;
assign v_23065 = v_5567 & v_23064;
assign v_23066 = v_5592 & v_5962;
assign v_23068 = v_5253 & v_23067;
assign v_23069 = v_5293 & ~v_5806;
assign v_23071 = v_5254 & v_23070;
assign v_23072 = v_5294 & v_5674;
assign v_23074 = v_4969 & v_23073;
assign v_23075 = v_4997 & v_5524;
assign v_23077 = v_4970 & v_23076;
assign v_23078 = v_4998 & v_5392;
assign v_23080 = v_4677 & v_23079;
assign v_23081 = v_4705 & v_5212;
assign v_23083 = v_4678 & v_23082;
assign v_23084 = v_4706 & v_5080;
assign v_23086 = v_4396 & v_23085;
assign v_23087 = v_4421 & v_4924;
assign v_23089 = v_4397 & v_23088;
assign v_23090 = v_4422 & v_4792;
assign v_23092 = v_4099 & v_23091;
assign v_23093 = v_4131 & v_4636;
assign v_23095 = v_4100 & v_23094;
assign v_23096 = v_4132 & v_4504;
assign v_23098 = v_3817 & v_23097;
assign v_23099 = v_3843 & v_4354;
assign v_23101 = v_3818 & v_23100;
assign v_23102 = v_3844 & v_4222;
assign v_23104 = v_3527 & v_23103;
assign v_23105 = v_3555 & v_4058;
assign v_23107 = v_3528 & v_23106;
assign v_23108 = v_3556 & v_3926;
assign v_23110 = v_3246 & v_23109;
assign v_23111 = v_3271 & v_3774;
assign v_23113 = v_3247 & v_23112;
assign v_23114 = v_3272 & v_3642;
assign v_23116 = v_2941 & v_23115;
assign v_23117 = v_2977 & v_3486;
assign v_23119 = v_2942 & v_23118;
assign v_23120 = v_2978 & v_3354;
assign v_23122 = v_2658 & v_23121;
assign v_23123 = v_2685 & ~v_3204;
assign v_23125 = v_2659 & v_23124;
assign v_23126 = v_2686 & v_3072;
assign v_23128 = v_2367 & v_23127;
assign v_23129 = v_2395 & v_2900;
assign v_23131 = v_2368 & v_23130;
assign v_23132 = v_2396 & v_2768;
assign v_23134 = v_2086 & v_23133;
assign v_23135 = v_2111 & v_2614;
assign v_23137 = v_2087 & v_23136;
assign v_23138 = v_2112 & v_2482;
assign v_23140 = v_1789 & v_23139;
assign v_23141 = v_1821 & v_2326;
assign v_23143 = v_1790 & v_23142;
assign v_23144 = v_1822 & v_2194;
assign v_23146 = v_1507 & v_23145;
assign v_23147 = v_1533 & v_2044;
assign v_23149 = v_1508 & v_23148;
assign v_23150 = v_1534 & v_1912;
assign v_23152 = v_1217 & v_23151;
assign v_23153 = v_1245 & v_1748;
assign v_23155 = v_1218 & v_23154;
assign v_23156 = v_1246 & v_1616;
assign v_23158 = v_936 & v_23157;
assign v_23159 = v_961 & v_1464;
assign v_23161 = v_937 & v_23160;
assign v_23162 = v_962 & v_1332;
assign v_23164 = v_92 & v_23163;
assign v_23165 = v_591 & v_1176;
assign v_23167 = v_94 & v_23166;
assign v_23168 = v_593 & v_1044;
assign v_23170 = v_806 & v_23169;
assign v_23171 = v_823 & v_898;
assign v_23177 = v_9903 & v_23176;
assign v_23178 = v_9601 & v_9844;
assign v_23179 = v_9630 & v_9712;
assign v_23181 = v_9307 & v_23180;
assign v_23182 = v_9335 & v_9554;
assign v_23184 = v_9308 & v_23183;
assign v_23185 = v_9336 & v_9422;
assign v_23187 = v_9026 & v_23186;
assign v_23188 = v_9051 & v_9266;
assign v_23190 = v_9027 & v_23189;
assign v_23191 = v_9052 & v_9134;
assign v_23193 = v_8729 & v_23192;
assign v_23194 = v_8761 & v_8984;
assign v_23196 = v_8730 & v_23195;
assign v_23197 = v_8762 & v_8852;
assign v_23199 = v_8447 & v_23198;
assign v_23200 = v_8473 & v_8688;
assign v_23202 = v_8448 & v_23201;
assign v_23203 = v_8474 & v_8556;
assign v_23205 = v_8157 & v_23204;
assign v_23206 = v_8185 & v_8404;
assign v_23208 = v_8158 & v_23207;
assign v_23209 = v_8186 & v_8272;
assign v_23211 = v_7876 & v_23210;
assign v_23212 = v_7901 & v_8116;
assign v_23214 = v_7877 & v_23213;
assign v_23215 = v_7902 & v_7984;
assign v_23217 = v_7571 & v_23216;
assign v_23218 = v_7607 & v_7834;
assign v_23220 = v_7572 & v_23219;
assign v_23221 = v_7608 & v_7702;
assign v_23223 = v_7288 & v_23222;
assign v_23224 = v_7315 & v_7530;
assign v_23226 = v_7289 & v_23225;
assign v_23227 = v_7316 & v_7398;
assign v_23229 = v_6997 & v_23228;
assign v_23230 = v_7025 & v_7244;
assign v_23232 = v_6998 & v_23231;
assign v_23233 = v_7026 & v_7112;
assign v_23235 = v_6716 & v_23234;
assign v_23236 = v_6741 & v_6956;
assign v_23238 = v_6717 & v_23237;
assign v_23239 = v_6742 & ~v_6824;
assign v_23241 = v_6419 & v_23240;
assign v_23242 = v_6451 & v_6674;
assign v_23244 = v_6420 & v_23243;
assign v_23245 = v_6452 & v_6542;
assign v_23247 = v_6137 & v_23246;
assign v_23248 = v_6163 & v_6378;
assign v_23250 = v_6138 & v_23249;
assign v_23251 = v_6164 & v_6246;
assign v_23253 = v_5847 & v_23252;
assign v_23254 = v_5875 & ~v_6094;
assign v_23256 = v_5848 & v_23255;
assign v_23257 = v_5876 & v_5962;
assign v_23259 = v_5566 & v_23258;
assign v_23260 = v_5591 & ~v_5806;
assign v_23262 = v_5567 & v_23261;
assign v_23263 = v_5592 & v_5674;
assign v_23265 = v_5253 & v_23264;
assign v_23266 = v_5293 & v_5524;
assign v_23268 = v_5254 & v_23267;
assign v_23269 = v_5294 & v_5392;
assign v_23271 = v_4969 & v_23270;
assign v_23272 = v_4997 & v_5212;
assign v_23274 = v_4970 & v_23273;
assign v_23275 = v_4998 & v_5080;
assign v_23277 = v_4677 & v_23276;
assign v_23278 = v_4705 & v_4924;
assign v_23280 = v_4678 & v_23279;
assign v_23281 = v_4706 & v_4792;
assign v_23283 = v_4396 & v_23282;
assign v_23284 = v_4421 & v_4636;
assign v_23286 = v_4397 & v_23285;
assign v_23287 = v_4422 & v_4504;
assign v_23289 = v_4099 & v_23288;
assign v_23290 = v_4131 & v_4354;
assign v_23292 = v_4100 & v_23291;
assign v_23293 = v_4132 & v_4222;
assign v_23295 = v_3817 & v_23294;
assign v_23296 = v_3843 & v_4058;
assign v_23298 = v_3818 & v_23297;
assign v_23299 = v_3844 & v_3926;
assign v_23301 = v_3527 & v_23300;
assign v_23302 = v_3555 & v_3774;
assign v_23304 = v_3528 & v_23303;
assign v_23305 = v_3556 & v_3642;
assign v_23307 = v_3246 & v_23306;
assign v_23308 = v_3271 & v_3486;
assign v_23310 = v_3247 & v_23309;
assign v_23311 = v_3272 & v_3354;
assign v_23313 = v_2941 & v_23312;
assign v_23314 = v_2977 & ~v_3204;
assign v_23316 = v_2942 & v_23315;
assign v_23317 = v_2978 & v_3072;
assign v_23319 = v_2658 & v_23318;
assign v_23320 = v_2685 & v_2900;
assign v_23322 = v_2659 & v_23321;
assign v_23323 = v_2686 & v_2768;
assign v_23325 = v_2367 & v_23324;
assign v_23326 = v_2395 & v_2614;
assign v_23328 = v_2368 & v_23327;
assign v_23329 = v_2396 & v_2482;
assign v_23331 = v_2086 & v_23330;
assign v_23332 = v_2111 & v_2326;
assign v_23334 = v_2087 & v_23333;
assign v_23335 = v_2112 & v_2194;
assign v_23337 = v_1789 & v_23336;
assign v_23338 = v_1821 & v_2044;
assign v_23340 = v_1790 & v_23339;
assign v_23341 = v_1822 & v_1912;
assign v_23343 = v_1507 & v_23342;
assign v_23344 = v_1533 & v_1748;
assign v_23346 = v_1508 & v_23345;
assign v_23347 = v_1534 & v_1616;
assign v_23349 = v_1217 & v_23348;
assign v_23350 = v_1245 & v_1464;
assign v_23352 = v_1218 & v_23351;
assign v_23353 = v_1246 & v_1332;
assign v_23355 = v_936 & v_23354;
assign v_23356 = v_961 & v_1176;
assign v_23358 = v_937 & v_23357;
assign v_23359 = v_962 & v_1044;
assign v_23361 = v_92 & v_23360;
assign v_23362 = v_591 & v_898;
assign v_23364 = v_94 & v_23363;
assign v_23365 = v_593 & v_771;
assign v_23371 = v_9884 & v_23370;
assign v_23405 = v_10415 & v_23404;
assign v_23427 = v_23425 & v_23426;
assign v_23428 = v_23424 & v_23427;
assign v_23429 = v_23423 & v_23428;
assign v_23430 = v_23422 & v_23429;
assign v_23431 = v_23421 & v_23430;
assign v_23432 = v_23420 & v_23431;
assign v_23433 = v_23419 & v_23432;
assign v_23437 = v_23435 & v_23436;
assign v_23440 = v_23438 & v_23439;
assign v_23443 = v_23441 & v_23442;
assign v_23446 = v_23444 & v_23445;
assign v_23449 = v_23447 & v_23448;
assign v_23452 = v_23450 & v_23451;
assign v_23455 = v_23453 & v_23454;
assign v_23458 = v_23456 & v_23457;
assign v_23461 = v_23459 & v_23460;
assign v_23464 = v_23462 & v_23463;
assign v_23467 = v_23465 & v_23466;
assign v_23470 = v_23468 & v_23469;
assign v_23473 = v_23471 & v_23472;
assign v_23476 = v_23474 & v_23475;
assign v_23479 = v_23477 & v_23478;
assign v_23482 = v_23480 & v_23481;
assign v_23485 = v_23483 & v_23484;
assign v_23488 = v_23486 & v_23487;
assign v_23491 = v_23489 & v_23490;
assign v_23494 = v_23492 & v_23493;
assign v_23497 = v_23495 & v_23496;
assign v_23500 = v_23498 & v_23499;
assign v_23503 = v_23501 & v_23502;
assign v_23506 = v_23504 & v_23505;
assign v_23509 = v_23507 & v_23508;
assign v_23512 = v_23510 & v_23511;
assign v_23515 = v_23513 & v_23514;
assign v_23518 = v_23516 & v_23517;
assign v_23521 = v_23519 & v_23520;
assign v_23524 = v_23522 & v_23523;
assign v_23527 = v_23525 & v_23526;
assign v_23530 = v_23528 & v_23529;
assign v_23533 = v_23531 & v_23532;
assign v_23536 = v_23534 & v_23535;
assign v_23539 = v_23537 & v_23538;
assign v_23542 = v_23540 & v_23541;
assign v_23545 = v_23543 & v_23544;
assign v_23548 = v_23546 & v_23547;
assign v_23551 = v_23549 & v_23550;
assign v_23554 = v_23552 & v_23553;
assign v_23557 = v_23555 & v_23556;
assign v_23560 = v_23558 & v_23559;
assign v_23563 = v_23561 & v_23562;
assign v_23566 = v_23564 & v_23565;
assign v_23569 = v_23567 & v_23568;
assign v_23572 = v_23570 & v_23571;
assign v_23575 = v_23573 & v_23574;
assign v_23578 = v_23576 & v_23577;
assign v_23581 = v_23579 & v_23580;
assign v_23584 = v_23582 & v_23583;
assign v_23587 = v_23585 & v_23586;
assign v_23590 = v_23588 & v_23589;
assign v_23593 = v_23591 & v_23592;
assign v_23596 = v_23594 & v_23595;
assign v_23599 = v_23597 & v_23598;
assign v_23602 = v_23600 & v_23601;
assign v_23605 = v_23603 & v_23604;
assign v_23608 = v_23606 & v_23607;
assign v_23611 = v_23609 & v_23610;
assign v_23614 = v_23612 & v_23613;
assign v_23617 = v_23615 & v_23616;
assign v_23620 = v_23618 & v_23619;
assign v_23623 = v_23621 & v_23622;
assign v_23626 = v_23624 & v_23625;
assign v_23629 = v_23627 & v_23628;
assign v_23632 = v_23630 & v_23631;
assign v_23635 = v_23633 & v_23634;
assign v_23638 = v_23636 & v_23637;
assign v_23641 = v_23639 & v_23640;
assign v_23644 = v_23642 & v_23643;
assign v_23647 = v_23645 & v_23646;
assign v_23650 = v_23648 & v_23649;
assign v_23653 = v_23651 & v_23652;
assign v_23656 = v_23654 & v_23655;
assign v_23659 = v_23657 & v_23658;
assign v_23662 = v_23660 & v_23661;
assign v_23665 = v_23663 & v_23664;
assign v_23668 = v_23666 & v_23667;
assign v_23671 = v_23669 & v_23670;
assign v_23674 = v_23672 & v_23673;
assign v_23677 = v_23675 & v_23676;
assign v_23680 = v_23678 & v_23679;
assign v_23683 = v_23681 & v_23682;
assign v_23686 = v_23684 & v_23685;
assign v_23689 = v_23687 & v_23688;
assign v_23692 = v_23690 & v_23691;
assign v_23695 = v_23693 & v_23694;
assign v_23698 = v_23696 & v_23697;
assign v_23701 = v_23699 & v_23700;
assign v_23704 = v_23702 & v_23703;
assign v_23707 = v_23705 & v_23706;
assign v_23710 = v_23708 & v_23709;
assign v_23713 = v_23711 & v_23712;
assign v_23716 = v_23714 & v_23715;
assign v_23719 = v_23717 & v_23718;
assign v_23722 = v_23720 & v_23721;
assign v_23725 = v_23723 & v_23724;
assign v_23728 = v_23726 & v_23727;
assign v_23731 = v_23729 & v_23730;
assign v_23734 = v_23732 & v_23733;
assign v_23737 = v_23735 & v_23736;
assign v_23740 = v_23738 & v_23739;
assign v_23743 = v_23741 & v_23742;
assign v_23746 = v_23744 & v_23745;
assign v_23749 = v_23747 & v_23748;
assign v_23752 = v_23750 & v_23751;
assign v_23755 = v_23753 & v_23754;
assign v_23758 = v_23756 & v_23757;
assign v_23761 = v_23759 & v_23760;
assign v_23764 = v_23762 & v_23763;
assign v_23767 = v_23765 & v_23766;
assign v_23770 = v_23768 & v_23769;
assign v_23773 = v_23771 & v_23772;
assign v_23776 = v_23774 & v_23775;
assign v_23779 = v_23777 & v_23778;
assign v_23782 = v_23780 & v_23781;
assign v_23785 = v_23783 & v_23784;
assign v_23788 = v_23786 & v_23787;
assign v_23791 = v_23789 & v_23790;
assign v_23794 = v_23792 & v_23793;
assign v_23797 = v_23795 & v_23796;
assign v_23800 = v_23798 & v_23799;
assign v_23803 = v_23801 & v_23802;
assign v_23806 = v_23804 & v_23805;
assign v_23809 = v_23807 & v_23808;
assign v_23812 = v_23810 & v_23811;
assign v_23813 = v_23623 & v_23812;
assign v_23816 = v_23814 & v_23815;
assign v_23819 = v_23817 & v_23818;
assign v_23822 = v_23820 & v_23821;
assign v_23825 = v_23823 & v_23824;
assign v_23828 = v_23826 & v_23827;
assign v_23831 = v_23829 & v_23830;
assign v_23834 = v_23832 & v_23833;
assign v_23837 = v_23835 & v_23836;
assign v_23840 = v_23838 & v_23839;
assign v_23843 = v_23841 & v_23842;
assign v_23846 = v_23844 & v_23845;
assign v_23849 = v_23847 & v_23848;
assign v_23852 = v_23850 & v_23851;
assign v_23855 = v_23853 & v_23854;
assign v_23858 = v_23856 & v_23857;
assign v_23861 = v_23859 & v_23860;
assign v_23864 = v_23862 & v_23863;
assign v_23867 = v_23865 & v_23866;
assign v_23870 = v_23868 & v_23869;
assign v_23873 = v_23871 & v_23872;
assign v_23876 = v_23874 & v_23875;
assign v_23879 = v_23877 & v_23878;
assign v_23882 = v_23880 & v_23881;
assign v_23885 = v_23883 & v_23884;
assign v_23888 = v_23886 & v_23887;
assign v_23891 = v_23889 & v_23890;
assign v_23894 = v_23892 & v_23893;
assign v_23897 = v_23895 & v_23896;
assign v_23900 = v_23898 & v_23899;
assign v_23903 = v_23901 & v_23902;
assign v_23906 = v_23904 & v_23905;
assign v_23909 = v_23907 & v_23908;
assign v_23912 = v_23910 & v_23911;
assign v_23915 = v_23913 & v_23914;
assign v_23918 = v_23916 & v_23917;
assign v_23921 = v_23919 & v_23920;
assign v_23924 = v_23922 & v_23923;
assign v_23927 = v_23925 & v_23926;
assign v_23930 = v_23928 & v_23929;
assign v_23933 = v_23931 & v_23932;
assign v_23936 = v_23934 & v_23935;
assign v_23939 = v_23937 & v_23938;
assign v_23942 = v_23940 & v_23941;
assign v_23945 = v_23943 & v_23944;
assign v_23948 = v_23946 & v_23947;
assign v_23951 = v_23949 & v_23950;
assign v_23954 = v_23952 & v_23953;
assign v_23957 = v_23955 & v_23956;
assign v_23960 = v_23958 & v_23959;
assign v_23963 = v_23961 & v_23962;
assign v_23966 = v_23964 & v_23965;
assign v_23969 = v_23967 & v_23968;
assign v_23972 = v_23970 & v_23971;
assign v_23975 = v_23973 & v_23974;
assign v_23978 = v_23976 & v_23977;
assign v_23981 = v_23979 & v_23980;
assign v_23984 = v_23982 & v_23983;
assign v_23987 = v_23985 & v_23986;
assign v_23990 = v_23988 & v_23989;
assign v_23993 = v_23991 & v_23992;
assign v_23996 = v_23994 & v_23995;
assign v_23999 = v_23997 & v_23998;
assign v_24002 = v_24000 & v_24001;
assign v_24003 = v_23813 & v_24002;
assign v_24006 = v_24004 & v_24005;
assign v_24009 = v_24007 & v_24008;
assign v_24012 = v_24010 & v_24011;
assign v_24015 = v_24013 & v_24014;
assign v_24018 = v_24016 & v_24017;
assign v_24021 = v_24019 & v_24020;
assign v_24024 = v_24022 & v_24023;
assign v_24027 = v_24025 & v_24026;
assign v_24030 = v_24028 & v_24029;
assign v_24033 = v_24031 & v_24032;
assign v_24036 = v_24034 & v_24035;
assign v_24039 = v_24037 & v_24038;
assign v_24042 = v_24040 & v_24041;
assign v_24045 = v_24043 & v_24044;
assign v_24048 = v_24046 & v_24047;
assign v_24051 = v_24049 & v_24050;
assign v_24054 = v_24052 & v_24053;
assign v_24057 = v_24055 & v_24056;
assign v_24060 = v_24058 & v_24059;
assign v_24063 = v_24061 & v_24062;
assign v_24066 = v_24064 & v_24065;
assign v_24069 = v_24067 & v_24068;
assign v_24072 = v_24070 & v_24071;
assign v_24075 = v_24073 & v_24074;
assign v_24078 = v_24076 & v_24077;
assign v_24081 = v_24079 & v_24080;
assign v_24084 = v_24082 & v_24083;
assign v_24087 = v_24085 & v_24086;
assign v_24090 = v_24088 & v_24089;
assign v_24093 = v_24091 & v_24092;
assign v_24096 = v_24094 & v_24095;
assign v_24099 = v_24097 & v_24098;
assign v_24102 = v_24100 & v_24101;
assign v_24105 = v_24103 & v_24104;
assign v_24108 = v_24106 & v_24107;
assign v_24111 = v_24109 & v_24110;
assign v_24114 = v_24112 & v_24113;
assign v_24117 = v_24115 & v_24116;
assign v_24120 = v_24118 & v_24119;
assign v_24123 = v_24121 & v_24122;
assign v_24126 = v_24124 & v_24125;
assign v_24129 = v_24127 & v_24128;
assign v_24132 = v_24130 & v_24131;
assign v_24135 = v_24133 & v_24134;
assign v_24138 = v_24136 & v_24137;
assign v_24141 = v_24139 & v_24140;
assign v_24144 = v_24142 & v_24143;
assign v_24147 = v_24145 & v_24146;
assign v_24150 = v_24148 & v_24149;
assign v_24153 = v_24151 & v_24152;
assign v_24156 = v_24154 & v_24155;
assign v_24159 = v_24157 & v_24158;
assign v_24162 = v_24160 & v_24161;
assign v_24165 = v_24163 & v_24164;
assign v_24168 = v_24166 & v_24167;
assign v_24171 = v_24169 & v_24170;
assign v_24174 = v_24172 & v_24173;
assign v_24177 = v_24175 & v_24176;
assign v_24180 = v_24178 & v_24179;
assign v_24183 = v_24181 & v_24182;
assign v_24186 = v_24184 & v_24185;
assign v_24189 = v_24187 & v_24188;
assign v_24192 = v_24190 & v_24191;
assign v_24193 = v_24003 & v_24192;
assign v_24196 = v_24194 & v_24195;
assign v_24199 = v_24197 & v_24198;
assign v_24202 = v_24200 & v_24201;
assign v_24205 = v_24203 & v_24204;
assign v_24208 = v_24206 & v_24207;
assign v_24211 = v_24209 & v_24210;
assign v_24214 = v_24212 & v_24213;
assign v_24217 = v_24215 & v_24216;
assign v_24220 = v_24218 & v_24219;
assign v_24223 = v_24221 & v_24222;
assign v_24226 = v_24224 & v_24225;
assign v_24229 = v_24227 & v_24228;
assign v_24232 = v_24230 & v_24231;
assign v_24235 = v_24233 & v_24234;
assign v_24238 = v_24236 & v_24237;
assign v_24241 = v_24239 & v_24240;
assign v_24244 = v_24242 & v_24243;
assign v_24247 = v_24245 & v_24246;
assign v_24250 = v_24248 & v_24249;
assign v_24253 = v_24251 & v_24252;
assign v_24256 = v_24254 & v_24255;
assign v_24259 = v_24257 & v_24258;
assign v_24262 = v_24260 & v_24261;
assign v_24265 = v_24263 & v_24264;
assign v_24268 = v_24266 & v_24267;
assign v_24271 = v_24269 & v_24270;
assign v_24274 = v_24272 & v_24273;
assign v_24277 = v_24275 & v_24276;
assign v_24280 = v_24278 & v_24279;
assign v_24283 = v_24281 & v_24282;
assign v_24286 = v_24284 & v_24285;
assign v_24289 = v_24287 & v_24288;
assign v_24292 = v_24290 & v_24291;
assign v_24295 = v_24293 & v_24294;
assign v_24298 = v_24296 & v_24297;
assign v_24301 = v_24299 & v_24300;
assign v_24304 = v_24302 & v_24303;
assign v_24307 = v_24305 & v_24306;
assign v_24310 = v_24308 & v_24309;
assign v_24313 = v_24311 & v_24312;
assign v_24316 = v_24314 & v_24315;
assign v_24319 = v_24317 & v_24318;
assign v_24322 = v_24320 & v_24321;
assign v_24325 = v_24323 & v_24324;
assign v_24328 = v_24326 & v_24327;
assign v_24331 = v_24329 & v_24330;
assign v_24334 = v_24332 & v_24333;
assign v_24337 = v_24335 & v_24336;
assign v_24340 = v_24338 & v_24339;
assign v_24343 = v_24341 & v_24342;
assign v_24346 = v_24344 & v_24345;
assign v_24349 = v_24347 & v_24348;
assign v_24352 = v_24350 & v_24351;
assign v_24355 = v_24353 & v_24354;
assign v_24358 = v_24356 & v_24357;
assign v_24361 = v_24359 & v_24360;
assign v_24364 = v_24362 & v_24363;
assign v_24367 = v_24365 & v_24366;
assign v_24370 = v_24368 & v_24369;
assign v_24373 = v_24371 & v_24372;
assign v_24376 = v_24374 & v_24375;
assign v_24379 = v_24377 & v_24378;
assign v_24382 = v_24380 & v_24381;
assign v_24383 = v_24193 & v_24382;
assign v_24386 = v_24384 & v_24385;
assign v_24389 = v_24387 & v_24388;
assign v_24392 = v_24390 & v_24391;
assign v_24395 = v_24393 & v_24394;
assign v_24398 = v_24396 & v_24397;
assign v_24401 = v_24399 & v_24400;
assign v_24404 = v_24402 & v_24403;
assign v_24407 = v_24405 & v_24406;
assign v_24410 = v_24408 & v_24409;
assign v_24413 = v_24411 & v_24412;
assign v_24416 = v_24414 & v_24415;
assign v_24419 = v_24417 & v_24418;
assign v_24422 = v_24420 & v_24421;
assign v_24425 = v_24423 & v_24424;
assign v_24428 = v_24426 & v_24427;
assign v_24431 = v_24429 & v_24430;
assign v_24434 = v_24432 & v_24433;
assign v_24437 = v_24435 & v_24436;
assign v_24440 = v_24438 & v_24439;
assign v_24443 = v_24441 & v_24442;
assign v_24446 = v_24444 & v_24445;
assign v_24449 = v_24447 & v_24448;
assign v_24452 = v_24450 & v_24451;
assign v_24455 = v_24453 & v_24454;
assign v_24458 = v_24456 & v_24457;
assign v_24461 = v_24459 & v_24460;
assign v_24464 = v_24462 & v_24463;
assign v_24467 = v_24465 & v_24466;
assign v_24470 = v_24468 & v_24469;
assign v_24473 = v_24471 & v_24472;
assign v_24476 = v_24474 & v_24475;
assign v_24479 = v_24477 & v_24478;
assign v_24482 = v_24480 & v_24481;
assign v_24485 = v_24483 & v_24484;
assign v_24488 = v_24486 & v_24487;
assign v_24491 = v_24489 & v_24490;
assign v_24494 = v_24492 & v_24493;
assign v_24497 = v_24495 & v_24496;
assign v_24500 = v_24498 & v_24499;
assign v_24503 = v_24501 & v_24502;
assign v_24506 = v_24504 & v_24505;
assign v_24509 = v_24507 & v_24508;
assign v_24512 = v_24510 & v_24511;
assign v_24515 = v_24513 & v_24514;
assign v_24518 = v_24516 & v_24517;
assign v_24521 = v_24519 & v_24520;
assign v_24524 = v_24522 & v_24523;
assign v_24527 = v_24525 & v_24526;
assign v_24530 = v_24528 & v_24529;
assign v_24533 = v_24531 & v_24532;
assign v_24536 = v_24534 & v_24535;
assign v_24539 = v_24537 & v_24538;
assign v_24542 = v_24540 & v_24541;
assign v_24545 = v_24543 & v_24544;
assign v_24548 = v_24546 & v_24547;
assign v_24551 = v_24549 & v_24550;
assign v_24554 = v_24552 & v_24553;
assign v_24557 = v_24555 & v_24556;
assign v_24560 = v_24558 & v_24559;
assign v_24563 = v_24561 & v_24562;
assign v_24566 = v_24564 & v_24565;
assign v_24569 = v_24567 & v_24568;
assign v_24572 = v_24570 & v_24571;
assign v_24573 = v_24383 & v_24572;
assign v_24576 = v_24574 & v_24575;
assign v_24579 = v_24577 & v_24578;
assign v_24582 = v_24580 & v_24581;
assign v_24585 = v_24583 & v_24584;
assign v_24588 = v_24586 & v_24587;
assign v_24591 = v_24589 & v_24590;
assign v_24594 = v_24592 & v_24593;
assign v_24597 = v_24595 & v_24596;
assign v_24600 = v_24598 & v_24599;
assign v_24603 = v_24601 & v_24602;
assign v_24606 = v_24604 & v_24605;
assign v_24609 = v_24607 & v_24608;
assign v_24612 = v_24610 & v_24611;
assign v_24615 = v_24613 & v_24614;
assign v_24618 = v_24616 & v_24617;
assign v_24621 = v_24619 & v_24620;
assign v_24624 = v_24622 & v_24623;
assign v_24627 = v_24625 & v_24626;
assign v_24630 = v_24628 & v_24629;
assign v_24633 = v_24631 & v_24632;
assign v_24636 = v_24634 & v_24635;
assign v_24639 = v_24637 & v_24638;
assign v_24642 = v_24640 & v_24641;
assign v_24645 = v_24643 & v_24644;
assign v_24648 = v_24646 & v_24647;
assign v_24651 = v_24649 & v_24650;
assign v_24654 = v_24652 & v_24653;
assign v_24657 = v_24655 & v_24656;
assign v_24660 = v_24658 & v_24659;
assign v_24663 = v_24661 & v_24662;
assign v_24666 = v_24664 & v_24665;
assign v_24669 = v_24667 & v_24668;
assign v_24672 = v_24670 & v_24671;
assign v_24675 = v_24673 & v_24674;
assign v_24678 = v_24676 & v_24677;
assign v_24681 = v_24679 & v_24680;
assign v_24684 = v_24682 & v_24683;
assign v_24687 = v_24685 & v_24686;
assign v_24690 = v_24688 & v_24689;
assign v_24693 = v_24691 & v_24692;
assign v_24696 = v_24694 & v_24695;
assign v_24699 = v_24697 & v_24698;
assign v_24702 = v_24700 & v_24701;
assign v_24705 = v_24703 & v_24704;
assign v_24708 = v_24706 & v_24707;
assign v_24711 = v_24709 & v_24710;
assign v_24714 = v_24712 & v_24713;
assign v_24717 = v_24715 & v_24716;
assign v_24720 = v_24718 & v_24719;
assign v_24723 = v_24721 & v_24722;
assign v_24726 = v_24724 & v_24725;
assign v_24729 = v_24727 & v_24728;
assign v_24732 = v_24730 & v_24731;
assign v_24735 = v_24733 & v_24734;
assign v_24738 = v_24736 & v_24737;
assign v_24741 = v_24739 & v_24740;
assign v_24744 = v_24742 & v_24743;
assign v_24747 = v_24745 & v_24746;
assign v_24750 = v_24748 & v_24749;
assign v_24753 = v_24751 & v_24752;
assign v_24756 = v_24754 & v_24755;
assign v_24759 = v_24757 & v_24758;
assign v_24762 = v_24760 & v_24761;
assign v_24763 = v_24573 & v_24762;
assign v_24766 = v_24764 & v_24765;
assign v_24769 = v_24767 & v_24768;
assign v_24772 = v_24770 & v_24771;
assign v_24775 = v_24773 & v_24774;
assign v_24778 = v_24776 & v_24777;
assign v_24781 = v_24779 & v_24780;
assign v_24784 = v_24782 & v_24783;
assign v_24787 = v_24785 & v_24786;
assign v_24790 = v_24788 & v_24789;
assign v_24793 = v_24791 & v_24792;
assign v_24796 = v_24794 & v_24795;
assign v_24799 = v_24797 & v_24798;
assign v_24802 = v_24800 & v_24801;
assign v_24805 = v_24803 & v_24804;
assign v_24808 = v_24806 & v_24807;
assign v_24811 = v_24809 & v_24810;
assign v_24814 = v_24812 & v_24813;
assign v_24817 = v_24815 & v_24816;
assign v_24820 = v_24818 & v_24819;
assign v_24823 = v_24821 & v_24822;
assign v_24826 = v_24824 & v_24825;
assign v_24829 = v_24827 & v_24828;
assign v_24832 = v_24830 & v_24831;
assign v_24835 = v_24833 & v_24834;
assign v_24838 = v_24836 & v_24837;
assign v_24841 = v_24839 & v_24840;
assign v_24844 = v_24842 & v_24843;
assign v_24847 = v_24845 & v_24846;
assign v_24850 = v_24848 & v_24849;
assign v_24853 = v_24851 & v_24852;
assign v_24856 = v_24854 & v_24855;
assign v_24859 = v_24857 & v_24858;
assign v_24862 = v_24860 & v_24861;
assign v_24865 = v_24863 & v_24864;
assign v_24868 = v_24866 & v_24867;
assign v_24871 = v_24869 & v_24870;
assign v_24874 = v_24872 & v_24873;
assign v_24877 = v_24875 & v_24876;
assign v_24880 = v_24878 & v_24879;
assign v_24883 = v_24881 & v_24882;
assign v_24886 = v_24884 & v_24885;
assign v_24889 = v_24887 & v_24888;
assign v_24892 = v_24890 & v_24891;
assign v_24895 = v_24893 & v_24894;
assign v_24898 = v_24896 & v_24897;
assign v_24901 = v_24899 & v_24900;
assign v_24904 = v_24902 & v_24903;
assign v_24907 = v_24905 & v_24906;
assign v_24910 = v_24908 & v_24909;
assign v_24913 = v_24911 & v_24912;
assign v_24916 = v_24914 & v_24915;
assign v_24919 = v_24917 & v_24918;
assign v_24922 = v_24920 & v_24921;
assign v_24925 = v_24923 & v_24924;
assign v_24928 = v_24926 & v_24927;
assign v_24931 = v_24929 & v_24930;
assign v_24934 = v_24932 & v_24933;
assign v_24937 = v_24935 & v_24936;
assign v_24940 = v_24938 & v_24939;
assign v_24943 = v_24941 & v_24942;
assign v_24946 = v_24944 & v_24945;
assign v_24949 = v_24947 & v_24948;
assign v_24952 = v_24950 & v_24951;
assign v_24953 = v_24763 & v_24952;
assign v_24956 = v_24954 & v_24955;
assign v_24959 = v_24957 & v_24958;
assign v_24962 = v_24960 & v_24961;
assign v_24965 = v_24963 & v_24964;
assign v_24968 = v_24966 & v_24967;
assign v_24971 = v_24969 & v_24970;
assign v_24974 = v_24972 & v_24973;
assign v_24977 = v_24975 & v_24976;
assign v_24980 = v_24978 & v_24979;
assign v_24983 = v_24981 & v_24982;
assign v_24986 = v_24984 & v_24985;
assign v_24989 = v_24987 & v_24988;
assign v_24992 = v_24990 & v_24991;
assign v_24995 = v_24993 & v_24994;
assign v_24998 = v_24996 & v_24997;
assign v_25001 = v_24999 & v_25000;
assign v_25004 = v_25002 & v_25003;
assign v_25007 = v_25005 & v_25006;
assign v_25010 = v_25008 & v_25009;
assign v_25013 = v_25011 & v_25012;
assign v_25016 = v_25014 & v_25015;
assign v_25019 = v_25017 & v_25018;
assign v_25022 = v_25020 & v_25021;
assign v_25025 = v_25023 & v_25024;
assign v_25028 = v_25026 & v_25027;
assign v_25031 = v_25029 & v_25030;
assign v_25034 = v_25032 & v_25033;
assign v_25037 = v_25035 & v_25036;
assign v_25040 = v_25038 & v_25039;
assign v_25043 = v_25041 & v_25042;
assign v_25046 = v_25044 & v_25045;
assign v_25049 = v_25047 & v_25048;
assign v_25052 = v_25050 & v_25051;
assign v_25055 = v_25053 & v_25054;
assign v_25058 = v_25056 & v_25057;
assign v_25061 = v_25059 & v_25060;
assign v_25064 = v_25062 & v_25063;
assign v_25067 = v_25065 & v_25066;
assign v_25070 = v_25068 & v_25069;
assign v_25073 = v_25071 & v_25072;
assign v_25076 = v_25074 & v_25075;
assign v_25079 = v_25077 & v_25078;
assign v_25082 = v_25080 & v_25081;
assign v_25085 = v_25083 & v_25084;
assign v_25088 = v_25086 & v_25087;
assign v_25091 = v_25089 & v_25090;
assign v_25094 = v_25092 & v_25093;
assign v_25097 = v_25095 & v_25096;
assign v_25100 = v_25098 & v_25099;
assign v_25103 = v_25101 & v_25102;
assign v_25106 = v_25104 & v_25105;
assign v_25109 = v_25107 & v_25108;
assign v_25112 = v_25110 & v_25111;
assign v_25115 = v_25113 & v_25114;
assign v_25118 = v_25116 & v_25117;
assign v_25121 = v_25119 & v_25120;
assign v_25124 = v_25122 & v_25123;
assign v_25127 = v_25125 & v_25126;
assign v_25130 = v_25128 & v_25129;
assign v_25133 = v_25131 & v_25132;
assign v_25136 = v_25134 & v_25135;
assign v_25139 = v_25137 & v_25138;
assign v_25142 = v_25140 & v_25141;
assign v_25145 = v_25143 & v_25144;
assign v_25148 = v_25146 & v_25147;
assign v_25151 = v_25149 & v_25150;
assign v_25154 = v_25152 & v_25153;
assign v_25157 = v_25155 & v_25156;
assign v_25160 = v_25158 & v_25159;
assign v_25163 = v_25161 & v_25162;
assign v_25166 = v_25164 & v_25165;
assign v_25169 = v_25167 & v_25168;
assign v_25172 = v_25170 & v_25171;
assign v_25175 = v_25173 & v_25174;
assign v_25178 = v_25176 & v_25177;
assign v_25181 = v_25179 & v_25180;
assign v_25184 = v_25182 & v_25183;
assign v_25187 = v_25185 & v_25186;
assign v_25190 = v_25188 & v_25189;
assign v_25193 = v_25191 & v_25192;
assign v_25196 = v_25194 & v_25195;
assign v_25199 = v_25197 & v_25198;
assign v_25202 = v_25200 & v_25201;
assign v_25205 = v_25203 & v_25204;
assign v_25208 = v_25206 & v_25207;
assign v_25211 = v_25209 & v_25210;
assign v_25214 = v_25212 & v_25213;
assign v_25217 = v_25215 & v_25216;
assign v_25220 = v_25218 & v_25219;
assign v_25223 = v_25221 & v_25222;
assign v_25226 = v_25224 & v_25225;
assign v_25229 = v_25227 & v_25228;
assign v_25232 = v_25230 & v_25231;
assign v_25235 = v_25233 & v_25234;
assign v_25238 = v_25236 & v_25237;
assign v_25241 = v_25239 & v_25240;
assign v_25244 = v_25242 & v_25243;
assign v_25247 = v_25245 & v_25246;
assign v_25250 = v_25248 & v_25249;
assign v_25253 = v_25251 & v_25252;
assign v_25256 = v_25254 & v_25255;
assign v_25259 = v_25257 & v_25258;
assign v_25262 = v_25260 & v_25261;
assign v_25265 = v_25263 & v_25264;
assign v_25268 = v_25266 & v_25267;
assign v_25271 = v_25269 & v_25270;
assign v_25274 = v_25272 & v_25273;
assign v_25277 = v_25275 & v_25276;
assign v_25280 = v_25278 & v_25279;
assign v_25283 = v_25281 & v_25282;
assign v_25286 = v_25284 & v_25285;
assign v_25289 = v_25287 & v_25288;
assign v_25292 = v_25290 & v_25291;
assign v_25295 = v_25293 & v_25294;
assign v_25298 = v_25296 & v_25297;
assign v_25301 = v_25299 & v_25300;
assign v_25304 = v_25302 & v_25303;
assign v_25307 = v_25305 & v_25306;
assign v_25310 = v_25308 & v_25309;
assign v_25313 = v_25311 & v_25312;
assign v_25316 = v_25314 & v_25315;
assign v_25319 = v_25317 & v_25318;
assign v_25322 = v_25320 & v_25321;
assign v_25325 = v_25323 & v_25324;
assign v_25328 = v_25326 & v_25327;
assign v_25331 = v_25329 & v_25330;
assign v_25332 = v_25142 & v_25331;
assign v_25335 = v_25333 & v_25334;
assign v_25338 = v_25336 & v_25337;
assign v_25341 = v_25339 & v_25340;
assign v_25344 = v_25342 & v_25343;
assign v_25347 = v_25345 & v_25346;
assign v_25350 = v_25348 & v_25349;
assign v_25353 = v_25351 & v_25352;
assign v_25356 = v_25354 & v_25355;
assign v_25359 = v_25357 & v_25358;
assign v_25362 = v_25360 & v_25361;
assign v_25365 = v_25363 & v_25364;
assign v_25368 = v_25366 & v_25367;
assign v_25371 = v_25369 & v_25370;
assign v_25374 = v_25372 & v_25373;
assign v_25377 = v_25375 & v_25376;
assign v_25380 = v_25378 & v_25379;
assign v_25383 = v_25381 & v_25382;
assign v_25386 = v_25384 & v_25385;
assign v_25389 = v_25387 & v_25388;
assign v_25392 = v_25390 & v_25391;
assign v_25395 = v_25393 & v_25394;
assign v_25398 = v_25396 & v_25397;
assign v_25401 = v_25399 & v_25400;
assign v_25404 = v_25402 & v_25403;
assign v_25407 = v_25405 & v_25406;
assign v_25410 = v_25408 & v_25409;
assign v_25413 = v_25411 & v_25412;
assign v_25416 = v_25414 & v_25415;
assign v_25419 = v_25417 & v_25418;
assign v_25422 = v_25420 & v_25421;
assign v_25425 = v_25423 & v_25424;
assign v_25428 = v_25426 & v_25427;
assign v_25431 = v_25429 & v_25430;
assign v_25434 = v_25432 & v_25433;
assign v_25437 = v_25435 & v_25436;
assign v_25440 = v_25438 & v_25439;
assign v_25443 = v_25441 & v_25442;
assign v_25446 = v_25444 & v_25445;
assign v_25449 = v_25447 & v_25448;
assign v_25452 = v_25450 & v_25451;
assign v_25455 = v_25453 & v_25454;
assign v_25458 = v_25456 & v_25457;
assign v_25461 = v_25459 & v_25460;
assign v_25464 = v_25462 & v_25463;
assign v_25467 = v_25465 & v_25466;
assign v_25470 = v_25468 & v_25469;
assign v_25473 = v_25471 & v_25472;
assign v_25476 = v_25474 & v_25475;
assign v_25479 = v_25477 & v_25478;
assign v_25482 = v_25480 & v_25481;
assign v_25485 = v_25483 & v_25484;
assign v_25488 = v_25486 & v_25487;
assign v_25491 = v_25489 & v_25490;
assign v_25494 = v_25492 & v_25493;
assign v_25497 = v_25495 & v_25496;
assign v_25500 = v_25498 & v_25499;
assign v_25503 = v_25501 & v_25502;
assign v_25506 = v_25504 & v_25505;
assign v_25509 = v_25507 & v_25508;
assign v_25512 = v_25510 & v_25511;
assign v_25515 = v_25513 & v_25514;
assign v_25518 = v_25516 & v_25517;
assign v_25521 = v_25519 & v_25520;
assign v_25522 = v_25332 & v_25521;
assign v_25525 = v_25523 & v_25524;
assign v_25528 = v_25526 & v_25527;
assign v_25531 = v_25529 & v_25530;
assign v_25534 = v_25532 & v_25533;
assign v_25537 = v_25535 & v_25536;
assign v_25540 = v_25538 & v_25539;
assign v_25543 = v_25541 & v_25542;
assign v_25546 = v_25544 & v_25545;
assign v_25549 = v_25547 & v_25548;
assign v_25552 = v_25550 & v_25551;
assign v_25555 = v_25553 & v_25554;
assign v_25558 = v_25556 & v_25557;
assign v_25561 = v_25559 & v_25560;
assign v_25564 = v_25562 & v_25563;
assign v_25567 = v_25565 & v_25566;
assign v_25570 = v_25568 & v_25569;
assign v_25573 = v_25571 & v_25572;
assign v_25576 = v_25574 & v_25575;
assign v_25579 = v_25577 & v_25578;
assign v_25582 = v_25580 & v_25581;
assign v_25585 = v_25583 & v_25584;
assign v_25588 = v_25586 & v_25587;
assign v_25591 = v_25589 & v_25590;
assign v_25594 = v_25592 & v_25593;
assign v_25597 = v_25595 & v_25596;
assign v_25600 = v_25598 & v_25599;
assign v_25603 = v_25601 & v_25602;
assign v_25606 = v_25604 & v_25605;
assign v_25609 = v_25607 & v_25608;
assign v_25612 = v_25610 & v_25611;
assign v_25615 = v_25613 & v_25614;
assign v_25618 = v_25616 & v_25617;
assign v_25621 = v_25619 & v_25620;
assign v_25624 = v_25622 & v_25623;
assign v_25627 = v_25625 & v_25626;
assign v_25630 = v_25628 & v_25629;
assign v_25633 = v_25631 & v_25632;
assign v_25636 = v_25634 & v_25635;
assign v_25639 = v_25637 & v_25638;
assign v_25642 = v_25640 & v_25641;
assign v_25645 = v_25643 & v_25644;
assign v_25648 = v_25646 & v_25647;
assign v_25651 = v_25649 & v_25650;
assign v_25654 = v_25652 & v_25653;
assign v_25657 = v_25655 & v_25656;
assign v_25660 = v_25658 & v_25659;
assign v_25663 = v_25661 & v_25662;
assign v_25666 = v_25664 & v_25665;
assign v_25669 = v_25667 & v_25668;
assign v_25672 = v_25670 & v_25671;
assign v_25675 = v_25673 & v_25674;
assign v_25678 = v_25676 & v_25677;
assign v_25681 = v_25679 & v_25680;
assign v_25684 = v_25682 & v_25683;
assign v_25687 = v_25685 & v_25686;
assign v_25690 = v_25688 & v_25689;
assign v_25693 = v_25691 & v_25692;
assign v_25696 = v_25694 & v_25695;
assign v_25699 = v_25697 & v_25698;
assign v_25702 = v_25700 & v_25701;
assign v_25705 = v_25703 & v_25704;
assign v_25708 = v_25706 & v_25707;
assign v_25711 = v_25709 & v_25710;
assign v_25712 = v_25522 & v_25711;
assign v_25715 = v_25713 & v_25714;
assign v_25718 = v_25716 & v_25717;
assign v_25721 = v_25719 & v_25720;
assign v_25724 = v_25722 & v_25723;
assign v_25727 = v_25725 & v_25726;
assign v_25730 = v_25728 & v_25729;
assign v_25733 = v_25731 & v_25732;
assign v_25736 = v_25734 & v_25735;
assign v_25739 = v_25737 & v_25738;
assign v_25742 = v_25740 & v_25741;
assign v_25745 = v_25743 & v_25744;
assign v_25748 = v_25746 & v_25747;
assign v_25751 = v_25749 & v_25750;
assign v_25754 = v_25752 & v_25753;
assign v_25757 = v_25755 & v_25756;
assign v_25760 = v_25758 & v_25759;
assign v_25763 = v_25761 & v_25762;
assign v_25766 = v_25764 & v_25765;
assign v_25769 = v_25767 & v_25768;
assign v_25772 = v_25770 & v_25771;
assign v_25775 = v_25773 & v_25774;
assign v_25778 = v_25776 & v_25777;
assign v_25781 = v_25779 & v_25780;
assign v_25784 = v_25782 & v_25783;
assign v_25787 = v_25785 & v_25786;
assign v_25790 = v_25788 & v_25789;
assign v_25793 = v_25791 & v_25792;
assign v_25796 = v_25794 & v_25795;
assign v_25799 = v_25797 & v_25798;
assign v_25802 = v_25800 & v_25801;
assign v_25805 = v_25803 & v_25804;
assign v_25808 = v_25806 & v_25807;
assign v_25811 = v_25809 & v_25810;
assign v_25814 = v_25812 & v_25813;
assign v_25817 = v_25815 & v_25816;
assign v_25820 = v_25818 & v_25819;
assign v_25823 = v_25821 & v_25822;
assign v_25826 = v_25824 & v_25825;
assign v_25829 = v_25827 & v_25828;
assign v_25832 = v_25830 & v_25831;
assign v_25835 = v_25833 & v_25834;
assign v_25838 = v_25836 & v_25837;
assign v_25841 = v_25839 & v_25840;
assign v_25844 = v_25842 & v_25843;
assign v_25847 = v_25845 & v_25846;
assign v_25850 = v_25848 & v_25849;
assign v_25853 = v_25851 & v_25852;
assign v_25856 = v_25854 & v_25855;
assign v_25859 = v_25857 & v_25858;
assign v_25862 = v_25860 & v_25861;
assign v_25865 = v_25863 & v_25864;
assign v_25868 = v_25866 & v_25867;
assign v_25871 = v_25869 & v_25870;
assign v_25874 = v_25872 & v_25873;
assign v_25877 = v_25875 & v_25876;
assign v_25880 = v_25878 & v_25879;
assign v_25883 = v_25881 & v_25882;
assign v_25886 = v_25884 & v_25885;
assign v_25889 = v_25887 & v_25888;
assign v_25892 = v_25890 & v_25891;
assign v_25895 = v_25893 & v_25894;
assign v_25898 = v_25896 & v_25897;
assign v_25901 = v_25899 & v_25900;
assign v_25902 = v_25712 & v_25901;
assign v_25905 = v_25903 & v_25904;
assign v_25908 = v_25906 & v_25907;
assign v_25911 = v_25909 & v_25910;
assign v_25914 = v_25912 & v_25913;
assign v_25917 = v_25915 & v_25916;
assign v_25920 = v_25918 & v_25919;
assign v_25923 = v_25921 & v_25922;
assign v_25926 = v_25924 & v_25925;
assign v_25929 = v_25927 & v_25928;
assign v_25932 = v_25930 & v_25931;
assign v_25935 = v_25933 & v_25934;
assign v_25938 = v_25936 & v_25937;
assign v_25941 = v_25939 & v_25940;
assign v_25944 = v_25942 & v_25943;
assign v_25947 = v_25945 & v_25946;
assign v_25950 = v_25948 & v_25949;
assign v_25953 = v_25951 & v_25952;
assign v_25956 = v_25954 & v_25955;
assign v_25959 = v_25957 & v_25958;
assign v_25962 = v_25960 & v_25961;
assign v_25965 = v_25963 & v_25964;
assign v_25968 = v_25966 & v_25967;
assign v_25971 = v_25969 & v_25970;
assign v_25974 = v_25972 & v_25973;
assign v_25977 = v_25975 & v_25976;
assign v_25980 = v_25978 & v_25979;
assign v_25983 = v_25981 & v_25982;
assign v_25986 = v_25984 & v_25985;
assign v_25989 = v_25987 & v_25988;
assign v_25992 = v_25990 & v_25991;
assign v_25995 = v_25993 & v_25994;
assign v_25998 = v_25996 & v_25997;
assign v_26001 = v_25999 & v_26000;
assign v_26004 = v_26002 & v_26003;
assign v_26007 = v_26005 & v_26006;
assign v_26010 = v_26008 & v_26009;
assign v_26013 = v_26011 & v_26012;
assign v_26016 = v_26014 & v_26015;
assign v_26019 = v_26017 & v_26018;
assign v_26022 = v_26020 & v_26021;
assign v_26025 = v_26023 & v_26024;
assign v_26028 = v_26026 & v_26027;
assign v_26031 = v_26029 & v_26030;
assign v_26034 = v_26032 & v_26033;
assign v_26037 = v_26035 & v_26036;
assign v_26040 = v_26038 & v_26039;
assign v_26043 = v_26041 & v_26042;
assign v_26046 = v_26044 & v_26045;
assign v_26049 = v_26047 & v_26048;
assign v_26052 = v_26050 & v_26051;
assign v_26055 = v_26053 & v_26054;
assign v_26058 = v_26056 & v_26057;
assign v_26061 = v_26059 & v_26060;
assign v_26064 = v_26062 & v_26063;
assign v_26067 = v_26065 & v_26066;
assign v_26070 = v_26068 & v_26069;
assign v_26073 = v_26071 & v_26072;
assign v_26076 = v_26074 & v_26075;
assign v_26079 = v_26077 & v_26078;
assign v_26082 = v_26080 & v_26081;
assign v_26085 = v_26083 & v_26084;
assign v_26088 = v_26086 & v_26087;
assign v_26091 = v_26089 & v_26090;
assign v_26092 = v_25902 & v_26091;
assign v_26093 = v_22787 & v_26092;
assign v_26096 = v_26094 & v_26095;
assign v_26099 = v_26097 & v_26098;
assign v_26102 = v_26100 & v_26101;
assign v_26105 = v_26103 & v_26104;
assign v_26108 = v_26106 & v_26107;
assign v_26111 = v_26109 & v_26110;
assign v_26114 = v_26112 & v_26113;
assign v_26117 = v_26115 & v_26116;
assign v_26120 = v_26118 & v_26119;
assign v_26123 = v_26121 & v_26122;
assign v_26126 = v_26124 & v_26125;
assign v_26129 = v_26127 & v_26128;
assign v_26132 = v_26130 & v_26131;
assign v_26135 = v_26133 & v_26134;
assign v_26138 = v_26136 & v_26137;
assign v_26141 = v_26139 & v_26140;
assign v_26144 = v_26142 & v_26143;
assign v_26147 = v_26145 & v_26146;
assign v_26150 = v_26148 & v_26149;
assign v_26153 = v_26151 & v_26152;
assign v_26156 = v_26154 & v_26155;
assign v_26159 = v_26157 & v_26158;
assign v_26162 = v_26160 & v_26161;
assign v_26165 = v_26163 & v_26164;
assign v_26168 = v_26166 & v_26167;
assign v_26171 = v_26169 & v_26170;
assign v_26174 = v_26172 & v_26173;
assign v_26177 = v_26175 & v_26176;
assign v_26180 = v_26178 & v_26179;
assign v_26183 = v_26181 & v_26182;
assign v_26186 = v_26184 & v_26185;
assign v_26189 = v_26187 & v_26188;
assign v_26192 = v_26190 & v_26191;
assign v_26195 = v_26193 & v_26194;
assign v_26198 = v_26196 & v_26197;
assign v_26201 = v_26199 & v_26200;
assign v_26204 = v_26202 & v_26203;
assign v_26207 = v_26205 & v_26206;
assign v_26210 = v_26208 & v_26209;
assign v_26213 = v_26211 & v_26212;
assign v_26216 = v_26214 & v_26215;
assign v_26219 = v_26217 & v_26218;
assign v_26222 = v_26220 & v_26221;
assign v_26225 = v_26223 & v_26224;
assign v_26228 = v_26226 & v_26227;
assign v_26231 = v_26229 & v_26230;
assign v_26234 = v_26232 & v_26233;
assign v_26237 = v_26235 & v_26236;
assign v_26240 = v_26238 & v_26239;
assign v_26243 = v_26241 & v_26242;
assign v_26246 = v_26244 & v_26245;
assign v_26249 = v_26247 & v_26248;
assign v_26252 = v_26250 & v_26251;
assign v_26255 = v_26253 & v_26254;
assign v_26258 = v_26256 & v_26257;
assign v_26261 = v_26259 & v_26260;
assign v_26264 = v_26262 & v_26263;
assign v_26267 = v_26265 & v_26266;
assign v_26270 = v_26268 & v_26269;
assign v_26273 = v_26271 & v_26272;
assign v_26276 = v_26274 & v_26275;
assign v_26279 = v_26277 & v_26278;
assign v_26282 = v_26280 & v_26281;
assign v_26283 = v_26093 & v_26282;
assign v_26284 = ~v_10414 & ~v_10421;
assign v_26285 = ~v_10427 & v_26284;
assign v_26286 = ~v_10433 & v_26285;
assign v_26287 = ~v_10439 & v_26286;
assign v_26288 = ~v_10445 & v_26287;
assign v_26289 = ~v_10451 & v_26288;
assign v_26290 = ~v_4 & v_26289;
assign v_26291 = v_26283 & v_26290;
assign v_26292 = v_24953 & v_26291;
assign v_26293 = ~v_10462 & v_26292;
assign v_26297 = v_26295 & v_26296;
assign v_26300 = v_26298 & v_26299;
assign v_26303 = v_26301 & v_26302;
assign v_26306 = v_26304 & v_26305;
assign v_26309 = v_26307 & v_26308;
assign v_26312 = v_26310 & v_26311;
assign v_26315 = v_26313 & v_26314;
assign v_26318 = v_26316 & v_26317;
assign v_26321 = v_26319 & v_26320;
assign v_26324 = v_26322 & v_26323;
assign v_26327 = v_26325 & v_26326;
assign v_26330 = v_26328 & v_26329;
assign v_26333 = v_26331 & v_26332;
assign v_26336 = v_26334 & v_26335;
assign v_26339 = v_26337 & v_26338;
assign v_26342 = v_26340 & v_26341;
assign v_26345 = v_26343 & v_26344;
assign v_26348 = v_26346 & v_26347;
assign v_26351 = v_26349 & v_26350;
assign v_26354 = v_26352 & v_26353;
assign v_26357 = v_26355 & v_26356;
assign v_26360 = v_26358 & v_26359;
assign v_26363 = v_26361 & v_26362;
assign v_26366 = v_26364 & v_26365;
assign v_26369 = v_26367 & v_26368;
assign v_26372 = v_26370 & v_26371;
assign v_26375 = v_26373 & v_26374;
assign v_26378 = v_26376 & v_26377;
assign v_26381 = v_26379 & v_26380;
assign v_26384 = v_26382 & v_26383;
assign v_26387 = v_26385 & v_26386;
assign v_26390 = v_26388 & v_26389;
assign v_26393 = v_26391 & v_26392;
assign v_26396 = v_26394 & v_26395;
assign v_26399 = v_26397 & v_26398;
assign v_26402 = v_26400 & v_26401;
assign v_26405 = v_26403 & v_26404;
assign v_26408 = v_26406 & v_26407;
assign v_26411 = v_26409 & v_26410;
assign v_26414 = v_26412 & v_26413;
assign v_26417 = v_26415 & v_26416;
assign v_26420 = v_26418 & v_26419;
assign v_26423 = v_26421 & v_26422;
assign v_26426 = v_26424 & v_26425;
assign v_26429 = v_26427 & v_26428;
assign v_26432 = v_26430 & v_26431;
assign v_26435 = v_26433 & v_26434;
assign v_26438 = v_26436 & v_26437;
assign v_26441 = v_26439 & v_26440;
assign v_26444 = v_26442 & v_26443;
assign v_26447 = v_26445 & v_26446;
assign v_26450 = v_26448 & v_26449;
assign v_26453 = v_26451 & v_26452;
assign v_26456 = v_26454 & v_26455;
assign v_26459 = v_26457 & v_26458;
assign v_26462 = v_26460 & v_26461;
assign v_26465 = v_26463 & v_26464;
assign v_26468 = v_26466 & v_26467;
assign v_26471 = v_26469 & v_26470;
assign v_26474 = v_26472 & v_26473;
assign v_26477 = v_26475 & v_26476;
assign v_26480 = v_26478 & v_26479;
assign v_26483 = v_26481 & v_26482;
assign v_26486 = v_26484 & v_26485;
assign v_26489 = v_26487 & v_26488;
assign v_26492 = v_26490 & v_26491;
assign v_26495 = v_26493 & v_26494;
assign v_26498 = v_26496 & v_26497;
assign v_26501 = v_26499 & v_26500;
assign v_26504 = v_26502 & v_26503;
assign v_26507 = v_26505 & v_26506;
assign v_26510 = v_26508 & v_26509;
assign v_26513 = v_26511 & v_26512;
assign v_26516 = v_26514 & v_26515;
assign v_26519 = v_26517 & v_26518;
assign v_26522 = v_26520 & v_26521;
assign v_26525 = v_26523 & v_26524;
assign v_26528 = v_26526 & v_26527;
assign v_26531 = v_26529 & v_26530;
assign v_26534 = v_26532 & v_26533;
assign v_26537 = v_26535 & v_26536;
assign v_26540 = v_26538 & v_26539;
assign v_26543 = v_26541 & v_26542;
assign v_26546 = v_26544 & v_26545;
assign v_26549 = v_26547 & v_26548;
assign v_26552 = v_26550 & v_26551;
assign v_26555 = v_26553 & v_26554;
assign v_26558 = v_26556 & v_26557;
assign v_26561 = v_26559 & v_26560;
assign v_26564 = v_26562 & v_26563;
assign v_26567 = v_26565 & v_26566;
assign v_26570 = v_26568 & v_26569;
assign v_26573 = v_26571 & v_26572;
assign v_26576 = v_26574 & v_26575;
assign v_26579 = v_26577 & v_26578;
assign v_26582 = v_26580 & v_26581;
assign v_26585 = v_26583 & v_26584;
assign v_26588 = v_26586 & v_26587;
assign v_26591 = v_26589 & v_26590;
assign v_26594 = v_26592 & v_26593;
assign v_26597 = v_26595 & v_26596;
assign v_26600 = v_26598 & v_26599;
assign v_26603 = v_26601 & v_26602;
assign v_26606 = v_26604 & v_26605;
assign v_26609 = v_26607 & v_26608;
assign v_26612 = v_26610 & v_26611;
assign v_26615 = v_26613 & v_26614;
assign v_26618 = v_26616 & v_26617;
assign v_26621 = v_26619 & v_26620;
assign v_26624 = v_26622 & v_26623;
assign v_26627 = v_26625 & v_26626;
assign v_26630 = v_26628 & v_26629;
assign v_26633 = v_26631 & v_26632;
assign v_26636 = v_26634 & v_26635;
assign v_26639 = v_26637 & v_26638;
assign v_26642 = v_26640 & v_26641;
assign v_26645 = v_26643 & v_26644;
assign v_26648 = v_26646 & v_26647;
assign v_26651 = v_26649 & v_26650;
assign v_26654 = v_26652 & v_26653;
assign v_26657 = v_26655 & v_26656;
assign v_26660 = v_26658 & v_26659;
assign v_26663 = v_26661 & v_26662;
assign v_26666 = v_26664 & v_26665;
assign v_26669 = v_26667 & v_26668;
assign v_26672 = v_26670 & v_26671;
assign v_26673 = v_26483 & v_26672;
assign v_26676 = v_26674 & v_26675;
assign v_26679 = v_26677 & v_26678;
assign v_26682 = v_26680 & v_26681;
assign v_26685 = v_26683 & v_26684;
assign v_26688 = v_26686 & v_26687;
assign v_26691 = v_26689 & v_26690;
assign v_26694 = v_26692 & v_26693;
assign v_26697 = v_26695 & v_26696;
assign v_26700 = v_26698 & v_26699;
assign v_26703 = v_26701 & v_26702;
assign v_26706 = v_26704 & v_26705;
assign v_26709 = v_26707 & v_26708;
assign v_26712 = v_26710 & v_26711;
assign v_26715 = v_26713 & v_26714;
assign v_26718 = v_26716 & v_26717;
assign v_26721 = v_26719 & v_26720;
assign v_26724 = v_26722 & v_26723;
assign v_26727 = v_26725 & v_26726;
assign v_26730 = v_26728 & v_26729;
assign v_26733 = v_26731 & v_26732;
assign v_26736 = v_26734 & v_26735;
assign v_26739 = v_26737 & v_26738;
assign v_26742 = v_26740 & v_26741;
assign v_26745 = v_26743 & v_26744;
assign v_26748 = v_26746 & v_26747;
assign v_26751 = v_26749 & v_26750;
assign v_26754 = v_26752 & v_26753;
assign v_26757 = v_26755 & v_26756;
assign v_26760 = v_26758 & v_26759;
assign v_26763 = v_26761 & v_26762;
assign v_26766 = v_26764 & v_26765;
assign v_26769 = v_26767 & v_26768;
assign v_26772 = v_26770 & v_26771;
assign v_26775 = v_26773 & v_26774;
assign v_26778 = v_26776 & v_26777;
assign v_26781 = v_26779 & v_26780;
assign v_26784 = v_26782 & v_26783;
assign v_26787 = v_26785 & v_26786;
assign v_26790 = v_26788 & v_26789;
assign v_26793 = v_26791 & v_26792;
assign v_26796 = v_26794 & v_26795;
assign v_26799 = v_26797 & v_26798;
assign v_26802 = v_26800 & v_26801;
assign v_26805 = v_26803 & v_26804;
assign v_26808 = v_26806 & v_26807;
assign v_26811 = v_26809 & v_26810;
assign v_26814 = v_26812 & v_26813;
assign v_26817 = v_26815 & v_26816;
assign v_26820 = v_26818 & v_26819;
assign v_26823 = v_26821 & v_26822;
assign v_26826 = v_26824 & v_26825;
assign v_26829 = v_26827 & v_26828;
assign v_26832 = v_26830 & v_26831;
assign v_26835 = v_26833 & v_26834;
assign v_26838 = v_26836 & v_26837;
assign v_26841 = v_26839 & v_26840;
assign v_26844 = v_26842 & v_26843;
assign v_26847 = v_26845 & v_26846;
assign v_26850 = v_26848 & v_26849;
assign v_26853 = v_26851 & v_26852;
assign v_26856 = v_26854 & v_26855;
assign v_26859 = v_26857 & v_26858;
assign v_26862 = v_26860 & v_26861;
assign v_26863 = v_26673 & v_26862;
assign v_26866 = v_26864 & v_26865;
assign v_26869 = v_26867 & v_26868;
assign v_26872 = v_26870 & v_26871;
assign v_26875 = v_26873 & v_26874;
assign v_26878 = v_26876 & v_26877;
assign v_26881 = v_26879 & v_26880;
assign v_26884 = v_26882 & v_26883;
assign v_26887 = v_26885 & v_26886;
assign v_26890 = v_26888 & v_26889;
assign v_26893 = v_26891 & v_26892;
assign v_26896 = v_26894 & v_26895;
assign v_26899 = v_26897 & v_26898;
assign v_26902 = v_26900 & v_26901;
assign v_26905 = v_26903 & v_26904;
assign v_26908 = v_26906 & v_26907;
assign v_26911 = v_26909 & v_26910;
assign v_26914 = v_26912 & v_26913;
assign v_26917 = v_26915 & v_26916;
assign v_26920 = v_26918 & v_26919;
assign v_26923 = v_26921 & v_26922;
assign v_26926 = v_26924 & v_26925;
assign v_26929 = v_26927 & v_26928;
assign v_26932 = v_26930 & v_26931;
assign v_26935 = v_26933 & v_26934;
assign v_26938 = v_26936 & v_26937;
assign v_26941 = v_26939 & v_26940;
assign v_26944 = v_26942 & v_26943;
assign v_26947 = v_26945 & v_26946;
assign v_26950 = v_26948 & v_26949;
assign v_26953 = v_26951 & v_26952;
assign v_26956 = v_26954 & v_26955;
assign v_26959 = v_26957 & v_26958;
assign v_26962 = v_26960 & v_26961;
assign v_26965 = v_26963 & v_26964;
assign v_26968 = v_26966 & v_26967;
assign v_26971 = v_26969 & v_26970;
assign v_26974 = v_26972 & v_26973;
assign v_26977 = v_26975 & v_26976;
assign v_26980 = v_26978 & v_26979;
assign v_26983 = v_26981 & v_26982;
assign v_26986 = v_26984 & v_26985;
assign v_26989 = v_26987 & v_26988;
assign v_26992 = v_26990 & v_26991;
assign v_26995 = v_26993 & v_26994;
assign v_26998 = v_26996 & v_26997;
assign v_27001 = v_26999 & v_27000;
assign v_27004 = v_27002 & v_27003;
assign v_27007 = v_27005 & v_27006;
assign v_27010 = v_27008 & v_27009;
assign v_27013 = v_27011 & v_27012;
assign v_27016 = v_27014 & v_27015;
assign v_27019 = v_27017 & v_27018;
assign v_27022 = v_27020 & v_27021;
assign v_27025 = v_27023 & v_27024;
assign v_27028 = v_27026 & v_27027;
assign v_27031 = v_27029 & v_27030;
assign v_27034 = v_27032 & v_27033;
assign v_27037 = v_27035 & v_27036;
assign v_27040 = v_27038 & v_27039;
assign v_27043 = v_27041 & v_27042;
assign v_27046 = v_27044 & v_27045;
assign v_27049 = v_27047 & v_27048;
assign v_27052 = v_27050 & v_27051;
assign v_27053 = v_26863 & v_27052;
assign v_27056 = v_27054 & v_27055;
assign v_27059 = v_27057 & v_27058;
assign v_27062 = v_27060 & v_27061;
assign v_27065 = v_27063 & v_27064;
assign v_27068 = v_27066 & v_27067;
assign v_27071 = v_27069 & v_27070;
assign v_27074 = v_27072 & v_27073;
assign v_27077 = v_27075 & v_27076;
assign v_27080 = v_27078 & v_27079;
assign v_27083 = v_27081 & v_27082;
assign v_27086 = v_27084 & v_27085;
assign v_27089 = v_27087 & v_27088;
assign v_27092 = v_27090 & v_27091;
assign v_27095 = v_27093 & v_27094;
assign v_27098 = v_27096 & v_27097;
assign v_27101 = v_27099 & v_27100;
assign v_27104 = v_27102 & v_27103;
assign v_27107 = v_27105 & v_27106;
assign v_27110 = v_27108 & v_27109;
assign v_27113 = v_27111 & v_27112;
assign v_27116 = v_27114 & v_27115;
assign v_27119 = v_27117 & v_27118;
assign v_27122 = v_27120 & v_27121;
assign v_27125 = v_27123 & v_27124;
assign v_27128 = v_27126 & v_27127;
assign v_27131 = v_27129 & v_27130;
assign v_27134 = v_27132 & v_27133;
assign v_27137 = v_27135 & v_27136;
assign v_27140 = v_27138 & v_27139;
assign v_27143 = v_27141 & v_27142;
assign v_27146 = v_27144 & v_27145;
assign v_27149 = v_27147 & v_27148;
assign v_27152 = v_27150 & v_27151;
assign v_27155 = v_27153 & v_27154;
assign v_27158 = v_27156 & v_27157;
assign v_27161 = v_27159 & v_27160;
assign v_27164 = v_27162 & v_27163;
assign v_27167 = v_27165 & v_27166;
assign v_27170 = v_27168 & v_27169;
assign v_27173 = v_27171 & v_27172;
assign v_27176 = v_27174 & v_27175;
assign v_27179 = v_27177 & v_27178;
assign v_27182 = v_27180 & v_27181;
assign v_27185 = v_27183 & v_27184;
assign v_27188 = v_27186 & v_27187;
assign v_27191 = v_27189 & v_27190;
assign v_27194 = v_27192 & v_27193;
assign v_27197 = v_27195 & v_27196;
assign v_27200 = v_27198 & v_27199;
assign v_27203 = v_27201 & v_27202;
assign v_27206 = v_27204 & v_27205;
assign v_27209 = v_27207 & v_27208;
assign v_27212 = v_27210 & v_27211;
assign v_27215 = v_27213 & v_27214;
assign v_27218 = v_27216 & v_27217;
assign v_27221 = v_27219 & v_27220;
assign v_27224 = v_27222 & v_27223;
assign v_27227 = v_27225 & v_27226;
assign v_27230 = v_27228 & v_27229;
assign v_27233 = v_27231 & v_27232;
assign v_27236 = v_27234 & v_27235;
assign v_27239 = v_27237 & v_27238;
assign v_27242 = v_27240 & v_27241;
assign v_27243 = v_27053 & v_27242;
assign v_27246 = v_27244 & v_27245;
assign v_27249 = v_27247 & v_27248;
assign v_27252 = v_27250 & v_27251;
assign v_27255 = v_27253 & v_27254;
assign v_27258 = v_27256 & v_27257;
assign v_27261 = v_27259 & v_27260;
assign v_27264 = v_27262 & v_27263;
assign v_27267 = v_27265 & v_27266;
assign v_27270 = v_27268 & v_27269;
assign v_27273 = v_27271 & v_27272;
assign v_27276 = v_27274 & v_27275;
assign v_27279 = v_27277 & v_27278;
assign v_27282 = v_27280 & v_27281;
assign v_27285 = v_27283 & v_27284;
assign v_27288 = v_27286 & v_27287;
assign v_27291 = v_27289 & v_27290;
assign v_27294 = v_27292 & v_27293;
assign v_27297 = v_27295 & v_27296;
assign v_27300 = v_27298 & v_27299;
assign v_27303 = v_27301 & v_27302;
assign v_27306 = v_27304 & v_27305;
assign v_27309 = v_27307 & v_27308;
assign v_27312 = v_27310 & v_27311;
assign v_27315 = v_27313 & v_27314;
assign v_27318 = v_27316 & v_27317;
assign v_27321 = v_27319 & v_27320;
assign v_27324 = v_27322 & v_27323;
assign v_27327 = v_27325 & v_27326;
assign v_27330 = v_27328 & v_27329;
assign v_27333 = v_27331 & v_27332;
assign v_27336 = v_27334 & v_27335;
assign v_27339 = v_27337 & v_27338;
assign v_27342 = v_27340 & v_27341;
assign v_27345 = v_27343 & v_27344;
assign v_27348 = v_27346 & v_27347;
assign v_27351 = v_27349 & v_27350;
assign v_27354 = v_27352 & v_27353;
assign v_27357 = v_27355 & v_27356;
assign v_27360 = v_27358 & v_27359;
assign v_27363 = v_27361 & v_27362;
assign v_27366 = v_27364 & v_27365;
assign v_27369 = v_27367 & v_27368;
assign v_27372 = v_27370 & v_27371;
assign v_27375 = v_27373 & v_27374;
assign v_27378 = v_27376 & v_27377;
assign v_27381 = v_27379 & v_27380;
assign v_27384 = v_27382 & v_27383;
assign v_27387 = v_27385 & v_27386;
assign v_27390 = v_27388 & v_27389;
assign v_27393 = v_27391 & v_27392;
assign v_27396 = v_27394 & v_27395;
assign v_27399 = v_27397 & v_27398;
assign v_27402 = v_27400 & v_27401;
assign v_27405 = v_27403 & v_27404;
assign v_27408 = v_27406 & v_27407;
assign v_27411 = v_27409 & v_27410;
assign v_27414 = v_27412 & v_27413;
assign v_27417 = v_27415 & v_27416;
assign v_27420 = v_27418 & v_27419;
assign v_27423 = v_27421 & v_27422;
assign v_27426 = v_27424 & v_27425;
assign v_27429 = v_27427 & v_27428;
assign v_27432 = v_27430 & v_27431;
assign v_27433 = v_27243 & v_27432;
assign v_27436 = v_27434 & v_27435;
assign v_27439 = v_27437 & v_27438;
assign v_27442 = v_27440 & v_27441;
assign v_27445 = v_27443 & v_27444;
assign v_27448 = v_27446 & v_27447;
assign v_27451 = v_27449 & v_27450;
assign v_27454 = v_27452 & v_27453;
assign v_27457 = v_27455 & v_27456;
assign v_27460 = v_27458 & v_27459;
assign v_27463 = v_27461 & v_27462;
assign v_27466 = v_27464 & v_27465;
assign v_27469 = v_27467 & v_27468;
assign v_27472 = v_27470 & v_27471;
assign v_27475 = v_27473 & v_27474;
assign v_27478 = v_27476 & v_27477;
assign v_27481 = v_27479 & v_27480;
assign v_27484 = v_27482 & v_27483;
assign v_27487 = v_27485 & v_27486;
assign v_27490 = v_27488 & v_27489;
assign v_27493 = v_27491 & v_27492;
assign v_27496 = v_27494 & v_27495;
assign v_27499 = v_27497 & v_27498;
assign v_27502 = v_27500 & v_27501;
assign v_27505 = v_27503 & v_27504;
assign v_27508 = v_27506 & v_27507;
assign v_27511 = v_27509 & v_27510;
assign v_27514 = v_27512 & v_27513;
assign v_27517 = v_27515 & v_27516;
assign v_27520 = v_27518 & v_27519;
assign v_27523 = v_27521 & v_27522;
assign v_27526 = v_27524 & v_27525;
assign v_27529 = v_27527 & v_27528;
assign v_27532 = v_27530 & v_27531;
assign v_27535 = v_27533 & v_27534;
assign v_27538 = v_27536 & v_27537;
assign v_27541 = v_27539 & v_27540;
assign v_27544 = v_27542 & v_27543;
assign v_27547 = v_27545 & v_27546;
assign v_27550 = v_27548 & v_27549;
assign v_27553 = v_27551 & v_27552;
assign v_27556 = v_27554 & v_27555;
assign v_27559 = v_27557 & v_27558;
assign v_27562 = v_27560 & v_27561;
assign v_27565 = v_27563 & v_27564;
assign v_27568 = v_27566 & v_27567;
assign v_27571 = v_27569 & v_27570;
assign v_27574 = v_27572 & v_27573;
assign v_27577 = v_27575 & v_27576;
assign v_27580 = v_27578 & v_27579;
assign v_27583 = v_27581 & v_27582;
assign v_27586 = v_27584 & v_27585;
assign v_27589 = v_27587 & v_27588;
assign v_27592 = v_27590 & v_27591;
assign v_27595 = v_27593 & v_27594;
assign v_27598 = v_27596 & v_27597;
assign v_27601 = v_27599 & v_27600;
assign v_27604 = v_27602 & v_27603;
assign v_27607 = v_27605 & v_27606;
assign v_27610 = v_27608 & v_27609;
assign v_27613 = v_27611 & v_27612;
assign v_27616 = v_27614 & v_27615;
assign v_27619 = v_27617 & v_27618;
assign v_27622 = v_27620 & v_27621;
assign v_27623 = v_27433 & v_27622;
assign v_27626 = v_27624 & v_27625;
assign v_27629 = v_27627 & v_27628;
assign v_27632 = v_27630 & v_27631;
assign v_27635 = v_27633 & v_27634;
assign v_27638 = v_27636 & v_27637;
assign v_27641 = v_27639 & v_27640;
assign v_27644 = v_27642 & v_27643;
assign v_27647 = v_27645 & v_27646;
assign v_27650 = v_27648 & v_27649;
assign v_27653 = v_27651 & v_27652;
assign v_27656 = v_27654 & v_27655;
assign v_27659 = v_27657 & v_27658;
assign v_27662 = v_27660 & v_27661;
assign v_27665 = v_27663 & v_27664;
assign v_27668 = v_27666 & v_27667;
assign v_27671 = v_27669 & v_27670;
assign v_27674 = v_27672 & v_27673;
assign v_27677 = v_27675 & v_27676;
assign v_27680 = v_27678 & v_27679;
assign v_27683 = v_27681 & v_27682;
assign v_27686 = v_27684 & v_27685;
assign v_27689 = v_27687 & v_27688;
assign v_27692 = v_27690 & v_27691;
assign v_27695 = v_27693 & v_27694;
assign v_27698 = v_27696 & v_27697;
assign v_27701 = v_27699 & v_27700;
assign v_27704 = v_27702 & v_27703;
assign v_27707 = v_27705 & v_27706;
assign v_27710 = v_27708 & v_27709;
assign v_27713 = v_27711 & v_27712;
assign v_27716 = v_27714 & v_27715;
assign v_27719 = v_27717 & v_27718;
assign v_27722 = v_27720 & v_27721;
assign v_27725 = v_27723 & v_27724;
assign v_27728 = v_27726 & v_27727;
assign v_27731 = v_27729 & v_27730;
assign v_27734 = v_27732 & v_27733;
assign v_27737 = v_27735 & v_27736;
assign v_27740 = v_27738 & v_27739;
assign v_27743 = v_27741 & v_27742;
assign v_27746 = v_27744 & v_27745;
assign v_27749 = v_27747 & v_27748;
assign v_27752 = v_27750 & v_27751;
assign v_27755 = v_27753 & v_27754;
assign v_27758 = v_27756 & v_27757;
assign v_27761 = v_27759 & v_27760;
assign v_27764 = v_27762 & v_27763;
assign v_27767 = v_27765 & v_27766;
assign v_27770 = v_27768 & v_27769;
assign v_27773 = v_27771 & v_27772;
assign v_27776 = v_27774 & v_27775;
assign v_27779 = v_27777 & v_27778;
assign v_27782 = v_27780 & v_27781;
assign v_27785 = v_27783 & v_27784;
assign v_27788 = v_27786 & v_27787;
assign v_27791 = v_27789 & v_27790;
assign v_27794 = v_27792 & v_27793;
assign v_27797 = v_27795 & v_27796;
assign v_27800 = v_27798 & v_27799;
assign v_27803 = v_27801 & v_27802;
assign v_27806 = v_27804 & v_27805;
assign v_27809 = v_27807 & v_27808;
assign v_27812 = v_27810 & v_27811;
assign v_27813 = v_27623 & v_27812;
assign v_27816 = v_27814 & v_27815;
assign v_27819 = v_27817 & v_27818;
assign v_27822 = v_27820 & v_27821;
assign v_27825 = v_27823 & v_27824;
assign v_27828 = v_27826 & v_27827;
assign v_27831 = v_27829 & v_27830;
assign v_27834 = v_27832 & v_27833;
assign v_27837 = v_27835 & v_27836;
assign v_27840 = v_27838 & v_27839;
assign v_27843 = v_27841 & v_27842;
assign v_27846 = v_27844 & v_27845;
assign v_27849 = v_27847 & v_27848;
assign v_27852 = v_27850 & v_27851;
assign v_27855 = v_27853 & v_27854;
assign v_27858 = v_27856 & v_27857;
assign v_27861 = v_27859 & v_27860;
assign v_27864 = v_27862 & v_27863;
assign v_27867 = v_27865 & v_27866;
assign v_27870 = v_27868 & v_27869;
assign v_27873 = v_27871 & v_27872;
assign v_27876 = v_27874 & v_27875;
assign v_27879 = v_27877 & v_27878;
assign v_27882 = v_27880 & v_27881;
assign v_27885 = v_27883 & v_27884;
assign v_27888 = v_27886 & v_27887;
assign v_27891 = v_27889 & v_27890;
assign v_27894 = v_27892 & v_27893;
assign v_27897 = v_27895 & v_27896;
assign v_27900 = v_27898 & v_27899;
assign v_27903 = v_27901 & v_27902;
assign v_27906 = v_27904 & v_27905;
assign v_27909 = v_27907 & v_27908;
assign v_27912 = v_27910 & v_27911;
assign v_27915 = v_27913 & v_27914;
assign v_27918 = v_27916 & v_27917;
assign v_27921 = v_27919 & v_27920;
assign v_27924 = v_27922 & v_27923;
assign v_27927 = v_27925 & v_27926;
assign v_27930 = v_27928 & v_27929;
assign v_27933 = v_27931 & v_27932;
assign v_27936 = v_27934 & v_27935;
assign v_27939 = v_27937 & v_27938;
assign v_27942 = v_27940 & v_27941;
assign v_27945 = v_27943 & v_27944;
assign v_27948 = v_27946 & v_27947;
assign v_27951 = v_27949 & v_27950;
assign v_27954 = v_27952 & v_27953;
assign v_27957 = v_27955 & v_27956;
assign v_27960 = v_27958 & v_27959;
assign v_27963 = v_27961 & v_27962;
assign v_27966 = v_27964 & v_27965;
assign v_27969 = v_27967 & v_27968;
assign v_27972 = v_27970 & v_27971;
assign v_27975 = v_27973 & v_27974;
assign v_27978 = v_27976 & v_27977;
assign v_27981 = v_27979 & v_27980;
assign v_27984 = v_27982 & v_27983;
assign v_27987 = v_27985 & v_27986;
assign v_27990 = v_27988 & v_27989;
assign v_27993 = v_27991 & v_27992;
assign v_27996 = v_27994 & v_27995;
assign v_27999 = v_27997 & v_27998;
assign v_28002 = v_28000 & v_28001;
assign v_28005 = v_28003 & v_28004;
assign v_28008 = v_28006 & v_28007;
assign v_28011 = v_28009 & v_28010;
assign v_28014 = v_28012 & v_28013;
assign v_28017 = v_28015 & v_28016;
assign v_28020 = v_28018 & v_28019;
assign v_28023 = v_28021 & v_28022;
assign v_28026 = v_28024 & v_28025;
assign v_28029 = v_28027 & v_28028;
assign v_28032 = v_28030 & v_28031;
assign v_28035 = v_28033 & v_28034;
assign v_28038 = v_28036 & v_28037;
assign v_28041 = v_28039 & v_28040;
assign v_28044 = v_28042 & v_28043;
assign v_28047 = v_28045 & v_28046;
assign v_28050 = v_28048 & v_28049;
assign v_28053 = v_28051 & v_28052;
assign v_28056 = v_28054 & v_28055;
assign v_28059 = v_28057 & v_28058;
assign v_28062 = v_28060 & v_28061;
assign v_28065 = v_28063 & v_28064;
assign v_28068 = v_28066 & v_28067;
assign v_28071 = v_28069 & v_28070;
assign v_28074 = v_28072 & v_28073;
assign v_28077 = v_28075 & v_28076;
assign v_28080 = v_28078 & v_28079;
assign v_28083 = v_28081 & v_28082;
assign v_28086 = v_28084 & v_28085;
assign v_28089 = v_28087 & v_28088;
assign v_28092 = v_28090 & v_28091;
assign v_28095 = v_28093 & v_28094;
assign v_28098 = v_28096 & v_28097;
assign v_28101 = v_28099 & v_28100;
assign v_28104 = v_28102 & v_28103;
assign v_28107 = v_28105 & v_28106;
assign v_28110 = v_28108 & v_28109;
assign v_28113 = v_28111 & v_28112;
assign v_28116 = v_28114 & v_28115;
assign v_28119 = v_28117 & v_28118;
assign v_28122 = v_28120 & v_28121;
assign v_28125 = v_28123 & v_28124;
assign v_28128 = v_28126 & v_28127;
assign v_28131 = v_28129 & v_28130;
assign v_28134 = v_28132 & v_28133;
assign v_28137 = v_28135 & v_28136;
assign v_28140 = v_28138 & v_28139;
assign v_28143 = v_28141 & v_28142;
assign v_28146 = v_28144 & v_28145;
assign v_28149 = v_28147 & v_28148;
assign v_28152 = v_28150 & v_28151;
assign v_28155 = v_28153 & v_28154;
assign v_28158 = v_28156 & v_28157;
assign v_28161 = v_28159 & v_28160;
assign v_28164 = v_28162 & v_28163;
assign v_28167 = v_28165 & v_28166;
assign v_28170 = v_28168 & v_28169;
assign v_28173 = v_28171 & v_28172;
assign v_28176 = v_28174 & v_28175;
assign v_28179 = v_28177 & v_28178;
assign v_28182 = v_28180 & v_28181;
assign v_28185 = v_28183 & v_28184;
assign v_28188 = v_28186 & v_28187;
assign v_28191 = v_28189 & v_28190;
assign v_28192 = v_28002 & v_28191;
assign v_28195 = v_28193 & v_28194;
assign v_28198 = v_28196 & v_28197;
assign v_28201 = v_28199 & v_28200;
assign v_28204 = v_28202 & v_28203;
assign v_28207 = v_28205 & v_28206;
assign v_28210 = v_28208 & v_28209;
assign v_28213 = v_28211 & v_28212;
assign v_28216 = v_28214 & v_28215;
assign v_28219 = v_28217 & v_28218;
assign v_28222 = v_28220 & v_28221;
assign v_28225 = v_28223 & v_28224;
assign v_28228 = v_28226 & v_28227;
assign v_28231 = v_28229 & v_28230;
assign v_28234 = v_28232 & v_28233;
assign v_28237 = v_28235 & v_28236;
assign v_28240 = v_28238 & v_28239;
assign v_28243 = v_28241 & v_28242;
assign v_28246 = v_28244 & v_28245;
assign v_28249 = v_28247 & v_28248;
assign v_28252 = v_28250 & v_28251;
assign v_28255 = v_28253 & v_28254;
assign v_28258 = v_28256 & v_28257;
assign v_28261 = v_28259 & v_28260;
assign v_28264 = v_28262 & v_28263;
assign v_28267 = v_28265 & v_28266;
assign v_28270 = v_28268 & v_28269;
assign v_28273 = v_28271 & v_28272;
assign v_28276 = v_28274 & v_28275;
assign v_28279 = v_28277 & v_28278;
assign v_28282 = v_28280 & v_28281;
assign v_28285 = v_28283 & v_28284;
assign v_28288 = v_28286 & v_28287;
assign v_28291 = v_28289 & v_28290;
assign v_28294 = v_28292 & v_28293;
assign v_28297 = v_28295 & v_28296;
assign v_28300 = v_28298 & v_28299;
assign v_28303 = v_28301 & v_28302;
assign v_28306 = v_28304 & v_28305;
assign v_28309 = v_28307 & v_28308;
assign v_28312 = v_28310 & v_28311;
assign v_28315 = v_28313 & v_28314;
assign v_28318 = v_28316 & v_28317;
assign v_28321 = v_28319 & v_28320;
assign v_28324 = v_28322 & v_28323;
assign v_28327 = v_28325 & v_28326;
assign v_28330 = v_28328 & v_28329;
assign v_28333 = v_28331 & v_28332;
assign v_28336 = v_28334 & v_28335;
assign v_28339 = v_28337 & v_28338;
assign v_28342 = v_28340 & v_28341;
assign v_28345 = v_28343 & v_28344;
assign v_28348 = v_28346 & v_28347;
assign v_28351 = v_28349 & v_28350;
assign v_28354 = v_28352 & v_28353;
assign v_28357 = v_28355 & v_28356;
assign v_28360 = v_28358 & v_28359;
assign v_28363 = v_28361 & v_28362;
assign v_28366 = v_28364 & v_28365;
assign v_28369 = v_28367 & v_28368;
assign v_28372 = v_28370 & v_28371;
assign v_28375 = v_28373 & v_28374;
assign v_28378 = v_28376 & v_28377;
assign v_28381 = v_28379 & v_28380;
assign v_28382 = v_28192 & v_28381;
assign v_28385 = v_28383 & v_28384;
assign v_28388 = v_28386 & v_28387;
assign v_28391 = v_28389 & v_28390;
assign v_28394 = v_28392 & v_28393;
assign v_28397 = v_28395 & v_28396;
assign v_28400 = v_28398 & v_28399;
assign v_28403 = v_28401 & v_28402;
assign v_28406 = v_28404 & v_28405;
assign v_28409 = v_28407 & v_28408;
assign v_28412 = v_28410 & v_28411;
assign v_28415 = v_28413 & v_28414;
assign v_28418 = v_28416 & v_28417;
assign v_28421 = v_28419 & v_28420;
assign v_28424 = v_28422 & v_28423;
assign v_28427 = v_28425 & v_28426;
assign v_28430 = v_28428 & v_28429;
assign v_28433 = v_28431 & v_28432;
assign v_28436 = v_28434 & v_28435;
assign v_28439 = v_28437 & v_28438;
assign v_28442 = v_28440 & v_28441;
assign v_28445 = v_28443 & v_28444;
assign v_28448 = v_28446 & v_28447;
assign v_28451 = v_28449 & v_28450;
assign v_28454 = v_28452 & v_28453;
assign v_28457 = v_28455 & v_28456;
assign v_28460 = v_28458 & v_28459;
assign v_28463 = v_28461 & v_28462;
assign v_28466 = v_28464 & v_28465;
assign v_28469 = v_28467 & v_28468;
assign v_28472 = v_28470 & v_28471;
assign v_28475 = v_28473 & v_28474;
assign v_28478 = v_28476 & v_28477;
assign v_28481 = v_28479 & v_28480;
assign v_28484 = v_28482 & v_28483;
assign v_28487 = v_28485 & v_28486;
assign v_28490 = v_28488 & v_28489;
assign v_28493 = v_28491 & v_28492;
assign v_28496 = v_28494 & v_28495;
assign v_28499 = v_28497 & v_28498;
assign v_28502 = v_28500 & v_28501;
assign v_28505 = v_28503 & v_28504;
assign v_28508 = v_28506 & v_28507;
assign v_28511 = v_28509 & v_28510;
assign v_28514 = v_28512 & v_28513;
assign v_28517 = v_28515 & v_28516;
assign v_28520 = v_28518 & v_28519;
assign v_28523 = v_28521 & v_28522;
assign v_28526 = v_28524 & v_28525;
assign v_28529 = v_28527 & v_28528;
assign v_28532 = v_28530 & v_28531;
assign v_28535 = v_28533 & v_28534;
assign v_28538 = v_28536 & v_28537;
assign v_28541 = v_28539 & v_28540;
assign v_28544 = v_28542 & v_28543;
assign v_28547 = v_28545 & v_28546;
assign v_28550 = v_28548 & v_28549;
assign v_28553 = v_28551 & v_28552;
assign v_28556 = v_28554 & v_28555;
assign v_28559 = v_28557 & v_28558;
assign v_28562 = v_28560 & v_28561;
assign v_28565 = v_28563 & v_28564;
assign v_28568 = v_28566 & v_28567;
assign v_28571 = v_28569 & v_28570;
assign v_28572 = v_28382 & v_28571;
assign v_28575 = v_28573 & v_28574;
assign v_28578 = v_28576 & v_28577;
assign v_28581 = v_28579 & v_28580;
assign v_28584 = v_28582 & v_28583;
assign v_28587 = v_28585 & v_28586;
assign v_28590 = v_28588 & v_28589;
assign v_28593 = v_28591 & v_28592;
assign v_28596 = v_28594 & v_28595;
assign v_28599 = v_28597 & v_28598;
assign v_28602 = v_28600 & v_28601;
assign v_28605 = v_28603 & v_28604;
assign v_28608 = v_28606 & v_28607;
assign v_28611 = v_28609 & v_28610;
assign v_28614 = v_28612 & v_28613;
assign v_28617 = v_28615 & v_28616;
assign v_28620 = v_28618 & v_28619;
assign v_28623 = v_28621 & v_28622;
assign v_28626 = v_28624 & v_28625;
assign v_28629 = v_28627 & v_28628;
assign v_28632 = v_28630 & v_28631;
assign v_28635 = v_28633 & v_28634;
assign v_28638 = v_28636 & v_28637;
assign v_28641 = v_28639 & v_28640;
assign v_28644 = v_28642 & v_28643;
assign v_28647 = v_28645 & v_28646;
assign v_28650 = v_28648 & v_28649;
assign v_28653 = v_28651 & v_28652;
assign v_28656 = v_28654 & v_28655;
assign v_28659 = v_28657 & v_28658;
assign v_28662 = v_28660 & v_28661;
assign v_28665 = v_28663 & v_28664;
assign v_28668 = v_28666 & v_28667;
assign v_28671 = v_28669 & v_28670;
assign v_28674 = v_28672 & v_28673;
assign v_28677 = v_28675 & v_28676;
assign v_28680 = v_28678 & v_28679;
assign v_28683 = v_28681 & v_28682;
assign v_28686 = v_28684 & v_28685;
assign v_28689 = v_28687 & v_28688;
assign v_28692 = v_28690 & v_28691;
assign v_28695 = v_28693 & v_28694;
assign v_28698 = v_28696 & v_28697;
assign v_28701 = v_28699 & v_28700;
assign v_28704 = v_28702 & v_28703;
assign v_28707 = v_28705 & v_28706;
assign v_28710 = v_28708 & v_28709;
assign v_28713 = v_28711 & v_28712;
assign v_28716 = v_28714 & v_28715;
assign v_28719 = v_28717 & v_28718;
assign v_28722 = v_28720 & v_28721;
assign v_28725 = v_28723 & v_28724;
assign v_28728 = v_28726 & v_28727;
assign v_28731 = v_28729 & v_28730;
assign v_28734 = v_28732 & v_28733;
assign v_28737 = v_28735 & v_28736;
assign v_28740 = v_28738 & v_28739;
assign v_28743 = v_28741 & v_28742;
assign v_28746 = v_28744 & v_28745;
assign v_28749 = v_28747 & v_28748;
assign v_28752 = v_28750 & v_28751;
assign v_28755 = v_28753 & v_28754;
assign v_28758 = v_28756 & v_28757;
assign v_28761 = v_28759 & v_28760;
assign v_28762 = v_28572 & v_28761;
assign v_28765 = v_28763 & v_28764;
assign v_28768 = v_28766 & v_28767;
assign v_28771 = v_28769 & v_28770;
assign v_28774 = v_28772 & v_28773;
assign v_28777 = v_28775 & v_28776;
assign v_28780 = v_28778 & v_28779;
assign v_28783 = v_28781 & v_28782;
assign v_28786 = v_28784 & v_28785;
assign v_28789 = v_28787 & v_28788;
assign v_28792 = v_28790 & v_28791;
assign v_28795 = v_28793 & v_28794;
assign v_28798 = v_28796 & v_28797;
assign v_28801 = v_28799 & v_28800;
assign v_28804 = v_28802 & v_28803;
assign v_28807 = v_28805 & v_28806;
assign v_28810 = v_28808 & v_28809;
assign v_28813 = v_28811 & v_28812;
assign v_28816 = v_28814 & v_28815;
assign v_28819 = v_28817 & v_28818;
assign v_28822 = v_28820 & v_28821;
assign v_28825 = v_28823 & v_28824;
assign v_28828 = v_28826 & v_28827;
assign v_28831 = v_28829 & v_28830;
assign v_28834 = v_28832 & v_28833;
assign v_28837 = v_28835 & v_28836;
assign v_28840 = v_28838 & v_28839;
assign v_28843 = v_28841 & v_28842;
assign v_28846 = v_28844 & v_28845;
assign v_28849 = v_28847 & v_28848;
assign v_28852 = v_28850 & v_28851;
assign v_28855 = v_28853 & v_28854;
assign v_28858 = v_28856 & v_28857;
assign v_28861 = v_28859 & v_28860;
assign v_28864 = v_28862 & v_28863;
assign v_28867 = v_28865 & v_28866;
assign v_28870 = v_28868 & v_28869;
assign v_28873 = v_28871 & v_28872;
assign v_28876 = v_28874 & v_28875;
assign v_28879 = v_28877 & v_28878;
assign v_28882 = v_28880 & v_28881;
assign v_28885 = v_28883 & v_28884;
assign v_28888 = v_28886 & v_28887;
assign v_28891 = v_28889 & v_28890;
assign v_28894 = v_28892 & v_28893;
assign v_28897 = v_28895 & v_28896;
assign v_28900 = v_28898 & v_28899;
assign v_28903 = v_28901 & v_28902;
assign v_28906 = v_28904 & v_28905;
assign v_28909 = v_28907 & v_28908;
assign v_28912 = v_28910 & v_28911;
assign v_28915 = v_28913 & v_28914;
assign v_28918 = v_28916 & v_28917;
assign v_28921 = v_28919 & v_28920;
assign v_28924 = v_28922 & v_28923;
assign v_28927 = v_28925 & v_28926;
assign v_28930 = v_28928 & v_28929;
assign v_28933 = v_28931 & v_28932;
assign v_28936 = v_28934 & v_28935;
assign v_28939 = v_28937 & v_28938;
assign v_28942 = v_28940 & v_28941;
assign v_28945 = v_28943 & v_28944;
assign v_28948 = v_28946 & v_28947;
assign v_28951 = v_28949 & v_28950;
assign v_28952 = v_28762 & v_28951;
assign v_28953 = v_22981 & v_28952;
assign v_28956 = v_28954 & v_28955;
assign v_28959 = v_28957 & v_28958;
assign v_28962 = v_28960 & v_28961;
assign v_28965 = v_28963 & v_28964;
assign v_28968 = v_28966 & v_28967;
assign v_28971 = v_28969 & v_28970;
assign v_28974 = v_28972 & v_28973;
assign v_28977 = v_28975 & v_28976;
assign v_28980 = v_28978 & v_28979;
assign v_28983 = v_28981 & v_28982;
assign v_28986 = v_28984 & v_28985;
assign v_28989 = v_28987 & v_28988;
assign v_28992 = v_28990 & v_28991;
assign v_28995 = v_28993 & v_28994;
assign v_28998 = v_28996 & v_28997;
assign v_29001 = v_28999 & v_29000;
assign v_29004 = v_29002 & v_29003;
assign v_29007 = v_29005 & v_29006;
assign v_29010 = v_29008 & v_29009;
assign v_29013 = v_29011 & v_29012;
assign v_29016 = v_29014 & v_29015;
assign v_29019 = v_29017 & v_29018;
assign v_29022 = v_29020 & v_29021;
assign v_29025 = v_29023 & v_29024;
assign v_29028 = v_29026 & v_29027;
assign v_29031 = v_29029 & v_29030;
assign v_29034 = v_29032 & v_29033;
assign v_29037 = v_29035 & v_29036;
assign v_29040 = v_29038 & v_29039;
assign v_29043 = v_29041 & v_29042;
assign v_29046 = v_29044 & v_29045;
assign v_29049 = v_29047 & v_29048;
assign v_29052 = v_29050 & v_29051;
assign v_29055 = v_29053 & v_29054;
assign v_29058 = v_29056 & v_29057;
assign v_29061 = v_29059 & v_29060;
assign v_29064 = v_29062 & v_29063;
assign v_29067 = v_29065 & v_29066;
assign v_29070 = v_29068 & v_29069;
assign v_29073 = v_29071 & v_29072;
assign v_29076 = v_29074 & v_29075;
assign v_29079 = v_29077 & v_29078;
assign v_29082 = v_29080 & v_29081;
assign v_29085 = v_29083 & v_29084;
assign v_29088 = v_29086 & v_29087;
assign v_29091 = v_29089 & v_29090;
assign v_29094 = v_29092 & v_29093;
assign v_29097 = v_29095 & v_29096;
assign v_29100 = v_29098 & v_29099;
assign v_29103 = v_29101 & v_29102;
assign v_29106 = v_29104 & v_29105;
assign v_29109 = v_29107 & v_29108;
assign v_29112 = v_29110 & v_29111;
assign v_29115 = v_29113 & v_29114;
assign v_29118 = v_29116 & v_29117;
assign v_29121 = v_29119 & v_29120;
assign v_29124 = v_29122 & v_29123;
assign v_29127 = v_29125 & v_29126;
assign v_29130 = v_29128 & v_29129;
assign v_29133 = v_29131 & v_29132;
assign v_29136 = v_29134 & v_29135;
assign v_29139 = v_29137 & v_29138;
assign v_29142 = v_29140 & v_29141;
assign v_29143 = v_28953 & v_29142;
assign v_29144 = v_26290 & v_29143;
assign v_29145 = v_27813 & v_29144;
assign v_29146 = ~v_10462 & v_29145;
assign v_29150 = v_29148 & v_29149;
assign v_29153 = v_29151 & v_29152;
assign v_29156 = v_29154 & v_29155;
assign v_29159 = v_29157 & v_29158;
assign v_29162 = v_29160 & v_29161;
assign v_29165 = v_29163 & v_29164;
assign v_29168 = v_29166 & v_29167;
assign v_29171 = v_29169 & v_29170;
assign v_29174 = v_29172 & v_29173;
assign v_29177 = v_29175 & v_29176;
assign v_29180 = v_29178 & v_29179;
assign v_29183 = v_29181 & v_29182;
assign v_29186 = v_29184 & v_29185;
assign v_29189 = v_29187 & v_29188;
assign v_29192 = v_29190 & v_29191;
assign v_29195 = v_29193 & v_29194;
assign v_29198 = v_29196 & v_29197;
assign v_29201 = v_29199 & v_29200;
assign v_29204 = v_29202 & v_29203;
assign v_29207 = v_29205 & v_29206;
assign v_29210 = v_29208 & v_29209;
assign v_29213 = v_29211 & v_29212;
assign v_29216 = v_29214 & v_29215;
assign v_29219 = v_29217 & v_29218;
assign v_29222 = v_29220 & v_29221;
assign v_29225 = v_29223 & v_29224;
assign v_29228 = v_29226 & v_29227;
assign v_29231 = v_29229 & v_29230;
assign v_29234 = v_29232 & v_29233;
assign v_29237 = v_29235 & v_29236;
assign v_29240 = v_29238 & v_29239;
assign v_29243 = v_29241 & v_29242;
assign v_29246 = v_29244 & v_29245;
assign v_29249 = v_29247 & v_29248;
assign v_29252 = v_29250 & v_29251;
assign v_29255 = v_29253 & v_29254;
assign v_29258 = v_29256 & v_29257;
assign v_29261 = v_29259 & v_29260;
assign v_29264 = v_29262 & v_29263;
assign v_29267 = v_29265 & v_29266;
assign v_29270 = v_29268 & v_29269;
assign v_29273 = v_29271 & v_29272;
assign v_29276 = v_29274 & v_29275;
assign v_29279 = v_29277 & v_29278;
assign v_29282 = v_29280 & v_29281;
assign v_29285 = v_29283 & v_29284;
assign v_29288 = v_29286 & v_29287;
assign v_29291 = v_29289 & v_29290;
assign v_29294 = v_29292 & v_29293;
assign v_29297 = v_29295 & v_29296;
assign v_29300 = v_29298 & v_29299;
assign v_29303 = v_29301 & v_29302;
assign v_29306 = v_29304 & v_29305;
assign v_29309 = v_29307 & v_29308;
assign v_29312 = v_29310 & v_29311;
assign v_29315 = v_29313 & v_29314;
assign v_29318 = v_29316 & v_29317;
assign v_29321 = v_29319 & v_29320;
assign v_29324 = v_29322 & v_29323;
assign v_29327 = v_29325 & v_29326;
assign v_29330 = v_29328 & v_29329;
assign v_29333 = v_29331 & v_29332;
assign v_29336 = v_29334 & v_29335;
assign v_29339 = v_29337 & v_29338;
assign v_29342 = v_29340 & v_29341;
assign v_29345 = v_29343 & v_29344;
assign v_29348 = v_29346 & v_29347;
assign v_29351 = v_29349 & v_29350;
assign v_29354 = v_29352 & v_29353;
assign v_29357 = v_29355 & v_29356;
assign v_29360 = v_29358 & v_29359;
assign v_29363 = v_29361 & v_29362;
assign v_29366 = v_29364 & v_29365;
assign v_29369 = v_29367 & v_29368;
assign v_29372 = v_29370 & v_29371;
assign v_29375 = v_29373 & v_29374;
assign v_29378 = v_29376 & v_29377;
assign v_29381 = v_29379 & v_29380;
assign v_29384 = v_29382 & v_29383;
assign v_29387 = v_29385 & v_29386;
assign v_29390 = v_29388 & v_29389;
assign v_29393 = v_29391 & v_29392;
assign v_29396 = v_29394 & v_29395;
assign v_29399 = v_29397 & v_29398;
assign v_29402 = v_29400 & v_29401;
assign v_29405 = v_29403 & v_29404;
assign v_29408 = v_29406 & v_29407;
assign v_29411 = v_29409 & v_29410;
assign v_29414 = v_29412 & v_29413;
assign v_29417 = v_29415 & v_29416;
assign v_29420 = v_29418 & v_29419;
assign v_29423 = v_29421 & v_29422;
assign v_29426 = v_29424 & v_29425;
assign v_29429 = v_29427 & v_29428;
assign v_29432 = v_29430 & v_29431;
assign v_29435 = v_29433 & v_29434;
assign v_29438 = v_29436 & v_29437;
assign v_29441 = v_29439 & v_29440;
assign v_29444 = v_29442 & v_29443;
assign v_29447 = v_29445 & v_29446;
assign v_29450 = v_29448 & v_29449;
assign v_29453 = v_29451 & v_29452;
assign v_29456 = v_29454 & v_29455;
assign v_29459 = v_29457 & v_29458;
assign v_29462 = v_29460 & v_29461;
assign v_29465 = v_29463 & v_29464;
assign v_29468 = v_29466 & v_29467;
assign v_29471 = v_29469 & v_29470;
assign v_29474 = v_29472 & v_29473;
assign v_29477 = v_29475 & v_29476;
assign v_29480 = v_29478 & v_29479;
assign v_29483 = v_29481 & v_29482;
assign v_29486 = v_29484 & v_29485;
assign v_29489 = v_29487 & v_29488;
assign v_29492 = v_29490 & v_29491;
assign v_29495 = v_29493 & v_29494;
assign v_29498 = v_29496 & v_29497;
assign v_29501 = v_29499 & v_29500;
assign v_29504 = v_29502 & v_29503;
assign v_29507 = v_29505 & v_29506;
assign v_29510 = v_29508 & v_29509;
assign v_29513 = v_29511 & v_29512;
assign v_29514 = v_29330 & v_29513;
assign v_29517 = v_29515 & v_29516;
assign v_29520 = v_29518 & v_29519;
assign v_29523 = v_29521 & v_29522;
assign v_29526 = v_29524 & v_29525;
assign v_29529 = v_29527 & v_29528;
assign v_29532 = v_29530 & v_29531;
assign v_29535 = v_29533 & v_29534;
assign v_29538 = v_29536 & v_29537;
assign v_29541 = v_29539 & v_29540;
assign v_29544 = v_29542 & v_29543;
assign v_29547 = v_29545 & v_29546;
assign v_29550 = v_29548 & v_29549;
assign v_29553 = v_29551 & v_29552;
assign v_29556 = v_29554 & v_29555;
assign v_29559 = v_29557 & v_29558;
assign v_29562 = v_29560 & v_29561;
assign v_29565 = v_29563 & v_29564;
assign v_29568 = v_29566 & v_29567;
assign v_29571 = v_29569 & v_29570;
assign v_29574 = v_29572 & v_29573;
assign v_29577 = v_29575 & v_29576;
assign v_29580 = v_29578 & v_29579;
assign v_29583 = v_29581 & v_29582;
assign v_29586 = v_29584 & v_29585;
assign v_29589 = v_29587 & v_29588;
assign v_29592 = v_29590 & v_29591;
assign v_29595 = v_29593 & v_29594;
assign v_29598 = v_29596 & v_29597;
assign v_29601 = v_29599 & v_29600;
assign v_29604 = v_29602 & v_29603;
assign v_29607 = v_29605 & v_29606;
assign v_29610 = v_29608 & v_29609;
assign v_29613 = v_29611 & v_29612;
assign v_29616 = v_29614 & v_29615;
assign v_29619 = v_29617 & v_29618;
assign v_29622 = v_29620 & v_29621;
assign v_29625 = v_29623 & v_29624;
assign v_29628 = v_29626 & v_29627;
assign v_29631 = v_29629 & v_29630;
assign v_29634 = v_29632 & v_29633;
assign v_29637 = v_29635 & v_29636;
assign v_29640 = v_29638 & v_29639;
assign v_29643 = v_29641 & v_29642;
assign v_29646 = v_29644 & v_29645;
assign v_29649 = v_29647 & v_29648;
assign v_29652 = v_29650 & v_29651;
assign v_29655 = v_29653 & v_29654;
assign v_29658 = v_29656 & v_29657;
assign v_29661 = v_29659 & v_29660;
assign v_29664 = v_29662 & v_29663;
assign v_29667 = v_29665 & v_29666;
assign v_29670 = v_29668 & v_29669;
assign v_29673 = v_29671 & v_29672;
assign v_29676 = v_29674 & v_29675;
assign v_29679 = v_29677 & v_29678;
assign v_29682 = v_29680 & v_29681;
assign v_29685 = v_29683 & v_29684;
assign v_29688 = v_29686 & v_29687;
assign v_29691 = v_29689 & v_29690;
assign v_29694 = v_29692 & v_29693;
assign v_29697 = v_29695 & v_29696;
assign v_29698 = v_29514 & v_29697;
assign v_29701 = v_29699 & v_29700;
assign v_29704 = v_29702 & v_29703;
assign v_29707 = v_29705 & v_29706;
assign v_29710 = v_29708 & v_29709;
assign v_29713 = v_29711 & v_29712;
assign v_29716 = v_29714 & v_29715;
assign v_29719 = v_29717 & v_29718;
assign v_29722 = v_29720 & v_29721;
assign v_29725 = v_29723 & v_29724;
assign v_29728 = v_29726 & v_29727;
assign v_29731 = v_29729 & v_29730;
assign v_29734 = v_29732 & v_29733;
assign v_29737 = v_29735 & v_29736;
assign v_29740 = v_29738 & v_29739;
assign v_29743 = v_29741 & v_29742;
assign v_29746 = v_29744 & v_29745;
assign v_29749 = v_29747 & v_29748;
assign v_29752 = v_29750 & v_29751;
assign v_29755 = v_29753 & v_29754;
assign v_29758 = v_29756 & v_29757;
assign v_29761 = v_29759 & v_29760;
assign v_29764 = v_29762 & v_29763;
assign v_29767 = v_29765 & v_29766;
assign v_29770 = v_29768 & v_29769;
assign v_29773 = v_29771 & v_29772;
assign v_29776 = v_29774 & v_29775;
assign v_29779 = v_29777 & v_29778;
assign v_29782 = v_29780 & v_29781;
assign v_29785 = v_29783 & v_29784;
assign v_29788 = v_29786 & v_29787;
assign v_29791 = v_29789 & v_29790;
assign v_29794 = v_29792 & v_29793;
assign v_29797 = v_29795 & v_29796;
assign v_29800 = v_29798 & v_29799;
assign v_29803 = v_29801 & v_29802;
assign v_29806 = v_29804 & v_29805;
assign v_29809 = v_29807 & v_29808;
assign v_29812 = v_29810 & v_29811;
assign v_29815 = v_29813 & v_29814;
assign v_29818 = v_29816 & v_29817;
assign v_29821 = v_29819 & v_29820;
assign v_29824 = v_29822 & v_29823;
assign v_29827 = v_29825 & v_29826;
assign v_29830 = v_29828 & v_29829;
assign v_29833 = v_29831 & v_29832;
assign v_29836 = v_29834 & v_29835;
assign v_29839 = v_29837 & v_29838;
assign v_29842 = v_29840 & v_29841;
assign v_29845 = v_29843 & v_29844;
assign v_29848 = v_29846 & v_29847;
assign v_29851 = v_29849 & v_29850;
assign v_29854 = v_29852 & v_29853;
assign v_29857 = v_29855 & v_29856;
assign v_29860 = v_29858 & v_29859;
assign v_29863 = v_29861 & v_29862;
assign v_29866 = v_29864 & v_29865;
assign v_29869 = v_29867 & v_29868;
assign v_29872 = v_29870 & v_29871;
assign v_29875 = v_29873 & v_29874;
assign v_29878 = v_29876 & v_29877;
assign v_29881 = v_29879 & v_29880;
assign v_29882 = v_29698 & v_29881;
assign v_29885 = v_29883 & v_29884;
assign v_29888 = v_29886 & v_29887;
assign v_29891 = v_29889 & v_29890;
assign v_29894 = v_29892 & v_29893;
assign v_29897 = v_29895 & v_29896;
assign v_29900 = v_29898 & v_29899;
assign v_29903 = v_29901 & v_29902;
assign v_29906 = v_29904 & v_29905;
assign v_29909 = v_29907 & v_29908;
assign v_29912 = v_29910 & v_29911;
assign v_29915 = v_29913 & v_29914;
assign v_29918 = v_29916 & v_29917;
assign v_29921 = v_29919 & v_29920;
assign v_29924 = v_29922 & v_29923;
assign v_29927 = v_29925 & v_29926;
assign v_29930 = v_29928 & v_29929;
assign v_29933 = v_29931 & v_29932;
assign v_29936 = v_29934 & v_29935;
assign v_29939 = v_29937 & v_29938;
assign v_29942 = v_29940 & v_29941;
assign v_29945 = v_29943 & v_29944;
assign v_29948 = v_29946 & v_29947;
assign v_29951 = v_29949 & v_29950;
assign v_29954 = v_29952 & v_29953;
assign v_29957 = v_29955 & v_29956;
assign v_29960 = v_29958 & v_29959;
assign v_29963 = v_29961 & v_29962;
assign v_29966 = v_29964 & v_29965;
assign v_29969 = v_29967 & v_29968;
assign v_29972 = v_29970 & v_29971;
assign v_29975 = v_29973 & v_29974;
assign v_29978 = v_29976 & v_29977;
assign v_29981 = v_29979 & v_29980;
assign v_29984 = v_29982 & v_29983;
assign v_29987 = v_29985 & v_29986;
assign v_29990 = v_29988 & v_29989;
assign v_29993 = v_29991 & v_29992;
assign v_29996 = v_29994 & v_29995;
assign v_29999 = v_29997 & v_29998;
assign v_30002 = v_30000 & v_30001;
assign v_30005 = v_30003 & v_30004;
assign v_30008 = v_30006 & v_30007;
assign v_30011 = v_30009 & v_30010;
assign v_30014 = v_30012 & v_30013;
assign v_30017 = v_30015 & v_30016;
assign v_30020 = v_30018 & v_30019;
assign v_30023 = v_30021 & v_30022;
assign v_30026 = v_30024 & v_30025;
assign v_30029 = v_30027 & v_30028;
assign v_30032 = v_30030 & v_30031;
assign v_30035 = v_30033 & v_30034;
assign v_30038 = v_30036 & v_30037;
assign v_30041 = v_30039 & v_30040;
assign v_30044 = v_30042 & v_30043;
assign v_30047 = v_30045 & v_30046;
assign v_30050 = v_30048 & v_30049;
assign v_30053 = v_30051 & v_30052;
assign v_30056 = v_30054 & v_30055;
assign v_30059 = v_30057 & v_30058;
assign v_30062 = v_30060 & v_30061;
assign v_30065 = v_30063 & v_30064;
assign v_30066 = v_29882 & v_30065;
assign v_30069 = v_30067 & v_30068;
assign v_30072 = v_30070 & v_30071;
assign v_30075 = v_30073 & v_30074;
assign v_30078 = v_30076 & v_30077;
assign v_30081 = v_30079 & v_30080;
assign v_30084 = v_30082 & v_30083;
assign v_30087 = v_30085 & v_30086;
assign v_30090 = v_30088 & v_30089;
assign v_30093 = v_30091 & v_30092;
assign v_30096 = v_30094 & v_30095;
assign v_30099 = v_30097 & v_30098;
assign v_30102 = v_30100 & v_30101;
assign v_30105 = v_30103 & v_30104;
assign v_30108 = v_30106 & v_30107;
assign v_30111 = v_30109 & v_30110;
assign v_30114 = v_30112 & v_30113;
assign v_30117 = v_30115 & v_30116;
assign v_30120 = v_30118 & v_30119;
assign v_30123 = v_30121 & v_30122;
assign v_30126 = v_30124 & v_30125;
assign v_30129 = v_30127 & v_30128;
assign v_30132 = v_30130 & v_30131;
assign v_30135 = v_30133 & v_30134;
assign v_30138 = v_30136 & v_30137;
assign v_30141 = v_30139 & v_30140;
assign v_30144 = v_30142 & v_30143;
assign v_30147 = v_30145 & v_30146;
assign v_30150 = v_30148 & v_30149;
assign v_30153 = v_30151 & v_30152;
assign v_30156 = v_30154 & v_30155;
assign v_30159 = v_30157 & v_30158;
assign v_30162 = v_30160 & v_30161;
assign v_30165 = v_30163 & v_30164;
assign v_30168 = v_30166 & v_30167;
assign v_30171 = v_30169 & v_30170;
assign v_30174 = v_30172 & v_30173;
assign v_30177 = v_30175 & v_30176;
assign v_30180 = v_30178 & v_30179;
assign v_30183 = v_30181 & v_30182;
assign v_30186 = v_30184 & v_30185;
assign v_30189 = v_30187 & v_30188;
assign v_30192 = v_30190 & v_30191;
assign v_30195 = v_30193 & v_30194;
assign v_30198 = v_30196 & v_30197;
assign v_30201 = v_30199 & v_30200;
assign v_30204 = v_30202 & v_30203;
assign v_30207 = v_30205 & v_30206;
assign v_30210 = v_30208 & v_30209;
assign v_30213 = v_30211 & v_30212;
assign v_30216 = v_30214 & v_30215;
assign v_30219 = v_30217 & v_30218;
assign v_30222 = v_30220 & v_30221;
assign v_30225 = v_30223 & v_30224;
assign v_30228 = v_30226 & v_30227;
assign v_30231 = v_30229 & v_30230;
assign v_30234 = v_30232 & v_30233;
assign v_30237 = v_30235 & v_30236;
assign v_30240 = v_30238 & v_30239;
assign v_30243 = v_30241 & v_30242;
assign v_30246 = v_30244 & v_30245;
assign v_30249 = v_30247 & v_30248;
assign v_30250 = v_30066 & v_30249;
assign v_30253 = v_30251 & v_30252;
assign v_30256 = v_30254 & v_30255;
assign v_30259 = v_30257 & v_30258;
assign v_30262 = v_30260 & v_30261;
assign v_30265 = v_30263 & v_30264;
assign v_30268 = v_30266 & v_30267;
assign v_30271 = v_30269 & v_30270;
assign v_30274 = v_30272 & v_30273;
assign v_30277 = v_30275 & v_30276;
assign v_30280 = v_30278 & v_30279;
assign v_30283 = v_30281 & v_30282;
assign v_30286 = v_30284 & v_30285;
assign v_30289 = v_30287 & v_30288;
assign v_30292 = v_30290 & v_30291;
assign v_30295 = v_30293 & v_30294;
assign v_30298 = v_30296 & v_30297;
assign v_30301 = v_30299 & v_30300;
assign v_30304 = v_30302 & v_30303;
assign v_30307 = v_30305 & v_30306;
assign v_30310 = v_30308 & v_30309;
assign v_30313 = v_30311 & v_30312;
assign v_30316 = v_30314 & v_30315;
assign v_30319 = v_30317 & v_30318;
assign v_30322 = v_30320 & v_30321;
assign v_30325 = v_30323 & v_30324;
assign v_30328 = v_30326 & v_30327;
assign v_30331 = v_30329 & v_30330;
assign v_30334 = v_30332 & v_30333;
assign v_30337 = v_30335 & v_30336;
assign v_30340 = v_30338 & v_30339;
assign v_30343 = v_30341 & v_30342;
assign v_30346 = v_30344 & v_30345;
assign v_30349 = v_30347 & v_30348;
assign v_30352 = v_30350 & v_30351;
assign v_30355 = v_30353 & v_30354;
assign v_30358 = v_30356 & v_30357;
assign v_30361 = v_30359 & v_30360;
assign v_30364 = v_30362 & v_30363;
assign v_30367 = v_30365 & v_30366;
assign v_30370 = v_30368 & v_30369;
assign v_30373 = v_30371 & v_30372;
assign v_30376 = v_30374 & v_30375;
assign v_30379 = v_30377 & v_30378;
assign v_30382 = v_30380 & v_30381;
assign v_30385 = v_30383 & v_30384;
assign v_30388 = v_30386 & v_30387;
assign v_30391 = v_30389 & v_30390;
assign v_30394 = v_30392 & v_30393;
assign v_30397 = v_30395 & v_30396;
assign v_30400 = v_30398 & v_30399;
assign v_30403 = v_30401 & v_30402;
assign v_30406 = v_30404 & v_30405;
assign v_30409 = v_30407 & v_30408;
assign v_30412 = v_30410 & v_30411;
assign v_30415 = v_30413 & v_30414;
assign v_30418 = v_30416 & v_30417;
assign v_30421 = v_30419 & v_30420;
assign v_30424 = v_30422 & v_30423;
assign v_30427 = v_30425 & v_30426;
assign v_30430 = v_30428 & v_30429;
assign v_30433 = v_30431 & v_30432;
assign v_30434 = v_30250 & v_30433;
assign v_30437 = v_30435 & v_30436;
assign v_30440 = v_30438 & v_30439;
assign v_30443 = v_30441 & v_30442;
assign v_30446 = v_30444 & v_30445;
assign v_30449 = v_30447 & v_30448;
assign v_30452 = v_30450 & v_30451;
assign v_30455 = v_30453 & v_30454;
assign v_30458 = v_30456 & v_30457;
assign v_30461 = v_30459 & v_30460;
assign v_30464 = v_30462 & v_30463;
assign v_30467 = v_30465 & v_30466;
assign v_30470 = v_30468 & v_30469;
assign v_30473 = v_30471 & v_30472;
assign v_30476 = v_30474 & v_30475;
assign v_30479 = v_30477 & v_30478;
assign v_30482 = v_30480 & v_30481;
assign v_30485 = v_30483 & v_30484;
assign v_30488 = v_30486 & v_30487;
assign v_30491 = v_30489 & v_30490;
assign v_30494 = v_30492 & v_30493;
assign v_30497 = v_30495 & v_30496;
assign v_30500 = v_30498 & v_30499;
assign v_30503 = v_30501 & v_30502;
assign v_30506 = v_30504 & v_30505;
assign v_30509 = v_30507 & v_30508;
assign v_30512 = v_30510 & v_30511;
assign v_30515 = v_30513 & v_30514;
assign v_30518 = v_30516 & v_30517;
assign v_30521 = v_30519 & v_30520;
assign v_30524 = v_30522 & v_30523;
assign v_30527 = v_30525 & v_30526;
assign v_30530 = v_30528 & v_30529;
assign v_30533 = v_30531 & v_30532;
assign v_30536 = v_30534 & v_30535;
assign v_30539 = v_30537 & v_30538;
assign v_30542 = v_30540 & v_30541;
assign v_30545 = v_30543 & v_30544;
assign v_30548 = v_30546 & v_30547;
assign v_30551 = v_30549 & v_30550;
assign v_30554 = v_30552 & v_30553;
assign v_30557 = v_30555 & v_30556;
assign v_30560 = v_30558 & v_30559;
assign v_30563 = v_30561 & v_30562;
assign v_30566 = v_30564 & v_30565;
assign v_30569 = v_30567 & v_30568;
assign v_30572 = v_30570 & v_30571;
assign v_30575 = v_30573 & v_30574;
assign v_30578 = v_30576 & v_30577;
assign v_30581 = v_30579 & v_30580;
assign v_30584 = v_30582 & v_30583;
assign v_30587 = v_30585 & v_30586;
assign v_30590 = v_30588 & v_30589;
assign v_30593 = v_30591 & v_30592;
assign v_30596 = v_30594 & v_30595;
assign v_30599 = v_30597 & v_30598;
assign v_30602 = v_30600 & v_30601;
assign v_30605 = v_30603 & v_30604;
assign v_30608 = v_30606 & v_30607;
assign v_30611 = v_30609 & v_30610;
assign v_30614 = v_30612 & v_30613;
assign v_30617 = v_30615 & v_30616;
assign v_30618 = v_30434 & v_30617;
assign v_30621 = v_30619 & v_30620;
assign v_30624 = v_30622 & v_30623;
assign v_30627 = v_30625 & v_30626;
assign v_30630 = v_30628 & v_30629;
assign v_30633 = v_30631 & v_30632;
assign v_30636 = v_30634 & v_30635;
assign v_30639 = v_30637 & v_30638;
assign v_30642 = v_30640 & v_30641;
assign v_30645 = v_30643 & v_30644;
assign v_30648 = v_30646 & v_30647;
assign v_30651 = v_30649 & v_30650;
assign v_30654 = v_30652 & v_30653;
assign v_30657 = v_30655 & v_30656;
assign v_30660 = v_30658 & v_30659;
assign v_30663 = v_30661 & v_30662;
assign v_30666 = v_30664 & v_30665;
assign v_30669 = v_30667 & v_30668;
assign v_30672 = v_30670 & v_30671;
assign v_30675 = v_30673 & v_30674;
assign v_30678 = v_30676 & v_30677;
assign v_30681 = v_30679 & v_30680;
assign v_30684 = v_30682 & v_30683;
assign v_30687 = v_30685 & v_30686;
assign v_30690 = v_30688 & v_30689;
assign v_30693 = v_30691 & v_30692;
assign v_30696 = v_30694 & v_30695;
assign v_30699 = v_30697 & v_30698;
assign v_30702 = v_30700 & v_30701;
assign v_30705 = v_30703 & v_30704;
assign v_30708 = v_30706 & v_30707;
assign v_30711 = v_30709 & v_30710;
assign v_30714 = v_30712 & v_30713;
assign v_30717 = v_30715 & v_30716;
assign v_30720 = v_30718 & v_30719;
assign v_30723 = v_30721 & v_30722;
assign v_30726 = v_30724 & v_30725;
assign v_30729 = v_30727 & v_30728;
assign v_30732 = v_30730 & v_30731;
assign v_30735 = v_30733 & v_30734;
assign v_30738 = v_30736 & v_30737;
assign v_30741 = v_30739 & v_30740;
assign v_30744 = v_30742 & v_30743;
assign v_30747 = v_30745 & v_30746;
assign v_30750 = v_30748 & v_30749;
assign v_30753 = v_30751 & v_30752;
assign v_30756 = v_30754 & v_30755;
assign v_30759 = v_30757 & v_30758;
assign v_30762 = v_30760 & v_30761;
assign v_30765 = v_30763 & v_30764;
assign v_30768 = v_30766 & v_30767;
assign v_30771 = v_30769 & v_30770;
assign v_30774 = v_30772 & v_30773;
assign v_30777 = v_30775 & v_30776;
assign v_30780 = v_30778 & v_30779;
assign v_30783 = v_30781 & v_30782;
assign v_30786 = v_30784 & v_30785;
assign v_30789 = v_30787 & v_30788;
assign v_30792 = v_30790 & v_30791;
assign v_30795 = v_30793 & v_30794;
assign v_30798 = v_30796 & v_30797;
assign v_30801 = v_30799 & v_30800;
assign v_30804 = v_30802 & v_30803;
assign v_30807 = v_30805 & v_30806;
assign v_30810 = v_30808 & v_30809;
assign v_30813 = v_30811 & v_30812;
assign v_30816 = v_30814 & v_30815;
assign v_30819 = v_30817 & v_30818;
assign v_30822 = v_30820 & v_30821;
assign v_30825 = v_30823 & v_30824;
assign v_30828 = v_30826 & v_30827;
assign v_30831 = v_30829 & v_30830;
assign v_30834 = v_30832 & v_30833;
assign v_30837 = v_30835 & v_30836;
assign v_30840 = v_30838 & v_30839;
assign v_30843 = v_30841 & v_30842;
assign v_30846 = v_30844 & v_30845;
assign v_30849 = v_30847 & v_30848;
assign v_30852 = v_30850 & v_30851;
assign v_30855 = v_30853 & v_30854;
assign v_30858 = v_30856 & v_30857;
assign v_30861 = v_30859 & v_30860;
assign v_30864 = v_30862 & v_30863;
assign v_30867 = v_30865 & v_30866;
assign v_30870 = v_30868 & v_30869;
assign v_30873 = v_30871 & v_30872;
assign v_30876 = v_30874 & v_30875;
assign v_30879 = v_30877 & v_30878;
assign v_30882 = v_30880 & v_30881;
assign v_30885 = v_30883 & v_30884;
assign v_30888 = v_30886 & v_30887;
assign v_30891 = v_30889 & v_30890;
assign v_30894 = v_30892 & v_30893;
assign v_30897 = v_30895 & v_30896;
assign v_30900 = v_30898 & v_30899;
assign v_30903 = v_30901 & v_30902;
assign v_30906 = v_30904 & v_30905;
assign v_30909 = v_30907 & v_30908;
assign v_30912 = v_30910 & v_30911;
assign v_30915 = v_30913 & v_30914;
assign v_30918 = v_30916 & v_30917;
assign v_30921 = v_30919 & v_30920;
assign v_30924 = v_30922 & v_30923;
assign v_30927 = v_30925 & v_30926;
assign v_30930 = v_30928 & v_30929;
assign v_30933 = v_30931 & v_30932;
assign v_30936 = v_30934 & v_30935;
assign v_30939 = v_30937 & v_30938;
assign v_30942 = v_30940 & v_30941;
assign v_30945 = v_30943 & v_30944;
assign v_30948 = v_30946 & v_30947;
assign v_30951 = v_30949 & v_30950;
assign v_30954 = v_30952 & v_30953;
assign v_30957 = v_30955 & v_30956;
assign v_30960 = v_30958 & v_30959;
assign v_30963 = v_30961 & v_30962;
assign v_30966 = v_30964 & v_30965;
assign v_30969 = v_30967 & v_30968;
assign v_30972 = v_30970 & v_30971;
assign v_30975 = v_30973 & v_30974;
assign v_30978 = v_30976 & v_30977;
assign v_30981 = v_30979 & v_30980;
assign v_30984 = v_30982 & v_30983;
assign v_30987 = v_30985 & v_30986;
assign v_30990 = v_30988 & v_30989;
assign v_30991 = v_30804 & v_30990;
assign v_30994 = v_30992 & v_30993;
assign v_30997 = v_30995 & v_30996;
assign v_31000 = v_30998 & v_30999;
assign v_31003 = v_31001 & v_31002;
assign v_31006 = v_31004 & v_31005;
assign v_31009 = v_31007 & v_31008;
assign v_31012 = v_31010 & v_31011;
assign v_31015 = v_31013 & v_31014;
assign v_31018 = v_31016 & v_31017;
assign v_31021 = v_31019 & v_31020;
assign v_31024 = v_31022 & v_31023;
assign v_31027 = v_31025 & v_31026;
assign v_31030 = v_31028 & v_31029;
assign v_31033 = v_31031 & v_31032;
assign v_31036 = v_31034 & v_31035;
assign v_31039 = v_31037 & v_31038;
assign v_31042 = v_31040 & v_31041;
assign v_31045 = v_31043 & v_31044;
assign v_31048 = v_31046 & v_31047;
assign v_31051 = v_31049 & v_31050;
assign v_31054 = v_31052 & v_31053;
assign v_31057 = v_31055 & v_31056;
assign v_31060 = v_31058 & v_31059;
assign v_31063 = v_31061 & v_31062;
assign v_31066 = v_31064 & v_31065;
assign v_31069 = v_31067 & v_31068;
assign v_31072 = v_31070 & v_31071;
assign v_31075 = v_31073 & v_31074;
assign v_31078 = v_31076 & v_31077;
assign v_31081 = v_31079 & v_31080;
assign v_31084 = v_31082 & v_31083;
assign v_31087 = v_31085 & v_31086;
assign v_31090 = v_31088 & v_31089;
assign v_31093 = v_31091 & v_31092;
assign v_31096 = v_31094 & v_31095;
assign v_31099 = v_31097 & v_31098;
assign v_31102 = v_31100 & v_31101;
assign v_31105 = v_31103 & v_31104;
assign v_31108 = v_31106 & v_31107;
assign v_31111 = v_31109 & v_31110;
assign v_31114 = v_31112 & v_31113;
assign v_31117 = v_31115 & v_31116;
assign v_31120 = v_31118 & v_31119;
assign v_31123 = v_31121 & v_31122;
assign v_31126 = v_31124 & v_31125;
assign v_31129 = v_31127 & v_31128;
assign v_31132 = v_31130 & v_31131;
assign v_31135 = v_31133 & v_31134;
assign v_31138 = v_31136 & v_31137;
assign v_31141 = v_31139 & v_31140;
assign v_31144 = v_31142 & v_31143;
assign v_31147 = v_31145 & v_31146;
assign v_31150 = v_31148 & v_31149;
assign v_31153 = v_31151 & v_31152;
assign v_31156 = v_31154 & v_31155;
assign v_31159 = v_31157 & v_31158;
assign v_31162 = v_31160 & v_31161;
assign v_31165 = v_31163 & v_31164;
assign v_31168 = v_31166 & v_31167;
assign v_31171 = v_31169 & v_31170;
assign v_31174 = v_31172 & v_31173;
assign v_31177 = v_31175 & v_31176;
assign v_31178 = v_30991 & v_31177;
assign v_31181 = v_31179 & v_31180;
assign v_31184 = v_31182 & v_31183;
assign v_31187 = v_31185 & v_31186;
assign v_31190 = v_31188 & v_31189;
assign v_31193 = v_31191 & v_31192;
assign v_31196 = v_31194 & v_31195;
assign v_31199 = v_31197 & v_31198;
assign v_31202 = v_31200 & v_31201;
assign v_31205 = v_31203 & v_31204;
assign v_31208 = v_31206 & v_31207;
assign v_31211 = v_31209 & v_31210;
assign v_31214 = v_31212 & v_31213;
assign v_31217 = v_31215 & v_31216;
assign v_31220 = v_31218 & v_31219;
assign v_31223 = v_31221 & v_31222;
assign v_31226 = v_31224 & v_31225;
assign v_31229 = v_31227 & v_31228;
assign v_31232 = v_31230 & v_31231;
assign v_31235 = v_31233 & v_31234;
assign v_31238 = v_31236 & v_31237;
assign v_31241 = v_31239 & v_31240;
assign v_31244 = v_31242 & v_31243;
assign v_31247 = v_31245 & v_31246;
assign v_31250 = v_31248 & v_31249;
assign v_31253 = v_31251 & v_31252;
assign v_31256 = v_31254 & v_31255;
assign v_31259 = v_31257 & v_31258;
assign v_31262 = v_31260 & v_31261;
assign v_31265 = v_31263 & v_31264;
assign v_31268 = v_31266 & v_31267;
assign v_31271 = v_31269 & v_31270;
assign v_31274 = v_31272 & v_31273;
assign v_31277 = v_31275 & v_31276;
assign v_31280 = v_31278 & v_31279;
assign v_31283 = v_31281 & v_31282;
assign v_31286 = v_31284 & v_31285;
assign v_31289 = v_31287 & v_31288;
assign v_31292 = v_31290 & v_31291;
assign v_31295 = v_31293 & v_31294;
assign v_31298 = v_31296 & v_31297;
assign v_31301 = v_31299 & v_31300;
assign v_31304 = v_31302 & v_31303;
assign v_31307 = v_31305 & v_31306;
assign v_31310 = v_31308 & v_31309;
assign v_31313 = v_31311 & v_31312;
assign v_31316 = v_31314 & v_31315;
assign v_31319 = v_31317 & v_31318;
assign v_31322 = v_31320 & v_31321;
assign v_31325 = v_31323 & v_31324;
assign v_31328 = v_31326 & v_31327;
assign v_31331 = v_31329 & v_31330;
assign v_31334 = v_31332 & v_31333;
assign v_31337 = v_31335 & v_31336;
assign v_31340 = v_31338 & v_31339;
assign v_31343 = v_31341 & v_31342;
assign v_31346 = v_31344 & v_31345;
assign v_31349 = v_31347 & v_31348;
assign v_31352 = v_31350 & v_31351;
assign v_31355 = v_31353 & v_31354;
assign v_31358 = v_31356 & v_31357;
assign v_31361 = v_31359 & v_31360;
assign v_31364 = v_31362 & v_31363;
assign v_31365 = v_31178 & v_31364;
assign v_31368 = v_31366 & v_31367;
assign v_31371 = v_31369 & v_31370;
assign v_31374 = v_31372 & v_31373;
assign v_31377 = v_31375 & v_31376;
assign v_31380 = v_31378 & v_31379;
assign v_31383 = v_31381 & v_31382;
assign v_31386 = v_31384 & v_31385;
assign v_31389 = v_31387 & v_31388;
assign v_31392 = v_31390 & v_31391;
assign v_31395 = v_31393 & v_31394;
assign v_31398 = v_31396 & v_31397;
assign v_31401 = v_31399 & v_31400;
assign v_31404 = v_31402 & v_31403;
assign v_31407 = v_31405 & v_31406;
assign v_31410 = v_31408 & v_31409;
assign v_31413 = v_31411 & v_31412;
assign v_31416 = v_31414 & v_31415;
assign v_31419 = v_31417 & v_31418;
assign v_31422 = v_31420 & v_31421;
assign v_31425 = v_31423 & v_31424;
assign v_31428 = v_31426 & v_31427;
assign v_31431 = v_31429 & v_31430;
assign v_31434 = v_31432 & v_31433;
assign v_31437 = v_31435 & v_31436;
assign v_31440 = v_31438 & v_31439;
assign v_31443 = v_31441 & v_31442;
assign v_31446 = v_31444 & v_31445;
assign v_31449 = v_31447 & v_31448;
assign v_31452 = v_31450 & v_31451;
assign v_31455 = v_31453 & v_31454;
assign v_31458 = v_31456 & v_31457;
assign v_31461 = v_31459 & v_31460;
assign v_31464 = v_31462 & v_31463;
assign v_31467 = v_31465 & v_31466;
assign v_31470 = v_31468 & v_31469;
assign v_31473 = v_31471 & v_31472;
assign v_31476 = v_31474 & v_31475;
assign v_31479 = v_31477 & v_31478;
assign v_31482 = v_31480 & v_31481;
assign v_31485 = v_31483 & v_31484;
assign v_31488 = v_31486 & v_31487;
assign v_31491 = v_31489 & v_31490;
assign v_31494 = v_31492 & v_31493;
assign v_31497 = v_31495 & v_31496;
assign v_31500 = v_31498 & v_31499;
assign v_31503 = v_31501 & v_31502;
assign v_31506 = v_31504 & v_31505;
assign v_31509 = v_31507 & v_31508;
assign v_31512 = v_31510 & v_31511;
assign v_31515 = v_31513 & v_31514;
assign v_31518 = v_31516 & v_31517;
assign v_31521 = v_31519 & v_31520;
assign v_31524 = v_31522 & v_31523;
assign v_31527 = v_31525 & v_31526;
assign v_31530 = v_31528 & v_31529;
assign v_31533 = v_31531 & v_31532;
assign v_31536 = v_31534 & v_31535;
assign v_31539 = v_31537 & v_31538;
assign v_31542 = v_31540 & v_31541;
assign v_31545 = v_31543 & v_31544;
assign v_31548 = v_31546 & v_31547;
assign v_31551 = v_31549 & v_31550;
assign v_31552 = v_31365 & v_31551;
assign v_31555 = v_31553 & v_31554;
assign v_31558 = v_31556 & v_31557;
assign v_31561 = v_31559 & v_31560;
assign v_31564 = v_31562 & v_31563;
assign v_31567 = v_31565 & v_31566;
assign v_31570 = v_31568 & v_31569;
assign v_31573 = v_31571 & v_31572;
assign v_31576 = v_31574 & v_31575;
assign v_31579 = v_31577 & v_31578;
assign v_31582 = v_31580 & v_31581;
assign v_31585 = v_31583 & v_31584;
assign v_31588 = v_31586 & v_31587;
assign v_31591 = v_31589 & v_31590;
assign v_31594 = v_31592 & v_31593;
assign v_31597 = v_31595 & v_31596;
assign v_31600 = v_31598 & v_31599;
assign v_31603 = v_31601 & v_31602;
assign v_31606 = v_31604 & v_31605;
assign v_31609 = v_31607 & v_31608;
assign v_31612 = v_31610 & v_31611;
assign v_31615 = v_31613 & v_31614;
assign v_31618 = v_31616 & v_31617;
assign v_31621 = v_31619 & v_31620;
assign v_31624 = v_31622 & v_31623;
assign v_31627 = v_31625 & v_31626;
assign v_31630 = v_31628 & v_31629;
assign v_31633 = v_31631 & v_31632;
assign v_31636 = v_31634 & v_31635;
assign v_31639 = v_31637 & v_31638;
assign v_31642 = v_31640 & v_31641;
assign v_31645 = v_31643 & v_31644;
assign v_31648 = v_31646 & v_31647;
assign v_31651 = v_31649 & v_31650;
assign v_31654 = v_31652 & v_31653;
assign v_31657 = v_31655 & v_31656;
assign v_31660 = v_31658 & v_31659;
assign v_31663 = v_31661 & v_31662;
assign v_31666 = v_31664 & v_31665;
assign v_31669 = v_31667 & v_31668;
assign v_31672 = v_31670 & v_31671;
assign v_31675 = v_31673 & v_31674;
assign v_31678 = v_31676 & v_31677;
assign v_31681 = v_31679 & v_31680;
assign v_31684 = v_31682 & v_31683;
assign v_31687 = v_31685 & v_31686;
assign v_31690 = v_31688 & v_31689;
assign v_31693 = v_31691 & v_31692;
assign v_31696 = v_31694 & v_31695;
assign v_31699 = v_31697 & v_31698;
assign v_31702 = v_31700 & v_31701;
assign v_31705 = v_31703 & v_31704;
assign v_31708 = v_31706 & v_31707;
assign v_31711 = v_31709 & v_31710;
assign v_31714 = v_31712 & v_31713;
assign v_31717 = v_31715 & v_31716;
assign v_31720 = v_31718 & v_31719;
assign v_31723 = v_31721 & v_31722;
assign v_31726 = v_31724 & v_31725;
assign v_31729 = v_31727 & v_31728;
assign v_31732 = v_31730 & v_31731;
assign v_31735 = v_31733 & v_31734;
assign v_31738 = v_31736 & v_31737;
assign v_31739 = v_31552 & v_31738;
assign v_31740 = v_23172 & v_31739;
assign v_31743 = v_31741 & v_31742;
assign v_31746 = v_31744 & v_31745;
assign v_31749 = v_31747 & v_31748;
assign v_31752 = v_31750 & v_31751;
assign v_31755 = v_31753 & v_31754;
assign v_31758 = v_31756 & v_31757;
assign v_31761 = v_31759 & v_31760;
assign v_31764 = v_31762 & v_31763;
assign v_31767 = v_31765 & v_31766;
assign v_31770 = v_31768 & v_31769;
assign v_31773 = v_31771 & v_31772;
assign v_31776 = v_31774 & v_31775;
assign v_31779 = v_31777 & v_31778;
assign v_31782 = v_31780 & v_31781;
assign v_31785 = v_31783 & v_31784;
assign v_31788 = v_31786 & v_31787;
assign v_31791 = v_31789 & v_31790;
assign v_31794 = v_31792 & v_31793;
assign v_31797 = v_31795 & v_31796;
assign v_31800 = v_31798 & v_31799;
assign v_31803 = v_31801 & v_31802;
assign v_31806 = v_31804 & v_31805;
assign v_31809 = v_31807 & v_31808;
assign v_31812 = v_31810 & v_31811;
assign v_31815 = v_31813 & v_31814;
assign v_31818 = v_31816 & v_31817;
assign v_31821 = v_31819 & v_31820;
assign v_31824 = v_31822 & v_31823;
assign v_31827 = v_31825 & v_31826;
assign v_31830 = v_31828 & v_31829;
assign v_31833 = v_31831 & v_31832;
assign v_31836 = v_31834 & v_31835;
assign v_31839 = v_31837 & v_31838;
assign v_31842 = v_31840 & v_31841;
assign v_31845 = v_31843 & v_31844;
assign v_31848 = v_31846 & v_31847;
assign v_31851 = v_31849 & v_31850;
assign v_31854 = v_31852 & v_31853;
assign v_31857 = v_31855 & v_31856;
assign v_31860 = v_31858 & v_31859;
assign v_31863 = v_31861 & v_31862;
assign v_31866 = v_31864 & v_31865;
assign v_31869 = v_31867 & v_31868;
assign v_31872 = v_31870 & v_31871;
assign v_31875 = v_31873 & v_31874;
assign v_31878 = v_31876 & v_31877;
assign v_31881 = v_31879 & v_31880;
assign v_31884 = v_31882 & v_31883;
assign v_31887 = v_31885 & v_31886;
assign v_31890 = v_31888 & v_31889;
assign v_31893 = v_31891 & v_31892;
assign v_31896 = v_31894 & v_31895;
assign v_31899 = v_31897 & v_31898;
assign v_31902 = v_31900 & v_31901;
assign v_31905 = v_31903 & v_31904;
assign v_31908 = v_31906 & v_31907;
assign v_31911 = v_31909 & v_31910;
assign v_31914 = v_31912 & v_31913;
assign v_31917 = v_31915 & v_31916;
assign v_31920 = v_31918 & v_31919;
assign v_31923 = v_31921 & v_31922;
assign v_31926 = v_31924 & v_31925;
assign v_31927 = v_31740 & v_31926;
assign v_31928 = v_26290 & v_31927;
assign v_31929 = v_30618 & v_31928;
assign v_31930 = ~v_10462 & v_31929;
assign v_31934 = v_31932 & v_31933;
assign v_31937 = v_31935 & v_31936;
assign v_31940 = v_31938 & v_31939;
assign v_31943 = v_31941 & v_31942;
assign v_31946 = v_31944 & v_31945;
assign v_31949 = v_31947 & v_31948;
assign v_31952 = v_31950 & v_31951;
assign v_31955 = v_31953 & v_31954;
assign v_31958 = v_31956 & v_31957;
assign v_31961 = v_31959 & v_31960;
assign v_31964 = v_31962 & v_31963;
assign v_31967 = v_31965 & v_31966;
assign v_31970 = v_31968 & v_31969;
assign v_31973 = v_31971 & v_31972;
assign v_31976 = v_31974 & v_31975;
assign v_31979 = v_31977 & v_31978;
assign v_31982 = v_31980 & v_31981;
assign v_31985 = v_31983 & v_31984;
assign v_31988 = v_31986 & v_31987;
assign v_31991 = v_31989 & v_31990;
assign v_31994 = v_31992 & v_31993;
assign v_31997 = v_31995 & v_31996;
assign v_32000 = v_31998 & v_31999;
assign v_32003 = v_32001 & v_32002;
assign v_32006 = v_32004 & v_32005;
assign v_32009 = v_32007 & v_32008;
assign v_32012 = v_32010 & v_32011;
assign v_32015 = v_32013 & v_32014;
assign v_32018 = v_32016 & v_32017;
assign v_32021 = v_32019 & v_32020;
assign v_32024 = v_32022 & v_32023;
assign v_32027 = v_32025 & v_32026;
assign v_32030 = v_32028 & v_32029;
assign v_32033 = v_32031 & v_32032;
assign v_32036 = v_32034 & v_32035;
assign v_32039 = v_32037 & v_32038;
assign v_32042 = v_32040 & v_32041;
assign v_32045 = v_32043 & v_32044;
assign v_32048 = v_32046 & v_32047;
assign v_32051 = v_32049 & v_32050;
assign v_32054 = v_32052 & v_32053;
assign v_32057 = v_32055 & v_32056;
assign v_32060 = v_32058 & v_32059;
assign v_32063 = v_32061 & v_32062;
assign v_32066 = v_32064 & v_32065;
assign v_32069 = v_32067 & v_32068;
assign v_32072 = v_32070 & v_32071;
assign v_32075 = v_32073 & v_32074;
assign v_32078 = v_32076 & v_32077;
assign v_32081 = v_32079 & v_32080;
assign v_32084 = v_32082 & v_32083;
assign v_32087 = v_32085 & v_32086;
assign v_32090 = v_32088 & v_32089;
assign v_32093 = v_32091 & v_32092;
assign v_32096 = v_32094 & v_32095;
assign v_32099 = v_32097 & v_32098;
assign v_32102 = v_32100 & v_32101;
assign v_32105 = v_32103 & v_32104;
assign v_32108 = v_32106 & v_32107;
assign v_32111 = v_32109 & v_32110;
assign v_32114 = v_32112 & v_32113;
assign v_32117 = v_32115 & v_32116;
assign v_32120 = v_32118 & v_32119;
assign v_32123 = v_32121 & v_32122;
assign v_32126 = v_32124 & v_32125;
assign v_32129 = v_32127 & v_32128;
assign v_32132 = v_32130 & v_32131;
assign v_32135 = v_32133 & v_32134;
assign v_32138 = v_32136 & v_32137;
assign v_32141 = v_32139 & v_32140;
assign v_32144 = v_32142 & v_32143;
assign v_32147 = v_32145 & v_32146;
assign v_32150 = v_32148 & v_32149;
assign v_32153 = v_32151 & v_32152;
assign v_32156 = v_32154 & v_32155;
assign v_32159 = v_32157 & v_32158;
assign v_32162 = v_32160 & v_32161;
assign v_32165 = v_32163 & v_32164;
assign v_32168 = v_32166 & v_32167;
assign v_32171 = v_32169 & v_32170;
assign v_32174 = v_32172 & v_32173;
assign v_32177 = v_32175 & v_32176;
assign v_32180 = v_32178 & v_32179;
assign v_32183 = v_32181 & v_32182;
assign v_32186 = v_32184 & v_32185;
assign v_32189 = v_32187 & v_32188;
assign v_32192 = v_32190 & v_32191;
assign v_32195 = v_32193 & v_32194;
assign v_32198 = v_32196 & v_32197;
assign v_32201 = v_32199 & v_32200;
assign v_32204 = v_32202 & v_32203;
assign v_32207 = v_32205 & v_32206;
assign v_32210 = v_32208 & v_32209;
assign v_32213 = v_32211 & v_32212;
assign v_32216 = v_32214 & v_32215;
assign v_32219 = v_32217 & v_32218;
assign v_32222 = v_32220 & v_32221;
assign v_32225 = v_32223 & v_32224;
assign v_32228 = v_32226 & v_32227;
assign v_32231 = v_32229 & v_32230;
assign v_32234 = v_32232 & v_32233;
assign v_32237 = v_32235 & v_32236;
assign v_32240 = v_32238 & v_32239;
assign v_32243 = v_32241 & v_32242;
assign v_32246 = v_32244 & v_32245;
assign v_32249 = v_32247 & v_32248;
assign v_32252 = v_32250 & v_32251;
assign v_32255 = v_32253 & v_32254;
assign v_32258 = v_32256 & v_32257;
assign v_32261 = v_32259 & v_32260;
assign v_32264 = v_32262 & v_32263;
assign v_32267 = v_32265 & v_32266;
assign v_32270 = v_32268 & v_32269;
assign v_32273 = v_32271 & v_32272;
assign v_32276 = v_32274 & v_32275;
assign v_32279 = v_32277 & v_32278;
assign v_32282 = v_32280 & v_32281;
assign v_32285 = v_32283 & v_32284;
assign v_32288 = v_32286 & v_32287;
assign v_32291 = v_32289 & v_32290;
assign v_32294 = v_32292 & v_32293;
assign v_32297 = v_32295 & v_32296;
assign v_32300 = v_32298 & v_32299;
assign v_32303 = v_32301 & v_32302;
assign v_32306 = v_32304 & v_32305;
assign v_32309 = v_32307 & v_32308;
assign v_32310 = v_32120 & v_32309;
assign v_32313 = v_32311 & v_32312;
assign v_32316 = v_32314 & v_32315;
assign v_32319 = v_32317 & v_32318;
assign v_32322 = v_32320 & v_32321;
assign v_32325 = v_32323 & v_32324;
assign v_32328 = v_32326 & v_32327;
assign v_32331 = v_32329 & v_32330;
assign v_32334 = v_32332 & v_32333;
assign v_32337 = v_32335 & v_32336;
assign v_32340 = v_32338 & v_32339;
assign v_32343 = v_32341 & v_32342;
assign v_32346 = v_32344 & v_32345;
assign v_32349 = v_32347 & v_32348;
assign v_32352 = v_32350 & v_32351;
assign v_32355 = v_32353 & v_32354;
assign v_32358 = v_32356 & v_32357;
assign v_32361 = v_32359 & v_32360;
assign v_32364 = v_32362 & v_32363;
assign v_32367 = v_32365 & v_32366;
assign v_32370 = v_32368 & v_32369;
assign v_32373 = v_32371 & v_32372;
assign v_32376 = v_32374 & v_32375;
assign v_32379 = v_32377 & v_32378;
assign v_32382 = v_32380 & v_32381;
assign v_32385 = v_32383 & v_32384;
assign v_32388 = v_32386 & v_32387;
assign v_32391 = v_32389 & v_32390;
assign v_32394 = v_32392 & v_32393;
assign v_32397 = v_32395 & v_32396;
assign v_32400 = v_32398 & v_32399;
assign v_32403 = v_32401 & v_32402;
assign v_32406 = v_32404 & v_32405;
assign v_32409 = v_32407 & v_32408;
assign v_32412 = v_32410 & v_32411;
assign v_32415 = v_32413 & v_32414;
assign v_32418 = v_32416 & v_32417;
assign v_32421 = v_32419 & v_32420;
assign v_32424 = v_32422 & v_32423;
assign v_32427 = v_32425 & v_32426;
assign v_32430 = v_32428 & v_32429;
assign v_32433 = v_32431 & v_32432;
assign v_32436 = v_32434 & v_32435;
assign v_32439 = v_32437 & v_32438;
assign v_32442 = v_32440 & v_32441;
assign v_32445 = v_32443 & v_32444;
assign v_32448 = v_32446 & v_32447;
assign v_32451 = v_32449 & v_32450;
assign v_32454 = v_32452 & v_32453;
assign v_32457 = v_32455 & v_32456;
assign v_32460 = v_32458 & v_32459;
assign v_32463 = v_32461 & v_32462;
assign v_32466 = v_32464 & v_32465;
assign v_32469 = v_32467 & v_32468;
assign v_32472 = v_32470 & v_32471;
assign v_32475 = v_32473 & v_32474;
assign v_32478 = v_32476 & v_32477;
assign v_32481 = v_32479 & v_32480;
assign v_32484 = v_32482 & v_32483;
assign v_32487 = v_32485 & v_32486;
assign v_32490 = v_32488 & v_32489;
assign v_32493 = v_32491 & v_32492;
assign v_32496 = v_32494 & v_32495;
assign v_32499 = v_32497 & v_32498;
assign v_32500 = v_32310 & v_32499;
assign v_32503 = v_32501 & v_32502;
assign v_32506 = v_32504 & v_32505;
assign v_32509 = v_32507 & v_32508;
assign v_32512 = v_32510 & v_32511;
assign v_32515 = v_32513 & v_32514;
assign v_32518 = v_32516 & v_32517;
assign v_32521 = v_32519 & v_32520;
assign v_32524 = v_32522 & v_32523;
assign v_32527 = v_32525 & v_32526;
assign v_32530 = v_32528 & v_32529;
assign v_32533 = v_32531 & v_32532;
assign v_32536 = v_32534 & v_32535;
assign v_32539 = v_32537 & v_32538;
assign v_32542 = v_32540 & v_32541;
assign v_32545 = v_32543 & v_32544;
assign v_32548 = v_32546 & v_32547;
assign v_32551 = v_32549 & v_32550;
assign v_32554 = v_32552 & v_32553;
assign v_32557 = v_32555 & v_32556;
assign v_32560 = v_32558 & v_32559;
assign v_32563 = v_32561 & v_32562;
assign v_32566 = v_32564 & v_32565;
assign v_32569 = v_32567 & v_32568;
assign v_32572 = v_32570 & v_32571;
assign v_32575 = v_32573 & v_32574;
assign v_32578 = v_32576 & v_32577;
assign v_32581 = v_32579 & v_32580;
assign v_32584 = v_32582 & v_32583;
assign v_32587 = v_32585 & v_32586;
assign v_32590 = v_32588 & v_32589;
assign v_32593 = v_32591 & v_32592;
assign v_32596 = v_32594 & v_32595;
assign v_32599 = v_32597 & v_32598;
assign v_32602 = v_32600 & v_32601;
assign v_32605 = v_32603 & v_32604;
assign v_32608 = v_32606 & v_32607;
assign v_32611 = v_32609 & v_32610;
assign v_32614 = v_32612 & v_32613;
assign v_32617 = v_32615 & v_32616;
assign v_32620 = v_32618 & v_32619;
assign v_32623 = v_32621 & v_32622;
assign v_32626 = v_32624 & v_32625;
assign v_32629 = v_32627 & v_32628;
assign v_32632 = v_32630 & v_32631;
assign v_32635 = v_32633 & v_32634;
assign v_32638 = v_32636 & v_32637;
assign v_32641 = v_32639 & v_32640;
assign v_32644 = v_32642 & v_32643;
assign v_32647 = v_32645 & v_32646;
assign v_32650 = v_32648 & v_32649;
assign v_32653 = v_32651 & v_32652;
assign v_32656 = v_32654 & v_32655;
assign v_32659 = v_32657 & v_32658;
assign v_32662 = v_32660 & v_32661;
assign v_32665 = v_32663 & v_32664;
assign v_32668 = v_32666 & v_32667;
assign v_32671 = v_32669 & v_32670;
assign v_32674 = v_32672 & v_32673;
assign v_32677 = v_32675 & v_32676;
assign v_32680 = v_32678 & v_32679;
assign v_32683 = v_32681 & v_32682;
assign v_32686 = v_32684 & v_32685;
assign v_32689 = v_32687 & v_32688;
assign v_32690 = v_32500 & v_32689;
assign v_32693 = v_32691 & v_32692;
assign v_32696 = v_32694 & v_32695;
assign v_32699 = v_32697 & v_32698;
assign v_32702 = v_32700 & v_32701;
assign v_32705 = v_32703 & v_32704;
assign v_32708 = v_32706 & v_32707;
assign v_32711 = v_32709 & v_32710;
assign v_32714 = v_32712 & v_32713;
assign v_32717 = v_32715 & v_32716;
assign v_32720 = v_32718 & v_32719;
assign v_32723 = v_32721 & v_32722;
assign v_32726 = v_32724 & v_32725;
assign v_32729 = v_32727 & v_32728;
assign v_32732 = v_32730 & v_32731;
assign v_32735 = v_32733 & v_32734;
assign v_32738 = v_32736 & v_32737;
assign v_32741 = v_32739 & v_32740;
assign v_32744 = v_32742 & v_32743;
assign v_32747 = v_32745 & v_32746;
assign v_32750 = v_32748 & v_32749;
assign v_32753 = v_32751 & v_32752;
assign v_32756 = v_32754 & v_32755;
assign v_32759 = v_32757 & v_32758;
assign v_32762 = v_32760 & v_32761;
assign v_32765 = v_32763 & v_32764;
assign v_32768 = v_32766 & v_32767;
assign v_32771 = v_32769 & v_32770;
assign v_32774 = v_32772 & v_32773;
assign v_32777 = v_32775 & v_32776;
assign v_32780 = v_32778 & v_32779;
assign v_32783 = v_32781 & v_32782;
assign v_32786 = v_32784 & v_32785;
assign v_32789 = v_32787 & v_32788;
assign v_32792 = v_32790 & v_32791;
assign v_32795 = v_32793 & v_32794;
assign v_32798 = v_32796 & v_32797;
assign v_32801 = v_32799 & v_32800;
assign v_32804 = v_32802 & v_32803;
assign v_32807 = v_32805 & v_32806;
assign v_32810 = v_32808 & v_32809;
assign v_32813 = v_32811 & v_32812;
assign v_32816 = v_32814 & v_32815;
assign v_32819 = v_32817 & v_32818;
assign v_32822 = v_32820 & v_32821;
assign v_32825 = v_32823 & v_32824;
assign v_32828 = v_32826 & v_32827;
assign v_32831 = v_32829 & v_32830;
assign v_32834 = v_32832 & v_32833;
assign v_32837 = v_32835 & v_32836;
assign v_32840 = v_32838 & v_32839;
assign v_32843 = v_32841 & v_32842;
assign v_32846 = v_32844 & v_32845;
assign v_32849 = v_32847 & v_32848;
assign v_32852 = v_32850 & v_32851;
assign v_32855 = v_32853 & v_32854;
assign v_32858 = v_32856 & v_32857;
assign v_32861 = v_32859 & v_32860;
assign v_32864 = v_32862 & v_32863;
assign v_32867 = v_32865 & v_32866;
assign v_32870 = v_32868 & v_32869;
assign v_32873 = v_32871 & v_32872;
assign v_32876 = v_32874 & v_32875;
assign v_32879 = v_32877 & v_32878;
assign v_32880 = v_32690 & v_32879;
assign v_32883 = v_32881 & v_32882;
assign v_32886 = v_32884 & v_32885;
assign v_32889 = v_32887 & v_32888;
assign v_32892 = v_32890 & v_32891;
assign v_32895 = v_32893 & v_32894;
assign v_32898 = v_32896 & v_32897;
assign v_32901 = v_32899 & v_32900;
assign v_32904 = v_32902 & v_32903;
assign v_32907 = v_32905 & v_32906;
assign v_32910 = v_32908 & v_32909;
assign v_32913 = v_32911 & v_32912;
assign v_32916 = v_32914 & v_32915;
assign v_32919 = v_32917 & v_32918;
assign v_32922 = v_32920 & v_32921;
assign v_32925 = v_32923 & v_32924;
assign v_32928 = v_32926 & v_32927;
assign v_32931 = v_32929 & v_32930;
assign v_32934 = v_32932 & v_32933;
assign v_32937 = v_32935 & v_32936;
assign v_32940 = v_32938 & v_32939;
assign v_32943 = v_32941 & v_32942;
assign v_32946 = v_32944 & v_32945;
assign v_32949 = v_32947 & v_32948;
assign v_32952 = v_32950 & v_32951;
assign v_32955 = v_32953 & v_32954;
assign v_32958 = v_32956 & v_32957;
assign v_32961 = v_32959 & v_32960;
assign v_32964 = v_32962 & v_32963;
assign v_32967 = v_32965 & v_32966;
assign v_32970 = v_32968 & v_32969;
assign v_32973 = v_32971 & v_32972;
assign v_32976 = v_32974 & v_32975;
assign v_32979 = v_32977 & v_32978;
assign v_32982 = v_32980 & v_32981;
assign v_32985 = v_32983 & v_32984;
assign v_32988 = v_32986 & v_32987;
assign v_32991 = v_32989 & v_32990;
assign v_32994 = v_32992 & v_32993;
assign v_32997 = v_32995 & v_32996;
assign v_33000 = v_32998 & v_32999;
assign v_33003 = v_33001 & v_33002;
assign v_33006 = v_33004 & v_33005;
assign v_33009 = v_33007 & v_33008;
assign v_33012 = v_33010 & v_33011;
assign v_33015 = v_33013 & v_33014;
assign v_33018 = v_33016 & v_33017;
assign v_33021 = v_33019 & v_33020;
assign v_33024 = v_33022 & v_33023;
assign v_33027 = v_33025 & v_33026;
assign v_33030 = v_33028 & v_33029;
assign v_33033 = v_33031 & v_33032;
assign v_33036 = v_33034 & v_33035;
assign v_33039 = v_33037 & v_33038;
assign v_33042 = v_33040 & v_33041;
assign v_33045 = v_33043 & v_33044;
assign v_33048 = v_33046 & v_33047;
assign v_33051 = v_33049 & v_33050;
assign v_33054 = v_33052 & v_33053;
assign v_33057 = v_33055 & v_33056;
assign v_33060 = v_33058 & v_33059;
assign v_33063 = v_33061 & v_33062;
assign v_33066 = v_33064 & v_33065;
assign v_33069 = v_33067 & v_33068;
assign v_33070 = v_32880 & v_33069;
assign v_33073 = v_33071 & v_33072;
assign v_33076 = v_33074 & v_33075;
assign v_33079 = v_33077 & v_33078;
assign v_33082 = v_33080 & v_33081;
assign v_33085 = v_33083 & v_33084;
assign v_33088 = v_33086 & v_33087;
assign v_33091 = v_33089 & v_33090;
assign v_33094 = v_33092 & v_33093;
assign v_33097 = v_33095 & v_33096;
assign v_33100 = v_33098 & v_33099;
assign v_33103 = v_33101 & v_33102;
assign v_33106 = v_33104 & v_33105;
assign v_33109 = v_33107 & v_33108;
assign v_33112 = v_33110 & v_33111;
assign v_33115 = v_33113 & v_33114;
assign v_33118 = v_33116 & v_33117;
assign v_33121 = v_33119 & v_33120;
assign v_33124 = v_33122 & v_33123;
assign v_33127 = v_33125 & v_33126;
assign v_33130 = v_33128 & v_33129;
assign v_33133 = v_33131 & v_33132;
assign v_33136 = v_33134 & v_33135;
assign v_33139 = v_33137 & v_33138;
assign v_33142 = v_33140 & v_33141;
assign v_33145 = v_33143 & v_33144;
assign v_33148 = v_33146 & v_33147;
assign v_33151 = v_33149 & v_33150;
assign v_33154 = v_33152 & v_33153;
assign v_33157 = v_33155 & v_33156;
assign v_33160 = v_33158 & v_33159;
assign v_33163 = v_33161 & v_33162;
assign v_33166 = v_33164 & v_33165;
assign v_33169 = v_33167 & v_33168;
assign v_33172 = v_33170 & v_33171;
assign v_33175 = v_33173 & v_33174;
assign v_33178 = v_33176 & v_33177;
assign v_33181 = v_33179 & v_33180;
assign v_33184 = v_33182 & v_33183;
assign v_33187 = v_33185 & v_33186;
assign v_33190 = v_33188 & v_33189;
assign v_33193 = v_33191 & v_33192;
assign v_33196 = v_33194 & v_33195;
assign v_33199 = v_33197 & v_33198;
assign v_33202 = v_33200 & v_33201;
assign v_33205 = v_33203 & v_33204;
assign v_33208 = v_33206 & v_33207;
assign v_33211 = v_33209 & v_33210;
assign v_33214 = v_33212 & v_33213;
assign v_33217 = v_33215 & v_33216;
assign v_33220 = v_33218 & v_33219;
assign v_33223 = v_33221 & v_33222;
assign v_33226 = v_33224 & v_33225;
assign v_33229 = v_33227 & v_33228;
assign v_33232 = v_33230 & v_33231;
assign v_33235 = v_33233 & v_33234;
assign v_33238 = v_33236 & v_33237;
assign v_33241 = v_33239 & v_33240;
assign v_33244 = v_33242 & v_33243;
assign v_33247 = v_33245 & v_33246;
assign v_33250 = v_33248 & v_33249;
assign v_33253 = v_33251 & v_33252;
assign v_33256 = v_33254 & v_33255;
assign v_33259 = v_33257 & v_33258;
assign v_33260 = v_33070 & v_33259;
assign v_33263 = v_33261 & v_33262;
assign v_33266 = v_33264 & v_33265;
assign v_33269 = v_33267 & v_33268;
assign v_33272 = v_33270 & v_33271;
assign v_33275 = v_33273 & v_33274;
assign v_33278 = v_33276 & v_33277;
assign v_33281 = v_33279 & v_33280;
assign v_33284 = v_33282 & v_33283;
assign v_33287 = v_33285 & v_33286;
assign v_33290 = v_33288 & v_33289;
assign v_33293 = v_33291 & v_33292;
assign v_33296 = v_33294 & v_33295;
assign v_33299 = v_33297 & v_33298;
assign v_33302 = v_33300 & v_33301;
assign v_33305 = v_33303 & v_33304;
assign v_33308 = v_33306 & v_33307;
assign v_33311 = v_33309 & v_33310;
assign v_33314 = v_33312 & v_33313;
assign v_33317 = v_33315 & v_33316;
assign v_33320 = v_33318 & v_33319;
assign v_33323 = v_33321 & v_33322;
assign v_33326 = v_33324 & v_33325;
assign v_33329 = v_33327 & v_33328;
assign v_33332 = v_33330 & v_33331;
assign v_33335 = v_33333 & v_33334;
assign v_33338 = v_33336 & v_33337;
assign v_33341 = v_33339 & v_33340;
assign v_33344 = v_33342 & v_33343;
assign v_33347 = v_33345 & v_33346;
assign v_33350 = v_33348 & v_33349;
assign v_33353 = v_33351 & v_33352;
assign v_33356 = v_33354 & v_33355;
assign v_33359 = v_33357 & v_33358;
assign v_33362 = v_33360 & v_33361;
assign v_33365 = v_33363 & v_33364;
assign v_33368 = v_33366 & v_33367;
assign v_33371 = v_33369 & v_33370;
assign v_33374 = v_33372 & v_33373;
assign v_33377 = v_33375 & v_33376;
assign v_33380 = v_33378 & v_33379;
assign v_33383 = v_33381 & v_33382;
assign v_33386 = v_33384 & v_33385;
assign v_33389 = v_33387 & v_33388;
assign v_33392 = v_33390 & v_33391;
assign v_33395 = v_33393 & v_33394;
assign v_33398 = v_33396 & v_33397;
assign v_33401 = v_33399 & v_33400;
assign v_33404 = v_33402 & v_33403;
assign v_33407 = v_33405 & v_33406;
assign v_33410 = v_33408 & v_33409;
assign v_33413 = v_33411 & v_33412;
assign v_33416 = v_33414 & v_33415;
assign v_33419 = v_33417 & v_33418;
assign v_33422 = v_33420 & v_33421;
assign v_33425 = v_33423 & v_33424;
assign v_33428 = v_33426 & v_33427;
assign v_33431 = v_33429 & v_33430;
assign v_33434 = v_33432 & v_33433;
assign v_33437 = v_33435 & v_33436;
assign v_33440 = v_33438 & v_33439;
assign v_33443 = v_33441 & v_33442;
assign v_33446 = v_33444 & v_33445;
assign v_33449 = v_33447 & v_33448;
assign v_33450 = v_33260 & v_33449;
assign v_33453 = v_33451 & v_33452;
assign v_33456 = v_33454 & v_33455;
assign v_33459 = v_33457 & v_33458;
assign v_33462 = v_33460 & v_33461;
assign v_33465 = v_33463 & v_33464;
assign v_33468 = v_33466 & v_33467;
assign v_33471 = v_33469 & v_33470;
assign v_33474 = v_33472 & v_33473;
assign v_33477 = v_33475 & v_33476;
assign v_33480 = v_33478 & v_33479;
assign v_33483 = v_33481 & v_33482;
assign v_33486 = v_33484 & v_33485;
assign v_33489 = v_33487 & v_33488;
assign v_33492 = v_33490 & v_33491;
assign v_33495 = v_33493 & v_33494;
assign v_33498 = v_33496 & v_33497;
assign v_33501 = v_33499 & v_33500;
assign v_33504 = v_33502 & v_33503;
assign v_33507 = v_33505 & v_33506;
assign v_33510 = v_33508 & v_33509;
assign v_33513 = v_33511 & v_33512;
assign v_33516 = v_33514 & v_33515;
assign v_33519 = v_33517 & v_33518;
assign v_33522 = v_33520 & v_33521;
assign v_33525 = v_33523 & v_33524;
assign v_33528 = v_33526 & v_33527;
assign v_33531 = v_33529 & v_33530;
assign v_33534 = v_33532 & v_33533;
assign v_33537 = v_33535 & v_33536;
assign v_33540 = v_33538 & v_33539;
assign v_33543 = v_33541 & v_33542;
assign v_33546 = v_33544 & v_33545;
assign v_33549 = v_33547 & v_33548;
assign v_33552 = v_33550 & v_33551;
assign v_33555 = v_33553 & v_33554;
assign v_33558 = v_33556 & v_33557;
assign v_33561 = v_33559 & v_33560;
assign v_33564 = v_33562 & v_33563;
assign v_33567 = v_33565 & v_33566;
assign v_33570 = v_33568 & v_33569;
assign v_33573 = v_33571 & v_33572;
assign v_33576 = v_33574 & v_33575;
assign v_33579 = v_33577 & v_33578;
assign v_33582 = v_33580 & v_33581;
assign v_33585 = v_33583 & v_33584;
assign v_33588 = v_33586 & v_33587;
assign v_33591 = v_33589 & v_33590;
assign v_33594 = v_33592 & v_33593;
assign v_33597 = v_33595 & v_33596;
assign v_33600 = v_33598 & v_33599;
assign v_33603 = v_33601 & v_33602;
assign v_33606 = v_33604 & v_33605;
assign v_33609 = v_33607 & v_33608;
assign v_33612 = v_33610 & v_33611;
assign v_33615 = v_33613 & v_33614;
assign v_33618 = v_33616 & v_33617;
assign v_33621 = v_33619 & v_33620;
assign v_33624 = v_33622 & v_33623;
assign v_33627 = v_33625 & v_33626;
assign v_33630 = v_33628 & v_33629;
assign v_33633 = v_33631 & v_33632;
assign v_33636 = v_33634 & v_33635;
assign v_33639 = v_33637 & v_33638;
assign v_33642 = v_33640 & v_33641;
assign v_33645 = v_33643 & v_33644;
assign v_33648 = v_33646 & v_33647;
assign v_33651 = v_33649 & v_33650;
assign v_33654 = v_33652 & v_33653;
assign v_33657 = v_33655 & v_33656;
assign v_33660 = v_33658 & v_33659;
assign v_33663 = v_33661 & v_33662;
assign v_33666 = v_33664 & v_33665;
assign v_33669 = v_33667 & v_33668;
assign v_33672 = v_33670 & v_33671;
assign v_33675 = v_33673 & v_33674;
assign v_33678 = v_33676 & v_33677;
assign v_33681 = v_33679 & v_33680;
assign v_33684 = v_33682 & v_33683;
assign v_33687 = v_33685 & v_33686;
assign v_33690 = v_33688 & v_33689;
assign v_33693 = v_33691 & v_33692;
assign v_33696 = v_33694 & v_33695;
assign v_33699 = v_33697 & v_33698;
assign v_33702 = v_33700 & v_33701;
assign v_33705 = v_33703 & v_33704;
assign v_33708 = v_33706 & v_33707;
assign v_33711 = v_33709 & v_33710;
assign v_33714 = v_33712 & v_33713;
assign v_33717 = v_33715 & v_33716;
assign v_33720 = v_33718 & v_33719;
assign v_33723 = v_33721 & v_33722;
assign v_33726 = v_33724 & v_33725;
assign v_33729 = v_33727 & v_33728;
assign v_33732 = v_33730 & v_33731;
assign v_33735 = v_33733 & v_33734;
assign v_33738 = v_33736 & v_33737;
assign v_33741 = v_33739 & v_33740;
assign v_33744 = v_33742 & v_33743;
assign v_33747 = v_33745 & v_33746;
assign v_33750 = v_33748 & v_33749;
assign v_33753 = v_33751 & v_33752;
assign v_33756 = v_33754 & v_33755;
assign v_33759 = v_33757 & v_33758;
assign v_33762 = v_33760 & v_33761;
assign v_33765 = v_33763 & v_33764;
assign v_33768 = v_33766 & v_33767;
assign v_33771 = v_33769 & v_33770;
assign v_33774 = v_33772 & v_33773;
assign v_33777 = v_33775 & v_33776;
assign v_33780 = v_33778 & v_33779;
assign v_33783 = v_33781 & v_33782;
assign v_33786 = v_33784 & v_33785;
assign v_33789 = v_33787 & v_33788;
assign v_33792 = v_33790 & v_33791;
assign v_33795 = v_33793 & v_33794;
assign v_33798 = v_33796 & v_33797;
assign v_33801 = v_33799 & v_33800;
assign v_33804 = v_33802 & v_33803;
assign v_33807 = v_33805 & v_33806;
assign v_33810 = v_33808 & v_33809;
assign v_33813 = v_33811 & v_33812;
assign v_33816 = v_33814 & v_33815;
assign v_33819 = v_33817 & v_33818;
assign v_33822 = v_33820 & v_33821;
assign v_33825 = v_33823 & v_33824;
assign v_33828 = v_33826 & v_33827;
assign v_33829 = v_33639 & v_33828;
assign v_33832 = v_33830 & v_33831;
assign v_33835 = v_33833 & v_33834;
assign v_33838 = v_33836 & v_33837;
assign v_33841 = v_33839 & v_33840;
assign v_33844 = v_33842 & v_33843;
assign v_33847 = v_33845 & v_33846;
assign v_33850 = v_33848 & v_33849;
assign v_33853 = v_33851 & v_33852;
assign v_33856 = v_33854 & v_33855;
assign v_33859 = v_33857 & v_33858;
assign v_33862 = v_33860 & v_33861;
assign v_33865 = v_33863 & v_33864;
assign v_33868 = v_33866 & v_33867;
assign v_33871 = v_33869 & v_33870;
assign v_33874 = v_33872 & v_33873;
assign v_33877 = v_33875 & v_33876;
assign v_33880 = v_33878 & v_33879;
assign v_33883 = v_33881 & v_33882;
assign v_33886 = v_33884 & v_33885;
assign v_33889 = v_33887 & v_33888;
assign v_33892 = v_33890 & v_33891;
assign v_33895 = v_33893 & v_33894;
assign v_33898 = v_33896 & v_33897;
assign v_33901 = v_33899 & v_33900;
assign v_33904 = v_33902 & v_33903;
assign v_33907 = v_33905 & v_33906;
assign v_33910 = v_33908 & v_33909;
assign v_33913 = v_33911 & v_33912;
assign v_33916 = v_33914 & v_33915;
assign v_33919 = v_33917 & v_33918;
assign v_33922 = v_33920 & v_33921;
assign v_33925 = v_33923 & v_33924;
assign v_33928 = v_33926 & v_33927;
assign v_33931 = v_33929 & v_33930;
assign v_33934 = v_33932 & v_33933;
assign v_33937 = v_33935 & v_33936;
assign v_33940 = v_33938 & v_33939;
assign v_33943 = v_33941 & v_33942;
assign v_33946 = v_33944 & v_33945;
assign v_33949 = v_33947 & v_33948;
assign v_33952 = v_33950 & v_33951;
assign v_33955 = v_33953 & v_33954;
assign v_33958 = v_33956 & v_33957;
assign v_33961 = v_33959 & v_33960;
assign v_33964 = v_33962 & v_33963;
assign v_33967 = v_33965 & v_33966;
assign v_33970 = v_33968 & v_33969;
assign v_33973 = v_33971 & v_33972;
assign v_33976 = v_33974 & v_33975;
assign v_33979 = v_33977 & v_33978;
assign v_33982 = v_33980 & v_33981;
assign v_33985 = v_33983 & v_33984;
assign v_33988 = v_33986 & v_33987;
assign v_33991 = v_33989 & v_33990;
assign v_33994 = v_33992 & v_33993;
assign v_33997 = v_33995 & v_33996;
assign v_34000 = v_33998 & v_33999;
assign v_34003 = v_34001 & v_34002;
assign v_34006 = v_34004 & v_34005;
assign v_34009 = v_34007 & v_34008;
assign v_34012 = v_34010 & v_34011;
assign v_34015 = v_34013 & v_34014;
assign v_34018 = v_34016 & v_34017;
assign v_34019 = v_33829 & v_34018;
assign v_34022 = v_34020 & v_34021;
assign v_34025 = v_34023 & v_34024;
assign v_34028 = v_34026 & v_34027;
assign v_34031 = v_34029 & v_34030;
assign v_34034 = v_34032 & v_34033;
assign v_34037 = v_34035 & v_34036;
assign v_34040 = v_34038 & v_34039;
assign v_34043 = v_34041 & v_34042;
assign v_34046 = v_34044 & v_34045;
assign v_34049 = v_34047 & v_34048;
assign v_34052 = v_34050 & v_34051;
assign v_34055 = v_34053 & v_34054;
assign v_34058 = v_34056 & v_34057;
assign v_34061 = v_34059 & v_34060;
assign v_34064 = v_34062 & v_34063;
assign v_34067 = v_34065 & v_34066;
assign v_34070 = v_34068 & v_34069;
assign v_34073 = v_34071 & v_34072;
assign v_34076 = v_34074 & v_34075;
assign v_34079 = v_34077 & v_34078;
assign v_34082 = v_34080 & v_34081;
assign v_34085 = v_34083 & v_34084;
assign v_34088 = v_34086 & v_34087;
assign v_34091 = v_34089 & v_34090;
assign v_34094 = v_34092 & v_34093;
assign v_34097 = v_34095 & v_34096;
assign v_34100 = v_34098 & v_34099;
assign v_34103 = v_34101 & v_34102;
assign v_34106 = v_34104 & v_34105;
assign v_34109 = v_34107 & v_34108;
assign v_34112 = v_34110 & v_34111;
assign v_34115 = v_34113 & v_34114;
assign v_34118 = v_34116 & v_34117;
assign v_34121 = v_34119 & v_34120;
assign v_34124 = v_34122 & v_34123;
assign v_34127 = v_34125 & v_34126;
assign v_34130 = v_34128 & v_34129;
assign v_34133 = v_34131 & v_34132;
assign v_34136 = v_34134 & v_34135;
assign v_34139 = v_34137 & v_34138;
assign v_34142 = v_34140 & v_34141;
assign v_34145 = v_34143 & v_34144;
assign v_34148 = v_34146 & v_34147;
assign v_34151 = v_34149 & v_34150;
assign v_34154 = v_34152 & v_34153;
assign v_34157 = v_34155 & v_34156;
assign v_34160 = v_34158 & v_34159;
assign v_34163 = v_34161 & v_34162;
assign v_34166 = v_34164 & v_34165;
assign v_34169 = v_34167 & v_34168;
assign v_34172 = v_34170 & v_34171;
assign v_34175 = v_34173 & v_34174;
assign v_34178 = v_34176 & v_34177;
assign v_34181 = v_34179 & v_34180;
assign v_34184 = v_34182 & v_34183;
assign v_34187 = v_34185 & v_34186;
assign v_34190 = v_34188 & v_34189;
assign v_34193 = v_34191 & v_34192;
assign v_34196 = v_34194 & v_34195;
assign v_34199 = v_34197 & v_34198;
assign v_34202 = v_34200 & v_34201;
assign v_34205 = v_34203 & v_34204;
assign v_34208 = v_34206 & v_34207;
assign v_34209 = v_34019 & v_34208;
assign v_34212 = v_34210 & v_34211;
assign v_34215 = v_34213 & v_34214;
assign v_34218 = v_34216 & v_34217;
assign v_34221 = v_34219 & v_34220;
assign v_34224 = v_34222 & v_34223;
assign v_34227 = v_34225 & v_34226;
assign v_34230 = v_34228 & v_34229;
assign v_34233 = v_34231 & v_34232;
assign v_34236 = v_34234 & v_34235;
assign v_34239 = v_34237 & v_34238;
assign v_34242 = v_34240 & v_34241;
assign v_34245 = v_34243 & v_34244;
assign v_34248 = v_34246 & v_34247;
assign v_34251 = v_34249 & v_34250;
assign v_34254 = v_34252 & v_34253;
assign v_34257 = v_34255 & v_34256;
assign v_34260 = v_34258 & v_34259;
assign v_34263 = v_34261 & v_34262;
assign v_34266 = v_34264 & v_34265;
assign v_34269 = v_34267 & v_34268;
assign v_34272 = v_34270 & v_34271;
assign v_34275 = v_34273 & v_34274;
assign v_34278 = v_34276 & v_34277;
assign v_34281 = v_34279 & v_34280;
assign v_34284 = v_34282 & v_34283;
assign v_34287 = v_34285 & v_34286;
assign v_34290 = v_34288 & v_34289;
assign v_34293 = v_34291 & v_34292;
assign v_34296 = v_34294 & v_34295;
assign v_34299 = v_34297 & v_34298;
assign v_34302 = v_34300 & v_34301;
assign v_34305 = v_34303 & v_34304;
assign v_34308 = v_34306 & v_34307;
assign v_34311 = v_34309 & v_34310;
assign v_34314 = v_34312 & v_34313;
assign v_34317 = v_34315 & v_34316;
assign v_34320 = v_34318 & v_34319;
assign v_34323 = v_34321 & v_34322;
assign v_34326 = v_34324 & v_34325;
assign v_34329 = v_34327 & v_34328;
assign v_34332 = v_34330 & v_34331;
assign v_34335 = v_34333 & v_34334;
assign v_34338 = v_34336 & v_34337;
assign v_34341 = v_34339 & v_34340;
assign v_34344 = v_34342 & v_34343;
assign v_34347 = v_34345 & v_34346;
assign v_34350 = v_34348 & v_34349;
assign v_34353 = v_34351 & v_34352;
assign v_34356 = v_34354 & v_34355;
assign v_34359 = v_34357 & v_34358;
assign v_34362 = v_34360 & v_34361;
assign v_34365 = v_34363 & v_34364;
assign v_34368 = v_34366 & v_34367;
assign v_34371 = v_34369 & v_34370;
assign v_34374 = v_34372 & v_34373;
assign v_34377 = v_34375 & v_34376;
assign v_34380 = v_34378 & v_34379;
assign v_34383 = v_34381 & v_34382;
assign v_34386 = v_34384 & v_34385;
assign v_34389 = v_34387 & v_34388;
assign v_34392 = v_34390 & v_34391;
assign v_34395 = v_34393 & v_34394;
assign v_34398 = v_34396 & v_34397;
assign v_34399 = v_34209 & v_34398;
assign v_34402 = v_34400 & v_34401;
assign v_34405 = v_34403 & v_34404;
assign v_34408 = v_34406 & v_34407;
assign v_34411 = v_34409 & v_34410;
assign v_34414 = v_34412 & v_34413;
assign v_34417 = v_34415 & v_34416;
assign v_34420 = v_34418 & v_34419;
assign v_34423 = v_34421 & v_34422;
assign v_34426 = v_34424 & v_34425;
assign v_34429 = v_34427 & v_34428;
assign v_34432 = v_34430 & v_34431;
assign v_34435 = v_34433 & v_34434;
assign v_34438 = v_34436 & v_34437;
assign v_34441 = v_34439 & v_34440;
assign v_34444 = v_34442 & v_34443;
assign v_34447 = v_34445 & v_34446;
assign v_34450 = v_34448 & v_34449;
assign v_34453 = v_34451 & v_34452;
assign v_34456 = v_34454 & v_34455;
assign v_34459 = v_34457 & v_34458;
assign v_34462 = v_34460 & v_34461;
assign v_34465 = v_34463 & v_34464;
assign v_34468 = v_34466 & v_34467;
assign v_34471 = v_34469 & v_34470;
assign v_34474 = v_34472 & v_34473;
assign v_34477 = v_34475 & v_34476;
assign v_34480 = v_34478 & v_34479;
assign v_34483 = v_34481 & v_34482;
assign v_34486 = v_34484 & v_34485;
assign v_34489 = v_34487 & v_34488;
assign v_34492 = v_34490 & v_34491;
assign v_34495 = v_34493 & v_34494;
assign v_34498 = v_34496 & v_34497;
assign v_34501 = v_34499 & v_34500;
assign v_34504 = v_34502 & v_34503;
assign v_34507 = v_34505 & v_34506;
assign v_34510 = v_34508 & v_34509;
assign v_34513 = v_34511 & v_34512;
assign v_34516 = v_34514 & v_34515;
assign v_34519 = v_34517 & v_34518;
assign v_34522 = v_34520 & v_34521;
assign v_34525 = v_34523 & v_34524;
assign v_34528 = v_34526 & v_34527;
assign v_34531 = v_34529 & v_34530;
assign v_34534 = v_34532 & v_34533;
assign v_34537 = v_34535 & v_34536;
assign v_34540 = v_34538 & v_34539;
assign v_34543 = v_34541 & v_34542;
assign v_34546 = v_34544 & v_34545;
assign v_34549 = v_34547 & v_34548;
assign v_34552 = v_34550 & v_34551;
assign v_34555 = v_34553 & v_34554;
assign v_34558 = v_34556 & v_34557;
assign v_34561 = v_34559 & v_34560;
assign v_34564 = v_34562 & v_34563;
assign v_34567 = v_34565 & v_34566;
assign v_34570 = v_34568 & v_34569;
assign v_34573 = v_34571 & v_34572;
assign v_34576 = v_34574 & v_34575;
assign v_34579 = v_34577 & v_34578;
assign v_34582 = v_34580 & v_34581;
assign v_34585 = v_34583 & v_34584;
assign v_34588 = v_34586 & v_34587;
assign v_34589 = v_34399 & v_34588;
assign v_34590 = v_23366 & v_34589;
assign v_34593 = v_34591 & v_34592;
assign v_34596 = v_34594 & v_34595;
assign v_34599 = v_34597 & v_34598;
assign v_34602 = v_34600 & v_34601;
assign v_34605 = v_34603 & v_34604;
assign v_34608 = v_34606 & v_34607;
assign v_34611 = v_34609 & v_34610;
assign v_34614 = v_34612 & v_34613;
assign v_34617 = v_34615 & v_34616;
assign v_34620 = v_34618 & v_34619;
assign v_34623 = v_34621 & v_34622;
assign v_34626 = v_34624 & v_34625;
assign v_34629 = v_34627 & v_34628;
assign v_34632 = v_34630 & v_34631;
assign v_34635 = v_34633 & v_34634;
assign v_34638 = v_34636 & v_34637;
assign v_34641 = v_34639 & v_34640;
assign v_34644 = v_34642 & v_34643;
assign v_34647 = v_34645 & v_34646;
assign v_34650 = v_34648 & v_34649;
assign v_34653 = v_34651 & v_34652;
assign v_34656 = v_34654 & v_34655;
assign v_34659 = v_34657 & v_34658;
assign v_34662 = v_34660 & v_34661;
assign v_34665 = v_34663 & v_34664;
assign v_34668 = v_34666 & v_34667;
assign v_34671 = v_34669 & v_34670;
assign v_34674 = v_34672 & v_34673;
assign v_34677 = v_34675 & v_34676;
assign v_34680 = v_34678 & v_34679;
assign v_34683 = v_34681 & v_34682;
assign v_34686 = v_34684 & v_34685;
assign v_34689 = v_34687 & v_34688;
assign v_34692 = v_34690 & v_34691;
assign v_34695 = v_34693 & v_34694;
assign v_34698 = v_34696 & v_34697;
assign v_34701 = v_34699 & v_34700;
assign v_34704 = v_34702 & v_34703;
assign v_34707 = v_34705 & v_34706;
assign v_34710 = v_34708 & v_34709;
assign v_34713 = v_34711 & v_34712;
assign v_34716 = v_34714 & v_34715;
assign v_34719 = v_34717 & v_34718;
assign v_34722 = v_34720 & v_34721;
assign v_34725 = v_34723 & v_34724;
assign v_34728 = v_34726 & v_34727;
assign v_34731 = v_34729 & v_34730;
assign v_34734 = v_34732 & v_34733;
assign v_34737 = v_34735 & v_34736;
assign v_34740 = v_34738 & v_34739;
assign v_34743 = v_34741 & v_34742;
assign v_34746 = v_34744 & v_34745;
assign v_34749 = v_34747 & v_34748;
assign v_34752 = v_34750 & v_34751;
assign v_34755 = v_34753 & v_34754;
assign v_34758 = v_34756 & v_34757;
assign v_34761 = v_34759 & v_34760;
assign v_34764 = v_34762 & v_34763;
assign v_34767 = v_34765 & v_34766;
assign v_34770 = v_34768 & v_34769;
assign v_34773 = v_34771 & v_34772;
assign v_34776 = v_34774 & v_34775;
assign v_34779 = v_34777 & v_34778;
assign v_34780 = v_34590 & v_34779;
assign v_34781 = v_26290 & v_34780;
assign v_34782 = v_33450 & v_34781;
assign v_34783 = ~v_10462 & v_34782;
assign v_34785 = v_13342 & v_26092;
assign v_34786 = v_26282 & v_34785;
assign v_34787 = v_26290 & v_34786;
assign v_34788 = ~v_10462 & v_34787;
assign v_34790 = v_16391 & v_28952;
assign v_34791 = v_29142 & v_34790;
assign v_34792 = v_26290 & v_34791;
assign v_34793 = ~v_10462 & v_34792;
assign v_34795 = v_19364 & v_31739;
assign v_34796 = v_31926 & v_34795;
assign v_34797 = v_26290 & v_34796;
assign v_34798 = ~v_10462 & v_34797;
assign v_34800 = v_22403 & v_34589;
assign v_34801 = v_34779 & v_34800;
assign v_34802 = v_26290 & v_34801;
assign v_34803 = ~v_10462 & v_34802;
assign v_34805 = ~v_6094 & ~v_6122;
assign v_34806 = ~v_6003 & ~v_6034;
assign v_34807 = ~v_6046 & v_34806;
assign v_34808 = ~v_6058 & v_34807;
assign v_34809 = ~v_6070 & v_34808;
assign v_34810 = ~v_6082 & v_34809;
assign v_34811 = v_34805 & v_34810;
assign v_34812 = ~v_6824 & ~v_6852;
assign v_34813 = ~v_6720 & ~v_6764;
assign v_34814 = ~v_6776 & v_34813;
assign v_34815 = ~v_6788 & v_34814;
assign v_34816 = ~v_6800 & v_34815;
assign v_34817 = ~v_6812 & v_34816;
assign v_34818 = v_34812 & v_34817;
assign v_34819 = ~v_5806 & ~v_5834;
assign v_34820 = ~v_5715 & ~v_5746;
assign v_34821 = ~v_5758 & v_34820;
assign v_34822 = ~v_5770 & v_34821;
assign v_34823 = ~v_5782 & v_34822;
assign v_34824 = ~v_5794 & v_34823;
assign v_34825 = v_34819 & v_34824;
assign v_34826 = ~v_4263 & ~v_4294;
assign v_34827 = ~v_4306 & v_34826;
assign v_34828 = ~v_4318 & v_34827;
assign v_34829 = ~v_4330 & v_34828;
assign v_34830 = ~v_4342 & v_34829;
assign v_34831 = v_4354 & v_34830;
assign v_34832 = ~v_4382 & v_34831;
assign v_34833 = v_26290 & v_34832;
assign v_34834 = v_34825 & v_34833;
assign v_34835 = v_34818 & v_34834;
assign v_34836 = v_34811 & v_34835;
assign v_34837 = ~v_10462 & v_34836;
assign v_34839 = ~v_10462 & v_34838;
assign v_34840 = v_34804 & v_34839;
assign v_34841 = v_34799 & v_34840;
assign v_34842 = v_34794 & v_34841;
assign v_34843 = v_34789 & v_34842;
assign v_34844 = v_34784 & v_34843;
assign v_34845 = v_31931 & v_34844;
assign v_34846 = v_29147 & v_34845;
assign v_34847 = v_26294 & v_34846;
assign v_34848 = v_23434 & v_34847;
assign v_34849 = v_23433 & v_34848;
assign v_34850 = ~v_3 & v_34849;
assign v_34853 = v_4 & v_26289;
assign v_34854 = ~v_3 & v_34853;
assign v_34859 = ~v_34852;
assign v_34861 = v_34859 & v_34860;
assign v_34862 = v_35133 & v_35134;
assign v_34864 = v_566 & v_719 & v_725 & v_729 & v_735;
assign v_34865 = v_739 & v_745 & v_749 & v_755 & v_759;
assign v_34866 = v_765 & v_769 & v_781 & v_791 & v_797;
assign v_34867 = v_801 & v_820 & v_836 & v_843 & v_848;
assign v_34868 = v_855 & v_860 & v_867 & v_872 & v_879;
assign v_34869 = v_884 & v_891 & v_896 & v_909 & v_920;
assign v_34870 = v_927 & v_932 & v_958 & v_982 & v_989;
assign v_34871 = v_994 & v_1001 & v_1006 & v_1013 & v_1018;
assign v_34872 = v_1025 & v_1030 & v_1037 & v_1042 & v_1057;
assign v_34873 = v_1070 & v_1077 & v_1082 & v_1099 & v_1114;
assign v_34874 = v_1121 & v_1126 & v_1133 & v_1138 & v_1145;
assign v_34875 = v_1150 & v_1157 & v_1162 & v_1169 & v_1174;
assign v_34876 = v_1189 & v_1202 & v_1209 & v_1214 & v_1243;
assign v_34877 = v_1270 & v_1277 & v_1282 & v_1289 & v_1294;
assign v_34878 = v_1301 & v_1306 & v_1313 & v_1318 & v_1325;
assign v_34879 = v_1330 & v_1345 & v_1358 & v_1365 & v_1370;
assign v_34880 = v_1387 & v_1402 & v_1409 & v_1414 & v_1421;
assign v_34881 = v_1426 & v_1433 & v_1438 & v_1445 & v_1450;
assign v_34882 = v_1457 & v_1462 & v_1477 & v_1490 & v_1497;
assign v_34883 = v_1502 & v_1529 & v_1554 & v_1561 & v_1566;
assign v_34884 = v_1573 & v_1578 & v_1585 & v_1590 & v_1597;
assign v_34885 = v_1602 & v_1609 & v_1614 & v_1629 & v_1642;
assign v_34886 = v_1649 & v_1654 & v_1671 & v_1686 & v_1693;
assign v_34887 = v_1698 & v_1705 & v_1710 & v_1717 & v_1722;
assign v_34888 = v_1729 & v_1734 & v_1741 & v_1746 & v_1761;
assign v_34889 = v_1774 & v_1781 & v_1786 & v_1819 & v_1850;
assign v_34890 = v_1857 & v_1862 & v_1869 & v_1874 & v_1881;
assign v_34891 = v_1886 & v_1893 & v_1898 & v_1905 & v_1910;
assign v_34892 = v_1925 & v_1938 & v_1945 & v_1950 & v_1967;
assign v_34893 = v_1982 & v_1989 & v_1994 & v_2001 & v_2006;
assign v_34894 = v_2013 & v_2018 & v_2025 & v_2030 & v_2037;
assign v_34895 = v_2042 & v_2057 & v_2070 & v_2077 & v_2082;
assign v_34896 = v_2108 & v_2132 & v_2139 & v_2144 & v_2151;
assign v_34897 = v_2156 & v_2163 & v_2168 & v_2175 & v_2180;
assign v_34898 = v_2187 & v_2192 & v_2207 & v_2220 & v_2227;
assign v_34899 = v_2232 & v_2249 & v_2264 & v_2271 & v_2276;
assign v_34900 = v_2283 & v_2288 & v_2295 & v_2300 & v_2307;
assign v_34901 = v_2312 & v_2319 & v_2324 & v_2339 & v_2352;
assign v_34902 = v_2359 & v_2364 & v_2393 & v_2420 & v_2427;
assign v_34903 = v_2432 & v_2439 & v_2444 & v_2451 & v_2456;
assign v_34904 = v_2463 & v_2468 & v_2475 & v_2480 & v_2495;
assign v_34905 = v_2508 & v_2515 & v_2520 & v_2537 & v_2552;
assign v_34906 = v_2559 & v_2564 & v_2571 & v_2576 & v_2583;
assign v_34907 = v_2588 & v_2595 & v_2600 & v_2607 & v_2612;
assign v_34908 = v_2627 & v_2640 & v_2647 & v_2652 & v_2680;
assign v_34909 = v_2706 & v_2713 & v_2718 & v_2725 & v_2730;
assign v_34910 = v_2737 & v_2742 & v_2749 & v_2754 & v_2761;
assign v_34911 = v_2766 & v_2781 & v_2794 & v_2801 & v_2806;
assign v_34912 = v_2823 & v_2838 & v_2845 & v_2850 & v_2857;
assign v_34913 = v_2862 & v_2869 & v_2874 & v_2881 & v_2886;
assign v_34914 = v_2893 & v_2898 & v_2913 & v_2926 & v_2933;
assign v_34915 = v_2938 & v_2975 & v_3010 & v_3017 & v_3022;
assign v_34916 = v_3029 & v_3034 & v_3041 & v_3046 & v_3053;
assign v_34917 = v_3058 & v_3065 & v_3070 & v_3085 & v_3098;
assign v_34918 = v_3105 & v_3110 & v_3127 & v_3142 & v_3149;
assign v_34919 = v_3154 & v_3161 & v_3166 & v_3173 & v_3178;
assign v_34920 = v_3185 & v_3190 & v_3197 & v_3202 & v_3217;
assign v_34921 = v_3230 & v_3237 & v_3242 & v_3268 & v_3292;
assign v_34922 = v_3299 & v_3304 & v_3311 & v_3316 & v_3323;
assign v_34923 = v_3328 & v_3335 & v_3340 & v_3347 & v_3352;
assign v_34924 = v_3367 & v_3380 & v_3387 & v_3392 & v_3409;
assign v_34925 = v_3424 & v_3431 & v_3436 & v_3443 & v_3448;
assign v_34926 = v_3455 & v_3460 & v_3467 & v_3472 & v_3479;
assign v_34927 = v_3484 & v_3499 & v_3512 & v_3519 & v_3524;
assign v_34928 = v_3553 & v_3580 & v_3587 & v_3592 & v_3599;
assign v_34929 = v_3604 & v_3611 & v_3616 & v_3623 & v_3628;
assign v_34930 = v_3635 & v_3640 & v_3655 & v_3668 & v_3675;
assign v_34931 = v_3680 & v_3697 & v_3712 & v_3719 & v_3724;
assign v_34932 = v_3731 & v_3736 & v_3743 & v_3748 & v_3755;
assign v_34933 = v_3760 & v_3767 & v_3772 & v_3787 & v_3800;
assign v_34934 = v_3807 & v_3812 & v_3839 & v_3864 & v_3871;
assign v_34935 = v_3876 & v_3883 & v_3888 & v_3895 & v_3900;
assign v_34936 = v_3907 & v_3912 & v_3919 & v_3924 & v_3939;
assign v_34937 = v_3952 & v_3959 & v_3964 & v_3981 & v_3996;
assign v_34938 = v_4003 & v_4008 & v_4015 & v_4020 & v_4027;
assign v_34939 = v_4032 & v_4039 & v_4044 & v_4051 & v_4056;
assign v_34940 = v_4071 & v_4084 & v_4091 & v_4096 & v_4129;
assign v_34941 = v_4160 & v_4167 & v_4172 & v_4179 & v_4184;
assign v_34942 = v_4191 & v_4196 & v_4203 & v_4208 & v_4215;
assign v_34943 = v_4220 & v_4235 & v_4248 & v_4255 & v_4260;
assign v_34944 = v_4277 & v_4292 & v_4299 & v_4304 & v_4311;
assign v_34945 = v_4316 & v_4323 & v_4328 & v_4335 & v_4340;
assign v_34946 = v_4347 & v_4352 & v_4367 & v_4380 & v_4387;
assign v_34947 = v_4392 & v_4418 & v_4442 & v_4449 & v_4454;
assign v_34948 = v_4461 & v_4466 & v_4473 & v_4478 & v_4485;
assign v_34949 = v_4490 & v_4497 & v_4502 & v_4517 & v_4530;
assign v_34950 = v_4537 & v_4542 & v_4559 & v_4574 & v_4581;
assign v_34951 = v_4586 & v_4593 & v_4598 & v_4605 & v_4610;
assign v_34952 = v_4617 & v_4622 & v_4629 & v_4634 & v_4649;
assign v_34953 = v_4662 & v_4669 & v_4674 & v_4703 & v_4730;
assign v_34954 = v_4737 & v_4742 & v_4749 & v_4754 & v_4761;
assign v_34955 = v_4766 & v_4773 & v_4778 & v_4785 & v_4790;
assign v_34956 = v_4805 & v_4818 & v_4825 & v_4830 & v_4847;
assign v_34957 = v_4862 & v_4869 & v_4874 & v_4881 & v_4886;
assign v_34958 = v_4893 & v_4898 & v_4905 & v_4910 & v_4917;
assign v_34959 = v_4922 & v_4937 & v_4950 & v_4957 & v_4962;
assign v_34960 = v_4991 & v_5018 & v_5025 & v_5030 & v_5037;
assign v_34961 = v_5042 & v_5049 & v_5054 & v_5061 & v_5066;
assign v_34962 = v_5073 & v_5078 & v_5093 & v_5106 & v_5113;
assign v_34963 = v_5118 & v_5135 & v_5150 & v_5157 & v_5162;
assign v_34964 = v_5169 & v_5174 & v_5181 & v_5186 & v_5193;
assign v_34965 = v_5198 & v_5205 & v_5210 & v_5225 & v_5238;
assign v_34966 = v_5245 & v_5250 & v_5291 & v_5330 & v_5337;
assign v_34967 = v_5342 & v_5349 & v_5354 & v_5361 & v_5366;
assign v_34968 = v_5373 & v_5378 & v_5385 & v_5390 & v_5405;
assign v_34969 = v_5418 & v_5425 & v_5430 & v_5447 & v_5462;
assign v_34970 = v_5469 & v_5474 & v_5481 & v_5486 & v_5493;
assign v_34971 = v_5498 & v_5505 & v_5510 & v_5517 & v_5522;
assign v_34972 = v_5537 & v_5550 & v_5557 & v_5562 & v_5588;
assign v_34973 = v_5612 & v_5619 & v_5624 & v_5631 & v_5636;
assign v_34974 = v_5643 & v_5648 & v_5655 & v_5660 & v_5667;
assign v_34975 = v_5672 & v_5687 & v_5700 & v_5707 & v_5712;
assign v_34976 = v_5729 & v_5744 & v_5751 & v_5756 & v_5763;
assign v_34977 = v_5768 & v_5775 & v_5780 & v_5787 & v_5792;
assign v_34978 = v_5799 & v_5804 & v_5819 & v_5832 & v_5839;
assign v_34979 = v_5844 & v_5873 & v_5900 & v_5907 & v_5912;
assign v_34980 = v_5919 & v_5924 & v_5931 & v_5936 & v_5943;
assign v_34981 = v_5948 & v_5955 & v_5960 & v_5975 & v_5988;
assign v_34982 = v_5995 & v_6000 & v_6017 & v_6032 & v_6039;
assign v_34983 = v_6044 & v_6051 & v_6056 & v_6063 & v_6068;
assign v_34984 = v_6075 & v_6080 & v_6087 & v_6092 & v_6107;
assign v_34985 = v_6120 & v_6127 & v_6132 & v_6159 & v_6184;
assign v_34986 = v_6191 & v_6196 & v_6203 & v_6208 & v_6215;
assign v_34987 = v_6220 & v_6227 & v_6232 & v_6239 & v_6244;
assign v_34988 = v_6259 & v_6272 & v_6279 & v_6284 & v_6301;
assign v_34989 = v_6316 & v_6323 & v_6328 & v_6335 & v_6340;
assign v_34990 = v_6347 & v_6352 & v_6359 & v_6364 & v_6371;
assign v_34991 = v_6376 & v_6391 & v_6404 & v_6411 & v_6416;
assign v_34992 = v_6449 & v_6480 & v_6487 & v_6492 & v_6499;
assign v_34993 = v_6504 & v_6511 & v_6516 & v_6523 & v_6528;
assign v_34994 = v_6535 & v_6540 & v_6555 & v_6568 & v_6575;
assign v_34995 = v_6580 & v_6597 & v_6612 & v_6619 & v_6624;
assign v_34996 = v_6631 & v_6636 & v_6643 & v_6648 & v_6655;
assign v_34997 = v_6660 & v_6667 & v_6672 & v_6687 & v_6700;
assign v_34998 = v_6707 & v_6712 & v_6738 & v_6762 & v_6769;
assign v_34999 = v_6774 & v_6781 & v_6786 & v_6793 & v_6798;
assign v_35000 = v_6805 & v_6810 & v_6817 & v_6822 & v_6837;
assign v_35001 = v_6850 & v_6857 & v_6862 & v_6879 & v_6894;
assign v_35002 = v_6901 & v_6906 & v_6913 & v_6918 & v_6925;
assign v_35003 = v_6930 & v_6937 & v_6942 & v_6949 & v_6954;
assign v_35004 = v_6969 & v_6982 & v_6989 & v_6994 & v_7023;
assign v_35005 = v_7050 & v_7057 & v_7062 & v_7069 & v_7074;
assign v_35006 = v_7081 & v_7086 & v_7093 & v_7098 & v_7105;
assign v_35007 = v_7110 & v_7125 & v_7138 & v_7145 & v_7150;
assign v_35008 = v_7167 & v_7182 & v_7189 & v_7194 & v_7201;
assign v_35009 = v_7206 & v_7213 & v_7218 & v_7225 & v_7230;
assign v_35010 = v_7237 & v_7242 & v_7257 & v_7270 & v_7277;
assign v_35011 = v_7282 & v_7310 & v_7336 & v_7343 & v_7348;
assign v_35012 = v_7355 & v_7360 & v_7367 & v_7372 & v_7379;
assign v_35013 = v_7384 & v_7391 & v_7396 & v_7411 & v_7424;
assign v_35014 = v_7431 & v_7436 & v_7453 & v_7468 & v_7475;
assign v_35015 = v_7480 & v_7487 & v_7492 & v_7499 & v_7504;
assign v_35016 = v_7511 & v_7516 & v_7523 & v_7528 & v_7543;
assign v_35017 = v_7556 & v_7563 & v_7568 & v_7605 & v_7640;
assign v_35018 = v_7647 & v_7652 & v_7659 & v_7664 & v_7671;
assign v_35019 = v_7676 & v_7683 & v_7688 & v_7695 & v_7700;
assign v_35020 = v_7715 & v_7728 & v_7735 & v_7740 & v_7757;
assign v_35021 = v_7772 & v_7779 & v_7784 & v_7791 & v_7796;
assign v_35022 = v_7803 & v_7808 & v_7815 & v_7820 & v_7827;
assign v_35023 = v_7832 & v_7847 & v_7860 & v_7867 & v_7872;
assign v_35024 = v_7898 & v_7922 & v_7929 & v_7934 & v_7941;
assign v_35025 = v_7946 & v_7953 & v_7958 & v_7965 & v_7970;
assign v_35026 = v_7977 & v_7982 & v_7997 & v_8010 & v_8017;
assign v_35027 = v_8022 & v_8039 & v_8054 & v_8061 & v_8066;
assign v_35028 = v_8073 & v_8078 & v_8085 & v_8090 & v_8097;
assign v_35029 = v_8102 & v_8109 & v_8114 & v_8129 & v_8142;
assign v_35030 = v_8149 & v_8154 & v_8183 & v_8210 & v_8217;
assign v_35031 = v_8222 & v_8229 & v_8234 & v_8241 & v_8246;
assign v_35032 = v_8253 & v_8258 & v_8265 & v_8270 & v_8285;
assign v_35033 = v_8298 & v_8305 & v_8310 & v_8327 & v_8342;
assign v_35034 = v_8349 & v_8354 & v_8361 & v_8366 & v_8373;
assign v_35035 = v_8378 & v_8385 & v_8390 & v_8397 & v_8402;
assign v_35036 = v_8417 & v_8430 & v_8437 & v_8442 & v_8469;
assign v_35037 = v_8494 & v_8501 & v_8506 & v_8513 & v_8518;
assign v_35038 = v_8525 & v_8530 & v_8537 & v_8542 & v_8549;
assign v_35039 = v_8554 & v_8569 & v_8582 & v_8589 & v_8594;
assign v_35040 = v_8611 & v_8626 & v_8633 & v_8638 & v_8645;
assign v_35041 = v_8650 & v_8657 & v_8662 & v_8669 & v_8674;
assign v_35042 = v_8681 & v_8686 & v_8701 & v_8714 & v_8721;
assign v_35043 = v_8726 & v_8759 & v_8790 & v_8797 & v_8802;
assign v_35044 = v_8809 & v_8814 & v_8821 & v_8826 & v_8833;
assign v_35045 = v_8838 & v_8845 & v_8850 & v_8865 & v_8878;
assign v_35046 = v_8885 & v_8890 & v_8907 & v_8922 & v_8929;
assign v_35047 = v_8934 & v_8941 & v_8946 & v_8953 & v_8958;
assign v_35048 = v_8965 & v_8970 & v_8977 & v_8982 & v_8997;
assign v_35049 = v_9010 & v_9017 & v_9022 & v_9048 & v_9072;
assign v_35050 = v_9079 & v_9084 & v_9091 & v_9096 & v_9103;
assign v_35051 = v_9108 & v_9115 & v_9120 & v_9127 & v_9132;
assign v_35052 = v_9147 & v_9160 & v_9167 & v_9172 & v_9189;
assign v_35053 = v_9204 & v_9211 & v_9216 & v_9223 & v_9228;
assign v_35054 = v_9235 & v_9240 & v_9247 & v_9252 & v_9259;
assign v_35055 = v_9264 & v_9279 & v_9292 & v_9299 & v_9304;
assign v_35056 = v_9333 & v_9360 & v_9367 & v_9372 & v_9379;
assign v_35057 = v_9384 & v_9391 & v_9396 & v_9403 & v_9408;
assign v_35058 = v_9415 & v_9420 & v_9435 & v_9448 & v_9455;
assign v_35059 = v_9460 & v_9477 & v_9492 & v_9499 & v_9504;
assign v_35060 = v_9511 & v_9516 & v_9523 & v_9528 & v_9535;
assign v_35061 = v_9540 & v_9547 & v_9552 & v_9567 & v_9580;
assign v_35062 = v_9587 & v_9592 & v_9622 & v_9650 & v_9657;
assign v_35063 = v_9662 & v_9669 & v_9674 & v_9681 & v_9686;
assign v_35064 = v_9693 & v_9698 & v_9705 & v_9710 & v_9725;
assign v_35065 = v_9738 & v_9745 & v_9750 & v_9767 & v_9782;
assign v_35066 = v_9789 & v_9794 & v_9801 & v_9806 & v_9813;
assign v_35067 = v_9818 & v_9825 & v_9830 & v_9837 & v_9842;
assign v_35068 = v_9857 & v_9870 & v_9877 & v_9882 & v_9928;
assign v_35069 = v_9947 & v_9966 & v_9984 & v_10003 & v_10021;
assign v_35070 = v_10040 & v_10058 & v_10077 & v_10095 & v_10114;
assign v_35071 = v_10132 & v_10150 & v_10167 & v_10181 & v_10194;
assign v_35072 = v_10210 & v_10223 & v_10237 & v_10250 & v_10264;
assign v_35073 = v_10277 & v_10291 & v_10304 & v_10318 & v_10331;
assign v_35074 = v_10345 & v_10358 & v_10372 & v_10385 & v_10399;
assign v_35075 = v_10412 & v_10417 & v_10419 & v_10423 & v_10425;
assign v_35076 = v_10429 & v_10431 & v_10435 & v_10437 & v_10441;
assign v_35077 = v_10443 & v_10447 & v_10449 & v_10453 & v_10455;
assign v_35078 = v_10458 & v_10460 & v_10463 & v_10464 & v_23418;
assign v_35079 = v_34851 & v_34855 & v_34858 & v_34861;
assign v_35080 = v_34864 & v_34865 & v_34866 & v_34867 & v_34868;
assign v_35081 = v_34869 & v_34870 & v_34871 & v_34872 & v_34873;
assign v_35082 = v_34874 & v_34875 & v_34876 & v_34877 & v_34878;
assign v_35083 = v_34879 & v_34880 & v_34881 & v_34882 & v_34883;
assign v_35084 = v_34884 & v_34885 & v_34886 & v_34887 & v_34888;
assign v_35085 = v_34889 & v_34890 & v_34891 & v_34892 & v_34893;
assign v_35086 = v_34894 & v_34895 & v_34896 & v_34897 & v_34898;
assign v_35087 = v_34899 & v_34900 & v_34901 & v_34902 & v_34903;
assign v_35088 = v_34904 & v_34905 & v_34906 & v_34907 & v_34908;
assign v_35089 = v_34909 & v_34910 & v_34911 & v_34912 & v_34913;
assign v_35090 = v_34914 & v_34915 & v_34916 & v_34917 & v_34918;
assign v_35091 = v_34919 & v_34920 & v_34921 & v_34922 & v_34923;
assign v_35092 = v_34924 & v_34925 & v_34926 & v_34927 & v_34928;
assign v_35093 = v_34929 & v_34930 & v_34931 & v_34932 & v_34933;
assign v_35094 = v_34934 & v_34935 & v_34936 & v_34937 & v_34938;
assign v_35095 = v_34939 & v_34940 & v_34941 & v_34942 & v_34943;
assign v_35096 = v_34944 & v_34945 & v_34946 & v_34947 & v_34948;
assign v_35097 = v_34949 & v_34950 & v_34951 & v_34952 & v_34953;
assign v_35098 = v_34954 & v_34955 & v_34956 & v_34957 & v_34958;
assign v_35099 = v_34959 & v_34960 & v_34961 & v_34962 & v_34963;
assign v_35100 = v_34964 & v_34965 & v_34966 & v_34967 & v_34968;
assign v_35101 = v_34969 & v_34970 & v_34971 & v_34972 & v_34973;
assign v_35102 = v_34974 & v_34975 & v_34976 & v_34977 & v_34978;
assign v_35103 = v_34979 & v_34980 & v_34981 & v_34982 & v_34983;
assign v_35104 = v_34984 & v_34985 & v_34986 & v_34987 & v_34988;
assign v_35105 = v_34989 & v_34990 & v_34991 & v_34992 & v_34993;
assign v_35106 = v_34994 & v_34995 & v_34996 & v_34997 & v_34998;
assign v_35107 = v_34999 & v_35000 & v_35001 & v_35002 & v_35003;
assign v_35108 = v_35004 & v_35005 & v_35006 & v_35007 & v_35008;
assign v_35109 = v_35009 & v_35010 & v_35011 & v_35012 & v_35013;
assign v_35110 = v_35014 & v_35015 & v_35016 & v_35017 & v_35018;
assign v_35111 = v_35019 & v_35020 & v_35021 & v_35022 & v_35023;
assign v_35112 = v_35024 & v_35025 & v_35026 & v_35027 & v_35028;
assign v_35113 = v_35029 & v_35030 & v_35031 & v_35032 & v_35033;
assign v_35114 = v_35034 & v_35035 & v_35036 & v_35037 & v_35038;
assign v_35115 = v_35039 & v_35040 & v_35041 & v_35042 & v_35043;
assign v_35116 = v_35044 & v_35045 & v_35046 & v_35047 & v_35048;
assign v_35117 = v_35049 & v_35050 & v_35051 & v_35052 & v_35053;
assign v_35118 = v_35054 & v_35055 & v_35056 & v_35057 & v_35058;
assign v_35119 = v_35059 & v_35060 & v_35061 & v_35062 & v_35063;
assign v_35120 = v_35064 & v_35065 & v_35066 & v_35067 & v_35068;
assign v_35121 = v_35069 & v_35070 & v_35071 & v_35072 & v_35073;
assign v_35122 = v_35074 & v_35075 & v_35076 & v_35077 & v_35078;
assign v_35123 = v_35079;
assign v_35124 = v_35080 & v_35081 & v_35082 & v_35083 & v_35084;
assign v_35125 = v_35085 & v_35086 & v_35087 & v_35088 & v_35089;
assign v_35126 = v_35090 & v_35091 & v_35092 & v_35093 & v_35094;
assign v_35127 = v_35095 & v_35096 & v_35097 & v_35098 & v_35099;
assign v_35128 = v_35100 & v_35101 & v_35102 & v_35103 & v_35104;
assign v_35129 = v_35105 & v_35106 & v_35107 & v_35108 & v_35109;
assign v_35130 = v_35110 & v_35111 & v_35112 & v_35113 & v_35114;
assign v_35131 = v_35115 & v_35116 & v_35117 & v_35118 & v_35119;
assign v_35132 = v_35120 & v_35121 & v_35122 & v_35123;
assign v_35133 = v_35124 & v_35125 & v_35126 & v_35127 & v_35128;
assign v_35134 = v_35129 & v_35130 & v_35131 & v_35132;
assign v_6 = v_2 | v_5;
assign v_10 = v_8 | v_9;
assign v_11 = ~v_8 | ~v_9;
assign v_15 = v_13 | v_14;
assign v_16 = ~v_13 | ~v_14;
assign v_20 = ~v_18 | v_19;
assign v_21 = v_18 | ~v_19;
assign v_25 = ~v_23 | v_24;
assign v_26 = v_23 | ~v_24;
assign v_33 = v_31 | v_32;
assign v_36 = v_34 | v_35;
assign v_39 = v_37 | v_38;
assign v_42 = v_40 | v_41;
assign v_48 = v_46 | v_47;
assign v_49 = v_44 | v_45;
assign v_50 = v_48 | v_49;
assign v_51 = v_42 | v_43;
assign v_53 = v_41 | v_52;
assign v_55 = v_38 | v_54;
assign v_57 = v_35 | v_56;
assign v_59 = v_32 | v_58;
assign v_60 = ~v_28 | ~v_29;
assign v_61 = v_59 | v_60;
assign v_63 = v_57 | v_62;
assign v_65 = v_55 | v_64;
assign v_67 = v_53 | v_66;
assign v_69 = ~v_43 | v_68;
assign v_71 = v_50 | v_70;
assign v_72 = v_12 | v_39;
assign v_74 = v_71 | v_73;
assign v_75 = v_17 | v_36;
assign v_77 = v_74 | v_76;
assign v_78 = v_22 | v_33;
assign v_80 = v_77 | v_79;
assign v_81 = v_27 | v_30;
assign v_83 = v_80 | v_82;
assign v_84 = v_28 | v_29;
assign v_86 = v_83 | v_85;
assign v_88 = v_86 | ~v_87;
assign v_90 = v_88 | ~v_89;
assign v_92 = v_90 | v_91;
assign v_93 = v_88 | v_89;
assign v_94 = ~v_91 | v_93;
assign v_97 = v_95 | ~v_96;
assign v_107 = ~v_18 | ~v_23;
assign v_108 = v_13 | v_107;
assign v_109 = v_8 | v_108;
assign v_110 = v_43 | v_109;
assign v_111 = v_45 | v_110;
assign v_113 = v_106 | v_112;
assign v_116 = v_114 | v_115;
assign v_119 = v_117 | v_118;
assign v_121 = ~v_8 | v_108;
assign v_122 = v_8 | v_101;
assign v_125 = v_120 | v_124;
assign v_128 = v_126 | v_127;
assign v_130 = ~v_13 | v_107;
assign v_131 = v_13 | v_100;
assign v_134 = v_129 | v_133;
assign v_137 = v_135 | v_136;
assign v_139 = v_18 | ~v_23;
assign v_140 = ~v_18 | v_23;
assign v_143 = v_138 | v_142;
assign v_146 = v_144 | v_145;
assign v_147 = v_60 | v_146;
assign v_148 = ~v_23 | ~v_24;
assign v_150 = v_143 | v_149;
assign v_151 = ~v_19 | v_137;
assign v_153 = v_134 | v_152;
assign v_154 = ~v_14 | v_128;
assign v_156 = v_125 | v_155;
assign v_157 = ~v_9 | v_119;
assign v_161 = v_159 | v_160;
assign v_162 = v_158 | v_161;
assign v_163 = v_116 | v_162;
assign v_164 = v_113 | v_163;
assign v_166 = ~v_47 | v_111;
assign v_167 = v_47 | v_104;
assign v_169 = ~v_45 | v_110;
assign v_170 = v_45 | v_103;
assign v_172 = v_9 | v_123;
assign v_174 = v_14 | v_132;
assign v_176 = v_19 | v_141;
assign v_178 = v_23 | v_24;
assign v_181 = v_145 | v_180;
assign v_183 = v_142 | v_182;
assign v_185 = v_133 | v_184;
assign v_187 = v_124 | v_186;
assign v_188 = ~v_43 | v_109;
assign v_189 = v_43 | v_102;
assign v_194 = v_105 | v_193;
assign v_195 = v_47 | v_111;
assign v_196 = v_164 | v_195;
assign v_198 = v_165 | v_197;
assign v_199 = v_168 | v_192;
assign v_201 = v_198 | v_200;
assign v_202 = v_171 | v_191;
assign v_204 = v_201 | v_203;
assign v_205 = v_187 | v_190;
assign v_207 = v_204 | v_206;
assign v_208 = v_173 | v_185;
assign v_210 = v_207 | v_209;
assign v_211 = v_175 | v_183;
assign v_213 = v_210 | v_212;
assign v_214 = v_177 | v_181;
assign v_216 = v_213 | v_215;
assign v_217 = v_30 | v_179;
assign v_219 = v_216 | v_218;
assign v_220 = v_85 | v_219;
assign v_221 = ~v_87 | v_220;
assign v_222 = v_89 | v_221;
assign v_223 = v_91 | v_222;
assign v_232 = ~v_23 | v_28;
assign v_233 = ~v_18 | v_232;
assign v_234 = v_13 | v_233;
assign v_235 = v_8 | v_234;
assign v_236 = v_43 | v_235;
assign v_237 = v_45 | v_236;
assign v_239 = v_231 | v_238;
assign v_242 = v_240 | v_241;
assign v_245 = v_243 | v_244;
assign v_247 = ~v_8 | v_234;
assign v_248 = v_8 | v_226;
assign v_251 = v_246 | v_250;
assign v_254 = v_252 | v_253;
assign v_256 = ~v_13 | v_233;
assign v_257 = v_13 | v_225;
assign v_260 = v_255 | v_259;
assign v_263 = v_261 | v_262;
assign v_265 = v_18 | v_232;
assign v_266 = ~v_18 | v_224;
assign v_269 = v_264 | v_268;
assign v_272 = v_270 | v_271;
assign v_274 = v_23 | v_28;
assign v_275 = ~v_23 | ~v_28;
assign v_278 = v_273 | v_277;
assign v_279 = v_28 | ~v_29;
assign v_280 = v_278 | v_279;
assign v_281 = ~v_24 | v_272;
assign v_283 = v_269 | v_282;
assign v_284 = ~v_19 | v_263;
assign v_286 = v_260 | v_285;
assign v_287 = ~v_14 | v_254;
assign v_289 = v_251 | v_288;
assign v_290 = ~v_9 | v_245;
assign v_294 = v_292 | v_293;
assign v_295 = v_291 | v_294;
assign v_296 = v_242 | v_295;
assign v_297 = v_239 | v_296;
assign v_299 = ~v_47 | v_237;
assign v_300 = v_47 | v_229;
assign v_302 = ~v_45 | v_236;
assign v_303 = v_45 | v_228;
assign v_305 = v_9 | v_249;
assign v_307 = v_14 | v_258;
assign v_309 = v_19 | v_267;
assign v_311 = v_24 | v_276;
assign v_315 = v_277 | v_314;
assign v_317 = v_268 | v_316;
assign v_319 = v_259 | v_318;
assign v_321 = v_250 | v_320;
assign v_322 = ~v_43 | v_235;
assign v_323 = v_43 | v_227;
assign v_328 = v_230 | v_327;
assign v_329 = v_47 | v_237;
assign v_330 = v_297 | v_329;
assign v_332 = v_298 | v_331;
assign v_333 = v_301 | v_326;
assign v_335 = v_332 | v_334;
assign v_336 = v_304 | v_325;
assign v_338 = v_335 | v_337;
assign v_339 = v_321 | v_324;
assign v_341 = v_338 | v_340;
assign v_342 = v_306 | v_319;
assign v_344 = v_341 | v_343;
assign v_345 = v_308 | v_317;
assign v_347 = v_344 | v_346;
assign v_348 = v_310 | v_315;
assign v_350 = v_347 | v_349;
assign v_351 = v_312 | v_313;
assign v_353 = v_350 | v_352;
assign v_354 = ~v_28 | v_29;
assign v_356 = v_353 | v_355;
assign v_357 = ~v_87 | v_356;
assign v_358 = v_89 | v_357;
assign v_359 = v_91 | v_358;
assign v_362 = v_360 | ~v_361;
assign v_369 = v_47 | v_368;
assign v_370 = v_18 | v_23;
assign v_371 = ~v_13 | v_370;
assign v_372 = ~v_8 | v_371;
assign v_373 = ~v_43 | v_372;
assign v_374 = ~v_45 | v_373;
assign v_375 = ~v_47 | v_374;
assign v_377 = v_45 | v_367;
assign v_379 = v_8 | v_365;
assign v_381 = v_9 | v_380;
assign v_383 = v_366 | v_382;
assign v_384 = ~v_9 | v_383;
assign v_386 = v_13 | v_364;
assign v_388 = v_14 | v_387;
assign v_390 = v_365 | v_389;
assign v_391 = ~v_14 | v_390;
assign v_394 = v_19 | v_393;
assign v_395 = v_100 | v_364;
assign v_396 = ~v_19 | v_395;
assign v_400 = v_398 | v_399;
assign v_403 = v_401 | v_402;
assign v_406 = v_404 | v_405;
assign v_407 = v_43 | v_366;
assign v_413 = v_411 | v_412;
assign v_414 = v_376 | v_410;
assign v_415 = v_413 | v_414;
assign v_416 = v_378 | v_409;
assign v_418 = v_368 | v_417;
assign v_420 = v_405 | v_419;
assign v_422 = v_402 | v_421;
assign v_424 = v_399 | v_423;
assign v_425 = v_149 | v_424;
assign v_427 = v_422 | v_426;
assign v_429 = v_420 | v_428;
assign v_432 = v_367 | v_431;
assign v_433 = v_430 | v_432;
assign v_434 = v_418 | v_433;
assign v_436 = v_415 | v_435;
assign v_437 = v_406 | v_408;
assign v_439 = v_436 | v_438;
assign v_440 = v_385 | v_403;
assign v_442 = v_439 | v_441;
assign v_443 = v_392 | v_400;
assign v_445 = v_442 | v_444;
assign v_446 = v_181 | v_397;
assign v_448 = v_445 | v_447;
assign v_449 = v_218 | v_448;
assign v_450 = v_85 | v_449;
assign v_451 = ~v_87 | v_450;
assign v_452 = v_89 | v_451;
assign v_453 = v_91 | v_452;
assign v_460 = v_47 | v_459;
assign v_461 = v_23 | ~v_28;
assign v_462 = v_18 | v_461;
assign v_463 = ~v_13 | v_462;
assign v_464 = ~v_8 | v_463;
assign v_465 = ~v_43 | v_464;
assign v_466 = ~v_45 | v_465;
assign v_467 = ~v_47 | v_466;
assign v_469 = v_45 | v_458;
assign v_471 = v_8 | v_456;
assign v_473 = v_9 | v_472;
assign v_475 = v_457 | v_474;
assign v_476 = ~v_9 | v_475;
assign v_478 = v_13 | v_455;
assign v_480 = v_14 | v_479;
assign v_482 = v_456 | v_481;
assign v_483 = ~v_14 | v_482;
assign v_485 = ~v_18 | v_454;
assign v_487 = v_19 | v_486;
assign v_489 = v_455 | v_488;
assign v_490 = ~v_19 | v_489;
assign v_493 = v_24 | v_492;
assign v_494 = v_224 | v_454;
assign v_495 = ~v_24 | v_494;
assign v_499 = v_497 | v_498;
assign v_502 = v_500 | v_501;
assign v_505 = v_503 | v_504;
assign v_508 = v_506 | v_507;
assign v_509 = v_43 | v_457;
assign v_515 = v_513 | v_514;
assign v_516 = v_468 | v_512;
assign v_517 = v_515 | v_516;
assign v_518 = v_470 | v_511;
assign v_520 = v_459 | v_519;
assign v_522 = v_507 | v_521;
assign v_524 = v_504 | v_523;
assign v_526 = v_501 | v_525;
assign v_528 = v_498 | v_527;
assign v_529 = v_279 | v_528;
assign v_531 = v_526 | v_530;
assign v_533 = v_524 | v_532;
assign v_535 = v_522 | v_534;
assign v_538 = v_458 | v_537;
assign v_539 = v_536 | v_538;
assign v_540 = v_520 | v_539;
assign v_542 = v_517 | v_541;
assign v_543 = v_508 | v_510;
assign v_545 = v_542 | v_544;
assign v_546 = v_477 | v_505;
assign v_548 = v_545 | v_547;
assign v_549 = v_484 | v_502;
assign v_551 = v_548 | v_550;
assign v_552 = v_491 | v_499;
assign v_554 = v_551 | v_553;
assign v_555 = v_313 | v_496;
assign v_557 = v_554 | v_556;
assign v_558 = v_355 | v_557;
assign v_559 = ~v_87 | v_558;
assign v_560 = v_89 | v_559;
assign v_561 = v_91 | v_560;
assign v_564 = v_562 | ~v_563;
assign v_566 = ~v_7 | v_565;
assign v_567 = ~v_45 | v_69;
assign v_572 = v_44 | v_571;
assign v_575 = v_40 | v_574;
assign v_578 = v_37 | v_577;
assign v_581 = v_34 | v_580;
assign v_584 = v_31 | v_583;
assign v_587 = v_30 | v_586;
assign v_594 = v_591 | v_593;
assign v_596 = ~v_98 | v_595;
assign v_597 = v_193 | v_195;
assign v_600 = v_598 | v_599;
assign v_603 = v_193 | v_602;
assign v_606 = v_192 | v_605;
assign v_609 = v_191 | v_608;
assign v_612 = v_186 | v_611;
assign v_615 = v_184 | v_614;
assign v_618 = v_182 | v_617;
assign v_621 = v_180 | v_620;
assign v_627 = v_327 | v_329;
assign v_630 = v_628 | v_629;
assign v_633 = v_327 | v_632;
assign v_636 = v_326 | v_635;
assign v_639 = v_325 | v_638;
assign v_642 = v_320 | v_641;
assign v_645 = v_318 | v_644;
assign v_648 = v_316 | v_647;
assign v_651 = v_314 | v_650;
assign v_654 = v_313 | v_653;
assign v_659 = v_626 | v_658;
assign v_661 = v_596 | v_660;
assign v_663 = v_412 | v_662;
assign v_664 = v_434 | v_663;
assign v_669 = v_410 | v_668;
assign v_672 = v_409 | v_671;
assign v_675 = v_404 | v_674;
assign v_678 = v_401 | v_677;
assign v_681 = v_398 | v_680;
assign v_689 = v_514 | v_688;
assign v_690 = v_540 | v_689;
assign v_695 = v_512 | v_694;
assign v_698 = v_511 | v_697;
assign v_701 = v_506 | v_700;
assign v_704 = v_503 | v_703;
assign v_707 = v_500 | v_706;
assign v_710 = v_497 | v_709;
assign v_716 = v_687 | v_715;
assign v_718 = v_661 | v_717;
assign v_719 = v_7 | v_718;
assign v_725 = ~v_720 | v_724;
assign v_726 = v_595 | ~v_721;
assign v_727 = v_660 | v_726;
assign v_728 = v_717 | v_727;
assign v_729 = v_720 | v_728;
assign v_735 = ~v_730 | v_734;
assign v_736 = v_595 | ~v_731;
assign v_737 = v_660 | v_736;
assign v_738 = v_717 | v_737;
assign v_739 = v_730 | v_738;
assign v_745 = ~v_740 | v_744;
assign v_746 = v_595 | ~v_741;
assign v_747 = v_660 | v_746;
assign v_748 = v_717 | v_747;
assign v_749 = v_740 | v_748;
assign v_755 = ~v_750 | v_754;
assign v_756 = v_595 | ~v_751;
assign v_757 = v_660 | v_756;
assign v_758 = v_717 | v_757;
assign v_759 = v_750 | v_758;
assign v_765 = ~v_760 | v_764;
assign v_766 = v_595 | ~v_761;
assign v_767 = v_660 | v_766;
assign v_768 = v_717 | v_767;
assign v_769 = v_760 | v_768;
assign v_774 = v_772 | v_773;
assign v_777 = v_775 | v_776;
assign v_780 = v_778 | v_779;
assign v_781 = ~v_770 | v_780;
assign v_782 = v_595 | ~v_771;
assign v_783 = v_97 | v_593;
assign v_785 = v_660 | v_784;
assign v_786 = v_362 | v_658;
assign v_788 = v_717 | v_787;
assign v_789 = v_564 | v_715;
assign v_791 = v_770 | v_790;
assign v_794 = v_595 | v_793;
assign v_795 = v_660 | v_794;
assign v_796 = v_717 | v_795;
assign v_797 = ~v_792 | v_796;
assign v_801 = v_792 | v_800;
assign v_803 = v_90 | ~v_96;
assign v_806 = v_91 | v_93;
assign v_808 = v_806 | ~v_807;
assign v_810 = ~v_91 | v_222;
assign v_811 = ~v_91 | v_358;
assign v_813 = ~v_361 | v_812;
assign v_815 = ~v_91 | v_452;
assign v_816 = ~v_91 | v_560;
assign v_818 = ~v_563 | v_817;
assign v_820 = ~v_802 | v_819;
assign v_822 = ~v_804 | v_821;
assign v_825 = v_822 | v_824;
assign v_828 = v_826 | v_827;
assign v_830 = v_825 | v_829;
assign v_833 = v_831 | v_832;
assign v_835 = v_830 | v_834;
assign v_836 = v_802 | v_835;
assign v_843 = ~v_837 | v_842;
assign v_844 = v_821 | ~v_838;
assign v_845 = v_824 | v_844;
assign v_846 = v_829 | v_845;
assign v_847 = v_834 | v_846;
assign v_848 = v_837 | v_847;
assign v_855 = ~v_849 | v_854;
assign v_856 = v_821 | ~v_850;
assign v_857 = v_824 | v_856;
assign v_858 = v_829 | v_857;
assign v_859 = v_834 | v_858;
assign v_860 = v_849 | v_859;
assign v_867 = ~v_861 | v_866;
assign v_868 = v_821 | ~v_862;
assign v_869 = v_824 | v_868;
assign v_870 = v_829 | v_869;
assign v_871 = v_834 | v_870;
assign v_872 = v_861 | v_871;
assign v_879 = ~v_873 | v_878;
assign v_880 = v_821 | ~v_874;
assign v_881 = v_824 | v_880;
assign v_882 = v_829 | v_881;
assign v_883 = v_834 | v_882;
assign v_884 = v_873 | v_883;
assign v_891 = ~v_885 | v_890;
assign v_892 = v_821 | ~v_886;
assign v_893 = v_824 | v_892;
assign v_894 = v_829 | v_893;
assign v_895 = v_834 | v_894;
assign v_896 = v_885 | v_895;
assign v_901 = v_899 | v_900;
assign v_905 = v_903 | v_904;
assign v_908 = v_906 | v_907;
assign v_909 = ~v_897 | v_908;
assign v_910 = v_821 | ~v_898;
assign v_911 = ~v_91 | v_803;
assign v_913 = v_824 | v_912;
assign v_914 = v_829 | v_913;
assign v_915 = v_813 | v_827;
assign v_917 = v_834 | v_916;
assign v_918 = v_818 | v_832;
assign v_920 = v_897 | v_919;
assign v_923 = v_821 | v_922;
assign v_924 = v_824 | v_923;
assign v_925 = v_829 | v_924;
assign v_926 = v_834 | v_925;
assign v_927 = ~v_921 | v_926;
assign v_932 = v_921 | v_931;
assign v_934 = v_86 | v_87;
assign v_935 = v_89 | v_934;
assign v_936 = v_91 | v_935;
assign v_937 = v_90 | ~v_91;
assign v_939 = ~v_96 | v_938;
assign v_942 = v_93 | ~v_807;
assign v_944 = ~v_89 | v_221;
assign v_945 = v_91 | v_944;
assign v_946 = ~v_89 | v_357;
assign v_947 = v_91 | v_946;
assign v_949 = ~v_361 | v_948;
assign v_951 = ~v_89 | v_451;
assign v_952 = v_91 | v_951;
assign v_953 = ~v_89 | v_559;
assign v_954 = v_91 | v_953;
assign v_956 = ~v_563 | v_955;
assign v_958 = ~v_933 | v_957;
assign v_963 = v_961 | v_962;
assign v_965 = ~v_940 | v_964;
assign v_967 = v_965 | v_966;
assign v_972 = v_969 | v_971;
assign v_974 = v_967 | v_973;
assign v_979 = v_976 | v_978;
assign v_981 = v_974 | v_980;
assign v_982 = v_933 | v_981;
assign v_989 = ~v_983 | v_988;
assign v_990 = v_964 | ~v_984;
assign v_991 = v_966 | v_990;
assign v_992 = v_973 | v_991;
assign v_993 = v_980 | v_992;
assign v_994 = v_983 | v_993;
assign v_1001 = ~v_995 | v_1000;
assign v_1002 = v_964 | ~v_996;
assign v_1003 = v_966 | v_1002;
assign v_1004 = v_973 | v_1003;
assign v_1005 = v_980 | v_1004;
assign v_1006 = v_995 | v_1005;
assign v_1013 = ~v_1007 | v_1012;
assign v_1014 = v_964 | ~v_1008;
assign v_1015 = v_966 | v_1014;
assign v_1016 = v_973 | v_1015;
assign v_1017 = v_980 | v_1016;
assign v_1018 = v_1007 | v_1017;
assign v_1025 = ~v_1019 | v_1024;
assign v_1026 = v_964 | ~v_1020;
assign v_1027 = v_966 | v_1026;
assign v_1028 = v_973 | v_1027;
assign v_1029 = v_980 | v_1028;
assign v_1030 = v_1019 | v_1029;
assign v_1037 = ~v_1031 | v_1036;
assign v_1038 = v_964 | ~v_1032;
assign v_1039 = v_966 | v_1038;
assign v_1040 = v_973 | v_1039;
assign v_1041 = v_980 | v_1040;
assign v_1042 = v_1031 | v_1041;
assign v_1047 = v_1045 | v_1046;
assign v_1050 = v_1048 | v_1049;
assign v_1053 = v_1051 | v_1052;
assign v_1056 = v_1054 | v_1055;
assign v_1057 = ~v_1043 | v_1056;
assign v_1058 = v_964 | ~v_1044;
assign v_1059 = v_939 | v_962;
assign v_1061 = v_966 | v_1060;
assign v_1062 = v_91 | v_942;
assign v_1064 = v_973 | v_1063;
assign v_1065 = v_949 | v_971;
assign v_1067 = v_980 | v_1066;
assign v_1068 = v_956 | v_978;
assign v_1070 = v_1043 | v_1069;
assign v_1073 = v_964 | v_1072;
assign v_1074 = v_966 | v_1073;
assign v_1075 = v_973 | v_1074;
assign v_1076 = v_980 | v_1075;
assign v_1077 = ~v_1071 | v_1076;
assign v_1082 = v_1071 | v_1081;
assign v_1084 = ~v_96 | v_935;
assign v_1087 = v_95 | ~v_807;
assign v_1089 = ~v_91 | v_944;
assign v_1090 = ~v_91 | v_946;
assign v_1092 = ~v_361 | v_1091;
assign v_1094 = ~v_91 | v_951;
assign v_1095 = ~v_91 | v_953;
assign v_1097 = ~v_563 | v_1096;
assign v_1099 = ~v_1083 | v_1098;
assign v_1101 = ~v_1085 | v_1100;
assign v_1103 = v_1101 | v_1102;
assign v_1106 = v_1104 | v_1105;
assign v_1108 = v_1103 | v_1107;
assign v_1111 = v_1109 | v_1110;
assign v_1113 = v_1108 | v_1112;
assign v_1114 = v_1083 | v_1113;
assign v_1121 = ~v_1115 | v_1120;
assign v_1122 = v_1100 | ~v_1116;
assign v_1123 = v_1102 | v_1122;
assign v_1124 = v_1107 | v_1123;
assign v_1125 = v_1112 | v_1124;
assign v_1126 = v_1115 | v_1125;
assign v_1133 = ~v_1127 | v_1132;
assign v_1134 = v_1100 | ~v_1128;
assign v_1135 = v_1102 | v_1134;
assign v_1136 = v_1107 | v_1135;
assign v_1137 = v_1112 | v_1136;
assign v_1138 = v_1127 | v_1137;
assign v_1145 = ~v_1139 | v_1144;
assign v_1146 = v_1100 | ~v_1140;
assign v_1147 = v_1102 | v_1146;
assign v_1148 = v_1107 | v_1147;
assign v_1149 = v_1112 | v_1148;
assign v_1150 = v_1139 | v_1149;
assign v_1157 = ~v_1151 | v_1156;
assign v_1158 = v_1100 | ~v_1152;
assign v_1159 = v_1102 | v_1158;
assign v_1160 = v_1107 | v_1159;
assign v_1161 = v_1112 | v_1160;
assign v_1162 = v_1151 | v_1161;
assign v_1169 = ~v_1163 | v_1168;
assign v_1170 = v_1100 | ~v_1164;
assign v_1171 = v_1102 | v_1170;
assign v_1172 = v_1107 | v_1171;
assign v_1173 = v_1112 | v_1172;
assign v_1174 = v_1163 | v_1173;
assign v_1179 = v_1177 | v_1178;
assign v_1182 = v_1180 | v_1181;
assign v_1185 = v_1183 | v_1184;
assign v_1188 = v_1186 | v_1187;
assign v_1189 = ~v_1175 | v_1188;
assign v_1190 = v_1100 | ~v_1176;
assign v_1191 = ~v_91 | v_1084;
assign v_1193 = v_1102 | v_1192;
assign v_1194 = v_591 | v_1087;
assign v_1196 = v_1107 | v_1195;
assign v_1197 = v_1092 | v_1105;
assign v_1199 = v_1112 | v_1198;
assign v_1200 = v_1097 | v_1110;
assign v_1202 = v_1175 | v_1201;
assign v_1205 = v_1100 | v_1204;
assign v_1206 = v_1102 | v_1205;
assign v_1207 = v_1107 | v_1206;
assign v_1208 = v_1112 | v_1207;
assign v_1209 = ~v_1203 | v_1208;
assign v_1214 = v_1203 | v_1213;
assign v_1216 = ~v_89 | v_934;
assign v_1217 = v_91 | v_1216;
assign v_1218 = ~v_91 | v_935;
assign v_1220 = ~v_96 | v_1219;
assign v_1223 = v_90 | ~v_807;
assign v_1225 = v_87 | v_220;
assign v_1226 = v_89 | v_1225;
assign v_1227 = v_91 | v_1226;
assign v_1228 = v_87 | v_356;
assign v_1229 = v_89 | v_1228;
assign v_1230 = v_91 | v_1229;
assign v_1232 = ~v_361 | v_1231;
assign v_1234 = v_87 | v_450;
assign v_1235 = v_89 | v_1234;
assign v_1236 = v_91 | v_1235;
assign v_1237 = v_87 | v_558;
assign v_1238 = v_89 | v_1237;
assign v_1239 = v_91 | v_1238;
assign v_1241 = ~v_563 | v_1240;
assign v_1243 = ~v_1215 | v_1242;
assign v_1247 = v_1245 | v_1246;
assign v_1249 = ~v_1221 | v_1248;
assign v_1251 = v_1249 | v_1250;
assign v_1258 = v_1254 | v_1257;
assign v_1260 = v_1251 | v_1259;
assign v_1267 = v_1263 | v_1266;
assign v_1269 = v_1260 | v_1268;
assign v_1270 = v_1215 | v_1269;
assign v_1277 = ~v_1271 | v_1276;
assign v_1278 = v_1248 | ~v_1272;
assign v_1279 = v_1250 | v_1278;
assign v_1280 = v_1259 | v_1279;
assign v_1281 = v_1268 | v_1280;
assign v_1282 = v_1271 | v_1281;
assign v_1289 = ~v_1283 | v_1288;
assign v_1290 = v_1248 | ~v_1284;
assign v_1291 = v_1250 | v_1290;
assign v_1292 = v_1259 | v_1291;
assign v_1293 = v_1268 | v_1292;
assign v_1294 = v_1283 | v_1293;
assign v_1301 = ~v_1295 | v_1300;
assign v_1302 = v_1248 | ~v_1296;
assign v_1303 = v_1250 | v_1302;
assign v_1304 = v_1259 | v_1303;
assign v_1305 = v_1268 | v_1304;
assign v_1306 = v_1295 | v_1305;
assign v_1313 = ~v_1307 | v_1312;
assign v_1314 = v_1248 | ~v_1308;
assign v_1315 = v_1250 | v_1314;
assign v_1316 = v_1259 | v_1315;
assign v_1317 = v_1268 | v_1316;
assign v_1318 = v_1307 | v_1317;
assign v_1325 = ~v_1319 | v_1324;
assign v_1326 = v_1248 | ~v_1320;
assign v_1327 = v_1250 | v_1326;
assign v_1328 = v_1259 | v_1327;
assign v_1329 = v_1268 | v_1328;
assign v_1330 = v_1319 | v_1329;
assign v_1335 = v_1333 | v_1334;
assign v_1338 = v_1336 | v_1337;
assign v_1341 = v_1339 | v_1340;
assign v_1344 = v_1342 | v_1343;
assign v_1345 = ~v_1331 | v_1344;
assign v_1346 = v_1248 | ~v_1332;
assign v_1347 = v_1220 | v_1246;
assign v_1349 = v_1250 | v_1348;
assign v_1350 = v_91 | v_1223;
assign v_1352 = v_1259 | v_1351;
assign v_1353 = v_1232 | v_1257;
assign v_1355 = v_1268 | v_1354;
assign v_1356 = v_1241 | v_1266;
assign v_1358 = v_1331 | v_1357;
assign v_1361 = v_1248 | v_1360;
assign v_1362 = v_1250 | v_1361;
assign v_1363 = v_1259 | v_1362;
assign v_1364 = v_1268 | v_1363;
assign v_1365 = ~v_1359 | v_1364;
assign v_1370 = v_1359 | v_1369;
assign v_1372 = ~v_96 | v_1216;
assign v_1375 = ~v_807 | v_938;
assign v_1377 = ~v_91 | v_1226;
assign v_1378 = ~v_91 | v_1229;
assign v_1380 = ~v_361 | v_1379;
assign v_1382 = ~v_91 | v_1235;
assign v_1383 = ~v_91 | v_1238;
assign v_1385 = ~v_563 | v_1384;
assign v_1387 = ~v_1371 | v_1386;
assign v_1389 = ~v_1373 | v_1388;
assign v_1391 = v_1389 | v_1390;
assign v_1394 = v_1392 | v_1393;
assign v_1396 = v_1391 | v_1395;
assign v_1399 = v_1397 | v_1398;
assign v_1401 = v_1396 | v_1400;
assign v_1402 = v_1371 | v_1401;
assign v_1409 = ~v_1403 | v_1408;
assign v_1410 = v_1388 | ~v_1404;
assign v_1411 = v_1390 | v_1410;
assign v_1412 = v_1395 | v_1411;
assign v_1413 = v_1400 | v_1412;
assign v_1414 = v_1403 | v_1413;
assign v_1421 = ~v_1415 | v_1420;
assign v_1422 = v_1388 | ~v_1416;
assign v_1423 = v_1390 | v_1422;
assign v_1424 = v_1395 | v_1423;
assign v_1425 = v_1400 | v_1424;
assign v_1426 = v_1415 | v_1425;
assign v_1433 = ~v_1427 | v_1432;
assign v_1434 = v_1388 | ~v_1428;
assign v_1435 = v_1390 | v_1434;
assign v_1436 = v_1395 | v_1435;
assign v_1437 = v_1400 | v_1436;
assign v_1438 = v_1427 | v_1437;
assign v_1445 = ~v_1439 | v_1444;
assign v_1446 = v_1388 | ~v_1440;
assign v_1447 = v_1390 | v_1446;
assign v_1448 = v_1395 | v_1447;
assign v_1449 = v_1400 | v_1448;
assign v_1450 = v_1439 | v_1449;
assign v_1457 = ~v_1451 | v_1456;
assign v_1458 = v_1388 | ~v_1452;
assign v_1459 = v_1390 | v_1458;
assign v_1460 = v_1395 | v_1459;
assign v_1461 = v_1400 | v_1460;
assign v_1462 = v_1451 | v_1461;
assign v_1467 = v_1465 | v_1466;
assign v_1470 = v_1468 | v_1469;
assign v_1473 = v_1471 | v_1472;
assign v_1476 = v_1474 | v_1475;
assign v_1477 = ~v_1463 | v_1476;
assign v_1478 = v_1388 | ~v_1464;
assign v_1479 = ~v_91 | v_1372;
assign v_1481 = v_1390 | v_1480;
assign v_1482 = v_961 | v_1375;
assign v_1484 = v_1395 | v_1483;
assign v_1485 = v_1380 | v_1393;
assign v_1487 = v_1400 | v_1486;
assign v_1488 = v_1385 | v_1398;
assign v_1490 = v_1463 | v_1489;
assign v_1493 = v_1388 | v_1492;
assign v_1494 = v_1390 | v_1493;
assign v_1495 = v_1395 | v_1494;
assign v_1496 = v_1400 | v_1495;
assign v_1497 = ~v_1491 | v_1496;
assign v_1502 = v_1491 | v_1501;
assign v_1504 = v_83 | v_587;
assign v_1505 = ~v_87 | v_1504;
assign v_1506 = v_89 | v_1505;
assign v_1507 = v_91 | v_1506;
assign v_1508 = ~v_91 | v_1216;
assign v_1510 = ~v_96 | v_1509;
assign v_1513 = ~v_807 | v_935;
assign v_1515 = ~v_89 | v_1225;
assign v_1516 = v_91 | v_1515;
assign v_1517 = ~v_89 | v_1228;
assign v_1518 = v_91 | v_1517;
assign v_1520 = ~v_361 | v_1519;
assign v_1522 = ~v_89 | v_1234;
assign v_1523 = v_91 | v_1522;
assign v_1524 = ~v_89 | v_1237;
assign v_1525 = v_91 | v_1524;
assign v_1527 = ~v_563 | v_1526;
assign v_1529 = ~v_1503 | v_1528;
assign v_1535 = v_1533 | v_1534;
assign v_1537 = ~v_1511 | v_1536;
assign v_1539 = v_1537 | v_1538;
assign v_1544 = v_1541 | v_1543;
assign v_1546 = v_1539 | v_1545;
assign v_1551 = v_1548 | v_1550;
assign v_1553 = v_1546 | v_1552;
assign v_1554 = v_1503 | v_1553;
assign v_1561 = ~v_1555 | v_1560;
assign v_1562 = v_1536 | ~v_1556;
assign v_1563 = v_1538 | v_1562;
assign v_1564 = v_1545 | v_1563;
assign v_1565 = v_1552 | v_1564;
assign v_1566 = v_1555 | v_1565;
assign v_1573 = ~v_1567 | v_1572;
assign v_1574 = v_1536 | ~v_1568;
assign v_1575 = v_1538 | v_1574;
assign v_1576 = v_1545 | v_1575;
assign v_1577 = v_1552 | v_1576;
assign v_1578 = v_1567 | v_1577;
assign v_1585 = ~v_1579 | v_1584;
assign v_1586 = v_1536 | ~v_1580;
assign v_1587 = v_1538 | v_1586;
assign v_1588 = v_1545 | v_1587;
assign v_1589 = v_1552 | v_1588;
assign v_1590 = v_1579 | v_1589;
assign v_1597 = ~v_1591 | v_1596;
assign v_1598 = v_1536 | ~v_1592;
assign v_1599 = v_1538 | v_1598;
assign v_1600 = v_1545 | v_1599;
assign v_1601 = v_1552 | v_1600;
assign v_1602 = v_1591 | v_1601;
assign v_1609 = ~v_1603 | v_1608;
assign v_1610 = v_1536 | ~v_1604;
assign v_1611 = v_1538 | v_1610;
assign v_1612 = v_1545 | v_1611;
assign v_1613 = v_1552 | v_1612;
assign v_1614 = v_1603 | v_1613;
assign v_1619 = v_1617 | v_1618;
assign v_1622 = v_1620 | v_1621;
assign v_1625 = v_1623 | v_1624;
assign v_1628 = v_1626 | v_1627;
assign v_1629 = ~v_1615 | v_1628;
assign v_1630 = v_1536 | ~v_1616;
assign v_1631 = v_1510 | v_1534;
assign v_1633 = v_1538 | v_1632;
assign v_1634 = v_91 | v_1513;
assign v_1636 = v_1545 | v_1635;
assign v_1637 = v_1520 | v_1543;
assign v_1639 = v_1552 | v_1638;
assign v_1640 = v_1527 | v_1550;
assign v_1642 = v_1615 | v_1641;
assign v_1645 = v_1536 | v_1644;
assign v_1646 = v_1538 | v_1645;
assign v_1647 = v_1545 | v_1646;
assign v_1648 = v_1552 | v_1647;
assign v_1649 = ~v_1643 | v_1648;
assign v_1654 = v_1643 | v_1653;
assign v_1656 = ~v_96 | v_1506;
assign v_1659 = ~v_807 | v_1219;
assign v_1661 = ~v_91 | v_1515;
assign v_1662 = ~v_91 | v_1517;
assign v_1664 = ~v_361 | v_1663;
assign v_1666 = ~v_91 | v_1522;
assign v_1667 = ~v_91 | v_1524;
assign v_1669 = ~v_563 | v_1668;
assign v_1671 = ~v_1655 | v_1670;
assign v_1673 = ~v_1657 | v_1672;
assign v_1675 = v_1673 | v_1674;
assign v_1678 = v_1676 | v_1677;
assign v_1680 = v_1675 | v_1679;
assign v_1683 = v_1681 | v_1682;
assign v_1685 = v_1680 | v_1684;
assign v_1686 = v_1655 | v_1685;
assign v_1693 = ~v_1687 | v_1692;
assign v_1694 = v_1672 | ~v_1688;
assign v_1695 = v_1674 | v_1694;
assign v_1696 = v_1679 | v_1695;
assign v_1697 = v_1684 | v_1696;
assign v_1698 = v_1687 | v_1697;
assign v_1705 = ~v_1699 | v_1704;
assign v_1706 = v_1672 | ~v_1700;
assign v_1707 = v_1674 | v_1706;
assign v_1708 = v_1679 | v_1707;
assign v_1709 = v_1684 | v_1708;
assign v_1710 = v_1699 | v_1709;
assign v_1717 = ~v_1711 | v_1716;
assign v_1718 = v_1672 | ~v_1712;
assign v_1719 = v_1674 | v_1718;
assign v_1720 = v_1679 | v_1719;
assign v_1721 = v_1684 | v_1720;
assign v_1722 = v_1711 | v_1721;
assign v_1729 = ~v_1723 | v_1728;
assign v_1730 = v_1672 | ~v_1724;
assign v_1731 = v_1674 | v_1730;
assign v_1732 = v_1679 | v_1731;
assign v_1733 = v_1684 | v_1732;
assign v_1734 = v_1723 | v_1733;
assign v_1741 = ~v_1735 | v_1740;
assign v_1742 = v_1672 | ~v_1736;
assign v_1743 = v_1674 | v_1742;
assign v_1744 = v_1679 | v_1743;
assign v_1745 = v_1684 | v_1744;
assign v_1746 = v_1735 | v_1745;
assign v_1751 = v_1749 | v_1750;
assign v_1754 = v_1752 | v_1753;
assign v_1757 = v_1755 | v_1756;
assign v_1760 = v_1758 | v_1759;
assign v_1761 = ~v_1747 | v_1760;
assign v_1762 = v_1672 | ~v_1748;
assign v_1763 = ~v_91 | v_1656;
assign v_1765 = v_1674 | v_1764;
assign v_1766 = v_1245 | v_1659;
assign v_1768 = v_1679 | v_1767;
assign v_1769 = v_1664 | v_1677;
assign v_1771 = v_1684 | v_1770;
assign v_1772 = v_1669 | v_1682;
assign v_1774 = v_1747 | v_1773;
assign v_1777 = v_1672 | v_1776;
assign v_1778 = v_1674 | v_1777;
assign v_1779 = v_1679 | v_1778;
assign v_1780 = v_1684 | v_1779;
assign v_1781 = ~v_1775 | v_1780;
assign v_1786 = v_1775 | v_1785;
assign v_1788 = ~v_89 | v_1505;
assign v_1789 = v_91 | v_1788;
assign v_1790 = ~v_91 | v_1506;
assign v_1792 = ~v_96 | v_1791;
assign v_1795 = ~v_807 | v_1216;
assign v_1797 = v_219 | v_587;
assign v_1798 = ~v_87 | v_1797;
assign v_1799 = v_89 | v_1798;
assign v_1800 = v_91 | v_1799;
assign v_1801 = v_353 | v_654;
assign v_1802 = ~v_87 | v_1801;
assign v_1803 = v_89 | v_1802;
assign v_1804 = v_91 | v_1803;
assign v_1806 = ~v_361 | v_1805;
assign v_1808 = v_449 | v_587;
assign v_1809 = ~v_87 | v_1808;
assign v_1810 = v_89 | v_1809;
assign v_1811 = v_91 | v_1810;
assign v_1812 = v_557 | v_654;
assign v_1813 = ~v_87 | v_1812;
assign v_1814 = v_89 | v_1813;
assign v_1815 = v_91 | v_1814;
assign v_1817 = ~v_563 | v_1816;
assign v_1819 = ~v_1787 | v_1818;
assign v_1823 = v_1821 | v_1822;
assign v_1825 = ~v_1793 | v_1824;
assign v_1827 = v_1825 | v_1826;
assign v_1836 = v_1831 | v_1835;
assign v_1838 = v_1827 | v_1837;
assign v_1847 = v_1842 | v_1846;
assign v_1849 = v_1838 | v_1848;
assign v_1850 = v_1787 | v_1849;
assign v_1857 = ~v_1851 | v_1856;
assign v_1858 = v_1824 | ~v_1852;
assign v_1859 = v_1826 | v_1858;
assign v_1860 = v_1837 | v_1859;
assign v_1861 = v_1848 | v_1860;
assign v_1862 = v_1851 | v_1861;
assign v_1869 = ~v_1863 | v_1868;
assign v_1870 = v_1824 | ~v_1864;
assign v_1871 = v_1826 | v_1870;
assign v_1872 = v_1837 | v_1871;
assign v_1873 = v_1848 | v_1872;
assign v_1874 = v_1863 | v_1873;
assign v_1881 = ~v_1875 | v_1880;
assign v_1882 = v_1824 | ~v_1876;
assign v_1883 = v_1826 | v_1882;
assign v_1884 = v_1837 | v_1883;
assign v_1885 = v_1848 | v_1884;
assign v_1886 = v_1875 | v_1885;
assign v_1893 = ~v_1887 | v_1892;
assign v_1894 = v_1824 | ~v_1888;
assign v_1895 = v_1826 | v_1894;
assign v_1896 = v_1837 | v_1895;
assign v_1897 = v_1848 | v_1896;
assign v_1898 = v_1887 | v_1897;
assign v_1905 = ~v_1899 | v_1904;
assign v_1906 = v_1824 | ~v_1900;
assign v_1907 = v_1826 | v_1906;
assign v_1908 = v_1837 | v_1907;
assign v_1909 = v_1848 | v_1908;
assign v_1910 = v_1899 | v_1909;
assign v_1915 = v_1913 | v_1914;
assign v_1918 = v_1916 | v_1917;
assign v_1921 = v_1919 | v_1920;
assign v_1924 = v_1922 | v_1923;
assign v_1925 = ~v_1911 | v_1924;
assign v_1926 = v_1824 | ~v_1912;
assign v_1927 = v_1792 | v_1822;
assign v_1929 = v_1826 | v_1928;
assign v_1930 = v_91 | v_1795;
assign v_1932 = v_1837 | v_1931;
assign v_1933 = v_1806 | v_1835;
assign v_1935 = v_1848 | v_1934;
assign v_1936 = v_1817 | v_1846;
assign v_1938 = v_1911 | v_1937;
assign v_1941 = v_1824 | v_1940;
assign v_1942 = v_1826 | v_1941;
assign v_1943 = v_1837 | v_1942;
assign v_1944 = v_1848 | v_1943;
assign v_1945 = ~v_1939 | v_1944;
assign v_1950 = v_1939 | v_1949;
assign v_1952 = ~v_96 | v_1788;
assign v_1955 = ~v_807 | v_1509;
assign v_1957 = ~v_91 | v_1799;
assign v_1958 = ~v_91 | v_1803;
assign v_1960 = ~v_361 | v_1959;
assign v_1962 = ~v_91 | v_1810;
assign v_1963 = ~v_91 | v_1814;
assign v_1965 = ~v_563 | v_1964;
assign v_1967 = ~v_1951 | v_1966;
assign v_1969 = ~v_1953 | v_1968;
assign v_1971 = v_1969 | v_1970;
assign v_1974 = v_1972 | v_1973;
assign v_1976 = v_1971 | v_1975;
assign v_1979 = v_1977 | v_1978;
assign v_1981 = v_1976 | v_1980;
assign v_1982 = v_1951 | v_1981;
assign v_1989 = ~v_1983 | v_1988;
assign v_1990 = v_1968 | ~v_1984;
assign v_1991 = v_1970 | v_1990;
assign v_1992 = v_1975 | v_1991;
assign v_1993 = v_1980 | v_1992;
assign v_1994 = v_1983 | v_1993;
assign v_2001 = ~v_1995 | v_2000;
assign v_2002 = v_1968 | ~v_1996;
assign v_2003 = v_1970 | v_2002;
assign v_2004 = v_1975 | v_2003;
assign v_2005 = v_1980 | v_2004;
assign v_2006 = v_1995 | v_2005;
assign v_2013 = ~v_2007 | v_2012;
assign v_2014 = v_1968 | ~v_2008;
assign v_2015 = v_1970 | v_2014;
assign v_2016 = v_1975 | v_2015;
assign v_2017 = v_1980 | v_2016;
assign v_2018 = v_2007 | v_2017;
assign v_2025 = ~v_2019 | v_2024;
assign v_2026 = v_1968 | ~v_2020;
assign v_2027 = v_1970 | v_2026;
assign v_2028 = v_1975 | v_2027;
assign v_2029 = v_1980 | v_2028;
assign v_2030 = v_2019 | v_2029;
assign v_2037 = ~v_2031 | v_2036;
assign v_2038 = v_1968 | ~v_2032;
assign v_2039 = v_1970 | v_2038;
assign v_2040 = v_1975 | v_2039;
assign v_2041 = v_1980 | v_2040;
assign v_2042 = v_2031 | v_2041;
assign v_2047 = v_2045 | v_2046;
assign v_2050 = v_2048 | v_2049;
assign v_2053 = v_2051 | v_2052;
assign v_2056 = v_2054 | v_2055;
assign v_2057 = ~v_2043 | v_2056;
assign v_2058 = v_1968 | ~v_2044;
assign v_2059 = ~v_91 | v_1952;
assign v_2061 = v_1970 | v_2060;
assign v_2062 = v_1533 | v_1955;
assign v_2064 = v_1975 | v_2063;
assign v_2065 = v_1960 | v_1973;
assign v_2067 = v_1980 | v_2066;
assign v_2068 = v_1965 | v_1978;
assign v_2070 = v_2043 | v_2069;
assign v_2077 = ~v_2071 | v_2076;
assign v_2078 = v_1968 | ~v_2072;
assign v_2079 = v_1970 | v_2078;
assign v_2080 = v_1975 | v_2079;
assign v_2081 = v_1980 | v_2080;
assign v_2082 = v_2071 | v_2081;
assign v_2084 = v_87 | v_1504;
assign v_2085 = v_89 | v_2084;
assign v_2086 = v_91 | v_2085;
assign v_2087 = ~v_91 | v_1788;
assign v_2089 = ~v_96 | v_2088;
assign v_2092 = ~v_807 | v_1506;
assign v_2094 = ~v_89 | v_1798;
assign v_2095 = v_91 | v_2094;
assign v_2096 = ~v_89 | v_1802;
assign v_2097 = v_91 | v_2096;
assign v_2099 = ~v_361 | v_2098;
assign v_2101 = ~v_89 | v_1809;
assign v_2102 = v_91 | v_2101;
assign v_2103 = ~v_89 | v_1813;
assign v_2104 = v_91 | v_2103;
assign v_2106 = ~v_563 | v_2105;
assign v_2108 = ~v_2083 | v_2107;
assign v_2113 = v_2111 | v_2112;
assign v_2115 = ~v_2090 | v_2114;
assign v_2117 = v_2115 | v_2116;
assign v_2122 = v_2119 | v_2121;
assign v_2124 = v_2117 | v_2123;
assign v_2129 = v_2126 | v_2128;
assign v_2131 = v_2124 | v_2130;
assign v_2132 = v_2083 | v_2131;
assign v_2139 = ~v_2133 | v_2138;
assign v_2140 = v_2114 | ~v_2134;
assign v_2141 = v_2116 | v_2140;
assign v_2142 = v_2123 | v_2141;
assign v_2143 = v_2130 | v_2142;
assign v_2144 = v_2133 | v_2143;
assign v_2151 = ~v_2145 | v_2150;
assign v_2152 = v_2114 | ~v_2146;
assign v_2153 = v_2116 | v_2152;
assign v_2154 = v_2123 | v_2153;
assign v_2155 = v_2130 | v_2154;
assign v_2156 = v_2145 | v_2155;
assign v_2163 = ~v_2157 | v_2162;
assign v_2164 = v_2114 | ~v_2158;
assign v_2165 = v_2116 | v_2164;
assign v_2166 = v_2123 | v_2165;
assign v_2167 = v_2130 | v_2166;
assign v_2168 = v_2157 | v_2167;
assign v_2175 = ~v_2169 | v_2174;
assign v_2176 = v_2114 | ~v_2170;
assign v_2177 = v_2116 | v_2176;
assign v_2178 = v_2123 | v_2177;
assign v_2179 = v_2130 | v_2178;
assign v_2180 = v_2169 | v_2179;
assign v_2187 = ~v_2181 | v_2186;
assign v_2188 = v_2114 | ~v_2182;
assign v_2189 = v_2116 | v_2188;
assign v_2190 = v_2123 | v_2189;
assign v_2191 = v_2130 | v_2190;
assign v_2192 = v_2181 | v_2191;
assign v_2197 = v_2195 | v_2196;
assign v_2200 = v_2198 | v_2199;
assign v_2203 = v_2201 | v_2202;
assign v_2206 = v_2204 | v_2205;
assign v_2207 = ~v_2193 | v_2206;
assign v_2208 = v_2114 | ~v_2194;
assign v_2209 = v_2089 | v_2112;
assign v_2211 = v_2116 | v_2210;
assign v_2212 = v_91 | v_2092;
assign v_2214 = v_2123 | v_2213;
assign v_2215 = v_2099 | v_2121;
assign v_2217 = v_2130 | v_2216;
assign v_2218 = v_2106 | v_2128;
assign v_2220 = v_2193 | v_2219;
assign v_2227 = ~v_2221 | v_2226;
assign v_2228 = v_2114 | ~v_2222;
assign v_2229 = v_2116 | v_2228;
assign v_2230 = v_2123 | v_2229;
assign v_2231 = v_2130 | v_2230;
assign v_2232 = v_2221 | v_2231;
assign v_2234 = ~v_96 | v_2085;
assign v_2237 = ~v_807 | v_1791;
assign v_2239 = ~v_91 | v_2094;
assign v_2240 = ~v_91 | v_2096;
assign v_2242 = ~v_361 | v_2241;
assign v_2244 = ~v_91 | v_2101;
assign v_2245 = ~v_91 | v_2103;
assign v_2247 = ~v_563 | v_2246;
assign v_2249 = ~v_2233 | v_2248;
assign v_2251 = ~v_2235 | v_2250;
assign v_2253 = v_2251 | v_2252;
assign v_2256 = v_2254 | v_2255;
assign v_2258 = v_2253 | v_2257;
assign v_2261 = v_2259 | v_2260;
assign v_2263 = v_2258 | v_2262;
assign v_2264 = v_2233 | v_2263;
assign v_2271 = ~v_2265 | v_2270;
assign v_2272 = v_2250 | ~v_2266;
assign v_2273 = v_2252 | v_2272;
assign v_2274 = v_2257 | v_2273;
assign v_2275 = v_2262 | v_2274;
assign v_2276 = v_2265 | v_2275;
assign v_2283 = ~v_2277 | v_2282;
assign v_2284 = v_2250 | ~v_2278;
assign v_2285 = v_2252 | v_2284;
assign v_2286 = v_2257 | v_2285;
assign v_2287 = v_2262 | v_2286;
assign v_2288 = v_2277 | v_2287;
assign v_2295 = ~v_2289 | v_2294;
assign v_2296 = v_2250 | ~v_2290;
assign v_2297 = v_2252 | v_2296;
assign v_2298 = v_2257 | v_2297;
assign v_2299 = v_2262 | v_2298;
assign v_2300 = v_2289 | v_2299;
assign v_2307 = ~v_2301 | v_2306;
assign v_2308 = v_2250 | ~v_2302;
assign v_2309 = v_2252 | v_2308;
assign v_2310 = v_2257 | v_2309;
assign v_2311 = v_2262 | v_2310;
assign v_2312 = v_2301 | v_2311;
assign v_2319 = ~v_2313 | v_2318;
assign v_2320 = v_2250 | ~v_2314;
assign v_2321 = v_2252 | v_2320;
assign v_2322 = v_2257 | v_2321;
assign v_2323 = v_2262 | v_2322;
assign v_2324 = v_2313 | v_2323;
assign v_2329 = v_2327 | v_2328;
assign v_2332 = v_2330 | v_2331;
assign v_2335 = v_2333 | v_2334;
assign v_2338 = v_2336 | v_2337;
assign v_2339 = ~v_2325 | v_2338;
assign v_2340 = v_2250 | ~v_2326;
assign v_2341 = ~v_91 | v_2234;
assign v_2343 = v_2252 | v_2342;
assign v_2344 = v_1821 | v_2237;
assign v_2346 = v_2257 | v_2345;
assign v_2347 = v_2242 | v_2255;
assign v_2349 = v_2262 | v_2348;
assign v_2350 = v_2247 | v_2260;
assign v_2352 = v_2325 | v_2351;
assign v_2359 = ~v_2353 | v_2358;
assign v_2360 = v_2250 | ~v_2354;
assign v_2361 = v_2252 | v_2360;
assign v_2362 = v_2257 | v_2361;
assign v_2363 = v_2262 | v_2362;
assign v_2364 = v_2353 | v_2363;
assign v_2366 = ~v_89 | v_2084;
assign v_2367 = v_91 | v_2366;
assign v_2368 = ~v_91 | v_2085;
assign v_2370 = ~v_96 | v_2369;
assign v_2373 = ~v_807 | v_1788;
assign v_2375 = v_87 | v_1797;
assign v_2376 = v_89 | v_2375;
assign v_2377 = v_91 | v_2376;
assign v_2378 = v_87 | v_1801;
assign v_2379 = v_89 | v_2378;
assign v_2380 = v_91 | v_2379;
assign v_2382 = ~v_361 | v_2381;
assign v_2384 = v_87 | v_1808;
assign v_2385 = v_89 | v_2384;
assign v_2386 = v_91 | v_2385;
assign v_2387 = v_87 | v_1812;
assign v_2388 = v_89 | v_2387;
assign v_2389 = v_91 | v_2388;
assign v_2391 = ~v_563 | v_2390;
assign v_2393 = ~v_2365 | v_2392;
assign v_2397 = v_2395 | v_2396;
assign v_2399 = ~v_2371 | v_2398;
assign v_2401 = v_2399 | v_2400;
assign v_2408 = v_2404 | v_2407;
assign v_2410 = v_2401 | v_2409;
assign v_2417 = v_2413 | v_2416;
assign v_2419 = v_2410 | v_2418;
assign v_2420 = v_2365 | v_2419;
assign v_2427 = ~v_2421 | v_2426;
assign v_2428 = v_2398 | ~v_2422;
assign v_2429 = v_2400 | v_2428;
assign v_2430 = v_2409 | v_2429;
assign v_2431 = v_2418 | v_2430;
assign v_2432 = v_2421 | v_2431;
assign v_2439 = ~v_2433 | v_2438;
assign v_2440 = v_2398 | ~v_2434;
assign v_2441 = v_2400 | v_2440;
assign v_2442 = v_2409 | v_2441;
assign v_2443 = v_2418 | v_2442;
assign v_2444 = v_2433 | v_2443;
assign v_2451 = ~v_2445 | v_2450;
assign v_2452 = v_2398 | ~v_2446;
assign v_2453 = v_2400 | v_2452;
assign v_2454 = v_2409 | v_2453;
assign v_2455 = v_2418 | v_2454;
assign v_2456 = v_2445 | v_2455;
assign v_2463 = ~v_2457 | v_2462;
assign v_2464 = v_2398 | ~v_2458;
assign v_2465 = v_2400 | v_2464;
assign v_2466 = v_2409 | v_2465;
assign v_2467 = v_2418 | v_2466;
assign v_2468 = v_2457 | v_2467;
assign v_2475 = ~v_2469 | v_2474;
assign v_2476 = v_2398 | ~v_2470;
assign v_2477 = v_2400 | v_2476;
assign v_2478 = v_2409 | v_2477;
assign v_2479 = v_2418 | v_2478;
assign v_2480 = v_2469 | v_2479;
assign v_2485 = v_2483 | v_2484;
assign v_2488 = v_2486 | v_2487;
assign v_2491 = v_2489 | v_2490;
assign v_2494 = v_2492 | v_2493;
assign v_2495 = ~v_2481 | v_2494;
assign v_2496 = v_2398 | ~v_2482;
assign v_2497 = v_2370 | v_2396;
assign v_2499 = v_2400 | v_2498;
assign v_2500 = v_91 | v_2373;
assign v_2502 = v_2409 | v_2501;
assign v_2503 = v_2382 | v_2407;
assign v_2505 = v_2418 | v_2504;
assign v_2506 = v_2391 | v_2416;
assign v_2508 = v_2481 | v_2507;
assign v_2511 = v_2398 | v_2510;
assign v_2512 = v_2400 | v_2511;
assign v_2513 = v_2409 | v_2512;
assign v_2514 = v_2418 | v_2513;
assign v_2515 = ~v_2509 | v_2514;
assign v_2520 = v_2509 | v_2519;
assign v_2522 = ~v_96 | v_2366;
assign v_2525 = ~v_807 | v_2088;
assign v_2527 = ~v_91 | v_2376;
assign v_2528 = ~v_91 | v_2379;
assign v_2530 = ~v_361 | v_2529;
assign v_2532 = ~v_91 | v_2385;
assign v_2533 = ~v_91 | v_2388;
assign v_2535 = ~v_563 | v_2534;
assign v_2537 = ~v_2521 | v_2536;
assign v_2539 = ~v_2523 | v_2538;
assign v_2541 = v_2539 | v_2540;
assign v_2544 = v_2542 | v_2543;
assign v_2546 = v_2541 | v_2545;
assign v_2549 = v_2547 | v_2548;
assign v_2551 = v_2546 | v_2550;
assign v_2552 = v_2521 | v_2551;
assign v_2559 = ~v_2553 | v_2558;
assign v_2560 = v_2538 | ~v_2554;
assign v_2561 = v_2540 | v_2560;
assign v_2562 = v_2545 | v_2561;
assign v_2563 = v_2550 | v_2562;
assign v_2564 = v_2553 | v_2563;
assign v_2571 = ~v_2565 | v_2570;
assign v_2572 = v_2538 | ~v_2566;
assign v_2573 = v_2540 | v_2572;
assign v_2574 = v_2545 | v_2573;
assign v_2575 = v_2550 | v_2574;
assign v_2576 = v_2565 | v_2575;
assign v_2583 = ~v_2577 | v_2582;
assign v_2584 = v_2538 | ~v_2578;
assign v_2585 = v_2540 | v_2584;
assign v_2586 = v_2545 | v_2585;
assign v_2587 = v_2550 | v_2586;
assign v_2588 = v_2577 | v_2587;
assign v_2595 = ~v_2589 | v_2594;
assign v_2596 = v_2538 | ~v_2590;
assign v_2597 = v_2540 | v_2596;
assign v_2598 = v_2545 | v_2597;
assign v_2599 = v_2550 | v_2598;
assign v_2600 = v_2589 | v_2599;
assign v_2607 = ~v_2601 | v_2606;
assign v_2608 = v_2538 | ~v_2602;
assign v_2609 = v_2540 | v_2608;
assign v_2610 = v_2545 | v_2609;
assign v_2611 = v_2550 | v_2610;
assign v_2612 = v_2601 | v_2611;
assign v_2617 = v_2615 | v_2616;
assign v_2620 = v_2618 | v_2619;
assign v_2623 = v_2621 | v_2622;
assign v_2626 = v_2624 | v_2625;
assign v_2627 = ~v_2613 | v_2626;
assign v_2628 = v_2538 | ~v_2614;
assign v_2629 = ~v_91 | v_2522;
assign v_2631 = v_2540 | v_2630;
assign v_2632 = v_2111 | v_2525;
assign v_2634 = v_2545 | v_2633;
assign v_2635 = v_2530 | v_2543;
assign v_2637 = v_2550 | v_2636;
assign v_2638 = v_2535 | v_2548;
assign v_2640 = v_2613 | v_2639;
assign v_2643 = v_2538 | v_2642;
assign v_2644 = v_2540 | v_2643;
assign v_2645 = v_2545 | v_2644;
assign v_2646 = v_2550 | v_2645;
assign v_2647 = ~v_2641 | v_2646;
assign v_2652 = v_2641 | v_2651;
assign v_2654 = v_80 | v_584;
assign v_2655 = v_85 | v_2654;
assign v_2656 = ~v_87 | v_2655;
assign v_2657 = v_89 | v_2656;
assign v_2658 = v_91 | v_2657;
assign v_2659 = ~v_91 | v_2366;
assign v_2661 = ~v_96 | v_2660;
assign v_2664 = ~v_807 | v_2085;
assign v_2666 = ~v_89 | v_2375;
assign v_2667 = v_91 | v_2666;
assign v_2668 = ~v_89 | v_2378;
assign v_2669 = v_91 | v_2668;
assign v_2671 = ~v_361 | v_2670;
assign v_2673 = ~v_89 | v_2384;
assign v_2674 = v_91 | v_2673;
assign v_2675 = ~v_89 | v_2387;
assign v_2676 = v_91 | v_2675;
assign v_2678 = ~v_563 | v_2677;
assign v_2680 = ~v_2653 | v_2679;
assign v_2687 = v_2685 | v_2686;
assign v_2689 = ~v_2662 | v_2688;
assign v_2691 = v_2689 | v_2690;
assign v_2696 = v_2693 | v_2695;
assign v_2698 = v_2691 | v_2697;
assign v_2703 = v_2700 | v_2702;
assign v_2705 = v_2698 | v_2704;
assign v_2706 = v_2653 | v_2705;
assign v_2713 = ~v_2707 | v_2712;
assign v_2714 = v_2688 | ~v_2708;
assign v_2715 = v_2690 | v_2714;
assign v_2716 = v_2697 | v_2715;
assign v_2717 = v_2704 | v_2716;
assign v_2718 = v_2707 | v_2717;
assign v_2725 = ~v_2719 | v_2724;
assign v_2726 = v_2688 | ~v_2720;
assign v_2727 = v_2690 | v_2726;
assign v_2728 = v_2697 | v_2727;
assign v_2729 = v_2704 | v_2728;
assign v_2730 = v_2719 | v_2729;
assign v_2737 = ~v_2731 | v_2736;
assign v_2738 = v_2688 | ~v_2732;
assign v_2739 = v_2690 | v_2738;
assign v_2740 = v_2697 | v_2739;
assign v_2741 = v_2704 | v_2740;
assign v_2742 = v_2731 | v_2741;
assign v_2749 = ~v_2743 | v_2748;
assign v_2750 = v_2688 | ~v_2744;
assign v_2751 = v_2690 | v_2750;
assign v_2752 = v_2697 | v_2751;
assign v_2753 = v_2704 | v_2752;
assign v_2754 = v_2743 | v_2753;
assign v_2761 = ~v_2755 | v_2760;
assign v_2762 = v_2688 | ~v_2756;
assign v_2763 = v_2690 | v_2762;
assign v_2764 = v_2697 | v_2763;
assign v_2765 = v_2704 | v_2764;
assign v_2766 = v_2755 | v_2765;
assign v_2771 = v_2769 | v_2770;
assign v_2774 = v_2772 | v_2773;
assign v_2777 = v_2775 | v_2776;
assign v_2780 = v_2778 | v_2779;
assign v_2781 = ~v_2767 | v_2780;
assign v_2782 = v_2688 | ~v_2768;
assign v_2783 = v_2661 | v_2686;
assign v_2785 = v_2690 | v_2784;
assign v_2786 = v_91 | v_2664;
assign v_2788 = v_2697 | v_2787;
assign v_2789 = v_2671 | v_2695;
assign v_2791 = v_2704 | v_2790;
assign v_2792 = v_2678 | v_2702;
assign v_2794 = v_2767 | v_2793;
assign v_2797 = v_2688 | v_2796;
assign v_2798 = v_2690 | v_2797;
assign v_2799 = v_2697 | v_2798;
assign v_2800 = v_2704 | v_2799;
assign v_2801 = ~v_2795 | v_2800;
assign v_2806 = v_2795 | v_2805;
assign v_2808 = ~v_96 | v_2657;
assign v_2811 = ~v_807 | v_2369;
assign v_2813 = ~v_91 | v_2666;
assign v_2814 = ~v_91 | v_2668;
assign v_2816 = ~v_361 | v_2815;
assign v_2818 = ~v_91 | v_2673;
assign v_2819 = ~v_91 | v_2675;
assign v_2821 = ~v_563 | v_2820;
assign v_2823 = ~v_2807 | v_2822;
assign v_2825 = ~v_2809 | v_2824;
assign v_2827 = v_2825 | v_2826;
assign v_2830 = v_2828 | v_2829;
assign v_2832 = v_2827 | v_2831;
assign v_2835 = v_2833 | v_2834;
assign v_2837 = v_2832 | v_2836;
assign v_2838 = v_2807 | v_2837;
assign v_2845 = ~v_2839 | v_2844;
assign v_2846 = v_2824 | ~v_2840;
assign v_2847 = v_2826 | v_2846;
assign v_2848 = v_2831 | v_2847;
assign v_2849 = v_2836 | v_2848;
assign v_2850 = v_2839 | v_2849;
assign v_2857 = ~v_2851 | v_2856;
assign v_2858 = v_2824 | ~v_2852;
assign v_2859 = v_2826 | v_2858;
assign v_2860 = v_2831 | v_2859;
assign v_2861 = v_2836 | v_2860;
assign v_2862 = v_2851 | v_2861;
assign v_2869 = ~v_2863 | v_2868;
assign v_2870 = v_2824 | ~v_2864;
assign v_2871 = v_2826 | v_2870;
assign v_2872 = v_2831 | v_2871;
assign v_2873 = v_2836 | v_2872;
assign v_2874 = v_2863 | v_2873;
assign v_2881 = ~v_2875 | v_2880;
assign v_2882 = v_2824 | ~v_2876;
assign v_2883 = v_2826 | v_2882;
assign v_2884 = v_2831 | v_2883;
assign v_2885 = v_2836 | v_2884;
assign v_2886 = v_2875 | v_2885;
assign v_2893 = ~v_2887 | v_2892;
assign v_2894 = v_2824 | ~v_2888;
assign v_2895 = v_2826 | v_2894;
assign v_2896 = v_2831 | v_2895;
assign v_2897 = v_2836 | v_2896;
assign v_2898 = v_2887 | v_2897;
assign v_2903 = v_2901 | v_2902;
assign v_2906 = v_2904 | v_2905;
assign v_2909 = v_2907 | v_2908;
assign v_2912 = v_2910 | v_2911;
assign v_2913 = ~v_2899 | v_2912;
assign v_2914 = v_2824 | ~v_2900;
assign v_2915 = ~v_91 | v_2808;
assign v_2917 = v_2826 | v_2916;
assign v_2918 = v_2395 | v_2811;
assign v_2920 = v_2831 | v_2919;
assign v_2921 = v_2816 | v_2829;
assign v_2923 = v_2836 | v_2922;
assign v_2924 = v_2821 | v_2834;
assign v_2926 = v_2899 | v_2925;
assign v_2929 = v_2824 | v_2928;
assign v_2930 = v_2826 | v_2929;
assign v_2931 = v_2831 | v_2930;
assign v_2932 = v_2836 | v_2931;
assign v_2933 = ~v_2927 | v_2932;
assign v_2938 = v_2927 | v_2937;
assign v_2940 = ~v_89 | v_2656;
assign v_2941 = v_91 | v_2940;
assign v_2942 = ~v_91 | v_2657;
assign v_2944 = ~v_96 | v_2943;
assign v_2947 = ~v_807 | v_2366;
assign v_2949 = v_216 | v_621;
assign v_2950 = v_85 | v_2949;
assign v_2951 = ~v_87 | v_2950;
assign v_2952 = v_89 | v_2951;
assign v_2953 = v_91 | v_2952;
assign v_2954 = v_350 | v_651;
assign v_2955 = v_355 | v_2954;
assign v_2956 = ~v_87 | v_2955;
assign v_2957 = v_89 | v_2956;
assign v_2958 = v_91 | v_2957;
assign v_2960 = ~v_361 | v_2959;
assign v_2962 = v_448 | v_621;
assign v_2963 = v_85 | v_2962;
assign v_2964 = ~v_87 | v_2963;
assign v_2965 = v_89 | v_2964;
assign v_2966 = v_91 | v_2965;
assign v_2967 = v_554 | v_710;
assign v_2968 = v_355 | v_2967;
assign v_2969 = ~v_87 | v_2968;
assign v_2970 = v_89 | v_2969;
assign v_2971 = v_91 | v_2970;
assign v_2973 = ~v_563 | v_2972;
assign v_2975 = ~v_2939 | v_2974;
assign v_2979 = v_2977 | v_2978;
assign v_2981 = ~v_2945 | v_2980;
assign v_2983 = v_2981 | v_2982;
assign v_2994 = v_2988 | v_2993;
assign v_2996 = v_2983 | v_2995;
assign v_3007 = v_3001 | v_3006;
assign v_3009 = v_2996 | v_3008;
assign v_3010 = v_2939 | v_3009;
assign v_3017 = ~v_3011 | v_3016;
assign v_3018 = v_2980 | ~v_3012;
assign v_3019 = v_2982 | v_3018;
assign v_3020 = v_2995 | v_3019;
assign v_3021 = v_3008 | v_3020;
assign v_3022 = v_3011 | v_3021;
assign v_3029 = ~v_3023 | v_3028;
assign v_3030 = v_2980 | ~v_3024;
assign v_3031 = v_2982 | v_3030;
assign v_3032 = v_2995 | v_3031;
assign v_3033 = v_3008 | v_3032;
assign v_3034 = v_3023 | v_3033;
assign v_3041 = ~v_3035 | v_3040;
assign v_3042 = v_2980 | ~v_3036;
assign v_3043 = v_2982 | v_3042;
assign v_3044 = v_2995 | v_3043;
assign v_3045 = v_3008 | v_3044;
assign v_3046 = v_3035 | v_3045;
assign v_3053 = ~v_3047 | v_3052;
assign v_3054 = v_2980 | ~v_3048;
assign v_3055 = v_2982 | v_3054;
assign v_3056 = v_2995 | v_3055;
assign v_3057 = v_3008 | v_3056;
assign v_3058 = v_3047 | v_3057;
assign v_3065 = ~v_3059 | v_3064;
assign v_3066 = v_2980 | ~v_3060;
assign v_3067 = v_2982 | v_3066;
assign v_3068 = v_2995 | v_3067;
assign v_3069 = v_3008 | v_3068;
assign v_3070 = v_3059 | v_3069;
assign v_3075 = v_3073 | v_3074;
assign v_3078 = v_3076 | v_3077;
assign v_3081 = v_3079 | v_3080;
assign v_3084 = v_3082 | v_3083;
assign v_3085 = ~v_3071 | v_3084;
assign v_3086 = v_2980 | ~v_3072;
assign v_3087 = v_2944 | v_2978;
assign v_3089 = v_2982 | v_3088;
assign v_3090 = v_91 | v_2947;
assign v_3092 = v_2995 | v_3091;
assign v_3093 = v_2960 | v_2993;
assign v_3095 = v_3008 | v_3094;
assign v_3096 = v_2973 | v_3006;
assign v_3098 = v_3071 | v_3097;
assign v_3101 = v_2980 | v_3100;
assign v_3102 = v_2982 | v_3101;
assign v_3103 = v_2995 | v_3102;
assign v_3104 = v_3008 | v_3103;
assign v_3105 = ~v_3099 | v_3104;
assign v_3110 = v_3099 | v_3109;
assign v_3112 = ~v_96 | v_2940;
assign v_3115 = ~v_807 | v_2660;
assign v_3117 = ~v_91 | v_2952;
assign v_3118 = ~v_91 | v_2957;
assign v_3120 = ~v_361 | v_3119;
assign v_3122 = ~v_91 | v_2965;
assign v_3123 = ~v_91 | v_2970;
assign v_3125 = ~v_563 | v_3124;
assign v_3127 = ~v_3111 | v_3126;
assign v_3129 = ~v_3113 | v_3128;
assign v_3131 = v_3129 | v_3130;
assign v_3134 = v_3132 | v_3133;
assign v_3136 = v_3131 | v_3135;
assign v_3139 = v_3137 | v_3138;
assign v_3141 = v_3136 | v_3140;
assign v_3142 = v_3111 | v_3141;
assign v_3149 = ~v_3143 | v_3148;
assign v_3150 = v_3128 | ~v_3144;
assign v_3151 = v_3130 | v_3150;
assign v_3152 = v_3135 | v_3151;
assign v_3153 = v_3140 | v_3152;
assign v_3154 = v_3143 | v_3153;
assign v_3161 = ~v_3155 | v_3160;
assign v_3162 = v_3128 | ~v_3156;
assign v_3163 = v_3130 | v_3162;
assign v_3164 = v_3135 | v_3163;
assign v_3165 = v_3140 | v_3164;
assign v_3166 = v_3155 | v_3165;
assign v_3173 = ~v_3167 | v_3172;
assign v_3174 = v_3128 | ~v_3168;
assign v_3175 = v_3130 | v_3174;
assign v_3176 = v_3135 | v_3175;
assign v_3177 = v_3140 | v_3176;
assign v_3178 = v_3167 | v_3177;
assign v_3185 = ~v_3179 | v_3184;
assign v_3186 = v_3128 | ~v_3180;
assign v_3187 = v_3130 | v_3186;
assign v_3188 = v_3135 | v_3187;
assign v_3189 = v_3140 | v_3188;
assign v_3190 = v_3179 | v_3189;
assign v_3197 = ~v_3191 | v_3196;
assign v_3198 = v_3128 | ~v_3192;
assign v_3199 = v_3130 | v_3198;
assign v_3200 = v_3135 | v_3199;
assign v_3201 = v_3140 | v_3200;
assign v_3202 = v_3191 | v_3201;
assign v_3205 = v_3128 | v_3204;
assign v_3206 = ~v_91 | v_3112;
assign v_3208 = v_3130 | v_3207;
assign v_3209 = v_2685 | v_3115;
assign v_3211 = v_3135 | v_3210;
assign v_3212 = v_3120 | v_3133;
assign v_3214 = v_3140 | v_3213;
assign v_3215 = v_3125 | v_3138;
assign v_3217 = ~v_3203 | v_3216;
assign v_3220 = v_3218 | v_3219;
assign v_3223 = v_3221 | v_3222;
assign v_3226 = v_3224 | v_3225;
assign v_3229 = v_3227 | v_3228;
assign v_3230 = v_3203 | v_3229;
assign v_3237 = ~v_3231 | v_3236;
assign v_3238 = v_3128 | ~v_3232;
assign v_3239 = v_3130 | v_3238;
assign v_3240 = v_3135 | v_3239;
assign v_3241 = v_3140 | v_3240;
assign v_3242 = v_3231 | v_3241;
assign v_3244 = v_87 | v_2655;
assign v_3245 = v_89 | v_3244;
assign v_3246 = v_91 | v_3245;
assign v_3247 = ~v_91 | v_2940;
assign v_3249 = ~v_96 | v_3248;
assign v_3252 = ~v_807 | v_2657;
assign v_3254 = ~v_89 | v_2951;
assign v_3255 = v_91 | v_3254;
assign v_3256 = ~v_89 | v_2956;
assign v_3257 = v_91 | v_3256;
assign v_3259 = ~v_361 | v_3258;
assign v_3261 = ~v_89 | v_2964;
assign v_3262 = v_91 | v_3261;
assign v_3263 = ~v_89 | v_2969;
assign v_3264 = v_91 | v_3263;
assign v_3266 = ~v_563 | v_3265;
assign v_3268 = ~v_3243 | v_3267;
assign v_3273 = v_3271 | v_3272;
assign v_3275 = ~v_3250 | v_3274;
assign v_3277 = v_3275 | v_3276;
assign v_3282 = v_3279 | v_3281;
assign v_3284 = v_3277 | v_3283;
assign v_3289 = v_3286 | v_3288;
assign v_3291 = v_3284 | v_3290;
assign v_3292 = v_3243 | v_3291;
assign v_3299 = ~v_3293 | v_3298;
assign v_3300 = v_3274 | ~v_3294;
assign v_3301 = v_3276 | v_3300;
assign v_3302 = v_3283 | v_3301;
assign v_3303 = v_3290 | v_3302;
assign v_3304 = v_3293 | v_3303;
assign v_3311 = ~v_3305 | v_3310;
assign v_3312 = v_3274 | ~v_3306;
assign v_3313 = v_3276 | v_3312;
assign v_3314 = v_3283 | v_3313;
assign v_3315 = v_3290 | v_3314;
assign v_3316 = v_3305 | v_3315;
assign v_3323 = ~v_3317 | v_3322;
assign v_3324 = v_3274 | ~v_3318;
assign v_3325 = v_3276 | v_3324;
assign v_3326 = v_3283 | v_3325;
assign v_3327 = v_3290 | v_3326;
assign v_3328 = v_3317 | v_3327;
assign v_3335 = ~v_3329 | v_3334;
assign v_3336 = v_3274 | ~v_3330;
assign v_3337 = v_3276 | v_3336;
assign v_3338 = v_3283 | v_3337;
assign v_3339 = v_3290 | v_3338;
assign v_3340 = v_3329 | v_3339;
assign v_3347 = ~v_3341 | v_3346;
assign v_3348 = v_3274 | ~v_3342;
assign v_3349 = v_3276 | v_3348;
assign v_3350 = v_3283 | v_3349;
assign v_3351 = v_3290 | v_3350;
assign v_3352 = v_3341 | v_3351;
assign v_3357 = v_3355 | v_3356;
assign v_3360 = v_3358 | v_3359;
assign v_3363 = v_3361 | v_3362;
assign v_3366 = v_3364 | v_3365;
assign v_3367 = ~v_3353 | v_3366;
assign v_3368 = v_3274 | ~v_3354;
assign v_3369 = v_3249 | v_3272;
assign v_3371 = v_3276 | v_3370;
assign v_3372 = v_91 | v_3252;
assign v_3374 = v_3283 | v_3373;
assign v_3375 = v_3259 | v_3281;
assign v_3377 = v_3290 | v_3376;
assign v_3378 = v_3266 | v_3288;
assign v_3380 = v_3353 | v_3379;
assign v_3383 = v_3274 | v_3382;
assign v_3384 = v_3276 | v_3383;
assign v_3385 = v_3283 | v_3384;
assign v_3386 = v_3290 | v_3385;
assign v_3387 = ~v_3381 | v_3386;
assign v_3392 = v_3381 | v_3391;
assign v_3394 = ~v_96 | v_3245;
assign v_3397 = ~v_807 | v_2943;
assign v_3399 = ~v_91 | v_3254;
assign v_3400 = ~v_91 | v_3256;
assign v_3402 = ~v_361 | v_3401;
assign v_3404 = ~v_91 | v_3261;
assign v_3405 = ~v_91 | v_3263;
assign v_3407 = ~v_563 | v_3406;
assign v_3409 = ~v_3393 | v_3408;
assign v_3411 = ~v_3395 | v_3410;
assign v_3413 = v_3411 | v_3412;
assign v_3416 = v_3414 | v_3415;
assign v_3418 = v_3413 | v_3417;
assign v_3421 = v_3419 | v_3420;
assign v_3423 = v_3418 | v_3422;
assign v_3424 = v_3393 | v_3423;
assign v_3431 = ~v_3425 | v_3430;
assign v_3432 = v_3410 | ~v_3426;
assign v_3433 = v_3412 | v_3432;
assign v_3434 = v_3417 | v_3433;
assign v_3435 = v_3422 | v_3434;
assign v_3436 = v_3425 | v_3435;
assign v_3443 = ~v_3437 | v_3442;
assign v_3444 = v_3410 | ~v_3438;
assign v_3445 = v_3412 | v_3444;
assign v_3446 = v_3417 | v_3445;
assign v_3447 = v_3422 | v_3446;
assign v_3448 = v_3437 | v_3447;
assign v_3455 = ~v_3449 | v_3454;
assign v_3456 = v_3410 | ~v_3450;
assign v_3457 = v_3412 | v_3456;
assign v_3458 = v_3417 | v_3457;
assign v_3459 = v_3422 | v_3458;
assign v_3460 = v_3449 | v_3459;
assign v_3467 = ~v_3461 | v_3466;
assign v_3468 = v_3410 | ~v_3462;
assign v_3469 = v_3412 | v_3468;
assign v_3470 = v_3417 | v_3469;
assign v_3471 = v_3422 | v_3470;
assign v_3472 = v_3461 | v_3471;
assign v_3479 = ~v_3473 | v_3478;
assign v_3480 = v_3410 | ~v_3474;
assign v_3481 = v_3412 | v_3480;
assign v_3482 = v_3417 | v_3481;
assign v_3483 = v_3422 | v_3482;
assign v_3484 = v_3473 | v_3483;
assign v_3489 = v_3487 | v_3488;
assign v_3492 = v_3490 | v_3491;
assign v_3495 = v_3493 | v_3494;
assign v_3498 = v_3496 | v_3497;
assign v_3499 = ~v_3485 | v_3498;
assign v_3500 = v_3410 | ~v_3486;
assign v_3501 = ~v_91 | v_3394;
assign v_3503 = v_3412 | v_3502;
assign v_3504 = v_2977 | v_3397;
assign v_3506 = v_3417 | v_3505;
assign v_3507 = v_3402 | v_3415;
assign v_3509 = v_3422 | v_3508;
assign v_3510 = v_3407 | v_3420;
assign v_3512 = v_3485 | v_3511;
assign v_3519 = ~v_3513 | v_3518;
assign v_3520 = v_3410 | ~v_3514;
assign v_3521 = v_3412 | v_3520;
assign v_3522 = v_3417 | v_3521;
assign v_3523 = v_3422 | v_3522;
assign v_3524 = v_3513 | v_3523;
assign v_3526 = ~v_89 | v_3244;
assign v_3527 = v_91 | v_3526;
assign v_3528 = ~v_91 | v_3245;
assign v_3530 = ~v_96 | v_3529;
assign v_3533 = ~v_807 | v_2940;
assign v_3535 = v_87 | v_2950;
assign v_3536 = v_89 | v_3535;
assign v_3537 = v_91 | v_3536;
assign v_3538 = v_87 | v_2955;
assign v_3539 = v_89 | v_3538;
assign v_3540 = v_91 | v_3539;
assign v_3542 = ~v_361 | v_3541;
assign v_3544 = v_87 | v_2963;
assign v_3545 = v_89 | v_3544;
assign v_3546 = v_91 | v_3545;
assign v_3547 = v_87 | v_2968;
assign v_3548 = v_89 | v_3547;
assign v_3549 = v_91 | v_3548;
assign v_3551 = ~v_563 | v_3550;
assign v_3553 = ~v_3525 | v_3552;
assign v_3557 = v_3555 | v_3556;
assign v_3559 = ~v_3531 | v_3558;
assign v_3561 = v_3559 | v_3560;
assign v_3568 = v_3564 | v_3567;
assign v_3570 = v_3561 | v_3569;
assign v_3577 = v_3573 | v_3576;
assign v_3579 = v_3570 | v_3578;
assign v_3580 = v_3525 | v_3579;
assign v_3587 = ~v_3581 | v_3586;
assign v_3588 = v_3558 | ~v_3582;
assign v_3589 = v_3560 | v_3588;
assign v_3590 = v_3569 | v_3589;
assign v_3591 = v_3578 | v_3590;
assign v_3592 = v_3581 | v_3591;
assign v_3599 = ~v_3593 | v_3598;
assign v_3600 = v_3558 | ~v_3594;
assign v_3601 = v_3560 | v_3600;
assign v_3602 = v_3569 | v_3601;
assign v_3603 = v_3578 | v_3602;
assign v_3604 = v_3593 | v_3603;
assign v_3611 = ~v_3605 | v_3610;
assign v_3612 = v_3558 | ~v_3606;
assign v_3613 = v_3560 | v_3612;
assign v_3614 = v_3569 | v_3613;
assign v_3615 = v_3578 | v_3614;
assign v_3616 = v_3605 | v_3615;
assign v_3623 = ~v_3617 | v_3622;
assign v_3624 = v_3558 | ~v_3618;
assign v_3625 = v_3560 | v_3624;
assign v_3626 = v_3569 | v_3625;
assign v_3627 = v_3578 | v_3626;
assign v_3628 = v_3617 | v_3627;
assign v_3635 = ~v_3629 | v_3634;
assign v_3636 = v_3558 | ~v_3630;
assign v_3637 = v_3560 | v_3636;
assign v_3638 = v_3569 | v_3637;
assign v_3639 = v_3578 | v_3638;
assign v_3640 = v_3629 | v_3639;
assign v_3645 = v_3643 | v_3644;
assign v_3648 = v_3646 | v_3647;
assign v_3651 = v_3649 | v_3650;
assign v_3654 = v_3652 | v_3653;
assign v_3655 = ~v_3641 | v_3654;
assign v_3656 = v_3558 | ~v_3642;
assign v_3657 = v_3530 | v_3556;
assign v_3659 = v_3560 | v_3658;
assign v_3660 = v_91 | v_3533;
assign v_3662 = v_3569 | v_3661;
assign v_3663 = v_3542 | v_3567;
assign v_3665 = v_3578 | v_3664;
assign v_3666 = v_3551 | v_3576;
assign v_3668 = v_3641 | v_3667;
assign v_3671 = v_3558 | v_3670;
assign v_3672 = v_3560 | v_3671;
assign v_3673 = v_3569 | v_3672;
assign v_3674 = v_3578 | v_3673;
assign v_3675 = ~v_3669 | v_3674;
assign v_3680 = v_3669 | v_3679;
assign v_3682 = ~v_96 | v_3526;
assign v_3685 = ~v_807 | v_3248;
assign v_3687 = ~v_91 | v_3536;
assign v_3688 = ~v_91 | v_3539;
assign v_3690 = ~v_361 | v_3689;
assign v_3692 = ~v_91 | v_3545;
assign v_3693 = ~v_91 | v_3548;
assign v_3695 = ~v_563 | v_3694;
assign v_3697 = ~v_3681 | v_3696;
assign v_3699 = ~v_3683 | v_3698;
assign v_3701 = v_3699 | v_3700;
assign v_3704 = v_3702 | v_3703;
assign v_3706 = v_3701 | v_3705;
assign v_3709 = v_3707 | v_3708;
assign v_3711 = v_3706 | v_3710;
assign v_3712 = v_3681 | v_3711;
assign v_3719 = ~v_3713 | v_3718;
assign v_3720 = v_3698 | ~v_3714;
assign v_3721 = v_3700 | v_3720;
assign v_3722 = v_3705 | v_3721;
assign v_3723 = v_3710 | v_3722;
assign v_3724 = v_3713 | v_3723;
assign v_3731 = ~v_3725 | v_3730;
assign v_3732 = v_3698 | ~v_3726;
assign v_3733 = v_3700 | v_3732;
assign v_3734 = v_3705 | v_3733;
assign v_3735 = v_3710 | v_3734;
assign v_3736 = v_3725 | v_3735;
assign v_3743 = ~v_3737 | v_3742;
assign v_3744 = v_3698 | ~v_3738;
assign v_3745 = v_3700 | v_3744;
assign v_3746 = v_3705 | v_3745;
assign v_3747 = v_3710 | v_3746;
assign v_3748 = v_3737 | v_3747;
assign v_3755 = ~v_3749 | v_3754;
assign v_3756 = v_3698 | ~v_3750;
assign v_3757 = v_3700 | v_3756;
assign v_3758 = v_3705 | v_3757;
assign v_3759 = v_3710 | v_3758;
assign v_3760 = v_3749 | v_3759;
assign v_3767 = ~v_3761 | v_3766;
assign v_3768 = v_3698 | ~v_3762;
assign v_3769 = v_3700 | v_3768;
assign v_3770 = v_3705 | v_3769;
assign v_3771 = v_3710 | v_3770;
assign v_3772 = v_3761 | v_3771;
assign v_3777 = v_3775 | v_3776;
assign v_3780 = v_3778 | v_3779;
assign v_3783 = v_3781 | v_3782;
assign v_3786 = v_3784 | v_3785;
assign v_3787 = ~v_3773 | v_3786;
assign v_3788 = v_3698 | ~v_3774;
assign v_3789 = ~v_91 | v_3682;
assign v_3791 = v_3700 | v_3790;
assign v_3792 = v_3271 | v_3685;
assign v_3794 = v_3705 | v_3793;
assign v_3795 = v_3690 | v_3703;
assign v_3797 = v_3710 | v_3796;
assign v_3798 = v_3695 | v_3708;
assign v_3800 = v_3773 | v_3799;
assign v_3803 = v_3698 | v_3802;
assign v_3804 = v_3700 | v_3803;
assign v_3805 = v_3705 | v_3804;
assign v_3806 = v_3710 | v_3805;
assign v_3807 = ~v_3801 | v_3806;
assign v_3812 = v_3801 | v_3811;
assign v_3814 = v_587 | v_2654;
assign v_3815 = ~v_87 | v_3814;
assign v_3816 = v_89 | v_3815;
assign v_3817 = v_91 | v_3816;
assign v_3818 = ~v_91 | v_3526;
assign v_3820 = ~v_96 | v_3819;
assign v_3823 = ~v_807 | v_3245;
assign v_3825 = ~v_89 | v_3535;
assign v_3826 = v_91 | v_3825;
assign v_3827 = ~v_89 | v_3538;
assign v_3828 = v_91 | v_3827;
assign v_3830 = ~v_361 | v_3829;
assign v_3832 = ~v_89 | v_3544;
assign v_3833 = v_91 | v_3832;
assign v_3834 = ~v_89 | v_3547;
assign v_3835 = v_91 | v_3834;
assign v_3837 = ~v_563 | v_3836;
assign v_3839 = ~v_3813 | v_3838;
assign v_3845 = v_3843 | v_3844;
assign v_3847 = ~v_3821 | v_3846;
assign v_3849 = v_3847 | v_3848;
assign v_3854 = v_3851 | v_3853;
assign v_3856 = v_3849 | v_3855;
assign v_3861 = v_3858 | v_3860;
assign v_3863 = v_3856 | v_3862;
assign v_3864 = v_3813 | v_3863;
assign v_3871 = ~v_3865 | v_3870;
assign v_3872 = v_3846 | ~v_3866;
assign v_3873 = v_3848 | v_3872;
assign v_3874 = v_3855 | v_3873;
assign v_3875 = v_3862 | v_3874;
assign v_3876 = v_3865 | v_3875;
assign v_3883 = ~v_3877 | v_3882;
assign v_3884 = v_3846 | ~v_3878;
assign v_3885 = v_3848 | v_3884;
assign v_3886 = v_3855 | v_3885;
assign v_3887 = v_3862 | v_3886;
assign v_3888 = v_3877 | v_3887;
assign v_3895 = ~v_3889 | v_3894;
assign v_3896 = v_3846 | ~v_3890;
assign v_3897 = v_3848 | v_3896;
assign v_3898 = v_3855 | v_3897;
assign v_3899 = v_3862 | v_3898;
assign v_3900 = v_3889 | v_3899;
assign v_3907 = ~v_3901 | v_3906;
assign v_3908 = v_3846 | ~v_3902;
assign v_3909 = v_3848 | v_3908;
assign v_3910 = v_3855 | v_3909;
assign v_3911 = v_3862 | v_3910;
assign v_3912 = v_3901 | v_3911;
assign v_3919 = ~v_3913 | v_3918;
assign v_3920 = v_3846 | ~v_3914;
assign v_3921 = v_3848 | v_3920;
assign v_3922 = v_3855 | v_3921;
assign v_3923 = v_3862 | v_3922;
assign v_3924 = v_3913 | v_3923;
assign v_3929 = v_3927 | v_3928;
assign v_3932 = v_3930 | v_3931;
assign v_3935 = v_3933 | v_3934;
assign v_3938 = v_3936 | v_3937;
assign v_3939 = ~v_3925 | v_3938;
assign v_3940 = v_3846 | ~v_3926;
assign v_3941 = v_3820 | v_3844;
assign v_3943 = v_3848 | v_3942;
assign v_3944 = v_91 | v_3823;
assign v_3946 = v_3855 | v_3945;
assign v_3947 = v_3830 | v_3853;
assign v_3949 = v_3862 | v_3948;
assign v_3950 = v_3837 | v_3860;
assign v_3952 = v_3925 | v_3951;
assign v_3955 = v_3846 | v_3954;
assign v_3956 = v_3848 | v_3955;
assign v_3957 = v_3855 | v_3956;
assign v_3958 = v_3862 | v_3957;
assign v_3959 = ~v_3953 | v_3958;
assign v_3964 = v_3953 | v_3963;
assign v_3966 = ~v_96 | v_3816;
assign v_3969 = ~v_807 | v_3529;
assign v_3971 = ~v_91 | v_3825;
assign v_3972 = ~v_91 | v_3827;
assign v_3974 = ~v_361 | v_3973;
assign v_3976 = ~v_91 | v_3832;
assign v_3977 = ~v_91 | v_3834;
assign v_3979 = ~v_563 | v_3978;
assign v_3981 = ~v_3965 | v_3980;
assign v_3983 = ~v_3967 | v_3982;
assign v_3985 = v_3983 | v_3984;
assign v_3988 = v_3986 | v_3987;
assign v_3990 = v_3985 | v_3989;
assign v_3993 = v_3991 | v_3992;
assign v_3995 = v_3990 | v_3994;
assign v_3996 = v_3965 | v_3995;
assign v_4003 = ~v_3997 | v_4002;
assign v_4004 = v_3982 | ~v_3998;
assign v_4005 = v_3984 | v_4004;
assign v_4006 = v_3989 | v_4005;
assign v_4007 = v_3994 | v_4006;
assign v_4008 = v_3997 | v_4007;
assign v_4015 = ~v_4009 | v_4014;
assign v_4016 = v_3982 | ~v_4010;
assign v_4017 = v_3984 | v_4016;
assign v_4018 = v_3989 | v_4017;
assign v_4019 = v_3994 | v_4018;
assign v_4020 = v_4009 | v_4019;
assign v_4027 = ~v_4021 | v_4026;
assign v_4028 = v_3982 | ~v_4022;
assign v_4029 = v_3984 | v_4028;
assign v_4030 = v_3989 | v_4029;
assign v_4031 = v_3994 | v_4030;
assign v_4032 = v_4021 | v_4031;
assign v_4039 = ~v_4033 | v_4038;
assign v_4040 = v_3982 | ~v_4034;
assign v_4041 = v_3984 | v_4040;
assign v_4042 = v_3989 | v_4041;
assign v_4043 = v_3994 | v_4042;
assign v_4044 = v_4033 | v_4043;
assign v_4051 = ~v_4045 | v_4050;
assign v_4052 = v_3982 | ~v_4046;
assign v_4053 = v_3984 | v_4052;
assign v_4054 = v_3989 | v_4053;
assign v_4055 = v_3994 | v_4054;
assign v_4056 = v_4045 | v_4055;
assign v_4061 = v_4059 | v_4060;
assign v_4064 = v_4062 | v_4063;
assign v_4067 = v_4065 | v_4066;
assign v_4070 = v_4068 | v_4069;
assign v_4071 = ~v_4057 | v_4070;
assign v_4072 = v_3982 | ~v_4058;
assign v_4073 = ~v_91 | v_3966;
assign v_4075 = v_3984 | v_4074;
assign v_4076 = v_3555 | v_3969;
assign v_4078 = v_3989 | v_4077;
assign v_4079 = v_3974 | v_3987;
assign v_4081 = v_3994 | v_4080;
assign v_4082 = v_3979 | v_3992;
assign v_4084 = v_4057 | v_4083;
assign v_4087 = v_3982 | v_4086;
assign v_4088 = v_3984 | v_4087;
assign v_4089 = v_3989 | v_4088;
assign v_4090 = v_3994 | v_4089;
assign v_4091 = ~v_4085 | v_4090;
assign v_4096 = v_4085 | v_4095;
assign v_4098 = ~v_89 | v_3815;
assign v_4099 = v_91 | v_4098;
assign v_4100 = ~v_91 | v_3816;
assign v_4102 = ~v_96 | v_4101;
assign v_4105 = ~v_807 | v_3526;
assign v_4107 = v_587 | v_2949;
assign v_4108 = ~v_87 | v_4107;
assign v_4109 = v_89 | v_4108;
assign v_4110 = v_91 | v_4109;
assign v_4111 = v_654 | v_2954;
assign v_4112 = ~v_87 | v_4111;
assign v_4113 = v_89 | v_4112;
assign v_4114 = v_91 | v_4113;
assign v_4116 = ~v_361 | v_4115;
assign v_4118 = v_587 | v_2962;
assign v_4119 = ~v_87 | v_4118;
assign v_4120 = v_89 | v_4119;
assign v_4121 = v_91 | v_4120;
assign v_4122 = v_654 | v_2967;
assign v_4123 = ~v_87 | v_4122;
assign v_4124 = v_89 | v_4123;
assign v_4125 = v_91 | v_4124;
assign v_4127 = ~v_563 | v_4126;
assign v_4129 = ~v_4097 | v_4128;
assign v_4133 = v_4131 | v_4132;
assign v_4135 = ~v_4103 | v_4134;
assign v_4137 = v_4135 | v_4136;
assign v_4146 = v_4141 | v_4145;
assign v_4148 = v_4137 | v_4147;
assign v_4157 = v_4152 | v_4156;
assign v_4159 = v_4148 | v_4158;
assign v_4160 = v_4097 | v_4159;
assign v_4167 = ~v_4161 | v_4166;
assign v_4168 = v_4134 | ~v_4162;
assign v_4169 = v_4136 | v_4168;
assign v_4170 = v_4147 | v_4169;
assign v_4171 = v_4158 | v_4170;
assign v_4172 = v_4161 | v_4171;
assign v_4179 = ~v_4173 | v_4178;
assign v_4180 = v_4134 | ~v_4174;
assign v_4181 = v_4136 | v_4180;
assign v_4182 = v_4147 | v_4181;
assign v_4183 = v_4158 | v_4182;
assign v_4184 = v_4173 | v_4183;
assign v_4191 = ~v_4185 | v_4190;
assign v_4192 = v_4134 | ~v_4186;
assign v_4193 = v_4136 | v_4192;
assign v_4194 = v_4147 | v_4193;
assign v_4195 = v_4158 | v_4194;
assign v_4196 = v_4185 | v_4195;
assign v_4203 = ~v_4197 | v_4202;
assign v_4204 = v_4134 | ~v_4198;
assign v_4205 = v_4136 | v_4204;
assign v_4206 = v_4147 | v_4205;
assign v_4207 = v_4158 | v_4206;
assign v_4208 = v_4197 | v_4207;
assign v_4215 = ~v_4209 | v_4214;
assign v_4216 = v_4134 | ~v_4210;
assign v_4217 = v_4136 | v_4216;
assign v_4218 = v_4147 | v_4217;
assign v_4219 = v_4158 | v_4218;
assign v_4220 = v_4209 | v_4219;
assign v_4225 = v_4223 | v_4224;
assign v_4228 = v_4226 | v_4227;
assign v_4231 = v_4229 | v_4230;
assign v_4234 = v_4232 | v_4233;
assign v_4235 = ~v_4221 | v_4234;
assign v_4236 = v_4134 | ~v_4222;
assign v_4237 = v_4102 | v_4132;
assign v_4239 = v_4136 | v_4238;
assign v_4240 = v_91 | v_4105;
assign v_4242 = v_4147 | v_4241;
assign v_4243 = v_4116 | v_4145;
assign v_4245 = v_4158 | v_4244;
assign v_4246 = v_4127 | v_4156;
assign v_4248 = v_4221 | v_4247;
assign v_4251 = v_4134 | v_4250;
assign v_4252 = v_4136 | v_4251;
assign v_4253 = v_4147 | v_4252;
assign v_4254 = v_4158 | v_4253;
assign v_4255 = ~v_4249 | v_4254;
assign v_4260 = v_4249 | v_4259;
assign v_4262 = ~v_96 | v_4098;
assign v_4265 = ~v_807 | v_3819;
assign v_4267 = ~v_91 | v_4109;
assign v_4268 = ~v_91 | v_4113;
assign v_4270 = ~v_361 | v_4269;
assign v_4272 = ~v_91 | v_4120;
assign v_4273 = ~v_91 | v_4124;
assign v_4275 = ~v_563 | v_4274;
assign v_4277 = ~v_4261 | v_4276;
assign v_4279 = ~v_4263 | v_4278;
assign v_4281 = v_4279 | v_4280;
assign v_4284 = v_4282 | v_4283;
assign v_4286 = v_4281 | v_4285;
assign v_4289 = v_4287 | v_4288;
assign v_4291 = v_4286 | v_4290;
assign v_4292 = v_4261 | v_4291;
assign v_4299 = ~v_4293 | v_4298;
assign v_4300 = v_4278 | ~v_4294;
assign v_4301 = v_4280 | v_4300;
assign v_4302 = v_4285 | v_4301;
assign v_4303 = v_4290 | v_4302;
assign v_4304 = v_4293 | v_4303;
assign v_4311 = ~v_4305 | v_4310;
assign v_4312 = v_4278 | ~v_4306;
assign v_4313 = v_4280 | v_4312;
assign v_4314 = v_4285 | v_4313;
assign v_4315 = v_4290 | v_4314;
assign v_4316 = v_4305 | v_4315;
assign v_4323 = ~v_4317 | v_4322;
assign v_4324 = v_4278 | ~v_4318;
assign v_4325 = v_4280 | v_4324;
assign v_4326 = v_4285 | v_4325;
assign v_4327 = v_4290 | v_4326;
assign v_4328 = v_4317 | v_4327;
assign v_4335 = ~v_4329 | v_4334;
assign v_4336 = v_4278 | ~v_4330;
assign v_4337 = v_4280 | v_4336;
assign v_4338 = v_4285 | v_4337;
assign v_4339 = v_4290 | v_4338;
assign v_4340 = v_4329 | v_4339;
assign v_4347 = ~v_4341 | v_4346;
assign v_4348 = v_4278 | ~v_4342;
assign v_4349 = v_4280 | v_4348;
assign v_4350 = v_4285 | v_4349;
assign v_4351 = v_4290 | v_4350;
assign v_4352 = v_4341 | v_4351;
assign v_4357 = v_4355 | v_4356;
assign v_4360 = v_4358 | v_4359;
assign v_4363 = v_4361 | v_4362;
assign v_4366 = v_4364 | v_4365;
assign v_4367 = ~v_4353 | v_4366;
assign v_4368 = v_4278 | ~v_4354;
assign v_4369 = ~v_91 | v_4262;
assign v_4371 = v_4280 | v_4370;
assign v_4372 = v_3843 | v_4265;
assign v_4374 = v_4285 | v_4373;
assign v_4375 = v_4270 | v_4283;
assign v_4377 = v_4290 | v_4376;
assign v_4378 = v_4275 | v_4288;
assign v_4380 = v_4353 | v_4379;
assign v_4387 = ~v_4381 | v_4386;
assign v_4388 = v_4278 | ~v_4382;
assign v_4389 = v_4280 | v_4388;
assign v_4390 = v_4285 | v_4389;
assign v_4391 = v_4290 | v_4390;
assign v_4392 = v_4381 | v_4391;
assign v_4394 = v_87 | v_3814;
assign v_4395 = v_89 | v_4394;
assign v_4396 = v_91 | v_4395;
assign v_4397 = ~v_91 | v_4098;
assign v_4399 = ~v_96 | v_4398;
assign v_4402 = ~v_807 | v_3816;
assign v_4404 = ~v_89 | v_4108;
assign v_4405 = v_91 | v_4404;
assign v_4406 = ~v_89 | v_4112;
assign v_4407 = v_91 | v_4406;
assign v_4409 = ~v_361 | v_4408;
assign v_4411 = ~v_89 | v_4119;
assign v_4412 = v_91 | v_4411;
assign v_4413 = ~v_89 | v_4123;
assign v_4414 = v_91 | v_4413;
assign v_4416 = ~v_563 | v_4415;
assign v_4418 = ~v_4393 | v_4417;
assign v_4423 = v_4421 | v_4422;
assign v_4425 = ~v_4400 | v_4424;
assign v_4427 = v_4425 | v_4426;
assign v_4432 = v_4429 | v_4431;
assign v_4434 = v_4427 | v_4433;
assign v_4439 = v_4436 | v_4438;
assign v_4441 = v_4434 | v_4440;
assign v_4442 = v_4393 | v_4441;
assign v_4449 = ~v_4443 | v_4448;
assign v_4450 = v_4424 | ~v_4444;
assign v_4451 = v_4426 | v_4450;
assign v_4452 = v_4433 | v_4451;
assign v_4453 = v_4440 | v_4452;
assign v_4454 = v_4443 | v_4453;
assign v_4461 = ~v_4455 | v_4460;
assign v_4462 = v_4424 | ~v_4456;
assign v_4463 = v_4426 | v_4462;
assign v_4464 = v_4433 | v_4463;
assign v_4465 = v_4440 | v_4464;
assign v_4466 = v_4455 | v_4465;
assign v_4473 = ~v_4467 | v_4472;
assign v_4474 = v_4424 | ~v_4468;
assign v_4475 = v_4426 | v_4474;
assign v_4476 = v_4433 | v_4475;
assign v_4477 = v_4440 | v_4476;
assign v_4478 = v_4467 | v_4477;
assign v_4485 = ~v_4479 | v_4484;
assign v_4486 = v_4424 | ~v_4480;
assign v_4487 = v_4426 | v_4486;
assign v_4488 = v_4433 | v_4487;
assign v_4489 = v_4440 | v_4488;
assign v_4490 = v_4479 | v_4489;
assign v_4497 = ~v_4491 | v_4496;
assign v_4498 = v_4424 | ~v_4492;
assign v_4499 = v_4426 | v_4498;
assign v_4500 = v_4433 | v_4499;
assign v_4501 = v_4440 | v_4500;
assign v_4502 = v_4491 | v_4501;
assign v_4507 = v_4505 | v_4506;
assign v_4510 = v_4508 | v_4509;
assign v_4513 = v_4511 | v_4512;
assign v_4516 = v_4514 | v_4515;
assign v_4517 = ~v_4503 | v_4516;
assign v_4518 = v_4424 | ~v_4504;
assign v_4519 = v_4399 | v_4422;
assign v_4521 = v_4426 | v_4520;
assign v_4522 = v_91 | v_4402;
assign v_4524 = v_4433 | v_4523;
assign v_4525 = v_4409 | v_4431;
assign v_4527 = v_4440 | v_4526;
assign v_4528 = v_4416 | v_4438;
assign v_4530 = v_4503 | v_4529;
assign v_4537 = ~v_4531 | v_4536;
assign v_4538 = v_4424 | ~v_4532;
assign v_4539 = v_4426 | v_4538;
assign v_4540 = v_4433 | v_4539;
assign v_4541 = v_4440 | v_4540;
assign v_4542 = v_4531 | v_4541;
assign v_4544 = ~v_96 | v_4395;
assign v_4547 = ~v_807 | v_4101;
assign v_4549 = ~v_91 | v_4404;
assign v_4550 = ~v_91 | v_4406;
assign v_4552 = ~v_361 | v_4551;
assign v_4554 = ~v_91 | v_4411;
assign v_4555 = ~v_91 | v_4413;
assign v_4557 = ~v_563 | v_4556;
assign v_4559 = ~v_4543 | v_4558;
assign v_4561 = ~v_4545 | v_4560;
assign v_4563 = v_4561 | v_4562;
assign v_4566 = v_4564 | v_4565;
assign v_4568 = v_4563 | v_4567;
assign v_4571 = v_4569 | v_4570;
assign v_4573 = v_4568 | v_4572;
assign v_4574 = v_4543 | v_4573;
assign v_4581 = ~v_4575 | v_4580;
assign v_4582 = v_4560 | ~v_4576;
assign v_4583 = v_4562 | v_4582;
assign v_4584 = v_4567 | v_4583;
assign v_4585 = v_4572 | v_4584;
assign v_4586 = v_4575 | v_4585;
assign v_4593 = ~v_4587 | v_4592;
assign v_4594 = v_4560 | ~v_4588;
assign v_4595 = v_4562 | v_4594;
assign v_4596 = v_4567 | v_4595;
assign v_4597 = v_4572 | v_4596;
assign v_4598 = v_4587 | v_4597;
assign v_4605 = ~v_4599 | v_4604;
assign v_4606 = v_4560 | ~v_4600;
assign v_4607 = v_4562 | v_4606;
assign v_4608 = v_4567 | v_4607;
assign v_4609 = v_4572 | v_4608;
assign v_4610 = v_4599 | v_4609;
assign v_4617 = ~v_4611 | v_4616;
assign v_4618 = v_4560 | ~v_4612;
assign v_4619 = v_4562 | v_4618;
assign v_4620 = v_4567 | v_4619;
assign v_4621 = v_4572 | v_4620;
assign v_4622 = v_4611 | v_4621;
assign v_4629 = ~v_4623 | v_4628;
assign v_4630 = v_4560 | ~v_4624;
assign v_4631 = v_4562 | v_4630;
assign v_4632 = v_4567 | v_4631;
assign v_4633 = v_4572 | v_4632;
assign v_4634 = v_4623 | v_4633;
assign v_4639 = v_4637 | v_4638;
assign v_4642 = v_4640 | v_4641;
assign v_4645 = v_4643 | v_4644;
assign v_4648 = v_4646 | v_4647;
assign v_4649 = ~v_4635 | v_4648;
assign v_4650 = v_4560 | ~v_4636;
assign v_4651 = ~v_91 | v_4544;
assign v_4653 = v_4562 | v_4652;
assign v_4654 = v_4131 | v_4547;
assign v_4656 = v_4567 | v_4655;
assign v_4657 = v_4552 | v_4565;
assign v_4659 = v_4572 | v_4658;
assign v_4660 = v_4557 | v_4570;
assign v_4662 = v_4635 | v_4661;
assign v_4669 = ~v_4663 | v_4668;
assign v_4670 = v_4560 | ~v_4664;
assign v_4671 = v_4562 | v_4670;
assign v_4672 = v_4567 | v_4671;
assign v_4673 = v_4572 | v_4672;
assign v_4674 = v_4663 | v_4673;
assign v_4676 = ~v_89 | v_4394;
assign v_4677 = v_91 | v_4676;
assign v_4678 = ~v_91 | v_4395;
assign v_4680 = ~v_96 | v_4679;
assign v_4683 = ~v_807 | v_4098;
assign v_4685 = v_87 | v_4107;
assign v_4686 = v_89 | v_4685;
assign v_4687 = v_91 | v_4686;
assign v_4688 = v_87 | v_4111;
assign v_4689 = v_89 | v_4688;
assign v_4690 = v_91 | v_4689;
assign v_4692 = ~v_361 | v_4691;
assign v_4694 = v_87 | v_4118;
assign v_4695 = v_89 | v_4694;
assign v_4696 = v_91 | v_4695;
assign v_4697 = v_87 | v_4122;
assign v_4698 = v_89 | v_4697;
assign v_4699 = v_91 | v_4698;
assign v_4701 = ~v_563 | v_4700;
assign v_4703 = ~v_4675 | v_4702;
assign v_4707 = v_4705 | v_4706;
assign v_4709 = ~v_4681 | v_4708;
assign v_4711 = v_4709 | v_4710;
assign v_4718 = v_4714 | v_4717;
assign v_4720 = v_4711 | v_4719;
assign v_4727 = v_4723 | v_4726;
assign v_4729 = v_4720 | v_4728;
assign v_4730 = v_4675 | v_4729;
assign v_4737 = ~v_4731 | v_4736;
assign v_4738 = v_4708 | ~v_4732;
assign v_4739 = v_4710 | v_4738;
assign v_4740 = v_4719 | v_4739;
assign v_4741 = v_4728 | v_4740;
assign v_4742 = v_4731 | v_4741;
assign v_4749 = ~v_4743 | v_4748;
assign v_4750 = v_4708 | ~v_4744;
assign v_4751 = v_4710 | v_4750;
assign v_4752 = v_4719 | v_4751;
assign v_4753 = v_4728 | v_4752;
assign v_4754 = v_4743 | v_4753;
assign v_4761 = ~v_4755 | v_4760;
assign v_4762 = v_4708 | ~v_4756;
assign v_4763 = v_4710 | v_4762;
assign v_4764 = v_4719 | v_4763;
assign v_4765 = v_4728 | v_4764;
assign v_4766 = v_4755 | v_4765;
assign v_4773 = ~v_4767 | v_4772;
assign v_4774 = v_4708 | ~v_4768;
assign v_4775 = v_4710 | v_4774;
assign v_4776 = v_4719 | v_4775;
assign v_4777 = v_4728 | v_4776;
assign v_4778 = v_4767 | v_4777;
assign v_4785 = ~v_4779 | v_4784;
assign v_4786 = v_4708 | ~v_4780;
assign v_4787 = v_4710 | v_4786;
assign v_4788 = v_4719 | v_4787;
assign v_4789 = v_4728 | v_4788;
assign v_4790 = v_4779 | v_4789;
assign v_4795 = v_4793 | v_4794;
assign v_4798 = v_4796 | v_4797;
assign v_4801 = v_4799 | v_4800;
assign v_4804 = v_4802 | v_4803;
assign v_4805 = ~v_4791 | v_4804;
assign v_4806 = v_4708 | ~v_4792;
assign v_4807 = v_4680 | v_4706;
assign v_4809 = v_4710 | v_4808;
assign v_4810 = v_91 | v_4683;
assign v_4812 = v_4719 | v_4811;
assign v_4813 = v_4692 | v_4717;
assign v_4815 = v_4728 | v_4814;
assign v_4816 = v_4701 | v_4726;
assign v_4818 = v_4791 | v_4817;
assign v_4825 = ~v_4819 | v_4824;
assign v_4826 = v_4708 | ~v_4820;
assign v_4827 = v_4710 | v_4826;
assign v_4828 = v_4719 | v_4827;
assign v_4829 = v_4728 | v_4828;
assign v_4830 = v_4819 | v_4829;
assign v_4832 = ~v_96 | v_4676;
assign v_4835 = ~v_807 | v_4398;
assign v_4837 = ~v_91 | v_4686;
assign v_4838 = ~v_91 | v_4689;
assign v_4840 = ~v_361 | v_4839;
assign v_4842 = ~v_91 | v_4695;
assign v_4843 = ~v_91 | v_4698;
assign v_4845 = ~v_563 | v_4844;
assign v_4847 = ~v_4831 | v_4846;
assign v_4849 = ~v_4833 | v_4848;
assign v_4851 = v_4849 | v_4850;
assign v_4854 = v_4852 | v_4853;
assign v_4856 = v_4851 | v_4855;
assign v_4859 = v_4857 | v_4858;
assign v_4861 = v_4856 | v_4860;
assign v_4862 = v_4831 | v_4861;
assign v_4869 = ~v_4863 | v_4868;
assign v_4870 = v_4848 | ~v_4864;
assign v_4871 = v_4850 | v_4870;
assign v_4872 = v_4855 | v_4871;
assign v_4873 = v_4860 | v_4872;
assign v_4874 = v_4863 | v_4873;
assign v_4881 = ~v_4875 | v_4880;
assign v_4882 = v_4848 | ~v_4876;
assign v_4883 = v_4850 | v_4882;
assign v_4884 = v_4855 | v_4883;
assign v_4885 = v_4860 | v_4884;
assign v_4886 = v_4875 | v_4885;
assign v_4893 = ~v_4887 | v_4892;
assign v_4894 = v_4848 | ~v_4888;
assign v_4895 = v_4850 | v_4894;
assign v_4896 = v_4855 | v_4895;
assign v_4897 = v_4860 | v_4896;
assign v_4898 = v_4887 | v_4897;
assign v_4905 = ~v_4899 | v_4904;
assign v_4906 = v_4848 | ~v_4900;
assign v_4907 = v_4850 | v_4906;
assign v_4908 = v_4855 | v_4907;
assign v_4909 = v_4860 | v_4908;
assign v_4910 = v_4899 | v_4909;
assign v_4917 = ~v_4911 | v_4916;
assign v_4918 = v_4848 | ~v_4912;
assign v_4919 = v_4850 | v_4918;
assign v_4920 = v_4855 | v_4919;
assign v_4921 = v_4860 | v_4920;
assign v_4922 = v_4911 | v_4921;
assign v_4927 = v_4925 | v_4926;
assign v_4930 = v_4928 | v_4929;
assign v_4933 = v_4931 | v_4932;
assign v_4936 = v_4934 | v_4935;
assign v_4937 = ~v_4923 | v_4936;
assign v_4938 = v_4848 | ~v_4924;
assign v_4939 = ~v_91 | v_4832;
assign v_4941 = v_4850 | v_4940;
assign v_4942 = v_4421 | v_4835;
assign v_4944 = v_4855 | v_4943;
assign v_4945 = v_4840 | v_4853;
assign v_4947 = v_4860 | v_4946;
assign v_4948 = v_4845 | v_4858;
assign v_4950 = v_4923 | v_4949;
assign v_4957 = ~v_4951 | v_4956;
assign v_4958 = v_4848 | ~v_4952;
assign v_4959 = v_4850 | v_4958;
assign v_4960 = v_4855 | v_4959;
assign v_4961 = v_4860 | v_4960;
assign v_4962 = v_4951 | v_4961;
assign v_4964 = v_77 | v_581;
assign v_4965 = v_82 | v_4964;
assign v_4966 = v_85 | v_4965;
assign v_4967 = ~v_87 | v_4966;
assign v_4968 = v_89 | v_4967;
assign v_4969 = v_91 | v_4968;
assign v_4970 = ~v_91 | v_4676;
assign v_4972 = ~v_96 | v_4971;
assign v_4975 = ~v_807 | v_4395;
assign v_4977 = ~v_89 | v_4685;
assign v_4978 = v_91 | v_4977;
assign v_4979 = ~v_89 | v_4688;
assign v_4980 = v_91 | v_4979;
assign v_4982 = ~v_361 | v_4981;
assign v_4984 = ~v_89 | v_4694;
assign v_4985 = v_91 | v_4984;
assign v_4986 = ~v_89 | v_4697;
assign v_4987 = v_91 | v_4986;
assign v_4989 = ~v_563 | v_4988;
assign v_4991 = ~v_4963 | v_4990;
assign v_4999 = v_4997 | v_4998;
assign v_5001 = ~v_4973 | v_5000;
assign v_5003 = v_5001 | v_5002;
assign v_5008 = v_5005 | v_5007;
assign v_5010 = v_5003 | v_5009;
assign v_5015 = v_5012 | v_5014;
assign v_5017 = v_5010 | v_5016;
assign v_5018 = v_4963 | v_5017;
assign v_5025 = ~v_5019 | v_5024;
assign v_5026 = v_5000 | ~v_5020;
assign v_5027 = v_5002 | v_5026;
assign v_5028 = v_5009 | v_5027;
assign v_5029 = v_5016 | v_5028;
assign v_5030 = v_5019 | v_5029;
assign v_5037 = ~v_5031 | v_5036;
assign v_5038 = v_5000 | ~v_5032;
assign v_5039 = v_5002 | v_5038;
assign v_5040 = v_5009 | v_5039;
assign v_5041 = v_5016 | v_5040;
assign v_5042 = v_5031 | v_5041;
assign v_5049 = ~v_5043 | v_5048;
assign v_5050 = v_5000 | ~v_5044;
assign v_5051 = v_5002 | v_5050;
assign v_5052 = v_5009 | v_5051;
assign v_5053 = v_5016 | v_5052;
assign v_5054 = v_5043 | v_5053;
assign v_5061 = ~v_5055 | v_5060;
assign v_5062 = v_5000 | ~v_5056;
assign v_5063 = v_5002 | v_5062;
assign v_5064 = v_5009 | v_5063;
assign v_5065 = v_5016 | v_5064;
assign v_5066 = v_5055 | v_5065;
assign v_5073 = ~v_5067 | v_5072;
assign v_5074 = v_5000 | ~v_5068;
assign v_5075 = v_5002 | v_5074;
assign v_5076 = v_5009 | v_5075;
assign v_5077 = v_5016 | v_5076;
assign v_5078 = v_5067 | v_5077;
assign v_5083 = v_5081 | v_5082;
assign v_5086 = v_5084 | v_5085;
assign v_5089 = v_5087 | v_5088;
assign v_5092 = v_5090 | v_5091;
assign v_5093 = ~v_5079 | v_5092;
assign v_5094 = v_5000 | ~v_5080;
assign v_5095 = v_4972 | v_4998;
assign v_5097 = v_5002 | v_5096;
assign v_5098 = v_91 | v_4975;
assign v_5100 = v_5009 | v_5099;
assign v_5101 = v_4982 | v_5007;
assign v_5103 = v_5016 | v_5102;
assign v_5104 = v_4989 | v_5014;
assign v_5106 = v_5079 | v_5105;
assign v_5113 = ~v_5107 | v_5112;
assign v_5114 = v_5000 | ~v_5108;
assign v_5115 = v_5002 | v_5114;
assign v_5116 = v_5009 | v_5115;
assign v_5117 = v_5016 | v_5116;
assign v_5118 = v_5107 | v_5117;
assign v_5120 = ~v_96 | v_4968;
assign v_5123 = ~v_807 | v_4679;
assign v_5125 = ~v_91 | v_4977;
assign v_5126 = ~v_91 | v_4979;
assign v_5128 = ~v_361 | v_5127;
assign v_5130 = ~v_91 | v_4984;
assign v_5131 = ~v_91 | v_4986;
assign v_5133 = ~v_563 | v_5132;
assign v_5135 = ~v_5119 | v_5134;
assign v_5137 = ~v_5121 | v_5136;
assign v_5139 = v_5137 | v_5138;
assign v_5142 = v_5140 | v_5141;
assign v_5144 = v_5139 | v_5143;
assign v_5147 = v_5145 | v_5146;
assign v_5149 = v_5144 | v_5148;
assign v_5150 = v_5119 | v_5149;
assign v_5157 = ~v_5151 | v_5156;
assign v_5158 = v_5136 | ~v_5152;
assign v_5159 = v_5138 | v_5158;
assign v_5160 = v_5143 | v_5159;
assign v_5161 = v_5148 | v_5160;
assign v_5162 = v_5151 | v_5161;
assign v_5169 = ~v_5163 | v_5168;
assign v_5170 = v_5136 | ~v_5164;
assign v_5171 = v_5138 | v_5170;
assign v_5172 = v_5143 | v_5171;
assign v_5173 = v_5148 | v_5172;
assign v_5174 = v_5163 | v_5173;
assign v_5181 = ~v_5175 | v_5180;
assign v_5182 = v_5136 | ~v_5176;
assign v_5183 = v_5138 | v_5182;
assign v_5184 = v_5143 | v_5183;
assign v_5185 = v_5148 | v_5184;
assign v_5186 = v_5175 | v_5185;
assign v_5193 = ~v_5187 | v_5192;
assign v_5194 = v_5136 | ~v_5188;
assign v_5195 = v_5138 | v_5194;
assign v_5196 = v_5143 | v_5195;
assign v_5197 = v_5148 | v_5196;
assign v_5198 = v_5187 | v_5197;
assign v_5205 = ~v_5199 | v_5204;
assign v_5206 = v_5136 | ~v_5200;
assign v_5207 = v_5138 | v_5206;
assign v_5208 = v_5143 | v_5207;
assign v_5209 = v_5148 | v_5208;
assign v_5210 = v_5199 | v_5209;
assign v_5215 = v_5213 | v_5214;
assign v_5218 = v_5216 | v_5217;
assign v_5221 = v_5219 | v_5220;
assign v_5224 = v_5222 | v_5223;
assign v_5225 = ~v_5211 | v_5224;
assign v_5226 = v_5136 | ~v_5212;
assign v_5227 = ~v_91 | v_5120;
assign v_5229 = v_5138 | v_5228;
assign v_5230 = v_4705 | v_5123;
assign v_5232 = v_5143 | v_5231;
assign v_5233 = v_5128 | v_5141;
assign v_5235 = v_5148 | v_5234;
assign v_5236 = v_5133 | v_5146;
assign v_5238 = v_5211 | v_5237;
assign v_5241 = v_5136 | v_5240;
assign v_5242 = v_5138 | v_5241;
assign v_5243 = v_5143 | v_5242;
assign v_5244 = v_5148 | v_5243;
assign v_5245 = ~v_5239 | v_5244;
assign v_5250 = v_5239 | v_5249;
assign v_5252 = ~v_89 | v_4967;
assign v_5253 = v_91 | v_5252;
assign v_5254 = ~v_91 | v_4968;
assign v_5256 = ~v_96 | v_5255;
assign v_5259 = ~v_807 | v_4676;
assign v_5261 = v_213 | v_618;
assign v_5262 = v_218 | v_5261;
assign v_5263 = v_85 | v_5262;
assign v_5264 = ~v_87 | v_5263;
assign v_5265 = v_89 | v_5264;
assign v_5266 = v_91 | v_5265;
assign v_5267 = v_347 | v_648;
assign v_5268 = v_352 | v_5267;
assign v_5269 = v_355 | v_5268;
assign v_5270 = ~v_87 | v_5269;
assign v_5271 = v_89 | v_5270;
assign v_5272 = v_91 | v_5271;
assign v_5274 = ~v_361 | v_5273;
assign v_5276 = v_445 | v_681;
assign v_5277 = v_218 | v_5276;
assign v_5278 = v_85 | v_5277;
assign v_5279 = ~v_87 | v_5278;
assign v_5280 = v_89 | v_5279;
assign v_5281 = v_91 | v_5280;
assign v_5282 = v_551 | v_707;
assign v_5283 = v_556 | v_5282;
assign v_5284 = v_355 | v_5283;
assign v_5285 = ~v_87 | v_5284;
assign v_5286 = v_89 | v_5285;
assign v_5287 = v_91 | v_5286;
assign v_5289 = ~v_563 | v_5288;
assign v_5291 = ~v_5251 | v_5290;
assign v_5295 = v_5293 | v_5294;
assign v_5297 = ~v_5257 | v_5296;
assign v_5299 = v_5297 | v_5298;
assign v_5312 = v_5305 | v_5311;
assign v_5314 = v_5299 | v_5313;
assign v_5327 = v_5320 | v_5326;
assign v_5329 = v_5314 | v_5328;
assign v_5330 = v_5251 | v_5329;
assign v_5337 = ~v_5331 | v_5336;
assign v_5338 = v_5296 | ~v_5332;
assign v_5339 = v_5298 | v_5338;
assign v_5340 = v_5313 | v_5339;
assign v_5341 = v_5328 | v_5340;
assign v_5342 = v_5331 | v_5341;
assign v_5349 = ~v_5343 | v_5348;
assign v_5350 = v_5296 | ~v_5344;
assign v_5351 = v_5298 | v_5350;
assign v_5352 = v_5313 | v_5351;
assign v_5353 = v_5328 | v_5352;
assign v_5354 = v_5343 | v_5353;
assign v_5361 = ~v_5355 | v_5360;
assign v_5362 = v_5296 | ~v_5356;
assign v_5363 = v_5298 | v_5362;
assign v_5364 = v_5313 | v_5363;
assign v_5365 = v_5328 | v_5364;
assign v_5366 = v_5355 | v_5365;
assign v_5373 = ~v_5367 | v_5372;
assign v_5374 = v_5296 | ~v_5368;
assign v_5375 = v_5298 | v_5374;
assign v_5376 = v_5313 | v_5375;
assign v_5377 = v_5328 | v_5376;
assign v_5378 = v_5367 | v_5377;
assign v_5385 = ~v_5379 | v_5384;
assign v_5386 = v_5296 | ~v_5380;
assign v_5387 = v_5298 | v_5386;
assign v_5388 = v_5313 | v_5387;
assign v_5389 = v_5328 | v_5388;
assign v_5390 = v_5379 | v_5389;
assign v_5395 = v_5393 | v_5394;
assign v_5398 = v_5396 | v_5397;
assign v_5401 = v_5399 | v_5400;
assign v_5404 = v_5402 | v_5403;
assign v_5405 = ~v_5391 | v_5404;
assign v_5406 = v_5296 | ~v_5392;
assign v_5407 = v_5256 | v_5294;
assign v_5409 = v_5298 | v_5408;
assign v_5410 = v_91 | v_5259;
assign v_5412 = v_5313 | v_5411;
assign v_5413 = v_5274 | v_5311;
assign v_5415 = v_5328 | v_5414;
assign v_5416 = v_5289 | v_5326;
assign v_5418 = v_5391 | v_5417;
assign v_5421 = v_5296 | v_5420;
assign v_5422 = v_5298 | v_5421;
assign v_5423 = v_5313 | v_5422;
assign v_5424 = v_5328 | v_5423;
assign v_5425 = ~v_5419 | v_5424;
assign v_5430 = v_5419 | v_5429;
assign v_5432 = ~v_96 | v_5252;
assign v_5435 = ~v_807 | v_4971;
assign v_5437 = ~v_91 | v_5265;
assign v_5438 = ~v_91 | v_5271;
assign v_5440 = ~v_361 | v_5439;
assign v_5442 = ~v_91 | v_5280;
assign v_5443 = ~v_91 | v_5286;
assign v_5445 = ~v_563 | v_5444;
assign v_5447 = ~v_5431 | v_5446;
assign v_5449 = ~v_5433 | v_5448;
assign v_5451 = v_5449 | v_5450;
assign v_5454 = v_5452 | v_5453;
assign v_5456 = v_5451 | v_5455;
assign v_5459 = v_5457 | v_5458;
assign v_5461 = v_5456 | v_5460;
assign v_5462 = v_5431 | v_5461;
assign v_5469 = ~v_5463 | v_5468;
assign v_5470 = v_5448 | ~v_5464;
assign v_5471 = v_5450 | v_5470;
assign v_5472 = v_5455 | v_5471;
assign v_5473 = v_5460 | v_5472;
assign v_5474 = v_5463 | v_5473;
assign v_5481 = ~v_5475 | v_5480;
assign v_5482 = v_5448 | ~v_5476;
assign v_5483 = v_5450 | v_5482;
assign v_5484 = v_5455 | v_5483;
assign v_5485 = v_5460 | v_5484;
assign v_5486 = v_5475 | v_5485;
assign v_5493 = ~v_5487 | v_5492;
assign v_5494 = v_5448 | ~v_5488;
assign v_5495 = v_5450 | v_5494;
assign v_5496 = v_5455 | v_5495;
assign v_5497 = v_5460 | v_5496;
assign v_5498 = v_5487 | v_5497;
assign v_5505 = ~v_5499 | v_5504;
assign v_5506 = v_5448 | ~v_5500;
assign v_5507 = v_5450 | v_5506;
assign v_5508 = v_5455 | v_5507;
assign v_5509 = v_5460 | v_5508;
assign v_5510 = v_5499 | v_5509;
assign v_5517 = ~v_5511 | v_5516;
assign v_5518 = v_5448 | ~v_5512;
assign v_5519 = v_5450 | v_5518;
assign v_5520 = v_5455 | v_5519;
assign v_5521 = v_5460 | v_5520;
assign v_5522 = v_5511 | v_5521;
assign v_5527 = v_5525 | v_5526;
assign v_5530 = v_5528 | v_5529;
assign v_5533 = v_5531 | v_5532;
assign v_5536 = v_5534 | v_5535;
assign v_5537 = ~v_5523 | v_5536;
assign v_5538 = v_5448 | ~v_5524;
assign v_5539 = ~v_91 | v_5432;
assign v_5541 = v_5450 | v_5540;
assign v_5542 = v_4997 | v_5435;
assign v_5544 = v_5455 | v_5543;
assign v_5545 = v_5440 | v_5453;
assign v_5547 = v_5460 | v_5546;
assign v_5548 = v_5445 | v_5458;
assign v_5550 = v_5523 | v_5549;
assign v_5557 = ~v_5551 | v_5556;
assign v_5558 = v_5448 | ~v_5552;
assign v_5559 = v_5450 | v_5558;
assign v_5560 = v_5455 | v_5559;
assign v_5561 = v_5460 | v_5560;
assign v_5562 = v_5551 | v_5561;
assign v_5564 = v_87 | v_4966;
assign v_5565 = v_89 | v_5564;
assign v_5566 = v_91 | v_5565;
assign v_5567 = ~v_91 | v_5252;
assign v_5569 = ~v_96 | v_5568;
assign v_5572 = ~v_807 | v_4968;
assign v_5574 = ~v_89 | v_5264;
assign v_5575 = v_91 | v_5574;
assign v_5576 = ~v_89 | v_5270;
assign v_5577 = v_91 | v_5576;
assign v_5579 = ~v_361 | v_5578;
assign v_5581 = ~v_89 | v_5279;
assign v_5582 = v_91 | v_5581;
assign v_5583 = ~v_89 | v_5285;
assign v_5584 = v_91 | v_5583;
assign v_5586 = ~v_563 | v_5585;
assign v_5588 = ~v_5563 | v_5587;
assign v_5593 = v_5591 | v_5592;
assign v_5595 = ~v_5570 | v_5594;
assign v_5597 = v_5595 | v_5596;
assign v_5602 = v_5599 | v_5601;
assign v_5604 = v_5597 | v_5603;
assign v_5609 = v_5606 | v_5608;
assign v_5611 = v_5604 | v_5610;
assign v_5612 = v_5563 | v_5611;
assign v_5619 = ~v_5613 | v_5618;
assign v_5620 = v_5594 | ~v_5614;
assign v_5621 = v_5596 | v_5620;
assign v_5622 = v_5603 | v_5621;
assign v_5623 = v_5610 | v_5622;
assign v_5624 = v_5613 | v_5623;
assign v_5631 = ~v_5625 | v_5630;
assign v_5632 = v_5594 | ~v_5626;
assign v_5633 = v_5596 | v_5632;
assign v_5634 = v_5603 | v_5633;
assign v_5635 = v_5610 | v_5634;
assign v_5636 = v_5625 | v_5635;
assign v_5643 = ~v_5637 | v_5642;
assign v_5644 = v_5594 | ~v_5638;
assign v_5645 = v_5596 | v_5644;
assign v_5646 = v_5603 | v_5645;
assign v_5647 = v_5610 | v_5646;
assign v_5648 = v_5637 | v_5647;
assign v_5655 = ~v_5649 | v_5654;
assign v_5656 = v_5594 | ~v_5650;
assign v_5657 = v_5596 | v_5656;
assign v_5658 = v_5603 | v_5657;
assign v_5659 = v_5610 | v_5658;
assign v_5660 = v_5649 | v_5659;
assign v_5667 = ~v_5661 | v_5666;
assign v_5668 = v_5594 | ~v_5662;
assign v_5669 = v_5596 | v_5668;
assign v_5670 = v_5603 | v_5669;
assign v_5671 = v_5610 | v_5670;
assign v_5672 = v_5661 | v_5671;
assign v_5677 = v_5675 | v_5676;
assign v_5680 = v_5678 | v_5679;
assign v_5683 = v_5681 | v_5682;
assign v_5686 = v_5684 | v_5685;
assign v_5687 = ~v_5673 | v_5686;
assign v_5688 = v_5594 | ~v_5674;
assign v_5689 = v_5569 | v_5592;
assign v_5691 = v_5596 | v_5690;
assign v_5692 = v_91 | v_5572;
assign v_5694 = v_5603 | v_5693;
assign v_5695 = v_5579 | v_5601;
assign v_5697 = v_5610 | v_5696;
assign v_5698 = v_5586 | v_5608;
assign v_5700 = v_5673 | v_5699;
assign v_5707 = ~v_5701 | v_5706;
assign v_5708 = v_5594 | ~v_5702;
assign v_5709 = v_5596 | v_5708;
assign v_5710 = v_5603 | v_5709;
assign v_5711 = v_5610 | v_5710;
assign v_5712 = v_5701 | v_5711;
assign v_5714 = ~v_96 | v_5565;
assign v_5717 = ~v_807 | v_5255;
assign v_5719 = ~v_91 | v_5574;
assign v_5720 = ~v_91 | v_5576;
assign v_5722 = ~v_361 | v_5721;
assign v_5724 = ~v_91 | v_5581;
assign v_5725 = ~v_91 | v_5583;
assign v_5727 = ~v_563 | v_5726;
assign v_5729 = ~v_5713 | v_5728;
assign v_5731 = ~v_5715 | v_5730;
assign v_5733 = v_5731 | v_5732;
assign v_5736 = v_5734 | v_5735;
assign v_5738 = v_5733 | v_5737;
assign v_5741 = v_5739 | v_5740;
assign v_5743 = v_5738 | v_5742;
assign v_5744 = v_5713 | v_5743;
assign v_5751 = ~v_5745 | v_5750;
assign v_5752 = v_5730 | ~v_5746;
assign v_5753 = v_5732 | v_5752;
assign v_5754 = v_5737 | v_5753;
assign v_5755 = v_5742 | v_5754;
assign v_5756 = v_5745 | v_5755;
assign v_5763 = ~v_5757 | v_5762;
assign v_5764 = v_5730 | ~v_5758;
assign v_5765 = v_5732 | v_5764;
assign v_5766 = v_5737 | v_5765;
assign v_5767 = v_5742 | v_5766;
assign v_5768 = v_5757 | v_5767;
assign v_5775 = ~v_5769 | v_5774;
assign v_5776 = v_5730 | ~v_5770;
assign v_5777 = v_5732 | v_5776;
assign v_5778 = v_5737 | v_5777;
assign v_5779 = v_5742 | v_5778;
assign v_5780 = v_5769 | v_5779;
assign v_5787 = ~v_5781 | v_5786;
assign v_5788 = v_5730 | ~v_5782;
assign v_5789 = v_5732 | v_5788;
assign v_5790 = v_5737 | v_5789;
assign v_5791 = v_5742 | v_5790;
assign v_5792 = v_5781 | v_5791;
assign v_5799 = ~v_5793 | v_5798;
assign v_5800 = v_5730 | ~v_5794;
assign v_5801 = v_5732 | v_5800;
assign v_5802 = v_5737 | v_5801;
assign v_5803 = v_5742 | v_5802;
assign v_5804 = v_5793 | v_5803;
assign v_5807 = v_5730 | v_5806;
assign v_5808 = ~v_91 | v_5714;
assign v_5810 = v_5732 | v_5809;
assign v_5811 = v_5293 | v_5717;
assign v_5813 = v_5737 | v_5812;
assign v_5814 = v_5722 | v_5735;
assign v_5816 = v_5742 | v_5815;
assign v_5817 = v_5727 | v_5740;
assign v_5819 = ~v_5805 | v_5818;
assign v_5822 = v_5820 | v_5821;
assign v_5825 = v_5823 | v_5824;
assign v_5828 = v_5826 | v_5827;
assign v_5831 = v_5829 | v_5830;
assign v_5832 = v_5805 | v_5831;
assign v_5839 = ~v_5833 | v_5838;
assign v_5840 = v_5730 | ~v_5834;
assign v_5841 = v_5732 | v_5840;
assign v_5842 = v_5737 | v_5841;
assign v_5843 = v_5742 | v_5842;
assign v_5844 = v_5833 | v_5843;
assign v_5846 = ~v_89 | v_5564;
assign v_5847 = v_91 | v_5846;
assign v_5848 = ~v_91 | v_5565;
assign v_5850 = ~v_96 | v_5849;
assign v_5853 = ~v_807 | v_5252;
assign v_5855 = v_87 | v_5263;
assign v_5856 = v_89 | v_5855;
assign v_5857 = v_91 | v_5856;
assign v_5858 = v_87 | v_5269;
assign v_5859 = v_89 | v_5858;
assign v_5860 = v_91 | v_5859;
assign v_5862 = ~v_361 | v_5861;
assign v_5864 = v_87 | v_5278;
assign v_5865 = v_89 | v_5864;
assign v_5866 = v_91 | v_5865;
assign v_5867 = v_87 | v_5284;
assign v_5868 = v_89 | v_5867;
assign v_5869 = v_91 | v_5868;
assign v_5871 = ~v_563 | v_5870;
assign v_5873 = ~v_5845 | v_5872;
assign v_5877 = v_5875 | v_5876;
assign v_5879 = ~v_5851 | v_5878;
assign v_5881 = v_5879 | v_5880;
assign v_5888 = v_5884 | v_5887;
assign v_5890 = v_5881 | v_5889;
assign v_5897 = v_5893 | v_5896;
assign v_5899 = v_5890 | v_5898;
assign v_5900 = v_5845 | v_5899;
assign v_5907 = ~v_5901 | v_5906;
assign v_5908 = v_5878 | ~v_5902;
assign v_5909 = v_5880 | v_5908;
assign v_5910 = v_5889 | v_5909;
assign v_5911 = v_5898 | v_5910;
assign v_5912 = v_5901 | v_5911;
assign v_5919 = ~v_5913 | v_5918;
assign v_5920 = v_5878 | ~v_5914;
assign v_5921 = v_5880 | v_5920;
assign v_5922 = v_5889 | v_5921;
assign v_5923 = v_5898 | v_5922;
assign v_5924 = v_5913 | v_5923;
assign v_5931 = ~v_5925 | v_5930;
assign v_5932 = v_5878 | ~v_5926;
assign v_5933 = v_5880 | v_5932;
assign v_5934 = v_5889 | v_5933;
assign v_5935 = v_5898 | v_5934;
assign v_5936 = v_5925 | v_5935;
assign v_5943 = ~v_5937 | v_5942;
assign v_5944 = v_5878 | ~v_5938;
assign v_5945 = v_5880 | v_5944;
assign v_5946 = v_5889 | v_5945;
assign v_5947 = v_5898 | v_5946;
assign v_5948 = v_5937 | v_5947;
assign v_5955 = ~v_5949 | v_5954;
assign v_5956 = v_5878 | ~v_5950;
assign v_5957 = v_5880 | v_5956;
assign v_5958 = v_5889 | v_5957;
assign v_5959 = v_5898 | v_5958;
assign v_5960 = v_5949 | v_5959;
assign v_5965 = v_5963 | v_5964;
assign v_5968 = v_5966 | v_5967;
assign v_5971 = v_5969 | v_5970;
assign v_5974 = v_5972 | v_5973;
assign v_5975 = ~v_5961 | v_5974;
assign v_5976 = v_5878 | ~v_5962;
assign v_5977 = v_5850 | v_5876;
assign v_5979 = v_5880 | v_5978;
assign v_5980 = v_91 | v_5853;
assign v_5982 = v_5889 | v_5981;
assign v_5983 = v_5862 | v_5887;
assign v_5985 = v_5898 | v_5984;
assign v_5986 = v_5871 | v_5896;
assign v_5988 = v_5961 | v_5987;
assign v_5995 = ~v_5989 | v_5994;
assign v_5996 = v_5878 | ~v_5990;
assign v_5997 = v_5880 | v_5996;
assign v_5998 = v_5889 | v_5997;
assign v_5999 = v_5898 | v_5998;
assign v_6000 = v_5989 | v_5999;
assign v_6002 = ~v_96 | v_5846;
assign v_6005 = ~v_807 | v_5568;
assign v_6007 = ~v_91 | v_5856;
assign v_6008 = ~v_91 | v_5859;
assign v_6010 = ~v_361 | v_6009;
assign v_6012 = ~v_91 | v_5865;
assign v_6013 = ~v_91 | v_5868;
assign v_6015 = ~v_563 | v_6014;
assign v_6017 = ~v_6001 | v_6016;
assign v_6019 = ~v_6003 | v_6018;
assign v_6021 = v_6019 | v_6020;
assign v_6024 = v_6022 | v_6023;
assign v_6026 = v_6021 | v_6025;
assign v_6029 = v_6027 | v_6028;
assign v_6031 = v_6026 | v_6030;
assign v_6032 = v_6001 | v_6031;
assign v_6039 = ~v_6033 | v_6038;
assign v_6040 = v_6018 | ~v_6034;
assign v_6041 = v_6020 | v_6040;
assign v_6042 = v_6025 | v_6041;
assign v_6043 = v_6030 | v_6042;
assign v_6044 = v_6033 | v_6043;
assign v_6051 = ~v_6045 | v_6050;
assign v_6052 = v_6018 | ~v_6046;
assign v_6053 = v_6020 | v_6052;
assign v_6054 = v_6025 | v_6053;
assign v_6055 = v_6030 | v_6054;
assign v_6056 = v_6045 | v_6055;
assign v_6063 = ~v_6057 | v_6062;
assign v_6064 = v_6018 | ~v_6058;
assign v_6065 = v_6020 | v_6064;
assign v_6066 = v_6025 | v_6065;
assign v_6067 = v_6030 | v_6066;
assign v_6068 = v_6057 | v_6067;
assign v_6075 = ~v_6069 | v_6074;
assign v_6076 = v_6018 | ~v_6070;
assign v_6077 = v_6020 | v_6076;
assign v_6078 = v_6025 | v_6077;
assign v_6079 = v_6030 | v_6078;
assign v_6080 = v_6069 | v_6079;
assign v_6087 = ~v_6081 | v_6086;
assign v_6088 = v_6018 | ~v_6082;
assign v_6089 = v_6020 | v_6088;
assign v_6090 = v_6025 | v_6089;
assign v_6091 = v_6030 | v_6090;
assign v_6092 = v_6081 | v_6091;
assign v_6095 = v_6018 | v_6094;
assign v_6096 = ~v_91 | v_6002;
assign v_6098 = v_6020 | v_6097;
assign v_6099 = v_5591 | v_6005;
assign v_6101 = v_6025 | v_6100;
assign v_6102 = v_6010 | v_6023;
assign v_6104 = v_6030 | v_6103;
assign v_6105 = v_6015 | v_6028;
assign v_6107 = ~v_6093 | v_6106;
assign v_6110 = v_6108 | v_6109;
assign v_6113 = v_6111 | v_6112;
assign v_6116 = v_6114 | v_6115;
assign v_6119 = v_6117 | v_6118;
assign v_6120 = v_6093 | v_6119;
assign v_6127 = ~v_6121 | v_6126;
assign v_6128 = v_6018 | ~v_6122;
assign v_6129 = v_6020 | v_6128;
assign v_6130 = v_6025 | v_6129;
assign v_6131 = v_6030 | v_6130;
assign v_6132 = v_6121 | v_6131;
assign v_6134 = v_587 | v_4965;
assign v_6135 = ~v_87 | v_6134;
assign v_6136 = v_89 | v_6135;
assign v_6137 = v_91 | v_6136;
assign v_6138 = ~v_91 | v_5846;
assign v_6140 = ~v_96 | v_6139;
assign v_6143 = ~v_807 | v_5565;
assign v_6145 = ~v_89 | v_5855;
assign v_6146 = v_91 | v_6145;
assign v_6147 = ~v_89 | v_5858;
assign v_6148 = v_91 | v_6147;
assign v_6150 = ~v_361 | v_6149;
assign v_6152 = ~v_89 | v_5864;
assign v_6153 = v_91 | v_6152;
assign v_6154 = ~v_89 | v_5867;
assign v_6155 = v_91 | v_6154;
assign v_6157 = ~v_563 | v_6156;
assign v_6159 = ~v_6133 | v_6158;
assign v_6165 = v_6163 | v_6164;
assign v_6167 = ~v_6141 | v_6166;
assign v_6169 = v_6167 | v_6168;
assign v_6174 = v_6171 | v_6173;
assign v_6176 = v_6169 | v_6175;
assign v_6181 = v_6178 | v_6180;
assign v_6183 = v_6176 | v_6182;
assign v_6184 = v_6133 | v_6183;
assign v_6191 = ~v_6185 | v_6190;
assign v_6192 = v_6166 | ~v_6186;
assign v_6193 = v_6168 | v_6192;
assign v_6194 = v_6175 | v_6193;
assign v_6195 = v_6182 | v_6194;
assign v_6196 = v_6185 | v_6195;
assign v_6203 = ~v_6197 | v_6202;
assign v_6204 = v_6166 | ~v_6198;
assign v_6205 = v_6168 | v_6204;
assign v_6206 = v_6175 | v_6205;
assign v_6207 = v_6182 | v_6206;
assign v_6208 = v_6197 | v_6207;
assign v_6215 = ~v_6209 | v_6214;
assign v_6216 = v_6166 | ~v_6210;
assign v_6217 = v_6168 | v_6216;
assign v_6218 = v_6175 | v_6217;
assign v_6219 = v_6182 | v_6218;
assign v_6220 = v_6209 | v_6219;
assign v_6227 = ~v_6221 | v_6226;
assign v_6228 = v_6166 | ~v_6222;
assign v_6229 = v_6168 | v_6228;
assign v_6230 = v_6175 | v_6229;
assign v_6231 = v_6182 | v_6230;
assign v_6232 = v_6221 | v_6231;
assign v_6239 = ~v_6233 | v_6238;
assign v_6240 = v_6166 | ~v_6234;
assign v_6241 = v_6168 | v_6240;
assign v_6242 = v_6175 | v_6241;
assign v_6243 = v_6182 | v_6242;
assign v_6244 = v_6233 | v_6243;
assign v_6249 = v_6247 | v_6248;
assign v_6252 = v_6250 | v_6251;
assign v_6255 = v_6253 | v_6254;
assign v_6258 = v_6256 | v_6257;
assign v_6259 = ~v_6245 | v_6258;
assign v_6260 = v_6166 | ~v_6246;
assign v_6261 = v_6140 | v_6164;
assign v_6263 = v_6168 | v_6262;
assign v_6264 = v_91 | v_6143;
assign v_6266 = v_6175 | v_6265;
assign v_6267 = v_6150 | v_6173;
assign v_6269 = v_6182 | v_6268;
assign v_6270 = v_6157 | v_6180;
assign v_6272 = v_6245 | v_6271;
assign v_6279 = ~v_6273 | v_6278;
assign v_6280 = v_6166 | ~v_6274;
assign v_6281 = v_6168 | v_6280;
assign v_6282 = v_6175 | v_6281;
assign v_6283 = v_6182 | v_6282;
assign v_6284 = v_6273 | v_6283;
assign v_6286 = ~v_96 | v_6136;
assign v_6289 = ~v_807 | v_5849;
assign v_6291 = ~v_91 | v_6145;
assign v_6292 = ~v_91 | v_6147;
assign v_6294 = ~v_361 | v_6293;
assign v_6296 = ~v_91 | v_6152;
assign v_6297 = ~v_91 | v_6154;
assign v_6299 = ~v_563 | v_6298;
assign v_6301 = ~v_6285 | v_6300;
assign v_6303 = ~v_6287 | v_6302;
assign v_6305 = v_6303 | v_6304;
assign v_6308 = v_6306 | v_6307;
assign v_6310 = v_6305 | v_6309;
assign v_6313 = v_6311 | v_6312;
assign v_6315 = v_6310 | v_6314;
assign v_6316 = v_6285 | v_6315;
assign v_6323 = ~v_6317 | v_6322;
assign v_6324 = v_6302 | ~v_6318;
assign v_6325 = v_6304 | v_6324;
assign v_6326 = v_6309 | v_6325;
assign v_6327 = v_6314 | v_6326;
assign v_6328 = v_6317 | v_6327;
assign v_6335 = ~v_6329 | v_6334;
assign v_6336 = v_6302 | ~v_6330;
assign v_6337 = v_6304 | v_6336;
assign v_6338 = v_6309 | v_6337;
assign v_6339 = v_6314 | v_6338;
assign v_6340 = v_6329 | v_6339;
assign v_6347 = ~v_6341 | v_6346;
assign v_6348 = v_6302 | ~v_6342;
assign v_6349 = v_6304 | v_6348;
assign v_6350 = v_6309 | v_6349;
assign v_6351 = v_6314 | v_6350;
assign v_6352 = v_6341 | v_6351;
assign v_6359 = ~v_6353 | v_6358;
assign v_6360 = v_6302 | ~v_6354;
assign v_6361 = v_6304 | v_6360;
assign v_6362 = v_6309 | v_6361;
assign v_6363 = v_6314 | v_6362;
assign v_6364 = v_6353 | v_6363;
assign v_6371 = ~v_6365 | v_6370;
assign v_6372 = v_6302 | ~v_6366;
assign v_6373 = v_6304 | v_6372;
assign v_6374 = v_6309 | v_6373;
assign v_6375 = v_6314 | v_6374;
assign v_6376 = v_6365 | v_6375;
assign v_6381 = v_6379 | v_6380;
assign v_6384 = v_6382 | v_6383;
assign v_6387 = v_6385 | v_6386;
assign v_6390 = v_6388 | v_6389;
assign v_6391 = ~v_6377 | v_6390;
assign v_6392 = v_6302 | ~v_6378;
assign v_6393 = ~v_91 | v_6286;
assign v_6395 = v_6304 | v_6394;
assign v_6396 = v_5875 | v_6289;
assign v_6398 = v_6309 | v_6397;
assign v_6399 = v_6294 | v_6307;
assign v_6401 = v_6314 | v_6400;
assign v_6402 = v_6299 | v_6312;
assign v_6404 = v_6377 | v_6403;
assign v_6407 = v_6302 | v_6406;
assign v_6408 = v_6304 | v_6407;
assign v_6409 = v_6309 | v_6408;
assign v_6410 = v_6314 | v_6409;
assign v_6411 = ~v_6405 | v_6410;
assign v_6416 = v_6405 | v_6415;
assign v_6418 = ~v_89 | v_6135;
assign v_6419 = v_91 | v_6418;
assign v_6420 = ~v_91 | v_6136;
assign v_6422 = ~v_96 | v_6421;
assign v_6425 = ~v_807 | v_5846;
assign v_6427 = v_587 | v_5262;
assign v_6428 = ~v_87 | v_6427;
assign v_6429 = v_89 | v_6428;
assign v_6430 = v_91 | v_6429;
assign v_6431 = v_654 | v_5268;
assign v_6432 = ~v_87 | v_6431;
assign v_6433 = v_89 | v_6432;
assign v_6434 = v_91 | v_6433;
assign v_6436 = ~v_361 | v_6435;
assign v_6438 = v_587 | v_5277;
assign v_6439 = ~v_87 | v_6438;
assign v_6440 = v_89 | v_6439;
assign v_6441 = v_91 | v_6440;
assign v_6442 = v_654 | v_5283;
assign v_6443 = ~v_87 | v_6442;
assign v_6444 = v_89 | v_6443;
assign v_6445 = v_91 | v_6444;
assign v_6447 = ~v_563 | v_6446;
assign v_6449 = ~v_6417 | v_6448;
assign v_6453 = v_6451 | v_6452;
assign v_6455 = ~v_6423 | v_6454;
assign v_6457 = v_6455 | v_6456;
assign v_6466 = v_6461 | v_6465;
assign v_6468 = v_6457 | v_6467;
assign v_6477 = v_6472 | v_6476;
assign v_6479 = v_6468 | v_6478;
assign v_6480 = v_6417 | v_6479;
assign v_6487 = ~v_6481 | v_6486;
assign v_6488 = v_6454 | ~v_6482;
assign v_6489 = v_6456 | v_6488;
assign v_6490 = v_6467 | v_6489;
assign v_6491 = v_6478 | v_6490;
assign v_6492 = v_6481 | v_6491;
assign v_6499 = ~v_6493 | v_6498;
assign v_6500 = v_6454 | ~v_6494;
assign v_6501 = v_6456 | v_6500;
assign v_6502 = v_6467 | v_6501;
assign v_6503 = v_6478 | v_6502;
assign v_6504 = v_6493 | v_6503;
assign v_6511 = ~v_6505 | v_6510;
assign v_6512 = v_6454 | ~v_6506;
assign v_6513 = v_6456 | v_6512;
assign v_6514 = v_6467 | v_6513;
assign v_6515 = v_6478 | v_6514;
assign v_6516 = v_6505 | v_6515;
assign v_6523 = ~v_6517 | v_6522;
assign v_6524 = v_6454 | ~v_6518;
assign v_6525 = v_6456 | v_6524;
assign v_6526 = v_6467 | v_6525;
assign v_6527 = v_6478 | v_6526;
assign v_6528 = v_6517 | v_6527;
assign v_6535 = ~v_6529 | v_6534;
assign v_6536 = v_6454 | ~v_6530;
assign v_6537 = v_6456 | v_6536;
assign v_6538 = v_6467 | v_6537;
assign v_6539 = v_6478 | v_6538;
assign v_6540 = v_6529 | v_6539;
assign v_6545 = v_6543 | v_6544;
assign v_6548 = v_6546 | v_6547;
assign v_6551 = v_6549 | v_6550;
assign v_6554 = v_6552 | v_6553;
assign v_6555 = ~v_6541 | v_6554;
assign v_6556 = v_6454 | ~v_6542;
assign v_6557 = v_6422 | v_6452;
assign v_6559 = v_6456 | v_6558;
assign v_6560 = v_91 | v_6425;
assign v_6562 = v_6467 | v_6561;
assign v_6563 = v_6436 | v_6465;
assign v_6565 = v_6478 | v_6564;
assign v_6566 = v_6447 | v_6476;
assign v_6568 = v_6541 | v_6567;
assign v_6571 = v_6454 | v_6570;
assign v_6572 = v_6456 | v_6571;
assign v_6573 = v_6467 | v_6572;
assign v_6574 = v_6478 | v_6573;
assign v_6575 = ~v_6569 | v_6574;
assign v_6580 = v_6569 | v_6579;
assign v_6582 = ~v_96 | v_6418;
assign v_6585 = ~v_807 | v_6139;
assign v_6587 = ~v_91 | v_6429;
assign v_6588 = ~v_91 | v_6433;
assign v_6590 = ~v_361 | v_6589;
assign v_6592 = ~v_91 | v_6440;
assign v_6593 = ~v_91 | v_6444;
assign v_6595 = ~v_563 | v_6594;
assign v_6597 = ~v_6581 | v_6596;
assign v_6599 = ~v_6583 | v_6598;
assign v_6601 = v_6599 | v_6600;
assign v_6604 = v_6602 | v_6603;
assign v_6606 = v_6601 | v_6605;
assign v_6609 = v_6607 | v_6608;
assign v_6611 = v_6606 | v_6610;
assign v_6612 = v_6581 | v_6611;
assign v_6619 = ~v_6613 | v_6618;
assign v_6620 = v_6598 | ~v_6614;
assign v_6621 = v_6600 | v_6620;
assign v_6622 = v_6605 | v_6621;
assign v_6623 = v_6610 | v_6622;
assign v_6624 = v_6613 | v_6623;
assign v_6631 = ~v_6625 | v_6630;
assign v_6632 = v_6598 | ~v_6626;
assign v_6633 = v_6600 | v_6632;
assign v_6634 = v_6605 | v_6633;
assign v_6635 = v_6610 | v_6634;
assign v_6636 = v_6625 | v_6635;
assign v_6643 = ~v_6637 | v_6642;
assign v_6644 = v_6598 | ~v_6638;
assign v_6645 = v_6600 | v_6644;
assign v_6646 = v_6605 | v_6645;
assign v_6647 = v_6610 | v_6646;
assign v_6648 = v_6637 | v_6647;
assign v_6655 = ~v_6649 | v_6654;
assign v_6656 = v_6598 | ~v_6650;
assign v_6657 = v_6600 | v_6656;
assign v_6658 = v_6605 | v_6657;
assign v_6659 = v_6610 | v_6658;
assign v_6660 = v_6649 | v_6659;
assign v_6667 = ~v_6661 | v_6666;
assign v_6668 = v_6598 | ~v_6662;
assign v_6669 = v_6600 | v_6668;
assign v_6670 = v_6605 | v_6669;
assign v_6671 = v_6610 | v_6670;
assign v_6672 = v_6661 | v_6671;
assign v_6677 = v_6675 | v_6676;
assign v_6680 = v_6678 | v_6679;
assign v_6683 = v_6681 | v_6682;
assign v_6686 = v_6684 | v_6685;
assign v_6687 = ~v_6673 | v_6686;
assign v_6688 = v_6598 | ~v_6674;
assign v_6689 = ~v_91 | v_6582;
assign v_6691 = v_6600 | v_6690;
assign v_6692 = v_6163 | v_6585;
assign v_6694 = v_6605 | v_6693;
assign v_6695 = v_6590 | v_6603;
assign v_6697 = v_6610 | v_6696;
assign v_6698 = v_6595 | v_6608;
assign v_6700 = v_6673 | v_6699;
assign v_6707 = ~v_6701 | v_6706;
assign v_6708 = v_6598 | ~v_6702;
assign v_6709 = v_6600 | v_6708;
assign v_6710 = v_6605 | v_6709;
assign v_6711 = v_6610 | v_6710;
assign v_6712 = v_6701 | v_6711;
assign v_6714 = v_87 | v_6134;
assign v_6715 = v_89 | v_6714;
assign v_6716 = v_91 | v_6715;
assign v_6717 = ~v_91 | v_6418;
assign v_6719 = ~v_96 | v_6718;
assign v_6722 = ~v_807 | v_6136;
assign v_6724 = ~v_89 | v_6428;
assign v_6725 = v_91 | v_6724;
assign v_6726 = ~v_89 | v_6432;
assign v_6727 = v_91 | v_6726;
assign v_6729 = ~v_361 | v_6728;
assign v_6731 = ~v_89 | v_6439;
assign v_6732 = v_91 | v_6731;
assign v_6733 = ~v_89 | v_6443;
assign v_6734 = v_91 | v_6733;
assign v_6736 = ~v_563 | v_6735;
assign v_6738 = ~v_6713 | v_6737;
assign v_6743 = v_6741 | v_6742;
assign v_6745 = ~v_6720 | v_6744;
assign v_6747 = v_6745 | v_6746;
assign v_6752 = v_6749 | v_6751;
assign v_6754 = v_6747 | v_6753;
assign v_6759 = v_6756 | v_6758;
assign v_6761 = v_6754 | v_6760;
assign v_6762 = v_6713 | v_6761;
assign v_6769 = ~v_6763 | v_6768;
assign v_6770 = v_6744 | ~v_6764;
assign v_6771 = v_6746 | v_6770;
assign v_6772 = v_6753 | v_6771;
assign v_6773 = v_6760 | v_6772;
assign v_6774 = v_6763 | v_6773;
assign v_6781 = ~v_6775 | v_6780;
assign v_6782 = v_6744 | ~v_6776;
assign v_6783 = v_6746 | v_6782;
assign v_6784 = v_6753 | v_6783;
assign v_6785 = v_6760 | v_6784;
assign v_6786 = v_6775 | v_6785;
assign v_6793 = ~v_6787 | v_6792;
assign v_6794 = v_6744 | ~v_6788;
assign v_6795 = v_6746 | v_6794;
assign v_6796 = v_6753 | v_6795;
assign v_6797 = v_6760 | v_6796;
assign v_6798 = v_6787 | v_6797;
assign v_6805 = ~v_6799 | v_6804;
assign v_6806 = v_6744 | ~v_6800;
assign v_6807 = v_6746 | v_6806;
assign v_6808 = v_6753 | v_6807;
assign v_6809 = v_6760 | v_6808;
assign v_6810 = v_6799 | v_6809;
assign v_6817 = ~v_6811 | v_6816;
assign v_6818 = v_6744 | ~v_6812;
assign v_6819 = v_6746 | v_6818;
assign v_6820 = v_6753 | v_6819;
assign v_6821 = v_6760 | v_6820;
assign v_6822 = v_6811 | v_6821;
assign v_6825 = v_6744 | v_6824;
assign v_6826 = v_6719 | v_6742;
assign v_6828 = v_6746 | v_6827;
assign v_6829 = v_91 | v_6722;
assign v_6831 = v_6753 | v_6830;
assign v_6832 = v_6729 | v_6751;
assign v_6834 = v_6760 | v_6833;
assign v_6835 = v_6736 | v_6758;
assign v_6837 = ~v_6823 | v_6836;
assign v_6840 = v_6838 | v_6839;
assign v_6843 = v_6841 | v_6842;
assign v_6846 = v_6844 | v_6845;
assign v_6849 = v_6847 | v_6848;
assign v_6850 = v_6823 | v_6849;
assign v_6857 = ~v_6851 | v_6856;
assign v_6858 = v_6744 | ~v_6852;
assign v_6859 = v_6746 | v_6858;
assign v_6860 = v_6753 | v_6859;
assign v_6861 = v_6760 | v_6860;
assign v_6862 = v_6851 | v_6861;
assign v_6864 = ~v_96 | v_6715;
assign v_6867 = ~v_807 | v_6421;
assign v_6869 = ~v_91 | v_6724;
assign v_6870 = ~v_91 | v_6726;
assign v_6872 = ~v_361 | v_6871;
assign v_6874 = ~v_91 | v_6731;
assign v_6875 = ~v_91 | v_6733;
assign v_6877 = ~v_563 | v_6876;
assign v_6879 = ~v_6863 | v_6878;
assign v_6881 = ~v_6865 | v_6880;
assign v_6883 = v_6881 | v_6882;
assign v_6886 = v_6884 | v_6885;
assign v_6888 = v_6883 | v_6887;
assign v_6891 = v_6889 | v_6890;
assign v_6893 = v_6888 | v_6892;
assign v_6894 = v_6863 | v_6893;
assign v_6901 = ~v_6895 | v_6900;
assign v_6902 = v_6880 | ~v_6896;
assign v_6903 = v_6882 | v_6902;
assign v_6904 = v_6887 | v_6903;
assign v_6905 = v_6892 | v_6904;
assign v_6906 = v_6895 | v_6905;
assign v_6913 = ~v_6907 | v_6912;
assign v_6914 = v_6880 | ~v_6908;
assign v_6915 = v_6882 | v_6914;
assign v_6916 = v_6887 | v_6915;
assign v_6917 = v_6892 | v_6916;
assign v_6918 = v_6907 | v_6917;
assign v_6925 = ~v_6919 | v_6924;
assign v_6926 = v_6880 | ~v_6920;
assign v_6927 = v_6882 | v_6926;
assign v_6928 = v_6887 | v_6927;
assign v_6929 = v_6892 | v_6928;
assign v_6930 = v_6919 | v_6929;
assign v_6937 = ~v_6931 | v_6936;
assign v_6938 = v_6880 | ~v_6932;
assign v_6939 = v_6882 | v_6938;
assign v_6940 = v_6887 | v_6939;
assign v_6941 = v_6892 | v_6940;
assign v_6942 = v_6931 | v_6941;
assign v_6949 = ~v_6943 | v_6948;
assign v_6950 = v_6880 | ~v_6944;
assign v_6951 = v_6882 | v_6950;
assign v_6952 = v_6887 | v_6951;
assign v_6953 = v_6892 | v_6952;
assign v_6954 = v_6943 | v_6953;
assign v_6959 = v_6957 | v_6958;
assign v_6962 = v_6960 | v_6961;
assign v_6965 = v_6963 | v_6964;
assign v_6968 = v_6966 | v_6967;
assign v_6969 = ~v_6955 | v_6968;
assign v_6970 = v_6880 | ~v_6956;
assign v_6971 = ~v_91 | v_6864;
assign v_6973 = v_6882 | v_6972;
assign v_6974 = v_6451 | v_6867;
assign v_6976 = v_6887 | v_6975;
assign v_6977 = v_6872 | v_6885;
assign v_6979 = v_6892 | v_6978;
assign v_6980 = v_6877 | v_6890;
assign v_6982 = v_6955 | v_6981;
assign v_6989 = ~v_6983 | v_6988;
assign v_6990 = v_6880 | ~v_6984;
assign v_6991 = v_6882 | v_6990;
assign v_6992 = v_6887 | v_6991;
assign v_6993 = v_6892 | v_6992;
assign v_6994 = v_6983 | v_6993;
assign v_6996 = ~v_89 | v_6714;
assign v_6997 = v_91 | v_6996;
assign v_6998 = ~v_91 | v_6715;
assign v_7000 = ~v_96 | v_6999;
assign v_7003 = ~v_807 | v_6418;
assign v_7005 = v_87 | v_6427;
assign v_7006 = v_89 | v_7005;
assign v_7007 = v_91 | v_7006;
assign v_7008 = v_87 | v_6431;
assign v_7009 = v_89 | v_7008;
assign v_7010 = v_91 | v_7009;
assign v_7012 = ~v_361 | v_7011;
assign v_7014 = v_87 | v_6438;
assign v_7015 = v_89 | v_7014;
assign v_7016 = v_91 | v_7015;
assign v_7017 = v_87 | v_6442;
assign v_7018 = v_89 | v_7017;
assign v_7019 = v_91 | v_7018;
assign v_7021 = ~v_563 | v_7020;
assign v_7023 = ~v_6995 | v_7022;
assign v_7027 = v_7025 | v_7026;
assign v_7029 = ~v_7001 | v_7028;
assign v_7031 = v_7029 | v_7030;
assign v_7038 = v_7034 | v_7037;
assign v_7040 = v_7031 | v_7039;
assign v_7047 = v_7043 | v_7046;
assign v_7049 = v_7040 | v_7048;
assign v_7050 = v_6995 | v_7049;
assign v_7057 = ~v_7051 | v_7056;
assign v_7058 = v_7028 | ~v_7052;
assign v_7059 = v_7030 | v_7058;
assign v_7060 = v_7039 | v_7059;
assign v_7061 = v_7048 | v_7060;
assign v_7062 = v_7051 | v_7061;
assign v_7069 = ~v_7063 | v_7068;
assign v_7070 = v_7028 | ~v_7064;
assign v_7071 = v_7030 | v_7070;
assign v_7072 = v_7039 | v_7071;
assign v_7073 = v_7048 | v_7072;
assign v_7074 = v_7063 | v_7073;
assign v_7081 = ~v_7075 | v_7080;
assign v_7082 = v_7028 | ~v_7076;
assign v_7083 = v_7030 | v_7082;
assign v_7084 = v_7039 | v_7083;
assign v_7085 = v_7048 | v_7084;
assign v_7086 = v_7075 | v_7085;
assign v_7093 = ~v_7087 | v_7092;
assign v_7094 = v_7028 | ~v_7088;
assign v_7095 = v_7030 | v_7094;
assign v_7096 = v_7039 | v_7095;
assign v_7097 = v_7048 | v_7096;
assign v_7098 = v_7087 | v_7097;
assign v_7105 = ~v_7099 | v_7104;
assign v_7106 = v_7028 | ~v_7100;
assign v_7107 = v_7030 | v_7106;
assign v_7108 = v_7039 | v_7107;
assign v_7109 = v_7048 | v_7108;
assign v_7110 = v_7099 | v_7109;
assign v_7115 = v_7113 | v_7114;
assign v_7118 = v_7116 | v_7117;
assign v_7121 = v_7119 | v_7120;
assign v_7124 = v_7122 | v_7123;
assign v_7125 = ~v_7111 | v_7124;
assign v_7126 = v_7028 | ~v_7112;
assign v_7127 = v_7000 | v_7026;
assign v_7129 = v_7030 | v_7128;
assign v_7130 = v_91 | v_7003;
assign v_7132 = v_7039 | v_7131;
assign v_7133 = v_7012 | v_7037;
assign v_7135 = v_7048 | v_7134;
assign v_7136 = v_7021 | v_7046;
assign v_7138 = v_7111 | v_7137;
assign v_7141 = v_7028 | v_7140;
assign v_7142 = v_7030 | v_7141;
assign v_7143 = v_7039 | v_7142;
assign v_7144 = v_7048 | v_7143;
assign v_7145 = ~v_7139 | v_7144;
assign v_7150 = v_7139 | v_7149;
assign v_7152 = ~v_96 | v_6996;
assign v_7155 = ~v_807 | v_6718;
assign v_7157 = ~v_91 | v_7006;
assign v_7158 = ~v_91 | v_7009;
assign v_7160 = ~v_361 | v_7159;
assign v_7162 = ~v_91 | v_7015;
assign v_7163 = ~v_91 | v_7018;
assign v_7165 = ~v_563 | v_7164;
assign v_7167 = ~v_7151 | v_7166;
assign v_7169 = ~v_7153 | v_7168;
assign v_7171 = v_7169 | v_7170;
assign v_7174 = v_7172 | v_7173;
assign v_7176 = v_7171 | v_7175;
assign v_7179 = v_7177 | v_7178;
assign v_7181 = v_7176 | v_7180;
assign v_7182 = v_7151 | v_7181;
assign v_7189 = ~v_7183 | v_7188;
assign v_7190 = v_7168 | ~v_7184;
assign v_7191 = v_7170 | v_7190;
assign v_7192 = v_7175 | v_7191;
assign v_7193 = v_7180 | v_7192;
assign v_7194 = v_7183 | v_7193;
assign v_7201 = ~v_7195 | v_7200;
assign v_7202 = v_7168 | ~v_7196;
assign v_7203 = v_7170 | v_7202;
assign v_7204 = v_7175 | v_7203;
assign v_7205 = v_7180 | v_7204;
assign v_7206 = v_7195 | v_7205;
assign v_7213 = ~v_7207 | v_7212;
assign v_7214 = v_7168 | ~v_7208;
assign v_7215 = v_7170 | v_7214;
assign v_7216 = v_7175 | v_7215;
assign v_7217 = v_7180 | v_7216;
assign v_7218 = v_7207 | v_7217;
assign v_7225 = ~v_7219 | v_7224;
assign v_7226 = v_7168 | ~v_7220;
assign v_7227 = v_7170 | v_7226;
assign v_7228 = v_7175 | v_7227;
assign v_7229 = v_7180 | v_7228;
assign v_7230 = v_7219 | v_7229;
assign v_7237 = ~v_7231 | v_7236;
assign v_7238 = v_7168 | ~v_7232;
assign v_7239 = v_7170 | v_7238;
assign v_7240 = v_7175 | v_7239;
assign v_7241 = v_7180 | v_7240;
assign v_7242 = v_7231 | v_7241;
assign v_7247 = v_7245 | v_7246;
assign v_7250 = v_7248 | v_7249;
assign v_7253 = v_7251 | v_7252;
assign v_7256 = v_7254 | v_7255;
assign v_7257 = ~v_7243 | v_7256;
assign v_7258 = v_7168 | ~v_7244;
assign v_7259 = ~v_91 | v_7152;
assign v_7261 = v_7170 | v_7260;
assign v_7262 = v_6741 | v_7155;
assign v_7264 = v_7175 | v_7263;
assign v_7265 = v_7160 | v_7173;
assign v_7267 = v_7180 | v_7266;
assign v_7268 = v_7165 | v_7178;
assign v_7270 = v_7243 | v_7269;
assign v_7277 = ~v_7271 | v_7276;
assign v_7278 = v_7168 | ~v_7272;
assign v_7279 = v_7170 | v_7278;
assign v_7280 = v_7175 | v_7279;
assign v_7281 = v_7180 | v_7280;
assign v_7282 = v_7271 | v_7281;
assign v_7284 = v_584 | v_4964;
assign v_7285 = v_85 | v_7284;
assign v_7286 = ~v_87 | v_7285;
assign v_7287 = v_89 | v_7286;
assign v_7288 = v_91 | v_7287;
assign v_7289 = ~v_91 | v_6996;
assign v_7291 = ~v_96 | v_7290;
assign v_7294 = ~v_807 | v_6715;
assign v_7296 = ~v_89 | v_7005;
assign v_7297 = v_91 | v_7296;
assign v_7298 = ~v_89 | v_7008;
assign v_7299 = v_91 | v_7298;
assign v_7301 = ~v_361 | v_7300;
assign v_7303 = ~v_89 | v_7014;
assign v_7304 = v_91 | v_7303;
assign v_7305 = ~v_89 | v_7017;
assign v_7306 = v_91 | v_7305;
assign v_7308 = ~v_563 | v_7307;
assign v_7310 = ~v_7283 | v_7309;
assign v_7317 = v_7315 | v_7316;
assign v_7319 = ~v_7292 | v_7318;
assign v_7321 = v_7319 | v_7320;
assign v_7326 = v_7323 | v_7325;
assign v_7328 = v_7321 | v_7327;
assign v_7333 = v_7330 | v_7332;
assign v_7335 = v_7328 | v_7334;
assign v_7336 = v_7283 | v_7335;
assign v_7343 = ~v_7337 | v_7342;
assign v_7344 = v_7318 | ~v_7338;
assign v_7345 = v_7320 | v_7344;
assign v_7346 = v_7327 | v_7345;
assign v_7347 = v_7334 | v_7346;
assign v_7348 = v_7337 | v_7347;
assign v_7355 = ~v_7349 | v_7354;
assign v_7356 = v_7318 | ~v_7350;
assign v_7357 = v_7320 | v_7356;
assign v_7358 = v_7327 | v_7357;
assign v_7359 = v_7334 | v_7358;
assign v_7360 = v_7349 | v_7359;
assign v_7367 = ~v_7361 | v_7366;
assign v_7368 = v_7318 | ~v_7362;
assign v_7369 = v_7320 | v_7368;
assign v_7370 = v_7327 | v_7369;
assign v_7371 = v_7334 | v_7370;
assign v_7372 = v_7361 | v_7371;
assign v_7379 = ~v_7373 | v_7378;
assign v_7380 = v_7318 | ~v_7374;
assign v_7381 = v_7320 | v_7380;
assign v_7382 = v_7327 | v_7381;
assign v_7383 = v_7334 | v_7382;
assign v_7384 = v_7373 | v_7383;
assign v_7391 = ~v_7385 | v_7390;
assign v_7392 = v_7318 | ~v_7386;
assign v_7393 = v_7320 | v_7392;
assign v_7394 = v_7327 | v_7393;
assign v_7395 = v_7334 | v_7394;
assign v_7396 = v_7385 | v_7395;
assign v_7401 = v_7399 | v_7400;
assign v_7404 = v_7402 | v_7403;
assign v_7407 = v_7405 | v_7406;
assign v_7410 = v_7408 | v_7409;
assign v_7411 = ~v_7397 | v_7410;
assign v_7412 = v_7318 | ~v_7398;
assign v_7413 = v_7291 | v_7316;
assign v_7415 = v_7320 | v_7414;
assign v_7416 = v_91 | v_7294;
assign v_7418 = v_7327 | v_7417;
assign v_7419 = v_7301 | v_7325;
assign v_7421 = v_7334 | v_7420;
assign v_7422 = v_7308 | v_7332;
assign v_7424 = v_7397 | v_7423;
assign v_7427 = v_7318 | v_7426;
assign v_7428 = v_7320 | v_7427;
assign v_7429 = v_7327 | v_7428;
assign v_7430 = v_7334 | v_7429;
assign v_7431 = ~v_7425 | v_7430;
assign v_7436 = v_7425 | v_7435;
assign v_7438 = ~v_96 | v_7287;
assign v_7441 = ~v_807 | v_6999;
assign v_7443 = ~v_91 | v_7296;
assign v_7444 = ~v_91 | v_7298;
assign v_7446 = ~v_361 | v_7445;
assign v_7448 = ~v_91 | v_7303;
assign v_7449 = ~v_91 | v_7305;
assign v_7451 = ~v_563 | v_7450;
assign v_7453 = ~v_7437 | v_7452;
assign v_7455 = ~v_7439 | v_7454;
assign v_7457 = v_7455 | v_7456;
assign v_7460 = v_7458 | v_7459;
assign v_7462 = v_7457 | v_7461;
assign v_7465 = v_7463 | v_7464;
assign v_7467 = v_7462 | v_7466;
assign v_7468 = v_7437 | v_7467;
assign v_7475 = ~v_7469 | v_7474;
assign v_7476 = v_7454 | ~v_7470;
assign v_7477 = v_7456 | v_7476;
assign v_7478 = v_7461 | v_7477;
assign v_7479 = v_7466 | v_7478;
assign v_7480 = v_7469 | v_7479;
assign v_7487 = ~v_7481 | v_7486;
assign v_7488 = v_7454 | ~v_7482;
assign v_7489 = v_7456 | v_7488;
assign v_7490 = v_7461 | v_7489;
assign v_7491 = v_7466 | v_7490;
assign v_7492 = v_7481 | v_7491;
assign v_7499 = ~v_7493 | v_7498;
assign v_7500 = v_7454 | ~v_7494;
assign v_7501 = v_7456 | v_7500;
assign v_7502 = v_7461 | v_7501;
assign v_7503 = v_7466 | v_7502;
assign v_7504 = v_7493 | v_7503;
assign v_7511 = ~v_7505 | v_7510;
assign v_7512 = v_7454 | ~v_7506;
assign v_7513 = v_7456 | v_7512;
assign v_7514 = v_7461 | v_7513;
assign v_7515 = v_7466 | v_7514;
assign v_7516 = v_7505 | v_7515;
assign v_7523 = ~v_7517 | v_7522;
assign v_7524 = v_7454 | ~v_7518;
assign v_7525 = v_7456 | v_7524;
assign v_7526 = v_7461 | v_7525;
assign v_7527 = v_7466 | v_7526;
assign v_7528 = v_7517 | v_7527;
assign v_7533 = v_7531 | v_7532;
assign v_7536 = v_7534 | v_7535;
assign v_7539 = v_7537 | v_7538;
assign v_7542 = v_7540 | v_7541;
assign v_7543 = ~v_7529 | v_7542;
assign v_7544 = v_7454 | ~v_7530;
assign v_7545 = ~v_91 | v_7438;
assign v_7547 = v_7456 | v_7546;
assign v_7548 = v_7025 | v_7441;
assign v_7550 = v_7461 | v_7549;
assign v_7551 = v_7446 | v_7459;
assign v_7553 = v_7466 | v_7552;
assign v_7554 = v_7451 | v_7464;
assign v_7556 = v_7529 | v_7555;
assign v_7559 = v_7454 | v_7558;
assign v_7560 = v_7456 | v_7559;
assign v_7561 = v_7461 | v_7560;
assign v_7562 = v_7466 | v_7561;
assign v_7563 = ~v_7557 | v_7562;
assign v_7568 = v_7557 | v_7567;
assign v_7570 = ~v_89 | v_7286;
assign v_7571 = v_91 | v_7570;
assign v_7572 = ~v_91 | v_7287;
assign v_7574 = ~v_96 | v_7573;
assign v_7577 = ~v_807 | v_6996;
assign v_7579 = v_621 | v_5261;
assign v_7580 = v_85 | v_7579;
assign v_7581 = ~v_87 | v_7580;
assign v_7582 = v_89 | v_7581;
assign v_7583 = v_91 | v_7582;
assign v_7584 = v_651 | v_5267;
assign v_7585 = v_355 | v_7584;
assign v_7586 = ~v_87 | v_7585;
assign v_7587 = v_89 | v_7586;
assign v_7588 = v_91 | v_7587;
assign v_7590 = ~v_361 | v_7589;
assign v_7592 = v_621 | v_5276;
assign v_7593 = v_85 | v_7592;
assign v_7594 = ~v_87 | v_7593;
assign v_7595 = v_89 | v_7594;
assign v_7596 = v_91 | v_7595;
assign v_7597 = v_710 | v_5282;
assign v_7598 = v_355 | v_7597;
assign v_7599 = ~v_87 | v_7598;
assign v_7600 = v_89 | v_7599;
assign v_7601 = v_91 | v_7600;
assign v_7603 = ~v_563 | v_7602;
assign v_7605 = ~v_7569 | v_7604;
assign v_7609 = v_7607 | v_7608;
assign v_7611 = ~v_7575 | v_7610;
assign v_7613 = v_7611 | v_7612;
assign v_7624 = v_7618 | v_7623;
assign v_7626 = v_7613 | v_7625;
assign v_7637 = v_7631 | v_7636;
assign v_7639 = v_7626 | v_7638;
assign v_7640 = v_7569 | v_7639;
assign v_7647 = ~v_7641 | v_7646;
assign v_7648 = v_7610 | ~v_7642;
assign v_7649 = v_7612 | v_7648;
assign v_7650 = v_7625 | v_7649;
assign v_7651 = v_7638 | v_7650;
assign v_7652 = v_7641 | v_7651;
assign v_7659 = ~v_7653 | v_7658;
assign v_7660 = v_7610 | ~v_7654;
assign v_7661 = v_7612 | v_7660;
assign v_7662 = v_7625 | v_7661;
assign v_7663 = v_7638 | v_7662;
assign v_7664 = v_7653 | v_7663;
assign v_7671 = ~v_7665 | v_7670;
assign v_7672 = v_7610 | ~v_7666;
assign v_7673 = v_7612 | v_7672;
assign v_7674 = v_7625 | v_7673;
assign v_7675 = v_7638 | v_7674;
assign v_7676 = v_7665 | v_7675;
assign v_7683 = ~v_7677 | v_7682;
assign v_7684 = v_7610 | ~v_7678;
assign v_7685 = v_7612 | v_7684;
assign v_7686 = v_7625 | v_7685;
assign v_7687 = v_7638 | v_7686;
assign v_7688 = v_7677 | v_7687;
assign v_7695 = ~v_7689 | v_7694;
assign v_7696 = v_7610 | ~v_7690;
assign v_7697 = v_7612 | v_7696;
assign v_7698 = v_7625 | v_7697;
assign v_7699 = v_7638 | v_7698;
assign v_7700 = v_7689 | v_7699;
assign v_7705 = v_7703 | v_7704;
assign v_7708 = v_7706 | v_7707;
assign v_7711 = v_7709 | v_7710;
assign v_7714 = v_7712 | v_7713;
assign v_7715 = ~v_7701 | v_7714;
assign v_7716 = v_7610 | ~v_7702;
assign v_7717 = v_7574 | v_7608;
assign v_7719 = v_7612 | v_7718;
assign v_7720 = v_91 | v_7577;
assign v_7722 = v_7625 | v_7721;
assign v_7723 = v_7590 | v_7623;
assign v_7725 = v_7638 | v_7724;
assign v_7726 = v_7603 | v_7636;
assign v_7728 = v_7701 | v_7727;
assign v_7731 = v_7610 | v_7730;
assign v_7732 = v_7612 | v_7731;
assign v_7733 = v_7625 | v_7732;
assign v_7734 = v_7638 | v_7733;
assign v_7735 = ~v_7729 | v_7734;
assign v_7740 = v_7729 | v_7739;
assign v_7742 = ~v_96 | v_7570;
assign v_7745 = ~v_807 | v_7290;
assign v_7747 = ~v_91 | v_7582;
assign v_7748 = ~v_91 | v_7587;
assign v_7750 = ~v_361 | v_7749;
assign v_7752 = ~v_91 | v_7595;
assign v_7753 = ~v_91 | v_7600;
assign v_7755 = ~v_563 | v_7754;
assign v_7757 = ~v_7741 | v_7756;
assign v_7759 = ~v_7743 | v_7758;
assign v_7761 = v_7759 | v_7760;
assign v_7764 = v_7762 | v_7763;
assign v_7766 = v_7761 | v_7765;
assign v_7769 = v_7767 | v_7768;
assign v_7771 = v_7766 | v_7770;
assign v_7772 = v_7741 | v_7771;
assign v_7779 = ~v_7773 | v_7778;
assign v_7780 = v_7758 | ~v_7774;
assign v_7781 = v_7760 | v_7780;
assign v_7782 = v_7765 | v_7781;
assign v_7783 = v_7770 | v_7782;
assign v_7784 = v_7773 | v_7783;
assign v_7791 = ~v_7785 | v_7790;
assign v_7792 = v_7758 | ~v_7786;
assign v_7793 = v_7760 | v_7792;
assign v_7794 = v_7765 | v_7793;
assign v_7795 = v_7770 | v_7794;
assign v_7796 = v_7785 | v_7795;
assign v_7803 = ~v_7797 | v_7802;
assign v_7804 = v_7758 | ~v_7798;
assign v_7805 = v_7760 | v_7804;
assign v_7806 = v_7765 | v_7805;
assign v_7807 = v_7770 | v_7806;
assign v_7808 = v_7797 | v_7807;
assign v_7815 = ~v_7809 | v_7814;
assign v_7816 = v_7758 | ~v_7810;
assign v_7817 = v_7760 | v_7816;
assign v_7818 = v_7765 | v_7817;
assign v_7819 = v_7770 | v_7818;
assign v_7820 = v_7809 | v_7819;
assign v_7827 = ~v_7821 | v_7826;
assign v_7828 = v_7758 | ~v_7822;
assign v_7829 = v_7760 | v_7828;
assign v_7830 = v_7765 | v_7829;
assign v_7831 = v_7770 | v_7830;
assign v_7832 = v_7821 | v_7831;
assign v_7837 = v_7835 | v_7836;
assign v_7840 = v_7838 | v_7839;
assign v_7843 = v_7841 | v_7842;
assign v_7846 = v_7844 | v_7845;
assign v_7847 = ~v_7833 | v_7846;
assign v_7848 = v_7758 | ~v_7834;
assign v_7849 = ~v_91 | v_7742;
assign v_7851 = v_7760 | v_7850;
assign v_7852 = v_7315 | v_7745;
assign v_7854 = v_7765 | v_7853;
assign v_7855 = v_7750 | v_7763;
assign v_7857 = v_7770 | v_7856;
assign v_7858 = v_7755 | v_7768;
assign v_7860 = v_7833 | v_7859;
assign v_7863 = v_7758 | v_7862;
assign v_7864 = v_7760 | v_7863;
assign v_7865 = v_7765 | v_7864;
assign v_7866 = v_7770 | v_7865;
assign v_7867 = ~v_7861 | v_7866;
assign v_7872 = v_7861 | v_7871;
assign v_7874 = v_87 | v_7285;
assign v_7875 = v_89 | v_7874;
assign v_7876 = v_91 | v_7875;
assign v_7877 = ~v_91 | v_7570;
assign v_7879 = ~v_96 | v_7878;
assign v_7882 = ~v_807 | v_7287;
assign v_7884 = ~v_89 | v_7581;
assign v_7885 = v_91 | v_7884;
assign v_7886 = ~v_89 | v_7586;
assign v_7887 = v_91 | v_7886;
assign v_7889 = ~v_361 | v_7888;
assign v_7891 = ~v_89 | v_7594;
assign v_7892 = v_91 | v_7891;
assign v_7893 = ~v_89 | v_7599;
assign v_7894 = v_91 | v_7893;
assign v_7896 = ~v_563 | v_7895;
assign v_7898 = ~v_7873 | v_7897;
assign v_7903 = v_7901 | v_7902;
assign v_7905 = ~v_7880 | v_7904;
assign v_7907 = v_7905 | v_7906;
assign v_7912 = v_7909 | v_7911;
assign v_7914 = v_7907 | v_7913;
assign v_7919 = v_7916 | v_7918;
assign v_7921 = v_7914 | v_7920;
assign v_7922 = v_7873 | v_7921;
assign v_7929 = ~v_7923 | v_7928;
assign v_7930 = v_7904 | ~v_7924;
assign v_7931 = v_7906 | v_7930;
assign v_7932 = v_7913 | v_7931;
assign v_7933 = v_7920 | v_7932;
assign v_7934 = v_7923 | v_7933;
assign v_7941 = ~v_7935 | v_7940;
assign v_7942 = v_7904 | ~v_7936;
assign v_7943 = v_7906 | v_7942;
assign v_7944 = v_7913 | v_7943;
assign v_7945 = v_7920 | v_7944;
assign v_7946 = v_7935 | v_7945;
assign v_7953 = ~v_7947 | v_7952;
assign v_7954 = v_7904 | ~v_7948;
assign v_7955 = v_7906 | v_7954;
assign v_7956 = v_7913 | v_7955;
assign v_7957 = v_7920 | v_7956;
assign v_7958 = v_7947 | v_7957;
assign v_7965 = ~v_7959 | v_7964;
assign v_7966 = v_7904 | ~v_7960;
assign v_7967 = v_7906 | v_7966;
assign v_7968 = v_7913 | v_7967;
assign v_7969 = v_7920 | v_7968;
assign v_7970 = v_7959 | v_7969;
assign v_7977 = ~v_7971 | v_7976;
assign v_7978 = v_7904 | ~v_7972;
assign v_7979 = v_7906 | v_7978;
assign v_7980 = v_7913 | v_7979;
assign v_7981 = v_7920 | v_7980;
assign v_7982 = v_7971 | v_7981;
assign v_7987 = v_7985 | v_7986;
assign v_7990 = v_7988 | v_7989;
assign v_7993 = v_7991 | v_7992;
assign v_7996 = v_7994 | v_7995;
assign v_7997 = ~v_7983 | v_7996;
assign v_7998 = v_7904 | ~v_7984;
assign v_7999 = v_7879 | v_7902;
assign v_8001 = v_7906 | v_8000;
assign v_8002 = v_91 | v_7882;
assign v_8004 = v_7913 | v_8003;
assign v_8005 = v_7889 | v_7911;
assign v_8007 = v_7920 | v_8006;
assign v_8008 = v_7896 | v_7918;
assign v_8010 = v_7983 | v_8009;
assign v_8013 = v_7904 | v_8012;
assign v_8014 = v_7906 | v_8013;
assign v_8015 = v_7913 | v_8014;
assign v_8016 = v_7920 | v_8015;
assign v_8017 = ~v_8011 | v_8016;
assign v_8022 = v_8011 | v_8021;
assign v_8024 = ~v_96 | v_7875;
assign v_8027 = ~v_807 | v_7573;
assign v_8029 = ~v_91 | v_7884;
assign v_8030 = ~v_91 | v_7886;
assign v_8032 = ~v_361 | v_8031;
assign v_8034 = ~v_91 | v_7891;
assign v_8035 = ~v_91 | v_7893;
assign v_8037 = ~v_563 | v_8036;
assign v_8039 = ~v_8023 | v_8038;
assign v_8041 = ~v_8025 | v_8040;
assign v_8043 = v_8041 | v_8042;
assign v_8046 = v_8044 | v_8045;
assign v_8048 = v_8043 | v_8047;
assign v_8051 = v_8049 | v_8050;
assign v_8053 = v_8048 | v_8052;
assign v_8054 = v_8023 | v_8053;
assign v_8061 = ~v_8055 | v_8060;
assign v_8062 = v_8040 | ~v_8056;
assign v_8063 = v_8042 | v_8062;
assign v_8064 = v_8047 | v_8063;
assign v_8065 = v_8052 | v_8064;
assign v_8066 = v_8055 | v_8065;
assign v_8073 = ~v_8067 | v_8072;
assign v_8074 = v_8040 | ~v_8068;
assign v_8075 = v_8042 | v_8074;
assign v_8076 = v_8047 | v_8075;
assign v_8077 = v_8052 | v_8076;
assign v_8078 = v_8067 | v_8077;
assign v_8085 = ~v_8079 | v_8084;
assign v_8086 = v_8040 | ~v_8080;
assign v_8087 = v_8042 | v_8086;
assign v_8088 = v_8047 | v_8087;
assign v_8089 = v_8052 | v_8088;
assign v_8090 = v_8079 | v_8089;
assign v_8097 = ~v_8091 | v_8096;
assign v_8098 = v_8040 | ~v_8092;
assign v_8099 = v_8042 | v_8098;
assign v_8100 = v_8047 | v_8099;
assign v_8101 = v_8052 | v_8100;
assign v_8102 = v_8091 | v_8101;
assign v_8109 = ~v_8103 | v_8108;
assign v_8110 = v_8040 | ~v_8104;
assign v_8111 = v_8042 | v_8110;
assign v_8112 = v_8047 | v_8111;
assign v_8113 = v_8052 | v_8112;
assign v_8114 = v_8103 | v_8113;
assign v_8119 = v_8117 | v_8118;
assign v_8122 = v_8120 | v_8121;
assign v_8125 = v_8123 | v_8124;
assign v_8128 = v_8126 | v_8127;
assign v_8129 = ~v_8115 | v_8128;
assign v_8130 = v_8040 | ~v_8116;
assign v_8131 = ~v_91 | v_8024;
assign v_8133 = v_8042 | v_8132;
assign v_8134 = v_7607 | v_8027;
assign v_8136 = v_8047 | v_8135;
assign v_8137 = v_8032 | v_8045;
assign v_8139 = v_8052 | v_8138;
assign v_8140 = v_8037 | v_8050;
assign v_8142 = v_8115 | v_8141;
assign v_8149 = ~v_8143 | v_8148;
assign v_8150 = v_8040 | ~v_8144;
assign v_8151 = v_8042 | v_8150;
assign v_8152 = v_8047 | v_8151;
assign v_8153 = v_8052 | v_8152;
assign v_8154 = v_8143 | v_8153;
assign v_8156 = ~v_89 | v_7874;
assign v_8157 = v_91 | v_8156;
assign v_8158 = ~v_91 | v_7875;
assign v_8160 = ~v_96 | v_8159;
assign v_8163 = ~v_807 | v_7570;
assign v_8165 = v_87 | v_7580;
assign v_8166 = v_89 | v_8165;
assign v_8167 = v_91 | v_8166;
assign v_8168 = v_87 | v_7585;
assign v_8169 = v_89 | v_8168;
assign v_8170 = v_91 | v_8169;
assign v_8172 = ~v_361 | v_8171;
assign v_8174 = v_87 | v_7593;
assign v_8175 = v_89 | v_8174;
assign v_8176 = v_91 | v_8175;
assign v_8177 = v_87 | v_7598;
assign v_8178 = v_89 | v_8177;
assign v_8179 = v_91 | v_8178;
assign v_8181 = ~v_563 | v_8180;
assign v_8183 = ~v_8155 | v_8182;
assign v_8187 = v_8185 | v_8186;
assign v_8189 = ~v_8161 | v_8188;
assign v_8191 = v_8189 | v_8190;
assign v_8198 = v_8194 | v_8197;
assign v_8200 = v_8191 | v_8199;
assign v_8207 = v_8203 | v_8206;
assign v_8209 = v_8200 | v_8208;
assign v_8210 = v_8155 | v_8209;
assign v_8217 = ~v_8211 | v_8216;
assign v_8218 = v_8188 | ~v_8212;
assign v_8219 = v_8190 | v_8218;
assign v_8220 = v_8199 | v_8219;
assign v_8221 = v_8208 | v_8220;
assign v_8222 = v_8211 | v_8221;
assign v_8229 = ~v_8223 | v_8228;
assign v_8230 = v_8188 | ~v_8224;
assign v_8231 = v_8190 | v_8230;
assign v_8232 = v_8199 | v_8231;
assign v_8233 = v_8208 | v_8232;
assign v_8234 = v_8223 | v_8233;
assign v_8241 = ~v_8235 | v_8240;
assign v_8242 = v_8188 | ~v_8236;
assign v_8243 = v_8190 | v_8242;
assign v_8244 = v_8199 | v_8243;
assign v_8245 = v_8208 | v_8244;
assign v_8246 = v_8235 | v_8245;
assign v_8253 = ~v_8247 | v_8252;
assign v_8254 = v_8188 | ~v_8248;
assign v_8255 = v_8190 | v_8254;
assign v_8256 = v_8199 | v_8255;
assign v_8257 = v_8208 | v_8256;
assign v_8258 = v_8247 | v_8257;
assign v_8265 = ~v_8259 | v_8264;
assign v_8266 = v_8188 | ~v_8260;
assign v_8267 = v_8190 | v_8266;
assign v_8268 = v_8199 | v_8267;
assign v_8269 = v_8208 | v_8268;
assign v_8270 = v_8259 | v_8269;
assign v_8275 = v_8273 | v_8274;
assign v_8278 = v_8276 | v_8277;
assign v_8281 = v_8279 | v_8280;
assign v_8284 = v_8282 | v_8283;
assign v_8285 = ~v_8271 | v_8284;
assign v_8286 = v_8188 | ~v_8272;
assign v_8287 = v_8160 | v_8186;
assign v_8289 = v_8190 | v_8288;
assign v_8290 = v_91 | v_8163;
assign v_8292 = v_8199 | v_8291;
assign v_8293 = v_8172 | v_8197;
assign v_8295 = v_8208 | v_8294;
assign v_8296 = v_8181 | v_8206;
assign v_8298 = v_8271 | v_8297;
assign v_8305 = ~v_8299 | v_8304;
assign v_8306 = v_8188 | ~v_8300;
assign v_8307 = v_8190 | v_8306;
assign v_8308 = v_8199 | v_8307;
assign v_8309 = v_8208 | v_8308;
assign v_8310 = v_8299 | v_8309;
assign v_8312 = ~v_96 | v_8156;
assign v_8315 = ~v_807 | v_7878;
assign v_8317 = ~v_91 | v_8166;
assign v_8318 = ~v_91 | v_8169;
assign v_8320 = ~v_361 | v_8319;
assign v_8322 = ~v_91 | v_8175;
assign v_8323 = ~v_91 | v_8178;
assign v_8325 = ~v_563 | v_8324;
assign v_8327 = ~v_8311 | v_8326;
assign v_8329 = ~v_8313 | v_8328;
assign v_8331 = v_8329 | v_8330;
assign v_8334 = v_8332 | v_8333;
assign v_8336 = v_8331 | v_8335;
assign v_8339 = v_8337 | v_8338;
assign v_8341 = v_8336 | v_8340;
assign v_8342 = v_8311 | v_8341;
assign v_8349 = ~v_8343 | v_8348;
assign v_8350 = v_8328 | ~v_8344;
assign v_8351 = v_8330 | v_8350;
assign v_8352 = v_8335 | v_8351;
assign v_8353 = v_8340 | v_8352;
assign v_8354 = v_8343 | v_8353;
assign v_8361 = ~v_8355 | v_8360;
assign v_8362 = v_8328 | ~v_8356;
assign v_8363 = v_8330 | v_8362;
assign v_8364 = v_8335 | v_8363;
assign v_8365 = v_8340 | v_8364;
assign v_8366 = v_8355 | v_8365;
assign v_8373 = ~v_8367 | v_8372;
assign v_8374 = v_8328 | ~v_8368;
assign v_8375 = v_8330 | v_8374;
assign v_8376 = v_8335 | v_8375;
assign v_8377 = v_8340 | v_8376;
assign v_8378 = v_8367 | v_8377;
assign v_8385 = ~v_8379 | v_8384;
assign v_8386 = v_8328 | ~v_8380;
assign v_8387 = v_8330 | v_8386;
assign v_8388 = v_8335 | v_8387;
assign v_8389 = v_8340 | v_8388;
assign v_8390 = v_8379 | v_8389;
assign v_8397 = ~v_8391 | v_8396;
assign v_8398 = v_8328 | ~v_8392;
assign v_8399 = v_8330 | v_8398;
assign v_8400 = v_8335 | v_8399;
assign v_8401 = v_8340 | v_8400;
assign v_8402 = v_8391 | v_8401;
assign v_8407 = v_8405 | v_8406;
assign v_8410 = v_8408 | v_8409;
assign v_8413 = v_8411 | v_8412;
assign v_8416 = v_8414 | v_8415;
assign v_8417 = ~v_8403 | v_8416;
assign v_8418 = v_8328 | ~v_8404;
assign v_8419 = ~v_91 | v_8312;
assign v_8421 = v_8330 | v_8420;
assign v_8422 = v_7901 | v_8315;
assign v_8424 = v_8335 | v_8423;
assign v_8425 = v_8320 | v_8333;
assign v_8427 = v_8340 | v_8426;
assign v_8428 = v_8325 | v_8338;
assign v_8430 = v_8403 | v_8429;
assign v_8437 = ~v_8431 | v_8436;
assign v_8438 = v_8328 | ~v_8432;
assign v_8439 = v_8330 | v_8438;
assign v_8440 = v_8335 | v_8439;
assign v_8441 = v_8340 | v_8440;
assign v_8442 = v_8431 | v_8441;
assign v_8444 = v_587 | v_7284;
assign v_8445 = ~v_87 | v_8444;
assign v_8446 = v_89 | v_8445;
assign v_8447 = v_91 | v_8446;
assign v_8448 = ~v_91 | v_8156;
assign v_8450 = ~v_96 | v_8449;
assign v_8453 = ~v_807 | v_7875;
assign v_8455 = ~v_89 | v_8165;
assign v_8456 = v_91 | v_8455;
assign v_8457 = ~v_89 | v_8168;
assign v_8458 = v_91 | v_8457;
assign v_8460 = ~v_361 | v_8459;
assign v_8462 = ~v_89 | v_8174;
assign v_8463 = v_91 | v_8462;
assign v_8464 = ~v_89 | v_8177;
assign v_8465 = v_91 | v_8464;
assign v_8467 = ~v_563 | v_8466;
assign v_8469 = ~v_8443 | v_8468;
assign v_8475 = v_8473 | v_8474;
assign v_8477 = ~v_8451 | v_8476;
assign v_8479 = v_8477 | v_8478;
assign v_8484 = v_8481 | v_8483;
assign v_8486 = v_8479 | v_8485;
assign v_8491 = v_8488 | v_8490;
assign v_8493 = v_8486 | v_8492;
assign v_8494 = v_8443 | v_8493;
assign v_8501 = ~v_8495 | v_8500;
assign v_8502 = v_8476 | ~v_8496;
assign v_8503 = v_8478 | v_8502;
assign v_8504 = v_8485 | v_8503;
assign v_8505 = v_8492 | v_8504;
assign v_8506 = v_8495 | v_8505;
assign v_8513 = ~v_8507 | v_8512;
assign v_8514 = v_8476 | ~v_8508;
assign v_8515 = v_8478 | v_8514;
assign v_8516 = v_8485 | v_8515;
assign v_8517 = v_8492 | v_8516;
assign v_8518 = v_8507 | v_8517;
assign v_8525 = ~v_8519 | v_8524;
assign v_8526 = v_8476 | ~v_8520;
assign v_8527 = v_8478 | v_8526;
assign v_8528 = v_8485 | v_8527;
assign v_8529 = v_8492 | v_8528;
assign v_8530 = v_8519 | v_8529;
assign v_8537 = ~v_8531 | v_8536;
assign v_8538 = v_8476 | ~v_8532;
assign v_8539 = v_8478 | v_8538;
assign v_8540 = v_8485 | v_8539;
assign v_8541 = v_8492 | v_8540;
assign v_8542 = v_8531 | v_8541;
assign v_8549 = ~v_8543 | v_8548;
assign v_8550 = v_8476 | ~v_8544;
assign v_8551 = v_8478 | v_8550;
assign v_8552 = v_8485 | v_8551;
assign v_8553 = v_8492 | v_8552;
assign v_8554 = v_8543 | v_8553;
assign v_8559 = v_8557 | v_8558;
assign v_8562 = v_8560 | v_8561;
assign v_8565 = v_8563 | v_8564;
assign v_8568 = v_8566 | v_8567;
assign v_8569 = ~v_8555 | v_8568;
assign v_8570 = v_8476 | ~v_8556;
assign v_8571 = v_8450 | v_8474;
assign v_8573 = v_8478 | v_8572;
assign v_8574 = v_91 | v_8453;
assign v_8576 = v_8485 | v_8575;
assign v_8577 = v_8460 | v_8483;
assign v_8579 = v_8492 | v_8578;
assign v_8580 = v_8467 | v_8490;
assign v_8582 = v_8555 | v_8581;
assign v_8585 = v_8476 | v_8584;
assign v_8586 = v_8478 | v_8585;
assign v_8587 = v_8485 | v_8586;
assign v_8588 = v_8492 | v_8587;
assign v_8589 = ~v_8583 | v_8588;
assign v_8594 = v_8583 | v_8593;
assign v_8596 = ~v_96 | v_8446;
assign v_8599 = ~v_807 | v_8159;
assign v_8601 = ~v_91 | v_8455;
assign v_8602 = ~v_91 | v_8457;
assign v_8604 = ~v_361 | v_8603;
assign v_8606 = ~v_91 | v_8462;
assign v_8607 = ~v_91 | v_8464;
assign v_8609 = ~v_563 | v_8608;
assign v_8611 = ~v_8595 | v_8610;
assign v_8613 = ~v_8597 | v_8612;
assign v_8615 = v_8613 | v_8614;
assign v_8618 = v_8616 | v_8617;
assign v_8620 = v_8615 | v_8619;
assign v_8623 = v_8621 | v_8622;
assign v_8625 = v_8620 | v_8624;
assign v_8626 = v_8595 | v_8625;
assign v_8633 = ~v_8627 | v_8632;
assign v_8634 = v_8612 | ~v_8628;
assign v_8635 = v_8614 | v_8634;
assign v_8636 = v_8619 | v_8635;
assign v_8637 = v_8624 | v_8636;
assign v_8638 = v_8627 | v_8637;
assign v_8645 = ~v_8639 | v_8644;
assign v_8646 = v_8612 | ~v_8640;
assign v_8647 = v_8614 | v_8646;
assign v_8648 = v_8619 | v_8647;
assign v_8649 = v_8624 | v_8648;
assign v_8650 = v_8639 | v_8649;
assign v_8657 = ~v_8651 | v_8656;
assign v_8658 = v_8612 | ~v_8652;
assign v_8659 = v_8614 | v_8658;
assign v_8660 = v_8619 | v_8659;
assign v_8661 = v_8624 | v_8660;
assign v_8662 = v_8651 | v_8661;
assign v_8669 = ~v_8663 | v_8668;
assign v_8670 = v_8612 | ~v_8664;
assign v_8671 = v_8614 | v_8670;
assign v_8672 = v_8619 | v_8671;
assign v_8673 = v_8624 | v_8672;
assign v_8674 = v_8663 | v_8673;
assign v_8681 = ~v_8675 | v_8680;
assign v_8682 = v_8612 | ~v_8676;
assign v_8683 = v_8614 | v_8682;
assign v_8684 = v_8619 | v_8683;
assign v_8685 = v_8624 | v_8684;
assign v_8686 = v_8675 | v_8685;
assign v_8691 = v_8689 | v_8690;
assign v_8694 = v_8692 | v_8693;
assign v_8697 = v_8695 | v_8696;
assign v_8700 = v_8698 | v_8699;
assign v_8701 = ~v_8687 | v_8700;
assign v_8702 = v_8612 | ~v_8688;
assign v_8703 = ~v_91 | v_8596;
assign v_8705 = v_8614 | v_8704;
assign v_8706 = v_8185 | v_8599;
assign v_8708 = v_8619 | v_8707;
assign v_8709 = v_8604 | v_8617;
assign v_8711 = v_8624 | v_8710;
assign v_8712 = v_8609 | v_8622;
assign v_8714 = v_8687 | v_8713;
assign v_8717 = v_8612 | v_8716;
assign v_8718 = v_8614 | v_8717;
assign v_8719 = v_8619 | v_8718;
assign v_8720 = v_8624 | v_8719;
assign v_8721 = ~v_8715 | v_8720;
assign v_8726 = v_8715 | v_8725;
assign v_8728 = ~v_89 | v_8445;
assign v_8729 = v_91 | v_8728;
assign v_8730 = ~v_91 | v_8446;
assign v_8732 = ~v_96 | v_8731;
assign v_8735 = ~v_807 | v_8156;
assign v_8737 = v_587 | v_7579;
assign v_8738 = ~v_87 | v_8737;
assign v_8739 = v_89 | v_8738;
assign v_8740 = v_91 | v_8739;
assign v_8741 = v_654 | v_7584;
assign v_8742 = ~v_87 | v_8741;
assign v_8743 = v_89 | v_8742;
assign v_8744 = v_91 | v_8743;
assign v_8746 = ~v_361 | v_8745;
assign v_8748 = v_587 | v_7592;
assign v_8749 = ~v_87 | v_8748;
assign v_8750 = v_89 | v_8749;
assign v_8751 = v_91 | v_8750;
assign v_8752 = v_654 | v_7597;
assign v_8753 = ~v_87 | v_8752;
assign v_8754 = v_89 | v_8753;
assign v_8755 = v_91 | v_8754;
assign v_8757 = ~v_563 | v_8756;
assign v_8759 = ~v_8727 | v_8758;
assign v_8763 = v_8761 | v_8762;
assign v_8765 = ~v_8733 | v_8764;
assign v_8767 = v_8765 | v_8766;
assign v_8776 = v_8771 | v_8775;
assign v_8778 = v_8767 | v_8777;
assign v_8787 = v_8782 | v_8786;
assign v_8789 = v_8778 | v_8788;
assign v_8790 = v_8727 | v_8789;
assign v_8797 = ~v_8791 | v_8796;
assign v_8798 = v_8764 | ~v_8792;
assign v_8799 = v_8766 | v_8798;
assign v_8800 = v_8777 | v_8799;
assign v_8801 = v_8788 | v_8800;
assign v_8802 = v_8791 | v_8801;
assign v_8809 = ~v_8803 | v_8808;
assign v_8810 = v_8764 | ~v_8804;
assign v_8811 = v_8766 | v_8810;
assign v_8812 = v_8777 | v_8811;
assign v_8813 = v_8788 | v_8812;
assign v_8814 = v_8803 | v_8813;
assign v_8821 = ~v_8815 | v_8820;
assign v_8822 = v_8764 | ~v_8816;
assign v_8823 = v_8766 | v_8822;
assign v_8824 = v_8777 | v_8823;
assign v_8825 = v_8788 | v_8824;
assign v_8826 = v_8815 | v_8825;
assign v_8833 = ~v_8827 | v_8832;
assign v_8834 = v_8764 | ~v_8828;
assign v_8835 = v_8766 | v_8834;
assign v_8836 = v_8777 | v_8835;
assign v_8837 = v_8788 | v_8836;
assign v_8838 = v_8827 | v_8837;
assign v_8845 = ~v_8839 | v_8844;
assign v_8846 = v_8764 | ~v_8840;
assign v_8847 = v_8766 | v_8846;
assign v_8848 = v_8777 | v_8847;
assign v_8849 = v_8788 | v_8848;
assign v_8850 = v_8839 | v_8849;
assign v_8855 = v_8853 | v_8854;
assign v_8858 = v_8856 | v_8857;
assign v_8861 = v_8859 | v_8860;
assign v_8864 = v_8862 | v_8863;
assign v_8865 = ~v_8851 | v_8864;
assign v_8866 = v_8764 | ~v_8852;
assign v_8867 = v_8732 | v_8762;
assign v_8869 = v_8766 | v_8868;
assign v_8870 = v_91 | v_8735;
assign v_8872 = v_8777 | v_8871;
assign v_8873 = v_8746 | v_8775;
assign v_8875 = v_8788 | v_8874;
assign v_8876 = v_8757 | v_8786;
assign v_8878 = v_8851 | v_8877;
assign v_8881 = v_8764 | v_8880;
assign v_8882 = v_8766 | v_8881;
assign v_8883 = v_8777 | v_8882;
assign v_8884 = v_8788 | v_8883;
assign v_8885 = ~v_8879 | v_8884;
assign v_8890 = v_8879 | v_8889;
assign v_8892 = ~v_96 | v_8728;
assign v_8895 = ~v_807 | v_8449;
assign v_8897 = ~v_91 | v_8739;
assign v_8898 = ~v_91 | v_8743;
assign v_8900 = ~v_361 | v_8899;
assign v_8902 = ~v_91 | v_8750;
assign v_8903 = ~v_91 | v_8754;
assign v_8905 = ~v_563 | v_8904;
assign v_8907 = ~v_8891 | v_8906;
assign v_8909 = ~v_8893 | v_8908;
assign v_8911 = v_8909 | v_8910;
assign v_8914 = v_8912 | v_8913;
assign v_8916 = v_8911 | v_8915;
assign v_8919 = v_8917 | v_8918;
assign v_8921 = v_8916 | v_8920;
assign v_8922 = v_8891 | v_8921;
assign v_8929 = ~v_8923 | v_8928;
assign v_8930 = v_8908 | ~v_8924;
assign v_8931 = v_8910 | v_8930;
assign v_8932 = v_8915 | v_8931;
assign v_8933 = v_8920 | v_8932;
assign v_8934 = v_8923 | v_8933;
assign v_8941 = ~v_8935 | v_8940;
assign v_8942 = v_8908 | ~v_8936;
assign v_8943 = v_8910 | v_8942;
assign v_8944 = v_8915 | v_8943;
assign v_8945 = v_8920 | v_8944;
assign v_8946 = v_8935 | v_8945;
assign v_8953 = ~v_8947 | v_8952;
assign v_8954 = v_8908 | ~v_8948;
assign v_8955 = v_8910 | v_8954;
assign v_8956 = v_8915 | v_8955;
assign v_8957 = v_8920 | v_8956;
assign v_8958 = v_8947 | v_8957;
assign v_8965 = ~v_8959 | v_8964;
assign v_8966 = v_8908 | ~v_8960;
assign v_8967 = v_8910 | v_8966;
assign v_8968 = v_8915 | v_8967;
assign v_8969 = v_8920 | v_8968;
assign v_8970 = v_8959 | v_8969;
assign v_8977 = ~v_8971 | v_8976;
assign v_8978 = v_8908 | ~v_8972;
assign v_8979 = v_8910 | v_8978;
assign v_8980 = v_8915 | v_8979;
assign v_8981 = v_8920 | v_8980;
assign v_8982 = v_8971 | v_8981;
assign v_8987 = v_8985 | v_8986;
assign v_8990 = v_8988 | v_8989;
assign v_8993 = v_8991 | v_8992;
assign v_8996 = v_8994 | v_8995;
assign v_8997 = ~v_8983 | v_8996;
assign v_8998 = v_8908 | ~v_8984;
assign v_8999 = ~v_91 | v_8892;
assign v_9001 = v_8910 | v_9000;
assign v_9002 = v_8473 | v_8895;
assign v_9004 = v_8915 | v_9003;
assign v_9005 = v_8900 | v_8913;
assign v_9007 = v_8920 | v_9006;
assign v_9008 = v_8905 | v_8918;
assign v_9010 = v_8983 | v_9009;
assign v_9013 = v_8908 | v_9012;
assign v_9014 = v_8910 | v_9013;
assign v_9015 = v_8915 | v_9014;
assign v_9016 = v_8920 | v_9015;
assign v_9017 = ~v_9011 | v_9016;
assign v_9022 = v_9011 | v_9021;
assign v_9024 = v_87 | v_8444;
assign v_9025 = v_89 | v_9024;
assign v_9026 = v_91 | v_9025;
assign v_9027 = ~v_91 | v_8728;
assign v_9029 = ~v_96 | v_9028;
assign v_9032 = ~v_807 | v_8446;
assign v_9034 = ~v_89 | v_8738;
assign v_9035 = v_91 | v_9034;
assign v_9036 = ~v_89 | v_8742;
assign v_9037 = v_91 | v_9036;
assign v_9039 = ~v_361 | v_9038;
assign v_9041 = ~v_89 | v_8749;
assign v_9042 = v_91 | v_9041;
assign v_9043 = ~v_89 | v_8753;
assign v_9044 = v_91 | v_9043;
assign v_9046 = ~v_563 | v_9045;
assign v_9048 = ~v_9023 | v_9047;
assign v_9053 = v_9051 | v_9052;
assign v_9055 = ~v_9030 | v_9054;
assign v_9057 = v_9055 | v_9056;
assign v_9062 = v_9059 | v_9061;
assign v_9064 = v_9057 | v_9063;
assign v_9069 = v_9066 | v_9068;
assign v_9071 = v_9064 | v_9070;
assign v_9072 = v_9023 | v_9071;
assign v_9079 = ~v_9073 | v_9078;
assign v_9080 = v_9054 | ~v_9074;
assign v_9081 = v_9056 | v_9080;
assign v_9082 = v_9063 | v_9081;
assign v_9083 = v_9070 | v_9082;
assign v_9084 = v_9073 | v_9083;
assign v_9091 = ~v_9085 | v_9090;
assign v_9092 = v_9054 | ~v_9086;
assign v_9093 = v_9056 | v_9092;
assign v_9094 = v_9063 | v_9093;
assign v_9095 = v_9070 | v_9094;
assign v_9096 = v_9085 | v_9095;
assign v_9103 = ~v_9097 | v_9102;
assign v_9104 = v_9054 | ~v_9098;
assign v_9105 = v_9056 | v_9104;
assign v_9106 = v_9063 | v_9105;
assign v_9107 = v_9070 | v_9106;
assign v_9108 = v_9097 | v_9107;
assign v_9115 = ~v_9109 | v_9114;
assign v_9116 = v_9054 | ~v_9110;
assign v_9117 = v_9056 | v_9116;
assign v_9118 = v_9063 | v_9117;
assign v_9119 = v_9070 | v_9118;
assign v_9120 = v_9109 | v_9119;
assign v_9127 = ~v_9121 | v_9126;
assign v_9128 = v_9054 | ~v_9122;
assign v_9129 = v_9056 | v_9128;
assign v_9130 = v_9063 | v_9129;
assign v_9131 = v_9070 | v_9130;
assign v_9132 = v_9121 | v_9131;
assign v_9137 = v_9135 | v_9136;
assign v_9140 = v_9138 | v_9139;
assign v_9143 = v_9141 | v_9142;
assign v_9146 = v_9144 | v_9145;
assign v_9147 = ~v_9133 | v_9146;
assign v_9148 = v_9054 | ~v_9134;
assign v_9149 = v_9029 | v_9052;
assign v_9151 = v_9056 | v_9150;
assign v_9152 = v_91 | v_9032;
assign v_9154 = v_9063 | v_9153;
assign v_9155 = v_9039 | v_9061;
assign v_9157 = v_9070 | v_9156;
assign v_9158 = v_9046 | v_9068;
assign v_9160 = v_9133 | v_9159;
assign v_9163 = v_9054 | v_9162;
assign v_9164 = v_9056 | v_9163;
assign v_9165 = v_9063 | v_9164;
assign v_9166 = v_9070 | v_9165;
assign v_9167 = ~v_9161 | v_9166;
assign v_9172 = v_9161 | v_9171;
assign v_9174 = ~v_96 | v_9025;
assign v_9177 = ~v_807 | v_8731;
assign v_9179 = ~v_91 | v_9034;
assign v_9180 = ~v_91 | v_9036;
assign v_9182 = ~v_361 | v_9181;
assign v_9184 = ~v_91 | v_9041;
assign v_9185 = ~v_91 | v_9043;
assign v_9187 = ~v_563 | v_9186;
assign v_9189 = ~v_9173 | v_9188;
assign v_9191 = ~v_9175 | v_9190;
assign v_9193 = v_9191 | v_9192;
assign v_9196 = v_9194 | v_9195;
assign v_9198 = v_9193 | v_9197;
assign v_9201 = v_9199 | v_9200;
assign v_9203 = v_9198 | v_9202;
assign v_9204 = v_9173 | v_9203;
assign v_9211 = ~v_9205 | v_9210;
assign v_9212 = v_9190 | ~v_9206;
assign v_9213 = v_9192 | v_9212;
assign v_9214 = v_9197 | v_9213;
assign v_9215 = v_9202 | v_9214;
assign v_9216 = v_9205 | v_9215;
assign v_9223 = ~v_9217 | v_9222;
assign v_9224 = v_9190 | ~v_9218;
assign v_9225 = v_9192 | v_9224;
assign v_9226 = v_9197 | v_9225;
assign v_9227 = v_9202 | v_9226;
assign v_9228 = v_9217 | v_9227;
assign v_9235 = ~v_9229 | v_9234;
assign v_9236 = v_9190 | ~v_9230;
assign v_9237 = v_9192 | v_9236;
assign v_9238 = v_9197 | v_9237;
assign v_9239 = v_9202 | v_9238;
assign v_9240 = v_9229 | v_9239;
assign v_9247 = ~v_9241 | v_9246;
assign v_9248 = v_9190 | ~v_9242;
assign v_9249 = v_9192 | v_9248;
assign v_9250 = v_9197 | v_9249;
assign v_9251 = v_9202 | v_9250;
assign v_9252 = v_9241 | v_9251;
assign v_9259 = ~v_9253 | v_9258;
assign v_9260 = v_9190 | ~v_9254;
assign v_9261 = v_9192 | v_9260;
assign v_9262 = v_9197 | v_9261;
assign v_9263 = v_9202 | v_9262;
assign v_9264 = v_9253 | v_9263;
assign v_9269 = v_9267 | v_9268;
assign v_9272 = v_9270 | v_9271;
assign v_9275 = v_9273 | v_9274;
assign v_9278 = v_9276 | v_9277;
assign v_9279 = ~v_9265 | v_9278;
assign v_9280 = v_9190 | ~v_9266;
assign v_9281 = ~v_91 | v_9174;
assign v_9283 = v_9192 | v_9282;
assign v_9284 = v_8761 | v_9177;
assign v_9286 = v_9197 | v_9285;
assign v_9287 = v_9182 | v_9195;
assign v_9289 = v_9202 | v_9288;
assign v_9290 = v_9187 | v_9200;
assign v_9292 = v_9265 | v_9291;
assign v_9295 = v_9190 | v_9294;
assign v_9296 = v_9192 | v_9295;
assign v_9297 = v_9197 | v_9296;
assign v_9298 = v_9202 | v_9297;
assign v_9299 = ~v_9293 | v_9298;
assign v_9304 = v_9293 | v_9303;
assign v_9306 = ~v_89 | v_9024;
assign v_9307 = v_91 | v_9306;
assign v_9308 = ~v_91 | v_9025;
assign v_9310 = ~v_96 | v_9309;
assign v_9313 = ~v_807 | v_8728;
assign v_9315 = v_87 | v_8737;
assign v_9316 = v_89 | v_9315;
assign v_9317 = v_91 | v_9316;
assign v_9318 = v_87 | v_8741;
assign v_9319 = v_89 | v_9318;
assign v_9320 = v_91 | v_9319;
assign v_9322 = ~v_361 | v_9321;
assign v_9324 = v_87 | v_8748;
assign v_9325 = v_89 | v_9324;
assign v_9326 = v_91 | v_9325;
assign v_9327 = v_87 | v_8752;
assign v_9328 = v_89 | v_9327;
assign v_9329 = v_91 | v_9328;
assign v_9331 = ~v_563 | v_9330;
assign v_9333 = ~v_9305 | v_9332;
assign v_9337 = v_9335 | v_9336;
assign v_9339 = ~v_9311 | v_9338;
assign v_9341 = v_9339 | v_9340;
assign v_9348 = v_9344 | v_9347;
assign v_9350 = v_9341 | v_9349;
assign v_9357 = v_9353 | v_9356;
assign v_9359 = v_9350 | v_9358;
assign v_9360 = v_9305 | v_9359;
assign v_9367 = ~v_9361 | v_9366;
assign v_9368 = v_9338 | ~v_9362;
assign v_9369 = v_9340 | v_9368;
assign v_9370 = v_9349 | v_9369;
assign v_9371 = v_9358 | v_9370;
assign v_9372 = v_9361 | v_9371;
assign v_9379 = ~v_9373 | v_9378;
assign v_9380 = v_9338 | ~v_9374;
assign v_9381 = v_9340 | v_9380;
assign v_9382 = v_9349 | v_9381;
assign v_9383 = v_9358 | v_9382;
assign v_9384 = v_9373 | v_9383;
assign v_9391 = ~v_9385 | v_9390;
assign v_9392 = v_9338 | ~v_9386;
assign v_9393 = v_9340 | v_9392;
assign v_9394 = v_9349 | v_9393;
assign v_9395 = v_9358 | v_9394;
assign v_9396 = v_9385 | v_9395;
assign v_9403 = ~v_9397 | v_9402;
assign v_9404 = v_9338 | ~v_9398;
assign v_9405 = v_9340 | v_9404;
assign v_9406 = v_9349 | v_9405;
assign v_9407 = v_9358 | v_9406;
assign v_9408 = v_9397 | v_9407;
assign v_9415 = ~v_9409 | v_9414;
assign v_9416 = v_9338 | ~v_9410;
assign v_9417 = v_9340 | v_9416;
assign v_9418 = v_9349 | v_9417;
assign v_9419 = v_9358 | v_9418;
assign v_9420 = v_9409 | v_9419;
assign v_9425 = v_9423 | v_9424;
assign v_9428 = v_9426 | v_9427;
assign v_9431 = v_9429 | v_9430;
assign v_9434 = v_9432 | v_9433;
assign v_9435 = ~v_9421 | v_9434;
assign v_9436 = v_9338 | ~v_9422;
assign v_9437 = v_9310 | v_9336;
assign v_9439 = v_9340 | v_9438;
assign v_9440 = v_91 | v_9313;
assign v_9442 = v_9349 | v_9441;
assign v_9443 = v_9322 | v_9347;
assign v_9445 = v_9358 | v_9444;
assign v_9446 = v_9331 | v_9356;
assign v_9448 = v_9421 | v_9447;
assign v_9451 = v_9338 | v_9450;
assign v_9452 = v_9340 | v_9451;
assign v_9453 = v_9349 | v_9452;
assign v_9454 = v_9358 | v_9453;
assign v_9455 = ~v_9449 | v_9454;
assign v_9460 = v_9449 | v_9459;
assign v_9462 = ~v_96 | v_9306;
assign v_9465 = ~v_807 | v_9028;
assign v_9467 = ~v_91 | v_9316;
assign v_9468 = ~v_91 | v_9319;
assign v_9470 = ~v_361 | v_9469;
assign v_9472 = ~v_91 | v_9325;
assign v_9473 = ~v_91 | v_9328;
assign v_9475 = ~v_563 | v_9474;
assign v_9477 = ~v_9461 | v_9476;
assign v_9479 = ~v_9463 | v_9478;
assign v_9481 = v_9479 | v_9480;
assign v_9484 = v_9482 | v_9483;
assign v_9486 = v_9481 | v_9485;
assign v_9489 = v_9487 | v_9488;
assign v_9491 = v_9486 | v_9490;
assign v_9492 = v_9461 | v_9491;
assign v_9499 = ~v_9493 | v_9498;
assign v_9500 = v_9478 | ~v_9494;
assign v_9501 = v_9480 | v_9500;
assign v_9502 = v_9485 | v_9501;
assign v_9503 = v_9490 | v_9502;
assign v_9504 = v_9493 | v_9503;
assign v_9511 = ~v_9505 | v_9510;
assign v_9512 = v_9478 | ~v_9506;
assign v_9513 = v_9480 | v_9512;
assign v_9514 = v_9485 | v_9513;
assign v_9515 = v_9490 | v_9514;
assign v_9516 = v_9505 | v_9515;
assign v_9523 = ~v_9517 | v_9522;
assign v_9524 = v_9478 | ~v_9518;
assign v_9525 = v_9480 | v_9524;
assign v_9526 = v_9485 | v_9525;
assign v_9527 = v_9490 | v_9526;
assign v_9528 = v_9517 | v_9527;
assign v_9535 = ~v_9529 | v_9534;
assign v_9536 = v_9478 | ~v_9530;
assign v_9537 = v_9480 | v_9536;
assign v_9538 = v_9485 | v_9537;
assign v_9539 = v_9490 | v_9538;
assign v_9540 = v_9529 | v_9539;
assign v_9547 = ~v_9541 | v_9546;
assign v_9548 = v_9478 | ~v_9542;
assign v_9549 = v_9480 | v_9548;
assign v_9550 = v_9485 | v_9549;
assign v_9551 = v_9490 | v_9550;
assign v_9552 = v_9541 | v_9551;
assign v_9557 = v_9555 | v_9556;
assign v_9560 = v_9558 | v_9559;
assign v_9563 = v_9561 | v_9562;
assign v_9566 = v_9564 | v_9565;
assign v_9567 = ~v_9553 | v_9566;
assign v_9568 = v_9478 | ~v_9554;
assign v_9569 = ~v_91 | v_9462;
assign v_9571 = v_9480 | v_9570;
assign v_9572 = v_9051 | v_9465;
assign v_9574 = v_9485 | v_9573;
assign v_9575 = v_9470 | v_9483;
assign v_9577 = v_9490 | v_9576;
assign v_9578 = v_9475 | v_9488;
assign v_9580 = v_9553 | v_9579;
assign v_9583 = v_9478 | v_9582;
assign v_9584 = v_9480 | v_9583;
assign v_9585 = v_9485 | v_9584;
assign v_9586 = v_9490 | v_9585;
assign v_9587 = ~v_9581 | v_9586;
assign v_9592 = v_9581 | v_9591;
assign v_9594 = v_74 | v_578;
assign v_9595 = v_79 | v_9594;
assign v_9596 = v_82 | v_9595;
assign v_9597 = v_85 | v_9596;
assign v_9598 = ~v_87 | v_9597;
assign v_9599 = v_89 | v_9598;
assign v_9600 = v_91 | v_9599;
assign v_9601 = ~v_91 | v_9306;
assign v_9603 = ~v_96 | v_9602;
assign v_9606 = ~v_807 | v_9025;
assign v_9608 = ~v_89 | v_9315;
assign v_9609 = v_91 | v_9608;
assign v_9610 = ~v_89 | v_9318;
assign v_9611 = v_91 | v_9610;
assign v_9613 = ~v_361 | v_9612;
assign v_9615 = ~v_89 | v_9324;
assign v_9616 = v_91 | v_9615;
assign v_9617 = ~v_89 | v_9327;
assign v_9618 = v_91 | v_9617;
assign v_9620 = ~v_563 | v_9619;
assign v_9622 = ~v_9593 | v_9621;
assign v_9631 = v_9629 | v_9630;
assign v_9633 = ~v_9604 | v_9632;
assign v_9635 = v_9633 | v_9634;
assign v_9640 = v_9637 | v_9639;
assign v_9642 = v_9635 | v_9641;
assign v_9647 = v_9644 | v_9646;
assign v_9649 = v_9642 | v_9648;
assign v_9650 = v_9593 | v_9649;
assign v_9657 = ~v_9651 | v_9656;
assign v_9658 = v_9632 | ~v_9652;
assign v_9659 = v_9634 | v_9658;
assign v_9660 = v_9641 | v_9659;
assign v_9661 = v_9648 | v_9660;
assign v_9662 = v_9651 | v_9661;
assign v_9669 = ~v_9663 | v_9668;
assign v_9670 = v_9632 | ~v_9664;
assign v_9671 = v_9634 | v_9670;
assign v_9672 = v_9641 | v_9671;
assign v_9673 = v_9648 | v_9672;
assign v_9674 = v_9663 | v_9673;
assign v_9681 = ~v_9675 | v_9680;
assign v_9682 = v_9632 | ~v_9676;
assign v_9683 = v_9634 | v_9682;
assign v_9684 = v_9641 | v_9683;
assign v_9685 = v_9648 | v_9684;
assign v_9686 = v_9675 | v_9685;
assign v_9693 = ~v_9687 | v_9692;
assign v_9694 = v_9632 | ~v_9688;
assign v_9695 = v_9634 | v_9694;
assign v_9696 = v_9641 | v_9695;
assign v_9697 = v_9648 | v_9696;
assign v_9698 = v_9687 | v_9697;
assign v_9705 = ~v_9699 | v_9704;
assign v_9706 = v_9632 | ~v_9700;
assign v_9707 = v_9634 | v_9706;
assign v_9708 = v_9641 | v_9707;
assign v_9709 = v_9648 | v_9708;
assign v_9710 = v_9699 | v_9709;
assign v_9715 = v_9713 | v_9714;
assign v_9718 = v_9716 | v_9717;
assign v_9721 = v_9719 | v_9720;
assign v_9724 = v_9722 | v_9723;
assign v_9725 = ~v_9711 | v_9724;
assign v_9726 = v_9632 | ~v_9712;
assign v_9727 = v_9603 | v_9630;
assign v_9729 = v_9634 | v_9728;
assign v_9730 = v_91 | v_9606;
assign v_9732 = v_9641 | v_9731;
assign v_9733 = v_9613 | v_9639;
assign v_9735 = v_9648 | v_9734;
assign v_9736 = v_9620 | v_9646;
assign v_9738 = v_9711 | v_9737;
assign v_9741 = v_9632 | v_9740;
assign v_9742 = v_9634 | v_9741;
assign v_9743 = v_9641 | v_9742;
assign v_9744 = v_9648 | v_9743;
assign v_9745 = ~v_9739 | v_9744;
assign v_9750 = v_9739 | v_9749;
assign v_9752 = ~v_96 | v_9599;
assign v_9755 = ~v_807 | v_9309;
assign v_9757 = ~v_91 | v_9608;
assign v_9758 = ~v_91 | v_9610;
assign v_9760 = ~v_361 | v_9759;
assign v_9762 = ~v_91 | v_9615;
assign v_9763 = ~v_91 | v_9617;
assign v_9765 = ~v_563 | v_9764;
assign v_9767 = ~v_9751 | v_9766;
assign v_9769 = ~v_9753 | v_9768;
assign v_9771 = v_9769 | v_9770;
assign v_9774 = v_9772 | v_9773;
assign v_9776 = v_9771 | v_9775;
assign v_9779 = v_9777 | v_9778;
assign v_9781 = v_9776 | v_9780;
assign v_9782 = v_9751 | v_9781;
assign v_9789 = ~v_9783 | v_9788;
assign v_9790 = v_9768 | ~v_9784;
assign v_9791 = v_9770 | v_9790;
assign v_9792 = v_9775 | v_9791;
assign v_9793 = v_9780 | v_9792;
assign v_9794 = v_9783 | v_9793;
assign v_9801 = ~v_9795 | v_9800;
assign v_9802 = v_9768 | ~v_9796;
assign v_9803 = v_9770 | v_9802;
assign v_9804 = v_9775 | v_9803;
assign v_9805 = v_9780 | v_9804;
assign v_9806 = v_9795 | v_9805;
assign v_9813 = ~v_9807 | v_9812;
assign v_9814 = v_9768 | ~v_9808;
assign v_9815 = v_9770 | v_9814;
assign v_9816 = v_9775 | v_9815;
assign v_9817 = v_9780 | v_9816;
assign v_9818 = v_9807 | v_9817;
assign v_9825 = ~v_9819 | v_9824;
assign v_9826 = v_9768 | ~v_9820;
assign v_9827 = v_9770 | v_9826;
assign v_9828 = v_9775 | v_9827;
assign v_9829 = v_9780 | v_9828;
assign v_9830 = v_9819 | v_9829;
assign v_9837 = ~v_9831 | v_9836;
assign v_9838 = v_9768 | ~v_9832;
assign v_9839 = v_9770 | v_9838;
assign v_9840 = v_9775 | v_9839;
assign v_9841 = v_9780 | v_9840;
assign v_9842 = v_9831 | v_9841;
assign v_9847 = v_9845 | v_9846;
assign v_9850 = v_9848 | v_9849;
assign v_9853 = v_9851 | v_9852;
assign v_9856 = v_9854 | v_9855;
assign v_9857 = ~v_9843 | v_9856;
assign v_9858 = v_9768 | ~v_9844;
assign v_9859 = ~v_91 | v_9752;
assign v_9861 = v_9770 | v_9860;
assign v_9862 = v_9335 | v_9755;
assign v_9864 = v_9775 | v_9863;
assign v_9865 = v_9760 | v_9773;
assign v_9867 = v_9780 | v_9866;
assign v_9868 = v_9765 | v_9778;
assign v_9870 = v_9843 | v_9869;
assign v_9873 = v_9768 | v_9872;
assign v_9874 = v_9770 | v_9873;
assign v_9875 = v_9775 | v_9874;
assign v_9876 = v_9780 | v_9875;
assign v_9877 = ~v_9871 | v_9876;
assign v_9882 = v_9871 | v_9881;
assign v_9886 = v_89 | v_91;
assign v_9887 = ~v_87 | v_9886;
assign v_9888 = v_29 | v_9887;
assign v_9889 = v_24 | v_9888;
assign v_9890 = v_19 | v_9889;
assign v_9891 = v_14 | v_9890;
assign v_9892 = ~v_9 | v_9891;
assign v_9899 = v_9 | v_9898;
assign v_9902 = v_9885 | v_9901;
assign v_9911 = v_9 | v_9910;
assign v_9912 = ~v_89 | ~v_91;
assign v_9913 = v_87 | v_9912;
assign v_9914 = ~v_29 | v_9913;
assign v_9915 = ~v_24 | v_9914;
assign v_9916 = ~v_19 | v_9915;
assign v_9917 = ~v_14 | v_9916;
assign v_9918 = ~v_9 | v_9917;
assign v_9921 = v_9904 | v_9920;
assign v_9924 = v_9922 | v_9923;
assign v_9927 = v_9925 | v_9926;
assign v_9928 = ~v_9883 | v_9927;
assign v_9929 = ~v_9 | v_9884;
assign v_9932 = v_9930 | v_9931;
assign v_9933 = ~v_9884 | v_9932;
assign v_9935 = v_9903 | v_9934;
assign v_9938 = v_9936 | v_9937;
assign v_9939 = ~v_9903 | v_9938;
assign v_9941 = v_96 | v_9940;
assign v_9942 = ~v_96 | v_9932;
assign v_9944 = v_807 | v_9943;
assign v_9945 = ~v_807 | v_9938;
assign v_9947 = v_9883 | v_9946;
assign v_9950 = ~v_14 | v_9890;
assign v_9951 = v_14 | v_9897;
assign v_9954 = v_9949 | v_9953;
assign v_9956 = v_14 | v_9909;
assign v_9959 = v_9955 | v_9958;
assign v_9962 = v_9960 | v_9961;
assign v_9965 = v_9963 | v_9964;
assign v_9966 = ~v_9948 | v_9965;
assign v_9967 = ~v_14 | v_9884;
assign v_9970 = v_9968 | v_9969;
assign v_9971 = ~v_9884 | v_9970;
assign v_9973 = v_9903 | v_9972;
assign v_9975 = v_9910 | v_9974;
assign v_9976 = ~v_9903 | v_9975;
assign v_9978 = v_96 | v_9977;
assign v_9979 = ~v_96 | v_9970;
assign v_9981 = v_807 | v_9980;
assign v_9982 = ~v_807 | v_9975;
assign v_9984 = v_9948 | v_9983;
assign v_9987 = ~v_19 | v_9889;
assign v_9988 = v_19 | v_9896;
assign v_9991 = v_9986 | v_9990;
assign v_9993 = v_19 | v_9908;
assign v_9996 = v_9992 | v_9995;
assign v_9999 = v_9997 | v_9998;
assign v_10002 = v_10000 | v_10001;
assign v_10003 = ~v_9985 | v_10002;
assign v_10004 = ~v_19 | v_9884;
assign v_10007 = v_10005 | v_10006;
assign v_10008 = ~v_9884 | v_10007;
assign v_10010 = v_9903 | v_10009;
assign v_10012 = v_9909 | v_10011;
assign v_10013 = ~v_9903 | v_10012;
assign v_10015 = v_96 | v_10014;
assign v_10016 = ~v_96 | v_10007;
assign v_10018 = v_807 | v_10017;
assign v_10019 = ~v_807 | v_10012;
assign v_10021 = v_9985 | v_10020;
assign v_10024 = ~v_24 | v_9888;
assign v_10025 = v_24 | v_9895;
assign v_10028 = v_10023 | v_10027;
assign v_10030 = v_24 | v_9907;
assign v_10033 = v_10029 | v_10032;
assign v_10036 = v_10034 | v_10035;
assign v_10039 = v_10037 | v_10038;
assign v_10040 = ~v_10022 | v_10039;
assign v_10041 = ~v_24 | v_9884;
assign v_10044 = v_10042 | v_10043;
assign v_10045 = ~v_9884 | v_10044;
assign v_10047 = v_9903 | v_10046;
assign v_10049 = v_9908 | v_10048;
assign v_10050 = ~v_9903 | v_10049;
assign v_10052 = v_96 | v_10051;
assign v_10053 = ~v_96 | v_10044;
assign v_10055 = v_807 | v_10054;
assign v_10056 = ~v_807 | v_10049;
assign v_10058 = v_10022 | v_10057;
assign v_10061 = ~v_29 | v_9887;
assign v_10062 = v_29 | v_9894;
assign v_10065 = v_10060 | v_10064;
assign v_10067 = v_29 | v_9906;
assign v_10070 = v_10066 | v_10069;
assign v_10073 = v_10071 | v_10072;
assign v_10076 = v_10074 | v_10075;
assign v_10077 = ~v_10059 | v_10076;
assign v_10078 = ~v_29 | v_9884;
assign v_10081 = v_10079 | v_10080;
assign v_10082 = ~v_9884 | v_10081;
assign v_10084 = v_9903 | v_10083;
assign v_10086 = v_9907 | v_10085;
assign v_10087 = ~v_9903 | v_10086;
assign v_10089 = v_96 | v_10088;
assign v_10090 = ~v_96 | v_10081;
assign v_10092 = v_807 | v_10091;
assign v_10093 = ~v_807 | v_10086;
assign v_10095 = v_10059 | v_10094;
assign v_10097 = v_87 | v_9884;
assign v_10100 = v_10098 | v_10099;
assign v_10101 = ~v_9884 | v_10100;
assign v_10103 = v_9903 | v_10102;
assign v_10105 = v_9906 | v_10104;
assign v_10106 = ~v_9903 | v_10105;
assign v_10108 = v_96 | v_10107;
assign v_10109 = ~v_96 | v_10100;
assign v_10111 = v_807 | v_10110;
assign v_10112 = ~v_807 | v_10105;
assign v_10114 = ~v_10096 | v_10113;
assign v_10116 = v_87 | v_9886;
assign v_10117 = ~v_87 | v_9893;
assign v_10120 = v_10115 | v_10119;
assign v_10122 = ~v_87 | v_9905;
assign v_10125 = v_10121 | v_10124;
assign v_10128 = v_10126 | v_10127;
assign v_10131 = v_10129 | v_10130;
assign v_10132 = v_10096 | v_10131;
assign v_10135 = ~v_89 | v_91;
assign v_10136 = v_89 | ~v_91;
assign v_10139 = v_10134 | v_10138;
assign v_10143 = v_10140 | v_10142;
assign v_10146 = v_10144 | v_10145;
assign v_10149 = v_10147 | v_10148;
assign v_10150 = ~v_10133 | v_10149;
assign v_10151 = ~v_89 | v_9884;
assign v_10154 = v_10152 | v_10153;
assign v_10155 = ~v_9884 | v_10154;
assign v_10157 = v_9903 | v_10156;
assign v_10158 = v_9893 | v_9905;
assign v_10159 = ~v_9903 | v_10158;
assign v_10161 = v_96 | v_10160;
assign v_10162 = ~v_96 | v_10154;
assign v_10164 = v_807 | v_10163;
assign v_10165 = ~v_807 | v_10158;
assign v_10167 = v_10133 | v_10166;
assign v_10171 = v_10169 | v_10170;
assign v_10174 = v_10172 | v_10173;
assign v_10177 = v_10175 | v_10176;
assign v_10180 = v_10178 | v_10179;
assign v_10181 = ~v_10168 | v_10180;
assign v_10182 = ~v_91 | v_9884;
assign v_10183 = v_91 | ~v_9884;
assign v_10185 = v_9903 | v_10184;
assign v_10186 = v_91 | ~v_9903;
assign v_10188 = v_96 | v_10187;
assign v_10189 = v_91 | ~v_96;
assign v_10191 = v_807 | v_10190;
assign v_10192 = v_91 | ~v_807;
assign v_10194 = v_10168 | v_10193;
assign v_10199 = v_10197 | v_10198;
assign v_10203 = v_10201 | v_10202;
assign v_10206 = v_10204 | v_10205;
assign v_10209 = v_10207 | v_10208;
assign v_10210 = ~v_10195 | v_10209;
assign v_10211 = ~v_47 | v_10196;
assign v_10212 = v_239 | ~v_10196;
assign v_10214 = v_10200 | v_10213;
assign v_10215 = v_689 | ~v_10200;
assign v_10217 = v_361 | v_10216;
assign v_10218 = v_239 | ~v_361;
assign v_10220 = v_563 | v_10219;
assign v_10221 = ~v_563 | v_689;
assign v_10223 = v_10195 | v_10222;
assign v_10227 = v_10225 | v_10226;
assign v_10230 = v_10228 | v_10229;
assign v_10233 = v_10231 | v_10232;
assign v_10236 = v_10234 | v_10235;
assign v_10237 = ~v_10224 | v_10236;
assign v_10238 = ~v_45 | v_10196;
assign v_10239 = v_242 | ~v_10196;
assign v_10241 = v_10200 | v_10240;
assign v_10242 = v_520 | ~v_10200;
assign v_10244 = v_361 | v_10243;
assign v_10245 = v_242 | ~v_361;
assign v_10247 = v_563 | v_10246;
assign v_10248 = v_520 | ~v_563;
assign v_10250 = v_10224 | v_10249;
assign v_10254 = v_10252 | v_10253;
assign v_10257 = v_10255 | v_10256;
assign v_10260 = v_10258 | v_10259;
assign v_10263 = v_10261 | v_10262;
assign v_10264 = ~v_10251 | v_10263;
assign v_10265 = ~v_43 | v_10196;
assign v_10266 = v_294 | ~v_10196;
assign v_10268 = v_10200 | v_10267;
assign v_10269 = v_538 | ~v_10200;
assign v_10271 = v_361 | v_10270;
assign v_10272 = v_294 | ~v_361;
assign v_10274 = v_563 | v_10273;
assign v_10275 = v_538 | ~v_563;
assign v_10277 = v_10251 | v_10276;
assign v_10281 = v_10279 | v_10280;
assign v_10284 = v_10282 | v_10283;
assign v_10287 = v_10285 | v_10286;
assign v_10290 = v_10288 | v_10289;
assign v_10291 = ~v_10278 | v_10290;
assign v_10292 = ~v_8 | v_10196;
assign v_10293 = v_245 | ~v_10196;
assign v_10295 = v_10200 | v_10294;
assign v_10296 = v_475 | ~v_10200;
assign v_10298 = v_361 | v_10297;
assign v_10299 = v_245 | ~v_361;
assign v_10301 = v_563 | v_10300;
assign v_10302 = v_475 | ~v_563;
assign v_10304 = v_10278 | v_10303;
assign v_10308 = v_10306 | v_10307;
assign v_10311 = v_10309 | v_10310;
assign v_10314 = v_10312 | v_10313;
assign v_10317 = v_10315 | v_10316;
assign v_10318 = ~v_10305 | v_10317;
assign v_10319 = ~v_13 | v_10196;
assign v_10320 = v_254 | ~v_10196;
assign v_10322 = v_10200 | v_10321;
assign v_10323 = v_482 | ~v_10200;
assign v_10325 = v_361 | v_10324;
assign v_10326 = v_254 | ~v_361;
assign v_10328 = v_563 | v_10327;
assign v_10329 = v_482 | ~v_563;
assign v_10331 = v_10305 | v_10330;
assign v_10333 = v_18 | v_10196;
assign v_10334 = v_263 | ~v_10196;
assign v_10336 = v_10200 | v_10335;
assign v_10337 = v_489 | ~v_10200;
assign v_10339 = v_361 | v_10338;
assign v_10340 = v_263 | ~v_361;
assign v_10342 = v_563 | v_10341;
assign v_10343 = v_489 | ~v_563;
assign v_10345 = ~v_10332 | v_10344;
assign v_10348 = v_10346 | v_10347;
assign v_10351 = v_10349 | v_10350;
assign v_10354 = v_10352 | v_10353;
assign v_10357 = v_10355 | v_10356;
assign v_10358 = v_10332 | v_10357;
assign v_10360 = v_23 | v_10196;
assign v_10361 = v_272 | ~v_10196;
assign v_10363 = v_10200 | v_10362;
assign v_10364 = v_494 | ~v_10200;
assign v_10366 = v_361 | v_10365;
assign v_10367 = v_272 | ~v_361;
assign v_10369 = v_563 | v_10368;
assign v_10370 = v_494 | ~v_563;
assign v_10372 = ~v_10359 | v_10371;
assign v_10375 = v_10373 | v_10374;
assign v_10378 = v_10376 | v_10377;
assign v_10381 = v_10379 | v_10380;
assign v_10384 = v_10382 | v_10383;
assign v_10385 = v_10359 | v_10384;
assign v_10389 = v_10387 | v_10388;
assign v_10392 = v_10390 | v_10391;
assign v_10395 = v_10393 | v_10394;
assign v_10398 = v_10396 | v_10397;
assign v_10399 = ~v_10386 | v_10398;
assign v_10400 = ~v_28 | v_10196;
assign v_10401 = v_28 | ~v_10196;
assign v_10403 = v_10200 | v_10402;
assign v_10404 = v_28 | ~v_10200;
assign v_10406 = v_361 | v_10405;
assign v_10407 = v_28 | ~v_361;
assign v_10409 = v_563 | v_10408;
assign v_10410 = v_28 | ~v_563;
assign v_10412 = v_10386 | v_10411;
assign v_10417 = ~v_10413 | v_10416;
assign v_10418 = ~v_10414 | v_10415;
assign v_10419 = v_10413 | v_10418;
assign v_10423 = ~v_10420 | v_10422;
assign v_10424 = v_10415 | ~v_10421;
assign v_10425 = v_10420 | v_10424;
assign v_10429 = ~v_10426 | v_10428;
assign v_10430 = v_10415 | ~v_10427;
assign v_10431 = v_10426 | v_10430;
assign v_10435 = ~v_10432 | v_10434;
assign v_10436 = v_10415 | ~v_10433;
assign v_10437 = v_10432 | v_10436;
assign v_10441 = ~v_10438 | v_10440;
assign v_10442 = v_10415 | ~v_10439;
assign v_10443 = v_10438 | v_10442;
assign v_10447 = ~v_10444 | v_10446;
assign v_10448 = v_10415 | ~v_10445;
assign v_10449 = v_10444 | v_10448;
assign v_10453 = ~v_10450 | v_10452;
assign v_10454 = v_10415 | ~v_10451;
assign v_10455 = v_10450 | v_10454;
assign v_10457 = v_4 | v_10415;
assign v_10458 = ~v_10456 | v_10457;
assign v_10460 = v_10456 | v_10459;
assign v_10463 = ~v_10461 | v_10462;
assign v_10464 = v_10461 | ~v_10462;
assign v_10466 = v_9884 | v_10415;
assign v_10467 = v_9903 | v_10466;
assign v_10468 = v_10196 | v_10467;
assign v_10469 = v_10200 | v_10468;
assign v_10470 = v_96 | v_10469;
assign v_10471 = v_807 | v_10470;
assign v_10472 = v_361 | v_10471;
assign v_10481 = v_10479 | v_10480;
assign v_10482 = v_10478 | v_10481;
assign v_10483 = v_10477 | v_10482;
assign v_10484 = v_10476 | v_10483;
assign v_10485 = v_10475 | v_10484;
assign v_10486 = v_10474 | v_10485;
assign v_10487 = v_10473 | v_10486;
assign v_10498 = v_10496 | v_10497;
assign v_10501 = v_10499 | v_10500;
assign v_10504 = v_10502 | v_10503;
assign v_10507 = v_10505 | v_10506;
assign v_10510 = v_10508 | v_10509;
assign v_10513 = v_10511 | v_10512;
assign v_10516 = v_10514 | v_10515;
assign v_10519 = v_10517 | v_10518;
assign v_10522 = v_10520 | v_10521;
assign v_10525 = v_10523 | v_10524;
assign v_10528 = v_10526 | v_10527;
assign v_10531 = v_10529 | v_10530;
assign v_10534 = v_10532 | v_10533;
assign v_10537 = v_10535 | v_10536;
assign v_10540 = v_10538 | v_10539;
assign v_10543 = v_10541 | v_10542;
assign v_10546 = v_10544 | v_10545;
assign v_10549 = v_10547 | v_10548;
assign v_10552 = v_10550 | v_10551;
assign v_10555 = v_10553 | v_10554;
assign v_10558 = v_10556 | v_10557;
assign v_10561 = v_10559 | v_10560;
assign v_10564 = v_10562 | v_10563;
assign v_10567 = v_10565 | v_10566;
assign v_10570 = v_10568 | v_10569;
assign v_10573 = v_10571 | v_10572;
assign v_10576 = v_10574 | v_10575;
assign v_10579 = v_10577 | v_10578;
assign v_10582 = v_10580 | v_10581;
assign v_10585 = v_10583 | v_10584;
assign v_10588 = v_10586 | v_10587;
assign v_10591 = v_10589 | v_10590;
assign v_10594 = v_10592 | v_10593;
assign v_10597 = v_10595 | v_10596;
assign v_10600 = v_10598 | v_10599;
assign v_10603 = v_10601 | v_10602;
assign v_10606 = v_10604 | v_10605;
assign v_10609 = v_10607 | v_10608;
assign v_10612 = v_10610 | v_10611;
assign v_10615 = v_10613 | v_10614;
assign v_10618 = v_10616 | v_10617;
assign v_10621 = v_10619 | v_10620;
assign v_10624 = v_10622 | v_10623;
assign v_10627 = v_10625 | v_10626;
assign v_10630 = v_10628 | v_10629;
assign v_10633 = v_10631 | v_10632;
assign v_10636 = v_10634 | v_10635;
assign v_10639 = v_10637 | v_10638;
assign v_10642 = v_10640 | v_10641;
assign v_10645 = v_10643 | v_10644;
assign v_10648 = v_10646 | v_10647;
assign v_10651 = v_10649 | v_10650;
assign v_10654 = v_10652 | v_10653;
assign v_10657 = v_10655 | v_10656;
assign v_10660 = v_10658 | v_10659;
assign v_10663 = v_10661 | v_10662;
assign v_10666 = v_10664 | v_10665;
assign v_10669 = v_10667 | v_10668;
assign v_10672 = v_10670 | v_10671;
assign v_10675 = v_10673 | v_10674;
assign v_10678 = v_10676 | v_10677;
assign v_10681 = v_10679 | v_10680;
assign v_10684 = v_10682 | v_10683;
assign v_10687 = v_10685 | v_10686;
assign v_10690 = v_10688 | v_10689;
assign v_10693 = v_10691 | v_10692;
assign v_10696 = v_10694 | v_10695;
assign v_10699 = v_10697 | v_10698;
assign v_10702 = v_10700 | v_10701;
assign v_10705 = v_10703 | v_10704;
assign v_10708 = v_10706 | v_10707;
assign v_10711 = v_10709 | v_10710;
assign v_10714 = v_10712 | v_10713;
assign v_10717 = v_10715 | v_10716;
assign v_10720 = v_10718 | v_10719;
assign v_10723 = v_10721 | v_10722;
assign v_10726 = v_10724 | v_10725;
assign v_10729 = v_10727 | v_10728;
assign v_10732 = v_10730 | v_10731;
assign v_10735 = v_10733 | v_10734;
assign v_10738 = v_10736 | v_10737;
assign v_10741 = v_10739 | v_10740;
assign v_10744 = v_10742 | v_10743;
assign v_10747 = v_10745 | v_10746;
assign v_10750 = v_10748 | v_10749;
assign v_10753 = v_10751 | v_10752;
assign v_10756 = v_10754 | v_10755;
assign v_10759 = v_10757 | v_10758;
assign v_10762 = v_10760 | v_10761;
assign v_10765 = v_10763 | v_10764;
assign v_10768 = v_10766 | v_10767;
assign v_10771 = v_10769 | v_10770;
assign v_10774 = v_10772 | v_10773;
assign v_10777 = v_10775 | v_10776;
assign v_10780 = v_10778 | v_10779;
assign v_10783 = v_10781 | v_10782;
assign v_10786 = v_10784 | v_10785;
assign v_10789 = v_10787 | v_10788;
assign v_10792 = v_10790 | v_10791;
assign v_10795 = v_10793 | v_10794;
assign v_10798 = v_10796 | v_10797;
assign v_10801 = v_10799 | v_10800;
assign v_10804 = v_10802 | v_10803;
assign v_10807 = v_10805 | v_10806;
assign v_10810 = v_10808 | v_10809;
assign v_10813 = v_10811 | v_10812;
assign v_10816 = v_10814 | v_10815;
assign v_10819 = v_10817 | v_10818;
assign v_10822 = v_10820 | v_10821;
assign v_10825 = v_10823 | v_10824;
assign v_10828 = v_10826 | v_10827;
assign v_10831 = v_10829 | v_10830;
assign v_10834 = v_10832 | v_10833;
assign v_10837 = v_10835 | v_10836;
assign v_10840 = v_10838 | v_10839;
assign v_10843 = v_10841 | v_10842;
assign v_10846 = v_10844 | v_10845;
assign v_10849 = v_10847 | v_10848;
assign v_10852 = v_10850 | v_10851;
assign v_10855 = v_10853 | v_10854;
assign v_10858 = v_10856 | v_10857;
assign v_10861 = v_10859 | v_10860;
assign v_10864 = v_10862 | v_10863;
assign v_10867 = v_10865 | v_10866;
assign v_10870 = v_10868 | v_10869;
assign v_10873 = v_10871 | v_10872;
assign v_10874 = v_10684 | v_10873;
assign v_10877 = v_10875 | v_10876;
assign v_10880 = v_10878 | v_10879;
assign v_10883 = v_10881 | v_10882;
assign v_10886 = v_10884 | v_10885;
assign v_10889 = v_10887 | v_10888;
assign v_10892 = v_10890 | v_10891;
assign v_10895 = v_10893 | v_10894;
assign v_10898 = v_10896 | v_10897;
assign v_10901 = v_10899 | v_10900;
assign v_10904 = v_10902 | v_10903;
assign v_10907 = v_10905 | v_10906;
assign v_10910 = v_10908 | v_10909;
assign v_10913 = v_10911 | v_10912;
assign v_10916 = v_10914 | v_10915;
assign v_10919 = v_10917 | v_10918;
assign v_10922 = v_10920 | v_10921;
assign v_10925 = v_10923 | v_10924;
assign v_10928 = v_10926 | v_10927;
assign v_10931 = v_10929 | v_10930;
assign v_10934 = v_10932 | v_10933;
assign v_10937 = v_10935 | v_10936;
assign v_10940 = v_10938 | v_10939;
assign v_10943 = v_10941 | v_10942;
assign v_10946 = v_10944 | v_10945;
assign v_10949 = v_10947 | v_10948;
assign v_10952 = v_10950 | v_10951;
assign v_10955 = v_10953 | v_10954;
assign v_10958 = v_10956 | v_10957;
assign v_10961 = v_10959 | v_10960;
assign v_10964 = v_10962 | v_10963;
assign v_10967 = v_10965 | v_10966;
assign v_10970 = v_10968 | v_10969;
assign v_10973 = v_10971 | v_10972;
assign v_10976 = v_10974 | v_10975;
assign v_10979 = v_10977 | v_10978;
assign v_10982 = v_10980 | v_10981;
assign v_10985 = v_10983 | v_10984;
assign v_10988 = v_10986 | v_10987;
assign v_10991 = v_10989 | v_10990;
assign v_10994 = v_10992 | v_10993;
assign v_10997 = v_10995 | v_10996;
assign v_11000 = v_10998 | v_10999;
assign v_11003 = v_11001 | v_11002;
assign v_11006 = v_11004 | v_11005;
assign v_11009 = v_11007 | v_11008;
assign v_11012 = v_11010 | v_11011;
assign v_11015 = v_11013 | v_11014;
assign v_11018 = v_11016 | v_11017;
assign v_11021 = v_11019 | v_11020;
assign v_11024 = v_11022 | v_11023;
assign v_11027 = v_11025 | v_11026;
assign v_11030 = v_11028 | v_11029;
assign v_11033 = v_11031 | v_11032;
assign v_11036 = v_11034 | v_11035;
assign v_11039 = v_11037 | v_11038;
assign v_11042 = v_11040 | v_11041;
assign v_11045 = v_11043 | v_11044;
assign v_11048 = v_11046 | v_11047;
assign v_11051 = v_11049 | v_11050;
assign v_11054 = v_11052 | v_11053;
assign v_11057 = v_11055 | v_11056;
assign v_11060 = v_11058 | v_11059;
assign v_11063 = v_11061 | v_11062;
assign v_11064 = v_10874 | v_11063;
assign v_11067 = v_11065 | v_11066;
assign v_11070 = v_11068 | v_11069;
assign v_11073 = v_11071 | v_11072;
assign v_11076 = v_11074 | v_11075;
assign v_11079 = v_11077 | v_11078;
assign v_11082 = v_11080 | v_11081;
assign v_11085 = v_11083 | v_11084;
assign v_11088 = v_11086 | v_11087;
assign v_11091 = v_11089 | v_11090;
assign v_11094 = v_11092 | v_11093;
assign v_11097 = v_11095 | v_11096;
assign v_11100 = v_11098 | v_11099;
assign v_11103 = v_11101 | v_11102;
assign v_11106 = v_11104 | v_11105;
assign v_11109 = v_11107 | v_11108;
assign v_11112 = v_11110 | v_11111;
assign v_11115 = v_11113 | v_11114;
assign v_11118 = v_11116 | v_11117;
assign v_11121 = v_11119 | v_11120;
assign v_11124 = v_11122 | v_11123;
assign v_11127 = v_11125 | v_11126;
assign v_11130 = v_11128 | v_11129;
assign v_11133 = v_11131 | v_11132;
assign v_11136 = v_11134 | v_11135;
assign v_11139 = v_11137 | v_11138;
assign v_11142 = v_11140 | v_11141;
assign v_11145 = v_11143 | v_11144;
assign v_11148 = v_11146 | v_11147;
assign v_11151 = v_11149 | v_11150;
assign v_11154 = v_11152 | v_11153;
assign v_11157 = v_11155 | v_11156;
assign v_11160 = v_11158 | v_11159;
assign v_11163 = v_11161 | v_11162;
assign v_11166 = v_11164 | v_11165;
assign v_11169 = v_11167 | v_11168;
assign v_11172 = v_11170 | v_11171;
assign v_11175 = v_11173 | v_11174;
assign v_11178 = v_11176 | v_11177;
assign v_11181 = v_11179 | v_11180;
assign v_11184 = v_11182 | v_11183;
assign v_11187 = v_11185 | v_11186;
assign v_11190 = v_11188 | v_11189;
assign v_11193 = v_11191 | v_11192;
assign v_11196 = v_11194 | v_11195;
assign v_11199 = v_11197 | v_11198;
assign v_11202 = v_11200 | v_11201;
assign v_11205 = v_11203 | v_11204;
assign v_11208 = v_11206 | v_11207;
assign v_11211 = v_11209 | v_11210;
assign v_11214 = v_11212 | v_11213;
assign v_11217 = v_11215 | v_11216;
assign v_11220 = v_11218 | v_11219;
assign v_11223 = v_11221 | v_11222;
assign v_11226 = v_11224 | v_11225;
assign v_11229 = v_11227 | v_11228;
assign v_11232 = v_11230 | v_11231;
assign v_11235 = v_11233 | v_11234;
assign v_11238 = v_11236 | v_11237;
assign v_11241 = v_11239 | v_11240;
assign v_11244 = v_11242 | v_11243;
assign v_11247 = v_11245 | v_11246;
assign v_11250 = v_11248 | v_11249;
assign v_11253 = v_11251 | v_11252;
assign v_11254 = v_11064 | v_11253;
assign v_11257 = v_11255 | v_11256;
assign v_11260 = v_11258 | v_11259;
assign v_11263 = v_11261 | v_11262;
assign v_11266 = v_11264 | v_11265;
assign v_11269 = v_11267 | v_11268;
assign v_11272 = v_11270 | v_11271;
assign v_11275 = v_11273 | v_11274;
assign v_11278 = v_11276 | v_11277;
assign v_11281 = v_11279 | v_11280;
assign v_11284 = v_11282 | v_11283;
assign v_11287 = v_11285 | v_11286;
assign v_11290 = v_11288 | v_11289;
assign v_11293 = v_11291 | v_11292;
assign v_11296 = v_11294 | v_11295;
assign v_11299 = v_11297 | v_11298;
assign v_11302 = v_11300 | v_11301;
assign v_11305 = v_11303 | v_11304;
assign v_11308 = v_11306 | v_11307;
assign v_11311 = v_11309 | v_11310;
assign v_11314 = v_11312 | v_11313;
assign v_11317 = v_11315 | v_11316;
assign v_11320 = v_11318 | v_11319;
assign v_11323 = v_11321 | v_11322;
assign v_11326 = v_11324 | v_11325;
assign v_11329 = v_11327 | v_11328;
assign v_11332 = v_11330 | v_11331;
assign v_11335 = v_11333 | v_11334;
assign v_11338 = v_11336 | v_11337;
assign v_11341 = v_11339 | v_11340;
assign v_11344 = v_11342 | v_11343;
assign v_11347 = v_11345 | v_11346;
assign v_11350 = v_11348 | v_11349;
assign v_11353 = v_11351 | v_11352;
assign v_11356 = v_11354 | v_11355;
assign v_11359 = v_11357 | v_11358;
assign v_11362 = v_11360 | v_11361;
assign v_11365 = v_11363 | v_11364;
assign v_11368 = v_11366 | v_11367;
assign v_11371 = v_11369 | v_11370;
assign v_11374 = v_11372 | v_11373;
assign v_11377 = v_11375 | v_11376;
assign v_11380 = v_11378 | v_11379;
assign v_11383 = v_11381 | v_11382;
assign v_11386 = v_11384 | v_11385;
assign v_11389 = v_11387 | v_11388;
assign v_11392 = v_11390 | v_11391;
assign v_11395 = v_11393 | v_11394;
assign v_11398 = v_11396 | v_11397;
assign v_11401 = v_11399 | v_11400;
assign v_11404 = v_11402 | v_11403;
assign v_11407 = v_11405 | v_11406;
assign v_11410 = v_11408 | v_11409;
assign v_11413 = v_11411 | v_11412;
assign v_11416 = v_11414 | v_11415;
assign v_11419 = v_11417 | v_11418;
assign v_11422 = v_11420 | v_11421;
assign v_11425 = v_11423 | v_11424;
assign v_11428 = v_11426 | v_11427;
assign v_11431 = v_11429 | v_11430;
assign v_11434 = v_11432 | v_11433;
assign v_11437 = v_11435 | v_11436;
assign v_11440 = v_11438 | v_11439;
assign v_11443 = v_11441 | v_11442;
assign v_11444 = v_11254 | v_11443;
assign v_11447 = v_11445 | v_11446;
assign v_11450 = v_11448 | v_11449;
assign v_11453 = v_11451 | v_11452;
assign v_11456 = v_11454 | v_11455;
assign v_11459 = v_11457 | v_11458;
assign v_11462 = v_11460 | v_11461;
assign v_11465 = v_11463 | v_11464;
assign v_11468 = v_11466 | v_11467;
assign v_11471 = v_11469 | v_11470;
assign v_11474 = v_11472 | v_11473;
assign v_11477 = v_11475 | v_11476;
assign v_11480 = v_11478 | v_11479;
assign v_11483 = v_11481 | v_11482;
assign v_11486 = v_11484 | v_11485;
assign v_11489 = v_11487 | v_11488;
assign v_11492 = v_11490 | v_11491;
assign v_11495 = v_11493 | v_11494;
assign v_11498 = v_11496 | v_11497;
assign v_11501 = v_11499 | v_11500;
assign v_11504 = v_11502 | v_11503;
assign v_11507 = v_11505 | v_11506;
assign v_11510 = v_11508 | v_11509;
assign v_11513 = v_11511 | v_11512;
assign v_11516 = v_11514 | v_11515;
assign v_11519 = v_11517 | v_11518;
assign v_11522 = v_11520 | v_11521;
assign v_11525 = v_11523 | v_11524;
assign v_11528 = v_11526 | v_11527;
assign v_11531 = v_11529 | v_11530;
assign v_11534 = v_11532 | v_11533;
assign v_11537 = v_11535 | v_11536;
assign v_11540 = v_11538 | v_11539;
assign v_11543 = v_11541 | v_11542;
assign v_11546 = v_11544 | v_11545;
assign v_11549 = v_11547 | v_11548;
assign v_11552 = v_11550 | v_11551;
assign v_11555 = v_11553 | v_11554;
assign v_11558 = v_11556 | v_11557;
assign v_11561 = v_11559 | v_11560;
assign v_11564 = v_11562 | v_11563;
assign v_11567 = v_11565 | v_11566;
assign v_11570 = v_11568 | v_11569;
assign v_11573 = v_11571 | v_11572;
assign v_11576 = v_11574 | v_11575;
assign v_11579 = v_11577 | v_11578;
assign v_11582 = v_11580 | v_11581;
assign v_11585 = v_11583 | v_11584;
assign v_11588 = v_11586 | v_11587;
assign v_11591 = v_11589 | v_11590;
assign v_11594 = v_11592 | v_11593;
assign v_11597 = v_11595 | v_11596;
assign v_11600 = v_11598 | v_11599;
assign v_11603 = v_11601 | v_11602;
assign v_11606 = v_11604 | v_11605;
assign v_11609 = v_11607 | v_11608;
assign v_11612 = v_11610 | v_11611;
assign v_11615 = v_11613 | v_11614;
assign v_11618 = v_11616 | v_11617;
assign v_11621 = v_11619 | v_11620;
assign v_11624 = v_11622 | v_11623;
assign v_11627 = v_11625 | v_11626;
assign v_11630 = v_11628 | v_11629;
assign v_11633 = v_11631 | v_11632;
assign v_11634 = v_11444 | v_11633;
assign v_11637 = v_11635 | v_11636;
assign v_11640 = v_11638 | v_11639;
assign v_11643 = v_11641 | v_11642;
assign v_11646 = v_11644 | v_11645;
assign v_11649 = v_11647 | v_11648;
assign v_11652 = v_11650 | v_11651;
assign v_11655 = v_11653 | v_11654;
assign v_11658 = v_11656 | v_11657;
assign v_11661 = v_11659 | v_11660;
assign v_11664 = v_11662 | v_11663;
assign v_11667 = v_11665 | v_11666;
assign v_11670 = v_11668 | v_11669;
assign v_11673 = v_11671 | v_11672;
assign v_11676 = v_11674 | v_11675;
assign v_11679 = v_11677 | v_11678;
assign v_11682 = v_11680 | v_11681;
assign v_11685 = v_11683 | v_11684;
assign v_11688 = v_11686 | v_11687;
assign v_11691 = v_11689 | v_11690;
assign v_11694 = v_11692 | v_11693;
assign v_11697 = v_11695 | v_11696;
assign v_11700 = v_11698 | v_11699;
assign v_11703 = v_11701 | v_11702;
assign v_11706 = v_11704 | v_11705;
assign v_11709 = v_11707 | v_11708;
assign v_11712 = v_11710 | v_11711;
assign v_11715 = v_11713 | v_11714;
assign v_11718 = v_11716 | v_11717;
assign v_11721 = v_11719 | v_11720;
assign v_11724 = v_11722 | v_11723;
assign v_11727 = v_11725 | v_11726;
assign v_11730 = v_11728 | v_11729;
assign v_11733 = v_11731 | v_11732;
assign v_11736 = v_11734 | v_11735;
assign v_11739 = v_11737 | v_11738;
assign v_11742 = v_11740 | v_11741;
assign v_11745 = v_11743 | v_11744;
assign v_11748 = v_11746 | v_11747;
assign v_11751 = v_11749 | v_11750;
assign v_11754 = v_11752 | v_11753;
assign v_11757 = v_11755 | v_11756;
assign v_11760 = v_11758 | v_11759;
assign v_11763 = v_11761 | v_11762;
assign v_11766 = v_11764 | v_11765;
assign v_11769 = v_11767 | v_11768;
assign v_11772 = v_11770 | v_11771;
assign v_11775 = v_11773 | v_11774;
assign v_11778 = v_11776 | v_11777;
assign v_11781 = v_11779 | v_11780;
assign v_11784 = v_11782 | v_11783;
assign v_11787 = v_11785 | v_11786;
assign v_11790 = v_11788 | v_11789;
assign v_11793 = v_11791 | v_11792;
assign v_11796 = v_11794 | v_11795;
assign v_11799 = v_11797 | v_11798;
assign v_11802 = v_11800 | v_11801;
assign v_11805 = v_11803 | v_11804;
assign v_11808 = v_11806 | v_11807;
assign v_11811 = v_11809 | v_11810;
assign v_11814 = v_11812 | v_11813;
assign v_11817 = v_11815 | v_11816;
assign v_11820 = v_11818 | v_11819;
assign v_11823 = v_11821 | v_11822;
assign v_11824 = v_11634 | v_11823;
assign v_11827 = v_11825 | v_11826;
assign v_11830 = v_11828 | v_11829;
assign v_11833 = v_11831 | v_11832;
assign v_11836 = v_11834 | v_11835;
assign v_11839 = v_11837 | v_11838;
assign v_11842 = v_11840 | v_11841;
assign v_11845 = v_11843 | v_11844;
assign v_11848 = v_11846 | v_11847;
assign v_11851 = v_11849 | v_11850;
assign v_11854 = v_11852 | v_11853;
assign v_11857 = v_11855 | v_11856;
assign v_11860 = v_11858 | v_11859;
assign v_11863 = v_11861 | v_11862;
assign v_11866 = v_11864 | v_11865;
assign v_11869 = v_11867 | v_11868;
assign v_11872 = v_11870 | v_11871;
assign v_11875 = v_11873 | v_11874;
assign v_11878 = v_11876 | v_11877;
assign v_11881 = v_11879 | v_11880;
assign v_11884 = v_11882 | v_11883;
assign v_11887 = v_11885 | v_11886;
assign v_11890 = v_11888 | v_11889;
assign v_11893 = v_11891 | v_11892;
assign v_11896 = v_11894 | v_11895;
assign v_11899 = v_11897 | v_11898;
assign v_11902 = v_11900 | v_11901;
assign v_11905 = v_11903 | v_11904;
assign v_11908 = v_11906 | v_11907;
assign v_11911 = v_11909 | v_11910;
assign v_11914 = v_11912 | v_11913;
assign v_11917 = v_11915 | v_11916;
assign v_11920 = v_11918 | v_11919;
assign v_11923 = v_11921 | v_11922;
assign v_11926 = v_11924 | v_11925;
assign v_11929 = v_11927 | v_11928;
assign v_11932 = v_11930 | v_11931;
assign v_11935 = v_11933 | v_11934;
assign v_11938 = v_11936 | v_11937;
assign v_11941 = v_11939 | v_11940;
assign v_11944 = v_11942 | v_11943;
assign v_11947 = v_11945 | v_11946;
assign v_11950 = v_11948 | v_11949;
assign v_11953 = v_11951 | v_11952;
assign v_11956 = v_11954 | v_11955;
assign v_11959 = v_11957 | v_11958;
assign v_11962 = v_11960 | v_11961;
assign v_11965 = v_11963 | v_11964;
assign v_11968 = v_11966 | v_11967;
assign v_11971 = v_11969 | v_11970;
assign v_11974 = v_11972 | v_11973;
assign v_11977 = v_11975 | v_11976;
assign v_11980 = v_11978 | v_11979;
assign v_11983 = v_11981 | v_11982;
assign v_11986 = v_11984 | v_11985;
assign v_11989 = v_11987 | v_11988;
assign v_11992 = v_11990 | v_11991;
assign v_11995 = v_11993 | v_11994;
assign v_11998 = v_11996 | v_11997;
assign v_12001 = v_11999 | v_12000;
assign v_12004 = v_12002 | v_12003;
assign v_12007 = v_12005 | v_12006;
assign v_12010 = v_12008 | v_12009;
assign v_12013 = v_12011 | v_12012;
assign v_12014 = v_11824 | v_12013;
assign v_12017 = v_12015 | v_12016;
assign v_12020 = v_12018 | v_12019;
assign v_12023 = v_12021 | v_12022;
assign v_12026 = v_12024 | v_12025;
assign v_12029 = v_12027 | v_12028;
assign v_12032 = v_12030 | v_12031;
assign v_12035 = v_12033 | v_12034;
assign v_12038 = v_12036 | v_12037;
assign v_12041 = v_12039 | v_12040;
assign v_12044 = v_12042 | v_12043;
assign v_12047 = v_12045 | v_12046;
assign v_12050 = v_12048 | v_12049;
assign v_12053 = v_12051 | v_12052;
assign v_12056 = v_12054 | v_12055;
assign v_12059 = v_12057 | v_12058;
assign v_12062 = v_12060 | v_12061;
assign v_12065 = v_12063 | v_12064;
assign v_12068 = v_12066 | v_12067;
assign v_12071 = v_12069 | v_12070;
assign v_12074 = v_12072 | v_12073;
assign v_12077 = v_12075 | v_12076;
assign v_12080 = v_12078 | v_12079;
assign v_12083 = v_12081 | v_12082;
assign v_12086 = v_12084 | v_12085;
assign v_12089 = v_12087 | v_12088;
assign v_12092 = v_12090 | v_12091;
assign v_12095 = v_12093 | v_12094;
assign v_12098 = v_12096 | v_12097;
assign v_12101 = v_12099 | v_12100;
assign v_12104 = v_12102 | v_12103;
assign v_12107 = v_12105 | v_12106;
assign v_12110 = v_12108 | v_12109;
assign v_12113 = v_12111 | v_12112;
assign v_12116 = v_12114 | v_12115;
assign v_12119 = v_12117 | v_12118;
assign v_12122 = v_12120 | v_12121;
assign v_12125 = v_12123 | v_12124;
assign v_12128 = v_12126 | v_12127;
assign v_12131 = v_12129 | v_12130;
assign v_12134 = v_12132 | v_12133;
assign v_12137 = v_12135 | v_12136;
assign v_12140 = v_12138 | v_12139;
assign v_12143 = v_12141 | v_12142;
assign v_12146 = v_12144 | v_12145;
assign v_12149 = v_12147 | v_12148;
assign v_12152 = v_12150 | v_12151;
assign v_12155 = v_12153 | v_12154;
assign v_12158 = v_12156 | v_12157;
assign v_12161 = v_12159 | v_12160;
assign v_12164 = v_12162 | v_12163;
assign v_12167 = v_12165 | v_12166;
assign v_12170 = v_12168 | v_12169;
assign v_12173 = v_12171 | v_12172;
assign v_12176 = v_12174 | v_12175;
assign v_12179 = v_12177 | v_12178;
assign v_12182 = v_12180 | v_12181;
assign v_12185 = v_12183 | v_12184;
assign v_12188 = v_12186 | v_12187;
assign v_12191 = v_12189 | v_12190;
assign v_12194 = v_12192 | v_12193;
assign v_12197 = v_12195 | v_12196;
assign v_12200 = v_12198 | v_12199;
assign v_12203 = v_12201 | v_12202;
assign v_12206 = v_12204 | v_12205;
assign v_12209 = v_12207 | v_12208;
assign v_12212 = v_12210 | v_12211;
assign v_12215 = v_12213 | v_12214;
assign v_12218 = v_12216 | v_12217;
assign v_12221 = v_12219 | v_12220;
assign v_12224 = v_12222 | v_12223;
assign v_12227 = v_12225 | v_12226;
assign v_12230 = v_12228 | v_12229;
assign v_12233 = v_12231 | v_12232;
assign v_12236 = v_12234 | v_12235;
assign v_12239 = v_12237 | v_12238;
assign v_12242 = v_12240 | v_12241;
assign v_12245 = v_12243 | v_12244;
assign v_12248 = v_12246 | v_12247;
assign v_12251 = v_12249 | v_12250;
assign v_12254 = v_12252 | v_12253;
assign v_12257 = v_12255 | v_12256;
assign v_12260 = v_12258 | v_12259;
assign v_12263 = v_12261 | v_12262;
assign v_12266 = v_12264 | v_12265;
assign v_12269 = v_12267 | v_12268;
assign v_12272 = v_12270 | v_12271;
assign v_12275 = v_12273 | v_12274;
assign v_12278 = v_12276 | v_12277;
assign v_12281 = v_12279 | v_12280;
assign v_12284 = v_12282 | v_12283;
assign v_12287 = v_12285 | v_12286;
assign v_12290 = v_12288 | v_12289;
assign v_12293 = v_12291 | v_12292;
assign v_12296 = v_12294 | v_12295;
assign v_12299 = v_12297 | v_12298;
assign v_12302 = v_12300 | v_12301;
assign v_12305 = v_12303 | v_12304;
assign v_12308 = v_12306 | v_12307;
assign v_12311 = v_12309 | v_12310;
assign v_12314 = v_12312 | v_12313;
assign v_12317 = v_12315 | v_12316;
assign v_12320 = v_12318 | v_12319;
assign v_12323 = v_12321 | v_12322;
assign v_12326 = v_12324 | v_12325;
assign v_12329 = v_12327 | v_12328;
assign v_12332 = v_12330 | v_12331;
assign v_12335 = v_12333 | v_12334;
assign v_12338 = v_12336 | v_12337;
assign v_12341 = v_12339 | v_12340;
assign v_12344 = v_12342 | v_12343;
assign v_12347 = v_12345 | v_12346;
assign v_12350 = v_12348 | v_12349;
assign v_12353 = v_12351 | v_12352;
assign v_12356 = v_12354 | v_12355;
assign v_12359 = v_12357 | v_12358;
assign v_12362 = v_12360 | v_12361;
assign v_12365 = v_12363 | v_12364;
assign v_12368 = v_12366 | v_12367;
assign v_12371 = v_12369 | v_12370;
assign v_12374 = v_12372 | v_12373;
assign v_12377 = v_12375 | v_12376;
assign v_12380 = v_12378 | v_12379;
assign v_12383 = v_12381 | v_12382;
assign v_12386 = v_12384 | v_12385;
assign v_12389 = v_12387 | v_12388;
assign v_12392 = v_12390 | v_12391;
assign v_12393 = v_12203 | v_12392;
assign v_12396 = v_12394 | v_12395;
assign v_12399 = v_12397 | v_12398;
assign v_12402 = v_12400 | v_12401;
assign v_12405 = v_12403 | v_12404;
assign v_12408 = v_12406 | v_12407;
assign v_12411 = v_12409 | v_12410;
assign v_12414 = v_12412 | v_12413;
assign v_12417 = v_12415 | v_12416;
assign v_12420 = v_12418 | v_12419;
assign v_12423 = v_12421 | v_12422;
assign v_12426 = v_12424 | v_12425;
assign v_12429 = v_12427 | v_12428;
assign v_12432 = v_12430 | v_12431;
assign v_12435 = v_12433 | v_12434;
assign v_12438 = v_12436 | v_12437;
assign v_12441 = v_12439 | v_12440;
assign v_12444 = v_12442 | v_12443;
assign v_12447 = v_12445 | v_12446;
assign v_12450 = v_12448 | v_12449;
assign v_12453 = v_12451 | v_12452;
assign v_12456 = v_12454 | v_12455;
assign v_12459 = v_12457 | v_12458;
assign v_12462 = v_12460 | v_12461;
assign v_12465 = v_12463 | v_12464;
assign v_12468 = v_12466 | v_12467;
assign v_12471 = v_12469 | v_12470;
assign v_12474 = v_12472 | v_12473;
assign v_12477 = v_12475 | v_12476;
assign v_12480 = v_12478 | v_12479;
assign v_12483 = v_12481 | v_12482;
assign v_12486 = v_12484 | v_12485;
assign v_12489 = v_12487 | v_12488;
assign v_12492 = v_12490 | v_12491;
assign v_12495 = v_12493 | v_12494;
assign v_12498 = v_12496 | v_12497;
assign v_12501 = v_12499 | v_12500;
assign v_12504 = v_12502 | v_12503;
assign v_12507 = v_12505 | v_12506;
assign v_12510 = v_12508 | v_12509;
assign v_12513 = v_12511 | v_12512;
assign v_12516 = v_12514 | v_12515;
assign v_12519 = v_12517 | v_12518;
assign v_12522 = v_12520 | v_12521;
assign v_12525 = v_12523 | v_12524;
assign v_12528 = v_12526 | v_12527;
assign v_12531 = v_12529 | v_12530;
assign v_12534 = v_12532 | v_12533;
assign v_12537 = v_12535 | v_12536;
assign v_12540 = v_12538 | v_12539;
assign v_12543 = v_12541 | v_12542;
assign v_12546 = v_12544 | v_12545;
assign v_12549 = v_12547 | v_12548;
assign v_12552 = v_12550 | v_12551;
assign v_12555 = v_12553 | v_12554;
assign v_12558 = v_12556 | v_12557;
assign v_12561 = v_12559 | v_12560;
assign v_12564 = v_12562 | v_12563;
assign v_12567 = v_12565 | v_12566;
assign v_12570 = v_12568 | v_12569;
assign v_12573 = v_12571 | v_12572;
assign v_12576 = v_12574 | v_12575;
assign v_12579 = v_12577 | v_12578;
assign v_12582 = v_12580 | v_12581;
assign v_12583 = v_12393 | v_12582;
assign v_12586 = v_12584 | v_12585;
assign v_12589 = v_12587 | v_12588;
assign v_12592 = v_12590 | v_12591;
assign v_12595 = v_12593 | v_12594;
assign v_12598 = v_12596 | v_12597;
assign v_12601 = v_12599 | v_12600;
assign v_12604 = v_12602 | v_12603;
assign v_12607 = v_12605 | v_12606;
assign v_12610 = v_12608 | v_12609;
assign v_12613 = v_12611 | v_12612;
assign v_12616 = v_12614 | v_12615;
assign v_12619 = v_12617 | v_12618;
assign v_12622 = v_12620 | v_12621;
assign v_12625 = v_12623 | v_12624;
assign v_12628 = v_12626 | v_12627;
assign v_12631 = v_12629 | v_12630;
assign v_12634 = v_12632 | v_12633;
assign v_12637 = v_12635 | v_12636;
assign v_12640 = v_12638 | v_12639;
assign v_12643 = v_12641 | v_12642;
assign v_12646 = v_12644 | v_12645;
assign v_12649 = v_12647 | v_12648;
assign v_12652 = v_12650 | v_12651;
assign v_12655 = v_12653 | v_12654;
assign v_12658 = v_12656 | v_12657;
assign v_12661 = v_12659 | v_12660;
assign v_12664 = v_12662 | v_12663;
assign v_12667 = v_12665 | v_12666;
assign v_12670 = v_12668 | v_12669;
assign v_12673 = v_12671 | v_12672;
assign v_12676 = v_12674 | v_12675;
assign v_12679 = v_12677 | v_12678;
assign v_12682 = v_12680 | v_12681;
assign v_12685 = v_12683 | v_12684;
assign v_12688 = v_12686 | v_12687;
assign v_12691 = v_12689 | v_12690;
assign v_12694 = v_12692 | v_12693;
assign v_12697 = v_12695 | v_12696;
assign v_12700 = v_12698 | v_12699;
assign v_12703 = v_12701 | v_12702;
assign v_12706 = v_12704 | v_12705;
assign v_12709 = v_12707 | v_12708;
assign v_12712 = v_12710 | v_12711;
assign v_12715 = v_12713 | v_12714;
assign v_12718 = v_12716 | v_12717;
assign v_12721 = v_12719 | v_12720;
assign v_12724 = v_12722 | v_12723;
assign v_12727 = v_12725 | v_12726;
assign v_12730 = v_12728 | v_12729;
assign v_12733 = v_12731 | v_12732;
assign v_12736 = v_12734 | v_12735;
assign v_12739 = v_12737 | v_12738;
assign v_12742 = v_12740 | v_12741;
assign v_12745 = v_12743 | v_12744;
assign v_12748 = v_12746 | v_12747;
assign v_12751 = v_12749 | v_12750;
assign v_12754 = v_12752 | v_12753;
assign v_12757 = v_12755 | v_12756;
assign v_12760 = v_12758 | v_12759;
assign v_12763 = v_12761 | v_12762;
assign v_12766 = v_12764 | v_12765;
assign v_12769 = v_12767 | v_12768;
assign v_12772 = v_12770 | v_12771;
assign v_12773 = v_12583 | v_12772;
assign v_12776 = v_12774 | v_12775;
assign v_12779 = v_12777 | v_12778;
assign v_12782 = v_12780 | v_12781;
assign v_12785 = v_12783 | v_12784;
assign v_12788 = v_12786 | v_12787;
assign v_12791 = v_12789 | v_12790;
assign v_12794 = v_12792 | v_12793;
assign v_12797 = v_12795 | v_12796;
assign v_12800 = v_12798 | v_12799;
assign v_12803 = v_12801 | v_12802;
assign v_12806 = v_12804 | v_12805;
assign v_12809 = v_12807 | v_12808;
assign v_12812 = v_12810 | v_12811;
assign v_12815 = v_12813 | v_12814;
assign v_12818 = v_12816 | v_12817;
assign v_12821 = v_12819 | v_12820;
assign v_12824 = v_12822 | v_12823;
assign v_12827 = v_12825 | v_12826;
assign v_12830 = v_12828 | v_12829;
assign v_12833 = v_12831 | v_12832;
assign v_12836 = v_12834 | v_12835;
assign v_12839 = v_12837 | v_12838;
assign v_12842 = v_12840 | v_12841;
assign v_12845 = v_12843 | v_12844;
assign v_12848 = v_12846 | v_12847;
assign v_12851 = v_12849 | v_12850;
assign v_12854 = v_12852 | v_12853;
assign v_12857 = v_12855 | v_12856;
assign v_12860 = v_12858 | v_12859;
assign v_12863 = v_12861 | v_12862;
assign v_12866 = v_12864 | v_12865;
assign v_12869 = v_12867 | v_12868;
assign v_12872 = v_12870 | v_12871;
assign v_12875 = v_12873 | v_12874;
assign v_12878 = v_12876 | v_12877;
assign v_12881 = v_12879 | v_12880;
assign v_12884 = v_12882 | v_12883;
assign v_12887 = v_12885 | v_12886;
assign v_12890 = v_12888 | v_12889;
assign v_12893 = v_12891 | v_12892;
assign v_12896 = v_12894 | v_12895;
assign v_12899 = v_12897 | v_12898;
assign v_12902 = v_12900 | v_12901;
assign v_12905 = v_12903 | v_12904;
assign v_12908 = v_12906 | v_12907;
assign v_12911 = v_12909 | v_12910;
assign v_12914 = v_12912 | v_12913;
assign v_12917 = v_12915 | v_12916;
assign v_12920 = v_12918 | v_12919;
assign v_12923 = v_12921 | v_12922;
assign v_12926 = v_12924 | v_12925;
assign v_12929 = v_12927 | v_12928;
assign v_12932 = v_12930 | v_12931;
assign v_12935 = v_12933 | v_12934;
assign v_12938 = v_12936 | v_12937;
assign v_12941 = v_12939 | v_12940;
assign v_12944 = v_12942 | v_12943;
assign v_12947 = v_12945 | v_12946;
assign v_12950 = v_12948 | v_12949;
assign v_12953 = v_12951 | v_12952;
assign v_12956 = v_12954 | v_12955;
assign v_12959 = v_12957 | v_12958;
assign v_12962 = v_12960 | v_12961;
assign v_12963 = v_12773 | v_12962;
assign v_12966 = v_12964 | v_12965;
assign v_12969 = v_12967 | v_12968;
assign v_12972 = v_12970 | v_12971;
assign v_12975 = v_12973 | v_12974;
assign v_12978 = v_12976 | v_12977;
assign v_12981 = v_12979 | v_12980;
assign v_12984 = v_12982 | v_12983;
assign v_12987 = v_12985 | v_12986;
assign v_12990 = v_12988 | v_12989;
assign v_12993 = v_12991 | v_12992;
assign v_12996 = v_12994 | v_12995;
assign v_12999 = v_12997 | v_12998;
assign v_13002 = v_13000 | v_13001;
assign v_13005 = v_13003 | v_13004;
assign v_13008 = v_13006 | v_13007;
assign v_13011 = v_13009 | v_13010;
assign v_13014 = v_13012 | v_13013;
assign v_13017 = v_13015 | v_13016;
assign v_13020 = v_13018 | v_13019;
assign v_13023 = v_13021 | v_13022;
assign v_13026 = v_13024 | v_13025;
assign v_13029 = v_13027 | v_13028;
assign v_13032 = v_13030 | v_13031;
assign v_13035 = v_13033 | v_13034;
assign v_13038 = v_13036 | v_13037;
assign v_13041 = v_13039 | v_13040;
assign v_13044 = v_13042 | v_13043;
assign v_13047 = v_13045 | v_13046;
assign v_13050 = v_13048 | v_13049;
assign v_13053 = v_13051 | v_13052;
assign v_13056 = v_13054 | v_13055;
assign v_13059 = v_13057 | v_13058;
assign v_13062 = v_13060 | v_13061;
assign v_13065 = v_13063 | v_13064;
assign v_13068 = v_13066 | v_13067;
assign v_13071 = v_13069 | v_13070;
assign v_13074 = v_13072 | v_13073;
assign v_13077 = v_13075 | v_13076;
assign v_13080 = v_13078 | v_13079;
assign v_13083 = v_13081 | v_13082;
assign v_13086 = v_13084 | v_13085;
assign v_13089 = v_13087 | v_13088;
assign v_13092 = v_13090 | v_13091;
assign v_13095 = v_13093 | v_13094;
assign v_13098 = v_13096 | v_13097;
assign v_13101 = v_13099 | v_13100;
assign v_13104 = v_13102 | v_13103;
assign v_13107 = v_13105 | v_13106;
assign v_13110 = v_13108 | v_13109;
assign v_13113 = v_13111 | v_13112;
assign v_13116 = v_13114 | v_13115;
assign v_13119 = v_13117 | v_13118;
assign v_13122 = v_13120 | v_13121;
assign v_13125 = v_13123 | v_13124;
assign v_13128 = v_13126 | v_13127;
assign v_13131 = v_13129 | v_13130;
assign v_13134 = v_13132 | v_13133;
assign v_13137 = v_13135 | v_13136;
assign v_13140 = v_13138 | v_13139;
assign v_13143 = v_13141 | v_13142;
assign v_13146 = v_13144 | v_13145;
assign v_13149 = v_13147 | v_13148;
assign v_13152 = v_13150 | v_13151;
assign v_13153 = v_12963 | v_13152;
assign v_13154 = v_9646 | ~v_9844;
assign v_13155 = v_9618 | ~v_9712;
assign v_13157 = v_9488 | v_13156;
assign v_13158 = v_9473 | ~v_9554;
assign v_13160 = v_9356 | v_13159;
assign v_13161 = v_9329 | ~v_9422;
assign v_13163 = v_9200 | v_13162;
assign v_13164 = v_9185 | ~v_9266;
assign v_13166 = v_9068 | v_13165;
assign v_13167 = v_9044 | ~v_9134;
assign v_13169 = v_8918 | v_13168;
assign v_13170 = v_8903 | ~v_8984;
assign v_13172 = v_8786 | v_13171;
assign v_13173 = v_8755 | ~v_8852;
assign v_13175 = v_8622 | v_13174;
assign v_13176 = v_8607 | ~v_8688;
assign v_13178 = v_8490 | v_13177;
assign v_13179 = v_8465 | ~v_8556;
assign v_13181 = v_8338 | v_13180;
assign v_13182 = v_8323 | ~v_8404;
assign v_13184 = v_8206 | v_13183;
assign v_13185 = v_8179 | ~v_8272;
assign v_13187 = v_8050 | v_13186;
assign v_13188 = v_8035 | ~v_8116;
assign v_13190 = v_7918 | v_13189;
assign v_13191 = v_7894 | ~v_7984;
assign v_13193 = v_7768 | v_13192;
assign v_13194 = v_7753 | ~v_7834;
assign v_13196 = v_7636 | v_13195;
assign v_13197 = v_7601 | ~v_7702;
assign v_13199 = v_7464 | v_13198;
assign v_13200 = v_7449 | ~v_7530;
assign v_13202 = v_7332 | v_13201;
assign v_13203 = v_7306 | ~v_7398;
assign v_13205 = v_7178 | v_13204;
assign v_13206 = v_7163 | ~v_7244;
assign v_13208 = v_7046 | v_13207;
assign v_13209 = v_7019 | ~v_7112;
assign v_13211 = v_6890 | v_13210;
assign v_13212 = v_6875 | ~v_6956;
assign v_13214 = v_6758 | v_13213;
assign v_13215 = v_6734 | v_6824;
assign v_13217 = v_6608 | v_13216;
assign v_13218 = v_6593 | ~v_6674;
assign v_13220 = v_6476 | v_13219;
assign v_13221 = v_6445 | ~v_6542;
assign v_13223 = v_6312 | v_13222;
assign v_13224 = v_6297 | ~v_6378;
assign v_13226 = v_6180 | v_13225;
assign v_13227 = v_6155 | ~v_6246;
assign v_13229 = v_6028 | v_13228;
assign v_13230 = v_6013 | v_6094;
assign v_13232 = v_5896 | v_13231;
assign v_13233 = v_5869 | ~v_5962;
assign v_13235 = v_5740 | v_13234;
assign v_13236 = v_5725 | v_5806;
assign v_13238 = v_5608 | v_13237;
assign v_13239 = v_5584 | ~v_5674;
assign v_13241 = v_5458 | v_13240;
assign v_13242 = v_5443 | ~v_5524;
assign v_13244 = v_5326 | v_13243;
assign v_13245 = v_5287 | ~v_5392;
assign v_13247 = v_5146 | v_13246;
assign v_13248 = v_5131 | ~v_5212;
assign v_13250 = v_5014 | v_13249;
assign v_13251 = v_4987 | ~v_5080;
assign v_13253 = v_4858 | v_13252;
assign v_13254 = v_4843 | ~v_4924;
assign v_13256 = v_4726 | v_13255;
assign v_13257 = v_4699 | ~v_4792;
assign v_13259 = v_4570 | v_13258;
assign v_13260 = v_4555 | ~v_4636;
assign v_13262 = v_4438 | v_13261;
assign v_13263 = v_4414 | ~v_4504;
assign v_13265 = v_4288 | v_13264;
assign v_13266 = v_4273 | ~v_4354;
assign v_13268 = v_4156 | v_13267;
assign v_13269 = v_4125 | ~v_4222;
assign v_13271 = v_3992 | v_13270;
assign v_13272 = v_3977 | ~v_4058;
assign v_13274 = v_3860 | v_13273;
assign v_13275 = v_3835 | ~v_3926;
assign v_13277 = v_3708 | v_13276;
assign v_13278 = v_3693 | ~v_3774;
assign v_13280 = v_3576 | v_13279;
assign v_13281 = v_3549 | ~v_3642;
assign v_13283 = v_3420 | v_13282;
assign v_13284 = v_3405 | ~v_3486;
assign v_13286 = v_3288 | v_13285;
assign v_13287 = v_3264 | ~v_3354;
assign v_13289 = v_3138 | v_13288;
assign v_13290 = v_3123 | v_3204;
assign v_13292 = v_3006 | v_13291;
assign v_13293 = v_2971 | ~v_3072;
assign v_13295 = v_2834 | v_13294;
assign v_13296 = v_2819 | ~v_2900;
assign v_13298 = v_2702 | v_13297;
assign v_13299 = v_2676 | ~v_2768;
assign v_13301 = v_2548 | v_13300;
assign v_13302 = v_2533 | ~v_2614;
assign v_13304 = v_2416 | v_13303;
assign v_13305 = v_2389 | ~v_2482;
assign v_13307 = v_2260 | v_13306;
assign v_13308 = v_2245 | ~v_2326;
assign v_13310 = v_2128 | v_13309;
assign v_13311 = v_2104 | ~v_2194;
assign v_13313 = v_1978 | v_13312;
assign v_13314 = v_1963 | ~v_2044;
assign v_13316 = v_1846 | v_13315;
assign v_13317 = v_1815 | ~v_1912;
assign v_13319 = v_1682 | v_13318;
assign v_13320 = v_1667 | ~v_1748;
assign v_13322 = v_1550 | v_13321;
assign v_13323 = v_1525 | ~v_1616;
assign v_13325 = v_1398 | v_13324;
assign v_13326 = v_1383 | ~v_1464;
assign v_13328 = v_1266 | v_13327;
assign v_13329 = v_1239 | ~v_1332;
assign v_13331 = v_1110 | v_13330;
assign v_13332 = v_1095 | ~v_1176;
assign v_13334 = v_978 | v_13333;
assign v_13335 = v_954 | ~v_1044;
assign v_13337 = v_832 | v_13336;
assign v_13338 = v_816 | ~v_898;
assign v_13340 = v_715 | v_13339;
assign v_13341 = v_561 | ~v_771;
assign v_13343 = v_13153 | v_13342;
assign v_13346 = v_13344 | v_13345;
assign v_13349 = v_13347 | v_13348;
assign v_13352 = v_13350 | v_13351;
assign v_13355 = v_13353 | v_13354;
assign v_13358 = v_13356 | v_13357;
assign v_13361 = v_13359 | v_13360;
assign v_13364 = v_13362 | v_13363;
assign v_13367 = v_13365 | v_13366;
assign v_13370 = v_13368 | v_13369;
assign v_13373 = v_13371 | v_13372;
assign v_13376 = v_13374 | v_13375;
assign v_13379 = v_13377 | v_13378;
assign v_13382 = v_13380 | v_13381;
assign v_13385 = v_13383 | v_13384;
assign v_13388 = v_13386 | v_13387;
assign v_13391 = v_13389 | v_13390;
assign v_13394 = v_13392 | v_13393;
assign v_13397 = v_13395 | v_13396;
assign v_13400 = v_13398 | v_13399;
assign v_13403 = v_13401 | v_13402;
assign v_13406 = v_13404 | v_13405;
assign v_13409 = v_13407 | v_13408;
assign v_13412 = v_13410 | v_13411;
assign v_13415 = v_13413 | v_13414;
assign v_13418 = v_13416 | v_13417;
assign v_13421 = v_13419 | v_13420;
assign v_13424 = v_13422 | v_13423;
assign v_13427 = v_13425 | v_13426;
assign v_13430 = v_13428 | v_13429;
assign v_13433 = v_13431 | v_13432;
assign v_13436 = v_13434 | v_13435;
assign v_13439 = v_13437 | v_13438;
assign v_13442 = v_13440 | v_13441;
assign v_13445 = v_13443 | v_13444;
assign v_13448 = v_13446 | v_13447;
assign v_13451 = v_13449 | v_13450;
assign v_13454 = v_13452 | v_13453;
assign v_13457 = v_13455 | v_13456;
assign v_13460 = v_13458 | v_13459;
assign v_13463 = v_13461 | v_13462;
assign v_13466 = v_13464 | v_13465;
assign v_13469 = v_13467 | v_13468;
assign v_13472 = v_13470 | v_13471;
assign v_13475 = v_13473 | v_13474;
assign v_13478 = v_13476 | v_13477;
assign v_13481 = v_13479 | v_13480;
assign v_13484 = v_13482 | v_13483;
assign v_13487 = v_13485 | v_13486;
assign v_13490 = v_13488 | v_13489;
assign v_13493 = v_13491 | v_13492;
assign v_13496 = v_13494 | v_13495;
assign v_13499 = v_13497 | v_13498;
assign v_13502 = v_13500 | v_13501;
assign v_13505 = v_13503 | v_13504;
assign v_13508 = v_13506 | v_13507;
assign v_13511 = v_13509 | v_13510;
assign v_13514 = v_13512 | v_13513;
assign v_13517 = v_13515 | v_13516;
assign v_13520 = v_13518 | v_13519;
assign v_13523 = v_13521 | v_13522;
assign v_13526 = v_13524 | v_13525;
assign v_13529 = v_13527 | v_13528;
assign v_13532 = v_13530 | v_13531;
assign v_13533 = v_13343 | v_13532;
assign v_13534 = v_10414 | v_10421;
assign v_13535 = v_10427 | v_13534;
assign v_13536 = v_10433 | v_13535;
assign v_13537 = v_10439 | v_13536;
assign v_13538 = v_10445 | v_13537;
assign v_13539 = v_10451 | v_13538;
assign v_13540 = v_4 | v_13539;
assign v_13541 = v_13533 | v_13540;
assign v_13542 = v_12014 | v_13541;
assign v_13543 = v_10462 | v_13542;
assign v_13547 = v_13545 | v_13546;
assign v_13550 = v_13548 | v_13549;
assign v_13553 = v_13551 | v_13552;
assign v_13556 = v_13554 | v_13555;
assign v_13559 = v_13557 | v_13558;
assign v_13562 = v_13560 | v_13561;
assign v_13565 = v_13563 | v_13564;
assign v_13568 = v_13566 | v_13567;
assign v_13571 = v_13569 | v_13570;
assign v_13574 = v_13572 | v_13573;
assign v_13577 = v_13575 | v_13576;
assign v_13580 = v_13578 | v_13579;
assign v_13583 = v_13581 | v_13582;
assign v_13586 = v_13584 | v_13585;
assign v_13589 = v_13587 | v_13588;
assign v_13592 = v_13590 | v_13591;
assign v_13595 = v_13593 | v_13594;
assign v_13598 = v_13596 | v_13597;
assign v_13601 = v_13599 | v_13600;
assign v_13604 = v_13602 | v_13603;
assign v_13607 = v_13605 | v_13606;
assign v_13610 = v_13608 | v_13609;
assign v_13613 = v_13611 | v_13612;
assign v_13616 = v_13614 | v_13615;
assign v_13619 = v_13617 | v_13618;
assign v_13622 = v_13620 | v_13621;
assign v_13625 = v_13623 | v_13624;
assign v_13628 = v_13626 | v_13627;
assign v_13631 = v_13629 | v_13630;
assign v_13634 = v_13632 | v_13633;
assign v_13637 = v_13635 | v_13636;
assign v_13640 = v_13638 | v_13639;
assign v_13643 = v_13641 | v_13642;
assign v_13646 = v_13644 | v_13645;
assign v_13649 = v_13647 | v_13648;
assign v_13652 = v_13650 | v_13651;
assign v_13655 = v_13653 | v_13654;
assign v_13658 = v_13656 | v_13657;
assign v_13661 = v_13659 | v_13660;
assign v_13664 = v_13662 | v_13663;
assign v_13667 = v_13665 | v_13666;
assign v_13670 = v_13668 | v_13669;
assign v_13673 = v_13671 | v_13672;
assign v_13676 = v_13674 | v_13675;
assign v_13679 = v_13677 | v_13678;
assign v_13682 = v_13680 | v_13681;
assign v_13685 = v_13683 | v_13684;
assign v_13688 = v_13686 | v_13687;
assign v_13691 = v_13689 | v_13690;
assign v_13694 = v_13692 | v_13693;
assign v_13697 = v_13695 | v_13696;
assign v_13700 = v_13698 | v_13699;
assign v_13703 = v_13701 | v_13702;
assign v_13706 = v_13704 | v_13705;
assign v_13709 = v_13707 | v_13708;
assign v_13712 = v_13710 | v_13711;
assign v_13715 = v_13713 | v_13714;
assign v_13718 = v_13716 | v_13717;
assign v_13721 = v_13719 | v_13720;
assign v_13724 = v_13722 | v_13723;
assign v_13727 = v_13725 | v_13726;
assign v_13730 = v_13728 | v_13729;
assign v_13733 = v_13731 | v_13732;
assign v_13736 = v_13734 | v_13735;
assign v_13739 = v_13737 | v_13738;
assign v_13742 = v_13740 | v_13741;
assign v_13745 = v_13743 | v_13744;
assign v_13748 = v_13746 | v_13747;
assign v_13751 = v_13749 | v_13750;
assign v_13754 = v_13752 | v_13753;
assign v_13757 = v_13755 | v_13756;
assign v_13760 = v_13758 | v_13759;
assign v_13763 = v_13761 | v_13762;
assign v_13766 = v_13764 | v_13765;
assign v_13769 = v_13767 | v_13768;
assign v_13772 = v_13770 | v_13771;
assign v_13775 = v_13773 | v_13774;
assign v_13778 = v_13776 | v_13777;
assign v_13781 = v_13779 | v_13780;
assign v_13784 = v_13782 | v_13783;
assign v_13787 = v_13785 | v_13786;
assign v_13790 = v_13788 | v_13789;
assign v_13793 = v_13791 | v_13792;
assign v_13796 = v_13794 | v_13795;
assign v_13799 = v_13797 | v_13798;
assign v_13802 = v_13800 | v_13801;
assign v_13805 = v_13803 | v_13804;
assign v_13808 = v_13806 | v_13807;
assign v_13811 = v_13809 | v_13810;
assign v_13814 = v_13812 | v_13813;
assign v_13817 = v_13815 | v_13816;
assign v_13820 = v_13818 | v_13819;
assign v_13823 = v_13821 | v_13822;
assign v_13826 = v_13824 | v_13825;
assign v_13829 = v_13827 | v_13828;
assign v_13832 = v_13830 | v_13831;
assign v_13835 = v_13833 | v_13834;
assign v_13838 = v_13836 | v_13837;
assign v_13841 = v_13839 | v_13840;
assign v_13844 = v_13842 | v_13843;
assign v_13847 = v_13845 | v_13846;
assign v_13850 = v_13848 | v_13849;
assign v_13853 = v_13851 | v_13852;
assign v_13856 = v_13854 | v_13855;
assign v_13859 = v_13857 | v_13858;
assign v_13862 = v_13860 | v_13861;
assign v_13865 = v_13863 | v_13864;
assign v_13868 = v_13866 | v_13867;
assign v_13871 = v_13869 | v_13870;
assign v_13874 = v_13872 | v_13873;
assign v_13877 = v_13875 | v_13876;
assign v_13880 = v_13878 | v_13879;
assign v_13883 = v_13881 | v_13882;
assign v_13886 = v_13884 | v_13885;
assign v_13889 = v_13887 | v_13888;
assign v_13892 = v_13890 | v_13891;
assign v_13895 = v_13893 | v_13894;
assign v_13898 = v_13896 | v_13897;
assign v_13901 = v_13899 | v_13900;
assign v_13904 = v_13902 | v_13903;
assign v_13907 = v_13905 | v_13906;
assign v_13910 = v_13908 | v_13909;
assign v_13913 = v_13911 | v_13912;
assign v_13916 = v_13914 | v_13915;
assign v_13919 = v_13917 | v_13918;
assign v_13922 = v_13920 | v_13921;
assign v_13923 = v_13733 | v_13922;
assign v_13926 = v_13924 | v_13925;
assign v_13929 = v_13927 | v_13928;
assign v_13932 = v_13930 | v_13931;
assign v_13935 = v_13933 | v_13934;
assign v_13938 = v_13936 | v_13937;
assign v_13941 = v_13939 | v_13940;
assign v_13944 = v_13942 | v_13943;
assign v_13947 = v_13945 | v_13946;
assign v_13950 = v_13948 | v_13949;
assign v_13953 = v_13951 | v_13952;
assign v_13956 = v_13954 | v_13955;
assign v_13959 = v_13957 | v_13958;
assign v_13962 = v_13960 | v_13961;
assign v_13965 = v_13963 | v_13964;
assign v_13968 = v_13966 | v_13967;
assign v_13971 = v_13969 | v_13970;
assign v_13974 = v_13972 | v_13973;
assign v_13977 = v_13975 | v_13976;
assign v_13980 = v_13978 | v_13979;
assign v_13983 = v_13981 | v_13982;
assign v_13986 = v_13984 | v_13985;
assign v_13989 = v_13987 | v_13988;
assign v_13992 = v_13990 | v_13991;
assign v_13995 = v_13993 | v_13994;
assign v_13998 = v_13996 | v_13997;
assign v_14001 = v_13999 | v_14000;
assign v_14004 = v_14002 | v_14003;
assign v_14007 = v_14005 | v_14006;
assign v_14010 = v_14008 | v_14009;
assign v_14013 = v_14011 | v_14012;
assign v_14016 = v_14014 | v_14015;
assign v_14019 = v_14017 | v_14018;
assign v_14022 = v_14020 | v_14021;
assign v_14025 = v_14023 | v_14024;
assign v_14028 = v_14026 | v_14027;
assign v_14031 = v_14029 | v_14030;
assign v_14034 = v_14032 | v_14033;
assign v_14037 = v_14035 | v_14036;
assign v_14040 = v_14038 | v_14039;
assign v_14043 = v_14041 | v_14042;
assign v_14046 = v_14044 | v_14045;
assign v_14049 = v_14047 | v_14048;
assign v_14052 = v_14050 | v_14051;
assign v_14055 = v_14053 | v_14054;
assign v_14058 = v_14056 | v_14057;
assign v_14061 = v_14059 | v_14060;
assign v_14064 = v_14062 | v_14063;
assign v_14067 = v_14065 | v_14066;
assign v_14070 = v_14068 | v_14069;
assign v_14073 = v_14071 | v_14072;
assign v_14076 = v_14074 | v_14075;
assign v_14079 = v_14077 | v_14078;
assign v_14082 = v_14080 | v_14081;
assign v_14085 = v_14083 | v_14084;
assign v_14088 = v_14086 | v_14087;
assign v_14091 = v_14089 | v_14090;
assign v_14094 = v_14092 | v_14093;
assign v_14097 = v_14095 | v_14096;
assign v_14100 = v_14098 | v_14099;
assign v_14103 = v_14101 | v_14102;
assign v_14106 = v_14104 | v_14105;
assign v_14109 = v_14107 | v_14108;
assign v_14112 = v_14110 | v_14111;
assign v_14113 = v_13923 | v_14112;
assign v_14116 = v_14114 | v_14115;
assign v_14119 = v_14117 | v_14118;
assign v_14122 = v_14120 | v_14121;
assign v_14125 = v_14123 | v_14124;
assign v_14128 = v_14126 | v_14127;
assign v_14131 = v_14129 | v_14130;
assign v_14134 = v_14132 | v_14133;
assign v_14137 = v_14135 | v_14136;
assign v_14140 = v_14138 | v_14139;
assign v_14143 = v_14141 | v_14142;
assign v_14146 = v_14144 | v_14145;
assign v_14149 = v_14147 | v_14148;
assign v_14152 = v_14150 | v_14151;
assign v_14155 = v_14153 | v_14154;
assign v_14158 = v_14156 | v_14157;
assign v_14161 = v_14159 | v_14160;
assign v_14164 = v_14162 | v_14163;
assign v_14167 = v_14165 | v_14166;
assign v_14170 = v_14168 | v_14169;
assign v_14173 = v_14171 | v_14172;
assign v_14176 = v_14174 | v_14175;
assign v_14179 = v_14177 | v_14178;
assign v_14182 = v_14180 | v_14181;
assign v_14185 = v_14183 | v_14184;
assign v_14188 = v_14186 | v_14187;
assign v_14191 = v_14189 | v_14190;
assign v_14194 = v_14192 | v_14193;
assign v_14197 = v_14195 | v_14196;
assign v_14200 = v_14198 | v_14199;
assign v_14203 = v_14201 | v_14202;
assign v_14206 = v_14204 | v_14205;
assign v_14209 = v_14207 | v_14208;
assign v_14212 = v_14210 | v_14211;
assign v_14215 = v_14213 | v_14214;
assign v_14218 = v_14216 | v_14217;
assign v_14221 = v_14219 | v_14220;
assign v_14224 = v_14222 | v_14223;
assign v_14227 = v_14225 | v_14226;
assign v_14230 = v_14228 | v_14229;
assign v_14233 = v_14231 | v_14232;
assign v_14236 = v_14234 | v_14235;
assign v_14239 = v_14237 | v_14238;
assign v_14242 = v_14240 | v_14241;
assign v_14245 = v_14243 | v_14244;
assign v_14248 = v_14246 | v_14247;
assign v_14251 = v_14249 | v_14250;
assign v_14254 = v_14252 | v_14253;
assign v_14257 = v_14255 | v_14256;
assign v_14260 = v_14258 | v_14259;
assign v_14263 = v_14261 | v_14262;
assign v_14266 = v_14264 | v_14265;
assign v_14269 = v_14267 | v_14268;
assign v_14272 = v_14270 | v_14271;
assign v_14275 = v_14273 | v_14274;
assign v_14278 = v_14276 | v_14277;
assign v_14281 = v_14279 | v_14280;
assign v_14284 = v_14282 | v_14283;
assign v_14287 = v_14285 | v_14286;
assign v_14290 = v_14288 | v_14289;
assign v_14293 = v_14291 | v_14292;
assign v_14296 = v_14294 | v_14295;
assign v_14299 = v_14297 | v_14298;
assign v_14302 = v_14300 | v_14301;
assign v_14303 = v_14113 | v_14302;
assign v_14306 = v_14304 | v_14305;
assign v_14309 = v_14307 | v_14308;
assign v_14312 = v_14310 | v_14311;
assign v_14315 = v_14313 | v_14314;
assign v_14318 = v_14316 | v_14317;
assign v_14321 = v_14319 | v_14320;
assign v_14324 = v_14322 | v_14323;
assign v_14327 = v_14325 | v_14326;
assign v_14330 = v_14328 | v_14329;
assign v_14333 = v_14331 | v_14332;
assign v_14336 = v_14334 | v_14335;
assign v_14339 = v_14337 | v_14338;
assign v_14342 = v_14340 | v_14341;
assign v_14345 = v_14343 | v_14344;
assign v_14348 = v_14346 | v_14347;
assign v_14351 = v_14349 | v_14350;
assign v_14354 = v_14352 | v_14353;
assign v_14357 = v_14355 | v_14356;
assign v_14360 = v_14358 | v_14359;
assign v_14363 = v_14361 | v_14362;
assign v_14366 = v_14364 | v_14365;
assign v_14369 = v_14367 | v_14368;
assign v_14372 = v_14370 | v_14371;
assign v_14375 = v_14373 | v_14374;
assign v_14378 = v_14376 | v_14377;
assign v_14381 = v_14379 | v_14380;
assign v_14384 = v_14382 | v_14383;
assign v_14387 = v_14385 | v_14386;
assign v_14390 = v_14388 | v_14389;
assign v_14393 = v_14391 | v_14392;
assign v_14396 = v_14394 | v_14395;
assign v_14399 = v_14397 | v_14398;
assign v_14402 = v_14400 | v_14401;
assign v_14405 = v_14403 | v_14404;
assign v_14408 = v_14406 | v_14407;
assign v_14411 = v_14409 | v_14410;
assign v_14414 = v_14412 | v_14413;
assign v_14417 = v_14415 | v_14416;
assign v_14420 = v_14418 | v_14419;
assign v_14423 = v_14421 | v_14422;
assign v_14426 = v_14424 | v_14425;
assign v_14429 = v_14427 | v_14428;
assign v_14432 = v_14430 | v_14431;
assign v_14435 = v_14433 | v_14434;
assign v_14438 = v_14436 | v_14437;
assign v_14441 = v_14439 | v_14440;
assign v_14444 = v_14442 | v_14443;
assign v_14447 = v_14445 | v_14446;
assign v_14450 = v_14448 | v_14449;
assign v_14453 = v_14451 | v_14452;
assign v_14456 = v_14454 | v_14455;
assign v_14459 = v_14457 | v_14458;
assign v_14462 = v_14460 | v_14461;
assign v_14465 = v_14463 | v_14464;
assign v_14468 = v_14466 | v_14467;
assign v_14471 = v_14469 | v_14470;
assign v_14474 = v_14472 | v_14473;
assign v_14477 = v_14475 | v_14476;
assign v_14480 = v_14478 | v_14479;
assign v_14483 = v_14481 | v_14482;
assign v_14486 = v_14484 | v_14485;
assign v_14489 = v_14487 | v_14488;
assign v_14492 = v_14490 | v_14491;
assign v_14493 = v_14303 | v_14492;
assign v_14496 = v_14494 | v_14495;
assign v_14499 = v_14497 | v_14498;
assign v_14502 = v_14500 | v_14501;
assign v_14505 = v_14503 | v_14504;
assign v_14508 = v_14506 | v_14507;
assign v_14511 = v_14509 | v_14510;
assign v_14514 = v_14512 | v_14513;
assign v_14517 = v_14515 | v_14516;
assign v_14520 = v_14518 | v_14519;
assign v_14523 = v_14521 | v_14522;
assign v_14526 = v_14524 | v_14525;
assign v_14529 = v_14527 | v_14528;
assign v_14532 = v_14530 | v_14531;
assign v_14535 = v_14533 | v_14534;
assign v_14538 = v_14536 | v_14537;
assign v_14541 = v_14539 | v_14540;
assign v_14544 = v_14542 | v_14543;
assign v_14547 = v_14545 | v_14546;
assign v_14550 = v_14548 | v_14549;
assign v_14553 = v_14551 | v_14552;
assign v_14556 = v_14554 | v_14555;
assign v_14559 = v_14557 | v_14558;
assign v_14562 = v_14560 | v_14561;
assign v_14565 = v_14563 | v_14564;
assign v_14568 = v_14566 | v_14567;
assign v_14571 = v_14569 | v_14570;
assign v_14574 = v_14572 | v_14573;
assign v_14577 = v_14575 | v_14576;
assign v_14580 = v_14578 | v_14579;
assign v_14583 = v_14581 | v_14582;
assign v_14586 = v_14584 | v_14585;
assign v_14589 = v_14587 | v_14588;
assign v_14592 = v_14590 | v_14591;
assign v_14595 = v_14593 | v_14594;
assign v_14598 = v_14596 | v_14597;
assign v_14601 = v_14599 | v_14600;
assign v_14604 = v_14602 | v_14603;
assign v_14607 = v_14605 | v_14606;
assign v_14610 = v_14608 | v_14609;
assign v_14613 = v_14611 | v_14612;
assign v_14616 = v_14614 | v_14615;
assign v_14619 = v_14617 | v_14618;
assign v_14622 = v_14620 | v_14621;
assign v_14625 = v_14623 | v_14624;
assign v_14628 = v_14626 | v_14627;
assign v_14631 = v_14629 | v_14630;
assign v_14634 = v_14632 | v_14633;
assign v_14637 = v_14635 | v_14636;
assign v_14640 = v_14638 | v_14639;
assign v_14643 = v_14641 | v_14642;
assign v_14646 = v_14644 | v_14645;
assign v_14649 = v_14647 | v_14648;
assign v_14652 = v_14650 | v_14651;
assign v_14655 = v_14653 | v_14654;
assign v_14658 = v_14656 | v_14657;
assign v_14661 = v_14659 | v_14660;
assign v_14664 = v_14662 | v_14663;
assign v_14667 = v_14665 | v_14666;
assign v_14670 = v_14668 | v_14669;
assign v_14673 = v_14671 | v_14672;
assign v_14676 = v_14674 | v_14675;
assign v_14679 = v_14677 | v_14678;
assign v_14682 = v_14680 | v_14681;
assign v_14683 = v_14493 | v_14682;
assign v_14686 = v_14684 | v_14685;
assign v_14689 = v_14687 | v_14688;
assign v_14692 = v_14690 | v_14691;
assign v_14695 = v_14693 | v_14694;
assign v_14698 = v_14696 | v_14697;
assign v_14701 = v_14699 | v_14700;
assign v_14704 = v_14702 | v_14703;
assign v_14707 = v_14705 | v_14706;
assign v_14710 = v_14708 | v_14709;
assign v_14713 = v_14711 | v_14712;
assign v_14716 = v_14714 | v_14715;
assign v_14719 = v_14717 | v_14718;
assign v_14722 = v_14720 | v_14721;
assign v_14725 = v_14723 | v_14724;
assign v_14728 = v_14726 | v_14727;
assign v_14731 = v_14729 | v_14730;
assign v_14734 = v_14732 | v_14733;
assign v_14737 = v_14735 | v_14736;
assign v_14740 = v_14738 | v_14739;
assign v_14743 = v_14741 | v_14742;
assign v_14746 = v_14744 | v_14745;
assign v_14749 = v_14747 | v_14748;
assign v_14752 = v_14750 | v_14751;
assign v_14755 = v_14753 | v_14754;
assign v_14758 = v_14756 | v_14757;
assign v_14761 = v_14759 | v_14760;
assign v_14764 = v_14762 | v_14763;
assign v_14767 = v_14765 | v_14766;
assign v_14770 = v_14768 | v_14769;
assign v_14773 = v_14771 | v_14772;
assign v_14776 = v_14774 | v_14775;
assign v_14779 = v_14777 | v_14778;
assign v_14782 = v_14780 | v_14781;
assign v_14785 = v_14783 | v_14784;
assign v_14788 = v_14786 | v_14787;
assign v_14791 = v_14789 | v_14790;
assign v_14794 = v_14792 | v_14793;
assign v_14797 = v_14795 | v_14796;
assign v_14800 = v_14798 | v_14799;
assign v_14803 = v_14801 | v_14802;
assign v_14806 = v_14804 | v_14805;
assign v_14809 = v_14807 | v_14808;
assign v_14812 = v_14810 | v_14811;
assign v_14815 = v_14813 | v_14814;
assign v_14818 = v_14816 | v_14817;
assign v_14821 = v_14819 | v_14820;
assign v_14824 = v_14822 | v_14823;
assign v_14827 = v_14825 | v_14826;
assign v_14830 = v_14828 | v_14829;
assign v_14833 = v_14831 | v_14832;
assign v_14836 = v_14834 | v_14835;
assign v_14839 = v_14837 | v_14838;
assign v_14842 = v_14840 | v_14841;
assign v_14845 = v_14843 | v_14844;
assign v_14848 = v_14846 | v_14847;
assign v_14851 = v_14849 | v_14850;
assign v_14854 = v_14852 | v_14853;
assign v_14857 = v_14855 | v_14856;
assign v_14860 = v_14858 | v_14859;
assign v_14863 = v_14861 | v_14862;
assign v_14866 = v_14864 | v_14865;
assign v_14869 = v_14867 | v_14868;
assign v_14872 = v_14870 | v_14871;
assign v_14873 = v_14683 | v_14872;
assign v_14876 = v_14874 | v_14875;
assign v_14879 = v_14877 | v_14878;
assign v_14882 = v_14880 | v_14881;
assign v_14885 = v_14883 | v_14884;
assign v_14888 = v_14886 | v_14887;
assign v_14891 = v_14889 | v_14890;
assign v_14894 = v_14892 | v_14893;
assign v_14897 = v_14895 | v_14896;
assign v_14900 = v_14898 | v_14899;
assign v_14903 = v_14901 | v_14902;
assign v_14906 = v_14904 | v_14905;
assign v_14909 = v_14907 | v_14908;
assign v_14912 = v_14910 | v_14911;
assign v_14915 = v_14913 | v_14914;
assign v_14918 = v_14916 | v_14917;
assign v_14921 = v_14919 | v_14920;
assign v_14924 = v_14922 | v_14923;
assign v_14927 = v_14925 | v_14926;
assign v_14930 = v_14928 | v_14929;
assign v_14933 = v_14931 | v_14932;
assign v_14936 = v_14934 | v_14935;
assign v_14939 = v_14937 | v_14938;
assign v_14942 = v_14940 | v_14941;
assign v_14945 = v_14943 | v_14944;
assign v_14948 = v_14946 | v_14947;
assign v_14951 = v_14949 | v_14950;
assign v_14954 = v_14952 | v_14953;
assign v_14957 = v_14955 | v_14956;
assign v_14960 = v_14958 | v_14959;
assign v_14963 = v_14961 | v_14962;
assign v_14966 = v_14964 | v_14965;
assign v_14969 = v_14967 | v_14968;
assign v_14972 = v_14970 | v_14971;
assign v_14975 = v_14973 | v_14974;
assign v_14978 = v_14976 | v_14977;
assign v_14981 = v_14979 | v_14980;
assign v_14984 = v_14982 | v_14983;
assign v_14987 = v_14985 | v_14986;
assign v_14990 = v_14988 | v_14989;
assign v_14993 = v_14991 | v_14992;
assign v_14996 = v_14994 | v_14995;
assign v_14999 = v_14997 | v_14998;
assign v_15002 = v_15000 | v_15001;
assign v_15005 = v_15003 | v_15004;
assign v_15008 = v_15006 | v_15007;
assign v_15011 = v_15009 | v_15010;
assign v_15014 = v_15012 | v_15013;
assign v_15017 = v_15015 | v_15016;
assign v_15020 = v_15018 | v_15019;
assign v_15023 = v_15021 | v_15022;
assign v_15026 = v_15024 | v_15025;
assign v_15029 = v_15027 | v_15028;
assign v_15032 = v_15030 | v_15031;
assign v_15035 = v_15033 | v_15034;
assign v_15038 = v_15036 | v_15037;
assign v_15041 = v_15039 | v_15040;
assign v_15044 = v_15042 | v_15043;
assign v_15047 = v_15045 | v_15046;
assign v_15050 = v_15048 | v_15049;
assign v_15053 = v_15051 | v_15052;
assign v_15056 = v_15054 | v_15055;
assign v_15059 = v_15057 | v_15058;
assign v_15062 = v_15060 | v_15061;
assign v_15063 = v_14873 | v_15062;
assign v_15066 = v_15064 | v_15065;
assign v_15069 = v_15067 | v_15068;
assign v_15072 = v_15070 | v_15071;
assign v_15075 = v_15073 | v_15074;
assign v_15078 = v_15076 | v_15077;
assign v_15081 = v_15079 | v_15080;
assign v_15084 = v_15082 | v_15083;
assign v_15087 = v_15085 | v_15086;
assign v_15090 = v_15088 | v_15089;
assign v_15093 = v_15091 | v_15092;
assign v_15096 = v_15094 | v_15095;
assign v_15099 = v_15097 | v_15098;
assign v_15102 = v_15100 | v_15101;
assign v_15105 = v_15103 | v_15104;
assign v_15108 = v_15106 | v_15107;
assign v_15111 = v_15109 | v_15110;
assign v_15114 = v_15112 | v_15113;
assign v_15117 = v_15115 | v_15116;
assign v_15120 = v_15118 | v_15119;
assign v_15123 = v_15121 | v_15122;
assign v_15126 = v_15124 | v_15125;
assign v_15129 = v_15127 | v_15128;
assign v_15132 = v_15130 | v_15131;
assign v_15135 = v_15133 | v_15134;
assign v_15138 = v_15136 | v_15137;
assign v_15141 = v_15139 | v_15140;
assign v_15144 = v_15142 | v_15143;
assign v_15147 = v_15145 | v_15146;
assign v_15150 = v_15148 | v_15149;
assign v_15153 = v_15151 | v_15152;
assign v_15156 = v_15154 | v_15155;
assign v_15159 = v_15157 | v_15158;
assign v_15162 = v_15160 | v_15161;
assign v_15165 = v_15163 | v_15164;
assign v_15168 = v_15166 | v_15167;
assign v_15171 = v_15169 | v_15170;
assign v_15174 = v_15172 | v_15173;
assign v_15177 = v_15175 | v_15176;
assign v_15180 = v_15178 | v_15179;
assign v_15183 = v_15181 | v_15182;
assign v_15186 = v_15184 | v_15185;
assign v_15189 = v_15187 | v_15188;
assign v_15192 = v_15190 | v_15191;
assign v_15195 = v_15193 | v_15194;
assign v_15198 = v_15196 | v_15197;
assign v_15201 = v_15199 | v_15200;
assign v_15204 = v_15202 | v_15203;
assign v_15207 = v_15205 | v_15206;
assign v_15210 = v_15208 | v_15209;
assign v_15213 = v_15211 | v_15212;
assign v_15216 = v_15214 | v_15215;
assign v_15219 = v_15217 | v_15218;
assign v_15222 = v_15220 | v_15221;
assign v_15225 = v_15223 | v_15224;
assign v_15228 = v_15226 | v_15227;
assign v_15231 = v_15229 | v_15230;
assign v_15234 = v_15232 | v_15233;
assign v_15237 = v_15235 | v_15236;
assign v_15240 = v_15238 | v_15239;
assign v_15243 = v_15241 | v_15242;
assign v_15246 = v_15244 | v_15245;
assign v_15249 = v_15247 | v_15248;
assign v_15252 = v_15250 | v_15251;
assign v_15255 = v_15253 | v_15254;
assign v_15258 = v_15256 | v_15257;
assign v_15261 = v_15259 | v_15260;
assign v_15264 = v_15262 | v_15263;
assign v_15267 = v_15265 | v_15266;
assign v_15270 = v_15268 | v_15269;
assign v_15273 = v_15271 | v_15272;
assign v_15276 = v_15274 | v_15275;
assign v_15279 = v_15277 | v_15278;
assign v_15282 = v_15280 | v_15281;
assign v_15285 = v_15283 | v_15284;
assign v_15288 = v_15286 | v_15287;
assign v_15291 = v_15289 | v_15290;
assign v_15294 = v_15292 | v_15293;
assign v_15297 = v_15295 | v_15296;
assign v_15300 = v_15298 | v_15299;
assign v_15303 = v_15301 | v_15302;
assign v_15306 = v_15304 | v_15305;
assign v_15309 = v_15307 | v_15308;
assign v_15312 = v_15310 | v_15311;
assign v_15315 = v_15313 | v_15314;
assign v_15318 = v_15316 | v_15317;
assign v_15321 = v_15319 | v_15320;
assign v_15324 = v_15322 | v_15323;
assign v_15327 = v_15325 | v_15326;
assign v_15330 = v_15328 | v_15329;
assign v_15333 = v_15331 | v_15332;
assign v_15336 = v_15334 | v_15335;
assign v_15339 = v_15337 | v_15338;
assign v_15342 = v_15340 | v_15341;
assign v_15345 = v_15343 | v_15344;
assign v_15348 = v_15346 | v_15347;
assign v_15351 = v_15349 | v_15350;
assign v_15354 = v_15352 | v_15353;
assign v_15357 = v_15355 | v_15356;
assign v_15360 = v_15358 | v_15359;
assign v_15363 = v_15361 | v_15362;
assign v_15366 = v_15364 | v_15365;
assign v_15369 = v_15367 | v_15368;
assign v_15372 = v_15370 | v_15371;
assign v_15375 = v_15373 | v_15374;
assign v_15378 = v_15376 | v_15377;
assign v_15381 = v_15379 | v_15380;
assign v_15384 = v_15382 | v_15383;
assign v_15387 = v_15385 | v_15386;
assign v_15390 = v_15388 | v_15389;
assign v_15393 = v_15391 | v_15392;
assign v_15396 = v_15394 | v_15395;
assign v_15399 = v_15397 | v_15398;
assign v_15402 = v_15400 | v_15401;
assign v_15405 = v_15403 | v_15404;
assign v_15408 = v_15406 | v_15407;
assign v_15411 = v_15409 | v_15410;
assign v_15414 = v_15412 | v_15413;
assign v_15417 = v_15415 | v_15416;
assign v_15420 = v_15418 | v_15419;
assign v_15423 = v_15421 | v_15422;
assign v_15426 = v_15424 | v_15425;
assign v_15429 = v_15427 | v_15428;
assign v_15432 = v_15430 | v_15431;
assign v_15435 = v_15433 | v_15434;
assign v_15438 = v_15436 | v_15437;
assign v_15441 = v_15439 | v_15440;
assign v_15442 = v_15252 | v_15441;
assign v_15445 = v_15443 | v_15444;
assign v_15448 = v_15446 | v_15447;
assign v_15451 = v_15449 | v_15450;
assign v_15454 = v_15452 | v_15453;
assign v_15457 = v_15455 | v_15456;
assign v_15460 = v_15458 | v_15459;
assign v_15463 = v_15461 | v_15462;
assign v_15466 = v_15464 | v_15465;
assign v_15469 = v_15467 | v_15468;
assign v_15472 = v_15470 | v_15471;
assign v_15475 = v_15473 | v_15474;
assign v_15478 = v_15476 | v_15477;
assign v_15481 = v_15479 | v_15480;
assign v_15484 = v_15482 | v_15483;
assign v_15487 = v_15485 | v_15486;
assign v_15490 = v_15488 | v_15489;
assign v_15493 = v_15491 | v_15492;
assign v_15496 = v_15494 | v_15495;
assign v_15499 = v_15497 | v_15498;
assign v_15502 = v_15500 | v_15501;
assign v_15505 = v_15503 | v_15504;
assign v_15508 = v_15506 | v_15507;
assign v_15511 = v_15509 | v_15510;
assign v_15514 = v_15512 | v_15513;
assign v_15517 = v_15515 | v_15516;
assign v_15520 = v_15518 | v_15519;
assign v_15523 = v_15521 | v_15522;
assign v_15526 = v_15524 | v_15525;
assign v_15529 = v_15527 | v_15528;
assign v_15532 = v_15530 | v_15531;
assign v_15535 = v_15533 | v_15534;
assign v_15538 = v_15536 | v_15537;
assign v_15541 = v_15539 | v_15540;
assign v_15544 = v_15542 | v_15543;
assign v_15547 = v_15545 | v_15546;
assign v_15550 = v_15548 | v_15549;
assign v_15553 = v_15551 | v_15552;
assign v_15556 = v_15554 | v_15555;
assign v_15559 = v_15557 | v_15558;
assign v_15562 = v_15560 | v_15561;
assign v_15565 = v_15563 | v_15564;
assign v_15568 = v_15566 | v_15567;
assign v_15571 = v_15569 | v_15570;
assign v_15574 = v_15572 | v_15573;
assign v_15577 = v_15575 | v_15576;
assign v_15580 = v_15578 | v_15579;
assign v_15583 = v_15581 | v_15582;
assign v_15586 = v_15584 | v_15585;
assign v_15589 = v_15587 | v_15588;
assign v_15592 = v_15590 | v_15591;
assign v_15595 = v_15593 | v_15594;
assign v_15598 = v_15596 | v_15597;
assign v_15601 = v_15599 | v_15600;
assign v_15604 = v_15602 | v_15603;
assign v_15607 = v_15605 | v_15606;
assign v_15610 = v_15608 | v_15609;
assign v_15613 = v_15611 | v_15612;
assign v_15616 = v_15614 | v_15615;
assign v_15619 = v_15617 | v_15618;
assign v_15622 = v_15620 | v_15621;
assign v_15625 = v_15623 | v_15624;
assign v_15628 = v_15626 | v_15627;
assign v_15631 = v_15629 | v_15630;
assign v_15632 = v_15442 | v_15631;
assign v_15635 = v_15633 | v_15634;
assign v_15638 = v_15636 | v_15637;
assign v_15641 = v_15639 | v_15640;
assign v_15644 = v_15642 | v_15643;
assign v_15647 = v_15645 | v_15646;
assign v_15650 = v_15648 | v_15649;
assign v_15653 = v_15651 | v_15652;
assign v_15656 = v_15654 | v_15655;
assign v_15659 = v_15657 | v_15658;
assign v_15662 = v_15660 | v_15661;
assign v_15665 = v_15663 | v_15664;
assign v_15668 = v_15666 | v_15667;
assign v_15671 = v_15669 | v_15670;
assign v_15674 = v_15672 | v_15673;
assign v_15677 = v_15675 | v_15676;
assign v_15680 = v_15678 | v_15679;
assign v_15683 = v_15681 | v_15682;
assign v_15686 = v_15684 | v_15685;
assign v_15689 = v_15687 | v_15688;
assign v_15692 = v_15690 | v_15691;
assign v_15695 = v_15693 | v_15694;
assign v_15698 = v_15696 | v_15697;
assign v_15701 = v_15699 | v_15700;
assign v_15704 = v_15702 | v_15703;
assign v_15707 = v_15705 | v_15706;
assign v_15710 = v_15708 | v_15709;
assign v_15713 = v_15711 | v_15712;
assign v_15716 = v_15714 | v_15715;
assign v_15719 = v_15717 | v_15718;
assign v_15722 = v_15720 | v_15721;
assign v_15725 = v_15723 | v_15724;
assign v_15728 = v_15726 | v_15727;
assign v_15731 = v_15729 | v_15730;
assign v_15734 = v_15732 | v_15733;
assign v_15737 = v_15735 | v_15736;
assign v_15740 = v_15738 | v_15739;
assign v_15743 = v_15741 | v_15742;
assign v_15746 = v_15744 | v_15745;
assign v_15749 = v_15747 | v_15748;
assign v_15752 = v_15750 | v_15751;
assign v_15755 = v_15753 | v_15754;
assign v_15758 = v_15756 | v_15757;
assign v_15761 = v_15759 | v_15760;
assign v_15764 = v_15762 | v_15763;
assign v_15767 = v_15765 | v_15766;
assign v_15770 = v_15768 | v_15769;
assign v_15773 = v_15771 | v_15772;
assign v_15776 = v_15774 | v_15775;
assign v_15779 = v_15777 | v_15778;
assign v_15782 = v_15780 | v_15781;
assign v_15785 = v_15783 | v_15784;
assign v_15788 = v_15786 | v_15787;
assign v_15791 = v_15789 | v_15790;
assign v_15794 = v_15792 | v_15793;
assign v_15797 = v_15795 | v_15796;
assign v_15800 = v_15798 | v_15799;
assign v_15803 = v_15801 | v_15802;
assign v_15806 = v_15804 | v_15805;
assign v_15809 = v_15807 | v_15808;
assign v_15812 = v_15810 | v_15811;
assign v_15815 = v_15813 | v_15814;
assign v_15818 = v_15816 | v_15817;
assign v_15821 = v_15819 | v_15820;
assign v_15822 = v_15632 | v_15821;
assign v_15825 = v_15823 | v_15824;
assign v_15828 = v_15826 | v_15827;
assign v_15831 = v_15829 | v_15830;
assign v_15834 = v_15832 | v_15833;
assign v_15837 = v_15835 | v_15836;
assign v_15840 = v_15838 | v_15839;
assign v_15843 = v_15841 | v_15842;
assign v_15846 = v_15844 | v_15845;
assign v_15849 = v_15847 | v_15848;
assign v_15852 = v_15850 | v_15851;
assign v_15855 = v_15853 | v_15854;
assign v_15858 = v_15856 | v_15857;
assign v_15861 = v_15859 | v_15860;
assign v_15864 = v_15862 | v_15863;
assign v_15867 = v_15865 | v_15866;
assign v_15870 = v_15868 | v_15869;
assign v_15873 = v_15871 | v_15872;
assign v_15876 = v_15874 | v_15875;
assign v_15879 = v_15877 | v_15878;
assign v_15882 = v_15880 | v_15881;
assign v_15885 = v_15883 | v_15884;
assign v_15888 = v_15886 | v_15887;
assign v_15891 = v_15889 | v_15890;
assign v_15894 = v_15892 | v_15893;
assign v_15897 = v_15895 | v_15896;
assign v_15900 = v_15898 | v_15899;
assign v_15903 = v_15901 | v_15902;
assign v_15906 = v_15904 | v_15905;
assign v_15909 = v_15907 | v_15908;
assign v_15912 = v_15910 | v_15911;
assign v_15915 = v_15913 | v_15914;
assign v_15918 = v_15916 | v_15917;
assign v_15921 = v_15919 | v_15920;
assign v_15924 = v_15922 | v_15923;
assign v_15927 = v_15925 | v_15926;
assign v_15930 = v_15928 | v_15929;
assign v_15933 = v_15931 | v_15932;
assign v_15936 = v_15934 | v_15935;
assign v_15939 = v_15937 | v_15938;
assign v_15942 = v_15940 | v_15941;
assign v_15945 = v_15943 | v_15944;
assign v_15948 = v_15946 | v_15947;
assign v_15951 = v_15949 | v_15950;
assign v_15954 = v_15952 | v_15953;
assign v_15957 = v_15955 | v_15956;
assign v_15960 = v_15958 | v_15959;
assign v_15963 = v_15961 | v_15962;
assign v_15966 = v_15964 | v_15965;
assign v_15969 = v_15967 | v_15968;
assign v_15972 = v_15970 | v_15971;
assign v_15975 = v_15973 | v_15974;
assign v_15978 = v_15976 | v_15977;
assign v_15981 = v_15979 | v_15980;
assign v_15984 = v_15982 | v_15983;
assign v_15987 = v_15985 | v_15986;
assign v_15990 = v_15988 | v_15989;
assign v_15993 = v_15991 | v_15992;
assign v_15996 = v_15994 | v_15995;
assign v_15999 = v_15997 | v_15998;
assign v_16002 = v_16000 | v_16001;
assign v_16005 = v_16003 | v_16004;
assign v_16008 = v_16006 | v_16007;
assign v_16011 = v_16009 | v_16010;
assign v_16012 = v_15822 | v_16011;
assign v_16015 = v_16013 | v_16014;
assign v_16018 = v_16016 | v_16017;
assign v_16021 = v_16019 | v_16020;
assign v_16024 = v_16022 | v_16023;
assign v_16027 = v_16025 | v_16026;
assign v_16030 = v_16028 | v_16029;
assign v_16033 = v_16031 | v_16032;
assign v_16036 = v_16034 | v_16035;
assign v_16039 = v_16037 | v_16038;
assign v_16042 = v_16040 | v_16041;
assign v_16045 = v_16043 | v_16044;
assign v_16048 = v_16046 | v_16047;
assign v_16051 = v_16049 | v_16050;
assign v_16054 = v_16052 | v_16053;
assign v_16057 = v_16055 | v_16056;
assign v_16060 = v_16058 | v_16059;
assign v_16063 = v_16061 | v_16062;
assign v_16066 = v_16064 | v_16065;
assign v_16069 = v_16067 | v_16068;
assign v_16072 = v_16070 | v_16071;
assign v_16075 = v_16073 | v_16074;
assign v_16078 = v_16076 | v_16077;
assign v_16081 = v_16079 | v_16080;
assign v_16084 = v_16082 | v_16083;
assign v_16087 = v_16085 | v_16086;
assign v_16090 = v_16088 | v_16089;
assign v_16093 = v_16091 | v_16092;
assign v_16096 = v_16094 | v_16095;
assign v_16099 = v_16097 | v_16098;
assign v_16102 = v_16100 | v_16101;
assign v_16105 = v_16103 | v_16104;
assign v_16108 = v_16106 | v_16107;
assign v_16111 = v_16109 | v_16110;
assign v_16114 = v_16112 | v_16113;
assign v_16117 = v_16115 | v_16116;
assign v_16120 = v_16118 | v_16119;
assign v_16123 = v_16121 | v_16122;
assign v_16126 = v_16124 | v_16125;
assign v_16129 = v_16127 | v_16128;
assign v_16132 = v_16130 | v_16131;
assign v_16135 = v_16133 | v_16134;
assign v_16138 = v_16136 | v_16137;
assign v_16141 = v_16139 | v_16140;
assign v_16144 = v_16142 | v_16143;
assign v_16147 = v_16145 | v_16146;
assign v_16150 = v_16148 | v_16149;
assign v_16153 = v_16151 | v_16152;
assign v_16156 = v_16154 | v_16155;
assign v_16159 = v_16157 | v_16158;
assign v_16162 = v_16160 | v_16161;
assign v_16165 = v_16163 | v_16164;
assign v_16168 = v_16166 | v_16167;
assign v_16171 = v_16169 | v_16170;
assign v_16174 = v_16172 | v_16173;
assign v_16177 = v_16175 | v_16176;
assign v_16180 = v_16178 | v_16179;
assign v_16183 = v_16181 | v_16182;
assign v_16186 = v_16184 | v_16185;
assign v_16189 = v_16187 | v_16188;
assign v_16192 = v_16190 | v_16191;
assign v_16195 = v_16193 | v_16194;
assign v_16198 = v_16196 | v_16197;
assign v_16201 = v_16199 | v_16200;
assign v_16202 = v_16012 | v_16201;
assign v_16203 = v_9639 | ~v_9844;
assign v_16204 = v_9611 | ~v_9712;
assign v_16206 = v_9483 | v_16205;
assign v_16207 = v_9468 | ~v_9554;
assign v_16209 = v_9347 | v_16208;
assign v_16210 = v_9320 | ~v_9422;
assign v_16212 = v_9195 | v_16211;
assign v_16213 = v_9180 | ~v_9266;
assign v_16215 = v_9061 | v_16214;
assign v_16216 = v_9037 | ~v_9134;
assign v_16218 = v_8913 | v_16217;
assign v_16219 = v_8898 | ~v_8984;
assign v_16221 = v_8775 | v_16220;
assign v_16222 = v_8744 | ~v_8852;
assign v_16224 = v_8617 | v_16223;
assign v_16225 = v_8602 | ~v_8688;
assign v_16227 = v_8483 | v_16226;
assign v_16228 = v_8458 | ~v_8556;
assign v_16230 = v_8333 | v_16229;
assign v_16231 = v_8318 | ~v_8404;
assign v_16233 = v_8197 | v_16232;
assign v_16234 = v_8170 | ~v_8272;
assign v_16236 = v_8045 | v_16235;
assign v_16237 = v_8030 | ~v_8116;
assign v_16239 = v_7911 | v_16238;
assign v_16240 = v_7887 | ~v_7984;
assign v_16242 = v_7763 | v_16241;
assign v_16243 = v_7748 | ~v_7834;
assign v_16245 = v_7623 | v_16244;
assign v_16246 = v_7588 | ~v_7702;
assign v_16248 = v_7459 | v_16247;
assign v_16249 = v_7444 | ~v_7530;
assign v_16251 = v_7325 | v_16250;
assign v_16252 = v_7299 | ~v_7398;
assign v_16254 = v_7173 | v_16253;
assign v_16255 = v_7158 | ~v_7244;
assign v_16257 = v_7037 | v_16256;
assign v_16258 = v_7010 | ~v_7112;
assign v_16260 = v_6885 | v_16259;
assign v_16261 = v_6870 | ~v_6956;
assign v_16263 = v_6751 | v_16262;
assign v_16264 = v_6727 | v_6824;
assign v_16266 = v_6603 | v_16265;
assign v_16267 = v_6588 | ~v_6674;
assign v_16269 = v_6465 | v_16268;
assign v_16270 = v_6434 | ~v_6542;
assign v_16272 = v_6307 | v_16271;
assign v_16273 = v_6292 | ~v_6378;
assign v_16275 = v_6173 | v_16274;
assign v_16276 = v_6148 | ~v_6246;
assign v_16278 = v_6023 | v_16277;
assign v_16279 = v_6008 | v_6094;
assign v_16281 = v_5887 | v_16280;
assign v_16282 = v_5860 | ~v_5962;
assign v_16284 = v_5735 | v_16283;
assign v_16285 = v_5720 | v_5806;
assign v_16287 = v_5601 | v_16286;
assign v_16288 = v_5577 | ~v_5674;
assign v_16290 = v_5453 | v_16289;
assign v_16291 = v_5438 | ~v_5524;
assign v_16293 = v_5311 | v_16292;
assign v_16294 = v_5272 | ~v_5392;
assign v_16296 = v_5141 | v_16295;
assign v_16297 = v_5126 | ~v_5212;
assign v_16299 = v_5007 | v_16298;
assign v_16300 = v_4980 | ~v_5080;
assign v_16302 = v_4853 | v_16301;
assign v_16303 = v_4838 | ~v_4924;
assign v_16305 = v_4717 | v_16304;
assign v_16306 = v_4690 | ~v_4792;
assign v_16308 = v_4565 | v_16307;
assign v_16309 = v_4550 | ~v_4636;
assign v_16311 = v_4431 | v_16310;
assign v_16312 = v_4407 | ~v_4504;
assign v_16314 = v_4283 | v_16313;
assign v_16315 = v_4268 | ~v_4354;
assign v_16317 = v_4145 | v_16316;
assign v_16318 = v_4114 | ~v_4222;
assign v_16320 = v_3987 | v_16319;
assign v_16321 = v_3972 | ~v_4058;
assign v_16323 = v_3853 | v_16322;
assign v_16324 = v_3828 | ~v_3926;
assign v_16326 = v_3703 | v_16325;
assign v_16327 = v_3688 | ~v_3774;
assign v_16329 = v_3567 | v_16328;
assign v_16330 = v_3540 | ~v_3642;
assign v_16332 = v_3415 | v_16331;
assign v_16333 = v_3400 | ~v_3486;
assign v_16335 = v_3281 | v_16334;
assign v_16336 = v_3257 | ~v_3354;
assign v_16338 = v_3133 | v_16337;
assign v_16339 = v_3118 | v_3204;
assign v_16341 = v_2993 | v_16340;
assign v_16342 = v_2958 | ~v_3072;
assign v_16344 = v_2829 | v_16343;
assign v_16345 = v_2814 | ~v_2900;
assign v_16347 = v_2695 | v_16346;
assign v_16348 = v_2669 | ~v_2768;
assign v_16350 = v_2543 | v_16349;
assign v_16351 = v_2528 | ~v_2614;
assign v_16353 = v_2407 | v_16352;
assign v_16354 = v_2380 | ~v_2482;
assign v_16356 = v_2255 | v_16355;
assign v_16357 = v_2240 | ~v_2326;
assign v_16359 = v_2121 | v_16358;
assign v_16360 = v_2097 | ~v_2194;
assign v_16362 = v_1973 | v_16361;
assign v_16363 = v_1958 | ~v_2044;
assign v_16365 = v_1835 | v_16364;
assign v_16366 = v_1804 | ~v_1912;
assign v_16368 = v_1677 | v_16367;
assign v_16369 = v_1662 | ~v_1748;
assign v_16371 = v_1543 | v_16370;
assign v_16372 = v_1518 | ~v_1616;
assign v_16374 = v_1393 | v_16373;
assign v_16375 = v_1378 | ~v_1464;
assign v_16377 = v_1257 | v_16376;
assign v_16378 = v_1230 | ~v_1332;
assign v_16380 = v_1105 | v_16379;
assign v_16381 = v_1090 | ~v_1176;
assign v_16383 = v_971 | v_16382;
assign v_16384 = v_947 | ~v_1044;
assign v_16386 = v_827 | v_16385;
assign v_16387 = v_811 | ~v_898;
assign v_16389 = v_658 | v_16388;
assign v_16390 = v_359 | ~v_771;
assign v_16392 = v_16202 | v_16391;
assign v_16395 = v_16393 | v_16394;
assign v_16398 = v_16396 | v_16397;
assign v_16401 = v_16399 | v_16400;
assign v_16404 = v_16402 | v_16403;
assign v_16407 = v_16405 | v_16406;
assign v_16410 = v_16408 | v_16409;
assign v_16413 = v_16411 | v_16412;
assign v_16416 = v_16414 | v_16415;
assign v_16419 = v_16417 | v_16418;
assign v_16422 = v_16420 | v_16421;
assign v_16425 = v_16423 | v_16424;
assign v_16428 = v_16426 | v_16427;
assign v_16431 = v_16429 | v_16430;
assign v_16434 = v_16432 | v_16433;
assign v_16437 = v_16435 | v_16436;
assign v_16440 = v_16438 | v_16439;
assign v_16443 = v_16441 | v_16442;
assign v_16446 = v_16444 | v_16445;
assign v_16449 = v_16447 | v_16448;
assign v_16452 = v_16450 | v_16451;
assign v_16455 = v_16453 | v_16454;
assign v_16458 = v_16456 | v_16457;
assign v_16461 = v_16459 | v_16460;
assign v_16464 = v_16462 | v_16463;
assign v_16467 = v_16465 | v_16466;
assign v_16470 = v_16468 | v_16469;
assign v_16473 = v_16471 | v_16472;
assign v_16476 = v_16474 | v_16475;
assign v_16479 = v_16477 | v_16478;
assign v_16482 = v_16480 | v_16481;
assign v_16485 = v_16483 | v_16484;
assign v_16488 = v_16486 | v_16487;
assign v_16491 = v_16489 | v_16490;
assign v_16494 = v_16492 | v_16493;
assign v_16497 = v_16495 | v_16496;
assign v_16500 = v_16498 | v_16499;
assign v_16503 = v_16501 | v_16502;
assign v_16506 = v_16504 | v_16505;
assign v_16509 = v_16507 | v_16508;
assign v_16512 = v_16510 | v_16511;
assign v_16515 = v_16513 | v_16514;
assign v_16518 = v_16516 | v_16517;
assign v_16521 = v_16519 | v_16520;
assign v_16524 = v_16522 | v_16523;
assign v_16527 = v_16525 | v_16526;
assign v_16530 = v_16528 | v_16529;
assign v_16533 = v_16531 | v_16532;
assign v_16536 = v_16534 | v_16535;
assign v_16539 = v_16537 | v_16538;
assign v_16542 = v_16540 | v_16541;
assign v_16545 = v_16543 | v_16544;
assign v_16548 = v_16546 | v_16547;
assign v_16551 = v_16549 | v_16550;
assign v_16554 = v_16552 | v_16553;
assign v_16557 = v_16555 | v_16556;
assign v_16560 = v_16558 | v_16559;
assign v_16563 = v_16561 | v_16562;
assign v_16566 = v_16564 | v_16565;
assign v_16569 = v_16567 | v_16568;
assign v_16572 = v_16570 | v_16571;
assign v_16575 = v_16573 | v_16574;
assign v_16578 = v_16576 | v_16577;
assign v_16581 = v_16579 | v_16580;
assign v_16582 = v_16392 | v_16581;
assign v_16583 = v_13540 | v_16582;
assign v_16584 = v_15063 | v_16583;
assign v_16585 = v_10462 | v_16584;
assign v_16589 = v_16587 | v_16588;
assign v_16592 = v_16590 | v_16591;
assign v_16595 = v_16593 | v_16594;
assign v_16598 = v_16596 | v_16597;
assign v_16601 = v_16599 | v_16600;
assign v_16604 = v_16602 | v_16603;
assign v_16607 = v_16605 | v_16606;
assign v_16610 = v_16608 | v_16609;
assign v_16613 = v_16611 | v_16612;
assign v_16616 = v_16614 | v_16615;
assign v_16619 = v_16617 | v_16618;
assign v_16622 = v_16620 | v_16621;
assign v_16625 = v_16623 | v_16624;
assign v_16628 = v_16626 | v_16627;
assign v_16631 = v_16629 | v_16630;
assign v_16634 = v_16632 | v_16633;
assign v_16637 = v_16635 | v_16636;
assign v_16640 = v_16638 | v_16639;
assign v_16643 = v_16641 | v_16642;
assign v_16646 = v_16644 | v_16645;
assign v_16649 = v_16647 | v_16648;
assign v_16652 = v_16650 | v_16651;
assign v_16655 = v_16653 | v_16654;
assign v_16658 = v_16656 | v_16657;
assign v_16661 = v_16659 | v_16660;
assign v_16664 = v_16662 | v_16663;
assign v_16667 = v_16665 | v_16666;
assign v_16670 = v_16668 | v_16669;
assign v_16673 = v_16671 | v_16672;
assign v_16676 = v_16674 | v_16675;
assign v_16679 = v_16677 | v_16678;
assign v_16682 = v_16680 | v_16681;
assign v_16685 = v_16683 | v_16684;
assign v_16688 = v_16686 | v_16687;
assign v_16691 = v_16689 | v_16690;
assign v_16694 = v_16692 | v_16693;
assign v_16697 = v_16695 | v_16696;
assign v_16700 = v_16698 | v_16699;
assign v_16703 = v_16701 | v_16702;
assign v_16706 = v_16704 | v_16705;
assign v_16709 = v_16707 | v_16708;
assign v_16712 = v_16710 | v_16711;
assign v_16715 = v_16713 | v_16714;
assign v_16718 = v_16716 | v_16717;
assign v_16721 = v_16719 | v_16720;
assign v_16724 = v_16722 | v_16723;
assign v_16727 = v_16725 | v_16726;
assign v_16730 = v_16728 | v_16729;
assign v_16733 = v_16731 | v_16732;
assign v_16736 = v_16734 | v_16735;
assign v_16739 = v_16737 | v_16738;
assign v_16742 = v_16740 | v_16741;
assign v_16745 = v_16743 | v_16744;
assign v_16748 = v_16746 | v_16747;
assign v_16751 = v_16749 | v_16750;
assign v_16754 = v_16752 | v_16753;
assign v_16757 = v_16755 | v_16756;
assign v_16760 = v_16758 | v_16759;
assign v_16763 = v_16761 | v_16762;
assign v_16766 = v_16764 | v_16765;
assign v_16769 = v_16767 | v_16768;
assign v_16772 = v_16770 | v_16771;
assign v_16775 = v_16773 | v_16774;
assign v_16778 = v_16776 | v_16777;
assign v_16781 = v_16779 | v_16780;
assign v_16784 = v_16782 | v_16783;
assign v_16787 = v_16785 | v_16786;
assign v_16790 = v_16788 | v_16789;
assign v_16793 = v_16791 | v_16792;
assign v_16796 = v_16794 | v_16795;
assign v_16799 = v_16797 | v_16798;
assign v_16802 = v_16800 | v_16801;
assign v_16805 = v_16803 | v_16804;
assign v_16808 = v_16806 | v_16807;
assign v_16811 = v_16809 | v_16810;
assign v_16814 = v_16812 | v_16813;
assign v_16817 = v_16815 | v_16816;
assign v_16820 = v_16818 | v_16819;
assign v_16823 = v_16821 | v_16822;
assign v_16826 = v_16824 | v_16825;
assign v_16829 = v_16827 | v_16828;
assign v_16832 = v_16830 | v_16831;
assign v_16835 = v_16833 | v_16834;
assign v_16838 = v_16836 | v_16837;
assign v_16841 = v_16839 | v_16840;
assign v_16844 = v_16842 | v_16843;
assign v_16847 = v_16845 | v_16846;
assign v_16850 = v_16848 | v_16849;
assign v_16853 = v_16851 | v_16852;
assign v_16856 = v_16854 | v_16855;
assign v_16859 = v_16857 | v_16858;
assign v_16862 = v_16860 | v_16861;
assign v_16865 = v_16863 | v_16864;
assign v_16868 = v_16866 | v_16867;
assign v_16871 = v_16869 | v_16870;
assign v_16874 = v_16872 | v_16873;
assign v_16877 = v_16875 | v_16876;
assign v_16880 = v_16878 | v_16879;
assign v_16883 = v_16881 | v_16882;
assign v_16886 = v_16884 | v_16885;
assign v_16889 = v_16887 | v_16888;
assign v_16892 = v_16890 | v_16891;
assign v_16895 = v_16893 | v_16894;
assign v_16898 = v_16896 | v_16897;
assign v_16901 = v_16899 | v_16900;
assign v_16904 = v_16902 | v_16903;
assign v_16907 = v_16905 | v_16906;
assign v_16910 = v_16908 | v_16909;
assign v_16913 = v_16911 | v_16912;
assign v_16916 = v_16914 | v_16915;
assign v_16919 = v_16917 | v_16918;
assign v_16922 = v_16920 | v_16921;
assign v_16925 = v_16923 | v_16924;
assign v_16928 = v_16926 | v_16927;
assign v_16931 = v_16929 | v_16930;
assign v_16934 = v_16932 | v_16933;
assign v_16937 = v_16935 | v_16936;
assign v_16940 = v_16938 | v_16939;
assign v_16943 = v_16941 | v_16942;
assign v_16946 = v_16944 | v_16945;
assign v_16949 = v_16947 | v_16948;
assign v_16952 = v_16950 | v_16951;
assign v_16953 = v_16769 | v_16952;
assign v_16956 = v_16954 | v_16955;
assign v_16959 = v_16957 | v_16958;
assign v_16962 = v_16960 | v_16961;
assign v_16965 = v_16963 | v_16964;
assign v_16968 = v_16966 | v_16967;
assign v_16971 = v_16969 | v_16970;
assign v_16974 = v_16972 | v_16973;
assign v_16977 = v_16975 | v_16976;
assign v_16980 = v_16978 | v_16979;
assign v_16983 = v_16981 | v_16982;
assign v_16986 = v_16984 | v_16985;
assign v_16989 = v_16987 | v_16988;
assign v_16992 = v_16990 | v_16991;
assign v_16995 = v_16993 | v_16994;
assign v_16998 = v_16996 | v_16997;
assign v_17001 = v_16999 | v_17000;
assign v_17004 = v_17002 | v_17003;
assign v_17007 = v_17005 | v_17006;
assign v_17010 = v_17008 | v_17009;
assign v_17013 = v_17011 | v_17012;
assign v_17016 = v_17014 | v_17015;
assign v_17019 = v_17017 | v_17018;
assign v_17022 = v_17020 | v_17021;
assign v_17025 = v_17023 | v_17024;
assign v_17028 = v_17026 | v_17027;
assign v_17031 = v_17029 | v_17030;
assign v_17034 = v_17032 | v_17033;
assign v_17037 = v_17035 | v_17036;
assign v_17040 = v_17038 | v_17039;
assign v_17043 = v_17041 | v_17042;
assign v_17046 = v_17044 | v_17045;
assign v_17049 = v_17047 | v_17048;
assign v_17052 = v_17050 | v_17051;
assign v_17055 = v_17053 | v_17054;
assign v_17058 = v_17056 | v_17057;
assign v_17061 = v_17059 | v_17060;
assign v_17064 = v_17062 | v_17063;
assign v_17067 = v_17065 | v_17066;
assign v_17070 = v_17068 | v_17069;
assign v_17073 = v_17071 | v_17072;
assign v_17076 = v_17074 | v_17075;
assign v_17079 = v_17077 | v_17078;
assign v_17082 = v_17080 | v_17081;
assign v_17085 = v_17083 | v_17084;
assign v_17088 = v_17086 | v_17087;
assign v_17091 = v_17089 | v_17090;
assign v_17094 = v_17092 | v_17093;
assign v_17097 = v_17095 | v_17096;
assign v_17100 = v_17098 | v_17099;
assign v_17103 = v_17101 | v_17102;
assign v_17106 = v_17104 | v_17105;
assign v_17109 = v_17107 | v_17108;
assign v_17112 = v_17110 | v_17111;
assign v_17115 = v_17113 | v_17114;
assign v_17118 = v_17116 | v_17117;
assign v_17121 = v_17119 | v_17120;
assign v_17124 = v_17122 | v_17123;
assign v_17127 = v_17125 | v_17126;
assign v_17130 = v_17128 | v_17129;
assign v_17133 = v_17131 | v_17132;
assign v_17136 = v_17134 | v_17135;
assign v_17137 = v_16953 | v_17136;
assign v_17140 = v_17138 | v_17139;
assign v_17143 = v_17141 | v_17142;
assign v_17146 = v_17144 | v_17145;
assign v_17149 = v_17147 | v_17148;
assign v_17152 = v_17150 | v_17151;
assign v_17155 = v_17153 | v_17154;
assign v_17158 = v_17156 | v_17157;
assign v_17161 = v_17159 | v_17160;
assign v_17164 = v_17162 | v_17163;
assign v_17167 = v_17165 | v_17166;
assign v_17170 = v_17168 | v_17169;
assign v_17173 = v_17171 | v_17172;
assign v_17176 = v_17174 | v_17175;
assign v_17179 = v_17177 | v_17178;
assign v_17182 = v_17180 | v_17181;
assign v_17185 = v_17183 | v_17184;
assign v_17188 = v_17186 | v_17187;
assign v_17191 = v_17189 | v_17190;
assign v_17194 = v_17192 | v_17193;
assign v_17197 = v_17195 | v_17196;
assign v_17200 = v_17198 | v_17199;
assign v_17203 = v_17201 | v_17202;
assign v_17206 = v_17204 | v_17205;
assign v_17209 = v_17207 | v_17208;
assign v_17212 = v_17210 | v_17211;
assign v_17215 = v_17213 | v_17214;
assign v_17218 = v_17216 | v_17217;
assign v_17221 = v_17219 | v_17220;
assign v_17224 = v_17222 | v_17223;
assign v_17227 = v_17225 | v_17226;
assign v_17230 = v_17228 | v_17229;
assign v_17233 = v_17231 | v_17232;
assign v_17236 = v_17234 | v_17235;
assign v_17239 = v_17237 | v_17238;
assign v_17242 = v_17240 | v_17241;
assign v_17245 = v_17243 | v_17244;
assign v_17248 = v_17246 | v_17247;
assign v_17251 = v_17249 | v_17250;
assign v_17254 = v_17252 | v_17253;
assign v_17257 = v_17255 | v_17256;
assign v_17260 = v_17258 | v_17259;
assign v_17263 = v_17261 | v_17262;
assign v_17266 = v_17264 | v_17265;
assign v_17269 = v_17267 | v_17268;
assign v_17272 = v_17270 | v_17271;
assign v_17275 = v_17273 | v_17274;
assign v_17278 = v_17276 | v_17277;
assign v_17281 = v_17279 | v_17280;
assign v_17284 = v_17282 | v_17283;
assign v_17287 = v_17285 | v_17286;
assign v_17290 = v_17288 | v_17289;
assign v_17293 = v_17291 | v_17292;
assign v_17296 = v_17294 | v_17295;
assign v_17299 = v_17297 | v_17298;
assign v_17302 = v_17300 | v_17301;
assign v_17305 = v_17303 | v_17304;
assign v_17308 = v_17306 | v_17307;
assign v_17311 = v_17309 | v_17310;
assign v_17314 = v_17312 | v_17313;
assign v_17317 = v_17315 | v_17316;
assign v_17320 = v_17318 | v_17319;
assign v_17321 = v_17137 | v_17320;
assign v_17324 = v_17322 | v_17323;
assign v_17327 = v_17325 | v_17326;
assign v_17330 = v_17328 | v_17329;
assign v_17333 = v_17331 | v_17332;
assign v_17336 = v_17334 | v_17335;
assign v_17339 = v_17337 | v_17338;
assign v_17342 = v_17340 | v_17341;
assign v_17345 = v_17343 | v_17344;
assign v_17348 = v_17346 | v_17347;
assign v_17351 = v_17349 | v_17350;
assign v_17354 = v_17352 | v_17353;
assign v_17357 = v_17355 | v_17356;
assign v_17360 = v_17358 | v_17359;
assign v_17363 = v_17361 | v_17362;
assign v_17366 = v_17364 | v_17365;
assign v_17369 = v_17367 | v_17368;
assign v_17372 = v_17370 | v_17371;
assign v_17375 = v_17373 | v_17374;
assign v_17378 = v_17376 | v_17377;
assign v_17381 = v_17379 | v_17380;
assign v_17384 = v_17382 | v_17383;
assign v_17387 = v_17385 | v_17386;
assign v_17390 = v_17388 | v_17389;
assign v_17393 = v_17391 | v_17392;
assign v_17396 = v_17394 | v_17395;
assign v_17399 = v_17397 | v_17398;
assign v_17402 = v_17400 | v_17401;
assign v_17405 = v_17403 | v_17404;
assign v_17408 = v_17406 | v_17407;
assign v_17411 = v_17409 | v_17410;
assign v_17414 = v_17412 | v_17413;
assign v_17417 = v_17415 | v_17416;
assign v_17420 = v_17418 | v_17419;
assign v_17423 = v_17421 | v_17422;
assign v_17426 = v_17424 | v_17425;
assign v_17429 = v_17427 | v_17428;
assign v_17432 = v_17430 | v_17431;
assign v_17435 = v_17433 | v_17434;
assign v_17438 = v_17436 | v_17437;
assign v_17441 = v_17439 | v_17440;
assign v_17444 = v_17442 | v_17443;
assign v_17447 = v_17445 | v_17446;
assign v_17450 = v_17448 | v_17449;
assign v_17453 = v_17451 | v_17452;
assign v_17456 = v_17454 | v_17455;
assign v_17459 = v_17457 | v_17458;
assign v_17462 = v_17460 | v_17461;
assign v_17465 = v_17463 | v_17464;
assign v_17468 = v_17466 | v_17467;
assign v_17471 = v_17469 | v_17470;
assign v_17474 = v_17472 | v_17473;
assign v_17477 = v_17475 | v_17476;
assign v_17480 = v_17478 | v_17479;
assign v_17483 = v_17481 | v_17482;
assign v_17486 = v_17484 | v_17485;
assign v_17489 = v_17487 | v_17488;
assign v_17492 = v_17490 | v_17491;
assign v_17495 = v_17493 | v_17494;
assign v_17498 = v_17496 | v_17497;
assign v_17501 = v_17499 | v_17500;
assign v_17504 = v_17502 | v_17503;
assign v_17505 = v_17321 | v_17504;
assign v_17508 = v_17506 | v_17507;
assign v_17511 = v_17509 | v_17510;
assign v_17514 = v_17512 | v_17513;
assign v_17517 = v_17515 | v_17516;
assign v_17520 = v_17518 | v_17519;
assign v_17523 = v_17521 | v_17522;
assign v_17526 = v_17524 | v_17525;
assign v_17529 = v_17527 | v_17528;
assign v_17532 = v_17530 | v_17531;
assign v_17535 = v_17533 | v_17534;
assign v_17538 = v_17536 | v_17537;
assign v_17541 = v_17539 | v_17540;
assign v_17544 = v_17542 | v_17543;
assign v_17547 = v_17545 | v_17546;
assign v_17550 = v_17548 | v_17549;
assign v_17553 = v_17551 | v_17552;
assign v_17556 = v_17554 | v_17555;
assign v_17559 = v_17557 | v_17558;
assign v_17562 = v_17560 | v_17561;
assign v_17565 = v_17563 | v_17564;
assign v_17568 = v_17566 | v_17567;
assign v_17571 = v_17569 | v_17570;
assign v_17574 = v_17572 | v_17573;
assign v_17577 = v_17575 | v_17576;
assign v_17580 = v_17578 | v_17579;
assign v_17583 = v_17581 | v_17582;
assign v_17586 = v_17584 | v_17585;
assign v_17589 = v_17587 | v_17588;
assign v_17592 = v_17590 | v_17591;
assign v_17595 = v_17593 | v_17594;
assign v_17598 = v_17596 | v_17597;
assign v_17601 = v_17599 | v_17600;
assign v_17604 = v_17602 | v_17603;
assign v_17607 = v_17605 | v_17606;
assign v_17610 = v_17608 | v_17609;
assign v_17613 = v_17611 | v_17612;
assign v_17616 = v_17614 | v_17615;
assign v_17619 = v_17617 | v_17618;
assign v_17622 = v_17620 | v_17621;
assign v_17625 = v_17623 | v_17624;
assign v_17628 = v_17626 | v_17627;
assign v_17631 = v_17629 | v_17630;
assign v_17634 = v_17632 | v_17633;
assign v_17637 = v_17635 | v_17636;
assign v_17640 = v_17638 | v_17639;
assign v_17643 = v_17641 | v_17642;
assign v_17646 = v_17644 | v_17645;
assign v_17649 = v_17647 | v_17648;
assign v_17652 = v_17650 | v_17651;
assign v_17655 = v_17653 | v_17654;
assign v_17658 = v_17656 | v_17657;
assign v_17661 = v_17659 | v_17660;
assign v_17664 = v_17662 | v_17663;
assign v_17667 = v_17665 | v_17666;
assign v_17670 = v_17668 | v_17669;
assign v_17673 = v_17671 | v_17672;
assign v_17676 = v_17674 | v_17675;
assign v_17679 = v_17677 | v_17678;
assign v_17682 = v_17680 | v_17681;
assign v_17685 = v_17683 | v_17684;
assign v_17688 = v_17686 | v_17687;
assign v_17689 = v_17505 | v_17688;
assign v_17692 = v_17690 | v_17691;
assign v_17695 = v_17693 | v_17694;
assign v_17698 = v_17696 | v_17697;
assign v_17701 = v_17699 | v_17700;
assign v_17704 = v_17702 | v_17703;
assign v_17707 = v_17705 | v_17706;
assign v_17710 = v_17708 | v_17709;
assign v_17713 = v_17711 | v_17712;
assign v_17716 = v_17714 | v_17715;
assign v_17719 = v_17717 | v_17718;
assign v_17722 = v_17720 | v_17721;
assign v_17725 = v_17723 | v_17724;
assign v_17728 = v_17726 | v_17727;
assign v_17731 = v_17729 | v_17730;
assign v_17734 = v_17732 | v_17733;
assign v_17737 = v_17735 | v_17736;
assign v_17740 = v_17738 | v_17739;
assign v_17743 = v_17741 | v_17742;
assign v_17746 = v_17744 | v_17745;
assign v_17749 = v_17747 | v_17748;
assign v_17752 = v_17750 | v_17751;
assign v_17755 = v_17753 | v_17754;
assign v_17758 = v_17756 | v_17757;
assign v_17761 = v_17759 | v_17760;
assign v_17764 = v_17762 | v_17763;
assign v_17767 = v_17765 | v_17766;
assign v_17770 = v_17768 | v_17769;
assign v_17773 = v_17771 | v_17772;
assign v_17776 = v_17774 | v_17775;
assign v_17779 = v_17777 | v_17778;
assign v_17782 = v_17780 | v_17781;
assign v_17785 = v_17783 | v_17784;
assign v_17788 = v_17786 | v_17787;
assign v_17791 = v_17789 | v_17790;
assign v_17794 = v_17792 | v_17793;
assign v_17797 = v_17795 | v_17796;
assign v_17800 = v_17798 | v_17799;
assign v_17803 = v_17801 | v_17802;
assign v_17806 = v_17804 | v_17805;
assign v_17809 = v_17807 | v_17808;
assign v_17812 = v_17810 | v_17811;
assign v_17815 = v_17813 | v_17814;
assign v_17818 = v_17816 | v_17817;
assign v_17821 = v_17819 | v_17820;
assign v_17824 = v_17822 | v_17823;
assign v_17827 = v_17825 | v_17826;
assign v_17830 = v_17828 | v_17829;
assign v_17833 = v_17831 | v_17832;
assign v_17836 = v_17834 | v_17835;
assign v_17839 = v_17837 | v_17838;
assign v_17842 = v_17840 | v_17841;
assign v_17845 = v_17843 | v_17844;
assign v_17848 = v_17846 | v_17847;
assign v_17851 = v_17849 | v_17850;
assign v_17854 = v_17852 | v_17853;
assign v_17857 = v_17855 | v_17856;
assign v_17860 = v_17858 | v_17859;
assign v_17863 = v_17861 | v_17862;
assign v_17866 = v_17864 | v_17865;
assign v_17869 = v_17867 | v_17868;
assign v_17872 = v_17870 | v_17871;
assign v_17873 = v_17689 | v_17872;
assign v_17876 = v_17874 | v_17875;
assign v_17879 = v_17877 | v_17878;
assign v_17882 = v_17880 | v_17881;
assign v_17885 = v_17883 | v_17884;
assign v_17888 = v_17886 | v_17887;
assign v_17891 = v_17889 | v_17890;
assign v_17894 = v_17892 | v_17893;
assign v_17897 = v_17895 | v_17896;
assign v_17900 = v_17898 | v_17899;
assign v_17903 = v_17901 | v_17902;
assign v_17906 = v_17904 | v_17905;
assign v_17909 = v_17907 | v_17908;
assign v_17912 = v_17910 | v_17911;
assign v_17915 = v_17913 | v_17914;
assign v_17918 = v_17916 | v_17917;
assign v_17921 = v_17919 | v_17920;
assign v_17924 = v_17922 | v_17923;
assign v_17927 = v_17925 | v_17926;
assign v_17930 = v_17928 | v_17929;
assign v_17933 = v_17931 | v_17932;
assign v_17936 = v_17934 | v_17935;
assign v_17939 = v_17937 | v_17938;
assign v_17942 = v_17940 | v_17941;
assign v_17945 = v_17943 | v_17944;
assign v_17948 = v_17946 | v_17947;
assign v_17951 = v_17949 | v_17950;
assign v_17954 = v_17952 | v_17953;
assign v_17957 = v_17955 | v_17956;
assign v_17960 = v_17958 | v_17959;
assign v_17963 = v_17961 | v_17962;
assign v_17966 = v_17964 | v_17965;
assign v_17969 = v_17967 | v_17968;
assign v_17972 = v_17970 | v_17971;
assign v_17975 = v_17973 | v_17974;
assign v_17978 = v_17976 | v_17977;
assign v_17981 = v_17979 | v_17980;
assign v_17984 = v_17982 | v_17983;
assign v_17987 = v_17985 | v_17986;
assign v_17990 = v_17988 | v_17989;
assign v_17993 = v_17991 | v_17992;
assign v_17996 = v_17994 | v_17995;
assign v_17999 = v_17997 | v_17998;
assign v_18002 = v_18000 | v_18001;
assign v_18005 = v_18003 | v_18004;
assign v_18008 = v_18006 | v_18007;
assign v_18011 = v_18009 | v_18010;
assign v_18014 = v_18012 | v_18013;
assign v_18017 = v_18015 | v_18016;
assign v_18020 = v_18018 | v_18019;
assign v_18023 = v_18021 | v_18022;
assign v_18026 = v_18024 | v_18025;
assign v_18029 = v_18027 | v_18028;
assign v_18032 = v_18030 | v_18031;
assign v_18035 = v_18033 | v_18034;
assign v_18038 = v_18036 | v_18037;
assign v_18041 = v_18039 | v_18040;
assign v_18044 = v_18042 | v_18043;
assign v_18047 = v_18045 | v_18046;
assign v_18050 = v_18048 | v_18049;
assign v_18053 = v_18051 | v_18052;
assign v_18056 = v_18054 | v_18055;
assign v_18057 = v_17873 | v_18056;
assign v_18060 = v_18058 | v_18059;
assign v_18063 = v_18061 | v_18062;
assign v_18066 = v_18064 | v_18065;
assign v_18069 = v_18067 | v_18068;
assign v_18072 = v_18070 | v_18071;
assign v_18075 = v_18073 | v_18074;
assign v_18078 = v_18076 | v_18077;
assign v_18081 = v_18079 | v_18080;
assign v_18084 = v_18082 | v_18083;
assign v_18087 = v_18085 | v_18086;
assign v_18090 = v_18088 | v_18089;
assign v_18093 = v_18091 | v_18092;
assign v_18096 = v_18094 | v_18095;
assign v_18099 = v_18097 | v_18098;
assign v_18102 = v_18100 | v_18101;
assign v_18105 = v_18103 | v_18104;
assign v_18108 = v_18106 | v_18107;
assign v_18111 = v_18109 | v_18110;
assign v_18114 = v_18112 | v_18113;
assign v_18117 = v_18115 | v_18116;
assign v_18120 = v_18118 | v_18119;
assign v_18123 = v_18121 | v_18122;
assign v_18126 = v_18124 | v_18125;
assign v_18129 = v_18127 | v_18128;
assign v_18132 = v_18130 | v_18131;
assign v_18135 = v_18133 | v_18134;
assign v_18138 = v_18136 | v_18137;
assign v_18141 = v_18139 | v_18140;
assign v_18144 = v_18142 | v_18143;
assign v_18147 = v_18145 | v_18146;
assign v_18150 = v_18148 | v_18149;
assign v_18153 = v_18151 | v_18152;
assign v_18156 = v_18154 | v_18155;
assign v_18159 = v_18157 | v_18158;
assign v_18162 = v_18160 | v_18161;
assign v_18165 = v_18163 | v_18164;
assign v_18168 = v_18166 | v_18167;
assign v_18171 = v_18169 | v_18170;
assign v_18174 = v_18172 | v_18173;
assign v_18177 = v_18175 | v_18176;
assign v_18180 = v_18178 | v_18179;
assign v_18183 = v_18181 | v_18182;
assign v_18186 = v_18184 | v_18185;
assign v_18189 = v_18187 | v_18188;
assign v_18192 = v_18190 | v_18191;
assign v_18195 = v_18193 | v_18194;
assign v_18198 = v_18196 | v_18197;
assign v_18201 = v_18199 | v_18200;
assign v_18204 = v_18202 | v_18203;
assign v_18207 = v_18205 | v_18206;
assign v_18210 = v_18208 | v_18209;
assign v_18213 = v_18211 | v_18212;
assign v_18216 = v_18214 | v_18215;
assign v_18219 = v_18217 | v_18218;
assign v_18222 = v_18220 | v_18221;
assign v_18225 = v_18223 | v_18224;
assign v_18228 = v_18226 | v_18227;
assign v_18231 = v_18229 | v_18230;
assign v_18234 = v_18232 | v_18233;
assign v_18237 = v_18235 | v_18236;
assign v_18240 = v_18238 | v_18239;
assign v_18243 = v_18241 | v_18242;
assign v_18246 = v_18244 | v_18245;
assign v_18249 = v_18247 | v_18248;
assign v_18252 = v_18250 | v_18251;
assign v_18255 = v_18253 | v_18254;
assign v_18258 = v_18256 | v_18257;
assign v_18261 = v_18259 | v_18260;
assign v_18264 = v_18262 | v_18263;
assign v_18267 = v_18265 | v_18266;
assign v_18270 = v_18268 | v_18269;
assign v_18273 = v_18271 | v_18272;
assign v_18276 = v_18274 | v_18275;
assign v_18279 = v_18277 | v_18278;
assign v_18282 = v_18280 | v_18281;
assign v_18285 = v_18283 | v_18284;
assign v_18288 = v_18286 | v_18287;
assign v_18291 = v_18289 | v_18290;
assign v_18294 = v_18292 | v_18293;
assign v_18297 = v_18295 | v_18296;
assign v_18300 = v_18298 | v_18299;
assign v_18303 = v_18301 | v_18302;
assign v_18306 = v_18304 | v_18305;
assign v_18309 = v_18307 | v_18308;
assign v_18312 = v_18310 | v_18311;
assign v_18315 = v_18313 | v_18314;
assign v_18318 = v_18316 | v_18317;
assign v_18321 = v_18319 | v_18320;
assign v_18324 = v_18322 | v_18323;
assign v_18327 = v_18325 | v_18326;
assign v_18330 = v_18328 | v_18329;
assign v_18333 = v_18331 | v_18332;
assign v_18336 = v_18334 | v_18335;
assign v_18339 = v_18337 | v_18338;
assign v_18342 = v_18340 | v_18341;
assign v_18345 = v_18343 | v_18344;
assign v_18348 = v_18346 | v_18347;
assign v_18351 = v_18349 | v_18350;
assign v_18354 = v_18352 | v_18353;
assign v_18357 = v_18355 | v_18356;
assign v_18360 = v_18358 | v_18359;
assign v_18363 = v_18361 | v_18362;
assign v_18366 = v_18364 | v_18365;
assign v_18369 = v_18367 | v_18368;
assign v_18372 = v_18370 | v_18371;
assign v_18375 = v_18373 | v_18374;
assign v_18378 = v_18376 | v_18377;
assign v_18381 = v_18379 | v_18380;
assign v_18384 = v_18382 | v_18383;
assign v_18387 = v_18385 | v_18386;
assign v_18390 = v_18388 | v_18389;
assign v_18393 = v_18391 | v_18392;
assign v_18396 = v_18394 | v_18395;
assign v_18399 = v_18397 | v_18398;
assign v_18402 = v_18400 | v_18401;
assign v_18405 = v_18403 | v_18404;
assign v_18408 = v_18406 | v_18407;
assign v_18411 = v_18409 | v_18410;
assign v_18414 = v_18412 | v_18413;
assign v_18417 = v_18415 | v_18416;
assign v_18420 = v_18418 | v_18419;
assign v_18423 = v_18421 | v_18422;
assign v_18426 = v_18424 | v_18425;
assign v_18429 = v_18427 | v_18428;
assign v_18430 = v_18243 | v_18429;
assign v_18433 = v_18431 | v_18432;
assign v_18436 = v_18434 | v_18435;
assign v_18439 = v_18437 | v_18438;
assign v_18442 = v_18440 | v_18441;
assign v_18445 = v_18443 | v_18444;
assign v_18448 = v_18446 | v_18447;
assign v_18451 = v_18449 | v_18450;
assign v_18454 = v_18452 | v_18453;
assign v_18457 = v_18455 | v_18456;
assign v_18460 = v_18458 | v_18459;
assign v_18463 = v_18461 | v_18462;
assign v_18466 = v_18464 | v_18465;
assign v_18469 = v_18467 | v_18468;
assign v_18472 = v_18470 | v_18471;
assign v_18475 = v_18473 | v_18474;
assign v_18478 = v_18476 | v_18477;
assign v_18481 = v_18479 | v_18480;
assign v_18484 = v_18482 | v_18483;
assign v_18487 = v_18485 | v_18486;
assign v_18490 = v_18488 | v_18489;
assign v_18493 = v_18491 | v_18492;
assign v_18496 = v_18494 | v_18495;
assign v_18499 = v_18497 | v_18498;
assign v_18502 = v_18500 | v_18501;
assign v_18505 = v_18503 | v_18504;
assign v_18508 = v_18506 | v_18507;
assign v_18511 = v_18509 | v_18510;
assign v_18514 = v_18512 | v_18513;
assign v_18517 = v_18515 | v_18516;
assign v_18520 = v_18518 | v_18519;
assign v_18523 = v_18521 | v_18522;
assign v_18526 = v_18524 | v_18525;
assign v_18529 = v_18527 | v_18528;
assign v_18532 = v_18530 | v_18531;
assign v_18535 = v_18533 | v_18534;
assign v_18538 = v_18536 | v_18537;
assign v_18541 = v_18539 | v_18540;
assign v_18544 = v_18542 | v_18543;
assign v_18547 = v_18545 | v_18546;
assign v_18550 = v_18548 | v_18549;
assign v_18553 = v_18551 | v_18552;
assign v_18556 = v_18554 | v_18555;
assign v_18559 = v_18557 | v_18558;
assign v_18562 = v_18560 | v_18561;
assign v_18565 = v_18563 | v_18564;
assign v_18568 = v_18566 | v_18567;
assign v_18571 = v_18569 | v_18570;
assign v_18574 = v_18572 | v_18573;
assign v_18577 = v_18575 | v_18576;
assign v_18580 = v_18578 | v_18579;
assign v_18583 = v_18581 | v_18582;
assign v_18586 = v_18584 | v_18585;
assign v_18589 = v_18587 | v_18588;
assign v_18592 = v_18590 | v_18591;
assign v_18595 = v_18593 | v_18594;
assign v_18598 = v_18596 | v_18597;
assign v_18601 = v_18599 | v_18600;
assign v_18604 = v_18602 | v_18603;
assign v_18607 = v_18605 | v_18606;
assign v_18610 = v_18608 | v_18609;
assign v_18613 = v_18611 | v_18612;
assign v_18616 = v_18614 | v_18615;
assign v_18617 = v_18430 | v_18616;
assign v_18620 = v_18618 | v_18619;
assign v_18623 = v_18621 | v_18622;
assign v_18626 = v_18624 | v_18625;
assign v_18629 = v_18627 | v_18628;
assign v_18632 = v_18630 | v_18631;
assign v_18635 = v_18633 | v_18634;
assign v_18638 = v_18636 | v_18637;
assign v_18641 = v_18639 | v_18640;
assign v_18644 = v_18642 | v_18643;
assign v_18647 = v_18645 | v_18646;
assign v_18650 = v_18648 | v_18649;
assign v_18653 = v_18651 | v_18652;
assign v_18656 = v_18654 | v_18655;
assign v_18659 = v_18657 | v_18658;
assign v_18662 = v_18660 | v_18661;
assign v_18665 = v_18663 | v_18664;
assign v_18668 = v_18666 | v_18667;
assign v_18671 = v_18669 | v_18670;
assign v_18674 = v_18672 | v_18673;
assign v_18677 = v_18675 | v_18676;
assign v_18680 = v_18678 | v_18679;
assign v_18683 = v_18681 | v_18682;
assign v_18686 = v_18684 | v_18685;
assign v_18689 = v_18687 | v_18688;
assign v_18692 = v_18690 | v_18691;
assign v_18695 = v_18693 | v_18694;
assign v_18698 = v_18696 | v_18697;
assign v_18701 = v_18699 | v_18700;
assign v_18704 = v_18702 | v_18703;
assign v_18707 = v_18705 | v_18706;
assign v_18710 = v_18708 | v_18709;
assign v_18713 = v_18711 | v_18712;
assign v_18716 = v_18714 | v_18715;
assign v_18719 = v_18717 | v_18718;
assign v_18722 = v_18720 | v_18721;
assign v_18725 = v_18723 | v_18724;
assign v_18728 = v_18726 | v_18727;
assign v_18731 = v_18729 | v_18730;
assign v_18734 = v_18732 | v_18733;
assign v_18737 = v_18735 | v_18736;
assign v_18740 = v_18738 | v_18739;
assign v_18743 = v_18741 | v_18742;
assign v_18746 = v_18744 | v_18745;
assign v_18749 = v_18747 | v_18748;
assign v_18752 = v_18750 | v_18751;
assign v_18755 = v_18753 | v_18754;
assign v_18758 = v_18756 | v_18757;
assign v_18761 = v_18759 | v_18760;
assign v_18764 = v_18762 | v_18763;
assign v_18767 = v_18765 | v_18766;
assign v_18770 = v_18768 | v_18769;
assign v_18773 = v_18771 | v_18772;
assign v_18776 = v_18774 | v_18775;
assign v_18779 = v_18777 | v_18778;
assign v_18782 = v_18780 | v_18781;
assign v_18785 = v_18783 | v_18784;
assign v_18788 = v_18786 | v_18787;
assign v_18791 = v_18789 | v_18790;
assign v_18794 = v_18792 | v_18793;
assign v_18797 = v_18795 | v_18796;
assign v_18800 = v_18798 | v_18799;
assign v_18803 = v_18801 | v_18802;
assign v_18804 = v_18617 | v_18803;
assign v_18807 = v_18805 | v_18806;
assign v_18810 = v_18808 | v_18809;
assign v_18813 = v_18811 | v_18812;
assign v_18816 = v_18814 | v_18815;
assign v_18819 = v_18817 | v_18818;
assign v_18822 = v_18820 | v_18821;
assign v_18825 = v_18823 | v_18824;
assign v_18828 = v_18826 | v_18827;
assign v_18831 = v_18829 | v_18830;
assign v_18834 = v_18832 | v_18833;
assign v_18837 = v_18835 | v_18836;
assign v_18840 = v_18838 | v_18839;
assign v_18843 = v_18841 | v_18842;
assign v_18846 = v_18844 | v_18845;
assign v_18849 = v_18847 | v_18848;
assign v_18852 = v_18850 | v_18851;
assign v_18855 = v_18853 | v_18854;
assign v_18858 = v_18856 | v_18857;
assign v_18861 = v_18859 | v_18860;
assign v_18864 = v_18862 | v_18863;
assign v_18867 = v_18865 | v_18866;
assign v_18870 = v_18868 | v_18869;
assign v_18873 = v_18871 | v_18872;
assign v_18876 = v_18874 | v_18875;
assign v_18879 = v_18877 | v_18878;
assign v_18882 = v_18880 | v_18881;
assign v_18885 = v_18883 | v_18884;
assign v_18888 = v_18886 | v_18887;
assign v_18891 = v_18889 | v_18890;
assign v_18894 = v_18892 | v_18893;
assign v_18897 = v_18895 | v_18896;
assign v_18900 = v_18898 | v_18899;
assign v_18903 = v_18901 | v_18902;
assign v_18906 = v_18904 | v_18905;
assign v_18909 = v_18907 | v_18908;
assign v_18912 = v_18910 | v_18911;
assign v_18915 = v_18913 | v_18914;
assign v_18918 = v_18916 | v_18917;
assign v_18921 = v_18919 | v_18920;
assign v_18924 = v_18922 | v_18923;
assign v_18927 = v_18925 | v_18926;
assign v_18930 = v_18928 | v_18929;
assign v_18933 = v_18931 | v_18932;
assign v_18936 = v_18934 | v_18935;
assign v_18939 = v_18937 | v_18938;
assign v_18942 = v_18940 | v_18941;
assign v_18945 = v_18943 | v_18944;
assign v_18948 = v_18946 | v_18947;
assign v_18951 = v_18949 | v_18950;
assign v_18954 = v_18952 | v_18953;
assign v_18957 = v_18955 | v_18956;
assign v_18960 = v_18958 | v_18959;
assign v_18963 = v_18961 | v_18962;
assign v_18966 = v_18964 | v_18965;
assign v_18969 = v_18967 | v_18968;
assign v_18972 = v_18970 | v_18971;
assign v_18975 = v_18973 | v_18974;
assign v_18978 = v_18976 | v_18977;
assign v_18981 = v_18979 | v_18980;
assign v_18984 = v_18982 | v_18983;
assign v_18987 = v_18985 | v_18986;
assign v_18990 = v_18988 | v_18989;
assign v_18991 = v_18804 | v_18990;
assign v_18994 = v_18992 | v_18993;
assign v_18997 = v_18995 | v_18996;
assign v_19000 = v_18998 | v_18999;
assign v_19003 = v_19001 | v_19002;
assign v_19006 = v_19004 | v_19005;
assign v_19009 = v_19007 | v_19008;
assign v_19012 = v_19010 | v_19011;
assign v_19015 = v_19013 | v_19014;
assign v_19018 = v_19016 | v_19017;
assign v_19021 = v_19019 | v_19020;
assign v_19024 = v_19022 | v_19023;
assign v_19027 = v_19025 | v_19026;
assign v_19030 = v_19028 | v_19029;
assign v_19033 = v_19031 | v_19032;
assign v_19036 = v_19034 | v_19035;
assign v_19039 = v_19037 | v_19038;
assign v_19042 = v_19040 | v_19041;
assign v_19045 = v_19043 | v_19044;
assign v_19048 = v_19046 | v_19047;
assign v_19051 = v_19049 | v_19050;
assign v_19054 = v_19052 | v_19053;
assign v_19057 = v_19055 | v_19056;
assign v_19060 = v_19058 | v_19059;
assign v_19063 = v_19061 | v_19062;
assign v_19066 = v_19064 | v_19065;
assign v_19069 = v_19067 | v_19068;
assign v_19072 = v_19070 | v_19071;
assign v_19075 = v_19073 | v_19074;
assign v_19078 = v_19076 | v_19077;
assign v_19081 = v_19079 | v_19080;
assign v_19084 = v_19082 | v_19083;
assign v_19087 = v_19085 | v_19086;
assign v_19090 = v_19088 | v_19089;
assign v_19093 = v_19091 | v_19092;
assign v_19096 = v_19094 | v_19095;
assign v_19099 = v_19097 | v_19098;
assign v_19102 = v_19100 | v_19101;
assign v_19105 = v_19103 | v_19104;
assign v_19108 = v_19106 | v_19107;
assign v_19111 = v_19109 | v_19110;
assign v_19114 = v_19112 | v_19113;
assign v_19117 = v_19115 | v_19116;
assign v_19120 = v_19118 | v_19119;
assign v_19123 = v_19121 | v_19122;
assign v_19126 = v_19124 | v_19125;
assign v_19129 = v_19127 | v_19128;
assign v_19132 = v_19130 | v_19131;
assign v_19135 = v_19133 | v_19134;
assign v_19138 = v_19136 | v_19137;
assign v_19141 = v_19139 | v_19140;
assign v_19144 = v_19142 | v_19143;
assign v_19147 = v_19145 | v_19146;
assign v_19150 = v_19148 | v_19149;
assign v_19153 = v_19151 | v_19152;
assign v_19156 = v_19154 | v_19155;
assign v_19159 = v_19157 | v_19158;
assign v_19162 = v_19160 | v_19161;
assign v_19165 = v_19163 | v_19164;
assign v_19168 = v_19166 | v_19167;
assign v_19171 = v_19169 | v_19170;
assign v_19174 = v_19172 | v_19173;
assign v_19177 = v_19175 | v_19176;
assign v_19178 = v_18991 | v_19177;
assign v_19179 = v_9336 | ~v_9844;
assign v_19180 = v_9308 | ~v_9712;
assign v_19182 = v_9051 | v_19181;
assign v_19183 = v_9026 | ~v_9554;
assign v_19185 = v_9052 | v_19184;
assign v_19186 = v_9027 | ~v_9422;
assign v_19188 = v_8761 | v_19187;
assign v_19189 = v_8729 | ~v_9266;
assign v_19191 = v_8762 | v_19190;
assign v_19192 = v_8730 | ~v_9134;
assign v_19194 = v_8473 | v_19193;
assign v_19195 = v_8447 | ~v_8984;
assign v_19197 = v_8474 | v_19196;
assign v_19198 = v_8448 | ~v_8852;
assign v_19200 = v_8185 | v_19199;
assign v_19201 = v_8157 | ~v_8688;
assign v_19203 = v_8186 | v_19202;
assign v_19204 = v_8158 | ~v_8556;
assign v_19206 = v_7901 | v_19205;
assign v_19207 = v_7876 | ~v_8404;
assign v_19209 = v_7902 | v_19208;
assign v_19210 = v_7877 | ~v_8272;
assign v_19212 = v_7607 | v_19211;
assign v_19213 = v_7571 | ~v_8116;
assign v_19215 = v_7608 | v_19214;
assign v_19216 = v_7572 | ~v_7984;
assign v_19218 = v_7315 | v_19217;
assign v_19219 = v_7288 | ~v_7834;
assign v_19221 = v_7316 | v_19220;
assign v_19222 = v_7289 | ~v_7702;
assign v_19224 = v_7025 | v_19223;
assign v_19225 = v_6997 | ~v_7530;
assign v_19227 = v_7026 | v_19226;
assign v_19228 = v_6998 | ~v_7398;
assign v_19230 = v_6741 | v_19229;
assign v_19231 = v_6716 | ~v_7244;
assign v_19233 = v_6742 | v_19232;
assign v_19234 = v_6717 | ~v_7112;
assign v_19236 = v_6451 | v_19235;
assign v_19237 = v_6419 | ~v_6956;
assign v_19239 = v_6452 | v_19238;
assign v_19240 = v_6420 | v_6824;
assign v_19242 = v_6163 | v_19241;
assign v_19243 = v_6137 | ~v_6674;
assign v_19245 = v_6164 | v_19244;
assign v_19246 = v_6138 | ~v_6542;
assign v_19248 = v_5875 | v_19247;
assign v_19249 = v_5847 | ~v_6378;
assign v_19251 = v_5876 | v_19250;
assign v_19252 = v_5848 | ~v_6246;
assign v_19254 = v_5591 | v_19253;
assign v_19255 = v_5566 | v_6094;
assign v_19257 = v_5592 | v_19256;
assign v_19258 = v_5567 | ~v_5962;
assign v_19260 = v_5293 | v_19259;
assign v_19261 = v_5253 | v_5806;
assign v_19263 = v_5294 | v_19262;
assign v_19264 = v_5254 | ~v_5674;
assign v_19266 = v_4997 | v_19265;
assign v_19267 = v_4969 | ~v_5524;
assign v_19269 = v_4998 | v_19268;
assign v_19270 = v_4970 | ~v_5392;
assign v_19272 = v_4705 | v_19271;
assign v_19273 = v_4677 | ~v_5212;
assign v_19275 = v_4706 | v_19274;
assign v_19276 = v_4678 | ~v_5080;
assign v_19278 = v_4421 | v_19277;
assign v_19279 = v_4396 | ~v_4924;
assign v_19281 = v_4422 | v_19280;
assign v_19282 = v_4397 | ~v_4792;
assign v_19284 = v_4131 | v_19283;
assign v_19285 = v_4099 | ~v_4636;
assign v_19287 = v_4132 | v_19286;
assign v_19288 = v_4100 | ~v_4504;
assign v_19290 = v_3843 | v_19289;
assign v_19291 = v_3817 | ~v_4354;
assign v_19293 = v_3844 | v_19292;
assign v_19294 = v_3818 | ~v_4222;
assign v_19296 = v_3555 | v_19295;
assign v_19297 = v_3527 | ~v_4058;
assign v_19299 = v_3556 | v_19298;
assign v_19300 = v_3528 | ~v_3926;
assign v_19302 = v_3271 | v_19301;
assign v_19303 = v_3246 | ~v_3774;
assign v_19305 = v_3272 | v_19304;
assign v_19306 = v_3247 | ~v_3642;
assign v_19308 = v_2977 | v_19307;
assign v_19309 = v_2941 | ~v_3486;
assign v_19311 = v_2978 | v_19310;
assign v_19312 = v_2942 | ~v_3354;
assign v_19314 = v_2685 | v_19313;
assign v_19315 = v_2658 | v_3204;
assign v_19317 = v_2686 | v_19316;
assign v_19318 = v_2659 | ~v_3072;
assign v_19320 = v_2395 | v_19319;
assign v_19321 = v_2367 | ~v_2900;
assign v_19323 = v_2396 | v_19322;
assign v_19324 = v_2368 | ~v_2768;
assign v_19326 = v_2111 | v_19325;
assign v_19327 = v_2086 | ~v_2614;
assign v_19329 = v_2112 | v_19328;
assign v_19330 = v_2087 | ~v_2482;
assign v_19332 = v_1821 | v_19331;
assign v_19333 = v_1789 | ~v_2326;
assign v_19335 = v_1822 | v_19334;
assign v_19336 = v_1790 | ~v_2194;
assign v_19338 = v_1533 | v_19337;
assign v_19339 = v_1507 | ~v_2044;
assign v_19341 = v_1534 | v_19340;
assign v_19342 = v_1508 | ~v_1912;
assign v_19344 = v_1245 | v_19343;
assign v_19345 = v_1217 | ~v_1748;
assign v_19347 = v_1246 | v_19346;
assign v_19348 = v_1218 | ~v_1616;
assign v_19350 = v_961 | v_19349;
assign v_19351 = v_936 | ~v_1464;
assign v_19353 = v_962 | v_19352;
assign v_19354 = v_937 | ~v_1332;
assign v_19356 = v_591 | v_19355;
assign v_19357 = v_92 | ~v_1176;
assign v_19359 = v_593 | v_19358;
assign v_19360 = v_94 | ~v_1044;
assign v_19362 = v_823 | v_19361;
assign v_19363 = v_806 | ~v_898;
assign v_19365 = v_19178 | v_19364;
assign v_19368 = v_19366 | v_19367;
assign v_19371 = v_19369 | v_19370;
assign v_19374 = v_19372 | v_19373;
assign v_19377 = v_19375 | v_19376;
assign v_19380 = v_19378 | v_19379;
assign v_19383 = v_19381 | v_19382;
assign v_19386 = v_19384 | v_19385;
assign v_19389 = v_19387 | v_19388;
assign v_19392 = v_19390 | v_19391;
assign v_19395 = v_19393 | v_19394;
assign v_19398 = v_19396 | v_19397;
assign v_19401 = v_19399 | v_19400;
assign v_19404 = v_19402 | v_19403;
assign v_19407 = v_19405 | v_19406;
assign v_19410 = v_19408 | v_19409;
assign v_19413 = v_19411 | v_19412;
assign v_19416 = v_19414 | v_19415;
assign v_19419 = v_19417 | v_19418;
assign v_19422 = v_19420 | v_19421;
assign v_19425 = v_19423 | v_19424;
assign v_19428 = v_19426 | v_19427;
assign v_19431 = v_19429 | v_19430;
assign v_19434 = v_19432 | v_19433;
assign v_19437 = v_19435 | v_19436;
assign v_19440 = v_19438 | v_19439;
assign v_19443 = v_19441 | v_19442;
assign v_19446 = v_19444 | v_19445;
assign v_19449 = v_19447 | v_19448;
assign v_19452 = v_19450 | v_19451;
assign v_19455 = v_19453 | v_19454;
assign v_19458 = v_19456 | v_19457;
assign v_19461 = v_19459 | v_19460;
assign v_19464 = v_19462 | v_19463;
assign v_19467 = v_19465 | v_19466;
assign v_19470 = v_19468 | v_19469;
assign v_19473 = v_19471 | v_19472;
assign v_19476 = v_19474 | v_19475;
assign v_19479 = v_19477 | v_19478;
assign v_19482 = v_19480 | v_19481;
assign v_19485 = v_19483 | v_19484;
assign v_19488 = v_19486 | v_19487;
assign v_19491 = v_19489 | v_19490;
assign v_19494 = v_19492 | v_19493;
assign v_19497 = v_19495 | v_19496;
assign v_19500 = v_19498 | v_19499;
assign v_19503 = v_19501 | v_19502;
assign v_19506 = v_19504 | v_19505;
assign v_19509 = v_19507 | v_19508;
assign v_19512 = v_19510 | v_19511;
assign v_19515 = v_19513 | v_19514;
assign v_19518 = v_19516 | v_19517;
assign v_19521 = v_19519 | v_19520;
assign v_19524 = v_19522 | v_19523;
assign v_19527 = v_19525 | v_19526;
assign v_19530 = v_19528 | v_19529;
assign v_19533 = v_19531 | v_19532;
assign v_19536 = v_19534 | v_19535;
assign v_19539 = v_19537 | v_19538;
assign v_19542 = v_19540 | v_19541;
assign v_19545 = v_19543 | v_19544;
assign v_19548 = v_19546 | v_19547;
assign v_19551 = v_19549 | v_19550;
assign v_19552 = v_19365 | v_19551;
assign v_19553 = v_13540 | v_19552;
assign v_19554 = v_18057 | v_19553;
assign v_19555 = v_10462 | v_19554;
assign v_19559 = v_19557 | v_19558;
assign v_19562 = v_19560 | v_19561;
assign v_19565 = v_19563 | v_19564;
assign v_19568 = v_19566 | v_19567;
assign v_19571 = v_19569 | v_19570;
assign v_19574 = v_19572 | v_19573;
assign v_19577 = v_19575 | v_19576;
assign v_19580 = v_19578 | v_19579;
assign v_19583 = v_19581 | v_19582;
assign v_19586 = v_19584 | v_19585;
assign v_19589 = v_19587 | v_19588;
assign v_19592 = v_19590 | v_19591;
assign v_19595 = v_19593 | v_19594;
assign v_19598 = v_19596 | v_19597;
assign v_19601 = v_19599 | v_19600;
assign v_19604 = v_19602 | v_19603;
assign v_19607 = v_19605 | v_19606;
assign v_19610 = v_19608 | v_19609;
assign v_19613 = v_19611 | v_19612;
assign v_19616 = v_19614 | v_19615;
assign v_19619 = v_19617 | v_19618;
assign v_19622 = v_19620 | v_19621;
assign v_19625 = v_19623 | v_19624;
assign v_19628 = v_19626 | v_19627;
assign v_19631 = v_19629 | v_19630;
assign v_19634 = v_19632 | v_19633;
assign v_19637 = v_19635 | v_19636;
assign v_19640 = v_19638 | v_19639;
assign v_19643 = v_19641 | v_19642;
assign v_19646 = v_19644 | v_19645;
assign v_19649 = v_19647 | v_19648;
assign v_19652 = v_19650 | v_19651;
assign v_19655 = v_19653 | v_19654;
assign v_19658 = v_19656 | v_19657;
assign v_19661 = v_19659 | v_19660;
assign v_19664 = v_19662 | v_19663;
assign v_19667 = v_19665 | v_19666;
assign v_19670 = v_19668 | v_19669;
assign v_19673 = v_19671 | v_19672;
assign v_19676 = v_19674 | v_19675;
assign v_19679 = v_19677 | v_19678;
assign v_19682 = v_19680 | v_19681;
assign v_19685 = v_19683 | v_19684;
assign v_19688 = v_19686 | v_19687;
assign v_19691 = v_19689 | v_19690;
assign v_19694 = v_19692 | v_19693;
assign v_19697 = v_19695 | v_19696;
assign v_19700 = v_19698 | v_19699;
assign v_19703 = v_19701 | v_19702;
assign v_19706 = v_19704 | v_19705;
assign v_19709 = v_19707 | v_19708;
assign v_19712 = v_19710 | v_19711;
assign v_19715 = v_19713 | v_19714;
assign v_19718 = v_19716 | v_19717;
assign v_19721 = v_19719 | v_19720;
assign v_19724 = v_19722 | v_19723;
assign v_19727 = v_19725 | v_19726;
assign v_19730 = v_19728 | v_19729;
assign v_19733 = v_19731 | v_19732;
assign v_19736 = v_19734 | v_19735;
assign v_19739 = v_19737 | v_19738;
assign v_19742 = v_19740 | v_19741;
assign v_19745 = v_19743 | v_19744;
assign v_19748 = v_19746 | v_19747;
assign v_19751 = v_19749 | v_19750;
assign v_19754 = v_19752 | v_19753;
assign v_19757 = v_19755 | v_19756;
assign v_19760 = v_19758 | v_19759;
assign v_19763 = v_19761 | v_19762;
assign v_19766 = v_19764 | v_19765;
assign v_19769 = v_19767 | v_19768;
assign v_19772 = v_19770 | v_19771;
assign v_19775 = v_19773 | v_19774;
assign v_19778 = v_19776 | v_19777;
assign v_19781 = v_19779 | v_19780;
assign v_19784 = v_19782 | v_19783;
assign v_19787 = v_19785 | v_19786;
assign v_19790 = v_19788 | v_19789;
assign v_19793 = v_19791 | v_19792;
assign v_19796 = v_19794 | v_19795;
assign v_19799 = v_19797 | v_19798;
assign v_19802 = v_19800 | v_19801;
assign v_19805 = v_19803 | v_19804;
assign v_19808 = v_19806 | v_19807;
assign v_19811 = v_19809 | v_19810;
assign v_19814 = v_19812 | v_19813;
assign v_19817 = v_19815 | v_19816;
assign v_19820 = v_19818 | v_19819;
assign v_19823 = v_19821 | v_19822;
assign v_19826 = v_19824 | v_19825;
assign v_19829 = v_19827 | v_19828;
assign v_19832 = v_19830 | v_19831;
assign v_19835 = v_19833 | v_19834;
assign v_19838 = v_19836 | v_19837;
assign v_19841 = v_19839 | v_19840;
assign v_19844 = v_19842 | v_19843;
assign v_19847 = v_19845 | v_19846;
assign v_19850 = v_19848 | v_19849;
assign v_19853 = v_19851 | v_19852;
assign v_19856 = v_19854 | v_19855;
assign v_19859 = v_19857 | v_19858;
assign v_19862 = v_19860 | v_19861;
assign v_19865 = v_19863 | v_19864;
assign v_19868 = v_19866 | v_19867;
assign v_19871 = v_19869 | v_19870;
assign v_19874 = v_19872 | v_19873;
assign v_19877 = v_19875 | v_19876;
assign v_19880 = v_19878 | v_19879;
assign v_19883 = v_19881 | v_19882;
assign v_19886 = v_19884 | v_19885;
assign v_19889 = v_19887 | v_19888;
assign v_19892 = v_19890 | v_19891;
assign v_19895 = v_19893 | v_19894;
assign v_19898 = v_19896 | v_19897;
assign v_19901 = v_19899 | v_19900;
assign v_19904 = v_19902 | v_19903;
assign v_19907 = v_19905 | v_19906;
assign v_19910 = v_19908 | v_19909;
assign v_19913 = v_19911 | v_19912;
assign v_19916 = v_19914 | v_19915;
assign v_19919 = v_19917 | v_19918;
assign v_19922 = v_19920 | v_19921;
assign v_19925 = v_19923 | v_19924;
assign v_19928 = v_19926 | v_19927;
assign v_19931 = v_19929 | v_19930;
assign v_19934 = v_19932 | v_19933;
assign v_19935 = v_19745 | v_19934;
assign v_19938 = v_19936 | v_19937;
assign v_19941 = v_19939 | v_19940;
assign v_19944 = v_19942 | v_19943;
assign v_19947 = v_19945 | v_19946;
assign v_19950 = v_19948 | v_19949;
assign v_19953 = v_19951 | v_19952;
assign v_19956 = v_19954 | v_19955;
assign v_19959 = v_19957 | v_19958;
assign v_19962 = v_19960 | v_19961;
assign v_19965 = v_19963 | v_19964;
assign v_19968 = v_19966 | v_19967;
assign v_19971 = v_19969 | v_19970;
assign v_19974 = v_19972 | v_19973;
assign v_19977 = v_19975 | v_19976;
assign v_19980 = v_19978 | v_19979;
assign v_19983 = v_19981 | v_19982;
assign v_19986 = v_19984 | v_19985;
assign v_19989 = v_19987 | v_19988;
assign v_19992 = v_19990 | v_19991;
assign v_19995 = v_19993 | v_19994;
assign v_19998 = v_19996 | v_19997;
assign v_20001 = v_19999 | v_20000;
assign v_20004 = v_20002 | v_20003;
assign v_20007 = v_20005 | v_20006;
assign v_20010 = v_20008 | v_20009;
assign v_20013 = v_20011 | v_20012;
assign v_20016 = v_20014 | v_20015;
assign v_20019 = v_20017 | v_20018;
assign v_20022 = v_20020 | v_20021;
assign v_20025 = v_20023 | v_20024;
assign v_20028 = v_20026 | v_20027;
assign v_20031 = v_20029 | v_20030;
assign v_20034 = v_20032 | v_20033;
assign v_20037 = v_20035 | v_20036;
assign v_20040 = v_20038 | v_20039;
assign v_20043 = v_20041 | v_20042;
assign v_20046 = v_20044 | v_20045;
assign v_20049 = v_20047 | v_20048;
assign v_20052 = v_20050 | v_20051;
assign v_20055 = v_20053 | v_20054;
assign v_20058 = v_20056 | v_20057;
assign v_20061 = v_20059 | v_20060;
assign v_20064 = v_20062 | v_20063;
assign v_20067 = v_20065 | v_20066;
assign v_20070 = v_20068 | v_20069;
assign v_20073 = v_20071 | v_20072;
assign v_20076 = v_20074 | v_20075;
assign v_20079 = v_20077 | v_20078;
assign v_20082 = v_20080 | v_20081;
assign v_20085 = v_20083 | v_20084;
assign v_20088 = v_20086 | v_20087;
assign v_20091 = v_20089 | v_20090;
assign v_20094 = v_20092 | v_20093;
assign v_20097 = v_20095 | v_20096;
assign v_20100 = v_20098 | v_20099;
assign v_20103 = v_20101 | v_20102;
assign v_20106 = v_20104 | v_20105;
assign v_20109 = v_20107 | v_20108;
assign v_20112 = v_20110 | v_20111;
assign v_20115 = v_20113 | v_20114;
assign v_20118 = v_20116 | v_20117;
assign v_20121 = v_20119 | v_20120;
assign v_20124 = v_20122 | v_20123;
assign v_20125 = v_19935 | v_20124;
assign v_20128 = v_20126 | v_20127;
assign v_20131 = v_20129 | v_20130;
assign v_20134 = v_20132 | v_20133;
assign v_20137 = v_20135 | v_20136;
assign v_20140 = v_20138 | v_20139;
assign v_20143 = v_20141 | v_20142;
assign v_20146 = v_20144 | v_20145;
assign v_20149 = v_20147 | v_20148;
assign v_20152 = v_20150 | v_20151;
assign v_20155 = v_20153 | v_20154;
assign v_20158 = v_20156 | v_20157;
assign v_20161 = v_20159 | v_20160;
assign v_20164 = v_20162 | v_20163;
assign v_20167 = v_20165 | v_20166;
assign v_20170 = v_20168 | v_20169;
assign v_20173 = v_20171 | v_20172;
assign v_20176 = v_20174 | v_20175;
assign v_20179 = v_20177 | v_20178;
assign v_20182 = v_20180 | v_20181;
assign v_20185 = v_20183 | v_20184;
assign v_20188 = v_20186 | v_20187;
assign v_20191 = v_20189 | v_20190;
assign v_20194 = v_20192 | v_20193;
assign v_20197 = v_20195 | v_20196;
assign v_20200 = v_20198 | v_20199;
assign v_20203 = v_20201 | v_20202;
assign v_20206 = v_20204 | v_20205;
assign v_20209 = v_20207 | v_20208;
assign v_20212 = v_20210 | v_20211;
assign v_20215 = v_20213 | v_20214;
assign v_20218 = v_20216 | v_20217;
assign v_20221 = v_20219 | v_20220;
assign v_20224 = v_20222 | v_20223;
assign v_20227 = v_20225 | v_20226;
assign v_20230 = v_20228 | v_20229;
assign v_20233 = v_20231 | v_20232;
assign v_20236 = v_20234 | v_20235;
assign v_20239 = v_20237 | v_20238;
assign v_20242 = v_20240 | v_20241;
assign v_20245 = v_20243 | v_20244;
assign v_20248 = v_20246 | v_20247;
assign v_20251 = v_20249 | v_20250;
assign v_20254 = v_20252 | v_20253;
assign v_20257 = v_20255 | v_20256;
assign v_20260 = v_20258 | v_20259;
assign v_20263 = v_20261 | v_20262;
assign v_20266 = v_20264 | v_20265;
assign v_20269 = v_20267 | v_20268;
assign v_20272 = v_20270 | v_20271;
assign v_20275 = v_20273 | v_20274;
assign v_20278 = v_20276 | v_20277;
assign v_20281 = v_20279 | v_20280;
assign v_20284 = v_20282 | v_20283;
assign v_20287 = v_20285 | v_20286;
assign v_20290 = v_20288 | v_20289;
assign v_20293 = v_20291 | v_20292;
assign v_20296 = v_20294 | v_20295;
assign v_20299 = v_20297 | v_20298;
assign v_20302 = v_20300 | v_20301;
assign v_20305 = v_20303 | v_20304;
assign v_20308 = v_20306 | v_20307;
assign v_20311 = v_20309 | v_20310;
assign v_20314 = v_20312 | v_20313;
assign v_20315 = v_20125 | v_20314;
assign v_20318 = v_20316 | v_20317;
assign v_20321 = v_20319 | v_20320;
assign v_20324 = v_20322 | v_20323;
assign v_20327 = v_20325 | v_20326;
assign v_20330 = v_20328 | v_20329;
assign v_20333 = v_20331 | v_20332;
assign v_20336 = v_20334 | v_20335;
assign v_20339 = v_20337 | v_20338;
assign v_20342 = v_20340 | v_20341;
assign v_20345 = v_20343 | v_20344;
assign v_20348 = v_20346 | v_20347;
assign v_20351 = v_20349 | v_20350;
assign v_20354 = v_20352 | v_20353;
assign v_20357 = v_20355 | v_20356;
assign v_20360 = v_20358 | v_20359;
assign v_20363 = v_20361 | v_20362;
assign v_20366 = v_20364 | v_20365;
assign v_20369 = v_20367 | v_20368;
assign v_20372 = v_20370 | v_20371;
assign v_20375 = v_20373 | v_20374;
assign v_20378 = v_20376 | v_20377;
assign v_20381 = v_20379 | v_20380;
assign v_20384 = v_20382 | v_20383;
assign v_20387 = v_20385 | v_20386;
assign v_20390 = v_20388 | v_20389;
assign v_20393 = v_20391 | v_20392;
assign v_20396 = v_20394 | v_20395;
assign v_20399 = v_20397 | v_20398;
assign v_20402 = v_20400 | v_20401;
assign v_20405 = v_20403 | v_20404;
assign v_20408 = v_20406 | v_20407;
assign v_20411 = v_20409 | v_20410;
assign v_20414 = v_20412 | v_20413;
assign v_20417 = v_20415 | v_20416;
assign v_20420 = v_20418 | v_20419;
assign v_20423 = v_20421 | v_20422;
assign v_20426 = v_20424 | v_20425;
assign v_20429 = v_20427 | v_20428;
assign v_20432 = v_20430 | v_20431;
assign v_20435 = v_20433 | v_20434;
assign v_20438 = v_20436 | v_20437;
assign v_20441 = v_20439 | v_20440;
assign v_20444 = v_20442 | v_20443;
assign v_20447 = v_20445 | v_20446;
assign v_20450 = v_20448 | v_20449;
assign v_20453 = v_20451 | v_20452;
assign v_20456 = v_20454 | v_20455;
assign v_20459 = v_20457 | v_20458;
assign v_20462 = v_20460 | v_20461;
assign v_20465 = v_20463 | v_20464;
assign v_20468 = v_20466 | v_20467;
assign v_20471 = v_20469 | v_20470;
assign v_20474 = v_20472 | v_20473;
assign v_20477 = v_20475 | v_20476;
assign v_20480 = v_20478 | v_20479;
assign v_20483 = v_20481 | v_20482;
assign v_20486 = v_20484 | v_20485;
assign v_20489 = v_20487 | v_20488;
assign v_20492 = v_20490 | v_20491;
assign v_20495 = v_20493 | v_20494;
assign v_20498 = v_20496 | v_20497;
assign v_20501 = v_20499 | v_20500;
assign v_20504 = v_20502 | v_20503;
assign v_20505 = v_20315 | v_20504;
assign v_20508 = v_20506 | v_20507;
assign v_20511 = v_20509 | v_20510;
assign v_20514 = v_20512 | v_20513;
assign v_20517 = v_20515 | v_20516;
assign v_20520 = v_20518 | v_20519;
assign v_20523 = v_20521 | v_20522;
assign v_20526 = v_20524 | v_20525;
assign v_20529 = v_20527 | v_20528;
assign v_20532 = v_20530 | v_20531;
assign v_20535 = v_20533 | v_20534;
assign v_20538 = v_20536 | v_20537;
assign v_20541 = v_20539 | v_20540;
assign v_20544 = v_20542 | v_20543;
assign v_20547 = v_20545 | v_20546;
assign v_20550 = v_20548 | v_20549;
assign v_20553 = v_20551 | v_20552;
assign v_20556 = v_20554 | v_20555;
assign v_20559 = v_20557 | v_20558;
assign v_20562 = v_20560 | v_20561;
assign v_20565 = v_20563 | v_20564;
assign v_20568 = v_20566 | v_20567;
assign v_20571 = v_20569 | v_20570;
assign v_20574 = v_20572 | v_20573;
assign v_20577 = v_20575 | v_20576;
assign v_20580 = v_20578 | v_20579;
assign v_20583 = v_20581 | v_20582;
assign v_20586 = v_20584 | v_20585;
assign v_20589 = v_20587 | v_20588;
assign v_20592 = v_20590 | v_20591;
assign v_20595 = v_20593 | v_20594;
assign v_20598 = v_20596 | v_20597;
assign v_20601 = v_20599 | v_20600;
assign v_20604 = v_20602 | v_20603;
assign v_20607 = v_20605 | v_20606;
assign v_20610 = v_20608 | v_20609;
assign v_20613 = v_20611 | v_20612;
assign v_20616 = v_20614 | v_20615;
assign v_20619 = v_20617 | v_20618;
assign v_20622 = v_20620 | v_20621;
assign v_20625 = v_20623 | v_20624;
assign v_20628 = v_20626 | v_20627;
assign v_20631 = v_20629 | v_20630;
assign v_20634 = v_20632 | v_20633;
assign v_20637 = v_20635 | v_20636;
assign v_20640 = v_20638 | v_20639;
assign v_20643 = v_20641 | v_20642;
assign v_20646 = v_20644 | v_20645;
assign v_20649 = v_20647 | v_20648;
assign v_20652 = v_20650 | v_20651;
assign v_20655 = v_20653 | v_20654;
assign v_20658 = v_20656 | v_20657;
assign v_20661 = v_20659 | v_20660;
assign v_20664 = v_20662 | v_20663;
assign v_20667 = v_20665 | v_20666;
assign v_20670 = v_20668 | v_20669;
assign v_20673 = v_20671 | v_20672;
assign v_20676 = v_20674 | v_20675;
assign v_20679 = v_20677 | v_20678;
assign v_20682 = v_20680 | v_20681;
assign v_20685 = v_20683 | v_20684;
assign v_20688 = v_20686 | v_20687;
assign v_20691 = v_20689 | v_20690;
assign v_20694 = v_20692 | v_20693;
assign v_20695 = v_20505 | v_20694;
assign v_20698 = v_20696 | v_20697;
assign v_20701 = v_20699 | v_20700;
assign v_20704 = v_20702 | v_20703;
assign v_20707 = v_20705 | v_20706;
assign v_20710 = v_20708 | v_20709;
assign v_20713 = v_20711 | v_20712;
assign v_20716 = v_20714 | v_20715;
assign v_20719 = v_20717 | v_20718;
assign v_20722 = v_20720 | v_20721;
assign v_20725 = v_20723 | v_20724;
assign v_20728 = v_20726 | v_20727;
assign v_20731 = v_20729 | v_20730;
assign v_20734 = v_20732 | v_20733;
assign v_20737 = v_20735 | v_20736;
assign v_20740 = v_20738 | v_20739;
assign v_20743 = v_20741 | v_20742;
assign v_20746 = v_20744 | v_20745;
assign v_20749 = v_20747 | v_20748;
assign v_20752 = v_20750 | v_20751;
assign v_20755 = v_20753 | v_20754;
assign v_20758 = v_20756 | v_20757;
assign v_20761 = v_20759 | v_20760;
assign v_20764 = v_20762 | v_20763;
assign v_20767 = v_20765 | v_20766;
assign v_20770 = v_20768 | v_20769;
assign v_20773 = v_20771 | v_20772;
assign v_20776 = v_20774 | v_20775;
assign v_20779 = v_20777 | v_20778;
assign v_20782 = v_20780 | v_20781;
assign v_20785 = v_20783 | v_20784;
assign v_20788 = v_20786 | v_20787;
assign v_20791 = v_20789 | v_20790;
assign v_20794 = v_20792 | v_20793;
assign v_20797 = v_20795 | v_20796;
assign v_20800 = v_20798 | v_20799;
assign v_20803 = v_20801 | v_20802;
assign v_20806 = v_20804 | v_20805;
assign v_20809 = v_20807 | v_20808;
assign v_20812 = v_20810 | v_20811;
assign v_20815 = v_20813 | v_20814;
assign v_20818 = v_20816 | v_20817;
assign v_20821 = v_20819 | v_20820;
assign v_20824 = v_20822 | v_20823;
assign v_20827 = v_20825 | v_20826;
assign v_20830 = v_20828 | v_20829;
assign v_20833 = v_20831 | v_20832;
assign v_20836 = v_20834 | v_20835;
assign v_20839 = v_20837 | v_20838;
assign v_20842 = v_20840 | v_20841;
assign v_20845 = v_20843 | v_20844;
assign v_20848 = v_20846 | v_20847;
assign v_20851 = v_20849 | v_20850;
assign v_20854 = v_20852 | v_20853;
assign v_20857 = v_20855 | v_20856;
assign v_20860 = v_20858 | v_20859;
assign v_20863 = v_20861 | v_20862;
assign v_20866 = v_20864 | v_20865;
assign v_20869 = v_20867 | v_20868;
assign v_20872 = v_20870 | v_20871;
assign v_20875 = v_20873 | v_20874;
assign v_20878 = v_20876 | v_20877;
assign v_20881 = v_20879 | v_20880;
assign v_20884 = v_20882 | v_20883;
assign v_20885 = v_20695 | v_20884;
assign v_20888 = v_20886 | v_20887;
assign v_20891 = v_20889 | v_20890;
assign v_20894 = v_20892 | v_20893;
assign v_20897 = v_20895 | v_20896;
assign v_20900 = v_20898 | v_20899;
assign v_20903 = v_20901 | v_20902;
assign v_20906 = v_20904 | v_20905;
assign v_20909 = v_20907 | v_20908;
assign v_20912 = v_20910 | v_20911;
assign v_20915 = v_20913 | v_20914;
assign v_20918 = v_20916 | v_20917;
assign v_20921 = v_20919 | v_20920;
assign v_20924 = v_20922 | v_20923;
assign v_20927 = v_20925 | v_20926;
assign v_20930 = v_20928 | v_20929;
assign v_20933 = v_20931 | v_20932;
assign v_20936 = v_20934 | v_20935;
assign v_20939 = v_20937 | v_20938;
assign v_20942 = v_20940 | v_20941;
assign v_20945 = v_20943 | v_20944;
assign v_20948 = v_20946 | v_20947;
assign v_20951 = v_20949 | v_20950;
assign v_20954 = v_20952 | v_20953;
assign v_20957 = v_20955 | v_20956;
assign v_20960 = v_20958 | v_20959;
assign v_20963 = v_20961 | v_20962;
assign v_20966 = v_20964 | v_20965;
assign v_20969 = v_20967 | v_20968;
assign v_20972 = v_20970 | v_20971;
assign v_20975 = v_20973 | v_20974;
assign v_20978 = v_20976 | v_20977;
assign v_20981 = v_20979 | v_20980;
assign v_20984 = v_20982 | v_20983;
assign v_20987 = v_20985 | v_20986;
assign v_20990 = v_20988 | v_20989;
assign v_20993 = v_20991 | v_20992;
assign v_20996 = v_20994 | v_20995;
assign v_20999 = v_20997 | v_20998;
assign v_21002 = v_21000 | v_21001;
assign v_21005 = v_21003 | v_21004;
assign v_21008 = v_21006 | v_21007;
assign v_21011 = v_21009 | v_21010;
assign v_21014 = v_21012 | v_21013;
assign v_21017 = v_21015 | v_21016;
assign v_21020 = v_21018 | v_21019;
assign v_21023 = v_21021 | v_21022;
assign v_21026 = v_21024 | v_21025;
assign v_21029 = v_21027 | v_21028;
assign v_21032 = v_21030 | v_21031;
assign v_21035 = v_21033 | v_21034;
assign v_21038 = v_21036 | v_21037;
assign v_21041 = v_21039 | v_21040;
assign v_21044 = v_21042 | v_21043;
assign v_21047 = v_21045 | v_21046;
assign v_21050 = v_21048 | v_21049;
assign v_21053 = v_21051 | v_21052;
assign v_21056 = v_21054 | v_21055;
assign v_21059 = v_21057 | v_21058;
assign v_21062 = v_21060 | v_21061;
assign v_21065 = v_21063 | v_21064;
assign v_21068 = v_21066 | v_21067;
assign v_21071 = v_21069 | v_21070;
assign v_21074 = v_21072 | v_21073;
assign v_21075 = v_20885 | v_21074;
assign v_21078 = v_21076 | v_21077;
assign v_21081 = v_21079 | v_21080;
assign v_21084 = v_21082 | v_21083;
assign v_21087 = v_21085 | v_21086;
assign v_21090 = v_21088 | v_21089;
assign v_21093 = v_21091 | v_21092;
assign v_21096 = v_21094 | v_21095;
assign v_21099 = v_21097 | v_21098;
assign v_21102 = v_21100 | v_21101;
assign v_21105 = v_21103 | v_21104;
assign v_21108 = v_21106 | v_21107;
assign v_21111 = v_21109 | v_21110;
assign v_21114 = v_21112 | v_21113;
assign v_21117 = v_21115 | v_21116;
assign v_21120 = v_21118 | v_21119;
assign v_21123 = v_21121 | v_21122;
assign v_21126 = v_21124 | v_21125;
assign v_21129 = v_21127 | v_21128;
assign v_21132 = v_21130 | v_21131;
assign v_21135 = v_21133 | v_21134;
assign v_21138 = v_21136 | v_21137;
assign v_21141 = v_21139 | v_21140;
assign v_21144 = v_21142 | v_21143;
assign v_21147 = v_21145 | v_21146;
assign v_21150 = v_21148 | v_21149;
assign v_21153 = v_21151 | v_21152;
assign v_21156 = v_21154 | v_21155;
assign v_21159 = v_21157 | v_21158;
assign v_21162 = v_21160 | v_21161;
assign v_21165 = v_21163 | v_21164;
assign v_21168 = v_21166 | v_21167;
assign v_21171 = v_21169 | v_21170;
assign v_21174 = v_21172 | v_21173;
assign v_21177 = v_21175 | v_21176;
assign v_21180 = v_21178 | v_21179;
assign v_21183 = v_21181 | v_21182;
assign v_21186 = v_21184 | v_21185;
assign v_21189 = v_21187 | v_21188;
assign v_21192 = v_21190 | v_21191;
assign v_21195 = v_21193 | v_21194;
assign v_21198 = v_21196 | v_21197;
assign v_21201 = v_21199 | v_21200;
assign v_21204 = v_21202 | v_21203;
assign v_21207 = v_21205 | v_21206;
assign v_21210 = v_21208 | v_21209;
assign v_21213 = v_21211 | v_21212;
assign v_21216 = v_21214 | v_21215;
assign v_21219 = v_21217 | v_21218;
assign v_21222 = v_21220 | v_21221;
assign v_21225 = v_21223 | v_21224;
assign v_21228 = v_21226 | v_21227;
assign v_21231 = v_21229 | v_21230;
assign v_21234 = v_21232 | v_21233;
assign v_21237 = v_21235 | v_21236;
assign v_21240 = v_21238 | v_21239;
assign v_21243 = v_21241 | v_21242;
assign v_21246 = v_21244 | v_21245;
assign v_21249 = v_21247 | v_21248;
assign v_21252 = v_21250 | v_21251;
assign v_21255 = v_21253 | v_21254;
assign v_21258 = v_21256 | v_21257;
assign v_21261 = v_21259 | v_21260;
assign v_21264 = v_21262 | v_21263;
assign v_21267 = v_21265 | v_21266;
assign v_21270 = v_21268 | v_21269;
assign v_21273 = v_21271 | v_21272;
assign v_21276 = v_21274 | v_21275;
assign v_21279 = v_21277 | v_21278;
assign v_21282 = v_21280 | v_21281;
assign v_21285 = v_21283 | v_21284;
assign v_21288 = v_21286 | v_21287;
assign v_21291 = v_21289 | v_21290;
assign v_21294 = v_21292 | v_21293;
assign v_21297 = v_21295 | v_21296;
assign v_21300 = v_21298 | v_21299;
assign v_21303 = v_21301 | v_21302;
assign v_21306 = v_21304 | v_21305;
assign v_21309 = v_21307 | v_21308;
assign v_21312 = v_21310 | v_21311;
assign v_21315 = v_21313 | v_21314;
assign v_21318 = v_21316 | v_21317;
assign v_21321 = v_21319 | v_21320;
assign v_21324 = v_21322 | v_21323;
assign v_21327 = v_21325 | v_21326;
assign v_21330 = v_21328 | v_21329;
assign v_21333 = v_21331 | v_21332;
assign v_21336 = v_21334 | v_21335;
assign v_21339 = v_21337 | v_21338;
assign v_21342 = v_21340 | v_21341;
assign v_21345 = v_21343 | v_21344;
assign v_21348 = v_21346 | v_21347;
assign v_21351 = v_21349 | v_21350;
assign v_21354 = v_21352 | v_21353;
assign v_21357 = v_21355 | v_21356;
assign v_21360 = v_21358 | v_21359;
assign v_21363 = v_21361 | v_21362;
assign v_21366 = v_21364 | v_21365;
assign v_21369 = v_21367 | v_21368;
assign v_21372 = v_21370 | v_21371;
assign v_21375 = v_21373 | v_21374;
assign v_21378 = v_21376 | v_21377;
assign v_21381 = v_21379 | v_21380;
assign v_21384 = v_21382 | v_21383;
assign v_21387 = v_21385 | v_21386;
assign v_21390 = v_21388 | v_21389;
assign v_21393 = v_21391 | v_21392;
assign v_21396 = v_21394 | v_21395;
assign v_21399 = v_21397 | v_21398;
assign v_21402 = v_21400 | v_21401;
assign v_21405 = v_21403 | v_21404;
assign v_21408 = v_21406 | v_21407;
assign v_21411 = v_21409 | v_21410;
assign v_21414 = v_21412 | v_21413;
assign v_21417 = v_21415 | v_21416;
assign v_21420 = v_21418 | v_21419;
assign v_21423 = v_21421 | v_21422;
assign v_21426 = v_21424 | v_21425;
assign v_21429 = v_21427 | v_21428;
assign v_21432 = v_21430 | v_21431;
assign v_21435 = v_21433 | v_21434;
assign v_21438 = v_21436 | v_21437;
assign v_21441 = v_21439 | v_21440;
assign v_21444 = v_21442 | v_21443;
assign v_21447 = v_21445 | v_21446;
assign v_21450 = v_21448 | v_21449;
assign v_21453 = v_21451 | v_21452;
assign v_21454 = v_21264 | v_21453;
assign v_21457 = v_21455 | v_21456;
assign v_21460 = v_21458 | v_21459;
assign v_21463 = v_21461 | v_21462;
assign v_21466 = v_21464 | v_21465;
assign v_21469 = v_21467 | v_21468;
assign v_21472 = v_21470 | v_21471;
assign v_21475 = v_21473 | v_21474;
assign v_21478 = v_21476 | v_21477;
assign v_21481 = v_21479 | v_21480;
assign v_21484 = v_21482 | v_21483;
assign v_21487 = v_21485 | v_21486;
assign v_21490 = v_21488 | v_21489;
assign v_21493 = v_21491 | v_21492;
assign v_21496 = v_21494 | v_21495;
assign v_21499 = v_21497 | v_21498;
assign v_21502 = v_21500 | v_21501;
assign v_21505 = v_21503 | v_21504;
assign v_21508 = v_21506 | v_21507;
assign v_21511 = v_21509 | v_21510;
assign v_21514 = v_21512 | v_21513;
assign v_21517 = v_21515 | v_21516;
assign v_21520 = v_21518 | v_21519;
assign v_21523 = v_21521 | v_21522;
assign v_21526 = v_21524 | v_21525;
assign v_21529 = v_21527 | v_21528;
assign v_21532 = v_21530 | v_21531;
assign v_21535 = v_21533 | v_21534;
assign v_21538 = v_21536 | v_21537;
assign v_21541 = v_21539 | v_21540;
assign v_21544 = v_21542 | v_21543;
assign v_21547 = v_21545 | v_21546;
assign v_21550 = v_21548 | v_21549;
assign v_21553 = v_21551 | v_21552;
assign v_21556 = v_21554 | v_21555;
assign v_21559 = v_21557 | v_21558;
assign v_21562 = v_21560 | v_21561;
assign v_21565 = v_21563 | v_21564;
assign v_21568 = v_21566 | v_21567;
assign v_21571 = v_21569 | v_21570;
assign v_21574 = v_21572 | v_21573;
assign v_21577 = v_21575 | v_21576;
assign v_21580 = v_21578 | v_21579;
assign v_21583 = v_21581 | v_21582;
assign v_21586 = v_21584 | v_21585;
assign v_21589 = v_21587 | v_21588;
assign v_21592 = v_21590 | v_21591;
assign v_21595 = v_21593 | v_21594;
assign v_21598 = v_21596 | v_21597;
assign v_21601 = v_21599 | v_21600;
assign v_21604 = v_21602 | v_21603;
assign v_21607 = v_21605 | v_21606;
assign v_21610 = v_21608 | v_21609;
assign v_21613 = v_21611 | v_21612;
assign v_21616 = v_21614 | v_21615;
assign v_21619 = v_21617 | v_21618;
assign v_21622 = v_21620 | v_21621;
assign v_21625 = v_21623 | v_21624;
assign v_21628 = v_21626 | v_21627;
assign v_21631 = v_21629 | v_21630;
assign v_21634 = v_21632 | v_21633;
assign v_21637 = v_21635 | v_21636;
assign v_21640 = v_21638 | v_21639;
assign v_21643 = v_21641 | v_21642;
assign v_21644 = v_21454 | v_21643;
assign v_21647 = v_21645 | v_21646;
assign v_21650 = v_21648 | v_21649;
assign v_21653 = v_21651 | v_21652;
assign v_21656 = v_21654 | v_21655;
assign v_21659 = v_21657 | v_21658;
assign v_21662 = v_21660 | v_21661;
assign v_21665 = v_21663 | v_21664;
assign v_21668 = v_21666 | v_21667;
assign v_21671 = v_21669 | v_21670;
assign v_21674 = v_21672 | v_21673;
assign v_21677 = v_21675 | v_21676;
assign v_21680 = v_21678 | v_21679;
assign v_21683 = v_21681 | v_21682;
assign v_21686 = v_21684 | v_21685;
assign v_21689 = v_21687 | v_21688;
assign v_21692 = v_21690 | v_21691;
assign v_21695 = v_21693 | v_21694;
assign v_21698 = v_21696 | v_21697;
assign v_21701 = v_21699 | v_21700;
assign v_21704 = v_21702 | v_21703;
assign v_21707 = v_21705 | v_21706;
assign v_21710 = v_21708 | v_21709;
assign v_21713 = v_21711 | v_21712;
assign v_21716 = v_21714 | v_21715;
assign v_21719 = v_21717 | v_21718;
assign v_21722 = v_21720 | v_21721;
assign v_21725 = v_21723 | v_21724;
assign v_21728 = v_21726 | v_21727;
assign v_21731 = v_21729 | v_21730;
assign v_21734 = v_21732 | v_21733;
assign v_21737 = v_21735 | v_21736;
assign v_21740 = v_21738 | v_21739;
assign v_21743 = v_21741 | v_21742;
assign v_21746 = v_21744 | v_21745;
assign v_21749 = v_21747 | v_21748;
assign v_21752 = v_21750 | v_21751;
assign v_21755 = v_21753 | v_21754;
assign v_21758 = v_21756 | v_21757;
assign v_21761 = v_21759 | v_21760;
assign v_21764 = v_21762 | v_21763;
assign v_21767 = v_21765 | v_21766;
assign v_21770 = v_21768 | v_21769;
assign v_21773 = v_21771 | v_21772;
assign v_21776 = v_21774 | v_21775;
assign v_21779 = v_21777 | v_21778;
assign v_21782 = v_21780 | v_21781;
assign v_21785 = v_21783 | v_21784;
assign v_21788 = v_21786 | v_21787;
assign v_21791 = v_21789 | v_21790;
assign v_21794 = v_21792 | v_21793;
assign v_21797 = v_21795 | v_21796;
assign v_21800 = v_21798 | v_21799;
assign v_21803 = v_21801 | v_21802;
assign v_21806 = v_21804 | v_21805;
assign v_21809 = v_21807 | v_21808;
assign v_21812 = v_21810 | v_21811;
assign v_21815 = v_21813 | v_21814;
assign v_21818 = v_21816 | v_21817;
assign v_21821 = v_21819 | v_21820;
assign v_21824 = v_21822 | v_21823;
assign v_21827 = v_21825 | v_21826;
assign v_21830 = v_21828 | v_21829;
assign v_21833 = v_21831 | v_21832;
assign v_21834 = v_21644 | v_21833;
assign v_21837 = v_21835 | v_21836;
assign v_21840 = v_21838 | v_21839;
assign v_21843 = v_21841 | v_21842;
assign v_21846 = v_21844 | v_21845;
assign v_21849 = v_21847 | v_21848;
assign v_21852 = v_21850 | v_21851;
assign v_21855 = v_21853 | v_21854;
assign v_21858 = v_21856 | v_21857;
assign v_21861 = v_21859 | v_21860;
assign v_21864 = v_21862 | v_21863;
assign v_21867 = v_21865 | v_21866;
assign v_21870 = v_21868 | v_21869;
assign v_21873 = v_21871 | v_21872;
assign v_21876 = v_21874 | v_21875;
assign v_21879 = v_21877 | v_21878;
assign v_21882 = v_21880 | v_21881;
assign v_21885 = v_21883 | v_21884;
assign v_21888 = v_21886 | v_21887;
assign v_21891 = v_21889 | v_21890;
assign v_21894 = v_21892 | v_21893;
assign v_21897 = v_21895 | v_21896;
assign v_21900 = v_21898 | v_21899;
assign v_21903 = v_21901 | v_21902;
assign v_21906 = v_21904 | v_21905;
assign v_21909 = v_21907 | v_21908;
assign v_21912 = v_21910 | v_21911;
assign v_21915 = v_21913 | v_21914;
assign v_21918 = v_21916 | v_21917;
assign v_21921 = v_21919 | v_21920;
assign v_21924 = v_21922 | v_21923;
assign v_21927 = v_21925 | v_21926;
assign v_21930 = v_21928 | v_21929;
assign v_21933 = v_21931 | v_21932;
assign v_21936 = v_21934 | v_21935;
assign v_21939 = v_21937 | v_21938;
assign v_21942 = v_21940 | v_21941;
assign v_21945 = v_21943 | v_21944;
assign v_21948 = v_21946 | v_21947;
assign v_21951 = v_21949 | v_21950;
assign v_21954 = v_21952 | v_21953;
assign v_21957 = v_21955 | v_21956;
assign v_21960 = v_21958 | v_21959;
assign v_21963 = v_21961 | v_21962;
assign v_21966 = v_21964 | v_21965;
assign v_21969 = v_21967 | v_21968;
assign v_21972 = v_21970 | v_21971;
assign v_21975 = v_21973 | v_21974;
assign v_21978 = v_21976 | v_21977;
assign v_21981 = v_21979 | v_21980;
assign v_21984 = v_21982 | v_21983;
assign v_21987 = v_21985 | v_21986;
assign v_21990 = v_21988 | v_21989;
assign v_21993 = v_21991 | v_21992;
assign v_21996 = v_21994 | v_21995;
assign v_21999 = v_21997 | v_21998;
assign v_22002 = v_22000 | v_22001;
assign v_22005 = v_22003 | v_22004;
assign v_22008 = v_22006 | v_22007;
assign v_22011 = v_22009 | v_22010;
assign v_22014 = v_22012 | v_22013;
assign v_22017 = v_22015 | v_22016;
assign v_22020 = v_22018 | v_22019;
assign v_22023 = v_22021 | v_22022;
assign v_22024 = v_21834 | v_22023;
assign v_22027 = v_22025 | v_22026;
assign v_22030 = v_22028 | v_22029;
assign v_22033 = v_22031 | v_22032;
assign v_22036 = v_22034 | v_22035;
assign v_22039 = v_22037 | v_22038;
assign v_22042 = v_22040 | v_22041;
assign v_22045 = v_22043 | v_22044;
assign v_22048 = v_22046 | v_22047;
assign v_22051 = v_22049 | v_22050;
assign v_22054 = v_22052 | v_22053;
assign v_22057 = v_22055 | v_22056;
assign v_22060 = v_22058 | v_22059;
assign v_22063 = v_22061 | v_22062;
assign v_22066 = v_22064 | v_22065;
assign v_22069 = v_22067 | v_22068;
assign v_22072 = v_22070 | v_22071;
assign v_22075 = v_22073 | v_22074;
assign v_22078 = v_22076 | v_22077;
assign v_22081 = v_22079 | v_22080;
assign v_22084 = v_22082 | v_22083;
assign v_22087 = v_22085 | v_22086;
assign v_22090 = v_22088 | v_22089;
assign v_22093 = v_22091 | v_22092;
assign v_22096 = v_22094 | v_22095;
assign v_22099 = v_22097 | v_22098;
assign v_22102 = v_22100 | v_22101;
assign v_22105 = v_22103 | v_22104;
assign v_22108 = v_22106 | v_22107;
assign v_22111 = v_22109 | v_22110;
assign v_22114 = v_22112 | v_22113;
assign v_22117 = v_22115 | v_22116;
assign v_22120 = v_22118 | v_22119;
assign v_22123 = v_22121 | v_22122;
assign v_22126 = v_22124 | v_22125;
assign v_22129 = v_22127 | v_22128;
assign v_22132 = v_22130 | v_22131;
assign v_22135 = v_22133 | v_22134;
assign v_22138 = v_22136 | v_22137;
assign v_22141 = v_22139 | v_22140;
assign v_22144 = v_22142 | v_22143;
assign v_22147 = v_22145 | v_22146;
assign v_22150 = v_22148 | v_22149;
assign v_22153 = v_22151 | v_22152;
assign v_22156 = v_22154 | v_22155;
assign v_22159 = v_22157 | v_22158;
assign v_22162 = v_22160 | v_22161;
assign v_22165 = v_22163 | v_22164;
assign v_22168 = v_22166 | v_22167;
assign v_22171 = v_22169 | v_22170;
assign v_22174 = v_22172 | v_22173;
assign v_22177 = v_22175 | v_22176;
assign v_22180 = v_22178 | v_22179;
assign v_22183 = v_22181 | v_22182;
assign v_22186 = v_22184 | v_22185;
assign v_22189 = v_22187 | v_22188;
assign v_22192 = v_22190 | v_22191;
assign v_22195 = v_22193 | v_22194;
assign v_22198 = v_22196 | v_22197;
assign v_22201 = v_22199 | v_22200;
assign v_22204 = v_22202 | v_22203;
assign v_22207 = v_22205 | v_22206;
assign v_22210 = v_22208 | v_22209;
assign v_22213 = v_22211 | v_22212;
assign v_22214 = v_22024 | v_22213;
assign v_22215 = v_9630 | ~v_9844;
assign v_22216 = v_9601 | ~v_9712;
assign v_22218 = v_9335 | v_22217;
assign v_22219 = v_9307 | ~v_9554;
assign v_22221 = v_9336 | v_22220;
assign v_22222 = v_9308 | ~v_9422;
assign v_22224 = v_9051 | v_22223;
assign v_22225 = v_9026 | ~v_9266;
assign v_22227 = v_9052 | v_22226;
assign v_22228 = v_9027 | ~v_9134;
assign v_22230 = v_8761 | v_22229;
assign v_22231 = v_8729 | ~v_8984;
assign v_22233 = v_8762 | v_22232;
assign v_22234 = v_8730 | ~v_8852;
assign v_22236 = v_8473 | v_22235;
assign v_22237 = v_8447 | ~v_8688;
assign v_22239 = v_8474 | v_22238;
assign v_22240 = v_8448 | ~v_8556;
assign v_22242 = v_8185 | v_22241;
assign v_22243 = v_8157 | ~v_8404;
assign v_22245 = v_8186 | v_22244;
assign v_22246 = v_8158 | ~v_8272;
assign v_22248 = v_7901 | v_22247;
assign v_22249 = v_7876 | ~v_8116;
assign v_22251 = v_7902 | v_22250;
assign v_22252 = v_7877 | ~v_7984;
assign v_22254 = v_7607 | v_22253;
assign v_22255 = v_7571 | ~v_7834;
assign v_22257 = v_7608 | v_22256;
assign v_22258 = v_7572 | ~v_7702;
assign v_22260 = v_7315 | v_22259;
assign v_22261 = v_7288 | ~v_7530;
assign v_22263 = v_7316 | v_22262;
assign v_22264 = v_7289 | ~v_7398;
assign v_22266 = v_7025 | v_22265;
assign v_22267 = v_6997 | ~v_7244;
assign v_22269 = v_7026 | v_22268;
assign v_22270 = v_6998 | ~v_7112;
assign v_22272 = v_6741 | v_22271;
assign v_22273 = v_6716 | ~v_6956;
assign v_22275 = v_6742 | v_22274;
assign v_22276 = v_6717 | v_6824;
assign v_22278 = v_6451 | v_22277;
assign v_22279 = v_6419 | ~v_6674;
assign v_22281 = v_6452 | v_22280;
assign v_22282 = v_6420 | ~v_6542;
assign v_22284 = v_6163 | v_22283;
assign v_22285 = v_6137 | ~v_6378;
assign v_22287 = v_6164 | v_22286;
assign v_22288 = v_6138 | ~v_6246;
assign v_22290 = v_5875 | v_22289;
assign v_22291 = v_5847 | v_6094;
assign v_22293 = v_5876 | v_22292;
assign v_22294 = v_5848 | ~v_5962;
assign v_22296 = v_5591 | v_22295;
assign v_22297 = v_5566 | v_5806;
assign v_22299 = v_5592 | v_22298;
assign v_22300 = v_5567 | ~v_5674;
assign v_22302 = v_5293 | v_22301;
assign v_22303 = v_5253 | ~v_5524;
assign v_22305 = v_5294 | v_22304;
assign v_22306 = v_5254 | ~v_5392;
assign v_22308 = v_4997 | v_22307;
assign v_22309 = v_4969 | ~v_5212;
assign v_22311 = v_4998 | v_22310;
assign v_22312 = v_4970 | ~v_5080;
assign v_22314 = v_4705 | v_22313;
assign v_22315 = v_4677 | ~v_4924;
assign v_22317 = v_4706 | v_22316;
assign v_22318 = v_4678 | ~v_4792;
assign v_22320 = v_4421 | v_22319;
assign v_22321 = v_4396 | ~v_4636;
assign v_22323 = v_4422 | v_22322;
assign v_22324 = v_4397 | ~v_4504;
assign v_22326 = v_4131 | v_22325;
assign v_22327 = v_4099 | ~v_4354;
assign v_22329 = v_4132 | v_22328;
assign v_22330 = v_4100 | ~v_4222;
assign v_22332 = v_3843 | v_22331;
assign v_22333 = v_3817 | ~v_4058;
assign v_22335 = v_3844 | v_22334;
assign v_22336 = v_3818 | ~v_3926;
assign v_22338 = v_3555 | v_22337;
assign v_22339 = v_3527 | ~v_3774;
assign v_22341 = v_3556 | v_22340;
assign v_22342 = v_3528 | ~v_3642;
assign v_22344 = v_3271 | v_22343;
assign v_22345 = v_3246 | ~v_3486;
assign v_22347 = v_3272 | v_22346;
assign v_22348 = v_3247 | ~v_3354;
assign v_22350 = v_2977 | v_22349;
assign v_22351 = v_2941 | v_3204;
assign v_22353 = v_2978 | v_22352;
assign v_22354 = v_2942 | ~v_3072;
assign v_22356 = v_2685 | v_22355;
assign v_22357 = v_2658 | ~v_2900;
assign v_22359 = v_2686 | v_22358;
assign v_22360 = v_2659 | ~v_2768;
assign v_22362 = v_2395 | v_22361;
assign v_22363 = v_2367 | ~v_2614;
assign v_22365 = v_2396 | v_22364;
assign v_22366 = v_2368 | ~v_2482;
assign v_22368 = v_2111 | v_22367;
assign v_22369 = v_2086 | ~v_2326;
assign v_22371 = v_2112 | v_22370;
assign v_22372 = v_2087 | ~v_2194;
assign v_22374 = v_1821 | v_22373;
assign v_22375 = v_1789 | ~v_2044;
assign v_22377 = v_1822 | v_22376;
assign v_22378 = v_1790 | ~v_1912;
assign v_22380 = v_1533 | v_22379;
assign v_22381 = v_1507 | ~v_1748;
assign v_22383 = v_1534 | v_22382;
assign v_22384 = v_1508 | ~v_1616;
assign v_22386 = v_1245 | v_22385;
assign v_22387 = v_1217 | ~v_1464;
assign v_22389 = v_1246 | v_22388;
assign v_22390 = v_1218 | ~v_1332;
assign v_22392 = v_961 | v_22391;
assign v_22393 = v_936 | ~v_1176;
assign v_22395 = v_962 | v_22394;
assign v_22396 = v_937 | ~v_1044;
assign v_22398 = v_591 | v_22397;
assign v_22399 = v_92 | ~v_898;
assign v_22401 = v_593 | v_22400;
assign v_22402 = v_94 | ~v_771;
assign v_22404 = v_22214 | v_22403;
assign v_22407 = v_22405 | v_22406;
assign v_22410 = v_22408 | v_22409;
assign v_22413 = v_22411 | v_22412;
assign v_22416 = v_22414 | v_22415;
assign v_22419 = v_22417 | v_22418;
assign v_22422 = v_22420 | v_22421;
assign v_22425 = v_22423 | v_22424;
assign v_22428 = v_22426 | v_22427;
assign v_22431 = v_22429 | v_22430;
assign v_22434 = v_22432 | v_22433;
assign v_22437 = v_22435 | v_22436;
assign v_22440 = v_22438 | v_22439;
assign v_22443 = v_22441 | v_22442;
assign v_22446 = v_22444 | v_22445;
assign v_22449 = v_22447 | v_22448;
assign v_22452 = v_22450 | v_22451;
assign v_22455 = v_22453 | v_22454;
assign v_22458 = v_22456 | v_22457;
assign v_22461 = v_22459 | v_22460;
assign v_22464 = v_22462 | v_22463;
assign v_22467 = v_22465 | v_22466;
assign v_22470 = v_22468 | v_22469;
assign v_22473 = v_22471 | v_22472;
assign v_22476 = v_22474 | v_22475;
assign v_22479 = v_22477 | v_22478;
assign v_22482 = v_22480 | v_22481;
assign v_22485 = v_22483 | v_22484;
assign v_22488 = v_22486 | v_22487;
assign v_22491 = v_22489 | v_22490;
assign v_22494 = v_22492 | v_22493;
assign v_22497 = v_22495 | v_22496;
assign v_22500 = v_22498 | v_22499;
assign v_22503 = v_22501 | v_22502;
assign v_22506 = v_22504 | v_22505;
assign v_22509 = v_22507 | v_22508;
assign v_22512 = v_22510 | v_22511;
assign v_22515 = v_22513 | v_22514;
assign v_22518 = v_22516 | v_22517;
assign v_22521 = v_22519 | v_22520;
assign v_22524 = v_22522 | v_22523;
assign v_22527 = v_22525 | v_22526;
assign v_22530 = v_22528 | v_22529;
assign v_22533 = v_22531 | v_22532;
assign v_22536 = v_22534 | v_22535;
assign v_22539 = v_22537 | v_22538;
assign v_22542 = v_22540 | v_22541;
assign v_22545 = v_22543 | v_22544;
assign v_22548 = v_22546 | v_22547;
assign v_22551 = v_22549 | v_22550;
assign v_22554 = v_22552 | v_22553;
assign v_22557 = v_22555 | v_22556;
assign v_22560 = v_22558 | v_22559;
assign v_22563 = v_22561 | v_22562;
assign v_22566 = v_22564 | v_22565;
assign v_22569 = v_22567 | v_22568;
assign v_22572 = v_22570 | v_22571;
assign v_22575 = v_22573 | v_22574;
assign v_22578 = v_22576 | v_22577;
assign v_22581 = v_22579 | v_22580;
assign v_22584 = v_22582 | v_22583;
assign v_22587 = v_22585 | v_22586;
assign v_22590 = v_22588 | v_22589;
assign v_22593 = v_22591 | v_22592;
assign v_22594 = v_22404 | v_22593;
assign v_22595 = v_13540 | v_22594;
assign v_22596 = v_21075 | v_22595;
assign v_22597 = v_10462 | v_22596;
assign v_22601 = v_22599 | v_22600;
assign v_22604 = v_22602 | v_22603;
assign v_22607 = v_22605 | v_22606;
assign v_22610 = v_22608 | v_22609;
assign v_22613 = v_22611 | v_22612;
assign v_22616 = v_22614 | v_22615;
assign v_22619 = v_22617 | v_22618;
assign v_22622 = v_22620 | v_22621;
assign v_22625 = v_22623 | v_22624;
assign v_22628 = v_22626 | v_22627;
assign v_22631 = v_22629 | v_22630;
assign v_22634 = v_22632 | v_22633;
assign v_22637 = v_22635 | v_22636;
assign v_22640 = v_22638 | v_22639;
assign v_22643 = v_22641 | v_22642;
assign v_22646 = v_22644 | v_22645;
assign v_22649 = v_22647 | v_22648;
assign v_22652 = v_22650 | v_22651;
assign v_22655 = v_22653 | v_22654;
assign v_22658 = v_22656 | v_22657;
assign v_22661 = v_22659 | v_22660;
assign v_22664 = v_22662 | v_22663;
assign v_22667 = v_22665 | v_22666;
assign v_22670 = v_22668 | v_22669;
assign v_22673 = v_22671 | v_22672;
assign v_22676 = v_22674 | v_22675;
assign v_22679 = v_22677 | v_22678;
assign v_22682 = v_22680 | v_22681;
assign v_22685 = v_22683 | v_22684;
assign v_22688 = v_22686 | v_22687;
assign v_22691 = v_22689 | v_22690;
assign v_22694 = v_22692 | v_22693;
assign v_22697 = v_22695 | v_22696;
assign v_22700 = v_22698 | v_22699;
assign v_22703 = v_22701 | v_22702;
assign v_22706 = v_22704 | v_22705;
assign v_22709 = v_22707 | v_22708;
assign v_22712 = v_22710 | v_22711;
assign v_22715 = v_22713 | v_22714;
assign v_22718 = v_22716 | v_22717;
assign v_22721 = v_22719 | v_22720;
assign v_22724 = v_22722 | v_22723;
assign v_22727 = v_22725 | v_22726;
assign v_22730 = v_22728 | v_22729;
assign v_22733 = v_22731 | v_22732;
assign v_22736 = v_22734 | v_22735;
assign v_22739 = v_22737 | v_22738;
assign v_22742 = v_22740 | v_22741;
assign v_22745 = v_22743 | v_22744;
assign v_22748 = v_22746 | v_22747;
assign v_22751 = v_22749 | v_22750;
assign v_22754 = v_22752 | v_22753;
assign v_22757 = v_22755 | v_22756;
assign v_22760 = v_22758 | v_22759;
assign v_22763 = v_22761 | v_22762;
assign v_22766 = v_22764 | v_22765;
assign v_22769 = v_22767 | v_22768;
assign v_22772 = v_22770 | v_22771;
assign v_22775 = v_22773 | v_22774;
assign v_22778 = v_22776 | v_22777;
assign v_22781 = v_22779 | v_22780;
assign v_22784 = v_22782 | v_22783;
assign v_22787 = v_22785 | v_22786;
assign v_22788 = v_13153 | v_22787;
assign v_22789 = v_13532 | v_22788;
assign v_22790 = v_13540 | v_22789;
assign v_22791 = v_10462 | v_22790;
assign v_22795 = v_22793 | v_22794;
assign v_22798 = v_22796 | v_22797;
assign v_22801 = v_22799 | v_22800;
assign v_22804 = v_22802 | v_22803;
assign v_22807 = v_22805 | v_22806;
assign v_22810 = v_22808 | v_22809;
assign v_22813 = v_22811 | v_22812;
assign v_22816 = v_22814 | v_22815;
assign v_22819 = v_22817 | v_22818;
assign v_22822 = v_22820 | v_22821;
assign v_22825 = v_22823 | v_22824;
assign v_22828 = v_22826 | v_22827;
assign v_22831 = v_22829 | v_22830;
assign v_22834 = v_22832 | v_22833;
assign v_22837 = v_22835 | v_22836;
assign v_22840 = v_22838 | v_22839;
assign v_22843 = v_22841 | v_22842;
assign v_22846 = v_22844 | v_22845;
assign v_22849 = v_22847 | v_22848;
assign v_22852 = v_22850 | v_22851;
assign v_22855 = v_22853 | v_22854;
assign v_22858 = v_22856 | v_22857;
assign v_22861 = v_22859 | v_22860;
assign v_22864 = v_22862 | v_22863;
assign v_22867 = v_22865 | v_22866;
assign v_22870 = v_22868 | v_22869;
assign v_22873 = v_22871 | v_22872;
assign v_22876 = v_22874 | v_22875;
assign v_22879 = v_22877 | v_22878;
assign v_22882 = v_22880 | v_22881;
assign v_22885 = v_22883 | v_22884;
assign v_22888 = v_22886 | v_22887;
assign v_22891 = v_22889 | v_22890;
assign v_22894 = v_22892 | v_22893;
assign v_22897 = v_22895 | v_22896;
assign v_22900 = v_22898 | v_22899;
assign v_22903 = v_22901 | v_22902;
assign v_22906 = v_22904 | v_22905;
assign v_22909 = v_22907 | v_22908;
assign v_22912 = v_22910 | v_22911;
assign v_22915 = v_22913 | v_22914;
assign v_22918 = v_22916 | v_22917;
assign v_22921 = v_22919 | v_22920;
assign v_22924 = v_22922 | v_22923;
assign v_22927 = v_22925 | v_22926;
assign v_22930 = v_22928 | v_22929;
assign v_22933 = v_22931 | v_22932;
assign v_22936 = v_22934 | v_22935;
assign v_22939 = v_22937 | v_22938;
assign v_22942 = v_22940 | v_22941;
assign v_22945 = v_22943 | v_22944;
assign v_22948 = v_22946 | v_22947;
assign v_22951 = v_22949 | v_22950;
assign v_22954 = v_22952 | v_22953;
assign v_22957 = v_22955 | v_22956;
assign v_22960 = v_22958 | v_22959;
assign v_22963 = v_22961 | v_22962;
assign v_22966 = v_22964 | v_22965;
assign v_22969 = v_22967 | v_22968;
assign v_22972 = v_22970 | v_22971;
assign v_22975 = v_22973 | v_22974;
assign v_22978 = v_22976 | v_22977;
assign v_22981 = v_22979 | v_22980;
assign v_22982 = v_16202 | v_22981;
assign v_22983 = v_16581 | v_22982;
assign v_22984 = v_13540 | v_22983;
assign v_22985 = v_10462 | v_22984;
assign v_22989 = v_22987 | v_22988;
assign v_22992 = v_22990 | v_22991;
assign v_22995 = v_22993 | v_22994;
assign v_22998 = v_22996 | v_22997;
assign v_23001 = v_22999 | v_23000;
assign v_23004 = v_23002 | v_23003;
assign v_23007 = v_23005 | v_23006;
assign v_23010 = v_23008 | v_23009;
assign v_23013 = v_23011 | v_23012;
assign v_23016 = v_23014 | v_23015;
assign v_23019 = v_23017 | v_23018;
assign v_23022 = v_23020 | v_23021;
assign v_23025 = v_23023 | v_23024;
assign v_23028 = v_23026 | v_23027;
assign v_23031 = v_23029 | v_23030;
assign v_23034 = v_23032 | v_23033;
assign v_23037 = v_23035 | v_23036;
assign v_23040 = v_23038 | v_23039;
assign v_23043 = v_23041 | v_23042;
assign v_23046 = v_23044 | v_23045;
assign v_23049 = v_23047 | v_23048;
assign v_23052 = v_23050 | v_23051;
assign v_23055 = v_23053 | v_23054;
assign v_23058 = v_23056 | v_23057;
assign v_23061 = v_23059 | v_23060;
assign v_23064 = v_23062 | v_23063;
assign v_23067 = v_23065 | v_23066;
assign v_23070 = v_23068 | v_23069;
assign v_23073 = v_23071 | v_23072;
assign v_23076 = v_23074 | v_23075;
assign v_23079 = v_23077 | v_23078;
assign v_23082 = v_23080 | v_23081;
assign v_23085 = v_23083 | v_23084;
assign v_23088 = v_23086 | v_23087;
assign v_23091 = v_23089 | v_23090;
assign v_23094 = v_23092 | v_23093;
assign v_23097 = v_23095 | v_23096;
assign v_23100 = v_23098 | v_23099;
assign v_23103 = v_23101 | v_23102;
assign v_23106 = v_23104 | v_23105;
assign v_23109 = v_23107 | v_23108;
assign v_23112 = v_23110 | v_23111;
assign v_23115 = v_23113 | v_23114;
assign v_23118 = v_23116 | v_23117;
assign v_23121 = v_23119 | v_23120;
assign v_23124 = v_23122 | v_23123;
assign v_23127 = v_23125 | v_23126;
assign v_23130 = v_23128 | v_23129;
assign v_23133 = v_23131 | v_23132;
assign v_23136 = v_23134 | v_23135;
assign v_23139 = v_23137 | v_23138;
assign v_23142 = v_23140 | v_23141;
assign v_23145 = v_23143 | v_23144;
assign v_23148 = v_23146 | v_23147;
assign v_23151 = v_23149 | v_23150;
assign v_23154 = v_23152 | v_23153;
assign v_23157 = v_23155 | v_23156;
assign v_23160 = v_23158 | v_23159;
assign v_23163 = v_23161 | v_23162;
assign v_23166 = v_23164 | v_23165;
assign v_23169 = v_23167 | v_23168;
assign v_23172 = v_23170 | v_23171;
assign v_23173 = v_19178 | v_23172;
assign v_23174 = v_19551 | v_23173;
assign v_23175 = v_13540 | v_23174;
assign v_23176 = v_10462 | v_23175;
assign v_23180 = v_23178 | v_23179;
assign v_23183 = v_23181 | v_23182;
assign v_23186 = v_23184 | v_23185;
assign v_23189 = v_23187 | v_23188;
assign v_23192 = v_23190 | v_23191;
assign v_23195 = v_23193 | v_23194;
assign v_23198 = v_23196 | v_23197;
assign v_23201 = v_23199 | v_23200;
assign v_23204 = v_23202 | v_23203;
assign v_23207 = v_23205 | v_23206;
assign v_23210 = v_23208 | v_23209;
assign v_23213 = v_23211 | v_23212;
assign v_23216 = v_23214 | v_23215;
assign v_23219 = v_23217 | v_23218;
assign v_23222 = v_23220 | v_23221;
assign v_23225 = v_23223 | v_23224;
assign v_23228 = v_23226 | v_23227;
assign v_23231 = v_23229 | v_23230;
assign v_23234 = v_23232 | v_23233;
assign v_23237 = v_23235 | v_23236;
assign v_23240 = v_23238 | v_23239;
assign v_23243 = v_23241 | v_23242;
assign v_23246 = v_23244 | v_23245;
assign v_23249 = v_23247 | v_23248;
assign v_23252 = v_23250 | v_23251;
assign v_23255 = v_23253 | v_23254;
assign v_23258 = v_23256 | v_23257;
assign v_23261 = v_23259 | v_23260;
assign v_23264 = v_23262 | v_23263;
assign v_23267 = v_23265 | v_23266;
assign v_23270 = v_23268 | v_23269;
assign v_23273 = v_23271 | v_23272;
assign v_23276 = v_23274 | v_23275;
assign v_23279 = v_23277 | v_23278;
assign v_23282 = v_23280 | v_23281;
assign v_23285 = v_23283 | v_23284;
assign v_23288 = v_23286 | v_23287;
assign v_23291 = v_23289 | v_23290;
assign v_23294 = v_23292 | v_23293;
assign v_23297 = v_23295 | v_23296;
assign v_23300 = v_23298 | v_23299;
assign v_23303 = v_23301 | v_23302;
assign v_23306 = v_23304 | v_23305;
assign v_23309 = v_23307 | v_23308;
assign v_23312 = v_23310 | v_23311;
assign v_23315 = v_23313 | v_23314;
assign v_23318 = v_23316 | v_23317;
assign v_23321 = v_23319 | v_23320;
assign v_23324 = v_23322 | v_23323;
assign v_23327 = v_23325 | v_23326;
assign v_23330 = v_23328 | v_23329;
assign v_23333 = v_23331 | v_23332;
assign v_23336 = v_23334 | v_23335;
assign v_23339 = v_23337 | v_23338;
assign v_23342 = v_23340 | v_23341;
assign v_23345 = v_23343 | v_23344;
assign v_23348 = v_23346 | v_23347;
assign v_23351 = v_23349 | v_23350;
assign v_23354 = v_23352 | v_23353;
assign v_23357 = v_23355 | v_23356;
assign v_23360 = v_23358 | v_23359;
assign v_23363 = v_23361 | v_23362;
assign v_23366 = v_23364 | v_23365;
assign v_23367 = v_22214 | v_23366;
assign v_23368 = v_22593 | v_23367;
assign v_23369 = v_13540 | v_23368;
assign v_23370 = v_10462 | v_23369;
assign v_23372 = v_6094 | v_6122;
assign v_23373 = v_6003 | v_6034;
assign v_23374 = v_6046 | v_23373;
assign v_23375 = v_6058 | v_23374;
assign v_23376 = v_6070 | v_23375;
assign v_23377 = v_6082 | v_23376;
assign v_23378 = v_23372 | v_23377;
assign v_23379 = v_6824 | v_6852;
assign v_23380 = v_6720 | v_6764;
assign v_23381 = v_6776 | v_23380;
assign v_23382 = v_6788 | v_23381;
assign v_23383 = v_6800 | v_23382;
assign v_23384 = v_6812 | v_23383;
assign v_23385 = v_23379 | v_23384;
assign v_23386 = v_5806 | v_5834;
assign v_23387 = v_5715 | v_5746;
assign v_23388 = v_5758 | v_23387;
assign v_23389 = v_5770 | v_23388;
assign v_23390 = v_5782 | v_23389;
assign v_23391 = v_5794 | v_23390;
assign v_23392 = v_23386 | v_23391;
assign v_23393 = v_4263 | v_4294;
assign v_23394 = v_4306 | v_23393;
assign v_23395 = v_4318 | v_23394;
assign v_23396 = v_4330 | v_23395;
assign v_23397 = v_4342 | v_23396;
assign v_23398 = ~v_4354 | v_23397;
assign v_23399 = v_4382 | v_23398;
assign v_23400 = v_13540 | v_23399;
assign v_23401 = v_23392 | v_23400;
assign v_23402 = v_23385 | v_23401;
assign v_23403 = v_23378 | v_23402;
assign v_23404 = v_10462 | v_23403;
assign v_23406 = v_10462 | v_23405;
assign v_23407 = v_23371 | v_23406;
assign v_23408 = v_23177 | v_23407;
assign v_23409 = v_22986 | v_23408;
assign v_23410 = v_22792 | v_23409;
assign v_23411 = v_22598 | v_23410;
assign v_23412 = v_19556 | v_23411;
assign v_23413 = v_16586 | v_23412;
assign v_23414 = v_13544 | v_23413;
assign v_23415 = v_10495 | v_23414;
assign v_23416 = v_10487 | v_23415;
assign v_23417 = v_3 | v_23416;
assign v_23418 = ~v_10465 | v_23417;
assign v_23419 = ~v_563 | v_10494;
assign v_23420 = ~v_361 | v_10493;
assign v_23421 = ~v_807 | v_10492;
assign v_23422 = ~v_96 | v_10491;
assign v_23423 = ~v_10200 | v_10490;
assign v_23424 = ~v_10196 | v_10489;
assign v_23425 = ~v_9903 | v_10488;
assign v_23426 = ~v_9884 | ~v_10415;
assign v_23434 = v_563 | v_10472;
assign v_23435 = v_9644 | ~v_9784;
assign v_23436 = v_9616 | ~v_9652;
assign v_23438 = v_9487 | v_23437;
assign v_23439 = v_9472 | ~v_9494;
assign v_23441 = v_9353 | v_23440;
assign v_23442 = v_9326 | ~v_9362;
assign v_23444 = v_9199 | v_23443;
assign v_23445 = v_9184 | ~v_9206;
assign v_23447 = v_9066 | v_23446;
assign v_23448 = v_9042 | ~v_9074;
assign v_23450 = v_8917 | v_23449;
assign v_23451 = v_8902 | ~v_8924;
assign v_23453 = v_8782 | v_23452;
assign v_23454 = v_8751 | ~v_8792;
assign v_23456 = v_8621 | v_23455;
assign v_23457 = v_8606 | ~v_8628;
assign v_23459 = v_8488 | v_23458;
assign v_23460 = v_8463 | ~v_8496;
assign v_23462 = v_8337 | v_23461;
assign v_23463 = v_8322 | ~v_8344;
assign v_23465 = v_8203 | v_23464;
assign v_23466 = v_8176 | ~v_8212;
assign v_23468 = v_8049 | v_23467;
assign v_23469 = v_8034 | ~v_8056;
assign v_23471 = v_7916 | v_23470;
assign v_23472 = v_7892 | ~v_7924;
assign v_23474 = v_7767 | v_23473;
assign v_23475 = v_7752 | ~v_7774;
assign v_23477 = v_7631 | v_23476;
assign v_23478 = v_7596 | ~v_7642;
assign v_23480 = v_7463 | v_23479;
assign v_23481 = v_7448 | ~v_7470;
assign v_23483 = v_7330 | v_23482;
assign v_23484 = v_7304 | ~v_7338;
assign v_23486 = v_7177 | v_23485;
assign v_23487 = v_7162 | ~v_7184;
assign v_23489 = v_7043 | v_23488;
assign v_23490 = v_7016 | ~v_7052;
assign v_23492 = v_6889 | v_23491;
assign v_23493 = v_6874 | ~v_6896;
assign v_23495 = v_6756 | v_23494;
assign v_23496 = v_6732 | ~v_6764;
assign v_23498 = v_6607 | v_23497;
assign v_23499 = v_6592 | ~v_6614;
assign v_23501 = v_6472 | v_23500;
assign v_23502 = v_6441 | ~v_6482;
assign v_23504 = v_6311 | v_23503;
assign v_23505 = v_6296 | ~v_6318;
assign v_23507 = v_6178 | v_23506;
assign v_23508 = v_6153 | ~v_6186;
assign v_23510 = v_6027 | v_23509;
assign v_23511 = v_6012 | ~v_6034;
assign v_23513 = v_5893 | v_23512;
assign v_23514 = v_5866 | ~v_5902;
assign v_23516 = v_5739 | v_23515;
assign v_23517 = v_5724 | ~v_5746;
assign v_23519 = v_5606 | v_23518;
assign v_23520 = v_5582 | ~v_5614;
assign v_23522 = v_5457 | v_23521;
assign v_23523 = v_5442 | ~v_5464;
assign v_23525 = v_5320 | v_23524;
assign v_23526 = v_5281 | ~v_5332;
assign v_23528 = v_5145 | v_23527;
assign v_23529 = v_5130 | ~v_5152;
assign v_23531 = v_5012 | v_23530;
assign v_23532 = v_4985 | ~v_5020;
assign v_23534 = v_4857 | v_23533;
assign v_23535 = v_4842 | ~v_4864;
assign v_23537 = v_4723 | v_23536;
assign v_23538 = v_4696 | ~v_4732;
assign v_23540 = v_4569 | v_23539;
assign v_23541 = v_4554 | ~v_4576;
assign v_23543 = v_4436 | v_23542;
assign v_23544 = v_4412 | ~v_4444;
assign v_23546 = v_4287 | v_23545;
assign v_23547 = v_4272 | ~v_4294;
assign v_23549 = v_4152 | v_23548;
assign v_23550 = v_4121 | ~v_4162;
assign v_23552 = v_3991 | v_23551;
assign v_23553 = v_3976 | ~v_3998;
assign v_23555 = v_3858 | v_23554;
assign v_23556 = v_3833 | ~v_3866;
assign v_23558 = v_3707 | v_23557;
assign v_23559 = v_3692 | ~v_3714;
assign v_23561 = v_3573 | v_23560;
assign v_23562 = v_3546 | ~v_3582;
assign v_23564 = v_3419 | v_23563;
assign v_23565 = v_3404 | ~v_3426;
assign v_23567 = v_3286 | v_23566;
assign v_23568 = v_3262 | ~v_3294;
assign v_23570 = v_3137 | v_23569;
assign v_23571 = v_3122 | ~v_3144;
assign v_23573 = v_3001 | v_23572;
assign v_23574 = v_2966 | ~v_3012;
assign v_23576 = v_2833 | v_23575;
assign v_23577 = v_2818 | ~v_2840;
assign v_23579 = v_2700 | v_23578;
assign v_23580 = v_2674 | ~v_2708;
assign v_23582 = v_2547 | v_23581;
assign v_23583 = v_2532 | ~v_2554;
assign v_23585 = v_2413 | v_23584;
assign v_23586 = v_2386 | ~v_2422;
assign v_23588 = v_2259 | v_23587;
assign v_23589 = v_2244 | ~v_2266;
assign v_23591 = v_2126 | v_23590;
assign v_23592 = v_2102 | ~v_2134;
assign v_23594 = v_1977 | v_23593;
assign v_23595 = v_1962 | ~v_1984;
assign v_23597 = v_1842 | v_23596;
assign v_23598 = v_1811 | ~v_1852;
assign v_23600 = v_1681 | v_23599;
assign v_23601 = v_1666 | ~v_1688;
assign v_23603 = v_1548 | v_23602;
assign v_23604 = v_1523 | ~v_1556;
assign v_23606 = v_1397 | v_23605;
assign v_23607 = v_1382 | ~v_1404;
assign v_23609 = v_1263 | v_23608;
assign v_23610 = v_1236 | ~v_1272;
assign v_23612 = v_1109 | v_23611;
assign v_23613 = v_1094 | ~v_1116;
assign v_23615 = v_976 | v_23614;
assign v_23616 = v_952 | ~v_984;
assign v_23618 = v_831 | v_23617;
assign v_23619 = v_815 | ~v_838;
assign v_23621 = v_687 | v_23620;
assign v_23622 = v_453 | ~v_721;
assign v_23624 = v_9644 | ~v_9753;
assign v_23625 = ~v_9604 | v_9616;
assign v_23627 = v_9487 | v_23626;
assign v_23628 = ~v_9463 | v_9472;
assign v_23630 = v_9353 | v_23629;
assign v_23631 = ~v_9311 | v_9326;
assign v_23633 = v_9199 | v_23632;
assign v_23634 = ~v_9175 | v_9184;
assign v_23636 = v_9066 | v_23635;
assign v_23637 = ~v_9030 | v_9042;
assign v_23639 = v_8917 | v_23638;
assign v_23640 = ~v_8893 | v_8902;
assign v_23642 = v_8782 | v_23641;
assign v_23643 = ~v_8733 | v_8751;
assign v_23645 = v_8621 | v_23644;
assign v_23646 = ~v_8597 | v_8606;
assign v_23648 = v_8488 | v_23647;
assign v_23649 = ~v_8451 | v_8463;
assign v_23651 = v_8337 | v_23650;
assign v_23652 = ~v_8313 | v_8322;
assign v_23654 = v_8203 | v_23653;
assign v_23655 = ~v_8161 | v_8176;
assign v_23657 = v_8049 | v_23656;
assign v_23658 = ~v_8025 | v_8034;
assign v_23660 = v_7916 | v_23659;
assign v_23661 = ~v_7880 | v_7892;
assign v_23663 = v_7767 | v_23662;
assign v_23664 = ~v_7743 | v_7752;
assign v_23666 = v_7631 | v_23665;
assign v_23667 = ~v_7575 | v_7596;
assign v_23669 = v_7463 | v_23668;
assign v_23670 = ~v_7439 | v_7448;
assign v_23672 = v_7330 | v_23671;
assign v_23673 = ~v_7292 | v_7304;
assign v_23675 = v_7177 | v_23674;
assign v_23676 = ~v_7153 | v_7162;
assign v_23678 = v_7043 | v_23677;
assign v_23679 = ~v_7001 | v_7016;
assign v_23681 = v_6889 | v_23680;
assign v_23682 = ~v_6865 | v_6874;
assign v_23684 = v_6756 | v_23683;
assign v_23685 = ~v_6720 | v_6732;
assign v_23687 = v_6607 | v_23686;
assign v_23688 = ~v_6583 | v_6592;
assign v_23690 = v_6472 | v_23689;
assign v_23691 = ~v_6423 | v_6441;
assign v_23693 = v_6311 | v_23692;
assign v_23694 = ~v_6287 | v_6296;
assign v_23696 = v_6178 | v_23695;
assign v_23697 = ~v_6141 | v_6153;
assign v_23699 = v_6027 | v_23698;
assign v_23700 = ~v_6003 | v_6012;
assign v_23702 = v_5893 | v_23701;
assign v_23703 = ~v_5851 | v_5866;
assign v_23705 = v_5739 | v_23704;
assign v_23706 = ~v_5715 | v_5724;
assign v_23708 = v_5606 | v_23707;
assign v_23709 = ~v_5570 | v_5582;
assign v_23711 = v_5457 | v_23710;
assign v_23712 = ~v_5433 | v_5442;
assign v_23714 = v_5320 | v_23713;
assign v_23715 = ~v_5257 | v_5281;
assign v_23717 = v_5145 | v_23716;
assign v_23718 = ~v_5121 | v_5130;
assign v_23720 = v_5012 | v_23719;
assign v_23721 = ~v_4973 | v_4985;
assign v_23723 = v_4857 | v_23722;
assign v_23724 = ~v_4833 | v_4842;
assign v_23726 = v_4723 | v_23725;
assign v_23727 = ~v_4681 | v_4696;
assign v_23729 = v_4569 | v_23728;
assign v_23730 = ~v_4545 | v_4554;
assign v_23732 = v_4436 | v_23731;
assign v_23733 = ~v_4400 | v_4412;
assign v_23735 = v_4287 | v_23734;
assign v_23736 = ~v_4263 | v_4272;
assign v_23738 = v_4152 | v_23737;
assign v_23739 = ~v_4103 | v_4121;
assign v_23741 = v_3991 | v_23740;
assign v_23742 = ~v_3967 | v_3976;
assign v_23744 = v_3858 | v_23743;
assign v_23745 = ~v_3821 | v_3833;
assign v_23747 = v_3707 | v_23746;
assign v_23748 = ~v_3683 | v_3692;
assign v_23750 = v_3573 | v_23749;
assign v_23751 = ~v_3531 | v_3546;
assign v_23753 = v_3419 | v_23752;
assign v_23754 = ~v_3395 | v_3404;
assign v_23756 = v_3286 | v_23755;
assign v_23757 = ~v_3250 | v_3262;
assign v_23759 = v_3137 | v_23758;
assign v_23760 = ~v_3113 | v_3122;
assign v_23762 = v_3001 | v_23761;
assign v_23763 = ~v_2945 | v_2966;
assign v_23765 = v_2833 | v_23764;
assign v_23766 = ~v_2809 | v_2818;
assign v_23768 = v_2700 | v_23767;
assign v_23769 = ~v_2662 | v_2674;
assign v_23771 = v_2547 | v_23770;
assign v_23772 = ~v_2523 | v_2532;
assign v_23774 = v_2413 | v_23773;
assign v_23775 = ~v_2371 | v_2386;
assign v_23777 = v_2259 | v_23776;
assign v_23778 = ~v_2235 | v_2244;
assign v_23780 = v_2126 | v_23779;
assign v_23781 = ~v_2090 | v_2102;
assign v_23783 = v_1977 | v_23782;
assign v_23784 = ~v_1953 | v_1962;
assign v_23786 = v_1842 | v_23785;
assign v_23787 = ~v_1793 | v_1811;
assign v_23789 = v_1681 | v_23788;
assign v_23790 = ~v_1657 | v_1666;
assign v_23792 = v_1548 | v_23791;
assign v_23793 = ~v_1511 | v_1523;
assign v_23795 = v_1397 | v_23794;
assign v_23796 = ~v_1373 | v_1382;
assign v_23798 = v_1263 | v_23797;
assign v_23799 = ~v_1221 | v_1236;
assign v_23801 = v_1109 | v_23800;
assign v_23802 = ~v_1085 | v_1094;
assign v_23804 = v_976 | v_23803;
assign v_23805 = ~v_940 | v_952;
assign v_23807 = v_831 | v_23806;
assign v_23808 = ~v_804 | v_815;
assign v_23810 = v_687 | v_23809;
assign v_23811 = ~v_98 | v_453;
assign v_23814 = v_9644 | ~v_9796;
assign v_23815 = v_9616 | ~v_9664;
assign v_23817 = v_9487 | v_23816;
assign v_23818 = v_9472 | ~v_9506;
assign v_23820 = v_9353 | v_23819;
assign v_23821 = v_9326 | ~v_9374;
assign v_23823 = v_9199 | v_23822;
assign v_23824 = v_9184 | ~v_9218;
assign v_23826 = v_9066 | v_23825;
assign v_23827 = v_9042 | ~v_9086;
assign v_23829 = v_8917 | v_23828;
assign v_23830 = v_8902 | ~v_8936;
assign v_23832 = v_8782 | v_23831;
assign v_23833 = v_8751 | ~v_8804;
assign v_23835 = v_8621 | v_23834;
assign v_23836 = v_8606 | ~v_8640;
assign v_23838 = v_8488 | v_23837;
assign v_23839 = v_8463 | ~v_8508;
assign v_23841 = v_8337 | v_23840;
assign v_23842 = v_8322 | ~v_8356;
assign v_23844 = v_8203 | v_23843;
assign v_23845 = v_8176 | ~v_8224;
assign v_23847 = v_8049 | v_23846;
assign v_23848 = v_8034 | ~v_8068;
assign v_23850 = v_7916 | v_23849;
assign v_23851 = v_7892 | ~v_7936;
assign v_23853 = v_7767 | v_23852;
assign v_23854 = v_7752 | ~v_7786;
assign v_23856 = v_7631 | v_23855;
assign v_23857 = v_7596 | ~v_7654;
assign v_23859 = v_7463 | v_23858;
assign v_23860 = v_7448 | ~v_7482;
assign v_23862 = v_7330 | v_23861;
assign v_23863 = v_7304 | ~v_7350;
assign v_23865 = v_7177 | v_23864;
assign v_23866 = v_7162 | ~v_7196;
assign v_23868 = v_7043 | v_23867;
assign v_23869 = v_7016 | ~v_7064;
assign v_23871 = v_6889 | v_23870;
assign v_23872 = v_6874 | ~v_6908;
assign v_23874 = v_6756 | v_23873;
assign v_23875 = v_6732 | ~v_6776;
assign v_23877 = v_6607 | v_23876;
assign v_23878 = v_6592 | ~v_6626;
assign v_23880 = v_6472 | v_23879;
assign v_23881 = v_6441 | ~v_6494;
assign v_23883 = v_6311 | v_23882;
assign v_23884 = v_6296 | ~v_6330;
assign v_23886 = v_6178 | v_23885;
assign v_23887 = v_6153 | ~v_6198;
assign v_23889 = v_6027 | v_23888;
assign v_23890 = v_6012 | ~v_6046;
assign v_23892 = v_5893 | v_23891;
assign v_23893 = v_5866 | ~v_5914;
assign v_23895 = v_5739 | v_23894;
assign v_23896 = v_5724 | ~v_5758;
assign v_23898 = v_5606 | v_23897;
assign v_23899 = v_5582 | ~v_5626;
assign v_23901 = v_5457 | v_23900;
assign v_23902 = v_5442 | ~v_5476;
assign v_23904 = v_5320 | v_23903;
assign v_23905 = v_5281 | ~v_5344;
assign v_23907 = v_5145 | v_23906;
assign v_23908 = v_5130 | ~v_5164;
assign v_23910 = v_5012 | v_23909;
assign v_23911 = v_4985 | ~v_5032;
assign v_23913 = v_4857 | v_23912;
assign v_23914 = v_4842 | ~v_4876;
assign v_23916 = v_4723 | v_23915;
assign v_23917 = v_4696 | ~v_4744;
assign v_23919 = v_4569 | v_23918;
assign v_23920 = v_4554 | ~v_4588;
assign v_23922 = v_4436 | v_23921;
assign v_23923 = v_4412 | ~v_4456;
assign v_23925 = v_4287 | v_23924;
assign v_23926 = v_4272 | ~v_4306;
assign v_23928 = v_4152 | v_23927;
assign v_23929 = v_4121 | ~v_4174;
assign v_23931 = v_3991 | v_23930;
assign v_23932 = v_3976 | ~v_4010;
assign v_23934 = v_3858 | v_23933;
assign v_23935 = v_3833 | ~v_3878;
assign v_23937 = v_3707 | v_23936;
assign v_23938 = v_3692 | ~v_3726;
assign v_23940 = v_3573 | v_23939;
assign v_23941 = v_3546 | ~v_3594;
assign v_23943 = v_3419 | v_23942;
assign v_23944 = v_3404 | ~v_3438;
assign v_23946 = v_3286 | v_23945;
assign v_23947 = v_3262 | ~v_3306;
assign v_23949 = v_3137 | v_23948;
assign v_23950 = v_3122 | ~v_3156;
assign v_23952 = v_3001 | v_23951;
assign v_23953 = v_2966 | ~v_3024;
assign v_23955 = v_2833 | v_23954;
assign v_23956 = v_2818 | ~v_2852;
assign v_23958 = v_2700 | v_23957;
assign v_23959 = v_2674 | ~v_2720;
assign v_23961 = v_2547 | v_23960;
assign v_23962 = v_2532 | ~v_2566;
assign v_23964 = v_2413 | v_23963;
assign v_23965 = v_2386 | ~v_2434;
assign v_23967 = v_2259 | v_23966;
assign v_23968 = v_2244 | ~v_2278;
assign v_23970 = v_2126 | v_23969;
assign v_23971 = v_2102 | ~v_2146;
assign v_23973 = v_1977 | v_23972;
assign v_23974 = v_1962 | ~v_1996;
assign v_23976 = v_1842 | v_23975;
assign v_23977 = v_1811 | ~v_1864;
assign v_23979 = v_1681 | v_23978;
assign v_23980 = v_1666 | ~v_1700;
assign v_23982 = v_1548 | v_23981;
assign v_23983 = v_1523 | ~v_1568;
assign v_23985 = v_1397 | v_23984;
assign v_23986 = v_1382 | ~v_1416;
assign v_23988 = v_1263 | v_23987;
assign v_23989 = v_1236 | ~v_1284;
assign v_23991 = v_1109 | v_23990;
assign v_23992 = v_1094 | ~v_1128;
assign v_23994 = v_976 | v_23993;
assign v_23995 = v_952 | ~v_996;
assign v_23997 = v_831 | v_23996;
assign v_23998 = v_815 | ~v_850;
assign v_24000 = v_687 | v_23999;
assign v_24001 = v_453 | ~v_731;
assign v_24004 = v_9644 | ~v_9808;
assign v_24005 = v_9616 | ~v_9676;
assign v_24007 = v_9487 | v_24006;
assign v_24008 = v_9472 | ~v_9518;
assign v_24010 = v_9353 | v_24009;
assign v_24011 = v_9326 | ~v_9386;
assign v_24013 = v_9199 | v_24012;
assign v_24014 = v_9184 | ~v_9230;
assign v_24016 = v_9066 | v_24015;
assign v_24017 = v_9042 | ~v_9098;
assign v_24019 = v_8917 | v_24018;
assign v_24020 = v_8902 | ~v_8948;
assign v_24022 = v_8782 | v_24021;
assign v_24023 = v_8751 | ~v_8816;
assign v_24025 = v_8621 | v_24024;
assign v_24026 = v_8606 | ~v_8652;
assign v_24028 = v_8488 | v_24027;
assign v_24029 = v_8463 | ~v_8520;
assign v_24031 = v_8337 | v_24030;
assign v_24032 = v_8322 | ~v_8368;
assign v_24034 = v_8203 | v_24033;
assign v_24035 = v_8176 | ~v_8236;
assign v_24037 = v_8049 | v_24036;
assign v_24038 = v_8034 | ~v_8080;
assign v_24040 = v_7916 | v_24039;
assign v_24041 = v_7892 | ~v_7948;
assign v_24043 = v_7767 | v_24042;
assign v_24044 = v_7752 | ~v_7798;
assign v_24046 = v_7631 | v_24045;
assign v_24047 = v_7596 | ~v_7666;
assign v_24049 = v_7463 | v_24048;
assign v_24050 = v_7448 | ~v_7494;
assign v_24052 = v_7330 | v_24051;
assign v_24053 = v_7304 | ~v_7362;
assign v_24055 = v_7177 | v_24054;
assign v_24056 = v_7162 | ~v_7208;
assign v_24058 = v_7043 | v_24057;
assign v_24059 = v_7016 | ~v_7076;
assign v_24061 = v_6889 | v_24060;
assign v_24062 = v_6874 | ~v_6920;
assign v_24064 = v_6756 | v_24063;
assign v_24065 = v_6732 | ~v_6788;
assign v_24067 = v_6607 | v_24066;
assign v_24068 = v_6592 | ~v_6638;
assign v_24070 = v_6472 | v_24069;
assign v_24071 = v_6441 | ~v_6506;
assign v_24073 = v_6311 | v_24072;
assign v_24074 = v_6296 | ~v_6342;
assign v_24076 = v_6178 | v_24075;
assign v_24077 = v_6153 | ~v_6210;
assign v_24079 = v_6027 | v_24078;
assign v_24080 = v_6012 | ~v_6058;
assign v_24082 = v_5893 | v_24081;
assign v_24083 = v_5866 | ~v_5926;
assign v_24085 = v_5739 | v_24084;
assign v_24086 = v_5724 | ~v_5770;
assign v_24088 = v_5606 | v_24087;
assign v_24089 = v_5582 | ~v_5638;
assign v_24091 = v_5457 | v_24090;
assign v_24092 = v_5442 | ~v_5488;
assign v_24094 = v_5320 | v_24093;
assign v_24095 = v_5281 | ~v_5356;
assign v_24097 = v_5145 | v_24096;
assign v_24098 = v_5130 | ~v_5176;
assign v_24100 = v_5012 | v_24099;
assign v_24101 = v_4985 | ~v_5044;
assign v_24103 = v_4857 | v_24102;
assign v_24104 = v_4842 | ~v_4888;
assign v_24106 = v_4723 | v_24105;
assign v_24107 = v_4696 | ~v_4756;
assign v_24109 = v_4569 | v_24108;
assign v_24110 = v_4554 | ~v_4600;
assign v_24112 = v_4436 | v_24111;
assign v_24113 = v_4412 | ~v_4468;
assign v_24115 = v_4287 | v_24114;
assign v_24116 = v_4272 | ~v_4318;
assign v_24118 = v_4152 | v_24117;
assign v_24119 = v_4121 | ~v_4186;
assign v_24121 = v_3991 | v_24120;
assign v_24122 = v_3976 | ~v_4022;
assign v_24124 = v_3858 | v_24123;
assign v_24125 = v_3833 | ~v_3890;
assign v_24127 = v_3707 | v_24126;
assign v_24128 = v_3692 | ~v_3738;
assign v_24130 = v_3573 | v_24129;
assign v_24131 = v_3546 | ~v_3606;
assign v_24133 = v_3419 | v_24132;
assign v_24134 = v_3404 | ~v_3450;
assign v_24136 = v_3286 | v_24135;
assign v_24137 = v_3262 | ~v_3318;
assign v_24139 = v_3137 | v_24138;
assign v_24140 = v_3122 | ~v_3168;
assign v_24142 = v_3001 | v_24141;
assign v_24143 = v_2966 | ~v_3036;
assign v_24145 = v_2833 | v_24144;
assign v_24146 = v_2818 | ~v_2864;
assign v_24148 = v_2700 | v_24147;
assign v_24149 = v_2674 | ~v_2732;
assign v_24151 = v_2547 | v_24150;
assign v_24152 = v_2532 | ~v_2578;
assign v_24154 = v_2413 | v_24153;
assign v_24155 = v_2386 | ~v_2446;
assign v_24157 = v_2259 | v_24156;
assign v_24158 = v_2244 | ~v_2290;
assign v_24160 = v_2126 | v_24159;
assign v_24161 = v_2102 | ~v_2158;
assign v_24163 = v_1977 | v_24162;
assign v_24164 = v_1962 | ~v_2008;
assign v_24166 = v_1842 | v_24165;
assign v_24167 = v_1811 | ~v_1876;
assign v_24169 = v_1681 | v_24168;
assign v_24170 = v_1666 | ~v_1712;
assign v_24172 = v_1548 | v_24171;
assign v_24173 = v_1523 | ~v_1580;
assign v_24175 = v_1397 | v_24174;
assign v_24176 = v_1382 | ~v_1428;
assign v_24178 = v_1263 | v_24177;
assign v_24179 = v_1236 | ~v_1296;
assign v_24181 = v_1109 | v_24180;
assign v_24182 = v_1094 | ~v_1140;
assign v_24184 = v_976 | v_24183;
assign v_24185 = v_952 | ~v_1008;
assign v_24187 = v_831 | v_24186;
assign v_24188 = v_815 | ~v_862;
assign v_24190 = v_687 | v_24189;
assign v_24191 = v_453 | ~v_741;
assign v_24194 = v_9644 | ~v_9820;
assign v_24195 = v_9616 | ~v_9688;
assign v_24197 = v_9487 | v_24196;
assign v_24198 = v_9472 | ~v_9530;
assign v_24200 = v_9353 | v_24199;
assign v_24201 = v_9326 | ~v_9398;
assign v_24203 = v_9199 | v_24202;
assign v_24204 = v_9184 | ~v_9242;
assign v_24206 = v_9066 | v_24205;
assign v_24207 = v_9042 | ~v_9110;
assign v_24209 = v_8917 | v_24208;
assign v_24210 = v_8902 | ~v_8960;
assign v_24212 = v_8782 | v_24211;
assign v_24213 = v_8751 | ~v_8828;
assign v_24215 = v_8621 | v_24214;
assign v_24216 = v_8606 | ~v_8664;
assign v_24218 = v_8488 | v_24217;
assign v_24219 = v_8463 | ~v_8532;
assign v_24221 = v_8337 | v_24220;
assign v_24222 = v_8322 | ~v_8380;
assign v_24224 = v_8203 | v_24223;
assign v_24225 = v_8176 | ~v_8248;
assign v_24227 = v_8049 | v_24226;
assign v_24228 = v_8034 | ~v_8092;
assign v_24230 = v_7916 | v_24229;
assign v_24231 = v_7892 | ~v_7960;
assign v_24233 = v_7767 | v_24232;
assign v_24234 = v_7752 | ~v_7810;
assign v_24236 = v_7631 | v_24235;
assign v_24237 = v_7596 | ~v_7678;
assign v_24239 = v_7463 | v_24238;
assign v_24240 = v_7448 | ~v_7506;
assign v_24242 = v_7330 | v_24241;
assign v_24243 = v_7304 | ~v_7374;
assign v_24245 = v_7177 | v_24244;
assign v_24246 = v_7162 | ~v_7220;
assign v_24248 = v_7043 | v_24247;
assign v_24249 = v_7016 | ~v_7088;
assign v_24251 = v_6889 | v_24250;
assign v_24252 = v_6874 | ~v_6932;
assign v_24254 = v_6756 | v_24253;
assign v_24255 = v_6732 | ~v_6800;
assign v_24257 = v_6607 | v_24256;
assign v_24258 = v_6592 | ~v_6650;
assign v_24260 = v_6472 | v_24259;
assign v_24261 = v_6441 | ~v_6518;
assign v_24263 = v_6311 | v_24262;
assign v_24264 = v_6296 | ~v_6354;
assign v_24266 = v_6178 | v_24265;
assign v_24267 = v_6153 | ~v_6222;
assign v_24269 = v_6027 | v_24268;
assign v_24270 = v_6012 | ~v_6070;
assign v_24272 = v_5893 | v_24271;
assign v_24273 = v_5866 | ~v_5938;
assign v_24275 = v_5739 | v_24274;
assign v_24276 = v_5724 | ~v_5782;
assign v_24278 = v_5606 | v_24277;
assign v_24279 = v_5582 | ~v_5650;
assign v_24281 = v_5457 | v_24280;
assign v_24282 = v_5442 | ~v_5500;
assign v_24284 = v_5320 | v_24283;
assign v_24285 = v_5281 | ~v_5368;
assign v_24287 = v_5145 | v_24286;
assign v_24288 = v_5130 | ~v_5188;
assign v_24290 = v_5012 | v_24289;
assign v_24291 = v_4985 | ~v_5056;
assign v_24293 = v_4857 | v_24292;
assign v_24294 = v_4842 | ~v_4900;
assign v_24296 = v_4723 | v_24295;
assign v_24297 = v_4696 | ~v_4768;
assign v_24299 = v_4569 | v_24298;
assign v_24300 = v_4554 | ~v_4612;
assign v_24302 = v_4436 | v_24301;
assign v_24303 = v_4412 | ~v_4480;
assign v_24305 = v_4287 | v_24304;
assign v_24306 = v_4272 | ~v_4330;
assign v_24308 = v_4152 | v_24307;
assign v_24309 = v_4121 | ~v_4198;
assign v_24311 = v_3991 | v_24310;
assign v_24312 = v_3976 | ~v_4034;
assign v_24314 = v_3858 | v_24313;
assign v_24315 = v_3833 | ~v_3902;
assign v_24317 = v_3707 | v_24316;
assign v_24318 = v_3692 | ~v_3750;
assign v_24320 = v_3573 | v_24319;
assign v_24321 = v_3546 | ~v_3618;
assign v_24323 = v_3419 | v_24322;
assign v_24324 = v_3404 | ~v_3462;
assign v_24326 = v_3286 | v_24325;
assign v_24327 = v_3262 | ~v_3330;
assign v_24329 = v_3137 | v_24328;
assign v_24330 = v_3122 | ~v_3180;
assign v_24332 = v_3001 | v_24331;
assign v_24333 = v_2966 | ~v_3048;
assign v_24335 = v_2833 | v_24334;
assign v_24336 = v_2818 | ~v_2876;
assign v_24338 = v_2700 | v_24337;
assign v_24339 = v_2674 | ~v_2744;
assign v_24341 = v_2547 | v_24340;
assign v_24342 = v_2532 | ~v_2590;
assign v_24344 = v_2413 | v_24343;
assign v_24345 = v_2386 | ~v_2458;
assign v_24347 = v_2259 | v_24346;
assign v_24348 = v_2244 | ~v_2302;
assign v_24350 = v_2126 | v_24349;
assign v_24351 = v_2102 | ~v_2170;
assign v_24353 = v_1977 | v_24352;
assign v_24354 = v_1962 | ~v_2020;
assign v_24356 = v_1842 | v_24355;
assign v_24357 = v_1811 | ~v_1888;
assign v_24359 = v_1681 | v_24358;
assign v_24360 = v_1666 | ~v_1724;
assign v_24362 = v_1548 | v_24361;
assign v_24363 = v_1523 | ~v_1592;
assign v_24365 = v_1397 | v_24364;
assign v_24366 = v_1382 | ~v_1440;
assign v_24368 = v_1263 | v_24367;
assign v_24369 = v_1236 | ~v_1308;
assign v_24371 = v_1109 | v_24370;
assign v_24372 = v_1094 | ~v_1152;
assign v_24374 = v_976 | v_24373;
assign v_24375 = v_952 | ~v_1020;
assign v_24377 = v_831 | v_24376;
assign v_24378 = v_815 | ~v_874;
assign v_24380 = v_687 | v_24379;
assign v_24381 = v_453 | ~v_751;
assign v_24384 = v_9644 | ~v_9832;
assign v_24385 = v_9616 | ~v_9700;
assign v_24387 = v_9487 | v_24386;
assign v_24388 = v_9472 | ~v_9542;
assign v_24390 = v_9353 | v_24389;
assign v_24391 = v_9326 | ~v_9410;
assign v_24393 = v_9199 | v_24392;
assign v_24394 = v_9184 | ~v_9254;
assign v_24396 = v_9066 | v_24395;
assign v_24397 = v_9042 | ~v_9122;
assign v_24399 = v_8917 | v_24398;
assign v_24400 = v_8902 | ~v_8972;
assign v_24402 = v_8782 | v_24401;
assign v_24403 = v_8751 | ~v_8840;
assign v_24405 = v_8621 | v_24404;
assign v_24406 = v_8606 | ~v_8676;
assign v_24408 = v_8488 | v_24407;
assign v_24409 = v_8463 | ~v_8544;
assign v_24411 = v_8337 | v_24410;
assign v_24412 = v_8322 | ~v_8392;
assign v_24414 = v_8203 | v_24413;
assign v_24415 = v_8176 | ~v_8260;
assign v_24417 = v_8049 | v_24416;
assign v_24418 = v_8034 | ~v_8104;
assign v_24420 = v_7916 | v_24419;
assign v_24421 = v_7892 | ~v_7972;
assign v_24423 = v_7767 | v_24422;
assign v_24424 = v_7752 | ~v_7822;
assign v_24426 = v_7631 | v_24425;
assign v_24427 = v_7596 | ~v_7690;
assign v_24429 = v_7463 | v_24428;
assign v_24430 = v_7448 | ~v_7518;
assign v_24432 = v_7330 | v_24431;
assign v_24433 = v_7304 | ~v_7386;
assign v_24435 = v_7177 | v_24434;
assign v_24436 = v_7162 | ~v_7232;
assign v_24438 = v_7043 | v_24437;
assign v_24439 = v_7016 | ~v_7100;
assign v_24441 = v_6889 | v_24440;
assign v_24442 = v_6874 | ~v_6944;
assign v_24444 = v_6756 | v_24443;
assign v_24445 = v_6732 | ~v_6812;
assign v_24447 = v_6607 | v_24446;
assign v_24448 = v_6592 | ~v_6662;
assign v_24450 = v_6472 | v_24449;
assign v_24451 = v_6441 | ~v_6530;
assign v_24453 = v_6311 | v_24452;
assign v_24454 = v_6296 | ~v_6366;
assign v_24456 = v_6178 | v_24455;
assign v_24457 = v_6153 | ~v_6234;
assign v_24459 = v_6027 | v_24458;
assign v_24460 = v_6012 | ~v_6082;
assign v_24462 = v_5893 | v_24461;
assign v_24463 = v_5866 | ~v_5950;
assign v_24465 = v_5739 | v_24464;
assign v_24466 = v_5724 | ~v_5794;
assign v_24468 = v_5606 | v_24467;
assign v_24469 = v_5582 | ~v_5662;
assign v_24471 = v_5457 | v_24470;
assign v_24472 = v_5442 | ~v_5512;
assign v_24474 = v_5320 | v_24473;
assign v_24475 = v_5281 | ~v_5380;
assign v_24477 = v_5145 | v_24476;
assign v_24478 = v_5130 | ~v_5200;
assign v_24480 = v_5012 | v_24479;
assign v_24481 = v_4985 | ~v_5068;
assign v_24483 = v_4857 | v_24482;
assign v_24484 = v_4842 | ~v_4912;
assign v_24486 = v_4723 | v_24485;
assign v_24487 = v_4696 | ~v_4780;
assign v_24489 = v_4569 | v_24488;
assign v_24490 = v_4554 | ~v_4624;
assign v_24492 = v_4436 | v_24491;
assign v_24493 = v_4412 | ~v_4492;
assign v_24495 = v_4287 | v_24494;
assign v_24496 = v_4272 | ~v_4342;
assign v_24498 = v_4152 | v_24497;
assign v_24499 = v_4121 | ~v_4210;
assign v_24501 = v_3991 | v_24500;
assign v_24502 = v_3976 | ~v_4046;
assign v_24504 = v_3858 | v_24503;
assign v_24505 = v_3833 | ~v_3914;
assign v_24507 = v_3707 | v_24506;
assign v_24508 = v_3692 | ~v_3762;
assign v_24510 = v_3573 | v_24509;
assign v_24511 = v_3546 | ~v_3630;
assign v_24513 = v_3419 | v_24512;
assign v_24514 = v_3404 | ~v_3474;
assign v_24516 = v_3286 | v_24515;
assign v_24517 = v_3262 | ~v_3342;
assign v_24519 = v_3137 | v_24518;
assign v_24520 = v_3122 | ~v_3192;
assign v_24522 = v_3001 | v_24521;
assign v_24523 = v_2966 | ~v_3060;
assign v_24525 = v_2833 | v_24524;
assign v_24526 = v_2818 | ~v_2888;
assign v_24528 = v_2700 | v_24527;
assign v_24529 = v_2674 | ~v_2756;
assign v_24531 = v_2547 | v_24530;
assign v_24532 = v_2532 | ~v_2602;
assign v_24534 = v_2413 | v_24533;
assign v_24535 = v_2386 | ~v_2470;
assign v_24537 = v_2259 | v_24536;
assign v_24538 = v_2244 | ~v_2314;
assign v_24540 = v_2126 | v_24539;
assign v_24541 = v_2102 | ~v_2182;
assign v_24543 = v_1977 | v_24542;
assign v_24544 = v_1962 | ~v_2032;
assign v_24546 = v_1842 | v_24545;
assign v_24547 = v_1811 | ~v_1900;
assign v_24549 = v_1681 | v_24548;
assign v_24550 = v_1666 | ~v_1736;
assign v_24552 = v_1548 | v_24551;
assign v_24553 = v_1523 | ~v_1604;
assign v_24555 = v_1397 | v_24554;
assign v_24556 = v_1382 | ~v_1452;
assign v_24558 = v_1263 | v_24557;
assign v_24559 = v_1236 | ~v_1320;
assign v_24561 = v_1109 | v_24560;
assign v_24562 = v_1094 | ~v_1164;
assign v_24564 = v_976 | v_24563;
assign v_24565 = v_952 | ~v_1032;
assign v_24567 = v_831 | v_24566;
assign v_24568 = v_815 | ~v_886;
assign v_24570 = v_687 | v_24569;
assign v_24571 = v_453 | ~v_761;
assign v_24574 = v_9644 | ~v_9844;
assign v_24575 = v_9616 | ~v_9712;
assign v_24577 = v_9487 | v_24576;
assign v_24578 = v_9472 | ~v_9554;
assign v_24580 = v_9353 | v_24579;
assign v_24581 = v_9326 | ~v_9422;
assign v_24583 = v_9199 | v_24582;
assign v_24584 = v_9184 | ~v_9266;
assign v_24586 = v_9066 | v_24585;
assign v_24587 = v_9042 | ~v_9134;
assign v_24589 = v_8917 | v_24588;
assign v_24590 = v_8902 | ~v_8984;
assign v_24592 = v_8782 | v_24591;
assign v_24593 = v_8751 | ~v_8852;
assign v_24595 = v_8621 | v_24594;
assign v_24596 = v_8606 | ~v_8688;
assign v_24598 = v_8488 | v_24597;
assign v_24599 = v_8463 | ~v_8556;
assign v_24601 = v_8337 | v_24600;
assign v_24602 = v_8322 | ~v_8404;
assign v_24604 = v_8203 | v_24603;
assign v_24605 = v_8176 | ~v_8272;
assign v_24607 = v_8049 | v_24606;
assign v_24608 = v_8034 | ~v_8116;
assign v_24610 = v_7916 | v_24609;
assign v_24611 = v_7892 | ~v_7984;
assign v_24613 = v_7767 | v_24612;
assign v_24614 = v_7752 | ~v_7834;
assign v_24616 = v_7631 | v_24615;
assign v_24617 = v_7596 | ~v_7702;
assign v_24619 = v_7463 | v_24618;
assign v_24620 = v_7448 | ~v_7530;
assign v_24622 = v_7330 | v_24621;
assign v_24623 = v_7304 | ~v_7398;
assign v_24625 = v_7177 | v_24624;
assign v_24626 = v_7162 | ~v_7244;
assign v_24628 = v_7043 | v_24627;
assign v_24629 = v_7016 | ~v_7112;
assign v_24631 = v_6889 | v_24630;
assign v_24632 = v_6874 | ~v_6956;
assign v_24634 = v_6756 | v_24633;
assign v_24635 = v_6732 | v_6824;
assign v_24637 = v_6607 | v_24636;
assign v_24638 = v_6592 | ~v_6674;
assign v_24640 = v_6472 | v_24639;
assign v_24641 = v_6441 | ~v_6542;
assign v_24643 = v_6311 | v_24642;
assign v_24644 = v_6296 | ~v_6378;
assign v_24646 = v_6178 | v_24645;
assign v_24647 = v_6153 | ~v_6246;
assign v_24649 = v_6027 | v_24648;
assign v_24650 = v_6012 | v_6094;
assign v_24652 = v_5893 | v_24651;
assign v_24653 = v_5866 | ~v_5962;
assign v_24655 = v_5739 | v_24654;
assign v_24656 = v_5724 | v_5806;
assign v_24658 = v_5606 | v_24657;
assign v_24659 = v_5582 | ~v_5674;
assign v_24661 = v_5457 | v_24660;
assign v_24662 = v_5442 | ~v_5524;
assign v_24664 = v_5320 | v_24663;
assign v_24665 = v_5281 | ~v_5392;
assign v_24667 = v_5145 | v_24666;
assign v_24668 = v_5130 | ~v_5212;
assign v_24670 = v_5012 | v_24669;
assign v_24671 = v_4985 | ~v_5080;
assign v_24673 = v_4857 | v_24672;
assign v_24674 = v_4842 | ~v_4924;
assign v_24676 = v_4723 | v_24675;
assign v_24677 = v_4696 | ~v_4792;
assign v_24679 = v_4569 | v_24678;
assign v_24680 = v_4554 | ~v_4636;
assign v_24682 = v_4436 | v_24681;
assign v_24683 = v_4412 | ~v_4504;
assign v_24685 = v_4287 | v_24684;
assign v_24686 = v_4272 | ~v_4354;
assign v_24688 = v_4152 | v_24687;
assign v_24689 = v_4121 | ~v_4222;
assign v_24691 = v_3991 | v_24690;
assign v_24692 = v_3976 | ~v_4058;
assign v_24694 = v_3858 | v_24693;
assign v_24695 = v_3833 | ~v_3926;
assign v_24697 = v_3707 | v_24696;
assign v_24698 = v_3692 | ~v_3774;
assign v_24700 = v_3573 | v_24699;
assign v_24701 = v_3546 | ~v_3642;
assign v_24703 = v_3419 | v_24702;
assign v_24704 = v_3404 | ~v_3486;
assign v_24706 = v_3286 | v_24705;
assign v_24707 = v_3262 | ~v_3354;
assign v_24709 = v_3137 | v_24708;
assign v_24710 = v_3122 | v_3204;
assign v_24712 = v_3001 | v_24711;
assign v_24713 = v_2966 | ~v_3072;
assign v_24715 = v_2833 | v_24714;
assign v_24716 = v_2818 | ~v_2900;
assign v_24718 = v_2700 | v_24717;
assign v_24719 = v_2674 | ~v_2768;
assign v_24721 = v_2547 | v_24720;
assign v_24722 = v_2532 | ~v_2614;
assign v_24724 = v_2413 | v_24723;
assign v_24725 = v_2386 | ~v_2482;
assign v_24727 = v_2259 | v_24726;
assign v_24728 = v_2244 | ~v_2326;
assign v_24730 = v_2126 | v_24729;
assign v_24731 = v_2102 | ~v_2194;
assign v_24733 = v_1977 | v_24732;
assign v_24734 = v_1962 | ~v_2044;
assign v_24736 = v_1842 | v_24735;
assign v_24737 = v_1811 | ~v_1912;
assign v_24739 = v_1681 | v_24738;
assign v_24740 = v_1666 | ~v_1748;
assign v_24742 = v_1548 | v_24741;
assign v_24743 = v_1523 | ~v_1616;
assign v_24745 = v_1397 | v_24744;
assign v_24746 = v_1382 | ~v_1464;
assign v_24748 = v_1263 | v_24747;
assign v_24749 = v_1236 | ~v_1332;
assign v_24751 = v_1109 | v_24750;
assign v_24752 = v_1094 | ~v_1176;
assign v_24754 = v_976 | v_24753;
assign v_24755 = v_952 | ~v_1044;
assign v_24757 = v_831 | v_24756;
assign v_24758 = v_815 | ~v_898;
assign v_24760 = v_687 | v_24759;
assign v_24761 = v_453 | ~v_771;
assign v_24764 = v_9644 | v_9872;
assign v_24765 = v_9616 | v_9740;
assign v_24767 = v_9487 | v_24766;
assign v_24768 = v_9472 | v_9582;
assign v_24770 = v_9353 | v_24769;
assign v_24771 = v_9326 | v_9450;
assign v_24773 = v_9199 | v_24772;
assign v_24774 = v_9184 | v_9294;
assign v_24776 = v_9066 | v_24775;
assign v_24777 = v_9042 | v_9162;
assign v_24779 = v_8917 | v_24778;
assign v_24780 = v_8902 | v_9012;
assign v_24782 = v_8782 | v_24781;
assign v_24783 = v_8751 | v_8880;
assign v_24785 = v_8621 | v_24784;
assign v_24786 = v_8606 | v_8716;
assign v_24788 = v_8488 | v_24787;
assign v_24789 = v_8463 | v_8584;
assign v_24791 = v_8337 | v_24790;
assign v_24792 = v_8322 | ~v_8432;
assign v_24794 = v_8203 | v_24793;
assign v_24795 = v_8176 | ~v_8300;
assign v_24797 = v_8049 | v_24796;
assign v_24798 = v_8034 | ~v_8144;
assign v_24800 = v_7916 | v_24799;
assign v_24801 = v_7892 | v_8012;
assign v_24803 = v_7767 | v_24802;
assign v_24804 = v_7752 | v_7862;
assign v_24806 = v_7631 | v_24805;
assign v_24807 = v_7596 | v_7730;
assign v_24809 = v_7463 | v_24808;
assign v_24810 = v_7448 | v_7558;
assign v_24812 = v_7330 | v_24811;
assign v_24813 = v_7304 | v_7426;
assign v_24815 = v_7177 | v_24814;
assign v_24816 = v_7162 | ~v_7272;
assign v_24818 = v_7043 | v_24817;
assign v_24819 = v_7016 | v_7140;
assign v_24821 = v_6889 | v_24820;
assign v_24822 = v_6874 | ~v_6984;
assign v_24824 = v_6756 | v_24823;
assign v_24825 = v_6732 | ~v_6852;
assign v_24827 = v_6607 | v_24826;
assign v_24828 = v_6592 | ~v_6702;
assign v_24830 = v_6472 | v_24829;
assign v_24831 = v_6441 | v_6570;
assign v_24833 = v_6311 | v_24832;
assign v_24834 = v_6296 | v_6406;
assign v_24836 = v_6178 | v_24835;
assign v_24837 = v_6153 | ~v_6274;
assign v_24839 = v_6027 | v_24838;
assign v_24840 = v_6012 | ~v_6122;
assign v_24842 = v_5893 | v_24841;
assign v_24843 = v_5866 | ~v_5990;
assign v_24845 = v_5739 | v_24844;
assign v_24846 = v_5724 | ~v_5834;
assign v_24848 = v_5606 | v_24847;
assign v_24849 = v_5582 | ~v_5702;
assign v_24851 = v_5457 | v_24850;
assign v_24852 = v_5442 | ~v_5552;
assign v_24854 = v_5320 | v_24853;
assign v_24855 = v_5281 | v_5420;
assign v_24857 = v_5145 | v_24856;
assign v_24858 = v_5130 | v_5240;
assign v_24860 = v_5012 | v_24859;
assign v_24861 = v_4985 | ~v_5108;
assign v_24863 = v_4857 | v_24862;
assign v_24864 = v_4842 | ~v_4952;
assign v_24866 = v_4723 | v_24865;
assign v_24867 = v_4696 | ~v_4820;
assign v_24869 = v_4569 | v_24868;
assign v_24870 = v_4554 | ~v_4664;
assign v_24872 = v_4436 | v_24871;
assign v_24873 = v_4412 | ~v_4532;
assign v_24875 = v_4287 | v_24874;
assign v_24876 = v_4272 | ~v_4382;
assign v_24878 = v_4152 | v_24877;
assign v_24879 = v_4121 | v_4250;
assign v_24881 = v_3991 | v_24880;
assign v_24882 = v_3976 | v_4086;
assign v_24884 = v_3858 | v_24883;
assign v_24885 = v_3833 | v_3954;
assign v_24887 = v_3707 | v_24886;
assign v_24888 = v_3692 | v_3802;
assign v_24890 = v_3573 | v_24889;
assign v_24891 = v_3546 | v_3670;
assign v_24893 = v_3419 | v_24892;
assign v_24894 = v_3404 | ~v_3514;
assign v_24896 = v_3286 | v_24895;
assign v_24897 = v_3262 | v_3382;
assign v_24899 = v_3137 | v_24898;
assign v_24900 = v_3122 | ~v_3232;
assign v_24902 = v_3001 | v_24901;
assign v_24903 = v_2966 | v_3100;
assign v_24905 = v_2833 | v_24904;
assign v_24906 = v_2818 | v_2928;
assign v_24908 = v_2700 | v_24907;
assign v_24909 = v_2674 | v_2796;
assign v_24911 = v_2547 | v_24910;
assign v_24912 = v_2532 | v_2642;
assign v_24914 = v_2413 | v_24913;
assign v_24915 = v_2386 | v_2510;
assign v_24917 = v_2259 | v_24916;
assign v_24918 = v_2244 | ~v_2354;
assign v_24920 = v_2126 | v_24919;
assign v_24921 = v_2102 | ~v_2222;
assign v_24923 = v_1977 | v_24922;
assign v_24924 = v_1962 | ~v_2072;
assign v_24926 = v_1842 | v_24925;
assign v_24927 = v_1811 | v_1940;
assign v_24929 = v_1681 | v_24928;
assign v_24930 = v_1666 | v_1776;
assign v_24932 = v_1548 | v_24931;
assign v_24933 = v_1523 | v_1644;
assign v_24935 = v_1397 | v_24934;
assign v_24936 = v_1382 | v_1492;
assign v_24938 = v_1263 | v_24937;
assign v_24939 = v_1236 | v_1360;
assign v_24941 = v_1109 | v_24940;
assign v_24942 = v_1094 | v_1204;
assign v_24944 = v_976 | v_24943;
assign v_24945 = v_952 | v_1072;
assign v_24947 = v_831 | v_24946;
assign v_24948 = v_815 | v_922;
assign v_24950 = v_687 | v_24949;
assign v_24951 = v_453 | v_793;
assign v_24954 = v_9646 | ~v_9784;
assign v_24955 = v_9618 | ~v_9652;
assign v_24957 = v_9488 | v_24956;
assign v_24958 = v_9473 | ~v_9494;
assign v_24960 = v_9356 | v_24959;
assign v_24961 = v_9329 | ~v_9362;
assign v_24963 = v_9200 | v_24962;
assign v_24964 = v_9185 | ~v_9206;
assign v_24966 = v_9068 | v_24965;
assign v_24967 = v_9044 | ~v_9074;
assign v_24969 = v_8918 | v_24968;
assign v_24970 = v_8903 | ~v_8924;
assign v_24972 = v_8786 | v_24971;
assign v_24973 = v_8755 | ~v_8792;
assign v_24975 = v_8622 | v_24974;
assign v_24976 = v_8607 | ~v_8628;
assign v_24978 = v_8490 | v_24977;
assign v_24979 = v_8465 | ~v_8496;
assign v_24981 = v_8338 | v_24980;
assign v_24982 = v_8323 | ~v_8344;
assign v_24984 = v_8206 | v_24983;
assign v_24985 = v_8179 | ~v_8212;
assign v_24987 = v_8050 | v_24986;
assign v_24988 = v_8035 | ~v_8056;
assign v_24990 = v_7918 | v_24989;
assign v_24991 = v_7894 | ~v_7924;
assign v_24993 = v_7768 | v_24992;
assign v_24994 = v_7753 | ~v_7774;
assign v_24996 = v_7636 | v_24995;
assign v_24997 = v_7601 | ~v_7642;
assign v_24999 = v_7464 | v_24998;
assign v_25000 = v_7449 | ~v_7470;
assign v_25002 = v_7332 | v_25001;
assign v_25003 = v_7306 | ~v_7338;
assign v_25005 = v_7178 | v_25004;
assign v_25006 = v_7163 | ~v_7184;
assign v_25008 = v_7046 | v_25007;
assign v_25009 = v_7019 | ~v_7052;
assign v_25011 = v_6890 | v_25010;
assign v_25012 = v_6875 | ~v_6896;
assign v_25014 = v_6758 | v_25013;
assign v_25015 = v_6734 | ~v_6764;
assign v_25017 = v_6608 | v_25016;
assign v_25018 = v_6593 | ~v_6614;
assign v_25020 = v_6476 | v_25019;
assign v_25021 = v_6445 | ~v_6482;
assign v_25023 = v_6312 | v_25022;
assign v_25024 = v_6297 | ~v_6318;
assign v_25026 = v_6180 | v_25025;
assign v_25027 = v_6155 | ~v_6186;
assign v_25029 = v_6028 | v_25028;
assign v_25030 = v_6013 | ~v_6034;
assign v_25032 = v_5896 | v_25031;
assign v_25033 = v_5869 | ~v_5902;
assign v_25035 = v_5740 | v_25034;
assign v_25036 = v_5725 | ~v_5746;
assign v_25038 = v_5608 | v_25037;
assign v_25039 = v_5584 | ~v_5614;
assign v_25041 = v_5458 | v_25040;
assign v_25042 = v_5443 | ~v_5464;
assign v_25044 = v_5326 | v_25043;
assign v_25045 = v_5287 | ~v_5332;
assign v_25047 = v_5146 | v_25046;
assign v_25048 = v_5131 | ~v_5152;
assign v_25050 = v_5014 | v_25049;
assign v_25051 = v_4987 | ~v_5020;
assign v_25053 = v_4858 | v_25052;
assign v_25054 = v_4843 | ~v_4864;
assign v_25056 = v_4726 | v_25055;
assign v_25057 = v_4699 | ~v_4732;
assign v_25059 = v_4570 | v_25058;
assign v_25060 = v_4555 | ~v_4576;
assign v_25062 = v_4438 | v_25061;
assign v_25063 = v_4414 | ~v_4444;
assign v_25065 = v_4288 | v_25064;
assign v_25066 = v_4273 | ~v_4294;
assign v_25068 = v_4156 | v_25067;
assign v_25069 = v_4125 | ~v_4162;
assign v_25071 = v_3992 | v_25070;
assign v_25072 = v_3977 | ~v_3998;
assign v_25074 = v_3860 | v_25073;
assign v_25075 = v_3835 | ~v_3866;
assign v_25077 = v_3708 | v_25076;
assign v_25078 = v_3693 | ~v_3714;
assign v_25080 = v_3576 | v_25079;
assign v_25081 = v_3549 | ~v_3582;
assign v_25083 = v_3420 | v_25082;
assign v_25084 = v_3405 | ~v_3426;
assign v_25086 = v_3288 | v_25085;
assign v_25087 = v_3264 | ~v_3294;
assign v_25089 = v_3138 | v_25088;
assign v_25090 = v_3123 | ~v_3144;
assign v_25092 = v_3006 | v_25091;
assign v_25093 = v_2971 | ~v_3012;
assign v_25095 = v_2834 | v_25094;
assign v_25096 = v_2819 | ~v_2840;
assign v_25098 = v_2702 | v_25097;
assign v_25099 = v_2676 | ~v_2708;
assign v_25101 = v_2548 | v_25100;
assign v_25102 = v_2533 | ~v_2554;
assign v_25104 = v_2416 | v_25103;
assign v_25105 = v_2389 | ~v_2422;
assign v_25107 = v_2260 | v_25106;
assign v_25108 = v_2245 | ~v_2266;
assign v_25110 = v_2128 | v_25109;
assign v_25111 = v_2104 | ~v_2134;
assign v_25113 = v_1978 | v_25112;
assign v_25114 = v_1963 | ~v_1984;
assign v_25116 = v_1846 | v_25115;
assign v_25117 = v_1815 | ~v_1852;
assign v_25119 = v_1682 | v_25118;
assign v_25120 = v_1667 | ~v_1688;
assign v_25122 = v_1550 | v_25121;
assign v_25123 = v_1525 | ~v_1556;
assign v_25125 = v_1398 | v_25124;
assign v_25126 = v_1383 | ~v_1404;
assign v_25128 = v_1266 | v_25127;
assign v_25129 = v_1239 | ~v_1272;
assign v_25131 = v_1110 | v_25130;
assign v_25132 = v_1095 | ~v_1116;
assign v_25134 = v_978 | v_25133;
assign v_25135 = v_954 | ~v_984;
assign v_25137 = v_832 | v_25136;
assign v_25138 = v_816 | ~v_838;
assign v_25140 = v_715 | v_25139;
assign v_25141 = v_561 | ~v_721;
assign v_25143 = v_9646 | ~v_9753;
assign v_25144 = ~v_9604 | v_9618;
assign v_25146 = v_9488 | v_25145;
assign v_25147 = ~v_9463 | v_9473;
assign v_25149 = v_9356 | v_25148;
assign v_25150 = ~v_9311 | v_9329;
assign v_25152 = v_9200 | v_25151;
assign v_25153 = ~v_9175 | v_9185;
assign v_25155 = v_9068 | v_25154;
assign v_25156 = ~v_9030 | v_9044;
assign v_25158 = v_8918 | v_25157;
assign v_25159 = ~v_8893 | v_8903;
assign v_25161 = v_8786 | v_25160;
assign v_25162 = ~v_8733 | v_8755;
assign v_25164 = v_8622 | v_25163;
assign v_25165 = ~v_8597 | v_8607;
assign v_25167 = v_8490 | v_25166;
assign v_25168 = ~v_8451 | v_8465;
assign v_25170 = v_8338 | v_25169;
assign v_25171 = ~v_8313 | v_8323;
assign v_25173 = v_8206 | v_25172;
assign v_25174 = ~v_8161 | v_8179;
assign v_25176 = v_8050 | v_25175;
assign v_25177 = ~v_8025 | v_8035;
assign v_25179 = v_7918 | v_25178;
assign v_25180 = ~v_7880 | v_7894;
assign v_25182 = v_7768 | v_25181;
assign v_25183 = ~v_7743 | v_7753;
assign v_25185 = v_7636 | v_25184;
assign v_25186 = ~v_7575 | v_7601;
assign v_25188 = v_7464 | v_25187;
assign v_25189 = ~v_7439 | v_7449;
assign v_25191 = v_7332 | v_25190;
assign v_25192 = ~v_7292 | v_7306;
assign v_25194 = v_7178 | v_25193;
assign v_25195 = ~v_7153 | v_7163;
assign v_25197 = v_7046 | v_25196;
assign v_25198 = ~v_7001 | v_7019;
assign v_25200 = v_6890 | v_25199;
assign v_25201 = ~v_6865 | v_6875;
assign v_25203 = v_6758 | v_25202;
assign v_25204 = ~v_6720 | v_6734;
assign v_25206 = v_6608 | v_25205;
assign v_25207 = ~v_6583 | v_6593;
assign v_25209 = v_6476 | v_25208;
assign v_25210 = ~v_6423 | v_6445;
assign v_25212 = v_6312 | v_25211;
assign v_25213 = ~v_6287 | v_6297;
assign v_25215 = v_6180 | v_25214;
assign v_25216 = ~v_6141 | v_6155;
assign v_25218 = v_6028 | v_25217;
assign v_25219 = ~v_6003 | v_6013;
assign v_25221 = v_5896 | v_25220;
assign v_25222 = ~v_5851 | v_5869;
assign v_25224 = v_5740 | v_25223;
assign v_25225 = ~v_5715 | v_5725;
assign v_25227 = v_5608 | v_25226;
assign v_25228 = ~v_5570 | v_5584;
assign v_25230 = v_5458 | v_25229;
assign v_25231 = ~v_5433 | v_5443;
assign v_25233 = v_5326 | v_25232;
assign v_25234 = ~v_5257 | v_5287;
assign v_25236 = v_5146 | v_25235;
assign v_25237 = ~v_5121 | v_5131;
assign v_25239 = v_5014 | v_25238;
assign v_25240 = ~v_4973 | v_4987;
assign v_25242 = v_4858 | v_25241;
assign v_25243 = ~v_4833 | v_4843;
assign v_25245 = v_4726 | v_25244;
assign v_25246 = ~v_4681 | v_4699;
assign v_25248 = v_4570 | v_25247;
assign v_25249 = ~v_4545 | v_4555;
assign v_25251 = v_4438 | v_25250;
assign v_25252 = ~v_4400 | v_4414;
assign v_25254 = v_4288 | v_25253;
assign v_25255 = ~v_4263 | v_4273;
assign v_25257 = v_4156 | v_25256;
assign v_25258 = ~v_4103 | v_4125;
assign v_25260 = v_3992 | v_25259;
assign v_25261 = ~v_3967 | v_3977;
assign v_25263 = v_3860 | v_25262;
assign v_25264 = ~v_3821 | v_3835;
assign v_25266 = v_3708 | v_25265;
assign v_25267 = ~v_3683 | v_3693;
assign v_25269 = v_3576 | v_25268;
assign v_25270 = ~v_3531 | v_3549;
assign v_25272 = v_3420 | v_25271;
assign v_25273 = ~v_3395 | v_3405;
assign v_25275 = v_3288 | v_25274;
assign v_25276 = ~v_3250 | v_3264;
assign v_25278 = v_3138 | v_25277;
assign v_25279 = ~v_3113 | v_3123;
assign v_25281 = v_3006 | v_25280;
assign v_25282 = ~v_2945 | v_2971;
assign v_25284 = v_2834 | v_25283;
assign v_25285 = ~v_2809 | v_2819;
assign v_25287 = v_2702 | v_25286;
assign v_25288 = ~v_2662 | v_2676;
assign v_25290 = v_2548 | v_25289;
assign v_25291 = ~v_2523 | v_2533;
assign v_25293 = v_2416 | v_25292;
assign v_25294 = ~v_2371 | v_2389;
assign v_25296 = v_2260 | v_25295;
assign v_25297 = ~v_2235 | v_2245;
assign v_25299 = v_2128 | v_25298;
assign v_25300 = ~v_2090 | v_2104;
assign v_25302 = v_1978 | v_25301;
assign v_25303 = ~v_1953 | v_1963;
assign v_25305 = v_1846 | v_25304;
assign v_25306 = ~v_1793 | v_1815;
assign v_25308 = v_1682 | v_25307;
assign v_25309 = ~v_1657 | v_1667;
assign v_25311 = v_1550 | v_25310;
assign v_25312 = ~v_1511 | v_1525;
assign v_25314 = v_1398 | v_25313;
assign v_25315 = ~v_1373 | v_1383;
assign v_25317 = v_1266 | v_25316;
assign v_25318 = ~v_1221 | v_1239;
assign v_25320 = v_1110 | v_25319;
assign v_25321 = ~v_1085 | v_1095;
assign v_25323 = v_978 | v_25322;
assign v_25324 = ~v_940 | v_954;
assign v_25326 = v_832 | v_25325;
assign v_25327 = ~v_804 | v_816;
assign v_25329 = v_715 | v_25328;
assign v_25330 = ~v_98 | v_561;
assign v_25333 = v_9646 | ~v_9796;
assign v_25334 = v_9618 | ~v_9664;
assign v_25336 = v_9488 | v_25335;
assign v_25337 = v_9473 | ~v_9506;
assign v_25339 = v_9356 | v_25338;
assign v_25340 = v_9329 | ~v_9374;
assign v_25342 = v_9200 | v_25341;
assign v_25343 = v_9185 | ~v_9218;
assign v_25345 = v_9068 | v_25344;
assign v_25346 = v_9044 | ~v_9086;
assign v_25348 = v_8918 | v_25347;
assign v_25349 = v_8903 | ~v_8936;
assign v_25351 = v_8786 | v_25350;
assign v_25352 = v_8755 | ~v_8804;
assign v_25354 = v_8622 | v_25353;
assign v_25355 = v_8607 | ~v_8640;
assign v_25357 = v_8490 | v_25356;
assign v_25358 = v_8465 | ~v_8508;
assign v_25360 = v_8338 | v_25359;
assign v_25361 = v_8323 | ~v_8356;
assign v_25363 = v_8206 | v_25362;
assign v_25364 = v_8179 | ~v_8224;
assign v_25366 = v_8050 | v_25365;
assign v_25367 = v_8035 | ~v_8068;
assign v_25369 = v_7918 | v_25368;
assign v_25370 = v_7894 | ~v_7936;
assign v_25372 = v_7768 | v_25371;
assign v_25373 = v_7753 | ~v_7786;
assign v_25375 = v_7636 | v_25374;
assign v_25376 = v_7601 | ~v_7654;
assign v_25378 = v_7464 | v_25377;
assign v_25379 = v_7449 | ~v_7482;
assign v_25381 = v_7332 | v_25380;
assign v_25382 = v_7306 | ~v_7350;
assign v_25384 = v_7178 | v_25383;
assign v_25385 = v_7163 | ~v_7196;
assign v_25387 = v_7046 | v_25386;
assign v_25388 = v_7019 | ~v_7064;
assign v_25390 = v_6890 | v_25389;
assign v_25391 = v_6875 | ~v_6908;
assign v_25393 = v_6758 | v_25392;
assign v_25394 = v_6734 | ~v_6776;
assign v_25396 = v_6608 | v_25395;
assign v_25397 = v_6593 | ~v_6626;
assign v_25399 = v_6476 | v_25398;
assign v_25400 = v_6445 | ~v_6494;
assign v_25402 = v_6312 | v_25401;
assign v_25403 = v_6297 | ~v_6330;
assign v_25405 = v_6180 | v_25404;
assign v_25406 = v_6155 | ~v_6198;
assign v_25408 = v_6028 | v_25407;
assign v_25409 = v_6013 | ~v_6046;
assign v_25411 = v_5896 | v_25410;
assign v_25412 = v_5869 | ~v_5914;
assign v_25414 = v_5740 | v_25413;
assign v_25415 = v_5725 | ~v_5758;
assign v_25417 = v_5608 | v_25416;
assign v_25418 = v_5584 | ~v_5626;
assign v_25420 = v_5458 | v_25419;
assign v_25421 = v_5443 | ~v_5476;
assign v_25423 = v_5326 | v_25422;
assign v_25424 = v_5287 | ~v_5344;
assign v_25426 = v_5146 | v_25425;
assign v_25427 = v_5131 | ~v_5164;
assign v_25429 = v_5014 | v_25428;
assign v_25430 = v_4987 | ~v_5032;
assign v_25432 = v_4858 | v_25431;
assign v_25433 = v_4843 | ~v_4876;
assign v_25435 = v_4726 | v_25434;
assign v_25436 = v_4699 | ~v_4744;
assign v_25438 = v_4570 | v_25437;
assign v_25439 = v_4555 | ~v_4588;
assign v_25441 = v_4438 | v_25440;
assign v_25442 = v_4414 | ~v_4456;
assign v_25444 = v_4288 | v_25443;
assign v_25445 = v_4273 | ~v_4306;
assign v_25447 = v_4156 | v_25446;
assign v_25448 = v_4125 | ~v_4174;
assign v_25450 = v_3992 | v_25449;
assign v_25451 = v_3977 | ~v_4010;
assign v_25453 = v_3860 | v_25452;
assign v_25454 = v_3835 | ~v_3878;
assign v_25456 = v_3708 | v_25455;
assign v_25457 = v_3693 | ~v_3726;
assign v_25459 = v_3576 | v_25458;
assign v_25460 = v_3549 | ~v_3594;
assign v_25462 = v_3420 | v_25461;
assign v_25463 = v_3405 | ~v_3438;
assign v_25465 = v_3288 | v_25464;
assign v_25466 = v_3264 | ~v_3306;
assign v_25468 = v_3138 | v_25467;
assign v_25469 = v_3123 | ~v_3156;
assign v_25471 = v_3006 | v_25470;
assign v_25472 = v_2971 | ~v_3024;
assign v_25474 = v_2834 | v_25473;
assign v_25475 = v_2819 | ~v_2852;
assign v_25477 = v_2702 | v_25476;
assign v_25478 = v_2676 | ~v_2720;
assign v_25480 = v_2548 | v_25479;
assign v_25481 = v_2533 | ~v_2566;
assign v_25483 = v_2416 | v_25482;
assign v_25484 = v_2389 | ~v_2434;
assign v_25486 = v_2260 | v_25485;
assign v_25487 = v_2245 | ~v_2278;
assign v_25489 = v_2128 | v_25488;
assign v_25490 = v_2104 | ~v_2146;
assign v_25492 = v_1978 | v_25491;
assign v_25493 = v_1963 | ~v_1996;
assign v_25495 = v_1846 | v_25494;
assign v_25496 = v_1815 | ~v_1864;
assign v_25498 = v_1682 | v_25497;
assign v_25499 = v_1667 | ~v_1700;
assign v_25501 = v_1550 | v_25500;
assign v_25502 = v_1525 | ~v_1568;
assign v_25504 = v_1398 | v_25503;
assign v_25505 = v_1383 | ~v_1416;
assign v_25507 = v_1266 | v_25506;
assign v_25508 = v_1239 | ~v_1284;
assign v_25510 = v_1110 | v_25509;
assign v_25511 = v_1095 | ~v_1128;
assign v_25513 = v_978 | v_25512;
assign v_25514 = v_954 | ~v_996;
assign v_25516 = v_832 | v_25515;
assign v_25517 = v_816 | ~v_850;
assign v_25519 = v_715 | v_25518;
assign v_25520 = v_561 | ~v_731;
assign v_25523 = v_9646 | ~v_9808;
assign v_25524 = v_9618 | ~v_9676;
assign v_25526 = v_9488 | v_25525;
assign v_25527 = v_9473 | ~v_9518;
assign v_25529 = v_9356 | v_25528;
assign v_25530 = v_9329 | ~v_9386;
assign v_25532 = v_9200 | v_25531;
assign v_25533 = v_9185 | ~v_9230;
assign v_25535 = v_9068 | v_25534;
assign v_25536 = v_9044 | ~v_9098;
assign v_25538 = v_8918 | v_25537;
assign v_25539 = v_8903 | ~v_8948;
assign v_25541 = v_8786 | v_25540;
assign v_25542 = v_8755 | ~v_8816;
assign v_25544 = v_8622 | v_25543;
assign v_25545 = v_8607 | ~v_8652;
assign v_25547 = v_8490 | v_25546;
assign v_25548 = v_8465 | ~v_8520;
assign v_25550 = v_8338 | v_25549;
assign v_25551 = v_8323 | ~v_8368;
assign v_25553 = v_8206 | v_25552;
assign v_25554 = v_8179 | ~v_8236;
assign v_25556 = v_8050 | v_25555;
assign v_25557 = v_8035 | ~v_8080;
assign v_25559 = v_7918 | v_25558;
assign v_25560 = v_7894 | ~v_7948;
assign v_25562 = v_7768 | v_25561;
assign v_25563 = v_7753 | ~v_7798;
assign v_25565 = v_7636 | v_25564;
assign v_25566 = v_7601 | ~v_7666;
assign v_25568 = v_7464 | v_25567;
assign v_25569 = v_7449 | ~v_7494;
assign v_25571 = v_7332 | v_25570;
assign v_25572 = v_7306 | ~v_7362;
assign v_25574 = v_7178 | v_25573;
assign v_25575 = v_7163 | ~v_7208;
assign v_25577 = v_7046 | v_25576;
assign v_25578 = v_7019 | ~v_7076;
assign v_25580 = v_6890 | v_25579;
assign v_25581 = v_6875 | ~v_6920;
assign v_25583 = v_6758 | v_25582;
assign v_25584 = v_6734 | ~v_6788;
assign v_25586 = v_6608 | v_25585;
assign v_25587 = v_6593 | ~v_6638;
assign v_25589 = v_6476 | v_25588;
assign v_25590 = v_6445 | ~v_6506;
assign v_25592 = v_6312 | v_25591;
assign v_25593 = v_6297 | ~v_6342;
assign v_25595 = v_6180 | v_25594;
assign v_25596 = v_6155 | ~v_6210;
assign v_25598 = v_6028 | v_25597;
assign v_25599 = v_6013 | ~v_6058;
assign v_25601 = v_5896 | v_25600;
assign v_25602 = v_5869 | ~v_5926;
assign v_25604 = v_5740 | v_25603;
assign v_25605 = v_5725 | ~v_5770;
assign v_25607 = v_5608 | v_25606;
assign v_25608 = v_5584 | ~v_5638;
assign v_25610 = v_5458 | v_25609;
assign v_25611 = v_5443 | ~v_5488;
assign v_25613 = v_5326 | v_25612;
assign v_25614 = v_5287 | ~v_5356;
assign v_25616 = v_5146 | v_25615;
assign v_25617 = v_5131 | ~v_5176;
assign v_25619 = v_5014 | v_25618;
assign v_25620 = v_4987 | ~v_5044;
assign v_25622 = v_4858 | v_25621;
assign v_25623 = v_4843 | ~v_4888;
assign v_25625 = v_4726 | v_25624;
assign v_25626 = v_4699 | ~v_4756;
assign v_25628 = v_4570 | v_25627;
assign v_25629 = v_4555 | ~v_4600;
assign v_25631 = v_4438 | v_25630;
assign v_25632 = v_4414 | ~v_4468;
assign v_25634 = v_4288 | v_25633;
assign v_25635 = v_4273 | ~v_4318;
assign v_25637 = v_4156 | v_25636;
assign v_25638 = v_4125 | ~v_4186;
assign v_25640 = v_3992 | v_25639;
assign v_25641 = v_3977 | ~v_4022;
assign v_25643 = v_3860 | v_25642;
assign v_25644 = v_3835 | ~v_3890;
assign v_25646 = v_3708 | v_25645;
assign v_25647 = v_3693 | ~v_3738;
assign v_25649 = v_3576 | v_25648;
assign v_25650 = v_3549 | ~v_3606;
assign v_25652 = v_3420 | v_25651;
assign v_25653 = v_3405 | ~v_3450;
assign v_25655 = v_3288 | v_25654;
assign v_25656 = v_3264 | ~v_3318;
assign v_25658 = v_3138 | v_25657;
assign v_25659 = v_3123 | ~v_3168;
assign v_25661 = v_3006 | v_25660;
assign v_25662 = v_2971 | ~v_3036;
assign v_25664 = v_2834 | v_25663;
assign v_25665 = v_2819 | ~v_2864;
assign v_25667 = v_2702 | v_25666;
assign v_25668 = v_2676 | ~v_2732;
assign v_25670 = v_2548 | v_25669;
assign v_25671 = v_2533 | ~v_2578;
assign v_25673 = v_2416 | v_25672;
assign v_25674 = v_2389 | ~v_2446;
assign v_25676 = v_2260 | v_25675;
assign v_25677 = v_2245 | ~v_2290;
assign v_25679 = v_2128 | v_25678;
assign v_25680 = v_2104 | ~v_2158;
assign v_25682 = v_1978 | v_25681;
assign v_25683 = v_1963 | ~v_2008;
assign v_25685 = v_1846 | v_25684;
assign v_25686 = v_1815 | ~v_1876;
assign v_25688 = v_1682 | v_25687;
assign v_25689 = v_1667 | ~v_1712;
assign v_25691 = v_1550 | v_25690;
assign v_25692 = v_1525 | ~v_1580;
assign v_25694 = v_1398 | v_25693;
assign v_25695 = v_1383 | ~v_1428;
assign v_25697 = v_1266 | v_25696;
assign v_25698 = v_1239 | ~v_1296;
assign v_25700 = v_1110 | v_25699;
assign v_25701 = v_1095 | ~v_1140;
assign v_25703 = v_978 | v_25702;
assign v_25704 = v_954 | ~v_1008;
assign v_25706 = v_832 | v_25705;
assign v_25707 = v_816 | ~v_862;
assign v_25709 = v_715 | v_25708;
assign v_25710 = v_561 | ~v_741;
assign v_25713 = v_9646 | ~v_9820;
assign v_25714 = v_9618 | ~v_9688;
assign v_25716 = v_9488 | v_25715;
assign v_25717 = v_9473 | ~v_9530;
assign v_25719 = v_9356 | v_25718;
assign v_25720 = v_9329 | ~v_9398;
assign v_25722 = v_9200 | v_25721;
assign v_25723 = v_9185 | ~v_9242;
assign v_25725 = v_9068 | v_25724;
assign v_25726 = v_9044 | ~v_9110;
assign v_25728 = v_8918 | v_25727;
assign v_25729 = v_8903 | ~v_8960;
assign v_25731 = v_8786 | v_25730;
assign v_25732 = v_8755 | ~v_8828;
assign v_25734 = v_8622 | v_25733;
assign v_25735 = v_8607 | ~v_8664;
assign v_25737 = v_8490 | v_25736;
assign v_25738 = v_8465 | ~v_8532;
assign v_25740 = v_8338 | v_25739;
assign v_25741 = v_8323 | ~v_8380;
assign v_25743 = v_8206 | v_25742;
assign v_25744 = v_8179 | ~v_8248;
assign v_25746 = v_8050 | v_25745;
assign v_25747 = v_8035 | ~v_8092;
assign v_25749 = v_7918 | v_25748;
assign v_25750 = v_7894 | ~v_7960;
assign v_25752 = v_7768 | v_25751;
assign v_25753 = v_7753 | ~v_7810;
assign v_25755 = v_7636 | v_25754;
assign v_25756 = v_7601 | ~v_7678;
assign v_25758 = v_7464 | v_25757;
assign v_25759 = v_7449 | ~v_7506;
assign v_25761 = v_7332 | v_25760;
assign v_25762 = v_7306 | ~v_7374;
assign v_25764 = v_7178 | v_25763;
assign v_25765 = v_7163 | ~v_7220;
assign v_25767 = v_7046 | v_25766;
assign v_25768 = v_7019 | ~v_7088;
assign v_25770 = v_6890 | v_25769;
assign v_25771 = v_6875 | ~v_6932;
assign v_25773 = v_6758 | v_25772;
assign v_25774 = v_6734 | ~v_6800;
assign v_25776 = v_6608 | v_25775;
assign v_25777 = v_6593 | ~v_6650;
assign v_25779 = v_6476 | v_25778;
assign v_25780 = v_6445 | ~v_6518;
assign v_25782 = v_6312 | v_25781;
assign v_25783 = v_6297 | ~v_6354;
assign v_25785 = v_6180 | v_25784;
assign v_25786 = v_6155 | ~v_6222;
assign v_25788 = v_6028 | v_25787;
assign v_25789 = v_6013 | ~v_6070;
assign v_25791 = v_5896 | v_25790;
assign v_25792 = v_5869 | ~v_5938;
assign v_25794 = v_5740 | v_25793;
assign v_25795 = v_5725 | ~v_5782;
assign v_25797 = v_5608 | v_25796;
assign v_25798 = v_5584 | ~v_5650;
assign v_25800 = v_5458 | v_25799;
assign v_25801 = v_5443 | ~v_5500;
assign v_25803 = v_5326 | v_25802;
assign v_25804 = v_5287 | ~v_5368;
assign v_25806 = v_5146 | v_25805;
assign v_25807 = v_5131 | ~v_5188;
assign v_25809 = v_5014 | v_25808;
assign v_25810 = v_4987 | ~v_5056;
assign v_25812 = v_4858 | v_25811;
assign v_25813 = v_4843 | ~v_4900;
assign v_25815 = v_4726 | v_25814;
assign v_25816 = v_4699 | ~v_4768;
assign v_25818 = v_4570 | v_25817;
assign v_25819 = v_4555 | ~v_4612;
assign v_25821 = v_4438 | v_25820;
assign v_25822 = v_4414 | ~v_4480;
assign v_25824 = v_4288 | v_25823;
assign v_25825 = v_4273 | ~v_4330;
assign v_25827 = v_4156 | v_25826;
assign v_25828 = v_4125 | ~v_4198;
assign v_25830 = v_3992 | v_25829;
assign v_25831 = v_3977 | ~v_4034;
assign v_25833 = v_3860 | v_25832;
assign v_25834 = v_3835 | ~v_3902;
assign v_25836 = v_3708 | v_25835;
assign v_25837 = v_3693 | ~v_3750;
assign v_25839 = v_3576 | v_25838;
assign v_25840 = v_3549 | ~v_3618;
assign v_25842 = v_3420 | v_25841;
assign v_25843 = v_3405 | ~v_3462;
assign v_25845 = v_3288 | v_25844;
assign v_25846 = v_3264 | ~v_3330;
assign v_25848 = v_3138 | v_25847;
assign v_25849 = v_3123 | ~v_3180;
assign v_25851 = v_3006 | v_25850;
assign v_25852 = v_2971 | ~v_3048;
assign v_25854 = v_2834 | v_25853;
assign v_25855 = v_2819 | ~v_2876;
assign v_25857 = v_2702 | v_25856;
assign v_25858 = v_2676 | ~v_2744;
assign v_25860 = v_2548 | v_25859;
assign v_25861 = v_2533 | ~v_2590;
assign v_25863 = v_2416 | v_25862;
assign v_25864 = v_2389 | ~v_2458;
assign v_25866 = v_2260 | v_25865;
assign v_25867 = v_2245 | ~v_2302;
assign v_25869 = v_2128 | v_25868;
assign v_25870 = v_2104 | ~v_2170;
assign v_25872 = v_1978 | v_25871;
assign v_25873 = v_1963 | ~v_2020;
assign v_25875 = v_1846 | v_25874;
assign v_25876 = v_1815 | ~v_1888;
assign v_25878 = v_1682 | v_25877;
assign v_25879 = v_1667 | ~v_1724;
assign v_25881 = v_1550 | v_25880;
assign v_25882 = v_1525 | ~v_1592;
assign v_25884 = v_1398 | v_25883;
assign v_25885 = v_1383 | ~v_1440;
assign v_25887 = v_1266 | v_25886;
assign v_25888 = v_1239 | ~v_1308;
assign v_25890 = v_1110 | v_25889;
assign v_25891 = v_1095 | ~v_1152;
assign v_25893 = v_978 | v_25892;
assign v_25894 = v_954 | ~v_1020;
assign v_25896 = v_832 | v_25895;
assign v_25897 = v_816 | ~v_874;
assign v_25899 = v_715 | v_25898;
assign v_25900 = v_561 | ~v_751;
assign v_25903 = v_9646 | ~v_9832;
assign v_25904 = v_9618 | ~v_9700;
assign v_25906 = v_9488 | v_25905;
assign v_25907 = v_9473 | ~v_9542;
assign v_25909 = v_9356 | v_25908;
assign v_25910 = v_9329 | ~v_9410;
assign v_25912 = v_9200 | v_25911;
assign v_25913 = v_9185 | ~v_9254;
assign v_25915 = v_9068 | v_25914;
assign v_25916 = v_9044 | ~v_9122;
assign v_25918 = v_8918 | v_25917;
assign v_25919 = v_8903 | ~v_8972;
assign v_25921 = v_8786 | v_25920;
assign v_25922 = v_8755 | ~v_8840;
assign v_25924 = v_8622 | v_25923;
assign v_25925 = v_8607 | ~v_8676;
assign v_25927 = v_8490 | v_25926;
assign v_25928 = v_8465 | ~v_8544;
assign v_25930 = v_8338 | v_25929;
assign v_25931 = v_8323 | ~v_8392;
assign v_25933 = v_8206 | v_25932;
assign v_25934 = v_8179 | ~v_8260;
assign v_25936 = v_8050 | v_25935;
assign v_25937 = v_8035 | ~v_8104;
assign v_25939 = v_7918 | v_25938;
assign v_25940 = v_7894 | ~v_7972;
assign v_25942 = v_7768 | v_25941;
assign v_25943 = v_7753 | ~v_7822;
assign v_25945 = v_7636 | v_25944;
assign v_25946 = v_7601 | ~v_7690;
assign v_25948 = v_7464 | v_25947;
assign v_25949 = v_7449 | ~v_7518;
assign v_25951 = v_7332 | v_25950;
assign v_25952 = v_7306 | ~v_7386;
assign v_25954 = v_7178 | v_25953;
assign v_25955 = v_7163 | ~v_7232;
assign v_25957 = v_7046 | v_25956;
assign v_25958 = v_7019 | ~v_7100;
assign v_25960 = v_6890 | v_25959;
assign v_25961 = v_6875 | ~v_6944;
assign v_25963 = v_6758 | v_25962;
assign v_25964 = v_6734 | ~v_6812;
assign v_25966 = v_6608 | v_25965;
assign v_25967 = v_6593 | ~v_6662;
assign v_25969 = v_6476 | v_25968;
assign v_25970 = v_6445 | ~v_6530;
assign v_25972 = v_6312 | v_25971;
assign v_25973 = v_6297 | ~v_6366;
assign v_25975 = v_6180 | v_25974;
assign v_25976 = v_6155 | ~v_6234;
assign v_25978 = v_6028 | v_25977;
assign v_25979 = v_6013 | ~v_6082;
assign v_25981 = v_5896 | v_25980;
assign v_25982 = v_5869 | ~v_5950;
assign v_25984 = v_5740 | v_25983;
assign v_25985 = v_5725 | ~v_5794;
assign v_25987 = v_5608 | v_25986;
assign v_25988 = v_5584 | ~v_5662;
assign v_25990 = v_5458 | v_25989;
assign v_25991 = v_5443 | ~v_5512;
assign v_25993 = v_5326 | v_25992;
assign v_25994 = v_5287 | ~v_5380;
assign v_25996 = v_5146 | v_25995;
assign v_25997 = v_5131 | ~v_5200;
assign v_25999 = v_5014 | v_25998;
assign v_26000 = v_4987 | ~v_5068;
assign v_26002 = v_4858 | v_26001;
assign v_26003 = v_4843 | ~v_4912;
assign v_26005 = v_4726 | v_26004;
assign v_26006 = v_4699 | ~v_4780;
assign v_26008 = v_4570 | v_26007;
assign v_26009 = v_4555 | ~v_4624;
assign v_26011 = v_4438 | v_26010;
assign v_26012 = v_4414 | ~v_4492;
assign v_26014 = v_4288 | v_26013;
assign v_26015 = v_4273 | ~v_4342;
assign v_26017 = v_4156 | v_26016;
assign v_26018 = v_4125 | ~v_4210;
assign v_26020 = v_3992 | v_26019;
assign v_26021 = v_3977 | ~v_4046;
assign v_26023 = v_3860 | v_26022;
assign v_26024 = v_3835 | ~v_3914;
assign v_26026 = v_3708 | v_26025;
assign v_26027 = v_3693 | ~v_3762;
assign v_26029 = v_3576 | v_26028;
assign v_26030 = v_3549 | ~v_3630;
assign v_26032 = v_3420 | v_26031;
assign v_26033 = v_3405 | ~v_3474;
assign v_26035 = v_3288 | v_26034;
assign v_26036 = v_3264 | ~v_3342;
assign v_26038 = v_3138 | v_26037;
assign v_26039 = v_3123 | ~v_3192;
assign v_26041 = v_3006 | v_26040;
assign v_26042 = v_2971 | ~v_3060;
assign v_26044 = v_2834 | v_26043;
assign v_26045 = v_2819 | ~v_2888;
assign v_26047 = v_2702 | v_26046;
assign v_26048 = v_2676 | ~v_2756;
assign v_26050 = v_2548 | v_26049;
assign v_26051 = v_2533 | ~v_2602;
assign v_26053 = v_2416 | v_26052;
assign v_26054 = v_2389 | ~v_2470;
assign v_26056 = v_2260 | v_26055;
assign v_26057 = v_2245 | ~v_2314;
assign v_26059 = v_2128 | v_26058;
assign v_26060 = v_2104 | ~v_2182;
assign v_26062 = v_1978 | v_26061;
assign v_26063 = v_1963 | ~v_2032;
assign v_26065 = v_1846 | v_26064;
assign v_26066 = v_1815 | ~v_1900;
assign v_26068 = v_1682 | v_26067;
assign v_26069 = v_1667 | ~v_1736;
assign v_26071 = v_1550 | v_26070;
assign v_26072 = v_1525 | ~v_1604;
assign v_26074 = v_1398 | v_26073;
assign v_26075 = v_1383 | ~v_1452;
assign v_26077 = v_1266 | v_26076;
assign v_26078 = v_1239 | ~v_1320;
assign v_26080 = v_1110 | v_26079;
assign v_26081 = v_1095 | ~v_1164;
assign v_26083 = v_978 | v_26082;
assign v_26084 = v_954 | ~v_1032;
assign v_26086 = v_832 | v_26085;
assign v_26087 = v_816 | ~v_886;
assign v_26089 = v_715 | v_26088;
assign v_26090 = v_561 | ~v_761;
assign v_26094 = v_9646 | v_9872;
assign v_26095 = v_9618 | v_9740;
assign v_26097 = v_9488 | v_26096;
assign v_26098 = v_9473 | v_9582;
assign v_26100 = v_9356 | v_26099;
assign v_26101 = v_9329 | v_9450;
assign v_26103 = v_9200 | v_26102;
assign v_26104 = v_9185 | v_9294;
assign v_26106 = v_9068 | v_26105;
assign v_26107 = v_9044 | v_9162;
assign v_26109 = v_8918 | v_26108;
assign v_26110 = v_8903 | v_9012;
assign v_26112 = v_8786 | v_26111;
assign v_26113 = v_8755 | v_8880;
assign v_26115 = v_8622 | v_26114;
assign v_26116 = v_8607 | v_8716;
assign v_26118 = v_8490 | v_26117;
assign v_26119 = v_8465 | v_8584;
assign v_26121 = v_8338 | v_26120;
assign v_26122 = v_8323 | ~v_8432;
assign v_26124 = v_8206 | v_26123;
assign v_26125 = v_8179 | ~v_8300;
assign v_26127 = v_8050 | v_26126;
assign v_26128 = v_8035 | ~v_8144;
assign v_26130 = v_7918 | v_26129;
assign v_26131 = v_7894 | v_8012;
assign v_26133 = v_7768 | v_26132;
assign v_26134 = v_7753 | v_7862;
assign v_26136 = v_7636 | v_26135;
assign v_26137 = v_7601 | v_7730;
assign v_26139 = v_7464 | v_26138;
assign v_26140 = v_7449 | v_7558;
assign v_26142 = v_7332 | v_26141;
assign v_26143 = v_7306 | v_7426;
assign v_26145 = v_7178 | v_26144;
assign v_26146 = v_7163 | ~v_7272;
assign v_26148 = v_7046 | v_26147;
assign v_26149 = v_7019 | v_7140;
assign v_26151 = v_6890 | v_26150;
assign v_26152 = v_6875 | ~v_6984;
assign v_26154 = v_6758 | v_26153;
assign v_26155 = v_6734 | ~v_6852;
assign v_26157 = v_6608 | v_26156;
assign v_26158 = v_6593 | ~v_6702;
assign v_26160 = v_6476 | v_26159;
assign v_26161 = v_6445 | v_6570;
assign v_26163 = v_6312 | v_26162;
assign v_26164 = v_6297 | v_6406;
assign v_26166 = v_6180 | v_26165;
assign v_26167 = v_6155 | ~v_6274;
assign v_26169 = v_6028 | v_26168;
assign v_26170 = v_6013 | ~v_6122;
assign v_26172 = v_5896 | v_26171;
assign v_26173 = v_5869 | ~v_5990;
assign v_26175 = v_5740 | v_26174;
assign v_26176 = v_5725 | ~v_5834;
assign v_26178 = v_5608 | v_26177;
assign v_26179 = v_5584 | ~v_5702;
assign v_26181 = v_5458 | v_26180;
assign v_26182 = v_5443 | ~v_5552;
assign v_26184 = v_5326 | v_26183;
assign v_26185 = v_5287 | v_5420;
assign v_26187 = v_5146 | v_26186;
assign v_26188 = v_5131 | v_5240;
assign v_26190 = v_5014 | v_26189;
assign v_26191 = v_4987 | ~v_5108;
assign v_26193 = v_4858 | v_26192;
assign v_26194 = v_4843 | ~v_4952;
assign v_26196 = v_4726 | v_26195;
assign v_26197 = v_4699 | ~v_4820;
assign v_26199 = v_4570 | v_26198;
assign v_26200 = v_4555 | ~v_4664;
assign v_26202 = v_4438 | v_26201;
assign v_26203 = v_4414 | ~v_4532;
assign v_26205 = v_4288 | v_26204;
assign v_26206 = v_4273 | ~v_4382;
assign v_26208 = v_4156 | v_26207;
assign v_26209 = v_4125 | v_4250;
assign v_26211 = v_3992 | v_26210;
assign v_26212 = v_3977 | v_4086;
assign v_26214 = v_3860 | v_26213;
assign v_26215 = v_3835 | v_3954;
assign v_26217 = v_3708 | v_26216;
assign v_26218 = v_3693 | v_3802;
assign v_26220 = v_3576 | v_26219;
assign v_26221 = v_3549 | v_3670;
assign v_26223 = v_3420 | v_26222;
assign v_26224 = v_3405 | ~v_3514;
assign v_26226 = v_3288 | v_26225;
assign v_26227 = v_3264 | v_3382;
assign v_26229 = v_3138 | v_26228;
assign v_26230 = v_3123 | ~v_3232;
assign v_26232 = v_3006 | v_26231;
assign v_26233 = v_2971 | v_3100;
assign v_26235 = v_2834 | v_26234;
assign v_26236 = v_2819 | v_2928;
assign v_26238 = v_2702 | v_26237;
assign v_26239 = v_2676 | v_2796;
assign v_26241 = v_2548 | v_26240;
assign v_26242 = v_2533 | v_2642;
assign v_26244 = v_2416 | v_26243;
assign v_26245 = v_2389 | v_2510;
assign v_26247 = v_2260 | v_26246;
assign v_26248 = v_2245 | ~v_2354;
assign v_26250 = v_2128 | v_26249;
assign v_26251 = v_2104 | ~v_2222;
assign v_26253 = v_1978 | v_26252;
assign v_26254 = v_1963 | ~v_2072;
assign v_26256 = v_1846 | v_26255;
assign v_26257 = v_1815 | v_1940;
assign v_26259 = v_1682 | v_26258;
assign v_26260 = v_1667 | v_1776;
assign v_26262 = v_1550 | v_26261;
assign v_26263 = v_1525 | v_1644;
assign v_26265 = v_1398 | v_26264;
assign v_26266 = v_1383 | v_1492;
assign v_26268 = v_1266 | v_26267;
assign v_26269 = v_1239 | v_1360;
assign v_26271 = v_1110 | v_26270;
assign v_26272 = v_1095 | v_1204;
assign v_26274 = v_978 | v_26273;
assign v_26275 = v_954 | v_1072;
assign v_26277 = v_832 | v_26276;
assign v_26278 = v_816 | v_922;
assign v_26280 = v_715 | v_26279;
assign v_26281 = v_561 | v_793;
assign v_26294 = ~v_563 | v_26293;
assign v_26295 = v_9637 | ~v_9784;
assign v_26296 = v_9609 | ~v_9652;
assign v_26298 = v_9482 | v_26297;
assign v_26299 = v_9467 | ~v_9494;
assign v_26301 = v_9344 | v_26300;
assign v_26302 = v_9317 | ~v_9362;
assign v_26304 = v_9194 | v_26303;
assign v_26305 = v_9179 | ~v_9206;
assign v_26307 = v_9059 | v_26306;
assign v_26308 = v_9035 | ~v_9074;
assign v_26310 = v_8912 | v_26309;
assign v_26311 = v_8897 | ~v_8924;
assign v_26313 = v_8771 | v_26312;
assign v_26314 = v_8740 | ~v_8792;
assign v_26316 = v_8616 | v_26315;
assign v_26317 = v_8601 | ~v_8628;
assign v_26319 = v_8481 | v_26318;
assign v_26320 = v_8456 | ~v_8496;
assign v_26322 = v_8332 | v_26321;
assign v_26323 = v_8317 | ~v_8344;
assign v_26325 = v_8194 | v_26324;
assign v_26326 = v_8167 | ~v_8212;
assign v_26328 = v_8044 | v_26327;
assign v_26329 = v_8029 | ~v_8056;
assign v_26331 = v_7909 | v_26330;
assign v_26332 = v_7885 | ~v_7924;
assign v_26334 = v_7762 | v_26333;
assign v_26335 = v_7747 | ~v_7774;
assign v_26337 = v_7618 | v_26336;
assign v_26338 = v_7583 | ~v_7642;
assign v_26340 = v_7458 | v_26339;
assign v_26341 = v_7443 | ~v_7470;
assign v_26343 = v_7323 | v_26342;
assign v_26344 = v_7297 | ~v_7338;
assign v_26346 = v_7172 | v_26345;
assign v_26347 = v_7157 | ~v_7184;
assign v_26349 = v_7034 | v_26348;
assign v_26350 = v_7007 | ~v_7052;
assign v_26352 = v_6884 | v_26351;
assign v_26353 = v_6869 | ~v_6896;
assign v_26355 = v_6749 | v_26354;
assign v_26356 = v_6725 | ~v_6764;
assign v_26358 = v_6602 | v_26357;
assign v_26359 = v_6587 | ~v_6614;
assign v_26361 = v_6461 | v_26360;
assign v_26362 = v_6430 | ~v_6482;
assign v_26364 = v_6306 | v_26363;
assign v_26365 = v_6291 | ~v_6318;
assign v_26367 = v_6171 | v_26366;
assign v_26368 = v_6146 | ~v_6186;
assign v_26370 = v_6022 | v_26369;
assign v_26371 = v_6007 | ~v_6034;
assign v_26373 = v_5884 | v_26372;
assign v_26374 = v_5857 | ~v_5902;
assign v_26376 = v_5734 | v_26375;
assign v_26377 = v_5719 | ~v_5746;
assign v_26379 = v_5599 | v_26378;
assign v_26380 = v_5575 | ~v_5614;
assign v_26382 = v_5452 | v_26381;
assign v_26383 = v_5437 | ~v_5464;
assign v_26385 = v_5305 | v_26384;
assign v_26386 = v_5266 | ~v_5332;
assign v_26388 = v_5140 | v_26387;
assign v_26389 = v_5125 | ~v_5152;
assign v_26391 = v_5005 | v_26390;
assign v_26392 = v_4978 | ~v_5020;
assign v_26394 = v_4852 | v_26393;
assign v_26395 = v_4837 | ~v_4864;
assign v_26397 = v_4714 | v_26396;
assign v_26398 = v_4687 | ~v_4732;
assign v_26400 = v_4564 | v_26399;
assign v_26401 = v_4549 | ~v_4576;
assign v_26403 = v_4429 | v_26402;
assign v_26404 = v_4405 | ~v_4444;
assign v_26406 = v_4282 | v_26405;
assign v_26407 = v_4267 | ~v_4294;
assign v_26409 = v_4141 | v_26408;
assign v_26410 = v_4110 | ~v_4162;
assign v_26412 = v_3986 | v_26411;
assign v_26413 = v_3971 | ~v_3998;
assign v_26415 = v_3851 | v_26414;
assign v_26416 = v_3826 | ~v_3866;
assign v_26418 = v_3702 | v_26417;
assign v_26419 = v_3687 | ~v_3714;
assign v_26421 = v_3564 | v_26420;
assign v_26422 = v_3537 | ~v_3582;
assign v_26424 = v_3414 | v_26423;
assign v_26425 = v_3399 | ~v_3426;
assign v_26427 = v_3279 | v_26426;
assign v_26428 = v_3255 | ~v_3294;
assign v_26430 = v_3132 | v_26429;
assign v_26431 = v_3117 | ~v_3144;
assign v_26433 = v_2988 | v_26432;
assign v_26434 = v_2953 | ~v_3012;
assign v_26436 = v_2828 | v_26435;
assign v_26437 = v_2813 | ~v_2840;
assign v_26439 = v_2693 | v_26438;
assign v_26440 = v_2667 | ~v_2708;
assign v_26442 = v_2542 | v_26441;
assign v_26443 = v_2527 | ~v_2554;
assign v_26445 = v_2404 | v_26444;
assign v_26446 = v_2377 | ~v_2422;
assign v_26448 = v_2254 | v_26447;
assign v_26449 = v_2239 | ~v_2266;
assign v_26451 = v_2119 | v_26450;
assign v_26452 = v_2095 | ~v_2134;
assign v_26454 = v_1972 | v_26453;
assign v_26455 = v_1957 | ~v_1984;
assign v_26457 = v_1831 | v_26456;
assign v_26458 = v_1800 | ~v_1852;
assign v_26460 = v_1676 | v_26459;
assign v_26461 = v_1661 | ~v_1688;
assign v_26463 = v_1541 | v_26462;
assign v_26464 = v_1516 | ~v_1556;
assign v_26466 = v_1392 | v_26465;
assign v_26467 = v_1377 | ~v_1404;
assign v_26469 = v_1254 | v_26468;
assign v_26470 = v_1227 | ~v_1272;
assign v_26472 = v_1104 | v_26471;
assign v_26473 = v_1089 | ~v_1116;
assign v_26475 = v_969 | v_26474;
assign v_26476 = v_945 | ~v_984;
assign v_26478 = v_826 | v_26477;
assign v_26479 = v_810 | ~v_838;
assign v_26481 = v_626 | v_26480;
assign v_26482 = v_223 | ~v_721;
assign v_26484 = v_9637 | ~v_9753;
assign v_26485 = ~v_9604 | v_9609;
assign v_26487 = v_9482 | v_26486;
assign v_26488 = ~v_9463 | v_9467;
assign v_26490 = v_9344 | v_26489;
assign v_26491 = ~v_9311 | v_9317;
assign v_26493 = v_9194 | v_26492;
assign v_26494 = ~v_9175 | v_9179;
assign v_26496 = v_9059 | v_26495;
assign v_26497 = ~v_9030 | v_9035;
assign v_26499 = v_8912 | v_26498;
assign v_26500 = ~v_8893 | v_8897;
assign v_26502 = v_8771 | v_26501;
assign v_26503 = ~v_8733 | v_8740;
assign v_26505 = v_8616 | v_26504;
assign v_26506 = ~v_8597 | v_8601;
assign v_26508 = v_8481 | v_26507;
assign v_26509 = ~v_8451 | v_8456;
assign v_26511 = v_8332 | v_26510;
assign v_26512 = ~v_8313 | v_8317;
assign v_26514 = v_8194 | v_26513;
assign v_26515 = ~v_8161 | v_8167;
assign v_26517 = v_8044 | v_26516;
assign v_26518 = ~v_8025 | v_8029;
assign v_26520 = v_7909 | v_26519;
assign v_26521 = ~v_7880 | v_7885;
assign v_26523 = v_7762 | v_26522;
assign v_26524 = ~v_7743 | v_7747;
assign v_26526 = v_7618 | v_26525;
assign v_26527 = ~v_7575 | v_7583;
assign v_26529 = v_7458 | v_26528;
assign v_26530 = ~v_7439 | v_7443;
assign v_26532 = v_7323 | v_26531;
assign v_26533 = ~v_7292 | v_7297;
assign v_26535 = v_7172 | v_26534;
assign v_26536 = ~v_7153 | v_7157;
assign v_26538 = v_7034 | v_26537;
assign v_26539 = ~v_7001 | v_7007;
assign v_26541 = v_6884 | v_26540;
assign v_26542 = ~v_6865 | v_6869;
assign v_26544 = v_6749 | v_26543;
assign v_26545 = ~v_6720 | v_6725;
assign v_26547 = v_6602 | v_26546;
assign v_26548 = ~v_6583 | v_6587;
assign v_26550 = v_6461 | v_26549;
assign v_26551 = ~v_6423 | v_6430;
assign v_26553 = v_6306 | v_26552;
assign v_26554 = ~v_6287 | v_6291;
assign v_26556 = v_6171 | v_26555;
assign v_26557 = ~v_6141 | v_6146;
assign v_26559 = v_6022 | v_26558;
assign v_26560 = ~v_6003 | v_6007;
assign v_26562 = v_5884 | v_26561;
assign v_26563 = ~v_5851 | v_5857;
assign v_26565 = v_5734 | v_26564;
assign v_26566 = ~v_5715 | v_5719;
assign v_26568 = v_5599 | v_26567;
assign v_26569 = ~v_5570 | v_5575;
assign v_26571 = v_5452 | v_26570;
assign v_26572 = ~v_5433 | v_5437;
assign v_26574 = v_5305 | v_26573;
assign v_26575 = ~v_5257 | v_5266;
assign v_26577 = v_5140 | v_26576;
assign v_26578 = ~v_5121 | v_5125;
assign v_26580 = v_5005 | v_26579;
assign v_26581 = ~v_4973 | v_4978;
assign v_26583 = v_4852 | v_26582;
assign v_26584 = ~v_4833 | v_4837;
assign v_26586 = v_4714 | v_26585;
assign v_26587 = ~v_4681 | v_4687;
assign v_26589 = v_4564 | v_26588;
assign v_26590 = ~v_4545 | v_4549;
assign v_26592 = v_4429 | v_26591;
assign v_26593 = ~v_4400 | v_4405;
assign v_26595 = v_4282 | v_26594;
assign v_26596 = ~v_4263 | v_4267;
assign v_26598 = v_4141 | v_26597;
assign v_26599 = ~v_4103 | v_4110;
assign v_26601 = v_3986 | v_26600;
assign v_26602 = ~v_3967 | v_3971;
assign v_26604 = v_3851 | v_26603;
assign v_26605 = ~v_3821 | v_3826;
assign v_26607 = v_3702 | v_26606;
assign v_26608 = ~v_3683 | v_3687;
assign v_26610 = v_3564 | v_26609;
assign v_26611 = ~v_3531 | v_3537;
assign v_26613 = v_3414 | v_26612;
assign v_26614 = ~v_3395 | v_3399;
assign v_26616 = v_3279 | v_26615;
assign v_26617 = ~v_3250 | v_3255;
assign v_26619 = v_3132 | v_26618;
assign v_26620 = ~v_3113 | v_3117;
assign v_26622 = v_2988 | v_26621;
assign v_26623 = ~v_2945 | v_2953;
assign v_26625 = v_2828 | v_26624;
assign v_26626 = ~v_2809 | v_2813;
assign v_26628 = v_2693 | v_26627;
assign v_26629 = ~v_2662 | v_2667;
assign v_26631 = v_2542 | v_26630;
assign v_26632 = ~v_2523 | v_2527;
assign v_26634 = v_2404 | v_26633;
assign v_26635 = ~v_2371 | v_2377;
assign v_26637 = v_2254 | v_26636;
assign v_26638 = ~v_2235 | v_2239;
assign v_26640 = v_2119 | v_26639;
assign v_26641 = ~v_2090 | v_2095;
assign v_26643 = v_1972 | v_26642;
assign v_26644 = ~v_1953 | v_1957;
assign v_26646 = v_1831 | v_26645;
assign v_26647 = ~v_1793 | v_1800;
assign v_26649 = v_1676 | v_26648;
assign v_26650 = ~v_1657 | v_1661;
assign v_26652 = v_1541 | v_26651;
assign v_26653 = ~v_1511 | v_1516;
assign v_26655 = v_1392 | v_26654;
assign v_26656 = ~v_1373 | v_1377;
assign v_26658 = v_1254 | v_26657;
assign v_26659 = ~v_1221 | v_1227;
assign v_26661 = v_1104 | v_26660;
assign v_26662 = ~v_1085 | v_1089;
assign v_26664 = v_969 | v_26663;
assign v_26665 = ~v_940 | v_945;
assign v_26667 = v_826 | v_26666;
assign v_26668 = ~v_804 | v_810;
assign v_26670 = v_626 | v_26669;
assign v_26671 = ~v_98 | v_223;
assign v_26674 = v_9637 | ~v_9796;
assign v_26675 = v_9609 | ~v_9664;
assign v_26677 = v_9482 | v_26676;
assign v_26678 = v_9467 | ~v_9506;
assign v_26680 = v_9344 | v_26679;
assign v_26681 = v_9317 | ~v_9374;
assign v_26683 = v_9194 | v_26682;
assign v_26684 = v_9179 | ~v_9218;
assign v_26686 = v_9059 | v_26685;
assign v_26687 = v_9035 | ~v_9086;
assign v_26689 = v_8912 | v_26688;
assign v_26690 = v_8897 | ~v_8936;
assign v_26692 = v_8771 | v_26691;
assign v_26693 = v_8740 | ~v_8804;
assign v_26695 = v_8616 | v_26694;
assign v_26696 = v_8601 | ~v_8640;
assign v_26698 = v_8481 | v_26697;
assign v_26699 = v_8456 | ~v_8508;
assign v_26701 = v_8332 | v_26700;
assign v_26702 = v_8317 | ~v_8356;
assign v_26704 = v_8194 | v_26703;
assign v_26705 = v_8167 | ~v_8224;
assign v_26707 = v_8044 | v_26706;
assign v_26708 = v_8029 | ~v_8068;
assign v_26710 = v_7909 | v_26709;
assign v_26711 = v_7885 | ~v_7936;
assign v_26713 = v_7762 | v_26712;
assign v_26714 = v_7747 | ~v_7786;
assign v_26716 = v_7618 | v_26715;
assign v_26717 = v_7583 | ~v_7654;
assign v_26719 = v_7458 | v_26718;
assign v_26720 = v_7443 | ~v_7482;
assign v_26722 = v_7323 | v_26721;
assign v_26723 = v_7297 | ~v_7350;
assign v_26725 = v_7172 | v_26724;
assign v_26726 = v_7157 | ~v_7196;
assign v_26728 = v_7034 | v_26727;
assign v_26729 = v_7007 | ~v_7064;
assign v_26731 = v_6884 | v_26730;
assign v_26732 = v_6869 | ~v_6908;
assign v_26734 = v_6749 | v_26733;
assign v_26735 = v_6725 | ~v_6776;
assign v_26737 = v_6602 | v_26736;
assign v_26738 = v_6587 | ~v_6626;
assign v_26740 = v_6461 | v_26739;
assign v_26741 = v_6430 | ~v_6494;
assign v_26743 = v_6306 | v_26742;
assign v_26744 = v_6291 | ~v_6330;
assign v_26746 = v_6171 | v_26745;
assign v_26747 = v_6146 | ~v_6198;
assign v_26749 = v_6022 | v_26748;
assign v_26750 = v_6007 | ~v_6046;
assign v_26752 = v_5884 | v_26751;
assign v_26753 = v_5857 | ~v_5914;
assign v_26755 = v_5734 | v_26754;
assign v_26756 = v_5719 | ~v_5758;
assign v_26758 = v_5599 | v_26757;
assign v_26759 = v_5575 | ~v_5626;
assign v_26761 = v_5452 | v_26760;
assign v_26762 = v_5437 | ~v_5476;
assign v_26764 = v_5305 | v_26763;
assign v_26765 = v_5266 | ~v_5344;
assign v_26767 = v_5140 | v_26766;
assign v_26768 = v_5125 | ~v_5164;
assign v_26770 = v_5005 | v_26769;
assign v_26771 = v_4978 | ~v_5032;
assign v_26773 = v_4852 | v_26772;
assign v_26774 = v_4837 | ~v_4876;
assign v_26776 = v_4714 | v_26775;
assign v_26777 = v_4687 | ~v_4744;
assign v_26779 = v_4564 | v_26778;
assign v_26780 = v_4549 | ~v_4588;
assign v_26782 = v_4429 | v_26781;
assign v_26783 = v_4405 | ~v_4456;
assign v_26785 = v_4282 | v_26784;
assign v_26786 = v_4267 | ~v_4306;
assign v_26788 = v_4141 | v_26787;
assign v_26789 = v_4110 | ~v_4174;
assign v_26791 = v_3986 | v_26790;
assign v_26792 = v_3971 | ~v_4010;
assign v_26794 = v_3851 | v_26793;
assign v_26795 = v_3826 | ~v_3878;
assign v_26797 = v_3702 | v_26796;
assign v_26798 = v_3687 | ~v_3726;
assign v_26800 = v_3564 | v_26799;
assign v_26801 = v_3537 | ~v_3594;
assign v_26803 = v_3414 | v_26802;
assign v_26804 = v_3399 | ~v_3438;
assign v_26806 = v_3279 | v_26805;
assign v_26807 = v_3255 | ~v_3306;
assign v_26809 = v_3132 | v_26808;
assign v_26810 = v_3117 | ~v_3156;
assign v_26812 = v_2988 | v_26811;
assign v_26813 = v_2953 | ~v_3024;
assign v_26815 = v_2828 | v_26814;
assign v_26816 = v_2813 | ~v_2852;
assign v_26818 = v_2693 | v_26817;
assign v_26819 = v_2667 | ~v_2720;
assign v_26821 = v_2542 | v_26820;
assign v_26822 = v_2527 | ~v_2566;
assign v_26824 = v_2404 | v_26823;
assign v_26825 = v_2377 | ~v_2434;
assign v_26827 = v_2254 | v_26826;
assign v_26828 = v_2239 | ~v_2278;
assign v_26830 = v_2119 | v_26829;
assign v_26831 = v_2095 | ~v_2146;
assign v_26833 = v_1972 | v_26832;
assign v_26834 = v_1957 | ~v_1996;
assign v_26836 = v_1831 | v_26835;
assign v_26837 = v_1800 | ~v_1864;
assign v_26839 = v_1676 | v_26838;
assign v_26840 = v_1661 | ~v_1700;
assign v_26842 = v_1541 | v_26841;
assign v_26843 = v_1516 | ~v_1568;
assign v_26845 = v_1392 | v_26844;
assign v_26846 = v_1377 | ~v_1416;
assign v_26848 = v_1254 | v_26847;
assign v_26849 = v_1227 | ~v_1284;
assign v_26851 = v_1104 | v_26850;
assign v_26852 = v_1089 | ~v_1128;
assign v_26854 = v_969 | v_26853;
assign v_26855 = v_945 | ~v_996;
assign v_26857 = v_826 | v_26856;
assign v_26858 = v_810 | ~v_850;
assign v_26860 = v_626 | v_26859;
assign v_26861 = v_223 | ~v_731;
assign v_26864 = v_9637 | ~v_9808;
assign v_26865 = v_9609 | ~v_9676;
assign v_26867 = v_9482 | v_26866;
assign v_26868 = v_9467 | ~v_9518;
assign v_26870 = v_9344 | v_26869;
assign v_26871 = v_9317 | ~v_9386;
assign v_26873 = v_9194 | v_26872;
assign v_26874 = v_9179 | ~v_9230;
assign v_26876 = v_9059 | v_26875;
assign v_26877 = v_9035 | ~v_9098;
assign v_26879 = v_8912 | v_26878;
assign v_26880 = v_8897 | ~v_8948;
assign v_26882 = v_8771 | v_26881;
assign v_26883 = v_8740 | ~v_8816;
assign v_26885 = v_8616 | v_26884;
assign v_26886 = v_8601 | ~v_8652;
assign v_26888 = v_8481 | v_26887;
assign v_26889 = v_8456 | ~v_8520;
assign v_26891 = v_8332 | v_26890;
assign v_26892 = v_8317 | ~v_8368;
assign v_26894 = v_8194 | v_26893;
assign v_26895 = v_8167 | ~v_8236;
assign v_26897 = v_8044 | v_26896;
assign v_26898 = v_8029 | ~v_8080;
assign v_26900 = v_7909 | v_26899;
assign v_26901 = v_7885 | ~v_7948;
assign v_26903 = v_7762 | v_26902;
assign v_26904 = v_7747 | ~v_7798;
assign v_26906 = v_7618 | v_26905;
assign v_26907 = v_7583 | ~v_7666;
assign v_26909 = v_7458 | v_26908;
assign v_26910 = v_7443 | ~v_7494;
assign v_26912 = v_7323 | v_26911;
assign v_26913 = v_7297 | ~v_7362;
assign v_26915 = v_7172 | v_26914;
assign v_26916 = v_7157 | ~v_7208;
assign v_26918 = v_7034 | v_26917;
assign v_26919 = v_7007 | ~v_7076;
assign v_26921 = v_6884 | v_26920;
assign v_26922 = v_6869 | ~v_6920;
assign v_26924 = v_6749 | v_26923;
assign v_26925 = v_6725 | ~v_6788;
assign v_26927 = v_6602 | v_26926;
assign v_26928 = v_6587 | ~v_6638;
assign v_26930 = v_6461 | v_26929;
assign v_26931 = v_6430 | ~v_6506;
assign v_26933 = v_6306 | v_26932;
assign v_26934 = v_6291 | ~v_6342;
assign v_26936 = v_6171 | v_26935;
assign v_26937 = v_6146 | ~v_6210;
assign v_26939 = v_6022 | v_26938;
assign v_26940 = v_6007 | ~v_6058;
assign v_26942 = v_5884 | v_26941;
assign v_26943 = v_5857 | ~v_5926;
assign v_26945 = v_5734 | v_26944;
assign v_26946 = v_5719 | ~v_5770;
assign v_26948 = v_5599 | v_26947;
assign v_26949 = v_5575 | ~v_5638;
assign v_26951 = v_5452 | v_26950;
assign v_26952 = v_5437 | ~v_5488;
assign v_26954 = v_5305 | v_26953;
assign v_26955 = v_5266 | ~v_5356;
assign v_26957 = v_5140 | v_26956;
assign v_26958 = v_5125 | ~v_5176;
assign v_26960 = v_5005 | v_26959;
assign v_26961 = v_4978 | ~v_5044;
assign v_26963 = v_4852 | v_26962;
assign v_26964 = v_4837 | ~v_4888;
assign v_26966 = v_4714 | v_26965;
assign v_26967 = v_4687 | ~v_4756;
assign v_26969 = v_4564 | v_26968;
assign v_26970 = v_4549 | ~v_4600;
assign v_26972 = v_4429 | v_26971;
assign v_26973 = v_4405 | ~v_4468;
assign v_26975 = v_4282 | v_26974;
assign v_26976 = v_4267 | ~v_4318;
assign v_26978 = v_4141 | v_26977;
assign v_26979 = v_4110 | ~v_4186;
assign v_26981 = v_3986 | v_26980;
assign v_26982 = v_3971 | ~v_4022;
assign v_26984 = v_3851 | v_26983;
assign v_26985 = v_3826 | ~v_3890;
assign v_26987 = v_3702 | v_26986;
assign v_26988 = v_3687 | ~v_3738;
assign v_26990 = v_3564 | v_26989;
assign v_26991 = v_3537 | ~v_3606;
assign v_26993 = v_3414 | v_26992;
assign v_26994 = v_3399 | ~v_3450;
assign v_26996 = v_3279 | v_26995;
assign v_26997 = v_3255 | ~v_3318;
assign v_26999 = v_3132 | v_26998;
assign v_27000 = v_3117 | ~v_3168;
assign v_27002 = v_2988 | v_27001;
assign v_27003 = v_2953 | ~v_3036;
assign v_27005 = v_2828 | v_27004;
assign v_27006 = v_2813 | ~v_2864;
assign v_27008 = v_2693 | v_27007;
assign v_27009 = v_2667 | ~v_2732;
assign v_27011 = v_2542 | v_27010;
assign v_27012 = v_2527 | ~v_2578;
assign v_27014 = v_2404 | v_27013;
assign v_27015 = v_2377 | ~v_2446;
assign v_27017 = v_2254 | v_27016;
assign v_27018 = v_2239 | ~v_2290;
assign v_27020 = v_2119 | v_27019;
assign v_27021 = v_2095 | ~v_2158;
assign v_27023 = v_1972 | v_27022;
assign v_27024 = v_1957 | ~v_2008;
assign v_27026 = v_1831 | v_27025;
assign v_27027 = v_1800 | ~v_1876;
assign v_27029 = v_1676 | v_27028;
assign v_27030 = v_1661 | ~v_1712;
assign v_27032 = v_1541 | v_27031;
assign v_27033 = v_1516 | ~v_1580;
assign v_27035 = v_1392 | v_27034;
assign v_27036 = v_1377 | ~v_1428;
assign v_27038 = v_1254 | v_27037;
assign v_27039 = v_1227 | ~v_1296;
assign v_27041 = v_1104 | v_27040;
assign v_27042 = v_1089 | ~v_1140;
assign v_27044 = v_969 | v_27043;
assign v_27045 = v_945 | ~v_1008;
assign v_27047 = v_826 | v_27046;
assign v_27048 = v_810 | ~v_862;
assign v_27050 = v_626 | v_27049;
assign v_27051 = v_223 | ~v_741;
assign v_27054 = v_9637 | ~v_9820;
assign v_27055 = v_9609 | ~v_9688;
assign v_27057 = v_9482 | v_27056;
assign v_27058 = v_9467 | ~v_9530;
assign v_27060 = v_9344 | v_27059;
assign v_27061 = v_9317 | ~v_9398;
assign v_27063 = v_9194 | v_27062;
assign v_27064 = v_9179 | ~v_9242;
assign v_27066 = v_9059 | v_27065;
assign v_27067 = v_9035 | ~v_9110;
assign v_27069 = v_8912 | v_27068;
assign v_27070 = v_8897 | ~v_8960;
assign v_27072 = v_8771 | v_27071;
assign v_27073 = v_8740 | ~v_8828;
assign v_27075 = v_8616 | v_27074;
assign v_27076 = v_8601 | ~v_8664;
assign v_27078 = v_8481 | v_27077;
assign v_27079 = v_8456 | ~v_8532;
assign v_27081 = v_8332 | v_27080;
assign v_27082 = v_8317 | ~v_8380;
assign v_27084 = v_8194 | v_27083;
assign v_27085 = v_8167 | ~v_8248;
assign v_27087 = v_8044 | v_27086;
assign v_27088 = v_8029 | ~v_8092;
assign v_27090 = v_7909 | v_27089;
assign v_27091 = v_7885 | ~v_7960;
assign v_27093 = v_7762 | v_27092;
assign v_27094 = v_7747 | ~v_7810;
assign v_27096 = v_7618 | v_27095;
assign v_27097 = v_7583 | ~v_7678;
assign v_27099 = v_7458 | v_27098;
assign v_27100 = v_7443 | ~v_7506;
assign v_27102 = v_7323 | v_27101;
assign v_27103 = v_7297 | ~v_7374;
assign v_27105 = v_7172 | v_27104;
assign v_27106 = v_7157 | ~v_7220;
assign v_27108 = v_7034 | v_27107;
assign v_27109 = v_7007 | ~v_7088;
assign v_27111 = v_6884 | v_27110;
assign v_27112 = v_6869 | ~v_6932;
assign v_27114 = v_6749 | v_27113;
assign v_27115 = v_6725 | ~v_6800;
assign v_27117 = v_6602 | v_27116;
assign v_27118 = v_6587 | ~v_6650;
assign v_27120 = v_6461 | v_27119;
assign v_27121 = v_6430 | ~v_6518;
assign v_27123 = v_6306 | v_27122;
assign v_27124 = v_6291 | ~v_6354;
assign v_27126 = v_6171 | v_27125;
assign v_27127 = v_6146 | ~v_6222;
assign v_27129 = v_6022 | v_27128;
assign v_27130 = v_6007 | ~v_6070;
assign v_27132 = v_5884 | v_27131;
assign v_27133 = v_5857 | ~v_5938;
assign v_27135 = v_5734 | v_27134;
assign v_27136 = v_5719 | ~v_5782;
assign v_27138 = v_5599 | v_27137;
assign v_27139 = v_5575 | ~v_5650;
assign v_27141 = v_5452 | v_27140;
assign v_27142 = v_5437 | ~v_5500;
assign v_27144 = v_5305 | v_27143;
assign v_27145 = v_5266 | ~v_5368;
assign v_27147 = v_5140 | v_27146;
assign v_27148 = v_5125 | ~v_5188;
assign v_27150 = v_5005 | v_27149;
assign v_27151 = v_4978 | ~v_5056;
assign v_27153 = v_4852 | v_27152;
assign v_27154 = v_4837 | ~v_4900;
assign v_27156 = v_4714 | v_27155;
assign v_27157 = v_4687 | ~v_4768;
assign v_27159 = v_4564 | v_27158;
assign v_27160 = v_4549 | ~v_4612;
assign v_27162 = v_4429 | v_27161;
assign v_27163 = v_4405 | ~v_4480;
assign v_27165 = v_4282 | v_27164;
assign v_27166 = v_4267 | ~v_4330;
assign v_27168 = v_4141 | v_27167;
assign v_27169 = v_4110 | ~v_4198;
assign v_27171 = v_3986 | v_27170;
assign v_27172 = v_3971 | ~v_4034;
assign v_27174 = v_3851 | v_27173;
assign v_27175 = v_3826 | ~v_3902;
assign v_27177 = v_3702 | v_27176;
assign v_27178 = v_3687 | ~v_3750;
assign v_27180 = v_3564 | v_27179;
assign v_27181 = v_3537 | ~v_3618;
assign v_27183 = v_3414 | v_27182;
assign v_27184 = v_3399 | ~v_3462;
assign v_27186 = v_3279 | v_27185;
assign v_27187 = v_3255 | ~v_3330;
assign v_27189 = v_3132 | v_27188;
assign v_27190 = v_3117 | ~v_3180;
assign v_27192 = v_2988 | v_27191;
assign v_27193 = v_2953 | ~v_3048;
assign v_27195 = v_2828 | v_27194;
assign v_27196 = v_2813 | ~v_2876;
assign v_27198 = v_2693 | v_27197;
assign v_27199 = v_2667 | ~v_2744;
assign v_27201 = v_2542 | v_27200;
assign v_27202 = v_2527 | ~v_2590;
assign v_27204 = v_2404 | v_27203;
assign v_27205 = v_2377 | ~v_2458;
assign v_27207 = v_2254 | v_27206;
assign v_27208 = v_2239 | ~v_2302;
assign v_27210 = v_2119 | v_27209;
assign v_27211 = v_2095 | ~v_2170;
assign v_27213 = v_1972 | v_27212;
assign v_27214 = v_1957 | ~v_2020;
assign v_27216 = v_1831 | v_27215;
assign v_27217 = v_1800 | ~v_1888;
assign v_27219 = v_1676 | v_27218;
assign v_27220 = v_1661 | ~v_1724;
assign v_27222 = v_1541 | v_27221;
assign v_27223 = v_1516 | ~v_1592;
assign v_27225 = v_1392 | v_27224;
assign v_27226 = v_1377 | ~v_1440;
assign v_27228 = v_1254 | v_27227;
assign v_27229 = v_1227 | ~v_1308;
assign v_27231 = v_1104 | v_27230;
assign v_27232 = v_1089 | ~v_1152;
assign v_27234 = v_969 | v_27233;
assign v_27235 = v_945 | ~v_1020;
assign v_27237 = v_826 | v_27236;
assign v_27238 = v_810 | ~v_874;
assign v_27240 = v_626 | v_27239;
assign v_27241 = v_223 | ~v_751;
assign v_27244 = v_9637 | ~v_9832;
assign v_27245 = v_9609 | ~v_9700;
assign v_27247 = v_9482 | v_27246;
assign v_27248 = v_9467 | ~v_9542;
assign v_27250 = v_9344 | v_27249;
assign v_27251 = v_9317 | ~v_9410;
assign v_27253 = v_9194 | v_27252;
assign v_27254 = v_9179 | ~v_9254;
assign v_27256 = v_9059 | v_27255;
assign v_27257 = v_9035 | ~v_9122;
assign v_27259 = v_8912 | v_27258;
assign v_27260 = v_8897 | ~v_8972;
assign v_27262 = v_8771 | v_27261;
assign v_27263 = v_8740 | ~v_8840;
assign v_27265 = v_8616 | v_27264;
assign v_27266 = v_8601 | ~v_8676;
assign v_27268 = v_8481 | v_27267;
assign v_27269 = v_8456 | ~v_8544;
assign v_27271 = v_8332 | v_27270;
assign v_27272 = v_8317 | ~v_8392;
assign v_27274 = v_8194 | v_27273;
assign v_27275 = v_8167 | ~v_8260;
assign v_27277 = v_8044 | v_27276;
assign v_27278 = v_8029 | ~v_8104;
assign v_27280 = v_7909 | v_27279;
assign v_27281 = v_7885 | ~v_7972;
assign v_27283 = v_7762 | v_27282;
assign v_27284 = v_7747 | ~v_7822;
assign v_27286 = v_7618 | v_27285;
assign v_27287 = v_7583 | ~v_7690;
assign v_27289 = v_7458 | v_27288;
assign v_27290 = v_7443 | ~v_7518;
assign v_27292 = v_7323 | v_27291;
assign v_27293 = v_7297 | ~v_7386;
assign v_27295 = v_7172 | v_27294;
assign v_27296 = v_7157 | ~v_7232;
assign v_27298 = v_7034 | v_27297;
assign v_27299 = v_7007 | ~v_7100;
assign v_27301 = v_6884 | v_27300;
assign v_27302 = v_6869 | ~v_6944;
assign v_27304 = v_6749 | v_27303;
assign v_27305 = v_6725 | ~v_6812;
assign v_27307 = v_6602 | v_27306;
assign v_27308 = v_6587 | ~v_6662;
assign v_27310 = v_6461 | v_27309;
assign v_27311 = v_6430 | ~v_6530;
assign v_27313 = v_6306 | v_27312;
assign v_27314 = v_6291 | ~v_6366;
assign v_27316 = v_6171 | v_27315;
assign v_27317 = v_6146 | ~v_6234;
assign v_27319 = v_6022 | v_27318;
assign v_27320 = v_6007 | ~v_6082;
assign v_27322 = v_5884 | v_27321;
assign v_27323 = v_5857 | ~v_5950;
assign v_27325 = v_5734 | v_27324;
assign v_27326 = v_5719 | ~v_5794;
assign v_27328 = v_5599 | v_27327;
assign v_27329 = v_5575 | ~v_5662;
assign v_27331 = v_5452 | v_27330;
assign v_27332 = v_5437 | ~v_5512;
assign v_27334 = v_5305 | v_27333;
assign v_27335 = v_5266 | ~v_5380;
assign v_27337 = v_5140 | v_27336;
assign v_27338 = v_5125 | ~v_5200;
assign v_27340 = v_5005 | v_27339;
assign v_27341 = v_4978 | ~v_5068;
assign v_27343 = v_4852 | v_27342;
assign v_27344 = v_4837 | ~v_4912;
assign v_27346 = v_4714 | v_27345;
assign v_27347 = v_4687 | ~v_4780;
assign v_27349 = v_4564 | v_27348;
assign v_27350 = v_4549 | ~v_4624;
assign v_27352 = v_4429 | v_27351;
assign v_27353 = v_4405 | ~v_4492;
assign v_27355 = v_4282 | v_27354;
assign v_27356 = v_4267 | ~v_4342;
assign v_27358 = v_4141 | v_27357;
assign v_27359 = v_4110 | ~v_4210;
assign v_27361 = v_3986 | v_27360;
assign v_27362 = v_3971 | ~v_4046;
assign v_27364 = v_3851 | v_27363;
assign v_27365 = v_3826 | ~v_3914;
assign v_27367 = v_3702 | v_27366;
assign v_27368 = v_3687 | ~v_3762;
assign v_27370 = v_3564 | v_27369;
assign v_27371 = v_3537 | ~v_3630;
assign v_27373 = v_3414 | v_27372;
assign v_27374 = v_3399 | ~v_3474;
assign v_27376 = v_3279 | v_27375;
assign v_27377 = v_3255 | ~v_3342;
assign v_27379 = v_3132 | v_27378;
assign v_27380 = v_3117 | ~v_3192;
assign v_27382 = v_2988 | v_27381;
assign v_27383 = v_2953 | ~v_3060;
assign v_27385 = v_2828 | v_27384;
assign v_27386 = v_2813 | ~v_2888;
assign v_27388 = v_2693 | v_27387;
assign v_27389 = v_2667 | ~v_2756;
assign v_27391 = v_2542 | v_27390;
assign v_27392 = v_2527 | ~v_2602;
assign v_27394 = v_2404 | v_27393;
assign v_27395 = v_2377 | ~v_2470;
assign v_27397 = v_2254 | v_27396;
assign v_27398 = v_2239 | ~v_2314;
assign v_27400 = v_2119 | v_27399;
assign v_27401 = v_2095 | ~v_2182;
assign v_27403 = v_1972 | v_27402;
assign v_27404 = v_1957 | ~v_2032;
assign v_27406 = v_1831 | v_27405;
assign v_27407 = v_1800 | ~v_1900;
assign v_27409 = v_1676 | v_27408;
assign v_27410 = v_1661 | ~v_1736;
assign v_27412 = v_1541 | v_27411;
assign v_27413 = v_1516 | ~v_1604;
assign v_27415 = v_1392 | v_27414;
assign v_27416 = v_1377 | ~v_1452;
assign v_27418 = v_1254 | v_27417;
assign v_27419 = v_1227 | ~v_1320;
assign v_27421 = v_1104 | v_27420;
assign v_27422 = v_1089 | ~v_1164;
assign v_27424 = v_969 | v_27423;
assign v_27425 = v_945 | ~v_1032;
assign v_27427 = v_826 | v_27426;
assign v_27428 = v_810 | ~v_886;
assign v_27430 = v_626 | v_27429;
assign v_27431 = v_223 | ~v_761;
assign v_27434 = v_9637 | ~v_9844;
assign v_27435 = v_9609 | ~v_9712;
assign v_27437 = v_9482 | v_27436;
assign v_27438 = v_9467 | ~v_9554;
assign v_27440 = v_9344 | v_27439;
assign v_27441 = v_9317 | ~v_9422;
assign v_27443 = v_9194 | v_27442;
assign v_27444 = v_9179 | ~v_9266;
assign v_27446 = v_9059 | v_27445;
assign v_27447 = v_9035 | ~v_9134;
assign v_27449 = v_8912 | v_27448;
assign v_27450 = v_8897 | ~v_8984;
assign v_27452 = v_8771 | v_27451;
assign v_27453 = v_8740 | ~v_8852;
assign v_27455 = v_8616 | v_27454;
assign v_27456 = v_8601 | ~v_8688;
assign v_27458 = v_8481 | v_27457;
assign v_27459 = v_8456 | ~v_8556;
assign v_27461 = v_8332 | v_27460;
assign v_27462 = v_8317 | ~v_8404;
assign v_27464 = v_8194 | v_27463;
assign v_27465 = v_8167 | ~v_8272;
assign v_27467 = v_8044 | v_27466;
assign v_27468 = v_8029 | ~v_8116;
assign v_27470 = v_7909 | v_27469;
assign v_27471 = v_7885 | ~v_7984;
assign v_27473 = v_7762 | v_27472;
assign v_27474 = v_7747 | ~v_7834;
assign v_27476 = v_7618 | v_27475;
assign v_27477 = v_7583 | ~v_7702;
assign v_27479 = v_7458 | v_27478;
assign v_27480 = v_7443 | ~v_7530;
assign v_27482 = v_7323 | v_27481;
assign v_27483 = v_7297 | ~v_7398;
assign v_27485 = v_7172 | v_27484;
assign v_27486 = v_7157 | ~v_7244;
assign v_27488 = v_7034 | v_27487;
assign v_27489 = v_7007 | ~v_7112;
assign v_27491 = v_6884 | v_27490;
assign v_27492 = v_6869 | ~v_6956;
assign v_27494 = v_6749 | v_27493;
assign v_27495 = v_6725 | v_6824;
assign v_27497 = v_6602 | v_27496;
assign v_27498 = v_6587 | ~v_6674;
assign v_27500 = v_6461 | v_27499;
assign v_27501 = v_6430 | ~v_6542;
assign v_27503 = v_6306 | v_27502;
assign v_27504 = v_6291 | ~v_6378;
assign v_27506 = v_6171 | v_27505;
assign v_27507 = v_6146 | ~v_6246;
assign v_27509 = v_6022 | v_27508;
assign v_27510 = v_6007 | v_6094;
assign v_27512 = v_5884 | v_27511;
assign v_27513 = v_5857 | ~v_5962;
assign v_27515 = v_5734 | v_27514;
assign v_27516 = v_5719 | v_5806;
assign v_27518 = v_5599 | v_27517;
assign v_27519 = v_5575 | ~v_5674;
assign v_27521 = v_5452 | v_27520;
assign v_27522 = v_5437 | ~v_5524;
assign v_27524 = v_5305 | v_27523;
assign v_27525 = v_5266 | ~v_5392;
assign v_27527 = v_5140 | v_27526;
assign v_27528 = v_5125 | ~v_5212;
assign v_27530 = v_5005 | v_27529;
assign v_27531 = v_4978 | ~v_5080;
assign v_27533 = v_4852 | v_27532;
assign v_27534 = v_4837 | ~v_4924;
assign v_27536 = v_4714 | v_27535;
assign v_27537 = v_4687 | ~v_4792;
assign v_27539 = v_4564 | v_27538;
assign v_27540 = v_4549 | ~v_4636;
assign v_27542 = v_4429 | v_27541;
assign v_27543 = v_4405 | ~v_4504;
assign v_27545 = v_4282 | v_27544;
assign v_27546 = v_4267 | ~v_4354;
assign v_27548 = v_4141 | v_27547;
assign v_27549 = v_4110 | ~v_4222;
assign v_27551 = v_3986 | v_27550;
assign v_27552 = v_3971 | ~v_4058;
assign v_27554 = v_3851 | v_27553;
assign v_27555 = v_3826 | ~v_3926;
assign v_27557 = v_3702 | v_27556;
assign v_27558 = v_3687 | ~v_3774;
assign v_27560 = v_3564 | v_27559;
assign v_27561 = v_3537 | ~v_3642;
assign v_27563 = v_3414 | v_27562;
assign v_27564 = v_3399 | ~v_3486;
assign v_27566 = v_3279 | v_27565;
assign v_27567 = v_3255 | ~v_3354;
assign v_27569 = v_3132 | v_27568;
assign v_27570 = v_3117 | v_3204;
assign v_27572 = v_2988 | v_27571;
assign v_27573 = v_2953 | ~v_3072;
assign v_27575 = v_2828 | v_27574;
assign v_27576 = v_2813 | ~v_2900;
assign v_27578 = v_2693 | v_27577;
assign v_27579 = v_2667 | ~v_2768;
assign v_27581 = v_2542 | v_27580;
assign v_27582 = v_2527 | ~v_2614;
assign v_27584 = v_2404 | v_27583;
assign v_27585 = v_2377 | ~v_2482;
assign v_27587 = v_2254 | v_27586;
assign v_27588 = v_2239 | ~v_2326;
assign v_27590 = v_2119 | v_27589;
assign v_27591 = v_2095 | ~v_2194;
assign v_27593 = v_1972 | v_27592;
assign v_27594 = v_1957 | ~v_2044;
assign v_27596 = v_1831 | v_27595;
assign v_27597 = v_1800 | ~v_1912;
assign v_27599 = v_1676 | v_27598;
assign v_27600 = v_1661 | ~v_1748;
assign v_27602 = v_1541 | v_27601;
assign v_27603 = v_1516 | ~v_1616;
assign v_27605 = v_1392 | v_27604;
assign v_27606 = v_1377 | ~v_1464;
assign v_27608 = v_1254 | v_27607;
assign v_27609 = v_1227 | ~v_1332;
assign v_27611 = v_1104 | v_27610;
assign v_27612 = v_1089 | ~v_1176;
assign v_27614 = v_969 | v_27613;
assign v_27615 = v_945 | ~v_1044;
assign v_27617 = v_826 | v_27616;
assign v_27618 = v_810 | ~v_898;
assign v_27620 = v_626 | v_27619;
assign v_27621 = v_223 | ~v_771;
assign v_27624 = v_9637 | v_9872;
assign v_27625 = v_9609 | v_9740;
assign v_27627 = v_9482 | v_27626;
assign v_27628 = v_9467 | v_9582;
assign v_27630 = v_9344 | v_27629;
assign v_27631 = v_9317 | v_9450;
assign v_27633 = v_9194 | v_27632;
assign v_27634 = v_9179 | v_9294;
assign v_27636 = v_9059 | v_27635;
assign v_27637 = v_9035 | v_9162;
assign v_27639 = v_8912 | v_27638;
assign v_27640 = v_8897 | v_9012;
assign v_27642 = v_8771 | v_27641;
assign v_27643 = v_8740 | v_8880;
assign v_27645 = v_8616 | v_27644;
assign v_27646 = v_8601 | v_8716;
assign v_27648 = v_8481 | v_27647;
assign v_27649 = v_8456 | v_8584;
assign v_27651 = v_8332 | v_27650;
assign v_27652 = v_8317 | ~v_8432;
assign v_27654 = v_8194 | v_27653;
assign v_27655 = v_8167 | ~v_8300;
assign v_27657 = v_8044 | v_27656;
assign v_27658 = v_8029 | ~v_8144;
assign v_27660 = v_7909 | v_27659;
assign v_27661 = v_7885 | v_8012;
assign v_27663 = v_7762 | v_27662;
assign v_27664 = v_7747 | v_7862;
assign v_27666 = v_7618 | v_27665;
assign v_27667 = v_7583 | v_7730;
assign v_27669 = v_7458 | v_27668;
assign v_27670 = v_7443 | v_7558;
assign v_27672 = v_7323 | v_27671;
assign v_27673 = v_7297 | v_7426;
assign v_27675 = v_7172 | v_27674;
assign v_27676 = v_7157 | ~v_7272;
assign v_27678 = v_7034 | v_27677;
assign v_27679 = v_7007 | v_7140;
assign v_27681 = v_6884 | v_27680;
assign v_27682 = v_6869 | ~v_6984;
assign v_27684 = v_6749 | v_27683;
assign v_27685 = v_6725 | ~v_6852;
assign v_27687 = v_6602 | v_27686;
assign v_27688 = v_6587 | ~v_6702;
assign v_27690 = v_6461 | v_27689;
assign v_27691 = v_6430 | v_6570;
assign v_27693 = v_6306 | v_27692;
assign v_27694 = v_6291 | v_6406;
assign v_27696 = v_6171 | v_27695;
assign v_27697 = v_6146 | ~v_6274;
assign v_27699 = v_6022 | v_27698;
assign v_27700 = v_6007 | ~v_6122;
assign v_27702 = v_5884 | v_27701;
assign v_27703 = v_5857 | ~v_5990;
assign v_27705 = v_5734 | v_27704;
assign v_27706 = v_5719 | ~v_5834;
assign v_27708 = v_5599 | v_27707;
assign v_27709 = v_5575 | ~v_5702;
assign v_27711 = v_5452 | v_27710;
assign v_27712 = v_5437 | ~v_5552;
assign v_27714 = v_5305 | v_27713;
assign v_27715 = v_5266 | v_5420;
assign v_27717 = v_5140 | v_27716;
assign v_27718 = v_5125 | v_5240;
assign v_27720 = v_5005 | v_27719;
assign v_27721 = v_4978 | ~v_5108;
assign v_27723 = v_4852 | v_27722;
assign v_27724 = v_4837 | ~v_4952;
assign v_27726 = v_4714 | v_27725;
assign v_27727 = v_4687 | ~v_4820;
assign v_27729 = v_4564 | v_27728;
assign v_27730 = v_4549 | ~v_4664;
assign v_27732 = v_4429 | v_27731;
assign v_27733 = v_4405 | ~v_4532;
assign v_27735 = v_4282 | v_27734;
assign v_27736 = v_4267 | ~v_4382;
assign v_27738 = v_4141 | v_27737;
assign v_27739 = v_4110 | v_4250;
assign v_27741 = v_3986 | v_27740;
assign v_27742 = v_3971 | v_4086;
assign v_27744 = v_3851 | v_27743;
assign v_27745 = v_3826 | v_3954;
assign v_27747 = v_3702 | v_27746;
assign v_27748 = v_3687 | v_3802;
assign v_27750 = v_3564 | v_27749;
assign v_27751 = v_3537 | v_3670;
assign v_27753 = v_3414 | v_27752;
assign v_27754 = v_3399 | ~v_3514;
assign v_27756 = v_3279 | v_27755;
assign v_27757 = v_3255 | v_3382;
assign v_27759 = v_3132 | v_27758;
assign v_27760 = v_3117 | ~v_3232;
assign v_27762 = v_2988 | v_27761;
assign v_27763 = v_2953 | v_3100;
assign v_27765 = v_2828 | v_27764;
assign v_27766 = v_2813 | v_2928;
assign v_27768 = v_2693 | v_27767;
assign v_27769 = v_2667 | v_2796;
assign v_27771 = v_2542 | v_27770;
assign v_27772 = v_2527 | v_2642;
assign v_27774 = v_2404 | v_27773;
assign v_27775 = v_2377 | v_2510;
assign v_27777 = v_2254 | v_27776;
assign v_27778 = v_2239 | ~v_2354;
assign v_27780 = v_2119 | v_27779;
assign v_27781 = v_2095 | ~v_2222;
assign v_27783 = v_1972 | v_27782;
assign v_27784 = v_1957 | ~v_2072;
assign v_27786 = v_1831 | v_27785;
assign v_27787 = v_1800 | v_1940;
assign v_27789 = v_1676 | v_27788;
assign v_27790 = v_1661 | v_1776;
assign v_27792 = v_1541 | v_27791;
assign v_27793 = v_1516 | v_1644;
assign v_27795 = v_1392 | v_27794;
assign v_27796 = v_1377 | v_1492;
assign v_27798 = v_1254 | v_27797;
assign v_27799 = v_1227 | v_1360;
assign v_27801 = v_1104 | v_27800;
assign v_27802 = v_1089 | v_1204;
assign v_27804 = v_969 | v_27803;
assign v_27805 = v_945 | v_1072;
assign v_27807 = v_826 | v_27806;
assign v_27808 = v_810 | v_922;
assign v_27810 = v_626 | v_27809;
assign v_27811 = v_223 | v_793;
assign v_27814 = v_9639 | ~v_9784;
assign v_27815 = v_9611 | ~v_9652;
assign v_27817 = v_9483 | v_27816;
assign v_27818 = v_9468 | ~v_9494;
assign v_27820 = v_9347 | v_27819;
assign v_27821 = v_9320 | ~v_9362;
assign v_27823 = v_9195 | v_27822;
assign v_27824 = v_9180 | ~v_9206;
assign v_27826 = v_9061 | v_27825;
assign v_27827 = v_9037 | ~v_9074;
assign v_27829 = v_8913 | v_27828;
assign v_27830 = v_8898 | ~v_8924;
assign v_27832 = v_8775 | v_27831;
assign v_27833 = v_8744 | ~v_8792;
assign v_27835 = v_8617 | v_27834;
assign v_27836 = v_8602 | ~v_8628;
assign v_27838 = v_8483 | v_27837;
assign v_27839 = v_8458 | ~v_8496;
assign v_27841 = v_8333 | v_27840;
assign v_27842 = v_8318 | ~v_8344;
assign v_27844 = v_8197 | v_27843;
assign v_27845 = v_8170 | ~v_8212;
assign v_27847 = v_8045 | v_27846;
assign v_27848 = v_8030 | ~v_8056;
assign v_27850 = v_7911 | v_27849;
assign v_27851 = v_7887 | ~v_7924;
assign v_27853 = v_7763 | v_27852;
assign v_27854 = v_7748 | ~v_7774;
assign v_27856 = v_7623 | v_27855;
assign v_27857 = v_7588 | ~v_7642;
assign v_27859 = v_7459 | v_27858;
assign v_27860 = v_7444 | ~v_7470;
assign v_27862 = v_7325 | v_27861;
assign v_27863 = v_7299 | ~v_7338;
assign v_27865 = v_7173 | v_27864;
assign v_27866 = v_7158 | ~v_7184;
assign v_27868 = v_7037 | v_27867;
assign v_27869 = v_7010 | ~v_7052;
assign v_27871 = v_6885 | v_27870;
assign v_27872 = v_6870 | ~v_6896;
assign v_27874 = v_6751 | v_27873;
assign v_27875 = v_6727 | ~v_6764;
assign v_27877 = v_6603 | v_27876;
assign v_27878 = v_6588 | ~v_6614;
assign v_27880 = v_6465 | v_27879;
assign v_27881 = v_6434 | ~v_6482;
assign v_27883 = v_6307 | v_27882;
assign v_27884 = v_6292 | ~v_6318;
assign v_27886 = v_6173 | v_27885;
assign v_27887 = v_6148 | ~v_6186;
assign v_27889 = v_6023 | v_27888;
assign v_27890 = v_6008 | ~v_6034;
assign v_27892 = v_5887 | v_27891;
assign v_27893 = v_5860 | ~v_5902;
assign v_27895 = v_5735 | v_27894;
assign v_27896 = v_5720 | ~v_5746;
assign v_27898 = v_5601 | v_27897;
assign v_27899 = v_5577 | ~v_5614;
assign v_27901 = v_5453 | v_27900;
assign v_27902 = v_5438 | ~v_5464;
assign v_27904 = v_5311 | v_27903;
assign v_27905 = v_5272 | ~v_5332;
assign v_27907 = v_5141 | v_27906;
assign v_27908 = v_5126 | ~v_5152;
assign v_27910 = v_5007 | v_27909;
assign v_27911 = v_4980 | ~v_5020;
assign v_27913 = v_4853 | v_27912;
assign v_27914 = v_4838 | ~v_4864;
assign v_27916 = v_4717 | v_27915;
assign v_27917 = v_4690 | ~v_4732;
assign v_27919 = v_4565 | v_27918;
assign v_27920 = v_4550 | ~v_4576;
assign v_27922 = v_4431 | v_27921;
assign v_27923 = v_4407 | ~v_4444;
assign v_27925 = v_4283 | v_27924;
assign v_27926 = v_4268 | ~v_4294;
assign v_27928 = v_4145 | v_27927;
assign v_27929 = v_4114 | ~v_4162;
assign v_27931 = v_3987 | v_27930;
assign v_27932 = v_3972 | ~v_3998;
assign v_27934 = v_3853 | v_27933;
assign v_27935 = v_3828 | ~v_3866;
assign v_27937 = v_3703 | v_27936;
assign v_27938 = v_3688 | ~v_3714;
assign v_27940 = v_3567 | v_27939;
assign v_27941 = v_3540 | ~v_3582;
assign v_27943 = v_3415 | v_27942;
assign v_27944 = v_3400 | ~v_3426;
assign v_27946 = v_3281 | v_27945;
assign v_27947 = v_3257 | ~v_3294;
assign v_27949 = v_3133 | v_27948;
assign v_27950 = v_3118 | ~v_3144;
assign v_27952 = v_2993 | v_27951;
assign v_27953 = v_2958 | ~v_3012;
assign v_27955 = v_2829 | v_27954;
assign v_27956 = v_2814 | ~v_2840;
assign v_27958 = v_2695 | v_27957;
assign v_27959 = v_2669 | ~v_2708;
assign v_27961 = v_2543 | v_27960;
assign v_27962 = v_2528 | ~v_2554;
assign v_27964 = v_2407 | v_27963;
assign v_27965 = v_2380 | ~v_2422;
assign v_27967 = v_2255 | v_27966;
assign v_27968 = v_2240 | ~v_2266;
assign v_27970 = v_2121 | v_27969;
assign v_27971 = v_2097 | ~v_2134;
assign v_27973 = v_1973 | v_27972;
assign v_27974 = v_1958 | ~v_1984;
assign v_27976 = v_1835 | v_27975;
assign v_27977 = v_1804 | ~v_1852;
assign v_27979 = v_1677 | v_27978;
assign v_27980 = v_1662 | ~v_1688;
assign v_27982 = v_1543 | v_27981;
assign v_27983 = v_1518 | ~v_1556;
assign v_27985 = v_1393 | v_27984;
assign v_27986 = v_1378 | ~v_1404;
assign v_27988 = v_1257 | v_27987;
assign v_27989 = v_1230 | ~v_1272;
assign v_27991 = v_1105 | v_27990;
assign v_27992 = v_1090 | ~v_1116;
assign v_27994 = v_971 | v_27993;
assign v_27995 = v_947 | ~v_984;
assign v_27997 = v_827 | v_27996;
assign v_27998 = v_811 | ~v_838;
assign v_28000 = v_658 | v_27999;
assign v_28001 = v_359 | ~v_721;
assign v_28003 = v_9639 | ~v_9753;
assign v_28004 = ~v_9604 | v_9611;
assign v_28006 = v_9483 | v_28005;
assign v_28007 = ~v_9463 | v_9468;
assign v_28009 = v_9347 | v_28008;
assign v_28010 = ~v_9311 | v_9320;
assign v_28012 = v_9195 | v_28011;
assign v_28013 = ~v_9175 | v_9180;
assign v_28015 = v_9061 | v_28014;
assign v_28016 = ~v_9030 | v_9037;
assign v_28018 = v_8913 | v_28017;
assign v_28019 = ~v_8893 | v_8898;
assign v_28021 = v_8775 | v_28020;
assign v_28022 = ~v_8733 | v_8744;
assign v_28024 = v_8617 | v_28023;
assign v_28025 = ~v_8597 | v_8602;
assign v_28027 = v_8483 | v_28026;
assign v_28028 = ~v_8451 | v_8458;
assign v_28030 = v_8333 | v_28029;
assign v_28031 = ~v_8313 | v_8318;
assign v_28033 = v_8197 | v_28032;
assign v_28034 = ~v_8161 | v_8170;
assign v_28036 = v_8045 | v_28035;
assign v_28037 = ~v_8025 | v_8030;
assign v_28039 = v_7911 | v_28038;
assign v_28040 = ~v_7880 | v_7887;
assign v_28042 = v_7763 | v_28041;
assign v_28043 = ~v_7743 | v_7748;
assign v_28045 = v_7623 | v_28044;
assign v_28046 = ~v_7575 | v_7588;
assign v_28048 = v_7459 | v_28047;
assign v_28049 = ~v_7439 | v_7444;
assign v_28051 = v_7325 | v_28050;
assign v_28052 = ~v_7292 | v_7299;
assign v_28054 = v_7173 | v_28053;
assign v_28055 = ~v_7153 | v_7158;
assign v_28057 = v_7037 | v_28056;
assign v_28058 = ~v_7001 | v_7010;
assign v_28060 = v_6885 | v_28059;
assign v_28061 = ~v_6865 | v_6870;
assign v_28063 = v_6751 | v_28062;
assign v_28064 = ~v_6720 | v_6727;
assign v_28066 = v_6603 | v_28065;
assign v_28067 = ~v_6583 | v_6588;
assign v_28069 = v_6465 | v_28068;
assign v_28070 = ~v_6423 | v_6434;
assign v_28072 = v_6307 | v_28071;
assign v_28073 = ~v_6287 | v_6292;
assign v_28075 = v_6173 | v_28074;
assign v_28076 = ~v_6141 | v_6148;
assign v_28078 = v_6023 | v_28077;
assign v_28079 = ~v_6003 | v_6008;
assign v_28081 = v_5887 | v_28080;
assign v_28082 = ~v_5851 | v_5860;
assign v_28084 = v_5735 | v_28083;
assign v_28085 = ~v_5715 | v_5720;
assign v_28087 = v_5601 | v_28086;
assign v_28088 = ~v_5570 | v_5577;
assign v_28090 = v_5453 | v_28089;
assign v_28091 = ~v_5433 | v_5438;
assign v_28093 = v_5311 | v_28092;
assign v_28094 = ~v_5257 | v_5272;
assign v_28096 = v_5141 | v_28095;
assign v_28097 = ~v_5121 | v_5126;
assign v_28099 = v_5007 | v_28098;
assign v_28100 = ~v_4973 | v_4980;
assign v_28102 = v_4853 | v_28101;
assign v_28103 = ~v_4833 | v_4838;
assign v_28105 = v_4717 | v_28104;
assign v_28106 = ~v_4681 | v_4690;
assign v_28108 = v_4565 | v_28107;
assign v_28109 = ~v_4545 | v_4550;
assign v_28111 = v_4431 | v_28110;
assign v_28112 = ~v_4400 | v_4407;
assign v_28114 = v_4283 | v_28113;
assign v_28115 = ~v_4263 | v_4268;
assign v_28117 = v_4145 | v_28116;
assign v_28118 = ~v_4103 | v_4114;
assign v_28120 = v_3987 | v_28119;
assign v_28121 = ~v_3967 | v_3972;
assign v_28123 = v_3853 | v_28122;
assign v_28124 = ~v_3821 | v_3828;
assign v_28126 = v_3703 | v_28125;
assign v_28127 = ~v_3683 | v_3688;
assign v_28129 = v_3567 | v_28128;
assign v_28130 = ~v_3531 | v_3540;
assign v_28132 = v_3415 | v_28131;
assign v_28133 = ~v_3395 | v_3400;
assign v_28135 = v_3281 | v_28134;
assign v_28136 = ~v_3250 | v_3257;
assign v_28138 = v_3133 | v_28137;
assign v_28139 = ~v_3113 | v_3118;
assign v_28141 = v_2993 | v_28140;
assign v_28142 = ~v_2945 | v_2958;
assign v_28144 = v_2829 | v_28143;
assign v_28145 = ~v_2809 | v_2814;
assign v_28147 = v_2695 | v_28146;
assign v_28148 = ~v_2662 | v_2669;
assign v_28150 = v_2543 | v_28149;
assign v_28151 = ~v_2523 | v_2528;
assign v_28153 = v_2407 | v_28152;
assign v_28154 = ~v_2371 | v_2380;
assign v_28156 = v_2255 | v_28155;
assign v_28157 = ~v_2235 | v_2240;
assign v_28159 = v_2121 | v_28158;
assign v_28160 = ~v_2090 | v_2097;
assign v_28162 = v_1973 | v_28161;
assign v_28163 = ~v_1953 | v_1958;
assign v_28165 = v_1835 | v_28164;
assign v_28166 = ~v_1793 | v_1804;
assign v_28168 = v_1677 | v_28167;
assign v_28169 = ~v_1657 | v_1662;
assign v_28171 = v_1543 | v_28170;
assign v_28172 = ~v_1511 | v_1518;
assign v_28174 = v_1393 | v_28173;
assign v_28175 = ~v_1373 | v_1378;
assign v_28177 = v_1257 | v_28176;
assign v_28178 = ~v_1221 | v_1230;
assign v_28180 = v_1105 | v_28179;
assign v_28181 = ~v_1085 | v_1090;
assign v_28183 = v_971 | v_28182;
assign v_28184 = ~v_940 | v_947;
assign v_28186 = v_827 | v_28185;
assign v_28187 = ~v_804 | v_811;
assign v_28189 = v_658 | v_28188;
assign v_28190 = ~v_98 | v_359;
assign v_28193 = v_9639 | ~v_9796;
assign v_28194 = v_9611 | ~v_9664;
assign v_28196 = v_9483 | v_28195;
assign v_28197 = v_9468 | ~v_9506;
assign v_28199 = v_9347 | v_28198;
assign v_28200 = v_9320 | ~v_9374;
assign v_28202 = v_9195 | v_28201;
assign v_28203 = v_9180 | ~v_9218;
assign v_28205 = v_9061 | v_28204;
assign v_28206 = v_9037 | ~v_9086;
assign v_28208 = v_8913 | v_28207;
assign v_28209 = v_8898 | ~v_8936;
assign v_28211 = v_8775 | v_28210;
assign v_28212 = v_8744 | ~v_8804;
assign v_28214 = v_8617 | v_28213;
assign v_28215 = v_8602 | ~v_8640;
assign v_28217 = v_8483 | v_28216;
assign v_28218 = v_8458 | ~v_8508;
assign v_28220 = v_8333 | v_28219;
assign v_28221 = v_8318 | ~v_8356;
assign v_28223 = v_8197 | v_28222;
assign v_28224 = v_8170 | ~v_8224;
assign v_28226 = v_8045 | v_28225;
assign v_28227 = v_8030 | ~v_8068;
assign v_28229 = v_7911 | v_28228;
assign v_28230 = v_7887 | ~v_7936;
assign v_28232 = v_7763 | v_28231;
assign v_28233 = v_7748 | ~v_7786;
assign v_28235 = v_7623 | v_28234;
assign v_28236 = v_7588 | ~v_7654;
assign v_28238 = v_7459 | v_28237;
assign v_28239 = v_7444 | ~v_7482;
assign v_28241 = v_7325 | v_28240;
assign v_28242 = v_7299 | ~v_7350;
assign v_28244 = v_7173 | v_28243;
assign v_28245 = v_7158 | ~v_7196;
assign v_28247 = v_7037 | v_28246;
assign v_28248 = v_7010 | ~v_7064;
assign v_28250 = v_6885 | v_28249;
assign v_28251 = v_6870 | ~v_6908;
assign v_28253 = v_6751 | v_28252;
assign v_28254 = v_6727 | ~v_6776;
assign v_28256 = v_6603 | v_28255;
assign v_28257 = v_6588 | ~v_6626;
assign v_28259 = v_6465 | v_28258;
assign v_28260 = v_6434 | ~v_6494;
assign v_28262 = v_6307 | v_28261;
assign v_28263 = v_6292 | ~v_6330;
assign v_28265 = v_6173 | v_28264;
assign v_28266 = v_6148 | ~v_6198;
assign v_28268 = v_6023 | v_28267;
assign v_28269 = v_6008 | ~v_6046;
assign v_28271 = v_5887 | v_28270;
assign v_28272 = v_5860 | ~v_5914;
assign v_28274 = v_5735 | v_28273;
assign v_28275 = v_5720 | ~v_5758;
assign v_28277 = v_5601 | v_28276;
assign v_28278 = v_5577 | ~v_5626;
assign v_28280 = v_5453 | v_28279;
assign v_28281 = v_5438 | ~v_5476;
assign v_28283 = v_5311 | v_28282;
assign v_28284 = v_5272 | ~v_5344;
assign v_28286 = v_5141 | v_28285;
assign v_28287 = v_5126 | ~v_5164;
assign v_28289 = v_5007 | v_28288;
assign v_28290 = v_4980 | ~v_5032;
assign v_28292 = v_4853 | v_28291;
assign v_28293 = v_4838 | ~v_4876;
assign v_28295 = v_4717 | v_28294;
assign v_28296 = v_4690 | ~v_4744;
assign v_28298 = v_4565 | v_28297;
assign v_28299 = v_4550 | ~v_4588;
assign v_28301 = v_4431 | v_28300;
assign v_28302 = v_4407 | ~v_4456;
assign v_28304 = v_4283 | v_28303;
assign v_28305 = v_4268 | ~v_4306;
assign v_28307 = v_4145 | v_28306;
assign v_28308 = v_4114 | ~v_4174;
assign v_28310 = v_3987 | v_28309;
assign v_28311 = v_3972 | ~v_4010;
assign v_28313 = v_3853 | v_28312;
assign v_28314 = v_3828 | ~v_3878;
assign v_28316 = v_3703 | v_28315;
assign v_28317 = v_3688 | ~v_3726;
assign v_28319 = v_3567 | v_28318;
assign v_28320 = v_3540 | ~v_3594;
assign v_28322 = v_3415 | v_28321;
assign v_28323 = v_3400 | ~v_3438;
assign v_28325 = v_3281 | v_28324;
assign v_28326 = v_3257 | ~v_3306;
assign v_28328 = v_3133 | v_28327;
assign v_28329 = v_3118 | ~v_3156;
assign v_28331 = v_2993 | v_28330;
assign v_28332 = v_2958 | ~v_3024;
assign v_28334 = v_2829 | v_28333;
assign v_28335 = v_2814 | ~v_2852;
assign v_28337 = v_2695 | v_28336;
assign v_28338 = v_2669 | ~v_2720;
assign v_28340 = v_2543 | v_28339;
assign v_28341 = v_2528 | ~v_2566;
assign v_28343 = v_2407 | v_28342;
assign v_28344 = v_2380 | ~v_2434;
assign v_28346 = v_2255 | v_28345;
assign v_28347 = v_2240 | ~v_2278;
assign v_28349 = v_2121 | v_28348;
assign v_28350 = v_2097 | ~v_2146;
assign v_28352 = v_1973 | v_28351;
assign v_28353 = v_1958 | ~v_1996;
assign v_28355 = v_1835 | v_28354;
assign v_28356 = v_1804 | ~v_1864;
assign v_28358 = v_1677 | v_28357;
assign v_28359 = v_1662 | ~v_1700;
assign v_28361 = v_1543 | v_28360;
assign v_28362 = v_1518 | ~v_1568;
assign v_28364 = v_1393 | v_28363;
assign v_28365 = v_1378 | ~v_1416;
assign v_28367 = v_1257 | v_28366;
assign v_28368 = v_1230 | ~v_1284;
assign v_28370 = v_1105 | v_28369;
assign v_28371 = v_1090 | ~v_1128;
assign v_28373 = v_971 | v_28372;
assign v_28374 = v_947 | ~v_996;
assign v_28376 = v_827 | v_28375;
assign v_28377 = v_811 | ~v_850;
assign v_28379 = v_658 | v_28378;
assign v_28380 = v_359 | ~v_731;
assign v_28383 = v_9639 | ~v_9808;
assign v_28384 = v_9611 | ~v_9676;
assign v_28386 = v_9483 | v_28385;
assign v_28387 = v_9468 | ~v_9518;
assign v_28389 = v_9347 | v_28388;
assign v_28390 = v_9320 | ~v_9386;
assign v_28392 = v_9195 | v_28391;
assign v_28393 = v_9180 | ~v_9230;
assign v_28395 = v_9061 | v_28394;
assign v_28396 = v_9037 | ~v_9098;
assign v_28398 = v_8913 | v_28397;
assign v_28399 = v_8898 | ~v_8948;
assign v_28401 = v_8775 | v_28400;
assign v_28402 = v_8744 | ~v_8816;
assign v_28404 = v_8617 | v_28403;
assign v_28405 = v_8602 | ~v_8652;
assign v_28407 = v_8483 | v_28406;
assign v_28408 = v_8458 | ~v_8520;
assign v_28410 = v_8333 | v_28409;
assign v_28411 = v_8318 | ~v_8368;
assign v_28413 = v_8197 | v_28412;
assign v_28414 = v_8170 | ~v_8236;
assign v_28416 = v_8045 | v_28415;
assign v_28417 = v_8030 | ~v_8080;
assign v_28419 = v_7911 | v_28418;
assign v_28420 = v_7887 | ~v_7948;
assign v_28422 = v_7763 | v_28421;
assign v_28423 = v_7748 | ~v_7798;
assign v_28425 = v_7623 | v_28424;
assign v_28426 = v_7588 | ~v_7666;
assign v_28428 = v_7459 | v_28427;
assign v_28429 = v_7444 | ~v_7494;
assign v_28431 = v_7325 | v_28430;
assign v_28432 = v_7299 | ~v_7362;
assign v_28434 = v_7173 | v_28433;
assign v_28435 = v_7158 | ~v_7208;
assign v_28437 = v_7037 | v_28436;
assign v_28438 = v_7010 | ~v_7076;
assign v_28440 = v_6885 | v_28439;
assign v_28441 = v_6870 | ~v_6920;
assign v_28443 = v_6751 | v_28442;
assign v_28444 = v_6727 | ~v_6788;
assign v_28446 = v_6603 | v_28445;
assign v_28447 = v_6588 | ~v_6638;
assign v_28449 = v_6465 | v_28448;
assign v_28450 = v_6434 | ~v_6506;
assign v_28452 = v_6307 | v_28451;
assign v_28453 = v_6292 | ~v_6342;
assign v_28455 = v_6173 | v_28454;
assign v_28456 = v_6148 | ~v_6210;
assign v_28458 = v_6023 | v_28457;
assign v_28459 = v_6008 | ~v_6058;
assign v_28461 = v_5887 | v_28460;
assign v_28462 = v_5860 | ~v_5926;
assign v_28464 = v_5735 | v_28463;
assign v_28465 = v_5720 | ~v_5770;
assign v_28467 = v_5601 | v_28466;
assign v_28468 = v_5577 | ~v_5638;
assign v_28470 = v_5453 | v_28469;
assign v_28471 = v_5438 | ~v_5488;
assign v_28473 = v_5311 | v_28472;
assign v_28474 = v_5272 | ~v_5356;
assign v_28476 = v_5141 | v_28475;
assign v_28477 = v_5126 | ~v_5176;
assign v_28479 = v_5007 | v_28478;
assign v_28480 = v_4980 | ~v_5044;
assign v_28482 = v_4853 | v_28481;
assign v_28483 = v_4838 | ~v_4888;
assign v_28485 = v_4717 | v_28484;
assign v_28486 = v_4690 | ~v_4756;
assign v_28488 = v_4565 | v_28487;
assign v_28489 = v_4550 | ~v_4600;
assign v_28491 = v_4431 | v_28490;
assign v_28492 = v_4407 | ~v_4468;
assign v_28494 = v_4283 | v_28493;
assign v_28495 = v_4268 | ~v_4318;
assign v_28497 = v_4145 | v_28496;
assign v_28498 = v_4114 | ~v_4186;
assign v_28500 = v_3987 | v_28499;
assign v_28501 = v_3972 | ~v_4022;
assign v_28503 = v_3853 | v_28502;
assign v_28504 = v_3828 | ~v_3890;
assign v_28506 = v_3703 | v_28505;
assign v_28507 = v_3688 | ~v_3738;
assign v_28509 = v_3567 | v_28508;
assign v_28510 = v_3540 | ~v_3606;
assign v_28512 = v_3415 | v_28511;
assign v_28513 = v_3400 | ~v_3450;
assign v_28515 = v_3281 | v_28514;
assign v_28516 = v_3257 | ~v_3318;
assign v_28518 = v_3133 | v_28517;
assign v_28519 = v_3118 | ~v_3168;
assign v_28521 = v_2993 | v_28520;
assign v_28522 = v_2958 | ~v_3036;
assign v_28524 = v_2829 | v_28523;
assign v_28525 = v_2814 | ~v_2864;
assign v_28527 = v_2695 | v_28526;
assign v_28528 = v_2669 | ~v_2732;
assign v_28530 = v_2543 | v_28529;
assign v_28531 = v_2528 | ~v_2578;
assign v_28533 = v_2407 | v_28532;
assign v_28534 = v_2380 | ~v_2446;
assign v_28536 = v_2255 | v_28535;
assign v_28537 = v_2240 | ~v_2290;
assign v_28539 = v_2121 | v_28538;
assign v_28540 = v_2097 | ~v_2158;
assign v_28542 = v_1973 | v_28541;
assign v_28543 = v_1958 | ~v_2008;
assign v_28545 = v_1835 | v_28544;
assign v_28546 = v_1804 | ~v_1876;
assign v_28548 = v_1677 | v_28547;
assign v_28549 = v_1662 | ~v_1712;
assign v_28551 = v_1543 | v_28550;
assign v_28552 = v_1518 | ~v_1580;
assign v_28554 = v_1393 | v_28553;
assign v_28555 = v_1378 | ~v_1428;
assign v_28557 = v_1257 | v_28556;
assign v_28558 = v_1230 | ~v_1296;
assign v_28560 = v_1105 | v_28559;
assign v_28561 = v_1090 | ~v_1140;
assign v_28563 = v_971 | v_28562;
assign v_28564 = v_947 | ~v_1008;
assign v_28566 = v_827 | v_28565;
assign v_28567 = v_811 | ~v_862;
assign v_28569 = v_658 | v_28568;
assign v_28570 = v_359 | ~v_741;
assign v_28573 = v_9639 | ~v_9820;
assign v_28574 = v_9611 | ~v_9688;
assign v_28576 = v_9483 | v_28575;
assign v_28577 = v_9468 | ~v_9530;
assign v_28579 = v_9347 | v_28578;
assign v_28580 = v_9320 | ~v_9398;
assign v_28582 = v_9195 | v_28581;
assign v_28583 = v_9180 | ~v_9242;
assign v_28585 = v_9061 | v_28584;
assign v_28586 = v_9037 | ~v_9110;
assign v_28588 = v_8913 | v_28587;
assign v_28589 = v_8898 | ~v_8960;
assign v_28591 = v_8775 | v_28590;
assign v_28592 = v_8744 | ~v_8828;
assign v_28594 = v_8617 | v_28593;
assign v_28595 = v_8602 | ~v_8664;
assign v_28597 = v_8483 | v_28596;
assign v_28598 = v_8458 | ~v_8532;
assign v_28600 = v_8333 | v_28599;
assign v_28601 = v_8318 | ~v_8380;
assign v_28603 = v_8197 | v_28602;
assign v_28604 = v_8170 | ~v_8248;
assign v_28606 = v_8045 | v_28605;
assign v_28607 = v_8030 | ~v_8092;
assign v_28609 = v_7911 | v_28608;
assign v_28610 = v_7887 | ~v_7960;
assign v_28612 = v_7763 | v_28611;
assign v_28613 = v_7748 | ~v_7810;
assign v_28615 = v_7623 | v_28614;
assign v_28616 = v_7588 | ~v_7678;
assign v_28618 = v_7459 | v_28617;
assign v_28619 = v_7444 | ~v_7506;
assign v_28621 = v_7325 | v_28620;
assign v_28622 = v_7299 | ~v_7374;
assign v_28624 = v_7173 | v_28623;
assign v_28625 = v_7158 | ~v_7220;
assign v_28627 = v_7037 | v_28626;
assign v_28628 = v_7010 | ~v_7088;
assign v_28630 = v_6885 | v_28629;
assign v_28631 = v_6870 | ~v_6932;
assign v_28633 = v_6751 | v_28632;
assign v_28634 = v_6727 | ~v_6800;
assign v_28636 = v_6603 | v_28635;
assign v_28637 = v_6588 | ~v_6650;
assign v_28639 = v_6465 | v_28638;
assign v_28640 = v_6434 | ~v_6518;
assign v_28642 = v_6307 | v_28641;
assign v_28643 = v_6292 | ~v_6354;
assign v_28645 = v_6173 | v_28644;
assign v_28646 = v_6148 | ~v_6222;
assign v_28648 = v_6023 | v_28647;
assign v_28649 = v_6008 | ~v_6070;
assign v_28651 = v_5887 | v_28650;
assign v_28652 = v_5860 | ~v_5938;
assign v_28654 = v_5735 | v_28653;
assign v_28655 = v_5720 | ~v_5782;
assign v_28657 = v_5601 | v_28656;
assign v_28658 = v_5577 | ~v_5650;
assign v_28660 = v_5453 | v_28659;
assign v_28661 = v_5438 | ~v_5500;
assign v_28663 = v_5311 | v_28662;
assign v_28664 = v_5272 | ~v_5368;
assign v_28666 = v_5141 | v_28665;
assign v_28667 = v_5126 | ~v_5188;
assign v_28669 = v_5007 | v_28668;
assign v_28670 = v_4980 | ~v_5056;
assign v_28672 = v_4853 | v_28671;
assign v_28673 = v_4838 | ~v_4900;
assign v_28675 = v_4717 | v_28674;
assign v_28676 = v_4690 | ~v_4768;
assign v_28678 = v_4565 | v_28677;
assign v_28679 = v_4550 | ~v_4612;
assign v_28681 = v_4431 | v_28680;
assign v_28682 = v_4407 | ~v_4480;
assign v_28684 = v_4283 | v_28683;
assign v_28685 = v_4268 | ~v_4330;
assign v_28687 = v_4145 | v_28686;
assign v_28688 = v_4114 | ~v_4198;
assign v_28690 = v_3987 | v_28689;
assign v_28691 = v_3972 | ~v_4034;
assign v_28693 = v_3853 | v_28692;
assign v_28694 = v_3828 | ~v_3902;
assign v_28696 = v_3703 | v_28695;
assign v_28697 = v_3688 | ~v_3750;
assign v_28699 = v_3567 | v_28698;
assign v_28700 = v_3540 | ~v_3618;
assign v_28702 = v_3415 | v_28701;
assign v_28703 = v_3400 | ~v_3462;
assign v_28705 = v_3281 | v_28704;
assign v_28706 = v_3257 | ~v_3330;
assign v_28708 = v_3133 | v_28707;
assign v_28709 = v_3118 | ~v_3180;
assign v_28711 = v_2993 | v_28710;
assign v_28712 = v_2958 | ~v_3048;
assign v_28714 = v_2829 | v_28713;
assign v_28715 = v_2814 | ~v_2876;
assign v_28717 = v_2695 | v_28716;
assign v_28718 = v_2669 | ~v_2744;
assign v_28720 = v_2543 | v_28719;
assign v_28721 = v_2528 | ~v_2590;
assign v_28723 = v_2407 | v_28722;
assign v_28724 = v_2380 | ~v_2458;
assign v_28726 = v_2255 | v_28725;
assign v_28727 = v_2240 | ~v_2302;
assign v_28729 = v_2121 | v_28728;
assign v_28730 = v_2097 | ~v_2170;
assign v_28732 = v_1973 | v_28731;
assign v_28733 = v_1958 | ~v_2020;
assign v_28735 = v_1835 | v_28734;
assign v_28736 = v_1804 | ~v_1888;
assign v_28738 = v_1677 | v_28737;
assign v_28739 = v_1662 | ~v_1724;
assign v_28741 = v_1543 | v_28740;
assign v_28742 = v_1518 | ~v_1592;
assign v_28744 = v_1393 | v_28743;
assign v_28745 = v_1378 | ~v_1440;
assign v_28747 = v_1257 | v_28746;
assign v_28748 = v_1230 | ~v_1308;
assign v_28750 = v_1105 | v_28749;
assign v_28751 = v_1090 | ~v_1152;
assign v_28753 = v_971 | v_28752;
assign v_28754 = v_947 | ~v_1020;
assign v_28756 = v_827 | v_28755;
assign v_28757 = v_811 | ~v_874;
assign v_28759 = v_658 | v_28758;
assign v_28760 = v_359 | ~v_751;
assign v_28763 = v_9639 | ~v_9832;
assign v_28764 = v_9611 | ~v_9700;
assign v_28766 = v_9483 | v_28765;
assign v_28767 = v_9468 | ~v_9542;
assign v_28769 = v_9347 | v_28768;
assign v_28770 = v_9320 | ~v_9410;
assign v_28772 = v_9195 | v_28771;
assign v_28773 = v_9180 | ~v_9254;
assign v_28775 = v_9061 | v_28774;
assign v_28776 = v_9037 | ~v_9122;
assign v_28778 = v_8913 | v_28777;
assign v_28779 = v_8898 | ~v_8972;
assign v_28781 = v_8775 | v_28780;
assign v_28782 = v_8744 | ~v_8840;
assign v_28784 = v_8617 | v_28783;
assign v_28785 = v_8602 | ~v_8676;
assign v_28787 = v_8483 | v_28786;
assign v_28788 = v_8458 | ~v_8544;
assign v_28790 = v_8333 | v_28789;
assign v_28791 = v_8318 | ~v_8392;
assign v_28793 = v_8197 | v_28792;
assign v_28794 = v_8170 | ~v_8260;
assign v_28796 = v_8045 | v_28795;
assign v_28797 = v_8030 | ~v_8104;
assign v_28799 = v_7911 | v_28798;
assign v_28800 = v_7887 | ~v_7972;
assign v_28802 = v_7763 | v_28801;
assign v_28803 = v_7748 | ~v_7822;
assign v_28805 = v_7623 | v_28804;
assign v_28806 = v_7588 | ~v_7690;
assign v_28808 = v_7459 | v_28807;
assign v_28809 = v_7444 | ~v_7518;
assign v_28811 = v_7325 | v_28810;
assign v_28812 = v_7299 | ~v_7386;
assign v_28814 = v_7173 | v_28813;
assign v_28815 = v_7158 | ~v_7232;
assign v_28817 = v_7037 | v_28816;
assign v_28818 = v_7010 | ~v_7100;
assign v_28820 = v_6885 | v_28819;
assign v_28821 = v_6870 | ~v_6944;
assign v_28823 = v_6751 | v_28822;
assign v_28824 = v_6727 | ~v_6812;
assign v_28826 = v_6603 | v_28825;
assign v_28827 = v_6588 | ~v_6662;
assign v_28829 = v_6465 | v_28828;
assign v_28830 = v_6434 | ~v_6530;
assign v_28832 = v_6307 | v_28831;
assign v_28833 = v_6292 | ~v_6366;
assign v_28835 = v_6173 | v_28834;
assign v_28836 = v_6148 | ~v_6234;
assign v_28838 = v_6023 | v_28837;
assign v_28839 = v_6008 | ~v_6082;
assign v_28841 = v_5887 | v_28840;
assign v_28842 = v_5860 | ~v_5950;
assign v_28844 = v_5735 | v_28843;
assign v_28845 = v_5720 | ~v_5794;
assign v_28847 = v_5601 | v_28846;
assign v_28848 = v_5577 | ~v_5662;
assign v_28850 = v_5453 | v_28849;
assign v_28851 = v_5438 | ~v_5512;
assign v_28853 = v_5311 | v_28852;
assign v_28854 = v_5272 | ~v_5380;
assign v_28856 = v_5141 | v_28855;
assign v_28857 = v_5126 | ~v_5200;
assign v_28859 = v_5007 | v_28858;
assign v_28860 = v_4980 | ~v_5068;
assign v_28862 = v_4853 | v_28861;
assign v_28863 = v_4838 | ~v_4912;
assign v_28865 = v_4717 | v_28864;
assign v_28866 = v_4690 | ~v_4780;
assign v_28868 = v_4565 | v_28867;
assign v_28869 = v_4550 | ~v_4624;
assign v_28871 = v_4431 | v_28870;
assign v_28872 = v_4407 | ~v_4492;
assign v_28874 = v_4283 | v_28873;
assign v_28875 = v_4268 | ~v_4342;
assign v_28877 = v_4145 | v_28876;
assign v_28878 = v_4114 | ~v_4210;
assign v_28880 = v_3987 | v_28879;
assign v_28881 = v_3972 | ~v_4046;
assign v_28883 = v_3853 | v_28882;
assign v_28884 = v_3828 | ~v_3914;
assign v_28886 = v_3703 | v_28885;
assign v_28887 = v_3688 | ~v_3762;
assign v_28889 = v_3567 | v_28888;
assign v_28890 = v_3540 | ~v_3630;
assign v_28892 = v_3415 | v_28891;
assign v_28893 = v_3400 | ~v_3474;
assign v_28895 = v_3281 | v_28894;
assign v_28896 = v_3257 | ~v_3342;
assign v_28898 = v_3133 | v_28897;
assign v_28899 = v_3118 | ~v_3192;
assign v_28901 = v_2993 | v_28900;
assign v_28902 = v_2958 | ~v_3060;
assign v_28904 = v_2829 | v_28903;
assign v_28905 = v_2814 | ~v_2888;
assign v_28907 = v_2695 | v_28906;
assign v_28908 = v_2669 | ~v_2756;
assign v_28910 = v_2543 | v_28909;
assign v_28911 = v_2528 | ~v_2602;
assign v_28913 = v_2407 | v_28912;
assign v_28914 = v_2380 | ~v_2470;
assign v_28916 = v_2255 | v_28915;
assign v_28917 = v_2240 | ~v_2314;
assign v_28919 = v_2121 | v_28918;
assign v_28920 = v_2097 | ~v_2182;
assign v_28922 = v_1973 | v_28921;
assign v_28923 = v_1958 | ~v_2032;
assign v_28925 = v_1835 | v_28924;
assign v_28926 = v_1804 | ~v_1900;
assign v_28928 = v_1677 | v_28927;
assign v_28929 = v_1662 | ~v_1736;
assign v_28931 = v_1543 | v_28930;
assign v_28932 = v_1518 | ~v_1604;
assign v_28934 = v_1393 | v_28933;
assign v_28935 = v_1378 | ~v_1452;
assign v_28937 = v_1257 | v_28936;
assign v_28938 = v_1230 | ~v_1320;
assign v_28940 = v_1105 | v_28939;
assign v_28941 = v_1090 | ~v_1164;
assign v_28943 = v_971 | v_28942;
assign v_28944 = v_947 | ~v_1032;
assign v_28946 = v_827 | v_28945;
assign v_28947 = v_811 | ~v_886;
assign v_28949 = v_658 | v_28948;
assign v_28950 = v_359 | ~v_761;
assign v_28954 = v_9639 | v_9872;
assign v_28955 = v_9611 | v_9740;
assign v_28957 = v_9483 | v_28956;
assign v_28958 = v_9468 | v_9582;
assign v_28960 = v_9347 | v_28959;
assign v_28961 = v_9320 | v_9450;
assign v_28963 = v_9195 | v_28962;
assign v_28964 = v_9180 | v_9294;
assign v_28966 = v_9061 | v_28965;
assign v_28967 = v_9037 | v_9162;
assign v_28969 = v_8913 | v_28968;
assign v_28970 = v_8898 | v_9012;
assign v_28972 = v_8775 | v_28971;
assign v_28973 = v_8744 | v_8880;
assign v_28975 = v_8617 | v_28974;
assign v_28976 = v_8602 | v_8716;
assign v_28978 = v_8483 | v_28977;
assign v_28979 = v_8458 | v_8584;
assign v_28981 = v_8333 | v_28980;
assign v_28982 = v_8318 | ~v_8432;
assign v_28984 = v_8197 | v_28983;
assign v_28985 = v_8170 | ~v_8300;
assign v_28987 = v_8045 | v_28986;
assign v_28988 = v_8030 | ~v_8144;
assign v_28990 = v_7911 | v_28989;
assign v_28991 = v_7887 | v_8012;
assign v_28993 = v_7763 | v_28992;
assign v_28994 = v_7748 | v_7862;
assign v_28996 = v_7623 | v_28995;
assign v_28997 = v_7588 | v_7730;
assign v_28999 = v_7459 | v_28998;
assign v_29000 = v_7444 | v_7558;
assign v_29002 = v_7325 | v_29001;
assign v_29003 = v_7299 | v_7426;
assign v_29005 = v_7173 | v_29004;
assign v_29006 = v_7158 | ~v_7272;
assign v_29008 = v_7037 | v_29007;
assign v_29009 = v_7010 | v_7140;
assign v_29011 = v_6885 | v_29010;
assign v_29012 = v_6870 | ~v_6984;
assign v_29014 = v_6751 | v_29013;
assign v_29015 = v_6727 | ~v_6852;
assign v_29017 = v_6603 | v_29016;
assign v_29018 = v_6588 | ~v_6702;
assign v_29020 = v_6465 | v_29019;
assign v_29021 = v_6434 | v_6570;
assign v_29023 = v_6307 | v_29022;
assign v_29024 = v_6292 | v_6406;
assign v_29026 = v_6173 | v_29025;
assign v_29027 = v_6148 | ~v_6274;
assign v_29029 = v_6023 | v_29028;
assign v_29030 = v_6008 | ~v_6122;
assign v_29032 = v_5887 | v_29031;
assign v_29033 = v_5860 | ~v_5990;
assign v_29035 = v_5735 | v_29034;
assign v_29036 = v_5720 | ~v_5834;
assign v_29038 = v_5601 | v_29037;
assign v_29039 = v_5577 | ~v_5702;
assign v_29041 = v_5453 | v_29040;
assign v_29042 = v_5438 | ~v_5552;
assign v_29044 = v_5311 | v_29043;
assign v_29045 = v_5272 | v_5420;
assign v_29047 = v_5141 | v_29046;
assign v_29048 = v_5126 | v_5240;
assign v_29050 = v_5007 | v_29049;
assign v_29051 = v_4980 | ~v_5108;
assign v_29053 = v_4853 | v_29052;
assign v_29054 = v_4838 | ~v_4952;
assign v_29056 = v_4717 | v_29055;
assign v_29057 = v_4690 | ~v_4820;
assign v_29059 = v_4565 | v_29058;
assign v_29060 = v_4550 | ~v_4664;
assign v_29062 = v_4431 | v_29061;
assign v_29063 = v_4407 | ~v_4532;
assign v_29065 = v_4283 | v_29064;
assign v_29066 = v_4268 | ~v_4382;
assign v_29068 = v_4145 | v_29067;
assign v_29069 = v_4114 | v_4250;
assign v_29071 = v_3987 | v_29070;
assign v_29072 = v_3972 | v_4086;
assign v_29074 = v_3853 | v_29073;
assign v_29075 = v_3828 | v_3954;
assign v_29077 = v_3703 | v_29076;
assign v_29078 = v_3688 | v_3802;
assign v_29080 = v_3567 | v_29079;
assign v_29081 = v_3540 | v_3670;
assign v_29083 = v_3415 | v_29082;
assign v_29084 = v_3400 | ~v_3514;
assign v_29086 = v_3281 | v_29085;
assign v_29087 = v_3257 | v_3382;
assign v_29089 = v_3133 | v_29088;
assign v_29090 = v_3118 | ~v_3232;
assign v_29092 = v_2993 | v_29091;
assign v_29093 = v_2958 | v_3100;
assign v_29095 = v_2829 | v_29094;
assign v_29096 = v_2814 | v_2928;
assign v_29098 = v_2695 | v_29097;
assign v_29099 = v_2669 | v_2796;
assign v_29101 = v_2543 | v_29100;
assign v_29102 = v_2528 | v_2642;
assign v_29104 = v_2407 | v_29103;
assign v_29105 = v_2380 | v_2510;
assign v_29107 = v_2255 | v_29106;
assign v_29108 = v_2240 | ~v_2354;
assign v_29110 = v_2121 | v_29109;
assign v_29111 = v_2097 | ~v_2222;
assign v_29113 = v_1973 | v_29112;
assign v_29114 = v_1958 | ~v_2072;
assign v_29116 = v_1835 | v_29115;
assign v_29117 = v_1804 | v_1940;
assign v_29119 = v_1677 | v_29118;
assign v_29120 = v_1662 | v_1776;
assign v_29122 = v_1543 | v_29121;
assign v_29123 = v_1518 | v_1644;
assign v_29125 = v_1393 | v_29124;
assign v_29126 = v_1378 | v_1492;
assign v_29128 = v_1257 | v_29127;
assign v_29129 = v_1230 | v_1360;
assign v_29131 = v_1105 | v_29130;
assign v_29132 = v_1090 | v_1204;
assign v_29134 = v_971 | v_29133;
assign v_29135 = v_947 | v_1072;
assign v_29137 = v_827 | v_29136;
assign v_29138 = v_811 | v_922;
assign v_29140 = v_658 | v_29139;
assign v_29141 = v_359 | v_793;
assign v_29147 = ~v_361 | v_29146;
assign v_29148 = v_9051 | ~v_9784;
assign v_29149 = v_9026 | ~v_9652;
assign v_29151 = v_9052 | v_29150;
assign v_29152 = v_9027 | ~v_9494;
assign v_29154 = v_8761 | v_29153;
assign v_29155 = v_8729 | ~v_9362;
assign v_29157 = v_8762 | v_29156;
assign v_29158 = v_8730 | ~v_9206;
assign v_29160 = v_8473 | v_29159;
assign v_29161 = v_8447 | ~v_9074;
assign v_29163 = v_8474 | v_29162;
assign v_29164 = v_8448 | ~v_8924;
assign v_29166 = v_8185 | v_29165;
assign v_29167 = v_8157 | ~v_8792;
assign v_29169 = v_8186 | v_29168;
assign v_29170 = v_8158 | ~v_8628;
assign v_29172 = v_7901 | v_29171;
assign v_29173 = v_7876 | ~v_8496;
assign v_29175 = v_7902 | v_29174;
assign v_29176 = v_7877 | ~v_8344;
assign v_29178 = v_7607 | v_29177;
assign v_29179 = v_7571 | ~v_8212;
assign v_29181 = v_7608 | v_29180;
assign v_29182 = v_7572 | ~v_8056;
assign v_29184 = v_7315 | v_29183;
assign v_29185 = v_7288 | ~v_7924;
assign v_29187 = v_7316 | v_29186;
assign v_29188 = v_7289 | ~v_7774;
assign v_29190 = v_7025 | v_29189;
assign v_29191 = v_6997 | ~v_7642;
assign v_29193 = v_7026 | v_29192;
assign v_29194 = v_6998 | ~v_7470;
assign v_29196 = v_6741 | v_29195;
assign v_29197 = v_6716 | ~v_7338;
assign v_29199 = v_6742 | v_29198;
assign v_29200 = v_6717 | ~v_7184;
assign v_29202 = v_6451 | v_29201;
assign v_29203 = v_6419 | ~v_7052;
assign v_29205 = v_6452 | v_29204;
assign v_29206 = v_6420 | ~v_6896;
assign v_29208 = v_6163 | v_29207;
assign v_29209 = v_6137 | ~v_6764;
assign v_29211 = v_6164 | v_29210;
assign v_29212 = v_6138 | ~v_6614;
assign v_29214 = v_5875 | v_29213;
assign v_29215 = v_5847 | ~v_6482;
assign v_29217 = v_5876 | v_29216;
assign v_29218 = v_5848 | ~v_6318;
assign v_29220 = v_5591 | v_29219;
assign v_29221 = v_5566 | ~v_6186;
assign v_29223 = v_5592 | v_29222;
assign v_29224 = v_5567 | ~v_6034;
assign v_29226 = v_5293 | v_29225;
assign v_29227 = v_5253 | ~v_5902;
assign v_29229 = v_5294 | v_29228;
assign v_29230 = v_5254 | ~v_5746;
assign v_29232 = v_4997 | v_29231;
assign v_29233 = v_4969 | ~v_5614;
assign v_29235 = v_4998 | v_29234;
assign v_29236 = v_4970 | ~v_5464;
assign v_29238 = v_4705 | v_29237;
assign v_29239 = v_4677 | ~v_5332;
assign v_29241 = v_4706 | v_29240;
assign v_29242 = v_4678 | ~v_5152;
assign v_29244 = v_4421 | v_29243;
assign v_29245 = v_4396 | ~v_5020;
assign v_29247 = v_4422 | v_29246;
assign v_29248 = v_4397 | ~v_4864;
assign v_29250 = v_4131 | v_29249;
assign v_29251 = v_4099 | ~v_4732;
assign v_29253 = v_4132 | v_29252;
assign v_29254 = v_4100 | ~v_4576;
assign v_29256 = v_3843 | v_29255;
assign v_29257 = v_3817 | ~v_4444;
assign v_29259 = v_3844 | v_29258;
assign v_29260 = v_3818 | ~v_4294;
assign v_29262 = v_3555 | v_29261;
assign v_29263 = v_3527 | ~v_4162;
assign v_29265 = v_3556 | v_29264;
assign v_29266 = v_3528 | ~v_3998;
assign v_29268 = v_3271 | v_29267;
assign v_29269 = v_3246 | ~v_3866;
assign v_29271 = v_3272 | v_29270;
assign v_29272 = v_3247 | ~v_3714;
assign v_29274 = v_2977 | v_29273;
assign v_29275 = v_2941 | ~v_3582;
assign v_29277 = v_2978 | v_29276;
assign v_29278 = v_2942 | ~v_3426;
assign v_29280 = v_2685 | v_29279;
assign v_29281 = v_2658 | ~v_3294;
assign v_29283 = v_2686 | v_29282;
assign v_29284 = v_2659 | ~v_3144;
assign v_29286 = v_2395 | v_29285;
assign v_29287 = v_2367 | ~v_3012;
assign v_29289 = v_2396 | v_29288;
assign v_29290 = v_2368 | ~v_2840;
assign v_29292 = v_2111 | v_29291;
assign v_29293 = v_2086 | ~v_2708;
assign v_29295 = v_2112 | v_29294;
assign v_29296 = v_2087 | ~v_2554;
assign v_29298 = v_1821 | v_29297;
assign v_29299 = v_1789 | ~v_2422;
assign v_29301 = v_1822 | v_29300;
assign v_29302 = v_1790 | ~v_2266;
assign v_29304 = v_1533 | v_29303;
assign v_29305 = v_1507 | ~v_2134;
assign v_29307 = v_1534 | v_29306;
assign v_29308 = v_1508 | ~v_1984;
assign v_29310 = v_1245 | v_29309;
assign v_29311 = v_1217 | ~v_1852;
assign v_29313 = v_1246 | v_29312;
assign v_29314 = v_1218 | ~v_1688;
assign v_29316 = v_961 | v_29315;
assign v_29317 = v_936 | ~v_1556;
assign v_29319 = v_962 | v_29318;
assign v_29320 = v_937 | ~v_1404;
assign v_29322 = v_591 | v_29321;
assign v_29323 = v_92 | ~v_1272;
assign v_29325 = v_593 | v_29324;
assign v_29326 = v_94 | ~v_1116;
assign v_29328 = v_823 | v_29327;
assign v_29329 = v_806 | ~v_984;
assign v_29331 = v_9051 | ~v_9753;
assign v_29332 = v_9026 | ~v_9604;
assign v_29334 = v_9052 | v_29333;
assign v_29335 = v_9027 | ~v_9463;
assign v_29337 = v_8761 | v_29336;
assign v_29338 = v_8729 | ~v_9311;
assign v_29340 = v_8762 | v_29339;
assign v_29341 = v_8730 | ~v_9175;
assign v_29343 = v_8473 | v_29342;
assign v_29344 = v_8447 | ~v_9030;
assign v_29346 = v_8474 | v_29345;
assign v_29347 = v_8448 | ~v_8893;
assign v_29349 = v_8185 | v_29348;
assign v_29350 = v_8157 | ~v_8733;
assign v_29352 = v_8186 | v_29351;
assign v_29353 = v_8158 | ~v_8597;
assign v_29355 = v_7901 | v_29354;
assign v_29356 = v_7876 | ~v_8451;
assign v_29358 = v_7902 | v_29357;
assign v_29359 = v_7877 | ~v_8313;
assign v_29361 = v_7607 | v_29360;
assign v_29362 = v_7571 | ~v_8161;
assign v_29364 = v_7608 | v_29363;
assign v_29365 = v_7572 | ~v_8025;
assign v_29367 = v_7315 | v_29366;
assign v_29368 = v_7288 | ~v_7880;
assign v_29370 = v_7316 | v_29369;
assign v_29371 = v_7289 | ~v_7743;
assign v_29373 = v_7025 | v_29372;
assign v_29374 = v_6997 | ~v_7575;
assign v_29376 = v_7026 | v_29375;
assign v_29377 = v_6998 | ~v_7439;
assign v_29379 = v_6741 | v_29378;
assign v_29380 = v_6716 | ~v_7292;
assign v_29382 = v_6742 | v_29381;
assign v_29383 = v_6717 | ~v_7153;
assign v_29385 = v_6451 | v_29384;
assign v_29386 = v_6419 | ~v_7001;
assign v_29388 = v_6452 | v_29387;
assign v_29389 = v_6420 | ~v_6865;
assign v_29391 = v_6163 | v_29390;
assign v_29392 = v_6137 | ~v_6720;
assign v_29394 = v_6164 | v_29393;
assign v_29395 = v_6138 | ~v_6583;
assign v_29397 = v_5875 | v_29396;
assign v_29398 = v_5847 | ~v_6423;
assign v_29400 = v_5876 | v_29399;
assign v_29401 = v_5848 | ~v_6287;
assign v_29403 = v_5591 | v_29402;
assign v_29404 = v_5566 | ~v_6141;
assign v_29406 = v_5592 | v_29405;
assign v_29407 = v_5567 | ~v_6003;
assign v_29409 = v_5293 | v_29408;
assign v_29410 = v_5253 | ~v_5851;
assign v_29412 = v_5294 | v_29411;
assign v_29413 = v_5254 | ~v_5715;
assign v_29415 = v_4997 | v_29414;
assign v_29416 = v_4969 | ~v_5570;
assign v_29418 = v_4998 | v_29417;
assign v_29419 = v_4970 | ~v_5433;
assign v_29421 = v_4705 | v_29420;
assign v_29422 = v_4677 | ~v_5257;
assign v_29424 = v_4706 | v_29423;
assign v_29425 = v_4678 | ~v_5121;
assign v_29427 = v_4421 | v_29426;
assign v_29428 = v_4396 | ~v_4973;
assign v_29430 = v_4422 | v_29429;
assign v_29431 = v_4397 | ~v_4833;
assign v_29433 = v_4131 | v_29432;
assign v_29434 = v_4099 | ~v_4681;
assign v_29436 = v_4132 | v_29435;
assign v_29437 = v_4100 | ~v_4545;
assign v_29439 = v_3843 | v_29438;
assign v_29440 = v_3817 | ~v_4400;
assign v_29442 = v_3844 | v_29441;
assign v_29443 = v_3818 | ~v_4263;
assign v_29445 = v_3555 | v_29444;
assign v_29446 = v_3527 | ~v_4103;
assign v_29448 = v_3556 | v_29447;
assign v_29449 = v_3528 | ~v_3967;
assign v_29451 = v_3271 | v_29450;
assign v_29452 = v_3246 | ~v_3821;
assign v_29454 = v_3272 | v_29453;
assign v_29455 = v_3247 | ~v_3683;
assign v_29457 = v_2977 | v_29456;
assign v_29458 = v_2941 | ~v_3531;
assign v_29460 = v_2978 | v_29459;
assign v_29461 = v_2942 | ~v_3395;
assign v_29463 = v_2685 | v_29462;
assign v_29464 = v_2658 | ~v_3250;
assign v_29466 = v_2686 | v_29465;
assign v_29467 = v_2659 | ~v_3113;
assign v_29469 = v_2395 | v_29468;
assign v_29470 = v_2367 | ~v_2945;
assign v_29472 = v_2396 | v_29471;
assign v_29473 = v_2368 | ~v_2809;
assign v_29475 = v_2111 | v_29474;
assign v_29476 = v_2086 | ~v_2662;
assign v_29478 = v_2112 | v_29477;
assign v_29479 = v_2087 | ~v_2523;
assign v_29481 = v_1821 | v_29480;
assign v_29482 = v_1789 | ~v_2371;
assign v_29484 = v_1822 | v_29483;
assign v_29485 = v_1790 | ~v_2235;
assign v_29487 = v_1533 | v_29486;
assign v_29488 = v_1507 | ~v_2090;
assign v_29490 = v_1534 | v_29489;
assign v_29491 = v_1508 | ~v_1953;
assign v_29493 = v_1245 | v_29492;
assign v_29494 = v_1217 | ~v_1793;
assign v_29496 = v_1246 | v_29495;
assign v_29497 = v_1218 | ~v_1657;
assign v_29499 = v_961 | v_29498;
assign v_29500 = v_936 | ~v_1511;
assign v_29502 = v_962 | v_29501;
assign v_29503 = v_937 | ~v_1373;
assign v_29505 = v_591 | v_29504;
assign v_29506 = v_92 | ~v_1221;
assign v_29508 = v_593 | v_29507;
assign v_29509 = v_94 | ~v_1085;
assign v_29511 = v_823 | v_29510;
assign v_29512 = v_806 | ~v_940;
assign v_29515 = v_9051 | ~v_9796;
assign v_29516 = v_9026 | ~v_9664;
assign v_29518 = v_9052 | v_29517;
assign v_29519 = v_9027 | ~v_9506;
assign v_29521 = v_8761 | v_29520;
assign v_29522 = v_8729 | ~v_9374;
assign v_29524 = v_8762 | v_29523;
assign v_29525 = v_8730 | ~v_9218;
assign v_29527 = v_8473 | v_29526;
assign v_29528 = v_8447 | ~v_9086;
assign v_29530 = v_8474 | v_29529;
assign v_29531 = v_8448 | ~v_8936;
assign v_29533 = v_8185 | v_29532;
assign v_29534 = v_8157 | ~v_8804;
assign v_29536 = v_8186 | v_29535;
assign v_29537 = v_8158 | ~v_8640;
assign v_29539 = v_7901 | v_29538;
assign v_29540 = v_7876 | ~v_8508;
assign v_29542 = v_7902 | v_29541;
assign v_29543 = v_7877 | ~v_8356;
assign v_29545 = v_7607 | v_29544;
assign v_29546 = v_7571 | ~v_8224;
assign v_29548 = v_7608 | v_29547;
assign v_29549 = v_7572 | ~v_8068;
assign v_29551 = v_7315 | v_29550;
assign v_29552 = v_7288 | ~v_7936;
assign v_29554 = v_7316 | v_29553;
assign v_29555 = v_7289 | ~v_7786;
assign v_29557 = v_7025 | v_29556;
assign v_29558 = v_6997 | ~v_7654;
assign v_29560 = v_7026 | v_29559;
assign v_29561 = v_6998 | ~v_7482;
assign v_29563 = v_6741 | v_29562;
assign v_29564 = v_6716 | ~v_7350;
assign v_29566 = v_6742 | v_29565;
assign v_29567 = v_6717 | ~v_7196;
assign v_29569 = v_6451 | v_29568;
assign v_29570 = v_6419 | ~v_7064;
assign v_29572 = v_6452 | v_29571;
assign v_29573 = v_6420 | ~v_6908;
assign v_29575 = v_6163 | v_29574;
assign v_29576 = v_6137 | ~v_6776;
assign v_29578 = v_6164 | v_29577;
assign v_29579 = v_6138 | ~v_6626;
assign v_29581 = v_5875 | v_29580;
assign v_29582 = v_5847 | ~v_6494;
assign v_29584 = v_5876 | v_29583;
assign v_29585 = v_5848 | ~v_6330;
assign v_29587 = v_5591 | v_29586;
assign v_29588 = v_5566 | ~v_6198;
assign v_29590 = v_5592 | v_29589;
assign v_29591 = v_5567 | ~v_6046;
assign v_29593 = v_5293 | v_29592;
assign v_29594 = v_5253 | ~v_5914;
assign v_29596 = v_5294 | v_29595;
assign v_29597 = v_5254 | ~v_5758;
assign v_29599 = v_4997 | v_29598;
assign v_29600 = v_4969 | ~v_5626;
assign v_29602 = v_4998 | v_29601;
assign v_29603 = v_4970 | ~v_5476;
assign v_29605 = v_4705 | v_29604;
assign v_29606 = v_4677 | ~v_5344;
assign v_29608 = v_4706 | v_29607;
assign v_29609 = v_4678 | ~v_5164;
assign v_29611 = v_4421 | v_29610;
assign v_29612 = v_4396 | ~v_5032;
assign v_29614 = v_4422 | v_29613;
assign v_29615 = v_4397 | ~v_4876;
assign v_29617 = v_4131 | v_29616;
assign v_29618 = v_4099 | ~v_4744;
assign v_29620 = v_4132 | v_29619;
assign v_29621 = v_4100 | ~v_4588;
assign v_29623 = v_3843 | v_29622;
assign v_29624 = v_3817 | ~v_4456;
assign v_29626 = v_3844 | v_29625;
assign v_29627 = v_3818 | ~v_4306;
assign v_29629 = v_3555 | v_29628;
assign v_29630 = v_3527 | ~v_4174;
assign v_29632 = v_3556 | v_29631;
assign v_29633 = v_3528 | ~v_4010;
assign v_29635 = v_3271 | v_29634;
assign v_29636 = v_3246 | ~v_3878;
assign v_29638 = v_3272 | v_29637;
assign v_29639 = v_3247 | ~v_3726;
assign v_29641 = v_2977 | v_29640;
assign v_29642 = v_2941 | ~v_3594;
assign v_29644 = v_2978 | v_29643;
assign v_29645 = v_2942 | ~v_3438;
assign v_29647 = v_2685 | v_29646;
assign v_29648 = v_2658 | ~v_3306;
assign v_29650 = v_2686 | v_29649;
assign v_29651 = v_2659 | ~v_3156;
assign v_29653 = v_2395 | v_29652;
assign v_29654 = v_2367 | ~v_3024;
assign v_29656 = v_2396 | v_29655;
assign v_29657 = v_2368 | ~v_2852;
assign v_29659 = v_2111 | v_29658;
assign v_29660 = v_2086 | ~v_2720;
assign v_29662 = v_2112 | v_29661;
assign v_29663 = v_2087 | ~v_2566;
assign v_29665 = v_1821 | v_29664;
assign v_29666 = v_1789 | ~v_2434;
assign v_29668 = v_1822 | v_29667;
assign v_29669 = v_1790 | ~v_2278;
assign v_29671 = v_1533 | v_29670;
assign v_29672 = v_1507 | ~v_2146;
assign v_29674 = v_1534 | v_29673;
assign v_29675 = v_1508 | ~v_1996;
assign v_29677 = v_1245 | v_29676;
assign v_29678 = v_1217 | ~v_1864;
assign v_29680 = v_1246 | v_29679;
assign v_29681 = v_1218 | ~v_1700;
assign v_29683 = v_961 | v_29682;
assign v_29684 = v_936 | ~v_1568;
assign v_29686 = v_962 | v_29685;
assign v_29687 = v_937 | ~v_1416;
assign v_29689 = v_591 | v_29688;
assign v_29690 = v_92 | ~v_1284;
assign v_29692 = v_593 | v_29691;
assign v_29693 = v_94 | ~v_1128;
assign v_29695 = v_823 | v_29694;
assign v_29696 = v_806 | ~v_996;
assign v_29699 = v_9051 | ~v_9808;
assign v_29700 = v_9026 | ~v_9676;
assign v_29702 = v_9052 | v_29701;
assign v_29703 = v_9027 | ~v_9518;
assign v_29705 = v_8761 | v_29704;
assign v_29706 = v_8729 | ~v_9386;
assign v_29708 = v_8762 | v_29707;
assign v_29709 = v_8730 | ~v_9230;
assign v_29711 = v_8473 | v_29710;
assign v_29712 = v_8447 | ~v_9098;
assign v_29714 = v_8474 | v_29713;
assign v_29715 = v_8448 | ~v_8948;
assign v_29717 = v_8185 | v_29716;
assign v_29718 = v_8157 | ~v_8816;
assign v_29720 = v_8186 | v_29719;
assign v_29721 = v_8158 | ~v_8652;
assign v_29723 = v_7901 | v_29722;
assign v_29724 = v_7876 | ~v_8520;
assign v_29726 = v_7902 | v_29725;
assign v_29727 = v_7877 | ~v_8368;
assign v_29729 = v_7607 | v_29728;
assign v_29730 = v_7571 | ~v_8236;
assign v_29732 = v_7608 | v_29731;
assign v_29733 = v_7572 | ~v_8080;
assign v_29735 = v_7315 | v_29734;
assign v_29736 = v_7288 | ~v_7948;
assign v_29738 = v_7316 | v_29737;
assign v_29739 = v_7289 | ~v_7798;
assign v_29741 = v_7025 | v_29740;
assign v_29742 = v_6997 | ~v_7666;
assign v_29744 = v_7026 | v_29743;
assign v_29745 = v_6998 | ~v_7494;
assign v_29747 = v_6741 | v_29746;
assign v_29748 = v_6716 | ~v_7362;
assign v_29750 = v_6742 | v_29749;
assign v_29751 = v_6717 | ~v_7208;
assign v_29753 = v_6451 | v_29752;
assign v_29754 = v_6419 | ~v_7076;
assign v_29756 = v_6452 | v_29755;
assign v_29757 = v_6420 | ~v_6920;
assign v_29759 = v_6163 | v_29758;
assign v_29760 = v_6137 | ~v_6788;
assign v_29762 = v_6164 | v_29761;
assign v_29763 = v_6138 | ~v_6638;
assign v_29765 = v_5875 | v_29764;
assign v_29766 = v_5847 | ~v_6506;
assign v_29768 = v_5876 | v_29767;
assign v_29769 = v_5848 | ~v_6342;
assign v_29771 = v_5591 | v_29770;
assign v_29772 = v_5566 | ~v_6210;
assign v_29774 = v_5592 | v_29773;
assign v_29775 = v_5567 | ~v_6058;
assign v_29777 = v_5293 | v_29776;
assign v_29778 = v_5253 | ~v_5926;
assign v_29780 = v_5294 | v_29779;
assign v_29781 = v_5254 | ~v_5770;
assign v_29783 = v_4997 | v_29782;
assign v_29784 = v_4969 | ~v_5638;
assign v_29786 = v_4998 | v_29785;
assign v_29787 = v_4970 | ~v_5488;
assign v_29789 = v_4705 | v_29788;
assign v_29790 = v_4677 | ~v_5356;
assign v_29792 = v_4706 | v_29791;
assign v_29793 = v_4678 | ~v_5176;
assign v_29795 = v_4421 | v_29794;
assign v_29796 = v_4396 | ~v_5044;
assign v_29798 = v_4422 | v_29797;
assign v_29799 = v_4397 | ~v_4888;
assign v_29801 = v_4131 | v_29800;
assign v_29802 = v_4099 | ~v_4756;
assign v_29804 = v_4132 | v_29803;
assign v_29805 = v_4100 | ~v_4600;
assign v_29807 = v_3843 | v_29806;
assign v_29808 = v_3817 | ~v_4468;
assign v_29810 = v_3844 | v_29809;
assign v_29811 = v_3818 | ~v_4318;
assign v_29813 = v_3555 | v_29812;
assign v_29814 = v_3527 | ~v_4186;
assign v_29816 = v_3556 | v_29815;
assign v_29817 = v_3528 | ~v_4022;
assign v_29819 = v_3271 | v_29818;
assign v_29820 = v_3246 | ~v_3890;
assign v_29822 = v_3272 | v_29821;
assign v_29823 = v_3247 | ~v_3738;
assign v_29825 = v_2977 | v_29824;
assign v_29826 = v_2941 | ~v_3606;
assign v_29828 = v_2978 | v_29827;
assign v_29829 = v_2942 | ~v_3450;
assign v_29831 = v_2685 | v_29830;
assign v_29832 = v_2658 | ~v_3318;
assign v_29834 = v_2686 | v_29833;
assign v_29835 = v_2659 | ~v_3168;
assign v_29837 = v_2395 | v_29836;
assign v_29838 = v_2367 | ~v_3036;
assign v_29840 = v_2396 | v_29839;
assign v_29841 = v_2368 | ~v_2864;
assign v_29843 = v_2111 | v_29842;
assign v_29844 = v_2086 | ~v_2732;
assign v_29846 = v_2112 | v_29845;
assign v_29847 = v_2087 | ~v_2578;
assign v_29849 = v_1821 | v_29848;
assign v_29850 = v_1789 | ~v_2446;
assign v_29852 = v_1822 | v_29851;
assign v_29853 = v_1790 | ~v_2290;
assign v_29855 = v_1533 | v_29854;
assign v_29856 = v_1507 | ~v_2158;
assign v_29858 = v_1534 | v_29857;
assign v_29859 = v_1508 | ~v_2008;
assign v_29861 = v_1245 | v_29860;
assign v_29862 = v_1217 | ~v_1876;
assign v_29864 = v_1246 | v_29863;
assign v_29865 = v_1218 | ~v_1712;
assign v_29867 = v_961 | v_29866;
assign v_29868 = v_936 | ~v_1580;
assign v_29870 = v_962 | v_29869;
assign v_29871 = v_937 | ~v_1428;
assign v_29873 = v_591 | v_29872;
assign v_29874 = v_92 | ~v_1296;
assign v_29876 = v_593 | v_29875;
assign v_29877 = v_94 | ~v_1140;
assign v_29879 = v_823 | v_29878;
assign v_29880 = v_806 | ~v_1008;
assign v_29883 = v_9051 | ~v_9820;
assign v_29884 = v_9026 | ~v_9688;
assign v_29886 = v_9052 | v_29885;
assign v_29887 = v_9027 | ~v_9530;
assign v_29889 = v_8761 | v_29888;
assign v_29890 = v_8729 | ~v_9398;
assign v_29892 = v_8762 | v_29891;
assign v_29893 = v_8730 | ~v_9242;
assign v_29895 = v_8473 | v_29894;
assign v_29896 = v_8447 | ~v_9110;
assign v_29898 = v_8474 | v_29897;
assign v_29899 = v_8448 | ~v_8960;
assign v_29901 = v_8185 | v_29900;
assign v_29902 = v_8157 | ~v_8828;
assign v_29904 = v_8186 | v_29903;
assign v_29905 = v_8158 | ~v_8664;
assign v_29907 = v_7901 | v_29906;
assign v_29908 = v_7876 | ~v_8532;
assign v_29910 = v_7902 | v_29909;
assign v_29911 = v_7877 | ~v_8380;
assign v_29913 = v_7607 | v_29912;
assign v_29914 = v_7571 | ~v_8248;
assign v_29916 = v_7608 | v_29915;
assign v_29917 = v_7572 | ~v_8092;
assign v_29919 = v_7315 | v_29918;
assign v_29920 = v_7288 | ~v_7960;
assign v_29922 = v_7316 | v_29921;
assign v_29923 = v_7289 | ~v_7810;
assign v_29925 = v_7025 | v_29924;
assign v_29926 = v_6997 | ~v_7678;
assign v_29928 = v_7026 | v_29927;
assign v_29929 = v_6998 | ~v_7506;
assign v_29931 = v_6741 | v_29930;
assign v_29932 = v_6716 | ~v_7374;
assign v_29934 = v_6742 | v_29933;
assign v_29935 = v_6717 | ~v_7220;
assign v_29937 = v_6451 | v_29936;
assign v_29938 = v_6419 | ~v_7088;
assign v_29940 = v_6452 | v_29939;
assign v_29941 = v_6420 | ~v_6932;
assign v_29943 = v_6163 | v_29942;
assign v_29944 = v_6137 | ~v_6800;
assign v_29946 = v_6164 | v_29945;
assign v_29947 = v_6138 | ~v_6650;
assign v_29949 = v_5875 | v_29948;
assign v_29950 = v_5847 | ~v_6518;
assign v_29952 = v_5876 | v_29951;
assign v_29953 = v_5848 | ~v_6354;
assign v_29955 = v_5591 | v_29954;
assign v_29956 = v_5566 | ~v_6222;
assign v_29958 = v_5592 | v_29957;
assign v_29959 = v_5567 | ~v_6070;
assign v_29961 = v_5293 | v_29960;
assign v_29962 = v_5253 | ~v_5938;
assign v_29964 = v_5294 | v_29963;
assign v_29965 = v_5254 | ~v_5782;
assign v_29967 = v_4997 | v_29966;
assign v_29968 = v_4969 | ~v_5650;
assign v_29970 = v_4998 | v_29969;
assign v_29971 = v_4970 | ~v_5500;
assign v_29973 = v_4705 | v_29972;
assign v_29974 = v_4677 | ~v_5368;
assign v_29976 = v_4706 | v_29975;
assign v_29977 = v_4678 | ~v_5188;
assign v_29979 = v_4421 | v_29978;
assign v_29980 = v_4396 | ~v_5056;
assign v_29982 = v_4422 | v_29981;
assign v_29983 = v_4397 | ~v_4900;
assign v_29985 = v_4131 | v_29984;
assign v_29986 = v_4099 | ~v_4768;
assign v_29988 = v_4132 | v_29987;
assign v_29989 = v_4100 | ~v_4612;
assign v_29991 = v_3843 | v_29990;
assign v_29992 = v_3817 | ~v_4480;
assign v_29994 = v_3844 | v_29993;
assign v_29995 = v_3818 | ~v_4330;
assign v_29997 = v_3555 | v_29996;
assign v_29998 = v_3527 | ~v_4198;
assign v_30000 = v_3556 | v_29999;
assign v_30001 = v_3528 | ~v_4034;
assign v_30003 = v_3271 | v_30002;
assign v_30004 = v_3246 | ~v_3902;
assign v_30006 = v_3272 | v_30005;
assign v_30007 = v_3247 | ~v_3750;
assign v_30009 = v_2977 | v_30008;
assign v_30010 = v_2941 | ~v_3618;
assign v_30012 = v_2978 | v_30011;
assign v_30013 = v_2942 | ~v_3462;
assign v_30015 = v_2685 | v_30014;
assign v_30016 = v_2658 | ~v_3330;
assign v_30018 = v_2686 | v_30017;
assign v_30019 = v_2659 | ~v_3180;
assign v_30021 = v_2395 | v_30020;
assign v_30022 = v_2367 | ~v_3048;
assign v_30024 = v_2396 | v_30023;
assign v_30025 = v_2368 | ~v_2876;
assign v_30027 = v_2111 | v_30026;
assign v_30028 = v_2086 | ~v_2744;
assign v_30030 = v_2112 | v_30029;
assign v_30031 = v_2087 | ~v_2590;
assign v_30033 = v_1821 | v_30032;
assign v_30034 = v_1789 | ~v_2458;
assign v_30036 = v_1822 | v_30035;
assign v_30037 = v_1790 | ~v_2302;
assign v_30039 = v_1533 | v_30038;
assign v_30040 = v_1507 | ~v_2170;
assign v_30042 = v_1534 | v_30041;
assign v_30043 = v_1508 | ~v_2020;
assign v_30045 = v_1245 | v_30044;
assign v_30046 = v_1217 | ~v_1888;
assign v_30048 = v_1246 | v_30047;
assign v_30049 = v_1218 | ~v_1724;
assign v_30051 = v_961 | v_30050;
assign v_30052 = v_936 | ~v_1592;
assign v_30054 = v_962 | v_30053;
assign v_30055 = v_937 | ~v_1440;
assign v_30057 = v_591 | v_30056;
assign v_30058 = v_92 | ~v_1308;
assign v_30060 = v_593 | v_30059;
assign v_30061 = v_94 | ~v_1152;
assign v_30063 = v_823 | v_30062;
assign v_30064 = v_806 | ~v_1020;
assign v_30067 = v_9051 | ~v_9832;
assign v_30068 = v_9026 | ~v_9700;
assign v_30070 = v_9052 | v_30069;
assign v_30071 = v_9027 | ~v_9542;
assign v_30073 = v_8761 | v_30072;
assign v_30074 = v_8729 | ~v_9410;
assign v_30076 = v_8762 | v_30075;
assign v_30077 = v_8730 | ~v_9254;
assign v_30079 = v_8473 | v_30078;
assign v_30080 = v_8447 | ~v_9122;
assign v_30082 = v_8474 | v_30081;
assign v_30083 = v_8448 | ~v_8972;
assign v_30085 = v_8185 | v_30084;
assign v_30086 = v_8157 | ~v_8840;
assign v_30088 = v_8186 | v_30087;
assign v_30089 = v_8158 | ~v_8676;
assign v_30091 = v_7901 | v_30090;
assign v_30092 = v_7876 | ~v_8544;
assign v_30094 = v_7902 | v_30093;
assign v_30095 = v_7877 | ~v_8392;
assign v_30097 = v_7607 | v_30096;
assign v_30098 = v_7571 | ~v_8260;
assign v_30100 = v_7608 | v_30099;
assign v_30101 = v_7572 | ~v_8104;
assign v_30103 = v_7315 | v_30102;
assign v_30104 = v_7288 | ~v_7972;
assign v_30106 = v_7316 | v_30105;
assign v_30107 = v_7289 | ~v_7822;
assign v_30109 = v_7025 | v_30108;
assign v_30110 = v_6997 | ~v_7690;
assign v_30112 = v_7026 | v_30111;
assign v_30113 = v_6998 | ~v_7518;
assign v_30115 = v_6741 | v_30114;
assign v_30116 = v_6716 | ~v_7386;
assign v_30118 = v_6742 | v_30117;
assign v_30119 = v_6717 | ~v_7232;
assign v_30121 = v_6451 | v_30120;
assign v_30122 = v_6419 | ~v_7100;
assign v_30124 = v_6452 | v_30123;
assign v_30125 = v_6420 | ~v_6944;
assign v_30127 = v_6163 | v_30126;
assign v_30128 = v_6137 | ~v_6812;
assign v_30130 = v_6164 | v_30129;
assign v_30131 = v_6138 | ~v_6662;
assign v_30133 = v_5875 | v_30132;
assign v_30134 = v_5847 | ~v_6530;
assign v_30136 = v_5876 | v_30135;
assign v_30137 = v_5848 | ~v_6366;
assign v_30139 = v_5591 | v_30138;
assign v_30140 = v_5566 | ~v_6234;
assign v_30142 = v_5592 | v_30141;
assign v_30143 = v_5567 | ~v_6082;
assign v_30145 = v_5293 | v_30144;
assign v_30146 = v_5253 | ~v_5950;
assign v_30148 = v_5294 | v_30147;
assign v_30149 = v_5254 | ~v_5794;
assign v_30151 = v_4997 | v_30150;
assign v_30152 = v_4969 | ~v_5662;
assign v_30154 = v_4998 | v_30153;
assign v_30155 = v_4970 | ~v_5512;
assign v_30157 = v_4705 | v_30156;
assign v_30158 = v_4677 | ~v_5380;
assign v_30160 = v_4706 | v_30159;
assign v_30161 = v_4678 | ~v_5200;
assign v_30163 = v_4421 | v_30162;
assign v_30164 = v_4396 | ~v_5068;
assign v_30166 = v_4422 | v_30165;
assign v_30167 = v_4397 | ~v_4912;
assign v_30169 = v_4131 | v_30168;
assign v_30170 = v_4099 | ~v_4780;
assign v_30172 = v_4132 | v_30171;
assign v_30173 = v_4100 | ~v_4624;
assign v_30175 = v_3843 | v_30174;
assign v_30176 = v_3817 | ~v_4492;
assign v_30178 = v_3844 | v_30177;
assign v_30179 = v_3818 | ~v_4342;
assign v_30181 = v_3555 | v_30180;
assign v_30182 = v_3527 | ~v_4210;
assign v_30184 = v_3556 | v_30183;
assign v_30185 = v_3528 | ~v_4046;
assign v_30187 = v_3271 | v_30186;
assign v_30188 = v_3246 | ~v_3914;
assign v_30190 = v_3272 | v_30189;
assign v_30191 = v_3247 | ~v_3762;
assign v_30193 = v_2977 | v_30192;
assign v_30194 = v_2941 | ~v_3630;
assign v_30196 = v_2978 | v_30195;
assign v_30197 = v_2942 | ~v_3474;
assign v_30199 = v_2685 | v_30198;
assign v_30200 = v_2658 | ~v_3342;
assign v_30202 = v_2686 | v_30201;
assign v_30203 = v_2659 | ~v_3192;
assign v_30205 = v_2395 | v_30204;
assign v_30206 = v_2367 | ~v_3060;
assign v_30208 = v_2396 | v_30207;
assign v_30209 = v_2368 | ~v_2888;
assign v_30211 = v_2111 | v_30210;
assign v_30212 = v_2086 | ~v_2756;
assign v_30214 = v_2112 | v_30213;
assign v_30215 = v_2087 | ~v_2602;
assign v_30217 = v_1821 | v_30216;
assign v_30218 = v_1789 | ~v_2470;
assign v_30220 = v_1822 | v_30219;
assign v_30221 = v_1790 | ~v_2314;
assign v_30223 = v_1533 | v_30222;
assign v_30224 = v_1507 | ~v_2182;
assign v_30226 = v_1534 | v_30225;
assign v_30227 = v_1508 | ~v_2032;
assign v_30229 = v_1245 | v_30228;
assign v_30230 = v_1217 | ~v_1900;
assign v_30232 = v_1246 | v_30231;
assign v_30233 = v_1218 | ~v_1736;
assign v_30235 = v_961 | v_30234;
assign v_30236 = v_936 | ~v_1604;
assign v_30238 = v_962 | v_30237;
assign v_30239 = v_937 | ~v_1452;
assign v_30241 = v_591 | v_30240;
assign v_30242 = v_92 | ~v_1320;
assign v_30244 = v_593 | v_30243;
assign v_30245 = v_94 | ~v_1164;
assign v_30247 = v_823 | v_30246;
assign v_30248 = v_806 | ~v_1032;
assign v_30251 = v_9051 | ~v_9844;
assign v_30252 = v_9026 | ~v_9712;
assign v_30254 = v_9052 | v_30253;
assign v_30255 = v_9027 | ~v_9554;
assign v_30257 = v_8761 | v_30256;
assign v_30258 = v_8729 | ~v_9422;
assign v_30260 = v_8762 | v_30259;
assign v_30261 = v_8730 | ~v_9266;
assign v_30263 = v_8473 | v_30262;
assign v_30264 = v_8447 | ~v_9134;
assign v_30266 = v_8474 | v_30265;
assign v_30267 = v_8448 | ~v_8984;
assign v_30269 = v_8185 | v_30268;
assign v_30270 = v_8157 | ~v_8852;
assign v_30272 = v_8186 | v_30271;
assign v_30273 = v_8158 | ~v_8688;
assign v_30275 = v_7901 | v_30274;
assign v_30276 = v_7876 | ~v_8556;
assign v_30278 = v_7902 | v_30277;
assign v_30279 = v_7877 | ~v_8404;
assign v_30281 = v_7607 | v_30280;
assign v_30282 = v_7571 | ~v_8272;
assign v_30284 = v_7608 | v_30283;
assign v_30285 = v_7572 | ~v_8116;
assign v_30287 = v_7315 | v_30286;
assign v_30288 = v_7288 | ~v_7984;
assign v_30290 = v_7316 | v_30289;
assign v_30291 = v_7289 | ~v_7834;
assign v_30293 = v_7025 | v_30292;
assign v_30294 = v_6997 | ~v_7702;
assign v_30296 = v_7026 | v_30295;
assign v_30297 = v_6998 | ~v_7530;
assign v_30299 = v_6741 | v_30298;
assign v_30300 = v_6716 | ~v_7398;
assign v_30302 = v_6742 | v_30301;
assign v_30303 = v_6717 | ~v_7244;
assign v_30305 = v_6451 | v_30304;
assign v_30306 = v_6419 | ~v_7112;
assign v_30308 = v_6452 | v_30307;
assign v_30309 = v_6420 | ~v_6956;
assign v_30311 = v_6163 | v_30310;
assign v_30312 = v_6137 | v_6824;
assign v_30314 = v_6164 | v_30313;
assign v_30315 = v_6138 | ~v_6674;
assign v_30317 = v_5875 | v_30316;
assign v_30318 = v_5847 | ~v_6542;
assign v_30320 = v_5876 | v_30319;
assign v_30321 = v_5848 | ~v_6378;
assign v_30323 = v_5591 | v_30322;
assign v_30324 = v_5566 | ~v_6246;
assign v_30326 = v_5592 | v_30325;
assign v_30327 = v_5567 | v_6094;
assign v_30329 = v_5293 | v_30328;
assign v_30330 = v_5253 | ~v_5962;
assign v_30332 = v_5294 | v_30331;
assign v_30333 = v_5254 | v_5806;
assign v_30335 = v_4997 | v_30334;
assign v_30336 = v_4969 | ~v_5674;
assign v_30338 = v_4998 | v_30337;
assign v_30339 = v_4970 | ~v_5524;
assign v_30341 = v_4705 | v_30340;
assign v_30342 = v_4677 | ~v_5392;
assign v_30344 = v_4706 | v_30343;
assign v_30345 = v_4678 | ~v_5212;
assign v_30347 = v_4421 | v_30346;
assign v_30348 = v_4396 | ~v_5080;
assign v_30350 = v_4422 | v_30349;
assign v_30351 = v_4397 | ~v_4924;
assign v_30353 = v_4131 | v_30352;
assign v_30354 = v_4099 | ~v_4792;
assign v_30356 = v_4132 | v_30355;
assign v_30357 = v_4100 | ~v_4636;
assign v_30359 = v_3843 | v_30358;
assign v_30360 = v_3817 | ~v_4504;
assign v_30362 = v_3844 | v_30361;
assign v_30363 = v_3818 | ~v_4354;
assign v_30365 = v_3555 | v_30364;
assign v_30366 = v_3527 | ~v_4222;
assign v_30368 = v_3556 | v_30367;
assign v_30369 = v_3528 | ~v_4058;
assign v_30371 = v_3271 | v_30370;
assign v_30372 = v_3246 | ~v_3926;
assign v_30374 = v_3272 | v_30373;
assign v_30375 = v_3247 | ~v_3774;
assign v_30377 = v_2977 | v_30376;
assign v_30378 = v_2941 | ~v_3642;
assign v_30380 = v_2978 | v_30379;
assign v_30381 = v_2942 | ~v_3486;
assign v_30383 = v_2685 | v_30382;
assign v_30384 = v_2658 | ~v_3354;
assign v_30386 = v_2686 | v_30385;
assign v_30387 = v_2659 | v_3204;
assign v_30389 = v_2395 | v_30388;
assign v_30390 = v_2367 | ~v_3072;
assign v_30392 = v_2396 | v_30391;
assign v_30393 = v_2368 | ~v_2900;
assign v_30395 = v_2111 | v_30394;
assign v_30396 = v_2086 | ~v_2768;
assign v_30398 = v_2112 | v_30397;
assign v_30399 = v_2087 | ~v_2614;
assign v_30401 = v_1821 | v_30400;
assign v_30402 = v_1789 | ~v_2482;
assign v_30404 = v_1822 | v_30403;
assign v_30405 = v_1790 | ~v_2326;
assign v_30407 = v_1533 | v_30406;
assign v_30408 = v_1507 | ~v_2194;
assign v_30410 = v_1534 | v_30409;
assign v_30411 = v_1508 | ~v_2044;
assign v_30413 = v_1245 | v_30412;
assign v_30414 = v_1217 | ~v_1912;
assign v_30416 = v_1246 | v_30415;
assign v_30417 = v_1218 | ~v_1748;
assign v_30419 = v_961 | v_30418;
assign v_30420 = v_936 | ~v_1616;
assign v_30422 = v_962 | v_30421;
assign v_30423 = v_937 | ~v_1464;
assign v_30425 = v_591 | v_30424;
assign v_30426 = v_92 | ~v_1332;
assign v_30428 = v_593 | v_30427;
assign v_30429 = v_94 | ~v_1176;
assign v_30431 = v_823 | v_30430;
assign v_30432 = v_806 | ~v_1044;
assign v_30435 = v_9051 | v_9872;
assign v_30436 = v_9026 | v_9740;
assign v_30438 = v_9052 | v_30437;
assign v_30439 = v_9027 | v_9582;
assign v_30441 = v_8761 | v_30440;
assign v_30442 = v_8729 | v_9450;
assign v_30444 = v_8762 | v_30443;
assign v_30445 = v_8730 | v_9294;
assign v_30447 = v_8473 | v_30446;
assign v_30448 = v_8447 | v_9162;
assign v_30450 = v_8474 | v_30449;
assign v_30451 = v_8448 | v_9012;
assign v_30453 = v_8185 | v_30452;
assign v_30454 = v_8157 | v_8880;
assign v_30456 = v_8186 | v_30455;
assign v_30457 = v_8158 | v_8716;
assign v_30459 = v_7901 | v_30458;
assign v_30460 = v_7876 | v_8584;
assign v_30462 = v_7902 | v_30461;
assign v_30463 = v_7877 | ~v_8432;
assign v_30465 = v_7607 | v_30464;
assign v_30466 = v_7571 | ~v_8300;
assign v_30468 = v_7608 | v_30467;
assign v_30469 = v_7572 | ~v_8144;
assign v_30471 = v_7315 | v_30470;
assign v_30472 = v_7288 | v_8012;
assign v_30474 = v_7316 | v_30473;
assign v_30475 = v_7289 | v_7862;
assign v_30477 = v_7025 | v_30476;
assign v_30478 = v_6997 | v_7730;
assign v_30480 = v_7026 | v_30479;
assign v_30481 = v_6998 | v_7558;
assign v_30483 = v_6741 | v_30482;
assign v_30484 = v_6716 | v_7426;
assign v_30486 = v_6742 | v_30485;
assign v_30487 = v_6717 | ~v_7272;
assign v_30489 = v_6451 | v_30488;
assign v_30490 = v_6419 | v_7140;
assign v_30492 = v_6452 | v_30491;
assign v_30493 = v_6420 | ~v_6984;
assign v_30495 = v_6163 | v_30494;
assign v_30496 = v_6137 | ~v_6852;
assign v_30498 = v_6164 | v_30497;
assign v_30499 = v_6138 | ~v_6702;
assign v_30501 = v_5875 | v_30500;
assign v_30502 = v_5847 | v_6570;
assign v_30504 = v_5876 | v_30503;
assign v_30505 = v_5848 | v_6406;
assign v_30507 = v_5591 | v_30506;
assign v_30508 = v_5566 | ~v_6274;
assign v_30510 = v_5592 | v_30509;
assign v_30511 = v_5567 | ~v_6122;
assign v_30513 = v_5293 | v_30512;
assign v_30514 = v_5253 | ~v_5990;
assign v_30516 = v_5294 | v_30515;
assign v_30517 = v_5254 | ~v_5834;
assign v_30519 = v_4997 | v_30518;
assign v_30520 = v_4969 | ~v_5702;
assign v_30522 = v_4998 | v_30521;
assign v_30523 = v_4970 | ~v_5552;
assign v_30525 = v_4705 | v_30524;
assign v_30526 = v_4677 | v_5420;
assign v_30528 = v_4706 | v_30527;
assign v_30529 = v_4678 | v_5240;
assign v_30531 = v_4421 | v_30530;
assign v_30532 = v_4396 | ~v_5108;
assign v_30534 = v_4422 | v_30533;
assign v_30535 = v_4397 | ~v_4952;
assign v_30537 = v_4131 | v_30536;
assign v_30538 = v_4099 | ~v_4820;
assign v_30540 = v_4132 | v_30539;
assign v_30541 = v_4100 | ~v_4664;
assign v_30543 = v_3843 | v_30542;
assign v_30544 = v_3817 | ~v_4532;
assign v_30546 = v_3844 | v_30545;
assign v_30547 = v_3818 | ~v_4382;
assign v_30549 = v_3555 | v_30548;
assign v_30550 = v_3527 | v_4250;
assign v_30552 = v_3556 | v_30551;
assign v_30553 = v_3528 | v_4086;
assign v_30555 = v_3271 | v_30554;
assign v_30556 = v_3246 | v_3954;
assign v_30558 = v_3272 | v_30557;
assign v_30559 = v_3247 | v_3802;
assign v_30561 = v_2977 | v_30560;
assign v_30562 = v_2941 | v_3670;
assign v_30564 = v_2978 | v_30563;
assign v_30565 = v_2942 | ~v_3514;
assign v_30567 = v_2685 | v_30566;
assign v_30568 = v_2658 | v_3382;
assign v_30570 = v_2686 | v_30569;
assign v_30571 = v_2659 | ~v_3232;
assign v_30573 = v_2395 | v_30572;
assign v_30574 = v_2367 | v_3100;
assign v_30576 = v_2396 | v_30575;
assign v_30577 = v_2368 | v_2928;
assign v_30579 = v_2111 | v_30578;
assign v_30580 = v_2086 | v_2796;
assign v_30582 = v_2112 | v_30581;
assign v_30583 = v_2087 | v_2642;
assign v_30585 = v_1821 | v_30584;
assign v_30586 = v_1789 | v_2510;
assign v_30588 = v_1822 | v_30587;
assign v_30589 = v_1790 | ~v_2354;
assign v_30591 = v_1533 | v_30590;
assign v_30592 = v_1507 | ~v_2222;
assign v_30594 = v_1534 | v_30593;
assign v_30595 = v_1508 | ~v_2072;
assign v_30597 = v_1245 | v_30596;
assign v_30598 = v_1217 | v_1940;
assign v_30600 = v_1246 | v_30599;
assign v_30601 = v_1218 | v_1776;
assign v_30603 = v_961 | v_30602;
assign v_30604 = v_936 | v_1644;
assign v_30606 = v_962 | v_30605;
assign v_30607 = v_937 | v_1492;
assign v_30609 = v_591 | v_30608;
assign v_30610 = v_92 | v_1360;
assign v_30612 = v_593 | v_30611;
assign v_30613 = v_94 | v_1204;
assign v_30615 = v_823 | v_30614;
assign v_30616 = v_806 | v_1072;
assign v_30619 = v_9336 | ~v_9784;
assign v_30620 = v_9308 | ~v_9652;
assign v_30622 = v_9051 | v_30621;
assign v_30623 = v_9026 | ~v_9494;
assign v_30625 = v_9052 | v_30624;
assign v_30626 = v_9027 | ~v_9362;
assign v_30628 = v_8761 | v_30627;
assign v_30629 = v_8729 | ~v_9206;
assign v_30631 = v_8762 | v_30630;
assign v_30632 = v_8730 | ~v_9074;
assign v_30634 = v_8473 | v_30633;
assign v_30635 = v_8447 | ~v_8924;
assign v_30637 = v_8474 | v_30636;
assign v_30638 = v_8448 | ~v_8792;
assign v_30640 = v_8185 | v_30639;
assign v_30641 = v_8157 | ~v_8628;
assign v_30643 = v_8186 | v_30642;
assign v_30644 = v_8158 | ~v_8496;
assign v_30646 = v_7901 | v_30645;
assign v_30647 = v_7876 | ~v_8344;
assign v_30649 = v_7902 | v_30648;
assign v_30650 = v_7877 | ~v_8212;
assign v_30652 = v_7607 | v_30651;
assign v_30653 = v_7571 | ~v_8056;
assign v_30655 = v_7608 | v_30654;
assign v_30656 = v_7572 | ~v_7924;
assign v_30658 = v_7315 | v_30657;
assign v_30659 = v_7288 | ~v_7774;
assign v_30661 = v_7316 | v_30660;
assign v_30662 = v_7289 | ~v_7642;
assign v_30664 = v_7025 | v_30663;
assign v_30665 = v_6997 | ~v_7470;
assign v_30667 = v_7026 | v_30666;
assign v_30668 = v_6998 | ~v_7338;
assign v_30670 = v_6741 | v_30669;
assign v_30671 = v_6716 | ~v_7184;
assign v_30673 = v_6742 | v_30672;
assign v_30674 = v_6717 | ~v_7052;
assign v_30676 = v_6451 | v_30675;
assign v_30677 = v_6419 | ~v_6896;
assign v_30679 = v_6452 | v_30678;
assign v_30680 = v_6420 | ~v_6764;
assign v_30682 = v_6163 | v_30681;
assign v_30683 = v_6137 | ~v_6614;
assign v_30685 = v_6164 | v_30684;
assign v_30686 = v_6138 | ~v_6482;
assign v_30688 = v_5875 | v_30687;
assign v_30689 = v_5847 | ~v_6318;
assign v_30691 = v_5876 | v_30690;
assign v_30692 = v_5848 | ~v_6186;
assign v_30694 = v_5591 | v_30693;
assign v_30695 = v_5566 | ~v_6034;
assign v_30697 = v_5592 | v_30696;
assign v_30698 = v_5567 | ~v_5902;
assign v_30700 = v_5293 | v_30699;
assign v_30701 = v_5253 | ~v_5746;
assign v_30703 = v_5294 | v_30702;
assign v_30704 = v_5254 | ~v_5614;
assign v_30706 = v_4997 | v_30705;
assign v_30707 = v_4969 | ~v_5464;
assign v_30709 = v_4998 | v_30708;
assign v_30710 = v_4970 | ~v_5332;
assign v_30712 = v_4705 | v_30711;
assign v_30713 = v_4677 | ~v_5152;
assign v_30715 = v_4706 | v_30714;
assign v_30716 = v_4678 | ~v_5020;
assign v_30718 = v_4421 | v_30717;
assign v_30719 = v_4396 | ~v_4864;
assign v_30721 = v_4422 | v_30720;
assign v_30722 = v_4397 | ~v_4732;
assign v_30724 = v_4131 | v_30723;
assign v_30725 = v_4099 | ~v_4576;
assign v_30727 = v_4132 | v_30726;
assign v_30728 = v_4100 | ~v_4444;
assign v_30730 = v_3843 | v_30729;
assign v_30731 = v_3817 | ~v_4294;
assign v_30733 = v_3844 | v_30732;
assign v_30734 = v_3818 | ~v_4162;
assign v_30736 = v_3555 | v_30735;
assign v_30737 = v_3527 | ~v_3998;
assign v_30739 = v_3556 | v_30738;
assign v_30740 = v_3528 | ~v_3866;
assign v_30742 = v_3271 | v_30741;
assign v_30743 = v_3246 | ~v_3714;
assign v_30745 = v_3272 | v_30744;
assign v_30746 = v_3247 | ~v_3582;
assign v_30748 = v_2977 | v_30747;
assign v_30749 = v_2941 | ~v_3426;
assign v_30751 = v_2978 | v_30750;
assign v_30752 = v_2942 | ~v_3294;
assign v_30754 = v_2685 | v_30753;
assign v_30755 = v_2658 | ~v_3144;
assign v_30757 = v_2686 | v_30756;
assign v_30758 = v_2659 | ~v_3012;
assign v_30760 = v_2395 | v_30759;
assign v_30761 = v_2367 | ~v_2840;
assign v_30763 = v_2396 | v_30762;
assign v_30764 = v_2368 | ~v_2708;
assign v_30766 = v_2111 | v_30765;
assign v_30767 = v_2086 | ~v_2554;
assign v_30769 = v_2112 | v_30768;
assign v_30770 = v_2087 | ~v_2422;
assign v_30772 = v_1821 | v_30771;
assign v_30773 = v_1789 | ~v_2266;
assign v_30775 = v_1822 | v_30774;
assign v_30776 = v_1790 | ~v_2134;
assign v_30778 = v_1533 | v_30777;
assign v_30779 = v_1507 | ~v_1984;
assign v_30781 = v_1534 | v_30780;
assign v_30782 = v_1508 | ~v_1852;
assign v_30784 = v_1245 | v_30783;
assign v_30785 = v_1217 | ~v_1688;
assign v_30787 = v_1246 | v_30786;
assign v_30788 = v_1218 | ~v_1556;
assign v_30790 = v_961 | v_30789;
assign v_30791 = v_936 | ~v_1404;
assign v_30793 = v_962 | v_30792;
assign v_30794 = v_937 | ~v_1272;
assign v_30796 = v_591 | v_30795;
assign v_30797 = v_92 | ~v_1116;
assign v_30799 = v_593 | v_30798;
assign v_30800 = v_94 | ~v_984;
assign v_30802 = v_823 | v_30801;
assign v_30803 = v_806 | ~v_838;
assign v_30805 = v_9336 | ~v_9753;
assign v_30806 = v_9308 | ~v_9604;
assign v_30808 = v_9051 | v_30807;
assign v_30809 = v_9026 | ~v_9463;
assign v_30811 = v_9052 | v_30810;
assign v_30812 = v_9027 | ~v_9311;
assign v_30814 = v_8761 | v_30813;
assign v_30815 = v_8729 | ~v_9175;
assign v_30817 = v_8762 | v_30816;
assign v_30818 = v_8730 | ~v_9030;
assign v_30820 = v_8473 | v_30819;
assign v_30821 = v_8447 | ~v_8893;
assign v_30823 = v_8474 | v_30822;
assign v_30824 = v_8448 | ~v_8733;
assign v_30826 = v_8185 | v_30825;
assign v_30827 = v_8157 | ~v_8597;
assign v_30829 = v_8186 | v_30828;
assign v_30830 = v_8158 | ~v_8451;
assign v_30832 = v_7901 | v_30831;
assign v_30833 = v_7876 | ~v_8313;
assign v_30835 = v_7902 | v_30834;
assign v_30836 = v_7877 | ~v_8161;
assign v_30838 = v_7607 | v_30837;
assign v_30839 = v_7571 | ~v_8025;
assign v_30841 = v_7608 | v_30840;
assign v_30842 = v_7572 | ~v_7880;
assign v_30844 = v_7315 | v_30843;
assign v_30845 = v_7288 | ~v_7743;
assign v_30847 = v_7316 | v_30846;
assign v_30848 = v_7289 | ~v_7575;
assign v_30850 = v_7025 | v_30849;
assign v_30851 = v_6997 | ~v_7439;
assign v_30853 = v_7026 | v_30852;
assign v_30854 = v_6998 | ~v_7292;
assign v_30856 = v_6741 | v_30855;
assign v_30857 = v_6716 | ~v_7153;
assign v_30859 = v_6742 | v_30858;
assign v_30860 = v_6717 | ~v_7001;
assign v_30862 = v_6451 | v_30861;
assign v_30863 = v_6419 | ~v_6865;
assign v_30865 = v_6452 | v_30864;
assign v_30866 = v_6420 | ~v_6720;
assign v_30868 = v_6163 | v_30867;
assign v_30869 = v_6137 | ~v_6583;
assign v_30871 = v_6164 | v_30870;
assign v_30872 = v_6138 | ~v_6423;
assign v_30874 = v_5875 | v_30873;
assign v_30875 = v_5847 | ~v_6287;
assign v_30877 = v_5876 | v_30876;
assign v_30878 = v_5848 | ~v_6141;
assign v_30880 = v_5591 | v_30879;
assign v_30881 = v_5566 | ~v_6003;
assign v_30883 = v_5592 | v_30882;
assign v_30884 = v_5567 | ~v_5851;
assign v_30886 = v_5293 | v_30885;
assign v_30887 = v_5253 | ~v_5715;
assign v_30889 = v_5294 | v_30888;
assign v_30890 = v_5254 | ~v_5570;
assign v_30892 = v_4997 | v_30891;
assign v_30893 = v_4969 | ~v_5433;
assign v_30895 = v_4998 | v_30894;
assign v_30896 = v_4970 | ~v_5257;
assign v_30898 = v_4705 | v_30897;
assign v_30899 = v_4677 | ~v_5121;
assign v_30901 = v_4706 | v_30900;
assign v_30902 = v_4678 | ~v_4973;
assign v_30904 = v_4421 | v_30903;
assign v_30905 = v_4396 | ~v_4833;
assign v_30907 = v_4422 | v_30906;
assign v_30908 = v_4397 | ~v_4681;
assign v_30910 = v_4131 | v_30909;
assign v_30911 = v_4099 | ~v_4545;
assign v_30913 = v_4132 | v_30912;
assign v_30914 = v_4100 | ~v_4400;
assign v_30916 = v_3843 | v_30915;
assign v_30917 = v_3817 | ~v_4263;
assign v_30919 = v_3844 | v_30918;
assign v_30920 = v_3818 | ~v_4103;
assign v_30922 = v_3555 | v_30921;
assign v_30923 = v_3527 | ~v_3967;
assign v_30925 = v_3556 | v_30924;
assign v_30926 = v_3528 | ~v_3821;
assign v_30928 = v_3271 | v_30927;
assign v_30929 = v_3246 | ~v_3683;
assign v_30931 = v_3272 | v_30930;
assign v_30932 = v_3247 | ~v_3531;
assign v_30934 = v_2977 | v_30933;
assign v_30935 = v_2941 | ~v_3395;
assign v_30937 = v_2978 | v_30936;
assign v_30938 = v_2942 | ~v_3250;
assign v_30940 = v_2685 | v_30939;
assign v_30941 = v_2658 | ~v_3113;
assign v_30943 = v_2686 | v_30942;
assign v_30944 = v_2659 | ~v_2945;
assign v_30946 = v_2395 | v_30945;
assign v_30947 = v_2367 | ~v_2809;
assign v_30949 = v_2396 | v_30948;
assign v_30950 = v_2368 | ~v_2662;
assign v_30952 = v_2111 | v_30951;
assign v_30953 = v_2086 | ~v_2523;
assign v_30955 = v_2112 | v_30954;
assign v_30956 = v_2087 | ~v_2371;
assign v_30958 = v_1821 | v_30957;
assign v_30959 = v_1789 | ~v_2235;
assign v_30961 = v_1822 | v_30960;
assign v_30962 = v_1790 | ~v_2090;
assign v_30964 = v_1533 | v_30963;
assign v_30965 = v_1507 | ~v_1953;
assign v_30967 = v_1534 | v_30966;
assign v_30968 = v_1508 | ~v_1793;
assign v_30970 = v_1245 | v_30969;
assign v_30971 = v_1217 | ~v_1657;
assign v_30973 = v_1246 | v_30972;
assign v_30974 = v_1218 | ~v_1511;
assign v_30976 = v_961 | v_30975;
assign v_30977 = v_936 | ~v_1373;
assign v_30979 = v_962 | v_30978;
assign v_30980 = v_937 | ~v_1221;
assign v_30982 = v_591 | v_30981;
assign v_30983 = v_92 | ~v_1085;
assign v_30985 = v_593 | v_30984;
assign v_30986 = v_94 | ~v_940;
assign v_30988 = v_823 | v_30987;
assign v_30989 = ~v_804 | v_806;
assign v_30992 = v_9336 | ~v_9796;
assign v_30993 = v_9308 | ~v_9664;
assign v_30995 = v_9051 | v_30994;
assign v_30996 = v_9026 | ~v_9506;
assign v_30998 = v_9052 | v_30997;
assign v_30999 = v_9027 | ~v_9374;
assign v_31001 = v_8761 | v_31000;
assign v_31002 = v_8729 | ~v_9218;
assign v_31004 = v_8762 | v_31003;
assign v_31005 = v_8730 | ~v_9086;
assign v_31007 = v_8473 | v_31006;
assign v_31008 = v_8447 | ~v_8936;
assign v_31010 = v_8474 | v_31009;
assign v_31011 = v_8448 | ~v_8804;
assign v_31013 = v_8185 | v_31012;
assign v_31014 = v_8157 | ~v_8640;
assign v_31016 = v_8186 | v_31015;
assign v_31017 = v_8158 | ~v_8508;
assign v_31019 = v_7901 | v_31018;
assign v_31020 = v_7876 | ~v_8356;
assign v_31022 = v_7902 | v_31021;
assign v_31023 = v_7877 | ~v_8224;
assign v_31025 = v_7607 | v_31024;
assign v_31026 = v_7571 | ~v_8068;
assign v_31028 = v_7608 | v_31027;
assign v_31029 = v_7572 | ~v_7936;
assign v_31031 = v_7315 | v_31030;
assign v_31032 = v_7288 | ~v_7786;
assign v_31034 = v_7316 | v_31033;
assign v_31035 = v_7289 | ~v_7654;
assign v_31037 = v_7025 | v_31036;
assign v_31038 = v_6997 | ~v_7482;
assign v_31040 = v_7026 | v_31039;
assign v_31041 = v_6998 | ~v_7350;
assign v_31043 = v_6741 | v_31042;
assign v_31044 = v_6716 | ~v_7196;
assign v_31046 = v_6742 | v_31045;
assign v_31047 = v_6717 | ~v_7064;
assign v_31049 = v_6451 | v_31048;
assign v_31050 = v_6419 | ~v_6908;
assign v_31052 = v_6452 | v_31051;
assign v_31053 = v_6420 | ~v_6776;
assign v_31055 = v_6163 | v_31054;
assign v_31056 = v_6137 | ~v_6626;
assign v_31058 = v_6164 | v_31057;
assign v_31059 = v_6138 | ~v_6494;
assign v_31061 = v_5875 | v_31060;
assign v_31062 = v_5847 | ~v_6330;
assign v_31064 = v_5876 | v_31063;
assign v_31065 = v_5848 | ~v_6198;
assign v_31067 = v_5591 | v_31066;
assign v_31068 = v_5566 | ~v_6046;
assign v_31070 = v_5592 | v_31069;
assign v_31071 = v_5567 | ~v_5914;
assign v_31073 = v_5293 | v_31072;
assign v_31074 = v_5253 | ~v_5758;
assign v_31076 = v_5294 | v_31075;
assign v_31077 = v_5254 | ~v_5626;
assign v_31079 = v_4997 | v_31078;
assign v_31080 = v_4969 | ~v_5476;
assign v_31082 = v_4998 | v_31081;
assign v_31083 = v_4970 | ~v_5344;
assign v_31085 = v_4705 | v_31084;
assign v_31086 = v_4677 | ~v_5164;
assign v_31088 = v_4706 | v_31087;
assign v_31089 = v_4678 | ~v_5032;
assign v_31091 = v_4421 | v_31090;
assign v_31092 = v_4396 | ~v_4876;
assign v_31094 = v_4422 | v_31093;
assign v_31095 = v_4397 | ~v_4744;
assign v_31097 = v_4131 | v_31096;
assign v_31098 = v_4099 | ~v_4588;
assign v_31100 = v_4132 | v_31099;
assign v_31101 = v_4100 | ~v_4456;
assign v_31103 = v_3843 | v_31102;
assign v_31104 = v_3817 | ~v_4306;
assign v_31106 = v_3844 | v_31105;
assign v_31107 = v_3818 | ~v_4174;
assign v_31109 = v_3555 | v_31108;
assign v_31110 = v_3527 | ~v_4010;
assign v_31112 = v_3556 | v_31111;
assign v_31113 = v_3528 | ~v_3878;
assign v_31115 = v_3271 | v_31114;
assign v_31116 = v_3246 | ~v_3726;
assign v_31118 = v_3272 | v_31117;
assign v_31119 = v_3247 | ~v_3594;
assign v_31121 = v_2977 | v_31120;
assign v_31122 = v_2941 | ~v_3438;
assign v_31124 = v_2978 | v_31123;
assign v_31125 = v_2942 | ~v_3306;
assign v_31127 = v_2685 | v_31126;
assign v_31128 = v_2658 | ~v_3156;
assign v_31130 = v_2686 | v_31129;
assign v_31131 = v_2659 | ~v_3024;
assign v_31133 = v_2395 | v_31132;
assign v_31134 = v_2367 | ~v_2852;
assign v_31136 = v_2396 | v_31135;
assign v_31137 = v_2368 | ~v_2720;
assign v_31139 = v_2111 | v_31138;
assign v_31140 = v_2086 | ~v_2566;
assign v_31142 = v_2112 | v_31141;
assign v_31143 = v_2087 | ~v_2434;
assign v_31145 = v_1821 | v_31144;
assign v_31146 = v_1789 | ~v_2278;
assign v_31148 = v_1822 | v_31147;
assign v_31149 = v_1790 | ~v_2146;
assign v_31151 = v_1533 | v_31150;
assign v_31152 = v_1507 | ~v_1996;
assign v_31154 = v_1534 | v_31153;
assign v_31155 = v_1508 | ~v_1864;
assign v_31157 = v_1245 | v_31156;
assign v_31158 = v_1217 | ~v_1700;
assign v_31160 = v_1246 | v_31159;
assign v_31161 = v_1218 | ~v_1568;
assign v_31163 = v_961 | v_31162;
assign v_31164 = v_936 | ~v_1416;
assign v_31166 = v_962 | v_31165;
assign v_31167 = v_937 | ~v_1284;
assign v_31169 = v_591 | v_31168;
assign v_31170 = v_92 | ~v_1128;
assign v_31172 = v_593 | v_31171;
assign v_31173 = v_94 | ~v_996;
assign v_31175 = v_823 | v_31174;
assign v_31176 = v_806 | ~v_850;
assign v_31179 = v_9336 | ~v_9808;
assign v_31180 = v_9308 | ~v_9676;
assign v_31182 = v_9051 | v_31181;
assign v_31183 = v_9026 | ~v_9518;
assign v_31185 = v_9052 | v_31184;
assign v_31186 = v_9027 | ~v_9386;
assign v_31188 = v_8761 | v_31187;
assign v_31189 = v_8729 | ~v_9230;
assign v_31191 = v_8762 | v_31190;
assign v_31192 = v_8730 | ~v_9098;
assign v_31194 = v_8473 | v_31193;
assign v_31195 = v_8447 | ~v_8948;
assign v_31197 = v_8474 | v_31196;
assign v_31198 = v_8448 | ~v_8816;
assign v_31200 = v_8185 | v_31199;
assign v_31201 = v_8157 | ~v_8652;
assign v_31203 = v_8186 | v_31202;
assign v_31204 = v_8158 | ~v_8520;
assign v_31206 = v_7901 | v_31205;
assign v_31207 = v_7876 | ~v_8368;
assign v_31209 = v_7902 | v_31208;
assign v_31210 = v_7877 | ~v_8236;
assign v_31212 = v_7607 | v_31211;
assign v_31213 = v_7571 | ~v_8080;
assign v_31215 = v_7608 | v_31214;
assign v_31216 = v_7572 | ~v_7948;
assign v_31218 = v_7315 | v_31217;
assign v_31219 = v_7288 | ~v_7798;
assign v_31221 = v_7316 | v_31220;
assign v_31222 = v_7289 | ~v_7666;
assign v_31224 = v_7025 | v_31223;
assign v_31225 = v_6997 | ~v_7494;
assign v_31227 = v_7026 | v_31226;
assign v_31228 = v_6998 | ~v_7362;
assign v_31230 = v_6741 | v_31229;
assign v_31231 = v_6716 | ~v_7208;
assign v_31233 = v_6742 | v_31232;
assign v_31234 = v_6717 | ~v_7076;
assign v_31236 = v_6451 | v_31235;
assign v_31237 = v_6419 | ~v_6920;
assign v_31239 = v_6452 | v_31238;
assign v_31240 = v_6420 | ~v_6788;
assign v_31242 = v_6163 | v_31241;
assign v_31243 = v_6137 | ~v_6638;
assign v_31245 = v_6164 | v_31244;
assign v_31246 = v_6138 | ~v_6506;
assign v_31248 = v_5875 | v_31247;
assign v_31249 = v_5847 | ~v_6342;
assign v_31251 = v_5876 | v_31250;
assign v_31252 = v_5848 | ~v_6210;
assign v_31254 = v_5591 | v_31253;
assign v_31255 = v_5566 | ~v_6058;
assign v_31257 = v_5592 | v_31256;
assign v_31258 = v_5567 | ~v_5926;
assign v_31260 = v_5293 | v_31259;
assign v_31261 = v_5253 | ~v_5770;
assign v_31263 = v_5294 | v_31262;
assign v_31264 = v_5254 | ~v_5638;
assign v_31266 = v_4997 | v_31265;
assign v_31267 = v_4969 | ~v_5488;
assign v_31269 = v_4998 | v_31268;
assign v_31270 = v_4970 | ~v_5356;
assign v_31272 = v_4705 | v_31271;
assign v_31273 = v_4677 | ~v_5176;
assign v_31275 = v_4706 | v_31274;
assign v_31276 = v_4678 | ~v_5044;
assign v_31278 = v_4421 | v_31277;
assign v_31279 = v_4396 | ~v_4888;
assign v_31281 = v_4422 | v_31280;
assign v_31282 = v_4397 | ~v_4756;
assign v_31284 = v_4131 | v_31283;
assign v_31285 = v_4099 | ~v_4600;
assign v_31287 = v_4132 | v_31286;
assign v_31288 = v_4100 | ~v_4468;
assign v_31290 = v_3843 | v_31289;
assign v_31291 = v_3817 | ~v_4318;
assign v_31293 = v_3844 | v_31292;
assign v_31294 = v_3818 | ~v_4186;
assign v_31296 = v_3555 | v_31295;
assign v_31297 = v_3527 | ~v_4022;
assign v_31299 = v_3556 | v_31298;
assign v_31300 = v_3528 | ~v_3890;
assign v_31302 = v_3271 | v_31301;
assign v_31303 = v_3246 | ~v_3738;
assign v_31305 = v_3272 | v_31304;
assign v_31306 = v_3247 | ~v_3606;
assign v_31308 = v_2977 | v_31307;
assign v_31309 = v_2941 | ~v_3450;
assign v_31311 = v_2978 | v_31310;
assign v_31312 = v_2942 | ~v_3318;
assign v_31314 = v_2685 | v_31313;
assign v_31315 = v_2658 | ~v_3168;
assign v_31317 = v_2686 | v_31316;
assign v_31318 = v_2659 | ~v_3036;
assign v_31320 = v_2395 | v_31319;
assign v_31321 = v_2367 | ~v_2864;
assign v_31323 = v_2396 | v_31322;
assign v_31324 = v_2368 | ~v_2732;
assign v_31326 = v_2111 | v_31325;
assign v_31327 = v_2086 | ~v_2578;
assign v_31329 = v_2112 | v_31328;
assign v_31330 = v_2087 | ~v_2446;
assign v_31332 = v_1821 | v_31331;
assign v_31333 = v_1789 | ~v_2290;
assign v_31335 = v_1822 | v_31334;
assign v_31336 = v_1790 | ~v_2158;
assign v_31338 = v_1533 | v_31337;
assign v_31339 = v_1507 | ~v_2008;
assign v_31341 = v_1534 | v_31340;
assign v_31342 = v_1508 | ~v_1876;
assign v_31344 = v_1245 | v_31343;
assign v_31345 = v_1217 | ~v_1712;
assign v_31347 = v_1246 | v_31346;
assign v_31348 = v_1218 | ~v_1580;
assign v_31350 = v_961 | v_31349;
assign v_31351 = v_936 | ~v_1428;
assign v_31353 = v_962 | v_31352;
assign v_31354 = v_937 | ~v_1296;
assign v_31356 = v_591 | v_31355;
assign v_31357 = v_92 | ~v_1140;
assign v_31359 = v_593 | v_31358;
assign v_31360 = v_94 | ~v_1008;
assign v_31362 = v_823 | v_31361;
assign v_31363 = v_806 | ~v_862;
assign v_31366 = v_9336 | ~v_9820;
assign v_31367 = v_9308 | ~v_9688;
assign v_31369 = v_9051 | v_31368;
assign v_31370 = v_9026 | ~v_9530;
assign v_31372 = v_9052 | v_31371;
assign v_31373 = v_9027 | ~v_9398;
assign v_31375 = v_8761 | v_31374;
assign v_31376 = v_8729 | ~v_9242;
assign v_31378 = v_8762 | v_31377;
assign v_31379 = v_8730 | ~v_9110;
assign v_31381 = v_8473 | v_31380;
assign v_31382 = v_8447 | ~v_8960;
assign v_31384 = v_8474 | v_31383;
assign v_31385 = v_8448 | ~v_8828;
assign v_31387 = v_8185 | v_31386;
assign v_31388 = v_8157 | ~v_8664;
assign v_31390 = v_8186 | v_31389;
assign v_31391 = v_8158 | ~v_8532;
assign v_31393 = v_7901 | v_31392;
assign v_31394 = v_7876 | ~v_8380;
assign v_31396 = v_7902 | v_31395;
assign v_31397 = v_7877 | ~v_8248;
assign v_31399 = v_7607 | v_31398;
assign v_31400 = v_7571 | ~v_8092;
assign v_31402 = v_7608 | v_31401;
assign v_31403 = v_7572 | ~v_7960;
assign v_31405 = v_7315 | v_31404;
assign v_31406 = v_7288 | ~v_7810;
assign v_31408 = v_7316 | v_31407;
assign v_31409 = v_7289 | ~v_7678;
assign v_31411 = v_7025 | v_31410;
assign v_31412 = v_6997 | ~v_7506;
assign v_31414 = v_7026 | v_31413;
assign v_31415 = v_6998 | ~v_7374;
assign v_31417 = v_6741 | v_31416;
assign v_31418 = v_6716 | ~v_7220;
assign v_31420 = v_6742 | v_31419;
assign v_31421 = v_6717 | ~v_7088;
assign v_31423 = v_6451 | v_31422;
assign v_31424 = v_6419 | ~v_6932;
assign v_31426 = v_6452 | v_31425;
assign v_31427 = v_6420 | ~v_6800;
assign v_31429 = v_6163 | v_31428;
assign v_31430 = v_6137 | ~v_6650;
assign v_31432 = v_6164 | v_31431;
assign v_31433 = v_6138 | ~v_6518;
assign v_31435 = v_5875 | v_31434;
assign v_31436 = v_5847 | ~v_6354;
assign v_31438 = v_5876 | v_31437;
assign v_31439 = v_5848 | ~v_6222;
assign v_31441 = v_5591 | v_31440;
assign v_31442 = v_5566 | ~v_6070;
assign v_31444 = v_5592 | v_31443;
assign v_31445 = v_5567 | ~v_5938;
assign v_31447 = v_5293 | v_31446;
assign v_31448 = v_5253 | ~v_5782;
assign v_31450 = v_5294 | v_31449;
assign v_31451 = v_5254 | ~v_5650;
assign v_31453 = v_4997 | v_31452;
assign v_31454 = v_4969 | ~v_5500;
assign v_31456 = v_4998 | v_31455;
assign v_31457 = v_4970 | ~v_5368;
assign v_31459 = v_4705 | v_31458;
assign v_31460 = v_4677 | ~v_5188;
assign v_31462 = v_4706 | v_31461;
assign v_31463 = v_4678 | ~v_5056;
assign v_31465 = v_4421 | v_31464;
assign v_31466 = v_4396 | ~v_4900;
assign v_31468 = v_4422 | v_31467;
assign v_31469 = v_4397 | ~v_4768;
assign v_31471 = v_4131 | v_31470;
assign v_31472 = v_4099 | ~v_4612;
assign v_31474 = v_4132 | v_31473;
assign v_31475 = v_4100 | ~v_4480;
assign v_31477 = v_3843 | v_31476;
assign v_31478 = v_3817 | ~v_4330;
assign v_31480 = v_3844 | v_31479;
assign v_31481 = v_3818 | ~v_4198;
assign v_31483 = v_3555 | v_31482;
assign v_31484 = v_3527 | ~v_4034;
assign v_31486 = v_3556 | v_31485;
assign v_31487 = v_3528 | ~v_3902;
assign v_31489 = v_3271 | v_31488;
assign v_31490 = v_3246 | ~v_3750;
assign v_31492 = v_3272 | v_31491;
assign v_31493 = v_3247 | ~v_3618;
assign v_31495 = v_2977 | v_31494;
assign v_31496 = v_2941 | ~v_3462;
assign v_31498 = v_2978 | v_31497;
assign v_31499 = v_2942 | ~v_3330;
assign v_31501 = v_2685 | v_31500;
assign v_31502 = v_2658 | ~v_3180;
assign v_31504 = v_2686 | v_31503;
assign v_31505 = v_2659 | ~v_3048;
assign v_31507 = v_2395 | v_31506;
assign v_31508 = v_2367 | ~v_2876;
assign v_31510 = v_2396 | v_31509;
assign v_31511 = v_2368 | ~v_2744;
assign v_31513 = v_2111 | v_31512;
assign v_31514 = v_2086 | ~v_2590;
assign v_31516 = v_2112 | v_31515;
assign v_31517 = v_2087 | ~v_2458;
assign v_31519 = v_1821 | v_31518;
assign v_31520 = v_1789 | ~v_2302;
assign v_31522 = v_1822 | v_31521;
assign v_31523 = v_1790 | ~v_2170;
assign v_31525 = v_1533 | v_31524;
assign v_31526 = v_1507 | ~v_2020;
assign v_31528 = v_1534 | v_31527;
assign v_31529 = v_1508 | ~v_1888;
assign v_31531 = v_1245 | v_31530;
assign v_31532 = v_1217 | ~v_1724;
assign v_31534 = v_1246 | v_31533;
assign v_31535 = v_1218 | ~v_1592;
assign v_31537 = v_961 | v_31536;
assign v_31538 = v_936 | ~v_1440;
assign v_31540 = v_962 | v_31539;
assign v_31541 = v_937 | ~v_1308;
assign v_31543 = v_591 | v_31542;
assign v_31544 = v_92 | ~v_1152;
assign v_31546 = v_593 | v_31545;
assign v_31547 = v_94 | ~v_1020;
assign v_31549 = v_823 | v_31548;
assign v_31550 = v_806 | ~v_874;
assign v_31553 = v_9336 | ~v_9832;
assign v_31554 = v_9308 | ~v_9700;
assign v_31556 = v_9051 | v_31555;
assign v_31557 = v_9026 | ~v_9542;
assign v_31559 = v_9052 | v_31558;
assign v_31560 = v_9027 | ~v_9410;
assign v_31562 = v_8761 | v_31561;
assign v_31563 = v_8729 | ~v_9254;
assign v_31565 = v_8762 | v_31564;
assign v_31566 = v_8730 | ~v_9122;
assign v_31568 = v_8473 | v_31567;
assign v_31569 = v_8447 | ~v_8972;
assign v_31571 = v_8474 | v_31570;
assign v_31572 = v_8448 | ~v_8840;
assign v_31574 = v_8185 | v_31573;
assign v_31575 = v_8157 | ~v_8676;
assign v_31577 = v_8186 | v_31576;
assign v_31578 = v_8158 | ~v_8544;
assign v_31580 = v_7901 | v_31579;
assign v_31581 = v_7876 | ~v_8392;
assign v_31583 = v_7902 | v_31582;
assign v_31584 = v_7877 | ~v_8260;
assign v_31586 = v_7607 | v_31585;
assign v_31587 = v_7571 | ~v_8104;
assign v_31589 = v_7608 | v_31588;
assign v_31590 = v_7572 | ~v_7972;
assign v_31592 = v_7315 | v_31591;
assign v_31593 = v_7288 | ~v_7822;
assign v_31595 = v_7316 | v_31594;
assign v_31596 = v_7289 | ~v_7690;
assign v_31598 = v_7025 | v_31597;
assign v_31599 = v_6997 | ~v_7518;
assign v_31601 = v_7026 | v_31600;
assign v_31602 = v_6998 | ~v_7386;
assign v_31604 = v_6741 | v_31603;
assign v_31605 = v_6716 | ~v_7232;
assign v_31607 = v_6742 | v_31606;
assign v_31608 = v_6717 | ~v_7100;
assign v_31610 = v_6451 | v_31609;
assign v_31611 = v_6419 | ~v_6944;
assign v_31613 = v_6452 | v_31612;
assign v_31614 = v_6420 | ~v_6812;
assign v_31616 = v_6163 | v_31615;
assign v_31617 = v_6137 | ~v_6662;
assign v_31619 = v_6164 | v_31618;
assign v_31620 = v_6138 | ~v_6530;
assign v_31622 = v_5875 | v_31621;
assign v_31623 = v_5847 | ~v_6366;
assign v_31625 = v_5876 | v_31624;
assign v_31626 = v_5848 | ~v_6234;
assign v_31628 = v_5591 | v_31627;
assign v_31629 = v_5566 | ~v_6082;
assign v_31631 = v_5592 | v_31630;
assign v_31632 = v_5567 | ~v_5950;
assign v_31634 = v_5293 | v_31633;
assign v_31635 = v_5253 | ~v_5794;
assign v_31637 = v_5294 | v_31636;
assign v_31638 = v_5254 | ~v_5662;
assign v_31640 = v_4997 | v_31639;
assign v_31641 = v_4969 | ~v_5512;
assign v_31643 = v_4998 | v_31642;
assign v_31644 = v_4970 | ~v_5380;
assign v_31646 = v_4705 | v_31645;
assign v_31647 = v_4677 | ~v_5200;
assign v_31649 = v_4706 | v_31648;
assign v_31650 = v_4678 | ~v_5068;
assign v_31652 = v_4421 | v_31651;
assign v_31653 = v_4396 | ~v_4912;
assign v_31655 = v_4422 | v_31654;
assign v_31656 = v_4397 | ~v_4780;
assign v_31658 = v_4131 | v_31657;
assign v_31659 = v_4099 | ~v_4624;
assign v_31661 = v_4132 | v_31660;
assign v_31662 = v_4100 | ~v_4492;
assign v_31664 = v_3843 | v_31663;
assign v_31665 = v_3817 | ~v_4342;
assign v_31667 = v_3844 | v_31666;
assign v_31668 = v_3818 | ~v_4210;
assign v_31670 = v_3555 | v_31669;
assign v_31671 = v_3527 | ~v_4046;
assign v_31673 = v_3556 | v_31672;
assign v_31674 = v_3528 | ~v_3914;
assign v_31676 = v_3271 | v_31675;
assign v_31677 = v_3246 | ~v_3762;
assign v_31679 = v_3272 | v_31678;
assign v_31680 = v_3247 | ~v_3630;
assign v_31682 = v_2977 | v_31681;
assign v_31683 = v_2941 | ~v_3474;
assign v_31685 = v_2978 | v_31684;
assign v_31686 = v_2942 | ~v_3342;
assign v_31688 = v_2685 | v_31687;
assign v_31689 = v_2658 | ~v_3192;
assign v_31691 = v_2686 | v_31690;
assign v_31692 = v_2659 | ~v_3060;
assign v_31694 = v_2395 | v_31693;
assign v_31695 = v_2367 | ~v_2888;
assign v_31697 = v_2396 | v_31696;
assign v_31698 = v_2368 | ~v_2756;
assign v_31700 = v_2111 | v_31699;
assign v_31701 = v_2086 | ~v_2602;
assign v_31703 = v_2112 | v_31702;
assign v_31704 = v_2087 | ~v_2470;
assign v_31706 = v_1821 | v_31705;
assign v_31707 = v_1789 | ~v_2314;
assign v_31709 = v_1822 | v_31708;
assign v_31710 = v_1790 | ~v_2182;
assign v_31712 = v_1533 | v_31711;
assign v_31713 = v_1507 | ~v_2032;
assign v_31715 = v_1534 | v_31714;
assign v_31716 = v_1508 | ~v_1900;
assign v_31718 = v_1245 | v_31717;
assign v_31719 = v_1217 | ~v_1736;
assign v_31721 = v_1246 | v_31720;
assign v_31722 = v_1218 | ~v_1604;
assign v_31724 = v_961 | v_31723;
assign v_31725 = v_936 | ~v_1452;
assign v_31727 = v_962 | v_31726;
assign v_31728 = v_937 | ~v_1320;
assign v_31730 = v_591 | v_31729;
assign v_31731 = v_92 | ~v_1164;
assign v_31733 = v_593 | v_31732;
assign v_31734 = v_94 | ~v_1032;
assign v_31736 = v_823 | v_31735;
assign v_31737 = v_806 | ~v_886;
assign v_31741 = v_9336 | v_9872;
assign v_31742 = v_9308 | v_9740;
assign v_31744 = v_9051 | v_31743;
assign v_31745 = v_9026 | v_9582;
assign v_31747 = v_9052 | v_31746;
assign v_31748 = v_9027 | v_9450;
assign v_31750 = v_8761 | v_31749;
assign v_31751 = v_8729 | v_9294;
assign v_31753 = v_8762 | v_31752;
assign v_31754 = v_8730 | v_9162;
assign v_31756 = v_8473 | v_31755;
assign v_31757 = v_8447 | v_9012;
assign v_31759 = v_8474 | v_31758;
assign v_31760 = v_8448 | v_8880;
assign v_31762 = v_8185 | v_31761;
assign v_31763 = v_8157 | v_8716;
assign v_31765 = v_8186 | v_31764;
assign v_31766 = v_8158 | v_8584;
assign v_31768 = v_7901 | v_31767;
assign v_31769 = v_7876 | ~v_8432;
assign v_31771 = v_7902 | v_31770;
assign v_31772 = v_7877 | ~v_8300;
assign v_31774 = v_7607 | v_31773;
assign v_31775 = v_7571 | ~v_8144;
assign v_31777 = v_7608 | v_31776;
assign v_31778 = v_7572 | v_8012;
assign v_31780 = v_7315 | v_31779;
assign v_31781 = v_7288 | v_7862;
assign v_31783 = v_7316 | v_31782;
assign v_31784 = v_7289 | v_7730;
assign v_31786 = v_7025 | v_31785;
assign v_31787 = v_6997 | v_7558;
assign v_31789 = v_7026 | v_31788;
assign v_31790 = v_6998 | v_7426;
assign v_31792 = v_6741 | v_31791;
assign v_31793 = v_6716 | ~v_7272;
assign v_31795 = v_6742 | v_31794;
assign v_31796 = v_6717 | v_7140;
assign v_31798 = v_6451 | v_31797;
assign v_31799 = v_6419 | ~v_6984;
assign v_31801 = v_6452 | v_31800;
assign v_31802 = v_6420 | ~v_6852;
assign v_31804 = v_6163 | v_31803;
assign v_31805 = v_6137 | ~v_6702;
assign v_31807 = v_6164 | v_31806;
assign v_31808 = v_6138 | v_6570;
assign v_31810 = v_5875 | v_31809;
assign v_31811 = v_5847 | v_6406;
assign v_31813 = v_5876 | v_31812;
assign v_31814 = v_5848 | ~v_6274;
assign v_31816 = v_5591 | v_31815;
assign v_31817 = v_5566 | ~v_6122;
assign v_31819 = v_5592 | v_31818;
assign v_31820 = v_5567 | ~v_5990;
assign v_31822 = v_5293 | v_31821;
assign v_31823 = v_5253 | ~v_5834;
assign v_31825 = v_5294 | v_31824;
assign v_31826 = v_5254 | ~v_5702;
assign v_31828 = v_4997 | v_31827;
assign v_31829 = v_4969 | ~v_5552;
assign v_31831 = v_4998 | v_31830;
assign v_31832 = v_4970 | v_5420;
assign v_31834 = v_4705 | v_31833;
assign v_31835 = v_4677 | v_5240;
assign v_31837 = v_4706 | v_31836;
assign v_31838 = v_4678 | ~v_5108;
assign v_31840 = v_4421 | v_31839;
assign v_31841 = v_4396 | ~v_4952;
assign v_31843 = v_4422 | v_31842;
assign v_31844 = v_4397 | ~v_4820;
assign v_31846 = v_4131 | v_31845;
assign v_31847 = v_4099 | ~v_4664;
assign v_31849 = v_4132 | v_31848;
assign v_31850 = v_4100 | ~v_4532;
assign v_31852 = v_3843 | v_31851;
assign v_31853 = v_3817 | ~v_4382;
assign v_31855 = v_3844 | v_31854;
assign v_31856 = v_3818 | v_4250;
assign v_31858 = v_3555 | v_31857;
assign v_31859 = v_3527 | v_4086;
assign v_31861 = v_3556 | v_31860;
assign v_31862 = v_3528 | v_3954;
assign v_31864 = v_3271 | v_31863;
assign v_31865 = v_3246 | v_3802;
assign v_31867 = v_3272 | v_31866;
assign v_31868 = v_3247 | v_3670;
assign v_31870 = v_2977 | v_31869;
assign v_31871 = v_2941 | ~v_3514;
assign v_31873 = v_2978 | v_31872;
assign v_31874 = v_2942 | v_3382;
assign v_31876 = v_2685 | v_31875;
assign v_31877 = v_2658 | ~v_3232;
assign v_31879 = v_2686 | v_31878;
assign v_31880 = v_2659 | v_3100;
assign v_31882 = v_2395 | v_31881;
assign v_31883 = v_2367 | v_2928;
assign v_31885 = v_2396 | v_31884;
assign v_31886 = v_2368 | v_2796;
assign v_31888 = v_2111 | v_31887;
assign v_31889 = v_2086 | v_2642;
assign v_31891 = v_2112 | v_31890;
assign v_31892 = v_2087 | v_2510;
assign v_31894 = v_1821 | v_31893;
assign v_31895 = v_1789 | ~v_2354;
assign v_31897 = v_1822 | v_31896;
assign v_31898 = v_1790 | ~v_2222;
assign v_31900 = v_1533 | v_31899;
assign v_31901 = v_1507 | ~v_2072;
assign v_31903 = v_1534 | v_31902;
assign v_31904 = v_1508 | v_1940;
assign v_31906 = v_1245 | v_31905;
assign v_31907 = v_1217 | v_1776;
assign v_31909 = v_1246 | v_31908;
assign v_31910 = v_1218 | v_1644;
assign v_31912 = v_961 | v_31911;
assign v_31913 = v_936 | v_1492;
assign v_31915 = v_962 | v_31914;
assign v_31916 = v_937 | v_1360;
assign v_31918 = v_591 | v_31917;
assign v_31919 = v_92 | v_1204;
assign v_31921 = v_593 | v_31920;
assign v_31922 = v_94 | v_1072;
assign v_31924 = v_823 | v_31923;
assign v_31925 = v_806 | v_922;
assign v_31931 = ~v_807 | v_31930;
assign v_31932 = v_9629 | ~v_9784;
assign v_31933 = v_9600 | ~v_9652;
assign v_31935 = v_9630 | v_31934;
assign v_31936 = ~v_9494 | v_9601;
assign v_31938 = v_9335 | v_31937;
assign v_31939 = v_9307 | ~v_9362;
assign v_31941 = v_9336 | v_31940;
assign v_31942 = ~v_9206 | v_9308;
assign v_31944 = v_9051 | v_31943;
assign v_31945 = v_9026 | ~v_9074;
assign v_31947 = v_9052 | v_31946;
assign v_31948 = ~v_8924 | v_9027;
assign v_31950 = v_8761 | v_31949;
assign v_31951 = v_8729 | ~v_8792;
assign v_31953 = v_8762 | v_31952;
assign v_31954 = ~v_8628 | v_8730;
assign v_31956 = v_8473 | v_31955;
assign v_31957 = v_8447 | ~v_8496;
assign v_31959 = v_8474 | v_31958;
assign v_31960 = ~v_8344 | v_8448;
assign v_31962 = v_8185 | v_31961;
assign v_31963 = v_8157 | ~v_8212;
assign v_31965 = v_8186 | v_31964;
assign v_31966 = ~v_8056 | v_8158;
assign v_31968 = v_7901 | v_31967;
assign v_31969 = v_7876 | ~v_7924;
assign v_31971 = v_7902 | v_31970;
assign v_31972 = ~v_7774 | v_7877;
assign v_31974 = v_7607 | v_31973;
assign v_31975 = v_7571 | ~v_7642;
assign v_31977 = v_7608 | v_31976;
assign v_31978 = ~v_7470 | v_7572;
assign v_31980 = v_7315 | v_31979;
assign v_31981 = v_7288 | ~v_7338;
assign v_31983 = v_7316 | v_31982;
assign v_31984 = ~v_7184 | v_7289;
assign v_31986 = v_7025 | v_31985;
assign v_31987 = v_6997 | ~v_7052;
assign v_31989 = v_7026 | v_31988;
assign v_31990 = ~v_6896 | v_6998;
assign v_31992 = v_6741 | v_31991;
assign v_31993 = v_6716 | ~v_6764;
assign v_31995 = v_6742 | v_31994;
assign v_31996 = ~v_6614 | v_6717;
assign v_31998 = v_6451 | v_31997;
assign v_31999 = v_6419 | ~v_6482;
assign v_32001 = v_6452 | v_32000;
assign v_32002 = ~v_6318 | v_6420;
assign v_32004 = v_6163 | v_32003;
assign v_32005 = v_6137 | ~v_6186;
assign v_32007 = v_6164 | v_32006;
assign v_32008 = ~v_6034 | v_6138;
assign v_32010 = v_5875 | v_32009;
assign v_32011 = v_5847 | ~v_5902;
assign v_32013 = v_5876 | v_32012;
assign v_32014 = ~v_5746 | v_5848;
assign v_32016 = v_5591 | v_32015;
assign v_32017 = v_5566 | ~v_5614;
assign v_32019 = v_5592 | v_32018;
assign v_32020 = ~v_5464 | v_5567;
assign v_32022 = v_5293 | v_32021;
assign v_32023 = v_5253 | ~v_5332;
assign v_32025 = v_5294 | v_32024;
assign v_32026 = ~v_5152 | v_5254;
assign v_32028 = v_4997 | v_32027;
assign v_32029 = v_4969 | ~v_5020;
assign v_32031 = v_4998 | v_32030;
assign v_32032 = ~v_4864 | v_4970;
assign v_32034 = v_4705 | v_32033;
assign v_32035 = v_4677 | ~v_4732;
assign v_32037 = v_4706 | v_32036;
assign v_32038 = ~v_4576 | v_4678;
assign v_32040 = v_4421 | v_32039;
assign v_32041 = v_4396 | ~v_4444;
assign v_32043 = v_4422 | v_32042;
assign v_32044 = ~v_4294 | v_4397;
assign v_32046 = v_4131 | v_32045;
assign v_32047 = v_4099 | ~v_4162;
assign v_32049 = v_4132 | v_32048;
assign v_32050 = ~v_3998 | v_4100;
assign v_32052 = v_3843 | v_32051;
assign v_32053 = v_3817 | ~v_3866;
assign v_32055 = v_3844 | v_32054;
assign v_32056 = ~v_3714 | v_3818;
assign v_32058 = v_3555 | v_32057;
assign v_32059 = v_3527 | ~v_3582;
assign v_32061 = v_3556 | v_32060;
assign v_32062 = ~v_3426 | v_3528;
assign v_32064 = v_3271 | v_32063;
assign v_32065 = v_3246 | ~v_3294;
assign v_32067 = v_3272 | v_32066;
assign v_32068 = ~v_3144 | v_3247;
assign v_32070 = v_2977 | v_32069;
assign v_32071 = v_2941 | ~v_3012;
assign v_32073 = v_2978 | v_32072;
assign v_32074 = ~v_2840 | v_2942;
assign v_32076 = v_2685 | v_32075;
assign v_32077 = v_2658 | ~v_2708;
assign v_32079 = v_2686 | v_32078;
assign v_32080 = ~v_2554 | v_2659;
assign v_32082 = v_2395 | v_32081;
assign v_32083 = v_2367 | ~v_2422;
assign v_32085 = v_2396 | v_32084;
assign v_32086 = ~v_2266 | v_2368;
assign v_32088 = v_2111 | v_32087;
assign v_32089 = v_2086 | ~v_2134;
assign v_32091 = v_2112 | v_32090;
assign v_32092 = ~v_1984 | v_2087;
assign v_32094 = v_1821 | v_32093;
assign v_32095 = v_1789 | ~v_1852;
assign v_32097 = v_1822 | v_32096;
assign v_32098 = ~v_1688 | v_1790;
assign v_32100 = v_1533 | v_32099;
assign v_32101 = v_1507 | ~v_1556;
assign v_32103 = v_1534 | v_32102;
assign v_32104 = ~v_1404 | v_1508;
assign v_32106 = v_1245 | v_32105;
assign v_32107 = v_1217 | ~v_1272;
assign v_32109 = v_1246 | v_32108;
assign v_32110 = ~v_1116 | v_1218;
assign v_32112 = v_961 | v_32111;
assign v_32113 = v_936 | ~v_984;
assign v_32115 = v_962 | v_32114;
assign v_32116 = ~v_838 | v_937;
assign v_32118 = v_591 | v_32117;
assign v_32119 = v_92 | ~v_721;
assign v_32121 = v_9629 | ~v_9753;
assign v_32122 = v_9600 | ~v_9604;
assign v_32124 = v_9630 | v_32123;
assign v_32125 = ~v_9463 | v_9601;
assign v_32127 = v_9335 | v_32126;
assign v_32128 = v_9307 | ~v_9311;
assign v_32130 = v_9336 | v_32129;
assign v_32131 = ~v_9175 | v_9308;
assign v_32133 = v_9051 | v_32132;
assign v_32134 = v_9026 | ~v_9030;
assign v_32136 = v_9052 | v_32135;
assign v_32137 = ~v_8893 | v_9027;
assign v_32139 = v_8761 | v_32138;
assign v_32140 = v_8729 | ~v_8733;
assign v_32142 = v_8762 | v_32141;
assign v_32143 = ~v_8597 | v_8730;
assign v_32145 = v_8473 | v_32144;
assign v_32146 = v_8447 | ~v_8451;
assign v_32148 = v_8474 | v_32147;
assign v_32149 = ~v_8313 | v_8448;
assign v_32151 = v_8185 | v_32150;
assign v_32152 = v_8157 | ~v_8161;
assign v_32154 = v_8186 | v_32153;
assign v_32155 = ~v_8025 | v_8158;
assign v_32157 = v_7901 | v_32156;
assign v_32158 = v_7876 | ~v_7880;
assign v_32160 = v_7902 | v_32159;
assign v_32161 = ~v_7743 | v_7877;
assign v_32163 = v_7607 | v_32162;
assign v_32164 = v_7571 | ~v_7575;
assign v_32166 = v_7608 | v_32165;
assign v_32167 = ~v_7439 | v_7572;
assign v_32169 = v_7315 | v_32168;
assign v_32170 = v_7288 | ~v_7292;
assign v_32172 = v_7316 | v_32171;
assign v_32173 = ~v_7153 | v_7289;
assign v_32175 = v_7025 | v_32174;
assign v_32176 = v_6997 | ~v_7001;
assign v_32178 = v_7026 | v_32177;
assign v_32179 = ~v_6865 | v_6998;
assign v_32181 = v_6741 | v_32180;
assign v_32182 = v_6716 | ~v_6720;
assign v_32184 = v_6742 | v_32183;
assign v_32185 = ~v_6583 | v_6717;
assign v_32187 = v_6451 | v_32186;
assign v_32188 = v_6419 | ~v_6423;
assign v_32190 = v_6452 | v_32189;
assign v_32191 = ~v_6287 | v_6420;
assign v_32193 = v_6163 | v_32192;
assign v_32194 = v_6137 | ~v_6141;
assign v_32196 = v_6164 | v_32195;
assign v_32197 = ~v_6003 | v_6138;
assign v_32199 = v_5875 | v_32198;
assign v_32200 = v_5847 | ~v_5851;
assign v_32202 = v_5876 | v_32201;
assign v_32203 = ~v_5715 | v_5848;
assign v_32205 = v_5591 | v_32204;
assign v_32206 = v_5566 | ~v_5570;
assign v_32208 = v_5592 | v_32207;
assign v_32209 = ~v_5433 | v_5567;
assign v_32211 = v_5293 | v_32210;
assign v_32212 = v_5253 | ~v_5257;
assign v_32214 = v_5294 | v_32213;
assign v_32215 = ~v_5121 | v_5254;
assign v_32217 = v_4997 | v_32216;
assign v_32218 = v_4969 | ~v_4973;
assign v_32220 = v_4998 | v_32219;
assign v_32221 = ~v_4833 | v_4970;
assign v_32223 = v_4705 | v_32222;
assign v_32224 = v_4677 | ~v_4681;
assign v_32226 = v_4706 | v_32225;
assign v_32227 = ~v_4545 | v_4678;
assign v_32229 = v_4421 | v_32228;
assign v_32230 = v_4396 | ~v_4400;
assign v_32232 = v_4422 | v_32231;
assign v_32233 = ~v_4263 | v_4397;
assign v_32235 = v_4131 | v_32234;
assign v_32236 = v_4099 | ~v_4103;
assign v_32238 = v_4132 | v_32237;
assign v_32239 = ~v_3967 | v_4100;
assign v_32241 = v_3843 | v_32240;
assign v_32242 = v_3817 | ~v_3821;
assign v_32244 = v_3844 | v_32243;
assign v_32245 = ~v_3683 | v_3818;
assign v_32247 = v_3555 | v_32246;
assign v_32248 = v_3527 | ~v_3531;
assign v_32250 = v_3556 | v_32249;
assign v_32251 = ~v_3395 | v_3528;
assign v_32253 = v_3271 | v_32252;
assign v_32254 = v_3246 | ~v_3250;
assign v_32256 = v_3272 | v_32255;
assign v_32257 = ~v_3113 | v_3247;
assign v_32259 = v_2977 | v_32258;
assign v_32260 = v_2941 | ~v_2945;
assign v_32262 = v_2978 | v_32261;
assign v_32263 = ~v_2809 | v_2942;
assign v_32265 = v_2685 | v_32264;
assign v_32266 = v_2658 | ~v_2662;
assign v_32268 = v_2686 | v_32267;
assign v_32269 = ~v_2523 | v_2659;
assign v_32271 = v_2395 | v_32270;
assign v_32272 = v_2367 | ~v_2371;
assign v_32274 = v_2396 | v_32273;
assign v_32275 = ~v_2235 | v_2368;
assign v_32277 = v_2111 | v_32276;
assign v_32278 = v_2086 | ~v_2090;
assign v_32280 = v_2112 | v_32279;
assign v_32281 = ~v_1953 | v_2087;
assign v_32283 = v_1821 | v_32282;
assign v_32284 = v_1789 | ~v_1793;
assign v_32286 = v_1822 | v_32285;
assign v_32287 = ~v_1657 | v_1790;
assign v_32289 = v_1533 | v_32288;
assign v_32290 = v_1507 | ~v_1511;
assign v_32292 = v_1534 | v_32291;
assign v_32293 = ~v_1373 | v_1508;
assign v_32295 = v_1245 | v_32294;
assign v_32296 = v_1217 | ~v_1221;
assign v_32298 = v_1246 | v_32297;
assign v_32299 = ~v_1085 | v_1218;
assign v_32301 = v_961 | v_32300;
assign v_32302 = v_936 | ~v_940;
assign v_32304 = v_962 | v_32303;
assign v_32305 = ~v_804 | v_937;
assign v_32307 = v_591 | v_32306;
assign v_32308 = v_92 | ~v_98;
assign v_32311 = v_9629 | ~v_9796;
assign v_32312 = v_9600 | ~v_9664;
assign v_32314 = v_9630 | v_32313;
assign v_32315 = ~v_9506 | v_9601;
assign v_32317 = v_9335 | v_32316;
assign v_32318 = v_9307 | ~v_9374;
assign v_32320 = v_9336 | v_32319;
assign v_32321 = ~v_9218 | v_9308;
assign v_32323 = v_9051 | v_32322;
assign v_32324 = v_9026 | ~v_9086;
assign v_32326 = v_9052 | v_32325;
assign v_32327 = ~v_8936 | v_9027;
assign v_32329 = v_8761 | v_32328;
assign v_32330 = v_8729 | ~v_8804;
assign v_32332 = v_8762 | v_32331;
assign v_32333 = ~v_8640 | v_8730;
assign v_32335 = v_8473 | v_32334;
assign v_32336 = v_8447 | ~v_8508;
assign v_32338 = v_8474 | v_32337;
assign v_32339 = ~v_8356 | v_8448;
assign v_32341 = v_8185 | v_32340;
assign v_32342 = v_8157 | ~v_8224;
assign v_32344 = v_8186 | v_32343;
assign v_32345 = ~v_8068 | v_8158;
assign v_32347 = v_7901 | v_32346;
assign v_32348 = v_7876 | ~v_7936;
assign v_32350 = v_7902 | v_32349;
assign v_32351 = ~v_7786 | v_7877;
assign v_32353 = v_7607 | v_32352;
assign v_32354 = v_7571 | ~v_7654;
assign v_32356 = v_7608 | v_32355;
assign v_32357 = ~v_7482 | v_7572;
assign v_32359 = v_7315 | v_32358;
assign v_32360 = v_7288 | ~v_7350;
assign v_32362 = v_7316 | v_32361;
assign v_32363 = ~v_7196 | v_7289;
assign v_32365 = v_7025 | v_32364;
assign v_32366 = v_6997 | ~v_7064;
assign v_32368 = v_7026 | v_32367;
assign v_32369 = ~v_6908 | v_6998;
assign v_32371 = v_6741 | v_32370;
assign v_32372 = v_6716 | ~v_6776;
assign v_32374 = v_6742 | v_32373;
assign v_32375 = ~v_6626 | v_6717;
assign v_32377 = v_6451 | v_32376;
assign v_32378 = v_6419 | ~v_6494;
assign v_32380 = v_6452 | v_32379;
assign v_32381 = ~v_6330 | v_6420;
assign v_32383 = v_6163 | v_32382;
assign v_32384 = v_6137 | ~v_6198;
assign v_32386 = v_6164 | v_32385;
assign v_32387 = ~v_6046 | v_6138;
assign v_32389 = v_5875 | v_32388;
assign v_32390 = v_5847 | ~v_5914;
assign v_32392 = v_5876 | v_32391;
assign v_32393 = ~v_5758 | v_5848;
assign v_32395 = v_5591 | v_32394;
assign v_32396 = v_5566 | ~v_5626;
assign v_32398 = v_5592 | v_32397;
assign v_32399 = ~v_5476 | v_5567;
assign v_32401 = v_5293 | v_32400;
assign v_32402 = v_5253 | ~v_5344;
assign v_32404 = v_5294 | v_32403;
assign v_32405 = ~v_5164 | v_5254;
assign v_32407 = v_4997 | v_32406;
assign v_32408 = v_4969 | ~v_5032;
assign v_32410 = v_4998 | v_32409;
assign v_32411 = ~v_4876 | v_4970;
assign v_32413 = v_4705 | v_32412;
assign v_32414 = v_4677 | ~v_4744;
assign v_32416 = v_4706 | v_32415;
assign v_32417 = ~v_4588 | v_4678;
assign v_32419 = v_4421 | v_32418;
assign v_32420 = v_4396 | ~v_4456;
assign v_32422 = v_4422 | v_32421;
assign v_32423 = ~v_4306 | v_4397;
assign v_32425 = v_4131 | v_32424;
assign v_32426 = v_4099 | ~v_4174;
assign v_32428 = v_4132 | v_32427;
assign v_32429 = ~v_4010 | v_4100;
assign v_32431 = v_3843 | v_32430;
assign v_32432 = v_3817 | ~v_3878;
assign v_32434 = v_3844 | v_32433;
assign v_32435 = ~v_3726 | v_3818;
assign v_32437 = v_3555 | v_32436;
assign v_32438 = v_3527 | ~v_3594;
assign v_32440 = v_3556 | v_32439;
assign v_32441 = ~v_3438 | v_3528;
assign v_32443 = v_3271 | v_32442;
assign v_32444 = v_3246 | ~v_3306;
assign v_32446 = v_3272 | v_32445;
assign v_32447 = ~v_3156 | v_3247;
assign v_32449 = v_2977 | v_32448;
assign v_32450 = v_2941 | ~v_3024;
assign v_32452 = v_2978 | v_32451;
assign v_32453 = ~v_2852 | v_2942;
assign v_32455 = v_2685 | v_32454;
assign v_32456 = v_2658 | ~v_2720;
assign v_32458 = v_2686 | v_32457;
assign v_32459 = ~v_2566 | v_2659;
assign v_32461 = v_2395 | v_32460;
assign v_32462 = v_2367 | ~v_2434;
assign v_32464 = v_2396 | v_32463;
assign v_32465 = ~v_2278 | v_2368;
assign v_32467 = v_2111 | v_32466;
assign v_32468 = v_2086 | ~v_2146;
assign v_32470 = v_2112 | v_32469;
assign v_32471 = ~v_1996 | v_2087;
assign v_32473 = v_1821 | v_32472;
assign v_32474 = v_1789 | ~v_1864;
assign v_32476 = v_1822 | v_32475;
assign v_32477 = ~v_1700 | v_1790;
assign v_32479 = v_1533 | v_32478;
assign v_32480 = v_1507 | ~v_1568;
assign v_32482 = v_1534 | v_32481;
assign v_32483 = ~v_1416 | v_1508;
assign v_32485 = v_1245 | v_32484;
assign v_32486 = v_1217 | ~v_1284;
assign v_32488 = v_1246 | v_32487;
assign v_32489 = ~v_1128 | v_1218;
assign v_32491 = v_961 | v_32490;
assign v_32492 = v_936 | ~v_996;
assign v_32494 = v_962 | v_32493;
assign v_32495 = ~v_850 | v_937;
assign v_32497 = v_591 | v_32496;
assign v_32498 = v_92 | ~v_731;
assign v_32501 = v_9629 | ~v_9808;
assign v_32502 = v_9600 | ~v_9676;
assign v_32504 = v_9630 | v_32503;
assign v_32505 = ~v_9518 | v_9601;
assign v_32507 = v_9335 | v_32506;
assign v_32508 = v_9307 | ~v_9386;
assign v_32510 = v_9336 | v_32509;
assign v_32511 = ~v_9230 | v_9308;
assign v_32513 = v_9051 | v_32512;
assign v_32514 = v_9026 | ~v_9098;
assign v_32516 = v_9052 | v_32515;
assign v_32517 = ~v_8948 | v_9027;
assign v_32519 = v_8761 | v_32518;
assign v_32520 = v_8729 | ~v_8816;
assign v_32522 = v_8762 | v_32521;
assign v_32523 = ~v_8652 | v_8730;
assign v_32525 = v_8473 | v_32524;
assign v_32526 = v_8447 | ~v_8520;
assign v_32528 = v_8474 | v_32527;
assign v_32529 = ~v_8368 | v_8448;
assign v_32531 = v_8185 | v_32530;
assign v_32532 = v_8157 | ~v_8236;
assign v_32534 = v_8186 | v_32533;
assign v_32535 = ~v_8080 | v_8158;
assign v_32537 = v_7901 | v_32536;
assign v_32538 = v_7876 | ~v_7948;
assign v_32540 = v_7902 | v_32539;
assign v_32541 = ~v_7798 | v_7877;
assign v_32543 = v_7607 | v_32542;
assign v_32544 = v_7571 | ~v_7666;
assign v_32546 = v_7608 | v_32545;
assign v_32547 = ~v_7494 | v_7572;
assign v_32549 = v_7315 | v_32548;
assign v_32550 = v_7288 | ~v_7362;
assign v_32552 = v_7316 | v_32551;
assign v_32553 = ~v_7208 | v_7289;
assign v_32555 = v_7025 | v_32554;
assign v_32556 = v_6997 | ~v_7076;
assign v_32558 = v_7026 | v_32557;
assign v_32559 = ~v_6920 | v_6998;
assign v_32561 = v_6741 | v_32560;
assign v_32562 = v_6716 | ~v_6788;
assign v_32564 = v_6742 | v_32563;
assign v_32565 = ~v_6638 | v_6717;
assign v_32567 = v_6451 | v_32566;
assign v_32568 = v_6419 | ~v_6506;
assign v_32570 = v_6452 | v_32569;
assign v_32571 = ~v_6342 | v_6420;
assign v_32573 = v_6163 | v_32572;
assign v_32574 = v_6137 | ~v_6210;
assign v_32576 = v_6164 | v_32575;
assign v_32577 = ~v_6058 | v_6138;
assign v_32579 = v_5875 | v_32578;
assign v_32580 = v_5847 | ~v_5926;
assign v_32582 = v_5876 | v_32581;
assign v_32583 = ~v_5770 | v_5848;
assign v_32585 = v_5591 | v_32584;
assign v_32586 = v_5566 | ~v_5638;
assign v_32588 = v_5592 | v_32587;
assign v_32589 = ~v_5488 | v_5567;
assign v_32591 = v_5293 | v_32590;
assign v_32592 = v_5253 | ~v_5356;
assign v_32594 = v_5294 | v_32593;
assign v_32595 = ~v_5176 | v_5254;
assign v_32597 = v_4997 | v_32596;
assign v_32598 = v_4969 | ~v_5044;
assign v_32600 = v_4998 | v_32599;
assign v_32601 = ~v_4888 | v_4970;
assign v_32603 = v_4705 | v_32602;
assign v_32604 = v_4677 | ~v_4756;
assign v_32606 = v_4706 | v_32605;
assign v_32607 = ~v_4600 | v_4678;
assign v_32609 = v_4421 | v_32608;
assign v_32610 = v_4396 | ~v_4468;
assign v_32612 = v_4422 | v_32611;
assign v_32613 = ~v_4318 | v_4397;
assign v_32615 = v_4131 | v_32614;
assign v_32616 = v_4099 | ~v_4186;
assign v_32618 = v_4132 | v_32617;
assign v_32619 = ~v_4022 | v_4100;
assign v_32621 = v_3843 | v_32620;
assign v_32622 = v_3817 | ~v_3890;
assign v_32624 = v_3844 | v_32623;
assign v_32625 = ~v_3738 | v_3818;
assign v_32627 = v_3555 | v_32626;
assign v_32628 = v_3527 | ~v_3606;
assign v_32630 = v_3556 | v_32629;
assign v_32631 = ~v_3450 | v_3528;
assign v_32633 = v_3271 | v_32632;
assign v_32634 = v_3246 | ~v_3318;
assign v_32636 = v_3272 | v_32635;
assign v_32637 = ~v_3168 | v_3247;
assign v_32639 = v_2977 | v_32638;
assign v_32640 = v_2941 | ~v_3036;
assign v_32642 = v_2978 | v_32641;
assign v_32643 = ~v_2864 | v_2942;
assign v_32645 = v_2685 | v_32644;
assign v_32646 = v_2658 | ~v_2732;
assign v_32648 = v_2686 | v_32647;
assign v_32649 = ~v_2578 | v_2659;
assign v_32651 = v_2395 | v_32650;
assign v_32652 = v_2367 | ~v_2446;
assign v_32654 = v_2396 | v_32653;
assign v_32655 = ~v_2290 | v_2368;
assign v_32657 = v_2111 | v_32656;
assign v_32658 = v_2086 | ~v_2158;
assign v_32660 = v_2112 | v_32659;
assign v_32661 = ~v_2008 | v_2087;
assign v_32663 = v_1821 | v_32662;
assign v_32664 = v_1789 | ~v_1876;
assign v_32666 = v_1822 | v_32665;
assign v_32667 = ~v_1712 | v_1790;
assign v_32669 = v_1533 | v_32668;
assign v_32670 = v_1507 | ~v_1580;
assign v_32672 = v_1534 | v_32671;
assign v_32673 = ~v_1428 | v_1508;
assign v_32675 = v_1245 | v_32674;
assign v_32676 = v_1217 | ~v_1296;
assign v_32678 = v_1246 | v_32677;
assign v_32679 = ~v_1140 | v_1218;
assign v_32681 = v_961 | v_32680;
assign v_32682 = v_936 | ~v_1008;
assign v_32684 = v_962 | v_32683;
assign v_32685 = ~v_862 | v_937;
assign v_32687 = v_591 | v_32686;
assign v_32688 = v_92 | ~v_741;
assign v_32691 = v_9629 | ~v_9820;
assign v_32692 = v_9600 | ~v_9688;
assign v_32694 = v_9630 | v_32693;
assign v_32695 = ~v_9530 | v_9601;
assign v_32697 = v_9335 | v_32696;
assign v_32698 = v_9307 | ~v_9398;
assign v_32700 = v_9336 | v_32699;
assign v_32701 = ~v_9242 | v_9308;
assign v_32703 = v_9051 | v_32702;
assign v_32704 = v_9026 | ~v_9110;
assign v_32706 = v_9052 | v_32705;
assign v_32707 = ~v_8960 | v_9027;
assign v_32709 = v_8761 | v_32708;
assign v_32710 = v_8729 | ~v_8828;
assign v_32712 = v_8762 | v_32711;
assign v_32713 = ~v_8664 | v_8730;
assign v_32715 = v_8473 | v_32714;
assign v_32716 = v_8447 | ~v_8532;
assign v_32718 = v_8474 | v_32717;
assign v_32719 = ~v_8380 | v_8448;
assign v_32721 = v_8185 | v_32720;
assign v_32722 = v_8157 | ~v_8248;
assign v_32724 = v_8186 | v_32723;
assign v_32725 = ~v_8092 | v_8158;
assign v_32727 = v_7901 | v_32726;
assign v_32728 = v_7876 | ~v_7960;
assign v_32730 = v_7902 | v_32729;
assign v_32731 = ~v_7810 | v_7877;
assign v_32733 = v_7607 | v_32732;
assign v_32734 = v_7571 | ~v_7678;
assign v_32736 = v_7608 | v_32735;
assign v_32737 = ~v_7506 | v_7572;
assign v_32739 = v_7315 | v_32738;
assign v_32740 = v_7288 | ~v_7374;
assign v_32742 = v_7316 | v_32741;
assign v_32743 = ~v_7220 | v_7289;
assign v_32745 = v_7025 | v_32744;
assign v_32746 = v_6997 | ~v_7088;
assign v_32748 = v_7026 | v_32747;
assign v_32749 = ~v_6932 | v_6998;
assign v_32751 = v_6741 | v_32750;
assign v_32752 = v_6716 | ~v_6800;
assign v_32754 = v_6742 | v_32753;
assign v_32755 = ~v_6650 | v_6717;
assign v_32757 = v_6451 | v_32756;
assign v_32758 = v_6419 | ~v_6518;
assign v_32760 = v_6452 | v_32759;
assign v_32761 = ~v_6354 | v_6420;
assign v_32763 = v_6163 | v_32762;
assign v_32764 = v_6137 | ~v_6222;
assign v_32766 = v_6164 | v_32765;
assign v_32767 = ~v_6070 | v_6138;
assign v_32769 = v_5875 | v_32768;
assign v_32770 = v_5847 | ~v_5938;
assign v_32772 = v_5876 | v_32771;
assign v_32773 = ~v_5782 | v_5848;
assign v_32775 = v_5591 | v_32774;
assign v_32776 = v_5566 | ~v_5650;
assign v_32778 = v_5592 | v_32777;
assign v_32779 = ~v_5500 | v_5567;
assign v_32781 = v_5293 | v_32780;
assign v_32782 = v_5253 | ~v_5368;
assign v_32784 = v_5294 | v_32783;
assign v_32785 = ~v_5188 | v_5254;
assign v_32787 = v_4997 | v_32786;
assign v_32788 = v_4969 | ~v_5056;
assign v_32790 = v_4998 | v_32789;
assign v_32791 = ~v_4900 | v_4970;
assign v_32793 = v_4705 | v_32792;
assign v_32794 = v_4677 | ~v_4768;
assign v_32796 = v_4706 | v_32795;
assign v_32797 = ~v_4612 | v_4678;
assign v_32799 = v_4421 | v_32798;
assign v_32800 = v_4396 | ~v_4480;
assign v_32802 = v_4422 | v_32801;
assign v_32803 = ~v_4330 | v_4397;
assign v_32805 = v_4131 | v_32804;
assign v_32806 = v_4099 | ~v_4198;
assign v_32808 = v_4132 | v_32807;
assign v_32809 = ~v_4034 | v_4100;
assign v_32811 = v_3843 | v_32810;
assign v_32812 = v_3817 | ~v_3902;
assign v_32814 = v_3844 | v_32813;
assign v_32815 = ~v_3750 | v_3818;
assign v_32817 = v_3555 | v_32816;
assign v_32818 = v_3527 | ~v_3618;
assign v_32820 = v_3556 | v_32819;
assign v_32821 = ~v_3462 | v_3528;
assign v_32823 = v_3271 | v_32822;
assign v_32824 = v_3246 | ~v_3330;
assign v_32826 = v_3272 | v_32825;
assign v_32827 = ~v_3180 | v_3247;
assign v_32829 = v_2977 | v_32828;
assign v_32830 = v_2941 | ~v_3048;
assign v_32832 = v_2978 | v_32831;
assign v_32833 = ~v_2876 | v_2942;
assign v_32835 = v_2685 | v_32834;
assign v_32836 = v_2658 | ~v_2744;
assign v_32838 = v_2686 | v_32837;
assign v_32839 = ~v_2590 | v_2659;
assign v_32841 = v_2395 | v_32840;
assign v_32842 = v_2367 | ~v_2458;
assign v_32844 = v_2396 | v_32843;
assign v_32845 = ~v_2302 | v_2368;
assign v_32847 = v_2111 | v_32846;
assign v_32848 = v_2086 | ~v_2170;
assign v_32850 = v_2112 | v_32849;
assign v_32851 = ~v_2020 | v_2087;
assign v_32853 = v_1821 | v_32852;
assign v_32854 = v_1789 | ~v_1888;
assign v_32856 = v_1822 | v_32855;
assign v_32857 = ~v_1724 | v_1790;
assign v_32859 = v_1533 | v_32858;
assign v_32860 = v_1507 | ~v_1592;
assign v_32862 = v_1534 | v_32861;
assign v_32863 = ~v_1440 | v_1508;
assign v_32865 = v_1245 | v_32864;
assign v_32866 = v_1217 | ~v_1308;
assign v_32868 = v_1246 | v_32867;
assign v_32869 = ~v_1152 | v_1218;
assign v_32871 = v_961 | v_32870;
assign v_32872 = v_936 | ~v_1020;
assign v_32874 = v_962 | v_32873;
assign v_32875 = ~v_874 | v_937;
assign v_32877 = v_591 | v_32876;
assign v_32878 = v_92 | ~v_751;
assign v_32881 = v_9629 | ~v_9832;
assign v_32882 = v_9600 | ~v_9700;
assign v_32884 = v_9630 | v_32883;
assign v_32885 = ~v_9542 | v_9601;
assign v_32887 = v_9335 | v_32886;
assign v_32888 = v_9307 | ~v_9410;
assign v_32890 = v_9336 | v_32889;
assign v_32891 = ~v_9254 | v_9308;
assign v_32893 = v_9051 | v_32892;
assign v_32894 = v_9026 | ~v_9122;
assign v_32896 = v_9052 | v_32895;
assign v_32897 = ~v_8972 | v_9027;
assign v_32899 = v_8761 | v_32898;
assign v_32900 = v_8729 | ~v_8840;
assign v_32902 = v_8762 | v_32901;
assign v_32903 = ~v_8676 | v_8730;
assign v_32905 = v_8473 | v_32904;
assign v_32906 = v_8447 | ~v_8544;
assign v_32908 = v_8474 | v_32907;
assign v_32909 = ~v_8392 | v_8448;
assign v_32911 = v_8185 | v_32910;
assign v_32912 = v_8157 | ~v_8260;
assign v_32914 = v_8186 | v_32913;
assign v_32915 = ~v_8104 | v_8158;
assign v_32917 = v_7901 | v_32916;
assign v_32918 = v_7876 | ~v_7972;
assign v_32920 = v_7902 | v_32919;
assign v_32921 = ~v_7822 | v_7877;
assign v_32923 = v_7607 | v_32922;
assign v_32924 = v_7571 | ~v_7690;
assign v_32926 = v_7608 | v_32925;
assign v_32927 = ~v_7518 | v_7572;
assign v_32929 = v_7315 | v_32928;
assign v_32930 = v_7288 | ~v_7386;
assign v_32932 = v_7316 | v_32931;
assign v_32933 = ~v_7232 | v_7289;
assign v_32935 = v_7025 | v_32934;
assign v_32936 = v_6997 | ~v_7100;
assign v_32938 = v_7026 | v_32937;
assign v_32939 = ~v_6944 | v_6998;
assign v_32941 = v_6741 | v_32940;
assign v_32942 = v_6716 | ~v_6812;
assign v_32944 = v_6742 | v_32943;
assign v_32945 = ~v_6662 | v_6717;
assign v_32947 = v_6451 | v_32946;
assign v_32948 = v_6419 | ~v_6530;
assign v_32950 = v_6452 | v_32949;
assign v_32951 = ~v_6366 | v_6420;
assign v_32953 = v_6163 | v_32952;
assign v_32954 = v_6137 | ~v_6234;
assign v_32956 = v_6164 | v_32955;
assign v_32957 = ~v_6082 | v_6138;
assign v_32959 = v_5875 | v_32958;
assign v_32960 = v_5847 | ~v_5950;
assign v_32962 = v_5876 | v_32961;
assign v_32963 = ~v_5794 | v_5848;
assign v_32965 = v_5591 | v_32964;
assign v_32966 = v_5566 | ~v_5662;
assign v_32968 = v_5592 | v_32967;
assign v_32969 = ~v_5512 | v_5567;
assign v_32971 = v_5293 | v_32970;
assign v_32972 = v_5253 | ~v_5380;
assign v_32974 = v_5294 | v_32973;
assign v_32975 = ~v_5200 | v_5254;
assign v_32977 = v_4997 | v_32976;
assign v_32978 = v_4969 | ~v_5068;
assign v_32980 = v_4998 | v_32979;
assign v_32981 = ~v_4912 | v_4970;
assign v_32983 = v_4705 | v_32982;
assign v_32984 = v_4677 | ~v_4780;
assign v_32986 = v_4706 | v_32985;
assign v_32987 = ~v_4624 | v_4678;
assign v_32989 = v_4421 | v_32988;
assign v_32990 = v_4396 | ~v_4492;
assign v_32992 = v_4422 | v_32991;
assign v_32993 = ~v_4342 | v_4397;
assign v_32995 = v_4131 | v_32994;
assign v_32996 = v_4099 | ~v_4210;
assign v_32998 = v_4132 | v_32997;
assign v_32999 = ~v_4046 | v_4100;
assign v_33001 = v_3843 | v_33000;
assign v_33002 = v_3817 | ~v_3914;
assign v_33004 = v_3844 | v_33003;
assign v_33005 = ~v_3762 | v_3818;
assign v_33007 = v_3555 | v_33006;
assign v_33008 = v_3527 | ~v_3630;
assign v_33010 = v_3556 | v_33009;
assign v_33011 = ~v_3474 | v_3528;
assign v_33013 = v_3271 | v_33012;
assign v_33014 = v_3246 | ~v_3342;
assign v_33016 = v_3272 | v_33015;
assign v_33017 = ~v_3192 | v_3247;
assign v_33019 = v_2977 | v_33018;
assign v_33020 = v_2941 | ~v_3060;
assign v_33022 = v_2978 | v_33021;
assign v_33023 = ~v_2888 | v_2942;
assign v_33025 = v_2685 | v_33024;
assign v_33026 = v_2658 | ~v_2756;
assign v_33028 = v_2686 | v_33027;
assign v_33029 = ~v_2602 | v_2659;
assign v_33031 = v_2395 | v_33030;
assign v_33032 = v_2367 | ~v_2470;
assign v_33034 = v_2396 | v_33033;
assign v_33035 = ~v_2314 | v_2368;
assign v_33037 = v_2111 | v_33036;
assign v_33038 = v_2086 | ~v_2182;
assign v_33040 = v_2112 | v_33039;
assign v_33041 = ~v_2032 | v_2087;
assign v_33043 = v_1821 | v_33042;
assign v_33044 = v_1789 | ~v_1900;
assign v_33046 = v_1822 | v_33045;
assign v_33047 = ~v_1736 | v_1790;
assign v_33049 = v_1533 | v_33048;
assign v_33050 = v_1507 | ~v_1604;
assign v_33052 = v_1534 | v_33051;
assign v_33053 = ~v_1452 | v_1508;
assign v_33055 = v_1245 | v_33054;
assign v_33056 = v_1217 | ~v_1320;
assign v_33058 = v_1246 | v_33057;
assign v_33059 = ~v_1164 | v_1218;
assign v_33061 = v_961 | v_33060;
assign v_33062 = v_936 | ~v_1032;
assign v_33064 = v_962 | v_33063;
assign v_33065 = ~v_886 | v_937;
assign v_33067 = v_591 | v_33066;
assign v_33068 = v_92 | ~v_761;
assign v_33071 = v_9629 | ~v_9844;
assign v_33072 = v_9600 | ~v_9712;
assign v_33074 = v_9630 | v_33073;
assign v_33075 = ~v_9554 | v_9601;
assign v_33077 = v_9335 | v_33076;
assign v_33078 = v_9307 | ~v_9422;
assign v_33080 = v_9336 | v_33079;
assign v_33081 = ~v_9266 | v_9308;
assign v_33083 = v_9051 | v_33082;
assign v_33084 = v_9026 | ~v_9134;
assign v_33086 = v_9052 | v_33085;
assign v_33087 = ~v_8984 | v_9027;
assign v_33089 = v_8761 | v_33088;
assign v_33090 = v_8729 | ~v_8852;
assign v_33092 = v_8762 | v_33091;
assign v_33093 = ~v_8688 | v_8730;
assign v_33095 = v_8473 | v_33094;
assign v_33096 = v_8447 | ~v_8556;
assign v_33098 = v_8474 | v_33097;
assign v_33099 = ~v_8404 | v_8448;
assign v_33101 = v_8185 | v_33100;
assign v_33102 = v_8157 | ~v_8272;
assign v_33104 = v_8186 | v_33103;
assign v_33105 = ~v_8116 | v_8158;
assign v_33107 = v_7901 | v_33106;
assign v_33108 = v_7876 | ~v_7984;
assign v_33110 = v_7902 | v_33109;
assign v_33111 = ~v_7834 | v_7877;
assign v_33113 = v_7607 | v_33112;
assign v_33114 = v_7571 | ~v_7702;
assign v_33116 = v_7608 | v_33115;
assign v_33117 = ~v_7530 | v_7572;
assign v_33119 = v_7315 | v_33118;
assign v_33120 = v_7288 | ~v_7398;
assign v_33122 = v_7316 | v_33121;
assign v_33123 = ~v_7244 | v_7289;
assign v_33125 = v_7025 | v_33124;
assign v_33126 = v_6997 | ~v_7112;
assign v_33128 = v_7026 | v_33127;
assign v_33129 = ~v_6956 | v_6998;
assign v_33131 = v_6741 | v_33130;
assign v_33132 = v_6716 | v_6824;
assign v_33134 = v_6742 | v_33133;
assign v_33135 = ~v_6674 | v_6717;
assign v_33137 = v_6451 | v_33136;
assign v_33138 = v_6419 | ~v_6542;
assign v_33140 = v_6452 | v_33139;
assign v_33141 = ~v_6378 | v_6420;
assign v_33143 = v_6163 | v_33142;
assign v_33144 = v_6137 | ~v_6246;
assign v_33146 = v_6164 | v_33145;
assign v_33147 = v_6094 | v_6138;
assign v_33149 = v_5875 | v_33148;
assign v_33150 = v_5847 | ~v_5962;
assign v_33152 = v_5876 | v_33151;
assign v_33153 = v_5806 | v_5848;
assign v_33155 = v_5591 | v_33154;
assign v_33156 = v_5566 | ~v_5674;
assign v_33158 = v_5592 | v_33157;
assign v_33159 = ~v_5524 | v_5567;
assign v_33161 = v_5293 | v_33160;
assign v_33162 = v_5253 | ~v_5392;
assign v_33164 = v_5294 | v_33163;
assign v_33165 = ~v_5212 | v_5254;
assign v_33167 = v_4997 | v_33166;
assign v_33168 = v_4969 | ~v_5080;
assign v_33170 = v_4998 | v_33169;
assign v_33171 = ~v_4924 | v_4970;
assign v_33173 = v_4705 | v_33172;
assign v_33174 = v_4677 | ~v_4792;
assign v_33176 = v_4706 | v_33175;
assign v_33177 = ~v_4636 | v_4678;
assign v_33179 = v_4421 | v_33178;
assign v_33180 = v_4396 | ~v_4504;
assign v_33182 = v_4422 | v_33181;
assign v_33183 = ~v_4354 | v_4397;
assign v_33185 = v_4131 | v_33184;
assign v_33186 = v_4099 | ~v_4222;
assign v_33188 = v_4132 | v_33187;
assign v_33189 = ~v_4058 | v_4100;
assign v_33191 = v_3843 | v_33190;
assign v_33192 = v_3817 | ~v_3926;
assign v_33194 = v_3844 | v_33193;
assign v_33195 = ~v_3774 | v_3818;
assign v_33197 = v_3555 | v_33196;
assign v_33198 = v_3527 | ~v_3642;
assign v_33200 = v_3556 | v_33199;
assign v_33201 = ~v_3486 | v_3528;
assign v_33203 = v_3271 | v_33202;
assign v_33204 = v_3246 | ~v_3354;
assign v_33206 = v_3272 | v_33205;
assign v_33207 = v_3204 | v_3247;
assign v_33209 = v_2977 | v_33208;
assign v_33210 = v_2941 | ~v_3072;
assign v_33212 = v_2978 | v_33211;
assign v_33213 = ~v_2900 | v_2942;
assign v_33215 = v_2685 | v_33214;
assign v_33216 = v_2658 | ~v_2768;
assign v_33218 = v_2686 | v_33217;
assign v_33219 = ~v_2614 | v_2659;
assign v_33221 = v_2395 | v_33220;
assign v_33222 = v_2367 | ~v_2482;
assign v_33224 = v_2396 | v_33223;
assign v_33225 = ~v_2326 | v_2368;
assign v_33227 = v_2111 | v_33226;
assign v_33228 = v_2086 | ~v_2194;
assign v_33230 = v_2112 | v_33229;
assign v_33231 = ~v_2044 | v_2087;
assign v_33233 = v_1821 | v_33232;
assign v_33234 = v_1789 | ~v_1912;
assign v_33236 = v_1822 | v_33235;
assign v_33237 = ~v_1748 | v_1790;
assign v_33239 = v_1533 | v_33238;
assign v_33240 = v_1507 | ~v_1616;
assign v_33242 = v_1534 | v_33241;
assign v_33243 = ~v_1464 | v_1508;
assign v_33245 = v_1245 | v_33244;
assign v_33246 = v_1217 | ~v_1332;
assign v_33248 = v_1246 | v_33247;
assign v_33249 = ~v_1176 | v_1218;
assign v_33251 = v_961 | v_33250;
assign v_33252 = v_936 | ~v_1044;
assign v_33254 = v_962 | v_33253;
assign v_33255 = ~v_898 | v_937;
assign v_33257 = v_591 | v_33256;
assign v_33258 = v_92 | ~v_771;
assign v_33261 = v_9629 | v_9872;
assign v_33262 = v_9600 | v_9740;
assign v_33264 = v_9630 | v_33263;
assign v_33265 = v_9582 | v_9601;
assign v_33267 = v_9335 | v_33266;
assign v_33268 = v_9307 | v_9450;
assign v_33270 = v_9336 | v_33269;
assign v_33271 = v_9294 | v_9308;
assign v_33273 = v_9051 | v_33272;
assign v_33274 = v_9026 | v_9162;
assign v_33276 = v_9052 | v_33275;
assign v_33277 = v_9012 | v_9027;
assign v_33279 = v_8761 | v_33278;
assign v_33280 = v_8729 | v_8880;
assign v_33282 = v_8762 | v_33281;
assign v_33283 = v_8716 | v_8730;
assign v_33285 = v_8473 | v_33284;
assign v_33286 = v_8447 | v_8584;
assign v_33288 = v_8474 | v_33287;
assign v_33289 = ~v_8432 | v_8448;
assign v_33291 = v_8185 | v_33290;
assign v_33292 = v_8157 | ~v_8300;
assign v_33294 = v_8186 | v_33293;
assign v_33295 = ~v_8144 | v_8158;
assign v_33297 = v_7901 | v_33296;
assign v_33298 = v_7876 | v_8012;
assign v_33300 = v_7902 | v_33299;
assign v_33301 = v_7862 | v_7877;
assign v_33303 = v_7607 | v_33302;
assign v_33304 = v_7571 | v_7730;
assign v_33306 = v_7608 | v_33305;
assign v_33307 = v_7558 | v_7572;
assign v_33309 = v_7315 | v_33308;
assign v_33310 = v_7288 | v_7426;
assign v_33312 = v_7316 | v_33311;
assign v_33313 = ~v_7272 | v_7289;
assign v_33315 = v_7025 | v_33314;
assign v_33316 = v_6997 | v_7140;
assign v_33318 = v_7026 | v_33317;
assign v_33319 = ~v_6984 | v_6998;
assign v_33321 = v_6741 | v_33320;
assign v_33322 = v_6716 | ~v_6852;
assign v_33324 = v_6742 | v_33323;
assign v_33325 = ~v_6702 | v_6717;
assign v_33327 = v_6451 | v_33326;
assign v_33328 = v_6419 | v_6570;
assign v_33330 = v_6452 | v_33329;
assign v_33331 = v_6406 | v_6420;
assign v_33333 = v_6163 | v_33332;
assign v_33334 = v_6137 | ~v_6274;
assign v_33336 = v_6164 | v_33335;
assign v_33337 = ~v_6122 | v_6138;
assign v_33339 = v_5875 | v_33338;
assign v_33340 = v_5847 | ~v_5990;
assign v_33342 = v_5876 | v_33341;
assign v_33343 = ~v_5834 | v_5848;
assign v_33345 = v_5591 | v_33344;
assign v_33346 = v_5566 | ~v_5702;
assign v_33348 = v_5592 | v_33347;
assign v_33349 = ~v_5552 | v_5567;
assign v_33351 = v_5293 | v_33350;
assign v_33352 = v_5253 | v_5420;
assign v_33354 = v_5294 | v_33353;
assign v_33355 = v_5240 | v_5254;
assign v_33357 = v_4997 | v_33356;
assign v_33358 = v_4969 | ~v_5108;
assign v_33360 = v_4998 | v_33359;
assign v_33361 = ~v_4952 | v_4970;
assign v_33363 = v_4705 | v_33362;
assign v_33364 = v_4677 | ~v_4820;
assign v_33366 = v_4706 | v_33365;
assign v_33367 = ~v_4664 | v_4678;
assign v_33369 = v_4421 | v_33368;
assign v_33370 = v_4396 | ~v_4532;
assign v_33372 = v_4422 | v_33371;
assign v_33373 = ~v_4382 | v_4397;
assign v_33375 = v_4131 | v_33374;
assign v_33376 = v_4099 | v_4250;
assign v_33378 = v_4132 | v_33377;
assign v_33379 = v_4086 | v_4100;
assign v_33381 = v_3843 | v_33380;
assign v_33382 = v_3817 | v_3954;
assign v_33384 = v_3844 | v_33383;
assign v_33385 = v_3802 | v_3818;
assign v_33387 = v_3555 | v_33386;
assign v_33388 = v_3527 | v_3670;
assign v_33390 = v_3556 | v_33389;
assign v_33391 = ~v_3514 | v_3528;
assign v_33393 = v_3271 | v_33392;
assign v_33394 = v_3246 | v_3382;
assign v_33396 = v_3272 | v_33395;
assign v_33397 = ~v_3232 | v_3247;
assign v_33399 = v_2977 | v_33398;
assign v_33400 = v_2941 | v_3100;
assign v_33402 = v_2978 | v_33401;
assign v_33403 = v_2928 | v_2942;
assign v_33405 = v_2685 | v_33404;
assign v_33406 = v_2658 | v_2796;
assign v_33408 = v_2686 | v_33407;
assign v_33409 = v_2642 | v_2659;
assign v_33411 = v_2395 | v_33410;
assign v_33412 = v_2367 | v_2510;
assign v_33414 = v_2396 | v_33413;
assign v_33415 = ~v_2354 | v_2368;
assign v_33417 = v_2111 | v_33416;
assign v_33418 = v_2086 | ~v_2222;
assign v_33420 = v_2112 | v_33419;
assign v_33421 = ~v_2072 | v_2087;
assign v_33423 = v_1821 | v_33422;
assign v_33424 = v_1789 | v_1940;
assign v_33426 = v_1822 | v_33425;
assign v_33427 = v_1776 | v_1790;
assign v_33429 = v_1533 | v_33428;
assign v_33430 = v_1507 | v_1644;
assign v_33432 = v_1534 | v_33431;
assign v_33433 = v_1492 | v_1508;
assign v_33435 = v_1245 | v_33434;
assign v_33436 = v_1217 | v_1360;
assign v_33438 = v_1246 | v_33437;
assign v_33439 = v_1204 | v_1218;
assign v_33441 = v_961 | v_33440;
assign v_33442 = v_936 | v_1072;
assign v_33444 = v_962 | v_33443;
assign v_33445 = v_922 | v_937;
assign v_33447 = v_591 | v_33446;
assign v_33448 = v_92 | v_793;
assign v_33451 = v_9630 | ~v_9784;
assign v_33452 = v_9601 | ~v_9652;
assign v_33454 = v_9335 | v_33453;
assign v_33455 = v_9307 | ~v_9494;
assign v_33457 = v_9336 | v_33456;
assign v_33458 = v_9308 | ~v_9362;
assign v_33460 = v_9051 | v_33459;
assign v_33461 = v_9026 | ~v_9206;
assign v_33463 = v_9052 | v_33462;
assign v_33464 = v_9027 | ~v_9074;
assign v_33466 = v_8761 | v_33465;
assign v_33467 = v_8729 | ~v_8924;
assign v_33469 = v_8762 | v_33468;
assign v_33470 = v_8730 | ~v_8792;
assign v_33472 = v_8473 | v_33471;
assign v_33473 = v_8447 | ~v_8628;
assign v_33475 = v_8474 | v_33474;
assign v_33476 = v_8448 | ~v_8496;
assign v_33478 = v_8185 | v_33477;
assign v_33479 = v_8157 | ~v_8344;
assign v_33481 = v_8186 | v_33480;
assign v_33482 = v_8158 | ~v_8212;
assign v_33484 = v_7901 | v_33483;
assign v_33485 = v_7876 | ~v_8056;
assign v_33487 = v_7902 | v_33486;
assign v_33488 = v_7877 | ~v_7924;
assign v_33490 = v_7607 | v_33489;
assign v_33491 = v_7571 | ~v_7774;
assign v_33493 = v_7608 | v_33492;
assign v_33494 = v_7572 | ~v_7642;
assign v_33496 = v_7315 | v_33495;
assign v_33497 = v_7288 | ~v_7470;
assign v_33499 = v_7316 | v_33498;
assign v_33500 = v_7289 | ~v_7338;
assign v_33502 = v_7025 | v_33501;
assign v_33503 = v_6997 | ~v_7184;
assign v_33505 = v_7026 | v_33504;
assign v_33506 = v_6998 | ~v_7052;
assign v_33508 = v_6741 | v_33507;
assign v_33509 = v_6716 | ~v_6896;
assign v_33511 = v_6742 | v_33510;
assign v_33512 = v_6717 | ~v_6764;
assign v_33514 = v_6451 | v_33513;
assign v_33515 = v_6419 | ~v_6614;
assign v_33517 = v_6452 | v_33516;
assign v_33518 = v_6420 | ~v_6482;
assign v_33520 = v_6163 | v_33519;
assign v_33521 = v_6137 | ~v_6318;
assign v_33523 = v_6164 | v_33522;
assign v_33524 = v_6138 | ~v_6186;
assign v_33526 = v_5875 | v_33525;
assign v_33527 = v_5847 | ~v_6034;
assign v_33529 = v_5876 | v_33528;
assign v_33530 = v_5848 | ~v_5902;
assign v_33532 = v_5591 | v_33531;
assign v_33533 = v_5566 | ~v_5746;
assign v_33535 = v_5592 | v_33534;
assign v_33536 = v_5567 | ~v_5614;
assign v_33538 = v_5293 | v_33537;
assign v_33539 = v_5253 | ~v_5464;
assign v_33541 = v_5294 | v_33540;
assign v_33542 = v_5254 | ~v_5332;
assign v_33544 = v_4997 | v_33543;
assign v_33545 = v_4969 | ~v_5152;
assign v_33547 = v_4998 | v_33546;
assign v_33548 = v_4970 | ~v_5020;
assign v_33550 = v_4705 | v_33549;
assign v_33551 = v_4677 | ~v_4864;
assign v_33553 = v_4706 | v_33552;
assign v_33554 = v_4678 | ~v_4732;
assign v_33556 = v_4421 | v_33555;
assign v_33557 = v_4396 | ~v_4576;
assign v_33559 = v_4422 | v_33558;
assign v_33560 = v_4397 | ~v_4444;
assign v_33562 = v_4131 | v_33561;
assign v_33563 = v_4099 | ~v_4294;
assign v_33565 = v_4132 | v_33564;
assign v_33566 = v_4100 | ~v_4162;
assign v_33568 = v_3843 | v_33567;
assign v_33569 = v_3817 | ~v_3998;
assign v_33571 = v_3844 | v_33570;
assign v_33572 = v_3818 | ~v_3866;
assign v_33574 = v_3555 | v_33573;
assign v_33575 = v_3527 | ~v_3714;
assign v_33577 = v_3556 | v_33576;
assign v_33578 = v_3528 | ~v_3582;
assign v_33580 = v_3271 | v_33579;
assign v_33581 = v_3246 | ~v_3426;
assign v_33583 = v_3272 | v_33582;
assign v_33584 = v_3247 | ~v_3294;
assign v_33586 = v_2977 | v_33585;
assign v_33587 = v_2941 | ~v_3144;
assign v_33589 = v_2978 | v_33588;
assign v_33590 = v_2942 | ~v_3012;
assign v_33592 = v_2685 | v_33591;
assign v_33593 = v_2658 | ~v_2840;
assign v_33595 = v_2686 | v_33594;
assign v_33596 = v_2659 | ~v_2708;
assign v_33598 = v_2395 | v_33597;
assign v_33599 = v_2367 | ~v_2554;
assign v_33601 = v_2396 | v_33600;
assign v_33602 = v_2368 | ~v_2422;
assign v_33604 = v_2111 | v_33603;
assign v_33605 = v_2086 | ~v_2266;
assign v_33607 = v_2112 | v_33606;
assign v_33608 = v_2087 | ~v_2134;
assign v_33610 = v_1821 | v_33609;
assign v_33611 = v_1789 | ~v_1984;
assign v_33613 = v_1822 | v_33612;
assign v_33614 = v_1790 | ~v_1852;
assign v_33616 = v_1533 | v_33615;
assign v_33617 = v_1507 | ~v_1688;
assign v_33619 = v_1534 | v_33618;
assign v_33620 = v_1508 | ~v_1556;
assign v_33622 = v_1245 | v_33621;
assign v_33623 = v_1217 | ~v_1404;
assign v_33625 = v_1246 | v_33624;
assign v_33626 = v_1218 | ~v_1272;
assign v_33628 = v_961 | v_33627;
assign v_33629 = v_936 | ~v_1116;
assign v_33631 = v_962 | v_33630;
assign v_33632 = v_937 | ~v_984;
assign v_33634 = v_591 | v_33633;
assign v_33635 = v_92 | ~v_838;
assign v_33637 = v_593 | v_33636;
assign v_33638 = v_94 | ~v_721;
assign v_33640 = v_9630 | ~v_9753;
assign v_33641 = v_9601 | ~v_9604;
assign v_33643 = v_9335 | v_33642;
assign v_33644 = v_9307 | ~v_9463;
assign v_33646 = v_9336 | v_33645;
assign v_33647 = v_9308 | ~v_9311;
assign v_33649 = v_9051 | v_33648;
assign v_33650 = v_9026 | ~v_9175;
assign v_33652 = v_9052 | v_33651;
assign v_33653 = v_9027 | ~v_9030;
assign v_33655 = v_8761 | v_33654;
assign v_33656 = v_8729 | ~v_8893;
assign v_33658 = v_8762 | v_33657;
assign v_33659 = v_8730 | ~v_8733;
assign v_33661 = v_8473 | v_33660;
assign v_33662 = v_8447 | ~v_8597;
assign v_33664 = v_8474 | v_33663;
assign v_33665 = v_8448 | ~v_8451;
assign v_33667 = v_8185 | v_33666;
assign v_33668 = v_8157 | ~v_8313;
assign v_33670 = v_8186 | v_33669;
assign v_33671 = v_8158 | ~v_8161;
assign v_33673 = v_7901 | v_33672;
assign v_33674 = v_7876 | ~v_8025;
assign v_33676 = v_7902 | v_33675;
assign v_33677 = v_7877 | ~v_7880;
assign v_33679 = v_7607 | v_33678;
assign v_33680 = v_7571 | ~v_7743;
assign v_33682 = v_7608 | v_33681;
assign v_33683 = v_7572 | ~v_7575;
assign v_33685 = v_7315 | v_33684;
assign v_33686 = v_7288 | ~v_7439;
assign v_33688 = v_7316 | v_33687;
assign v_33689 = v_7289 | ~v_7292;
assign v_33691 = v_7025 | v_33690;
assign v_33692 = v_6997 | ~v_7153;
assign v_33694 = v_7026 | v_33693;
assign v_33695 = v_6998 | ~v_7001;
assign v_33697 = v_6741 | v_33696;
assign v_33698 = v_6716 | ~v_6865;
assign v_33700 = v_6742 | v_33699;
assign v_33701 = v_6717 | ~v_6720;
assign v_33703 = v_6451 | v_33702;
assign v_33704 = v_6419 | ~v_6583;
assign v_33706 = v_6452 | v_33705;
assign v_33707 = v_6420 | ~v_6423;
assign v_33709 = v_6163 | v_33708;
assign v_33710 = v_6137 | ~v_6287;
assign v_33712 = v_6164 | v_33711;
assign v_33713 = v_6138 | ~v_6141;
assign v_33715 = v_5875 | v_33714;
assign v_33716 = v_5847 | ~v_6003;
assign v_33718 = v_5876 | v_33717;
assign v_33719 = v_5848 | ~v_5851;
assign v_33721 = v_5591 | v_33720;
assign v_33722 = v_5566 | ~v_5715;
assign v_33724 = v_5592 | v_33723;
assign v_33725 = v_5567 | ~v_5570;
assign v_33727 = v_5293 | v_33726;
assign v_33728 = v_5253 | ~v_5433;
assign v_33730 = v_5294 | v_33729;
assign v_33731 = v_5254 | ~v_5257;
assign v_33733 = v_4997 | v_33732;
assign v_33734 = v_4969 | ~v_5121;
assign v_33736 = v_4998 | v_33735;
assign v_33737 = v_4970 | ~v_4973;
assign v_33739 = v_4705 | v_33738;
assign v_33740 = v_4677 | ~v_4833;
assign v_33742 = v_4706 | v_33741;
assign v_33743 = v_4678 | ~v_4681;
assign v_33745 = v_4421 | v_33744;
assign v_33746 = v_4396 | ~v_4545;
assign v_33748 = v_4422 | v_33747;
assign v_33749 = v_4397 | ~v_4400;
assign v_33751 = v_4131 | v_33750;
assign v_33752 = v_4099 | ~v_4263;
assign v_33754 = v_4132 | v_33753;
assign v_33755 = v_4100 | ~v_4103;
assign v_33757 = v_3843 | v_33756;
assign v_33758 = v_3817 | ~v_3967;
assign v_33760 = v_3844 | v_33759;
assign v_33761 = v_3818 | ~v_3821;
assign v_33763 = v_3555 | v_33762;
assign v_33764 = v_3527 | ~v_3683;
assign v_33766 = v_3556 | v_33765;
assign v_33767 = v_3528 | ~v_3531;
assign v_33769 = v_3271 | v_33768;
assign v_33770 = v_3246 | ~v_3395;
assign v_33772 = v_3272 | v_33771;
assign v_33773 = v_3247 | ~v_3250;
assign v_33775 = v_2977 | v_33774;
assign v_33776 = v_2941 | ~v_3113;
assign v_33778 = v_2978 | v_33777;
assign v_33779 = v_2942 | ~v_2945;
assign v_33781 = v_2685 | v_33780;
assign v_33782 = v_2658 | ~v_2809;
assign v_33784 = v_2686 | v_33783;
assign v_33785 = v_2659 | ~v_2662;
assign v_33787 = v_2395 | v_33786;
assign v_33788 = v_2367 | ~v_2523;
assign v_33790 = v_2396 | v_33789;
assign v_33791 = v_2368 | ~v_2371;
assign v_33793 = v_2111 | v_33792;
assign v_33794 = v_2086 | ~v_2235;
assign v_33796 = v_2112 | v_33795;
assign v_33797 = v_2087 | ~v_2090;
assign v_33799 = v_1821 | v_33798;
assign v_33800 = v_1789 | ~v_1953;
assign v_33802 = v_1822 | v_33801;
assign v_33803 = v_1790 | ~v_1793;
assign v_33805 = v_1533 | v_33804;
assign v_33806 = v_1507 | ~v_1657;
assign v_33808 = v_1534 | v_33807;
assign v_33809 = v_1508 | ~v_1511;
assign v_33811 = v_1245 | v_33810;
assign v_33812 = v_1217 | ~v_1373;
assign v_33814 = v_1246 | v_33813;
assign v_33815 = v_1218 | ~v_1221;
assign v_33817 = v_961 | v_33816;
assign v_33818 = v_936 | ~v_1085;
assign v_33820 = v_962 | v_33819;
assign v_33821 = v_937 | ~v_940;
assign v_33823 = v_591 | v_33822;
assign v_33824 = v_92 | ~v_804;
assign v_33826 = v_593 | v_33825;
assign v_33827 = v_94 | ~v_98;
assign v_33830 = v_9630 | ~v_9796;
assign v_33831 = v_9601 | ~v_9664;
assign v_33833 = v_9335 | v_33832;
assign v_33834 = v_9307 | ~v_9506;
assign v_33836 = v_9336 | v_33835;
assign v_33837 = v_9308 | ~v_9374;
assign v_33839 = v_9051 | v_33838;
assign v_33840 = v_9026 | ~v_9218;
assign v_33842 = v_9052 | v_33841;
assign v_33843 = v_9027 | ~v_9086;
assign v_33845 = v_8761 | v_33844;
assign v_33846 = v_8729 | ~v_8936;
assign v_33848 = v_8762 | v_33847;
assign v_33849 = v_8730 | ~v_8804;
assign v_33851 = v_8473 | v_33850;
assign v_33852 = v_8447 | ~v_8640;
assign v_33854 = v_8474 | v_33853;
assign v_33855 = v_8448 | ~v_8508;
assign v_33857 = v_8185 | v_33856;
assign v_33858 = v_8157 | ~v_8356;
assign v_33860 = v_8186 | v_33859;
assign v_33861 = v_8158 | ~v_8224;
assign v_33863 = v_7901 | v_33862;
assign v_33864 = v_7876 | ~v_8068;
assign v_33866 = v_7902 | v_33865;
assign v_33867 = v_7877 | ~v_7936;
assign v_33869 = v_7607 | v_33868;
assign v_33870 = v_7571 | ~v_7786;
assign v_33872 = v_7608 | v_33871;
assign v_33873 = v_7572 | ~v_7654;
assign v_33875 = v_7315 | v_33874;
assign v_33876 = v_7288 | ~v_7482;
assign v_33878 = v_7316 | v_33877;
assign v_33879 = v_7289 | ~v_7350;
assign v_33881 = v_7025 | v_33880;
assign v_33882 = v_6997 | ~v_7196;
assign v_33884 = v_7026 | v_33883;
assign v_33885 = v_6998 | ~v_7064;
assign v_33887 = v_6741 | v_33886;
assign v_33888 = v_6716 | ~v_6908;
assign v_33890 = v_6742 | v_33889;
assign v_33891 = v_6717 | ~v_6776;
assign v_33893 = v_6451 | v_33892;
assign v_33894 = v_6419 | ~v_6626;
assign v_33896 = v_6452 | v_33895;
assign v_33897 = v_6420 | ~v_6494;
assign v_33899 = v_6163 | v_33898;
assign v_33900 = v_6137 | ~v_6330;
assign v_33902 = v_6164 | v_33901;
assign v_33903 = v_6138 | ~v_6198;
assign v_33905 = v_5875 | v_33904;
assign v_33906 = v_5847 | ~v_6046;
assign v_33908 = v_5876 | v_33907;
assign v_33909 = v_5848 | ~v_5914;
assign v_33911 = v_5591 | v_33910;
assign v_33912 = v_5566 | ~v_5758;
assign v_33914 = v_5592 | v_33913;
assign v_33915 = v_5567 | ~v_5626;
assign v_33917 = v_5293 | v_33916;
assign v_33918 = v_5253 | ~v_5476;
assign v_33920 = v_5294 | v_33919;
assign v_33921 = v_5254 | ~v_5344;
assign v_33923 = v_4997 | v_33922;
assign v_33924 = v_4969 | ~v_5164;
assign v_33926 = v_4998 | v_33925;
assign v_33927 = v_4970 | ~v_5032;
assign v_33929 = v_4705 | v_33928;
assign v_33930 = v_4677 | ~v_4876;
assign v_33932 = v_4706 | v_33931;
assign v_33933 = v_4678 | ~v_4744;
assign v_33935 = v_4421 | v_33934;
assign v_33936 = v_4396 | ~v_4588;
assign v_33938 = v_4422 | v_33937;
assign v_33939 = v_4397 | ~v_4456;
assign v_33941 = v_4131 | v_33940;
assign v_33942 = v_4099 | ~v_4306;
assign v_33944 = v_4132 | v_33943;
assign v_33945 = v_4100 | ~v_4174;
assign v_33947 = v_3843 | v_33946;
assign v_33948 = v_3817 | ~v_4010;
assign v_33950 = v_3844 | v_33949;
assign v_33951 = v_3818 | ~v_3878;
assign v_33953 = v_3555 | v_33952;
assign v_33954 = v_3527 | ~v_3726;
assign v_33956 = v_3556 | v_33955;
assign v_33957 = v_3528 | ~v_3594;
assign v_33959 = v_3271 | v_33958;
assign v_33960 = v_3246 | ~v_3438;
assign v_33962 = v_3272 | v_33961;
assign v_33963 = v_3247 | ~v_3306;
assign v_33965 = v_2977 | v_33964;
assign v_33966 = v_2941 | ~v_3156;
assign v_33968 = v_2978 | v_33967;
assign v_33969 = v_2942 | ~v_3024;
assign v_33971 = v_2685 | v_33970;
assign v_33972 = v_2658 | ~v_2852;
assign v_33974 = v_2686 | v_33973;
assign v_33975 = v_2659 | ~v_2720;
assign v_33977 = v_2395 | v_33976;
assign v_33978 = v_2367 | ~v_2566;
assign v_33980 = v_2396 | v_33979;
assign v_33981 = v_2368 | ~v_2434;
assign v_33983 = v_2111 | v_33982;
assign v_33984 = v_2086 | ~v_2278;
assign v_33986 = v_2112 | v_33985;
assign v_33987 = v_2087 | ~v_2146;
assign v_33989 = v_1821 | v_33988;
assign v_33990 = v_1789 | ~v_1996;
assign v_33992 = v_1822 | v_33991;
assign v_33993 = v_1790 | ~v_1864;
assign v_33995 = v_1533 | v_33994;
assign v_33996 = v_1507 | ~v_1700;
assign v_33998 = v_1534 | v_33997;
assign v_33999 = v_1508 | ~v_1568;
assign v_34001 = v_1245 | v_34000;
assign v_34002 = v_1217 | ~v_1416;
assign v_34004 = v_1246 | v_34003;
assign v_34005 = v_1218 | ~v_1284;
assign v_34007 = v_961 | v_34006;
assign v_34008 = v_936 | ~v_1128;
assign v_34010 = v_962 | v_34009;
assign v_34011 = v_937 | ~v_996;
assign v_34013 = v_591 | v_34012;
assign v_34014 = v_92 | ~v_850;
assign v_34016 = v_593 | v_34015;
assign v_34017 = v_94 | ~v_731;
assign v_34020 = v_9630 | ~v_9808;
assign v_34021 = v_9601 | ~v_9676;
assign v_34023 = v_9335 | v_34022;
assign v_34024 = v_9307 | ~v_9518;
assign v_34026 = v_9336 | v_34025;
assign v_34027 = v_9308 | ~v_9386;
assign v_34029 = v_9051 | v_34028;
assign v_34030 = v_9026 | ~v_9230;
assign v_34032 = v_9052 | v_34031;
assign v_34033 = v_9027 | ~v_9098;
assign v_34035 = v_8761 | v_34034;
assign v_34036 = v_8729 | ~v_8948;
assign v_34038 = v_8762 | v_34037;
assign v_34039 = v_8730 | ~v_8816;
assign v_34041 = v_8473 | v_34040;
assign v_34042 = v_8447 | ~v_8652;
assign v_34044 = v_8474 | v_34043;
assign v_34045 = v_8448 | ~v_8520;
assign v_34047 = v_8185 | v_34046;
assign v_34048 = v_8157 | ~v_8368;
assign v_34050 = v_8186 | v_34049;
assign v_34051 = v_8158 | ~v_8236;
assign v_34053 = v_7901 | v_34052;
assign v_34054 = v_7876 | ~v_8080;
assign v_34056 = v_7902 | v_34055;
assign v_34057 = v_7877 | ~v_7948;
assign v_34059 = v_7607 | v_34058;
assign v_34060 = v_7571 | ~v_7798;
assign v_34062 = v_7608 | v_34061;
assign v_34063 = v_7572 | ~v_7666;
assign v_34065 = v_7315 | v_34064;
assign v_34066 = v_7288 | ~v_7494;
assign v_34068 = v_7316 | v_34067;
assign v_34069 = v_7289 | ~v_7362;
assign v_34071 = v_7025 | v_34070;
assign v_34072 = v_6997 | ~v_7208;
assign v_34074 = v_7026 | v_34073;
assign v_34075 = v_6998 | ~v_7076;
assign v_34077 = v_6741 | v_34076;
assign v_34078 = v_6716 | ~v_6920;
assign v_34080 = v_6742 | v_34079;
assign v_34081 = v_6717 | ~v_6788;
assign v_34083 = v_6451 | v_34082;
assign v_34084 = v_6419 | ~v_6638;
assign v_34086 = v_6452 | v_34085;
assign v_34087 = v_6420 | ~v_6506;
assign v_34089 = v_6163 | v_34088;
assign v_34090 = v_6137 | ~v_6342;
assign v_34092 = v_6164 | v_34091;
assign v_34093 = v_6138 | ~v_6210;
assign v_34095 = v_5875 | v_34094;
assign v_34096 = v_5847 | ~v_6058;
assign v_34098 = v_5876 | v_34097;
assign v_34099 = v_5848 | ~v_5926;
assign v_34101 = v_5591 | v_34100;
assign v_34102 = v_5566 | ~v_5770;
assign v_34104 = v_5592 | v_34103;
assign v_34105 = v_5567 | ~v_5638;
assign v_34107 = v_5293 | v_34106;
assign v_34108 = v_5253 | ~v_5488;
assign v_34110 = v_5294 | v_34109;
assign v_34111 = v_5254 | ~v_5356;
assign v_34113 = v_4997 | v_34112;
assign v_34114 = v_4969 | ~v_5176;
assign v_34116 = v_4998 | v_34115;
assign v_34117 = v_4970 | ~v_5044;
assign v_34119 = v_4705 | v_34118;
assign v_34120 = v_4677 | ~v_4888;
assign v_34122 = v_4706 | v_34121;
assign v_34123 = v_4678 | ~v_4756;
assign v_34125 = v_4421 | v_34124;
assign v_34126 = v_4396 | ~v_4600;
assign v_34128 = v_4422 | v_34127;
assign v_34129 = v_4397 | ~v_4468;
assign v_34131 = v_4131 | v_34130;
assign v_34132 = v_4099 | ~v_4318;
assign v_34134 = v_4132 | v_34133;
assign v_34135 = v_4100 | ~v_4186;
assign v_34137 = v_3843 | v_34136;
assign v_34138 = v_3817 | ~v_4022;
assign v_34140 = v_3844 | v_34139;
assign v_34141 = v_3818 | ~v_3890;
assign v_34143 = v_3555 | v_34142;
assign v_34144 = v_3527 | ~v_3738;
assign v_34146 = v_3556 | v_34145;
assign v_34147 = v_3528 | ~v_3606;
assign v_34149 = v_3271 | v_34148;
assign v_34150 = v_3246 | ~v_3450;
assign v_34152 = v_3272 | v_34151;
assign v_34153 = v_3247 | ~v_3318;
assign v_34155 = v_2977 | v_34154;
assign v_34156 = v_2941 | ~v_3168;
assign v_34158 = v_2978 | v_34157;
assign v_34159 = v_2942 | ~v_3036;
assign v_34161 = v_2685 | v_34160;
assign v_34162 = v_2658 | ~v_2864;
assign v_34164 = v_2686 | v_34163;
assign v_34165 = v_2659 | ~v_2732;
assign v_34167 = v_2395 | v_34166;
assign v_34168 = v_2367 | ~v_2578;
assign v_34170 = v_2396 | v_34169;
assign v_34171 = v_2368 | ~v_2446;
assign v_34173 = v_2111 | v_34172;
assign v_34174 = v_2086 | ~v_2290;
assign v_34176 = v_2112 | v_34175;
assign v_34177 = v_2087 | ~v_2158;
assign v_34179 = v_1821 | v_34178;
assign v_34180 = v_1789 | ~v_2008;
assign v_34182 = v_1822 | v_34181;
assign v_34183 = v_1790 | ~v_1876;
assign v_34185 = v_1533 | v_34184;
assign v_34186 = v_1507 | ~v_1712;
assign v_34188 = v_1534 | v_34187;
assign v_34189 = v_1508 | ~v_1580;
assign v_34191 = v_1245 | v_34190;
assign v_34192 = v_1217 | ~v_1428;
assign v_34194 = v_1246 | v_34193;
assign v_34195 = v_1218 | ~v_1296;
assign v_34197 = v_961 | v_34196;
assign v_34198 = v_936 | ~v_1140;
assign v_34200 = v_962 | v_34199;
assign v_34201 = v_937 | ~v_1008;
assign v_34203 = v_591 | v_34202;
assign v_34204 = v_92 | ~v_862;
assign v_34206 = v_593 | v_34205;
assign v_34207 = v_94 | ~v_741;
assign v_34210 = v_9630 | ~v_9820;
assign v_34211 = v_9601 | ~v_9688;
assign v_34213 = v_9335 | v_34212;
assign v_34214 = v_9307 | ~v_9530;
assign v_34216 = v_9336 | v_34215;
assign v_34217 = v_9308 | ~v_9398;
assign v_34219 = v_9051 | v_34218;
assign v_34220 = v_9026 | ~v_9242;
assign v_34222 = v_9052 | v_34221;
assign v_34223 = v_9027 | ~v_9110;
assign v_34225 = v_8761 | v_34224;
assign v_34226 = v_8729 | ~v_8960;
assign v_34228 = v_8762 | v_34227;
assign v_34229 = v_8730 | ~v_8828;
assign v_34231 = v_8473 | v_34230;
assign v_34232 = v_8447 | ~v_8664;
assign v_34234 = v_8474 | v_34233;
assign v_34235 = v_8448 | ~v_8532;
assign v_34237 = v_8185 | v_34236;
assign v_34238 = v_8157 | ~v_8380;
assign v_34240 = v_8186 | v_34239;
assign v_34241 = v_8158 | ~v_8248;
assign v_34243 = v_7901 | v_34242;
assign v_34244 = v_7876 | ~v_8092;
assign v_34246 = v_7902 | v_34245;
assign v_34247 = v_7877 | ~v_7960;
assign v_34249 = v_7607 | v_34248;
assign v_34250 = v_7571 | ~v_7810;
assign v_34252 = v_7608 | v_34251;
assign v_34253 = v_7572 | ~v_7678;
assign v_34255 = v_7315 | v_34254;
assign v_34256 = v_7288 | ~v_7506;
assign v_34258 = v_7316 | v_34257;
assign v_34259 = v_7289 | ~v_7374;
assign v_34261 = v_7025 | v_34260;
assign v_34262 = v_6997 | ~v_7220;
assign v_34264 = v_7026 | v_34263;
assign v_34265 = v_6998 | ~v_7088;
assign v_34267 = v_6741 | v_34266;
assign v_34268 = v_6716 | ~v_6932;
assign v_34270 = v_6742 | v_34269;
assign v_34271 = v_6717 | ~v_6800;
assign v_34273 = v_6451 | v_34272;
assign v_34274 = v_6419 | ~v_6650;
assign v_34276 = v_6452 | v_34275;
assign v_34277 = v_6420 | ~v_6518;
assign v_34279 = v_6163 | v_34278;
assign v_34280 = v_6137 | ~v_6354;
assign v_34282 = v_6164 | v_34281;
assign v_34283 = v_6138 | ~v_6222;
assign v_34285 = v_5875 | v_34284;
assign v_34286 = v_5847 | ~v_6070;
assign v_34288 = v_5876 | v_34287;
assign v_34289 = v_5848 | ~v_5938;
assign v_34291 = v_5591 | v_34290;
assign v_34292 = v_5566 | ~v_5782;
assign v_34294 = v_5592 | v_34293;
assign v_34295 = v_5567 | ~v_5650;
assign v_34297 = v_5293 | v_34296;
assign v_34298 = v_5253 | ~v_5500;
assign v_34300 = v_5294 | v_34299;
assign v_34301 = v_5254 | ~v_5368;
assign v_34303 = v_4997 | v_34302;
assign v_34304 = v_4969 | ~v_5188;
assign v_34306 = v_4998 | v_34305;
assign v_34307 = v_4970 | ~v_5056;
assign v_34309 = v_4705 | v_34308;
assign v_34310 = v_4677 | ~v_4900;
assign v_34312 = v_4706 | v_34311;
assign v_34313 = v_4678 | ~v_4768;
assign v_34315 = v_4421 | v_34314;
assign v_34316 = v_4396 | ~v_4612;
assign v_34318 = v_4422 | v_34317;
assign v_34319 = v_4397 | ~v_4480;
assign v_34321 = v_4131 | v_34320;
assign v_34322 = v_4099 | ~v_4330;
assign v_34324 = v_4132 | v_34323;
assign v_34325 = v_4100 | ~v_4198;
assign v_34327 = v_3843 | v_34326;
assign v_34328 = v_3817 | ~v_4034;
assign v_34330 = v_3844 | v_34329;
assign v_34331 = v_3818 | ~v_3902;
assign v_34333 = v_3555 | v_34332;
assign v_34334 = v_3527 | ~v_3750;
assign v_34336 = v_3556 | v_34335;
assign v_34337 = v_3528 | ~v_3618;
assign v_34339 = v_3271 | v_34338;
assign v_34340 = v_3246 | ~v_3462;
assign v_34342 = v_3272 | v_34341;
assign v_34343 = v_3247 | ~v_3330;
assign v_34345 = v_2977 | v_34344;
assign v_34346 = v_2941 | ~v_3180;
assign v_34348 = v_2978 | v_34347;
assign v_34349 = v_2942 | ~v_3048;
assign v_34351 = v_2685 | v_34350;
assign v_34352 = v_2658 | ~v_2876;
assign v_34354 = v_2686 | v_34353;
assign v_34355 = v_2659 | ~v_2744;
assign v_34357 = v_2395 | v_34356;
assign v_34358 = v_2367 | ~v_2590;
assign v_34360 = v_2396 | v_34359;
assign v_34361 = v_2368 | ~v_2458;
assign v_34363 = v_2111 | v_34362;
assign v_34364 = v_2086 | ~v_2302;
assign v_34366 = v_2112 | v_34365;
assign v_34367 = v_2087 | ~v_2170;
assign v_34369 = v_1821 | v_34368;
assign v_34370 = v_1789 | ~v_2020;
assign v_34372 = v_1822 | v_34371;
assign v_34373 = v_1790 | ~v_1888;
assign v_34375 = v_1533 | v_34374;
assign v_34376 = v_1507 | ~v_1724;
assign v_34378 = v_1534 | v_34377;
assign v_34379 = v_1508 | ~v_1592;
assign v_34381 = v_1245 | v_34380;
assign v_34382 = v_1217 | ~v_1440;
assign v_34384 = v_1246 | v_34383;
assign v_34385 = v_1218 | ~v_1308;
assign v_34387 = v_961 | v_34386;
assign v_34388 = v_936 | ~v_1152;
assign v_34390 = v_962 | v_34389;
assign v_34391 = v_937 | ~v_1020;
assign v_34393 = v_591 | v_34392;
assign v_34394 = v_92 | ~v_874;
assign v_34396 = v_593 | v_34395;
assign v_34397 = v_94 | ~v_751;
assign v_34400 = v_9630 | ~v_9832;
assign v_34401 = v_9601 | ~v_9700;
assign v_34403 = v_9335 | v_34402;
assign v_34404 = v_9307 | ~v_9542;
assign v_34406 = v_9336 | v_34405;
assign v_34407 = v_9308 | ~v_9410;
assign v_34409 = v_9051 | v_34408;
assign v_34410 = v_9026 | ~v_9254;
assign v_34412 = v_9052 | v_34411;
assign v_34413 = v_9027 | ~v_9122;
assign v_34415 = v_8761 | v_34414;
assign v_34416 = v_8729 | ~v_8972;
assign v_34418 = v_8762 | v_34417;
assign v_34419 = v_8730 | ~v_8840;
assign v_34421 = v_8473 | v_34420;
assign v_34422 = v_8447 | ~v_8676;
assign v_34424 = v_8474 | v_34423;
assign v_34425 = v_8448 | ~v_8544;
assign v_34427 = v_8185 | v_34426;
assign v_34428 = v_8157 | ~v_8392;
assign v_34430 = v_8186 | v_34429;
assign v_34431 = v_8158 | ~v_8260;
assign v_34433 = v_7901 | v_34432;
assign v_34434 = v_7876 | ~v_8104;
assign v_34436 = v_7902 | v_34435;
assign v_34437 = v_7877 | ~v_7972;
assign v_34439 = v_7607 | v_34438;
assign v_34440 = v_7571 | ~v_7822;
assign v_34442 = v_7608 | v_34441;
assign v_34443 = v_7572 | ~v_7690;
assign v_34445 = v_7315 | v_34444;
assign v_34446 = v_7288 | ~v_7518;
assign v_34448 = v_7316 | v_34447;
assign v_34449 = v_7289 | ~v_7386;
assign v_34451 = v_7025 | v_34450;
assign v_34452 = v_6997 | ~v_7232;
assign v_34454 = v_7026 | v_34453;
assign v_34455 = v_6998 | ~v_7100;
assign v_34457 = v_6741 | v_34456;
assign v_34458 = v_6716 | ~v_6944;
assign v_34460 = v_6742 | v_34459;
assign v_34461 = v_6717 | ~v_6812;
assign v_34463 = v_6451 | v_34462;
assign v_34464 = v_6419 | ~v_6662;
assign v_34466 = v_6452 | v_34465;
assign v_34467 = v_6420 | ~v_6530;
assign v_34469 = v_6163 | v_34468;
assign v_34470 = v_6137 | ~v_6366;
assign v_34472 = v_6164 | v_34471;
assign v_34473 = v_6138 | ~v_6234;
assign v_34475 = v_5875 | v_34474;
assign v_34476 = v_5847 | ~v_6082;
assign v_34478 = v_5876 | v_34477;
assign v_34479 = v_5848 | ~v_5950;
assign v_34481 = v_5591 | v_34480;
assign v_34482 = v_5566 | ~v_5794;
assign v_34484 = v_5592 | v_34483;
assign v_34485 = v_5567 | ~v_5662;
assign v_34487 = v_5293 | v_34486;
assign v_34488 = v_5253 | ~v_5512;
assign v_34490 = v_5294 | v_34489;
assign v_34491 = v_5254 | ~v_5380;
assign v_34493 = v_4997 | v_34492;
assign v_34494 = v_4969 | ~v_5200;
assign v_34496 = v_4998 | v_34495;
assign v_34497 = v_4970 | ~v_5068;
assign v_34499 = v_4705 | v_34498;
assign v_34500 = v_4677 | ~v_4912;
assign v_34502 = v_4706 | v_34501;
assign v_34503 = v_4678 | ~v_4780;
assign v_34505 = v_4421 | v_34504;
assign v_34506 = v_4396 | ~v_4624;
assign v_34508 = v_4422 | v_34507;
assign v_34509 = v_4397 | ~v_4492;
assign v_34511 = v_4131 | v_34510;
assign v_34512 = v_4099 | ~v_4342;
assign v_34514 = v_4132 | v_34513;
assign v_34515 = v_4100 | ~v_4210;
assign v_34517 = v_3843 | v_34516;
assign v_34518 = v_3817 | ~v_4046;
assign v_34520 = v_3844 | v_34519;
assign v_34521 = v_3818 | ~v_3914;
assign v_34523 = v_3555 | v_34522;
assign v_34524 = v_3527 | ~v_3762;
assign v_34526 = v_3556 | v_34525;
assign v_34527 = v_3528 | ~v_3630;
assign v_34529 = v_3271 | v_34528;
assign v_34530 = v_3246 | ~v_3474;
assign v_34532 = v_3272 | v_34531;
assign v_34533 = v_3247 | ~v_3342;
assign v_34535 = v_2977 | v_34534;
assign v_34536 = v_2941 | ~v_3192;
assign v_34538 = v_2978 | v_34537;
assign v_34539 = v_2942 | ~v_3060;
assign v_34541 = v_2685 | v_34540;
assign v_34542 = v_2658 | ~v_2888;
assign v_34544 = v_2686 | v_34543;
assign v_34545 = v_2659 | ~v_2756;
assign v_34547 = v_2395 | v_34546;
assign v_34548 = v_2367 | ~v_2602;
assign v_34550 = v_2396 | v_34549;
assign v_34551 = v_2368 | ~v_2470;
assign v_34553 = v_2111 | v_34552;
assign v_34554 = v_2086 | ~v_2314;
assign v_34556 = v_2112 | v_34555;
assign v_34557 = v_2087 | ~v_2182;
assign v_34559 = v_1821 | v_34558;
assign v_34560 = v_1789 | ~v_2032;
assign v_34562 = v_1822 | v_34561;
assign v_34563 = v_1790 | ~v_1900;
assign v_34565 = v_1533 | v_34564;
assign v_34566 = v_1507 | ~v_1736;
assign v_34568 = v_1534 | v_34567;
assign v_34569 = v_1508 | ~v_1604;
assign v_34571 = v_1245 | v_34570;
assign v_34572 = v_1217 | ~v_1452;
assign v_34574 = v_1246 | v_34573;
assign v_34575 = v_1218 | ~v_1320;
assign v_34577 = v_961 | v_34576;
assign v_34578 = v_936 | ~v_1164;
assign v_34580 = v_962 | v_34579;
assign v_34581 = v_937 | ~v_1032;
assign v_34583 = v_591 | v_34582;
assign v_34584 = v_92 | ~v_886;
assign v_34586 = v_593 | v_34585;
assign v_34587 = v_94 | ~v_761;
assign v_34591 = v_9630 | v_9872;
assign v_34592 = v_9601 | v_9740;
assign v_34594 = v_9335 | v_34593;
assign v_34595 = v_9307 | v_9582;
assign v_34597 = v_9336 | v_34596;
assign v_34598 = v_9308 | v_9450;
assign v_34600 = v_9051 | v_34599;
assign v_34601 = v_9026 | v_9294;
assign v_34603 = v_9052 | v_34602;
assign v_34604 = v_9027 | v_9162;
assign v_34606 = v_8761 | v_34605;
assign v_34607 = v_8729 | v_9012;
assign v_34609 = v_8762 | v_34608;
assign v_34610 = v_8730 | v_8880;
assign v_34612 = v_8473 | v_34611;
assign v_34613 = v_8447 | v_8716;
assign v_34615 = v_8474 | v_34614;
assign v_34616 = v_8448 | v_8584;
assign v_34618 = v_8185 | v_34617;
assign v_34619 = v_8157 | ~v_8432;
assign v_34621 = v_8186 | v_34620;
assign v_34622 = v_8158 | ~v_8300;
assign v_34624 = v_7901 | v_34623;
assign v_34625 = v_7876 | ~v_8144;
assign v_34627 = v_7902 | v_34626;
assign v_34628 = v_7877 | v_8012;
assign v_34630 = v_7607 | v_34629;
assign v_34631 = v_7571 | v_7862;
assign v_34633 = v_7608 | v_34632;
assign v_34634 = v_7572 | v_7730;
assign v_34636 = v_7315 | v_34635;
assign v_34637 = v_7288 | v_7558;
assign v_34639 = v_7316 | v_34638;
assign v_34640 = v_7289 | v_7426;
assign v_34642 = v_7025 | v_34641;
assign v_34643 = v_6997 | ~v_7272;
assign v_34645 = v_7026 | v_34644;
assign v_34646 = v_6998 | v_7140;
assign v_34648 = v_6741 | v_34647;
assign v_34649 = v_6716 | ~v_6984;
assign v_34651 = v_6742 | v_34650;
assign v_34652 = v_6717 | ~v_6852;
assign v_34654 = v_6451 | v_34653;
assign v_34655 = v_6419 | ~v_6702;
assign v_34657 = v_6452 | v_34656;
assign v_34658 = v_6420 | v_6570;
assign v_34660 = v_6163 | v_34659;
assign v_34661 = v_6137 | v_6406;
assign v_34663 = v_6164 | v_34662;
assign v_34664 = v_6138 | ~v_6274;
assign v_34666 = v_5875 | v_34665;
assign v_34667 = v_5847 | ~v_6122;
assign v_34669 = v_5876 | v_34668;
assign v_34670 = v_5848 | ~v_5990;
assign v_34672 = v_5591 | v_34671;
assign v_34673 = v_5566 | ~v_5834;
assign v_34675 = v_5592 | v_34674;
assign v_34676 = v_5567 | ~v_5702;
assign v_34678 = v_5293 | v_34677;
assign v_34679 = v_5253 | ~v_5552;
assign v_34681 = v_5294 | v_34680;
assign v_34682 = v_5254 | v_5420;
assign v_34684 = v_4997 | v_34683;
assign v_34685 = v_4969 | v_5240;
assign v_34687 = v_4998 | v_34686;
assign v_34688 = v_4970 | ~v_5108;
assign v_34690 = v_4705 | v_34689;
assign v_34691 = v_4677 | ~v_4952;
assign v_34693 = v_4706 | v_34692;
assign v_34694 = v_4678 | ~v_4820;
assign v_34696 = v_4421 | v_34695;
assign v_34697 = v_4396 | ~v_4664;
assign v_34699 = v_4422 | v_34698;
assign v_34700 = v_4397 | ~v_4532;
assign v_34702 = v_4131 | v_34701;
assign v_34703 = v_4099 | ~v_4382;
assign v_34705 = v_4132 | v_34704;
assign v_34706 = v_4100 | v_4250;
assign v_34708 = v_3843 | v_34707;
assign v_34709 = v_3817 | v_4086;
assign v_34711 = v_3844 | v_34710;
assign v_34712 = v_3818 | v_3954;
assign v_34714 = v_3555 | v_34713;
assign v_34715 = v_3527 | v_3802;
assign v_34717 = v_3556 | v_34716;
assign v_34718 = v_3528 | v_3670;
assign v_34720 = v_3271 | v_34719;
assign v_34721 = v_3246 | ~v_3514;
assign v_34723 = v_3272 | v_34722;
assign v_34724 = v_3247 | v_3382;
assign v_34726 = v_2977 | v_34725;
assign v_34727 = v_2941 | ~v_3232;
assign v_34729 = v_2978 | v_34728;
assign v_34730 = v_2942 | v_3100;
assign v_34732 = v_2685 | v_34731;
assign v_34733 = v_2658 | v_2928;
assign v_34735 = v_2686 | v_34734;
assign v_34736 = v_2659 | v_2796;
assign v_34738 = v_2395 | v_34737;
assign v_34739 = v_2367 | v_2642;
assign v_34741 = v_2396 | v_34740;
assign v_34742 = v_2368 | v_2510;
assign v_34744 = v_2111 | v_34743;
assign v_34745 = v_2086 | ~v_2354;
assign v_34747 = v_2112 | v_34746;
assign v_34748 = v_2087 | ~v_2222;
assign v_34750 = v_1821 | v_34749;
assign v_34751 = v_1789 | ~v_2072;
assign v_34753 = v_1822 | v_34752;
assign v_34754 = v_1790 | v_1940;
assign v_34756 = v_1533 | v_34755;
assign v_34757 = v_1507 | v_1776;
assign v_34759 = v_1534 | v_34758;
assign v_34760 = v_1508 | v_1644;
assign v_34762 = v_1245 | v_34761;
assign v_34763 = v_1217 | v_1492;
assign v_34765 = v_1246 | v_34764;
assign v_34766 = v_1218 | v_1360;
assign v_34768 = v_961 | v_34767;
assign v_34769 = v_936 | v_1204;
assign v_34771 = v_962 | v_34770;
assign v_34772 = v_937 | v_1072;
assign v_34774 = v_591 | v_34773;
assign v_34775 = v_92 | v_922;
assign v_34777 = v_593 | v_34776;
assign v_34778 = v_94 | v_793;
assign v_34784 = ~v_96 | v_34783;
assign v_34789 = ~v_10200 | v_34788;
assign v_34794 = ~v_10196 | v_34793;
assign v_34799 = ~v_9903 | v_34798;
assign v_34804 = ~v_9884 | v_34803;
assign v_34838 = ~v_10415 | v_34837;
assign v_34851 = v_10465 | v_34850;
assign v_34855 = ~v_34852 | v_34854;
assign v_34856 = ~v_4 | v_13539;
assign v_34857 = v_3 | v_34856;
assign v_34858 = v_34852 | v_34857;
assign v_34860 = ~v_10456 | v_10465;
assign x_1 = v_6 | v_34862;
assign o_1 = x_1;
endmodule
