module formula(v_1,v_2,v_3,v_4,v_5,v_6,v_7,v_8,v_9,v_10,v_11,v_12,v_13,v_14,v_15,v_16,v_17,v_18,v_19,v_20,v_21,v_22,v_23,v_24,v_25,v_26,v_27,v_28,v_29,v_30,v_31,v_32,v_33,v_34,v_35,v_36,v_37,v_38,v_39,v_40,v_41,v_42,v_43,v_44,v_45,v_46,v_47,v_48,v_49,v_50,v_51,v_52,v_53,v_54,v_55,v_56,v_57,v_58,v_59,v_60,v_61,v_62,v_63,v_64,v_65,v_66,v_67,v_68,v_69,v_70,v_71,v_72,v_73,v_74,v_75,v_76,v_77,v_78,v_79,v_80,v_81,v_82,v_83,v_84,v_85,v_86,v_87,v_88,v_89,v_90,v_91,v_92,v_93,v_94,v_95,v_96,v_97,v_98,v_99,v_100,v_101,v_102,v_103,v_104,v_105,v_106,v_107,v_108,v_109,v_110,v_111,v_112,v_113,v_114,v_115,v_116,v_117,v_118,v_119,v_120,v_121,v_122,v_123,v_124,v_125,v_126,v_127,v_128,v_129,v_130,v_131,v_132,v_133,v_134,v_135,v_136,v_137,v_138,v_139,v_140,v_141,v_142,v_143,v_144,v_145,v_146,v_147,v_148,v_149,v_150,v_151,v_152,v_153,v_154,v_155,v_156,v_157,v_158,v_159,v_160,v_161,v_162,v_163,v_164,v_165,v_166,v_167,v_168,o_1);
	input v_1;
	input v_2;
	input v_3;
	input v_4;
	input v_5;
	input v_6;
	input v_7;
	input v_8;
	input v_9;
	input v_10;
	input v_11;
	input v_12;
	input v_13;
	input v_14;
	input v_15;
	input v_16;
	input v_17;
	input v_18;
	input v_19;
	input v_20;
	input v_21;
	input v_22;
	input v_23;
	input v_24;
	input v_25;
	input v_26;
	input v_27;
	input v_28;
	input v_29;
	input v_30;
	input v_31;
	input v_32;
	input v_33;
	input v_34;
	input v_35;
	input v_36;
	input v_37;
	input v_38;
	input v_39;
	input v_40;
	input v_41;
	input v_42;
	input v_43;
	input v_44;
	input v_45;
	input v_46;
	input v_47;
	input v_48;
	input v_49;
	input v_50;
	input v_51;
	input v_52;
	input v_53;
	input v_54;
	input v_55;
	input v_56;
	input v_57;
	input v_58;
	input v_59;
	input v_60;
	input v_61;
	input v_62;
	input v_63;
	input v_64;
	input v_65;
	input v_66;
	input v_67;
	input v_68;
	input v_69;
	input v_70;
	input v_71;
	input v_72;
	input v_73;
	input v_74;
	input v_75;
	input v_76;
	input v_77;
	input v_78;
	input v_79;
	input v_80;
	input v_81;
	input v_82;
	input v_83;
	input v_84;
	input v_85;
	input v_86;
	input v_87;
	input v_88;
	input v_89;
	input v_90;
	input v_91;
	input v_92;
	input v_93;
	input v_94;
	input v_95;
	input v_96;
	input v_97;
	input v_98;
	input v_99;
	input v_100;
	input v_101;
	input v_102;
	input v_103;
	input v_104;
	input v_105;
	input v_106;
	input v_107;
	input v_108;
	input v_109;
	input v_110;
	input v_111;
	input v_112;
	input v_113;
	input v_114;
	input v_115;
	input v_116;
	input v_117;
	input v_118;
	input v_119;
	input v_120;
	input v_121;
	input v_122;
	input v_123;
	input v_124;
	input v_125;
	input v_126;
	input v_127;
	input v_128;
	input v_129;
	input v_130;
	input v_131;
	input v_132;
	input v_133;
	input v_134;
	input v_135;
	input v_136;
	input v_137;
	input v_138;
	input v_139;
	input v_140;
	input v_141;
	input v_142;
	input v_143;
	input v_144;
	input v_145;
	input v_146;
	input v_147;
	input v_148;
	input v_149;
	input v_150;
	input v_151;
	input v_152;
	input v_153;
	input v_154;
	input v_155;
	input v_156;
	input v_157;
	input v_158;
	input v_159;
	input v_160;
	input v_161;
	input v_162;
	input v_163;
	input v_164;
	input v_165;
	input v_166;
	input v_167;
	input v_168;
	wire v_169;
	wire v_170;
	wire v_171;
	wire v_172;
	wire v_173;
	wire v_174;
	wire v_175;
	wire v_176;
	wire v_177;
	wire v_178;
	wire v_179;
	wire v_180;
	wire v_181;
	wire v_182;
	wire v_183;
	wire v_184;
	wire v_185;
	wire v_186;
	wire v_187;
	wire v_188;
	wire v_189;
	wire v_190;
	wire v_191;
	wire v_192;
	wire v_193;
	wire v_194;
	wire v_195;
	wire v_196;
	wire v_197;
	wire v_198;
	wire v_199;
	wire v_200;
	wire v_201;
	wire v_202;
	wire v_203;
	wire v_204;
	wire v_205;
	wire v_206;
	wire v_207;
	wire v_208;
	wire v_209;
	wire v_210;
	wire v_211;
	wire v_212;
	wire v_213;
	wire v_214;
	wire v_215;
	wire v_216;
	wire v_217;
	wire v_218;
	wire v_219;
	wire v_220;
	wire v_221;
	wire v_222;
	wire v_223;
	wire v_224;
	wire v_225;
	wire v_226;
	wire v_227;
	wire v_228;
	wire v_229;
	wire v_230;
	wire v_231;
	wire v_232;
	wire v_233;
	wire v_234;
	wire v_235;
	wire v_236;
	wire v_237;
	wire v_238;
	wire v_239;
	wire v_240;
	wire v_241;
	wire v_242;
	wire v_243;
	wire v_244;
	wire v_245;
	wire v_246;
	wire v_247;
	wire v_248;
	wire v_249;
	wire v_250;
	wire v_251;
	wire v_252;
	wire v_253;
	wire v_254;
	wire v_255;
	wire v_256;
	wire v_257;
	wire v_258;
	wire v_259;
	wire v_260;
	wire v_261;
	wire v_262;
	wire v_263;
	wire v_264;
	wire v_265;
	wire v_266;
	wire v_267;
	wire v_268;
	wire v_269;
	wire v_270;
	wire v_271;
	wire v_272;
	wire v_273;
	wire v_274;
	wire v_275;
	wire v_276;
	wire v_277;
	wire v_278;
	wire v_279;
	wire v_280;
	wire v_281;
	wire v_282;
	wire v_283;
	wire v_284;
	wire v_285;
	wire v_286;
	wire v_287;
	wire v_288;
	wire v_289;
	wire v_290;
	wire v_291;
	wire v_292;
	wire v_293;
	wire v_294;
	wire v_295;
	wire v_296;
	wire v_297;
	wire v_298;
	wire v_299;
	wire v_300;
	wire v_301;
	wire v_302;
	wire v_303;
	wire v_304;
	wire v_305;
	wire v_306;
	wire v_307;
	wire v_308;
	wire v_309;
	wire v_310;
	wire v_311;
	wire v_312;
	wire v_313;
	wire v_314;
	wire v_315;
	wire v_316;
	wire v_317;
	wire v_318;
	wire v_319;
	wire v_320;
	wire v_321;
	wire v_322;
	wire v_323;
	wire v_324;
	wire v_325;
	wire v_326;
	wire v_327;
	wire v_328;
	wire v_329;
	wire v_330;
	wire v_331;
	wire v_332;
	wire v_333;
	wire v_334;
	wire v_335;
	wire v_336;
	wire v_337;
	wire v_338;
	wire v_339;
	wire v_340;
	wire v_341;
	wire v_342;
	wire v_343;
	wire v_344;
	wire v_345;
	wire v_346;
	wire v_347;
	wire v_348;
	wire v_349;
	wire v_350;
	wire v_351;
	wire v_352;
	wire v_353;
	wire v_354;
	wire v_355;
	wire v_356;
	wire v_357;
	wire v_358;
	wire v_359;
	wire v_360;
	wire v_361;
	wire v_362;
	wire v_363;
	wire v_364;
	wire v_365;
	wire v_366;
	wire v_367;
	wire v_368;
	wire v_369;
	wire v_370;
	wire v_371;
	wire v_372;
	wire v_373;
	wire v_374;
	wire v_375;
	wire v_376;
	wire v_377;
	wire v_378;
	wire v_379;
	wire v_380;
	wire v_381;
	wire v_382;
	wire v_383;
	wire v_384;
	wire v_385;
	wire v_386;
	wire v_387;
	wire v_388;
	wire v_389;
	wire v_390;
	wire v_391;
	wire v_392;
	wire v_393;
	wire v_394;
	wire v_395;
	wire v_396;
	wire v_397;
	wire v_398;
	wire v_399;
	wire v_400;
	wire v_401;
	wire v_402;
	wire v_403;
	wire v_404;
	wire v_405;
	wire v_406;
	wire v_407;
	wire v_408;
	wire v_409;
	wire v_410;
	wire v_411;
	wire v_412;
	wire v_413;
	wire v_414;
	wire v_415;
	wire v_416;
	wire v_417;
	wire v_418;
	wire v_419;
	wire v_420;
	wire v_421;
	wire v_422;
	wire v_423;
	wire v_424;
	wire v_425;
	wire v_426;
	wire v_427;
	wire v_428;
	wire v_429;
	wire v_430;
	wire v_431;
	wire v_432;
	wire v_433;
	wire v_434;
	wire v_435;
	wire v_436;
	wire v_437;
	wire v_438;
	wire v_439;
	wire v_440;
	wire v_441;
	wire v_442;
	wire v_443;
	wire v_444;
	wire v_445;
	wire v_446;
	wire v_447;
	wire v_448;
	wire v_449;
	wire v_450;
	wire v_451;
	wire v_452;
	wire v_453;
	wire v_454;
	wire v_455;
	wire v_456;
	wire v_457;
	wire v_458;
	wire v_459;
	wire v_460;
	wire v_461;
	wire v_462;
	wire v_463;
	wire v_464;
	wire v_465;
	wire v_466;
	wire v_467;
	wire v_468;
	wire v_469;
	wire v_470;
	wire v_471;
	wire v_472;
	wire v_473;
	wire v_474;
	wire v_475;
	wire v_476;
	wire v_477;
	wire v_478;
	wire v_479;
	wire v_480;
	wire v_481;
	wire v_482;
	wire v_483;
	wire v_484;
	wire v_485;
	wire v_486;
	wire v_487;
	wire v_488;
	wire v_489;
	wire v_490;
	wire v_491;
	wire v_492;
	wire v_493;
	wire v_494;
	wire v_495;
	wire v_496;
	wire v_497;
	wire v_498;
	wire v_499;
	wire v_500;
	wire v_501;
	wire v_502;
	wire v_503;
	wire v_504;
	wire v_505;
	wire v_506;
	wire v_507;
	wire v_508;
	wire v_509;
	wire v_510;
	wire v_511;
	wire v_512;
	wire v_513;
	wire v_514;
	wire v_515;
	wire v_516;
	wire v_517;
	wire v_518;
	wire v_519;
	wire v_520;
	wire v_521;
	wire v_522;
	wire v_523;
	wire v_524;
	wire v_525;
	wire v_526;
	wire v_527;
	wire v_528;
	wire v_529;
	wire v_530;
	wire v_531;
	wire v_532;
	wire v_533;
	wire v_534;
	wire v_535;
	wire v_536;
	wire v_537;
	wire v_538;
	wire v_539;
	wire v_540;
	wire v_541;
	wire v_542;
	wire v_543;
	wire v_544;
	wire v_545;
	wire v_546;
	wire v_547;
	wire v_548;
	wire v_549;
	wire v_550;
	wire v_551;
	wire v_552;
	wire v_553;
	wire v_554;
	wire v_555;
	wire v_556;
	wire v_557;
	wire v_558;
	wire v_559;
	wire v_560;
	wire v_561;
	wire v_562;
	wire v_563;
	wire v_564;
	wire v_565;
	wire v_566;
	wire v_567;
	wire v_568;
	wire v_569;
	wire v_570;
	wire v_571;
	wire v_572;
	wire v_573;
	wire v_574;
	wire v_575;
	wire v_576;
	wire v_577;
	wire v_578;
	wire v_579;
	wire v_580;
	wire v_581;
	wire v_582;
	wire v_583;
	wire v_584;
	wire v_585;
	wire v_586;
	wire v_587;
	wire v_588;
	wire v_589;
	wire v_590;
	wire v_591;
	wire v_592;
	wire v_593;
	wire v_594;
	wire v_595;
	wire v_596;
	wire v_597;
	wire v_598;
	wire v_599;
	wire v_600;
	wire v_601;
	wire v_602;
	wire v_603;
	wire v_604;
	wire v_605;
	wire v_606;
	wire v_607;
	wire v_608;
	wire v_609;
	wire v_610;
	wire v_611;
	wire v_612;
	wire v_613;
	wire v_614;
	wire v_615;
	wire v_616;
	wire v_617;
	wire v_618;
	wire v_619;
	wire v_620;
	wire v_621;
	wire v_622;
	wire v_623;
	wire v_624;
	wire v_625;
	wire v_626;
	wire v_627;
	wire v_628;
	wire v_629;
	wire v_630;
	wire v_631;
	wire v_632;
	wire v_633;
	wire v_634;
	wire v_635;
	wire v_636;
	wire v_637;
	wire v_638;
	wire v_639;
	wire v_640;
	wire v_641;
	wire v_642;
	wire v_643;
	wire v_644;
	wire v_645;
	wire v_646;
	wire v_647;
	wire v_648;
	wire v_649;
	wire v_650;
	wire v_651;
	wire v_652;
	wire v_653;
	wire v_654;
	wire v_655;
	wire v_656;
	wire v_657;
	wire v_658;
	wire v_659;
	wire v_660;
	wire v_661;
	wire v_662;
	wire v_663;
	wire v_664;
	wire v_665;
	wire v_666;
	wire v_667;
	wire v_668;
	wire v_669;
	wire v_670;
	wire v_671;
	wire v_672;
	wire v_673;
	wire v_674;
	wire v_675;
	wire v_676;
	wire v_677;
	wire v_678;
	wire v_679;
	wire v_680;
	wire v_681;
	wire v_682;
	wire v_683;
	wire v_684;
	wire v_685;
	wire v_686;
	wire v_687;
	wire v_688;
	wire v_689;
	wire v_690;
	wire v_691;
	wire v_692;
	wire v_693;
	wire v_694;
	wire v_695;
	wire v_696;
	wire v_697;
	wire v_698;
	wire v_699;
	wire v_700;
	wire v_701;
	wire v_702;
	wire v_703;
	wire v_704;
	wire v_705;
	wire v_706;
	wire v_707;
	wire v_708;
	wire v_709;
	wire v_710;
	wire v_711;
	wire v_712;
	wire v_713;
	wire v_714;
	wire v_715;
	wire v_716;
	wire v_717;
	wire v_718;
	wire v_719;
	wire v_720;
	wire v_721;
	wire v_722;
	wire v_723;
	wire v_724;
	wire v_725;
	wire v_726;
	wire v_727;
	wire v_728;
	wire v_729;
	wire v_730;
	wire v_731;
	wire v_732;
	wire v_733;
	wire v_734;
	wire v_735;
	wire v_736;
	wire v_737;
	wire v_738;
	wire v_739;
	wire v_740;
	wire v_741;
	wire v_742;
	wire v_743;
	wire v_744;
	wire v_745;
	wire v_746;
	wire v_747;
	wire v_748;
	wire v_749;
	wire v_750;
	wire v_751;
	wire v_752;
	wire v_753;
	wire v_754;
	wire v_755;
	wire v_756;
	wire v_757;
	wire v_758;
	wire v_759;
	wire v_760;
	wire v_761;
	wire v_762;
	wire v_763;
	wire v_764;
	wire v_765;
	wire v_766;
	wire v_767;
	wire v_768;
	wire v_769;
	wire v_770;
	wire v_771;
	wire v_772;
	wire v_773;
	wire v_774;
	wire v_775;
	wire v_776;
	wire v_777;
	wire v_778;
	wire v_779;
	wire v_780;
	wire v_781;
	wire v_782;
	wire v_783;
	wire v_784;
	wire v_785;
	wire v_786;
	wire v_787;
	wire v_788;
	wire v_789;
	wire v_790;
	wire v_791;
	wire v_792;
	wire v_793;
	wire v_794;
	wire v_795;
	wire v_796;
	wire v_797;
	wire v_798;
	wire v_799;
	wire v_800;
	wire v_801;
	wire v_802;
	wire v_803;
	wire v_804;
	wire v_805;
	wire v_806;
	wire v_807;
	wire v_808;
	wire v_809;
	wire v_810;
	wire v_811;
	wire v_812;
	wire v_813;
	wire v_814;
	wire v_815;
	wire v_816;
	wire v_817;
	wire v_818;
	wire v_819;
	wire v_820;
	wire v_821;
	wire v_822;
	wire v_823;
	wire v_824;
	wire v_825;
	wire v_826;
	wire v_827;
	wire v_828;
	wire v_829;
	wire v_830;
	wire v_831;
	wire v_832;
	wire v_833;
	wire v_834;
	wire v_835;
	wire v_836;
	wire v_837;
	wire v_838;
	wire v_839;
	wire v_840;
	wire v_841;
	wire v_842;
	wire v_843;
	wire v_844;
	wire v_845;
	wire v_846;
	wire v_847;
	wire v_848;
	wire v_849;
	wire v_850;
	wire v_851;
	wire v_852;
	wire v_853;
	wire v_854;
	wire v_855;
	wire v_856;
	wire v_857;
	wire v_858;
	wire v_859;
	wire v_860;
	wire v_861;
	wire v_862;
	wire v_863;
	wire v_864;
	wire v_865;
	wire v_866;
	wire v_867;
	wire v_868;
	wire v_869;
	wire v_870;
	wire v_871;
	wire v_872;
	wire v_873;
	wire v_874;
	wire v_875;
	wire v_876;
	wire v_877;
	wire v_878;
	wire v_879;
	wire v_880;
	wire v_881;
	wire v_882;
	wire v_883;
	wire v_884;
	wire v_885;
	wire v_886;
	wire v_887;
	wire v_888;
	wire v_889;
	wire v_890;
	wire v_891;
	wire v_892;
	wire v_893;
	wire v_894;
	wire v_895;
	wire v_896;
	wire v_897;
	wire v_898;
	wire v_899;
	wire v_900;
	wire v_901;
	wire v_902;
	wire v_903;
	wire v_904;
	wire v_905;
	wire v_906;
	wire v_907;
	wire v_908;
	wire v_909;
	wire v_910;
	wire v_911;
	wire v_912;
	wire v_913;
	wire v_914;
	wire v_915;
	wire v_916;
	wire v_917;
	wire v_918;
	wire v_919;
	wire v_920;
	wire v_921;
	wire v_922;
	wire v_923;
	wire v_924;
	wire v_925;
	wire v_926;
	wire v_927;
	wire v_928;
	wire v_929;
	wire v_930;
	wire v_931;
	wire v_932;
	wire v_933;
	wire v_934;
	wire v_935;
	wire v_936;
	wire v_937;
	wire v_938;
	wire v_939;
	wire v_940;
	wire v_941;
	wire v_942;
	wire v_943;
	wire v_944;
	wire v_945;
	wire v_946;
	wire v_947;
	wire v_948;
	wire v_949;
	wire v_950;
	wire v_951;
	wire v_952;
	wire v_953;
	wire v_954;
	wire v_955;
	wire v_956;
	wire v_957;
	wire v_958;
	wire v_959;
	wire v_960;
	wire v_961;
	wire v_962;
	wire v_963;
	wire v_964;
	wire v_965;
	wire v_966;
	wire v_967;
	wire v_968;
	wire v_969;
	wire v_970;
	wire v_971;
	wire v_972;
	wire v_973;
	wire v_974;
	wire v_975;
	wire v_976;
	wire v_977;
	wire v_978;
	wire v_979;
	wire v_980;
	wire v_981;
	wire v_982;
	wire v_983;
	wire v_984;
	wire v_985;
	wire v_986;
	wire v_987;
	wire v_988;
	wire v_989;
	wire v_990;
	wire v_991;
	wire v_992;
	wire v_993;
	wire v_994;
	wire v_995;
	wire v_996;
	wire v_997;
	wire v_998;
	wire v_999;
	wire v_1000;
	wire v_1001;
	wire v_1002;
	wire v_1003;
	wire v_1004;
	wire v_1005;
	wire v_1006;
	wire v_1007;
	wire v_1008;
	wire v_1009;
	wire v_1010;
	wire v_1011;
	wire v_1012;
	wire v_1013;
	wire v_1014;
	wire v_1015;
	wire v_1016;
	wire v_1017;
	wire v_1018;
	wire v_1019;
	wire v_1020;
	wire v_1021;
	wire v_1022;
	wire v_1023;
	wire v_1024;
	wire v_1025;
	wire v_1026;
	wire v_1027;
	wire v_1028;
	wire v_1029;
	wire v_1030;
	wire v_1031;
	wire v_1032;
	wire v_1033;
	wire v_1034;
	wire v_1035;
	wire v_1036;
	wire v_1037;
	wire v_1038;
	wire v_1039;
	wire v_1040;
	wire v_1041;
	wire v_1042;
	wire v_1043;
	wire v_1044;
	wire v_1045;
	wire v_1046;
	wire v_1047;
	wire v_1048;
	wire v_1049;
	wire v_1050;
	wire v_1051;
	wire v_1052;
	wire v_1053;
	wire v_1054;
	wire v_1055;
	wire v_1056;
	wire v_1057;
	wire v_1058;
	wire v_1059;
	wire v_1060;
	wire v_1061;
	wire v_1062;
	wire v_1063;
	wire v_1064;
	wire v_1065;
	wire v_1066;
	wire v_1067;
	wire v_1068;
	wire v_1069;
	wire v_1070;
	wire v_1071;
	wire v_1072;
	wire v_1073;
	wire v_1074;
	wire v_1075;
	wire v_1076;
	wire v_1077;
	wire v_1078;
	wire v_1079;
	wire v_1080;
	wire v_1081;
	wire v_1082;
	wire v_1083;
	wire v_1084;
	wire v_1085;
	wire v_1086;
	wire v_1087;
	wire v_1088;
	wire v_1089;
	wire v_1090;
	wire v_1091;
	wire v_1092;
	wire v_1093;
	wire v_1094;
	wire v_1095;
	wire v_1096;
	wire v_1097;
	wire v_1098;
	wire v_1099;
	wire v_1100;
	wire v_1101;
	wire v_1102;
	wire v_1103;
	wire v_1104;
	wire v_1105;
	wire v_1106;
	wire v_1107;
	wire v_1108;
	wire v_1109;
	wire v_1110;
	wire v_1111;
	wire v_1112;
	wire v_1113;
	wire v_1114;
	wire v_1115;
	wire v_1116;
	wire v_1117;
	wire v_1118;
	wire v_1119;
	wire v_1120;
	wire v_1121;
	wire v_1122;
	wire v_1123;
	wire v_1124;
	wire v_1125;
	wire v_1126;
	wire v_1127;
	wire v_1128;
	wire v_1129;
	wire v_1130;
	wire v_1131;
	wire x_1;
	output o_1;
	assign v_989 = v_156 ;
	assign v_969 = v_153 ;
	assign v_945 = v_148 ;
	assign v_925 = v_145 ;
	assign v_901 = v_140 ;
	assign v_881 = v_137 ;
	assign v_857 = v_132 ;
	assign v_837 = v_129 ;
	assign v_813 = v_124 ;
	assign v_793 = v_121 ;
	assign v_769 = v_116 ;
	assign v_749 = v_113 ;
	assign v_725 = v_108 ;
	assign v_705 = v_105 ;
	assign v_681 = v_100 ;
	assign v_661 = v_97 ;
	assign v_637 = v_92 ;
	assign v_617 = v_89 ;
	assign v_589 = v_76 ;
	assign v_569 = v_73 ;
	assign v_545 = v_68 ;
	assign v_525 = v_65 ;
	assign v_501 = v_60 ;
	assign v_481 = v_57 ;
	assign v_457 = v_52 ;
	assign v_437 = v_49 ;
	assign v_413 = v_44 ;
	assign v_393 = v_41 ;
	assign v_369 = v_36 ;
	assign v_349 = v_33 ;
	assign v_325 = v_28 ;
	assign v_305 = v_25 ;
	assign v_281 = v_20 ;
	assign v_261 = v_17 ;
	assign v_237 = v_12 ;
	assign v_217 = v_9 ;
	assign v_193 = v_4 ;
	assign v_173 = v_1 ;
	assign v_991 = (v_157 & v_989) ;
	assign v_971 = (v_154 & v_969) ;
	assign v_947 = (v_149 & v_945) ;
	assign v_927 = (v_146 & v_925) ;
	assign v_903 = (v_141 & v_901) ;
	assign v_883 = (v_138 & v_881) ;
	assign v_859 = (v_133 & v_857) ;
	assign v_839 = (v_130 & v_837) ;
	assign v_815 = (v_125 & v_813) ;
	assign v_795 = (v_122 & v_793) ;
	assign v_771 = (v_117 & v_769) ;
	assign v_751 = (v_114 & v_749) ;
	assign v_727 = (v_109 & v_725) ;
	assign v_707 = (v_106 & v_705) ;
	assign v_683 = (v_101 & v_681) ;
	assign v_663 = (v_98 & v_661) ;
	assign v_639 = (v_93 & v_637) ;
	assign v_619 = (v_90 & v_617) ;
	assign v_591 = (v_77 & v_589) ;
	assign v_571 = (v_74 & v_569) ;
	assign v_547 = (v_69 & v_545) ;
	assign v_527 = (v_66 & v_525) ;
	assign v_503 = (v_61 & v_501) ;
	assign v_483 = (v_58 & v_481) ;
	assign v_459 = (v_53 & v_457) ;
	assign v_439 = (v_50 & v_437) ;
	assign v_415 = (v_45 & v_413) ;
	assign v_395 = (v_42 & v_393) ;
	assign v_371 = (v_37 & v_369) ;
	assign v_351 = (v_34 & v_349) ;
	assign v_327 = (v_29 & v_325) ;
	assign v_307 = (v_26 & v_305) ;
	assign v_283 = (v_21 & v_281) ;
	assign v_263 = (v_18 & v_261) ;
	assign v_239 = (v_13 & v_237) ;
	assign v_219 = (v_10 & v_217) ;
	assign v_195 = (v_5 & v_193) ;
	assign v_175 = (v_2 & v_173) ;
	assign v_992 = v_991 ;
	assign v_972 = v_971 ;
	assign v_948 = v_947 ;
	assign v_928 = v_927 ;
	assign v_904 = v_903 ;
	assign v_884 = v_883 ;
	assign v_860 = v_859 ;
	assign v_840 = v_839 ;
	assign v_816 = v_815 ;
	assign v_796 = v_795 ;
	assign v_772 = v_771 ;
	assign v_752 = v_751 ;
	assign v_728 = v_727 ;
	assign v_708 = v_707 ;
	assign v_684 = v_683 ;
	assign v_664 = v_663 ;
	assign v_640 = v_639 ;
	assign v_620 = v_619 ;
	assign v_592 = v_591 ;
	assign v_572 = v_571 ;
	assign v_548 = v_547 ;
	assign v_528 = v_527 ;
	assign v_504 = v_503 ;
	assign v_484 = v_483 ;
	assign v_460 = v_459 ;
	assign v_440 = v_439 ;
	assign v_416 = v_415 ;
	assign v_396 = v_395 ;
	assign v_372 = v_371 ;
	assign v_352 = v_351 ;
	assign v_328 = v_327 ;
	assign v_308 = v_307 ;
	assign v_284 = v_283 ;
	assign v_264 = v_263 ;
	assign v_240 = v_239 ;
	assign v_220 = v_219 ;
	assign v_196 = v_195 ;
	assign v_176 = v_175 ;
	assign v_993 = (v_992 ^ v_158) ;
	assign v_968 = (v_160 ^ v_159) ;
	assign v_990 = (v_989 ^ v_157) ;
	assign v_973 = (v_972 ^ v_155) ;
	assign v_970 = (v_969 ^ v_154) ;
	assign v_949 = (v_948 ^ v_150) ;
	assign v_924 = (v_152 ^ v_151) ;
	assign v_946 = (v_945 ^ v_149) ;
	assign v_929 = (v_928 ^ v_147) ;
	assign v_926 = (v_925 ^ v_146) ;
	assign v_905 = (v_904 ^ v_142) ;
	assign v_880 = (v_144 ^ v_143) ;
	assign v_902 = (v_901 ^ v_141) ;
	assign v_885 = (v_884 ^ v_139) ;
	assign v_882 = (v_881 ^ v_138) ;
	assign v_861 = (v_860 ^ v_134) ;
	assign v_836 = (v_136 ^ v_135) ;
	assign v_858 = (v_857 ^ v_133) ;
	assign v_841 = (v_840 ^ v_131) ;
	assign v_838 = (v_837 ^ v_130) ;
	assign v_817 = (v_816 ^ v_126) ;
	assign v_792 = (v_128 ^ v_127) ;
	assign v_814 = (v_813 ^ v_125) ;
	assign v_797 = (v_796 ^ v_123) ;
	assign v_794 = (v_793 ^ v_122) ;
	assign v_773 = (v_772 ^ v_118) ;
	assign v_748 = (v_120 ^ v_119) ;
	assign v_770 = (v_769 ^ v_117) ;
	assign v_753 = (v_752 ^ v_115) ;
	assign v_750 = (v_749 ^ v_114) ;
	assign v_729 = (v_728 ^ v_110) ;
	assign v_704 = (v_112 ^ v_111) ;
	assign v_726 = (v_725 ^ v_109) ;
	assign v_709 = (v_708 ^ v_107) ;
	assign v_706 = (v_705 ^ v_106) ;
	assign v_685 = (v_684 ^ v_102) ;
	assign v_660 = (v_104 ^ v_103) ;
	assign v_682 = (v_681 ^ v_101) ;
	assign v_665 = (v_664 ^ v_99) ;
	assign v_662 = (v_661 ^ v_98) ;
	assign v_641 = (v_640 ^ v_94) ;
	assign v_616 = (v_96 ^ v_95) ;
	assign v_638 = (v_637 ^ v_93) ;
	assign v_621 = (v_620 ^ v_91) ;
	assign v_618 = (v_617 ^ v_90) ;
	assign v_593 = (v_592 ^ v_78) ;
	assign v_568 = (v_80 ^ v_79) ;
	assign v_590 = (v_589 ^ v_77) ;
	assign v_573 = (v_572 ^ v_75) ;
	assign v_570 = (v_569 ^ v_74) ;
	assign v_549 = (v_548 ^ v_70) ;
	assign v_524 = (v_72 ^ v_71) ;
	assign v_546 = (v_545 ^ v_69) ;
	assign v_529 = (v_528 ^ v_67) ;
	assign v_526 = (v_525 ^ v_66) ;
	assign v_505 = (v_504 ^ v_62) ;
	assign v_480 = (v_64 ^ v_63) ;
	assign v_502 = (v_501 ^ v_61) ;
	assign v_485 = (v_484 ^ v_59) ;
	assign v_482 = (v_481 ^ v_58) ;
	assign v_461 = (v_460 ^ v_54) ;
	assign v_436 = (v_56 ^ v_55) ;
	assign v_458 = (v_457 ^ v_53) ;
	assign v_441 = (v_440 ^ v_51) ;
	assign v_438 = (v_437 ^ v_50) ;
	assign v_417 = (v_416 ^ v_46) ;
	assign v_392 = (v_48 ^ v_47) ;
	assign v_414 = (v_413 ^ v_45) ;
	assign v_397 = (v_396 ^ v_43) ;
	assign v_394 = (v_393 ^ v_42) ;
	assign v_373 = (v_372 ^ v_38) ;
	assign v_348 = (v_40 ^ v_39) ;
	assign v_370 = (v_369 ^ v_37) ;
	assign v_353 = (v_352 ^ v_35) ;
	assign v_350 = (v_349 ^ v_34) ;
	assign v_329 = (v_328 ^ v_30) ;
	assign v_304 = (v_32 ^ v_31) ;
	assign v_326 = (v_325 ^ v_29) ;
	assign v_309 = (v_308 ^ v_27) ;
	assign v_306 = (v_305 ^ v_26) ;
	assign v_285 = (v_284 ^ v_22) ;
	assign v_260 = (v_24 ^ v_23) ;
	assign v_282 = (v_281 ^ v_21) ;
	assign v_265 = (v_264 ^ v_19) ;
	assign v_262 = (v_261 ^ v_18) ;
	assign v_241 = (v_240 ^ v_14) ;
	assign v_216 = (v_16 ^ v_15) ;
	assign v_238 = (v_237 ^ v_13) ;
	assign v_221 = (v_220 ^ v_11) ;
	assign v_218 = (v_217 ^ v_10) ;
	assign v_197 = (v_196 ^ v_6) ;
	assign v_172 = (v_8 ^ v_7) ;
	assign v_194 = (v_193 ^ v_5) ;
	assign v_177 = (v_176 ^ v_3) ;
	assign v_174 = (v_173 ^ v_2) ;
	assign v_1003 = (v_968 & v_993) ;
	assign v_1002 = (~v_968 & v_158) ;
	assign v_1000 = (v_968 & v_990) ;
	assign v_999 = (~v_968 & v_157) ;
	assign v_997 = (~v_156 & v_968) ;
	assign v_996 = (~v_968 & v_156) ;
	assign v_983 = (v_968 & v_155) ;
	assign v_982 = (~v_968 & v_973) ;
	assign v_980 = (v_968 & v_154) ;
	assign v_979 = (~v_968 & v_970) ;
	assign v_977 = (v_968 & v_153) ;
	assign v_976 = (~v_968 & ~v_153) ;
	assign v_959 = (v_924 & v_949) ;
	assign v_958 = (~v_924 & v_150) ;
	assign v_956 = (v_924 & v_946) ;
	assign v_955 = (~v_924 & v_149) ;
	assign v_953 = (~v_148 & v_924) ;
	assign v_952 = (~v_924 & v_148) ;
	assign v_939 = (v_924 & v_147) ;
	assign v_938 = (~v_924 & v_929) ;
	assign v_936 = (v_924 & v_146) ;
	assign v_935 = (~v_924 & v_926) ;
	assign v_933 = (v_924 & v_145) ;
	assign v_932 = (~v_924 & ~v_145) ;
	assign v_915 = (v_880 & v_905) ;
	assign v_914 = (~v_880 & v_142) ;
	assign v_912 = (v_880 & v_902) ;
	assign v_911 = (~v_880 & v_141) ;
	assign v_909 = (~v_140 & v_880) ;
	assign v_908 = (~v_880 & v_140) ;
	assign v_895 = (v_880 & v_139) ;
	assign v_894 = (~v_880 & v_885) ;
	assign v_892 = (v_880 & v_138) ;
	assign v_891 = (~v_880 & v_882) ;
	assign v_889 = (v_880 & v_137) ;
	assign v_888 = (~v_880 & ~v_137) ;
	assign v_871 = (v_836 & v_861) ;
	assign v_870 = (~v_836 & v_134) ;
	assign v_868 = (v_836 & v_858) ;
	assign v_867 = (~v_836 & v_133) ;
	assign v_865 = (~v_132 & v_836) ;
	assign v_864 = (~v_836 & v_132) ;
	assign v_851 = (v_836 & v_131) ;
	assign v_850 = (~v_836 & v_841) ;
	assign v_848 = (v_836 & v_130) ;
	assign v_847 = (~v_836 & v_838) ;
	assign v_845 = (v_836 & v_129) ;
	assign v_844 = (~v_836 & ~v_129) ;
	assign v_827 = (v_792 & v_817) ;
	assign v_826 = (~v_792 & v_126) ;
	assign v_824 = (v_792 & v_814) ;
	assign v_823 = (~v_792 & v_125) ;
	assign v_821 = (~v_124 & v_792) ;
	assign v_820 = (~v_792 & v_124) ;
	assign v_807 = (v_792 & v_123) ;
	assign v_806 = (~v_792 & v_797) ;
	assign v_804 = (v_792 & v_122) ;
	assign v_803 = (~v_792 & v_794) ;
	assign v_801 = (v_792 & v_121) ;
	assign v_800 = (~v_792 & ~v_121) ;
	assign v_783 = (v_748 & v_773) ;
	assign v_782 = (~v_748 & v_118) ;
	assign v_780 = (v_748 & v_770) ;
	assign v_779 = (~v_748 & v_117) ;
	assign v_777 = (~v_116 & v_748) ;
	assign v_776 = (~v_748 & v_116) ;
	assign v_763 = (v_748 & v_115) ;
	assign v_762 = (~v_748 & v_753) ;
	assign v_760 = (v_748 & v_114) ;
	assign v_759 = (~v_748 & v_750) ;
	assign v_757 = (v_748 & v_113) ;
	assign v_756 = (~v_748 & ~v_113) ;
	assign v_739 = (v_704 & v_729) ;
	assign v_738 = (~v_704 & v_110) ;
	assign v_736 = (v_704 & v_726) ;
	assign v_735 = (~v_704 & v_109) ;
	assign v_733 = (~v_108 & v_704) ;
	assign v_732 = (~v_704 & v_108) ;
	assign v_719 = (v_704 & v_107) ;
	assign v_718 = (~v_704 & v_709) ;
	assign v_716 = (v_704 & v_106) ;
	assign v_715 = (~v_704 & v_706) ;
	assign v_713 = (v_704 & v_105) ;
	assign v_712 = (~v_704 & ~v_105) ;
	assign v_695 = (v_660 & v_685) ;
	assign v_694 = (~v_660 & v_102) ;
	assign v_692 = (v_660 & v_682) ;
	assign v_691 = (~v_660 & v_101) ;
	assign v_689 = (~v_100 & v_660) ;
	assign v_688 = (~v_660 & v_100) ;
	assign v_675 = (v_660 & v_99) ;
	assign v_674 = (~v_660 & v_665) ;
	assign v_672 = (v_660 & v_98) ;
	assign v_671 = (~v_660 & v_662) ;
	assign v_669 = (v_660 & v_97) ;
	assign v_668 = (~v_660 & ~v_97) ;
	assign v_651 = (v_616 & v_641) ;
	assign v_650 = (~v_616 & v_94) ;
	assign v_648 = (v_616 & v_638) ;
	assign v_647 = (~v_616 & v_93) ;
	assign v_645 = (~v_92 & v_616) ;
	assign v_644 = (~v_616 & v_92) ;
	assign v_631 = (v_616 & v_91) ;
	assign v_630 = (~v_616 & v_621) ;
	assign v_628 = (v_616 & v_90) ;
	assign v_627 = (~v_616 & v_618) ;
	assign v_625 = (v_616 & v_89) ;
	assign v_624 = (~v_616 & ~v_89) ;
	assign v_603 = (v_568 & v_593) ;
	assign v_602 = (~v_568 & v_78) ;
	assign v_600 = (v_568 & v_590) ;
	assign v_599 = (~v_568 & v_77) ;
	assign v_597 = (~v_76 & v_568) ;
	assign v_596 = (~v_568 & v_76) ;
	assign v_583 = (v_568 & v_75) ;
	assign v_582 = (~v_568 & v_573) ;
	assign v_580 = (v_568 & v_74) ;
	assign v_579 = (~v_568 & v_570) ;
	assign v_577 = (v_568 & v_73) ;
	assign v_576 = (~v_568 & ~v_73) ;
	assign v_559 = (v_524 & v_549) ;
	assign v_558 = (~v_524 & v_70) ;
	assign v_556 = (v_524 & v_546) ;
	assign v_555 = (~v_524 & v_69) ;
	assign v_553 = (~v_68 & v_524) ;
	assign v_552 = (~v_524 & v_68) ;
	assign v_539 = (v_524 & v_67) ;
	assign v_538 = (~v_524 & v_529) ;
	assign v_536 = (v_524 & v_66) ;
	assign v_535 = (~v_524 & v_526) ;
	assign v_533 = (v_524 & v_65) ;
	assign v_532 = (~v_524 & ~v_65) ;
	assign v_515 = (v_480 & v_505) ;
	assign v_514 = (~v_480 & v_62) ;
	assign v_512 = (v_480 & v_502) ;
	assign v_511 = (~v_480 & v_61) ;
	assign v_509 = (~v_60 & v_480) ;
	assign v_508 = (~v_480 & v_60) ;
	assign v_495 = (v_480 & v_59) ;
	assign v_494 = (~v_480 & v_485) ;
	assign v_492 = (v_480 & v_58) ;
	assign v_491 = (~v_480 & v_482) ;
	assign v_489 = (v_480 & v_57) ;
	assign v_488 = (~v_480 & ~v_57) ;
	assign v_471 = (v_436 & v_461) ;
	assign v_470 = (~v_436 & v_54) ;
	assign v_468 = (v_436 & v_458) ;
	assign v_467 = (~v_436 & v_53) ;
	assign v_465 = (~v_52 & v_436) ;
	assign v_464 = (~v_436 & v_52) ;
	assign v_451 = (v_436 & v_51) ;
	assign v_450 = (~v_436 & v_441) ;
	assign v_448 = (v_436 & v_50) ;
	assign v_447 = (~v_436 & v_438) ;
	assign v_445 = (v_436 & v_49) ;
	assign v_444 = (~v_436 & ~v_49) ;
	assign v_427 = (v_392 & v_417) ;
	assign v_426 = (~v_392 & v_46) ;
	assign v_424 = (v_392 & v_414) ;
	assign v_423 = (~v_392 & v_45) ;
	assign v_421 = (~v_44 & v_392) ;
	assign v_420 = (~v_392 & v_44) ;
	assign v_407 = (v_392 & v_43) ;
	assign v_406 = (~v_392 & v_397) ;
	assign v_404 = (v_392 & v_42) ;
	assign v_403 = (~v_392 & v_394) ;
	assign v_401 = (v_392 & v_41) ;
	assign v_400 = (~v_392 & ~v_41) ;
	assign v_383 = (v_348 & v_373) ;
	assign v_382 = (~v_348 & v_38) ;
	assign v_380 = (v_348 & v_370) ;
	assign v_379 = (~v_348 & v_37) ;
	assign v_377 = (~v_36 & v_348) ;
	assign v_376 = (~v_348 & v_36) ;
	assign v_363 = (v_348 & v_35) ;
	assign v_362 = (~v_348 & v_353) ;
	assign v_360 = (v_348 & v_34) ;
	assign v_359 = (~v_348 & v_350) ;
	assign v_357 = (v_348 & v_33) ;
	assign v_356 = (~v_348 & ~v_33) ;
	assign v_339 = (v_304 & v_329) ;
	assign v_338 = (~v_304 & v_30) ;
	assign v_336 = (v_304 & v_326) ;
	assign v_335 = (~v_304 & v_29) ;
	assign v_333 = (~v_28 & v_304) ;
	assign v_332 = (~v_304 & v_28) ;
	assign v_319 = (v_304 & v_27) ;
	assign v_318 = (~v_304 & v_309) ;
	assign v_316 = (v_304 & v_26) ;
	assign v_315 = (~v_304 & v_306) ;
	assign v_313 = (v_304 & v_25) ;
	assign v_312 = (~v_304 & ~v_25) ;
	assign v_295 = (v_260 & v_285) ;
	assign v_294 = (~v_260 & v_22) ;
	assign v_292 = (v_260 & v_282) ;
	assign v_291 = (~v_260 & v_21) ;
	assign v_289 = (~v_20 & v_260) ;
	assign v_288 = (~v_260 & v_20) ;
	assign v_275 = (v_260 & v_19) ;
	assign v_274 = (~v_260 & v_265) ;
	assign v_272 = (v_260 & v_18) ;
	assign v_271 = (~v_260 & v_262) ;
	assign v_269 = (v_260 & v_17) ;
	assign v_268 = (~v_260 & ~v_17) ;
	assign v_251 = (v_216 & v_241) ;
	assign v_250 = (~v_216 & v_14) ;
	assign v_248 = (v_216 & v_238) ;
	assign v_247 = (~v_216 & v_13) ;
	assign v_245 = (~v_12 & v_216) ;
	assign v_244 = (~v_216 & v_12) ;
	assign v_231 = (v_216 & v_11) ;
	assign v_230 = (~v_216 & v_221) ;
	assign v_228 = (v_216 & v_10) ;
	assign v_227 = (~v_216 & v_218) ;
	assign v_225 = (v_216 & v_9) ;
	assign v_224 = (~v_216 & ~v_9) ;
	assign v_207 = (v_172 & v_197) ;
	assign v_206 = (~v_172 & v_6) ;
	assign v_204 = (v_172 & v_194) ;
	assign v_203 = (~v_172 & v_5) ;
	assign v_201 = (~v_4 & v_172) ;
	assign v_200 = (~v_172 & v_4) ;
	assign v_187 = (v_172 & v_3) ;
	assign v_186 = (~v_172 & v_177) ;
	assign v_184 = (v_172 & v_2) ;
	assign v_183 = (~v_172 & v_174) ;
	assign v_181 = (v_172 & v_1) ;
	assign v_180 = (~v_172 & ~v_1) ;
	assign v_1004 = (v_1002 | v_1003) ;
	assign v_1001 = (v_999 | v_1000) ;
	assign v_998 = (v_996 | v_997) ;
	assign v_984 = (v_982 | v_983) ;
	assign v_981 = (v_979 | v_980) ;
	assign v_978 = (v_976 | v_977) ;
	assign v_960 = (v_958 | v_959) ;
	assign v_957 = (v_955 | v_956) ;
	assign v_954 = (v_952 | v_953) ;
	assign v_940 = (v_938 | v_939) ;
	assign v_937 = (v_935 | v_936) ;
	assign v_934 = (v_932 | v_933) ;
	assign v_916 = (v_914 | v_915) ;
	assign v_913 = (v_911 | v_912) ;
	assign v_910 = (v_908 | v_909) ;
	assign v_896 = (v_894 | v_895) ;
	assign v_893 = (v_891 | v_892) ;
	assign v_890 = (v_888 | v_889) ;
	assign v_872 = (v_870 | v_871) ;
	assign v_869 = (v_867 | v_868) ;
	assign v_866 = (v_864 | v_865) ;
	assign v_852 = (v_850 | v_851) ;
	assign v_849 = (v_847 | v_848) ;
	assign v_846 = (v_844 | v_845) ;
	assign v_828 = (v_826 | v_827) ;
	assign v_825 = (v_823 | v_824) ;
	assign v_822 = (v_820 | v_821) ;
	assign v_808 = (v_806 | v_807) ;
	assign v_805 = (v_803 | v_804) ;
	assign v_802 = (v_800 | v_801) ;
	assign v_784 = (v_782 | v_783) ;
	assign v_781 = (v_779 | v_780) ;
	assign v_778 = (v_776 | v_777) ;
	assign v_764 = (v_762 | v_763) ;
	assign v_761 = (v_759 | v_760) ;
	assign v_758 = (v_756 | v_757) ;
	assign v_740 = (v_738 | v_739) ;
	assign v_737 = (v_735 | v_736) ;
	assign v_734 = (v_732 | v_733) ;
	assign v_720 = (v_718 | v_719) ;
	assign v_717 = (v_715 | v_716) ;
	assign v_714 = (v_712 | v_713) ;
	assign v_696 = (v_694 | v_695) ;
	assign v_693 = (v_691 | v_692) ;
	assign v_690 = (v_688 | v_689) ;
	assign v_676 = (v_674 | v_675) ;
	assign v_673 = (v_671 | v_672) ;
	assign v_670 = (v_668 | v_669) ;
	assign v_652 = (v_650 | v_651) ;
	assign v_649 = (v_647 | v_648) ;
	assign v_646 = (v_644 | v_645) ;
	assign v_632 = (v_630 | v_631) ;
	assign v_629 = (v_627 | v_628) ;
	assign v_626 = (v_624 | v_625) ;
	assign v_604 = (v_602 | v_603) ;
	assign v_601 = (v_599 | v_600) ;
	assign v_598 = (v_596 | v_597) ;
	assign v_584 = (v_582 | v_583) ;
	assign v_581 = (v_579 | v_580) ;
	assign v_578 = (v_576 | v_577) ;
	assign v_560 = (v_558 | v_559) ;
	assign v_557 = (v_555 | v_556) ;
	assign v_554 = (v_552 | v_553) ;
	assign v_540 = (v_538 | v_539) ;
	assign v_537 = (v_535 | v_536) ;
	assign v_534 = (v_532 | v_533) ;
	assign v_516 = (v_514 | v_515) ;
	assign v_513 = (v_511 | v_512) ;
	assign v_510 = (v_508 | v_509) ;
	assign v_496 = (v_494 | v_495) ;
	assign v_493 = (v_491 | v_492) ;
	assign v_490 = (v_488 | v_489) ;
	assign v_472 = (v_470 | v_471) ;
	assign v_469 = (v_467 | v_468) ;
	assign v_466 = (v_464 | v_465) ;
	assign v_452 = (v_450 | v_451) ;
	assign v_449 = (v_447 | v_448) ;
	assign v_446 = (v_444 | v_445) ;
	assign v_428 = (v_426 | v_427) ;
	assign v_425 = (v_423 | v_424) ;
	assign v_422 = (v_420 | v_421) ;
	assign v_408 = (v_406 | v_407) ;
	assign v_405 = (v_403 | v_404) ;
	assign v_402 = (v_400 | v_401) ;
	assign v_384 = (v_382 | v_383) ;
	assign v_381 = (v_379 | v_380) ;
	assign v_378 = (v_376 | v_377) ;
	assign v_364 = (v_362 | v_363) ;
	assign v_361 = (v_359 | v_360) ;
	assign v_358 = (v_356 | v_357) ;
	assign v_340 = (v_338 | v_339) ;
	assign v_337 = (v_335 | v_336) ;
	assign v_334 = (v_332 | v_333) ;
	assign v_320 = (v_318 | v_319) ;
	assign v_317 = (v_315 | v_316) ;
	assign v_314 = (v_312 | v_313) ;
	assign v_296 = (v_294 | v_295) ;
	assign v_293 = (v_291 | v_292) ;
	assign v_290 = (v_288 | v_289) ;
	assign v_276 = (v_274 | v_275) ;
	assign v_273 = (v_271 | v_272) ;
	assign v_270 = (v_268 | v_269) ;
	assign v_252 = (v_250 | v_251) ;
	assign v_249 = (v_247 | v_248) ;
	assign v_246 = (v_244 | v_245) ;
	assign v_232 = (v_230 | v_231) ;
	assign v_229 = (v_227 | v_228) ;
	assign v_226 = (v_224 | v_225) ;
	assign v_208 = (v_206 | v_207) ;
	assign v_205 = (v_203 | v_204) ;
	assign v_202 = (v_200 | v_201) ;
	assign v_188 = (v_186 | v_187) ;
	assign v_185 = (v_183 | v_184) ;
	assign v_182 = (v_180 | v_181) ;
	assign v_1118 = (v_166 ^ v_86) ;
	assign v_1117 = (v_165 ^ v_85) ;
	assign v_1116 = (v_164 ^ v_84) ;
	assign v_1114 = (v_163 ^ v_83) ;
	assign v_1113 = (v_162 ^ v_82) ;
	assign v_1112 = (v_161 ^ v_81) ;
	assign v_1107 = (v_158 ^ v_86) ;
	assign v_1106 = (v_157 ^ v_85) ;
	assign v_1105 = (v_156 ^ v_84) ;
	assign v_1103 = (v_155 ^ v_83) ;
	assign v_1102 = (v_154 ^ v_82) ;
	assign v_1101 = (v_153 ^ v_81) ;
	assign v_1096 = (v_150 ^ v_86) ;
	assign v_1095 = (v_149 ^ v_85) ;
	assign v_1094 = (v_148 ^ v_84) ;
	assign v_1092 = (v_147 ^ v_83) ;
	assign v_1091 = (v_146 ^ v_82) ;
	assign v_1090 = (v_145 ^ v_81) ;
	assign v_1085 = (v_142 ^ v_86) ;
	assign v_1084 = (v_141 ^ v_85) ;
	assign v_1083 = (v_140 ^ v_84) ;
	assign v_1081 = (v_139 ^ v_83) ;
	assign v_1080 = (v_138 ^ v_82) ;
	assign v_1079 = (v_137 ^ v_81) ;
	assign v_1074 = (v_134 ^ v_86) ;
	assign v_1073 = (v_133 ^ v_85) ;
	assign v_1072 = (v_132 ^ v_84) ;
	assign v_1070 = (v_131 ^ v_83) ;
	assign v_1069 = (v_130 ^ v_82) ;
	assign v_1068 = (v_129 ^ v_81) ;
	assign v_1063 = (v_126 ^ v_86) ;
	assign v_1062 = (v_125 ^ v_85) ;
	assign v_1061 = (v_124 ^ v_84) ;
	assign v_1059 = (v_123 ^ v_83) ;
	assign v_1058 = (v_122 ^ v_82) ;
	assign v_1057 = (v_121 ^ v_81) ;
	assign v_1052 = (v_118 ^ v_86) ;
	assign v_1051 = (v_117 ^ v_85) ;
	assign v_1050 = (v_116 ^ v_84) ;
	assign v_1048 = (v_115 ^ v_83) ;
	assign v_1047 = (v_114 ^ v_82) ;
	assign v_1046 = (v_113 ^ v_81) ;
	assign v_1041 = (v_110 ^ v_86) ;
	assign v_1040 = (v_109 ^ v_85) ;
	assign v_1039 = (v_108 ^ v_84) ;
	assign v_1037 = (v_107 ^ v_83) ;
	assign v_1036 = (v_106 ^ v_82) ;
	assign v_1035 = (v_105 ^ v_81) ;
	assign v_1030 = (v_102 ^ v_86) ;
	assign v_1029 = (v_101 ^ v_85) ;
	assign v_1028 = (v_100 ^ v_84) ;
	assign v_1026 = (v_99 ^ v_83) ;
	assign v_1025 = (v_98 ^ v_82) ;
	assign v_1024 = (v_97 ^ v_81) ;
	assign v_1019 = (v_94 ^ v_86) ;
	assign v_1018 = (v_93 ^ v_85) ;
	assign v_1017 = (v_92 ^ v_84) ;
	assign v_1015 = (v_91 ^ v_83) ;
	assign v_1014 = (v_90 ^ v_82) ;
	assign v_1013 = (v_89 ^ v_81) ;
	assign v_1007 = (v_1004 ^ v_166) ;
	assign v_1006 = (v_1001 ^ v_165) ;
	assign v_1005 = (v_998 ^ v_164) ;
	assign v_987 = (v_984 ^ v_163) ;
	assign v_986 = (v_981 ^ v_162) ;
	assign v_985 = (v_978 ^ v_161) ;
	assign v_963 = (v_960 ^ v_158) ;
	assign v_962 = (v_957 ^ v_157) ;
	assign v_961 = (v_954 ^ v_156) ;
	assign v_943 = (v_940 ^ v_155) ;
	assign v_942 = (v_937 ^ v_154) ;
	assign v_941 = (v_934 ^ v_153) ;
	assign v_919 = (v_916 ^ v_150) ;
	assign v_918 = (v_913 ^ v_149) ;
	assign v_917 = (v_910 ^ v_148) ;
	assign v_899 = (v_896 ^ v_147) ;
	assign v_898 = (v_893 ^ v_146) ;
	assign v_897 = (v_890 ^ v_145) ;
	assign v_875 = (v_872 ^ v_142) ;
	assign v_874 = (v_869 ^ v_141) ;
	assign v_873 = (v_866 ^ v_140) ;
	assign v_855 = (v_852 ^ v_139) ;
	assign v_854 = (v_849 ^ v_138) ;
	assign v_853 = (v_846 ^ v_137) ;
	assign v_831 = (v_828 ^ v_134) ;
	assign v_830 = (v_825 ^ v_133) ;
	assign v_829 = (v_822 ^ v_132) ;
	assign v_811 = (v_808 ^ v_131) ;
	assign v_810 = (v_805 ^ v_130) ;
	assign v_809 = (v_802 ^ v_129) ;
	assign v_787 = (v_784 ^ v_126) ;
	assign v_786 = (v_781 ^ v_125) ;
	assign v_785 = (v_778 ^ v_124) ;
	assign v_767 = (v_764 ^ v_123) ;
	assign v_766 = (v_761 ^ v_122) ;
	assign v_765 = (v_758 ^ v_121) ;
	assign v_743 = (v_740 ^ v_118) ;
	assign v_742 = (v_737 ^ v_117) ;
	assign v_741 = (v_734 ^ v_116) ;
	assign v_723 = (v_720 ^ v_115) ;
	assign v_722 = (v_717 ^ v_114) ;
	assign v_721 = (v_714 ^ v_113) ;
	assign v_699 = (v_696 ^ v_110) ;
	assign v_698 = (v_693 ^ v_109) ;
	assign v_697 = (v_690 ^ v_108) ;
	assign v_679 = (v_676 ^ v_107) ;
	assign v_678 = (v_673 ^ v_106) ;
	assign v_677 = (v_670 ^ v_105) ;
	assign v_655 = (v_652 ^ v_102) ;
	assign v_654 = (v_649 ^ v_101) ;
	assign v_653 = (v_646 ^ v_100) ;
	assign v_635 = (v_632 ^ v_99) ;
	assign v_634 = (v_629 ^ v_98) ;
	assign v_633 = (v_626 ^ v_97) ;
	assign v_607 = (v_604 ^ v_86) ;
	assign v_606 = (v_601 ^ v_85) ;
	assign v_605 = (v_598 ^ v_84) ;
	assign v_587 = (v_584 ^ v_83) ;
	assign v_586 = (v_581 ^ v_82) ;
	assign v_585 = (v_578 ^ v_81) ;
	assign v_563 = (v_560 ^ v_78) ;
	assign v_562 = (v_557 ^ v_77) ;
	assign v_561 = (v_554 ^ v_76) ;
	assign v_543 = (v_540 ^ v_75) ;
	assign v_542 = (v_537 ^ v_74) ;
	assign v_541 = (v_534 ^ v_73) ;
	assign v_519 = (v_516 ^ v_70) ;
	assign v_518 = (v_513 ^ v_69) ;
	assign v_517 = (v_510 ^ v_68) ;
	assign v_499 = (v_496 ^ v_67) ;
	assign v_498 = (v_493 ^ v_66) ;
	assign v_497 = (v_490 ^ v_65) ;
	assign v_475 = (v_472 ^ v_62) ;
	assign v_474 = (v_469 ^ v_61) ;
	assign v_473 = (v_466 ^ v_60) ;
	assign v_455 = (v_452 ^ v_59) ;
	assign v_454 = (v_449 ^ v_58) ;
	assign v_453 = (v_446 ^ v_57) ;
	assign v_431 = (v_428 ^ v_54) ;
	assign v_430 = (v_425 ^ v_53) ;
	assign v_429 = (v_422 ^ v_52) ;
	assign v_411 = (v_408 ^ v_51) ;
	assign v_410 = (v_405 ^ v_50) ;
	assign v_409 = (v_402 ^ v_49) ;
	assign v_387 = (v_384 ^ v_46) ;
	assign v_386 = (v_381 ^ v_45) ;
	assign v_385 = (v_378 ^ v_44) ;
	assign v_367 = (v_364 ^ v_43) ;
	assign v_366 = (v_361 ^ v_42) ;
	assign v_365 = (v_358 ^ v_41) ;
	assign v_343 = (v_340 ^ v_38) ;
	assign v_342 = (v_337 ^ v_37) ;
	assign v_341 = (v_334 ^ v_36) ;
	assign v_323 = (v_320 ^ v_35) ;
	assign v_322 = (v_317 ^ v_34) ;
	assign v_321 = (v_314 ^ v_33) ;
	assign v_299 = (v_296 ^ v_30) ;
	assign v_298 = (v_293 ^ v_29) ;
	assign v_297 = (v_290 ^ v_28) ;
	assign v_279 = (v_276 ^ v_27) ;
	assign v_278 = (v_273 ^ v_26) ;
	assign v_277 = (v_270 ^ v_25) ;
	assign v_255 = (v_252 ^ v_22) ;
	assign v_254 = (v_249 ^ v_21) ;
	assign v_253 = (v_246 ^ v_20) ;
	assign v_235 = (v_232 ^ v_19) ;
	assign v_234 = (v_229 ^ v_18) ;
	assign v_233 = (v_226 ^ v_17) ;
	assign v_211 = (v_208 ^ v_14) ;
	assign v_210 = (v_205 ^ v_13) ;
	assign v_209 = (v_202 ^ v_12) ;
	assign v_191 = (v_188 ^ v_11) ;
	assign v_190 = (v_185 ^ v_10) ;
	assign v_189 = (v_182 ^ v_9) ;
	assign v_1119 = ((~v_1116 & ~v_1117) & ~v_1118) ;
	assign v_1115 = ((~v_1112 & ~v_1113) & ~v_1114) ;
	assign v_1121 = (v_168 ^ v_88) ;
	assign v_1120 = (v_167 ^ v_87) ;
	assign v_1108 = ((~v_1105 & ~v_1106) & ~v_1107) ;
	assign v_1104 = ((~v_1101 & ~v_1102) & ~v_1103) ;
	assign v_1110 = (v_160 ^ v_88) ;
	assign v_1109 = (v_159 ^ v_87) ;
	assign v_1097 = ((~v_1094 & ~v_1095) & ~v_1096) ;
	assign v_1093 = ((~v_1090 & ~v_1091) & ~v_1092) ;
	assign v_1099 = (v_152 ^ v_88) ;
	assign v_1098 = (v_151 ^ v_87) ;
	assign v_1086 = ((~v_1083 & ~v_1084) & ~v_1085) ;
	assign v_1082 = ((~v_1079 & ~v_1080) & ~v_1081) ;
	assign v_1088 = (v_144 ^ v_88) ;
	assign v_1087 = (v_143 ^ v_87) ;
	assign v_1075 = ((~v_1072 & ~v_1073) & ~v_1074) ;
	assign v_1071 = ((~v_1068 & ~v_1069) & ~v_1070) ;
	assign v_1077 = (v_136 ^ v_88) ;
	assign v_1076 = (v_135 ^ v_87) ;
	assign v_1064 = ((~v_1061 & ~v_1062) & ~v_1063) ;
	assign v_1060 = ((~v_1057 & ~v_1058) & ~v_1059) ;
	assign v_1066 = (v_128 ^ v_88) ;
	assign v_1065 = (v_127 ^ v_87) ;
	assign v_1053 = ((~v_1050 & ~v_1051) & ~v_1052) ;
	assign v_1049 = ((~v_1046 & ~v_1047) & ~v_1048) ;
	assign v_1055 = (v_120 ^ v_88) ;
	assign v_1054 = (v_119 ^ v_87) ;
	assign v_1042 = ((~v_1039 & ~v_1040) & ~v_1041) ;
	assign v_1038 = ((~v_1035 & ~v_1036) & ~v_1037) ;
	assign v_1044 = (v_112 ^ v_88) ;
	assign v_1043 = (v_111 ^ v_87) ;
	assign v_1031 = ((~v_1028 & ~v_1029) & ~v_1030) ;
	assign v_1027 = ((~v_1024 & ~v_1025) & ~v_1026) ;
	assign v_1033 = (v_104 ^ v_88) ;
	assign v_1032 = (v_103 ^ v_87) ;
	assign v_1020 = ((~v_1017 & ~v_1018) & ~v_1019) ;
	assign v_1016 = ((~v_1013 & ~v_1014) & ~v_1015) ;
	assign v_1022 = (v_96 ^ v_88) ;
	assign v_1021 = (v_95 ^ v_87) ;
	assign v_1008 = ((~v_1005 & ~v_1006) & ~v_1007) ;
	assign v_988 = ((~v_985 & ~v_986) & ~v_987) ;
	assign v_1010 = (v_159 ^ v_168) ;
	assign v_1009 = (~v_167 ^ v_160) ;
	assign v_964 = ((~v_961 & ~v_962) & ~v_963) ;
	assign v_944 = ((~v_941 & ~v_942) & ~v_943) ;
	assign v_966 = (v_151 ^ v_160) ;
	assign v_965 = (~v_159 ^ v_152) ;
	assign v_920 = ((~v_917 & ~v_918) & ~v_919) ;
	assign v_900 = ((~v_897 & ~v_898) & ~v_899) ;
	assign v_922 = (v_143 ^ v_152) ;
	assign v_921 = (~v_151 ^ v_144) ;
	assign v_876 = ((~v_873 & ~v_874) & ~v_875) ;
	assign v_856 = ((~v_853 & ~v_854) & ~v_855) ;
	assign v_878 = (v_135 ^ v_144) ;
	assign v_877 = (~v_143 ^ v_136) ;
	assign v_832 = ((~v_829 & ~v_830) & ~v_831) ;
	assign v_812 = ((~v_809 & ~v_810) & ~v_811) ;
	assign v_834 = (v_127 ^ v_136) ;
	assign v_833 = (~v_135 ^ v_128) ;
	assign v_788 = ((~v_785 & ~v_786) & ~v_787) ;
	assign v_768 = ((~v_765 & ~v_766) & ~v_767) ;
	assign v_790 = (v_119 ^ v_128) ;
	assign v_789 = (~v_127 ^ v_120) ;
	assign v_744 = ((~v_741 & ~v_742) & ~v_743) ;
	assign v_724 = ((~v_721 & ~v_722) & ~v_723) ;
	assign v_746 = (v_111 ^ v_120) ;
	assign v_745 = (~v_119 ^ v_112) ;
	assign v_700 = ((~v_697 & ~v_698) & ~v_699) ;
	assign v_680 = ((~v_677 & ~v_678) & ~v_679) ;
	assign v_702 = (v_103 ^ v_112) ;
	assign v_701 = (~v_111 ^ v_104) ;
	assign v_656 = ((~v_653 & ~v_654) & ~v_655) ;
	assign v_636 = ((~v_633 & ~v_634) & ~v_635) ;
	assign v_658 = (v_95 ^ v_104) ;
	assign v_657 = (~v_103 ^ v_96) ;
	assign v_614 = ((~v_92 & ~v_93) & ~v_94) ;
	assign v_613 = ((~v_89 & ~v_90) & ~v_91) ;
	assign v_608 = ((~v_605 & ~v_606) & ~v_607) ;
	assign v_588 = ((~v_585 & ~v_586) & ~v_587) ;
	assign v_610 = (v_79 ^ v_88) ;
	assign v_609 = (~v_87 ^ v_80) ;
	assign v_564 = ((~v_561 & ~v_562) & ~v_563) ;
	assign v_544 = ((~v_541 & ~v_542) & ~v_543) ;
	assign v_566 = (v_71 ^ v_80) ;
	assign v_565 = (~v_79 ^ v_72) ;
	assign v_520 = ((~v_517 & ~v_518) & ~v_519) ;
	assign v_500 = ((~v_497 & ~v_498) & ~v_499) ;
	assign v_522 = (v_63 ^ v_72) ;
	assign v_521 = (~v_71 ^ v_64) ;
	assign v_476 = ((~v_473 & ~v_474) & ~v_475) ;
	assign v_456 = ((~v_453 & ~v_454) & ~v_455) ;
	assign v_478 = (v_55 ^ v_64) ;
	assign v_477 = (~v_63 ^ v_56) ;
	assign v_432 = ((~v_429 & ~v_430) & ~v_431) ;
	assign v_412 = ((~v_409 & ~v_410) & ~v_411) ;
	assign v_434 = (v_47 ^ v_56) ;
	assign v_433 = (~v_55 ^ v_48) ;
	assign v_388 = ((~v_385 & ~v_386) & ~v_387) ;
	assign v_368 = ((~v_365 & ~v_366) & ~v_367) ;
	assign v_390 = (v_39 ^ v_48) ;
	assign v_389 = (~v_47 ^ v_40) ;
	assign v_344 = ((~v_341 & ~v_342) & ~v_343) ;
	assign v_324 = ((~v_321 & ~v_322) & ~v_323) ;
	assign v_346 = (v_31 ^ v_40) ;
	assign v_345 = (~v_39 ^ v_32) ;
	assign v_300 = ((~v_297 & ~v_298) & ~v_299) ;
	assign v_280 = ((~v_277 & ~v_278) & ~v_279) ;
	assign v_302 = (v_23 ^ v_32) ;
	assign v_301 = (~v_31 ^ v_24) ;
	assign v_256 = ((~v_253 & ~v_254) & ~v_255) ;
	assign v_236 = ((~v_233 & ~v_234) & ~v_235) ;
	assign v_258 = (v_15 ^ v_24) ;
	assign v_257 = (~v_23 ^ v_16) ;
	assign v_212 = ((~v_209 & ~v_210) & ~v_211) ;
	assign v_192 = ((~v_189 & ~v_190) & ~v_191) ;
	assign v_214 = (v_7 ^ v_16) ;
	assign v_213 = (~v_15 ^ v_8) ;
	assign v_170 = ((~v_4 & ~v_5) & ~v_6) ;
	assign v_169 = ((~v_1 & ~v_2) & ~v_3) ;
	assign v_1122 = (((~v_1120 & ~v_1121) & v_1115) & v_1119) ;
	assign v_1111 = (((~v_1109 & ~v_1110) & v_1104) & v_1108) ;
	assign v_1100 = (((~v_1098 & ~v_1099) & v_1093) & v_1097) ;
	assign v_1089 = (((~v_1087 & ~v_1088) & v_1082) & v_1086) ;
	assign v_1078 = (((~v_1076 & ~v_1077) & v_1071) & v_1075) ;
	assign v_1067 = (((~v_1065 & ~v_1066) & v_1060) & v_1064) ;
	assign v_1056 = (((~v_1054 & ~v_1055) & v_1049) & v_1053) ;
	assign v_1045 = (((~v_1043 & ~v_1044) & v_1038) & v_1042) ;
	assign v_1034 = (((~v_1032 & ~v_1033) & v_1027) & v_1031) ;
	assign v_1023 = (((~v_1021 & ~v_1022) & v_1016) & v_1020) ;
	assign v_1011 = (((~v_1009 & ~v_1010) & v_988) & v_1008) ;
	assign v_967 = (((~v_965 & ~v_966) & v_944) & v_964) ;
	assign v_923 = (((~v_921 & ~v_922) & v_900) & v_920) ;
	assign v_879 = (((~v_877 & ~v_878) & v_856) & v_876) ;
	assign v_835 = (((~v_833 & ~v_834) & v_812) & v_832) ;
	assign v_791 = (((~v_789 & ~v_790) & v_768) & v_788) ;
	assign v_747 = (((~v_745 & ~v_746) & v_724) & v_744) ;
	assign v_703 = (((~v_701 & ~v_702) & v_680) & v_700) ;
	assign v_659 = (((~v_657 & ~v_658) & v_636) & v_656) ;
	assign v_615 = (((~v_95 & ~v_96) & v_613) & v_614) ;
	assign v_611 = (((~v_609 & ~v_610) & v_588) & v_608) ;
	assign v_567 = (((~v_565 & ~v_566) & v_544) & v_564) ;
	assign v_523 = (((~v_521 & ~v_522) & v_500) & v_520) ;
	assign v_479 = (((~v_477 & ~v_478) & v_456) & v_476) ;
	assign v_435 = (((~v_433 & ~v_434) & v_412) & v_432) ;
	assign v_391 = (((~v_389 & ~v_390) & v_368) & v_388) ;
	assign v_347 = (((~v_345 & ~v_346) & v_324) & v_344) ;
	assign v_303 = (((~v_301 & ~v_302) & v_280) & v_300) ;
	assign v_259 = (((~v_257 & ~v_258) & v_236) & v_256) ;
	assign v_215 = (((~v_213 & ~v_214) & v_192) & v_212) ;
	assign v_171 = (((~v_7 & ~v_8) & v_169) & v_170) ;
	assign v_1131 = ((((v_1078 | v_1089) | v_1100) | v_1111) | v_1122) ;
	assign v_1130 = ((((v_1023 | v_1034) | v_1045) | v_1056) | v_1067) ;
	assign v_1129 = ((((v_835 & v_879) & v_923) & v_967) & v_1011) ;
	assign v_1128 = ((((v_615 & v_659) & v_703) & v_747) & v_791) ;
	assign v_1127 = v_611 ;
	assign v_1126 = ((((v_391 & v_435) & v_479) & v_523) & v_567) ;
	assign v_1125 = ((((v_171 & v_215) & v_259) & v_303) & v_347) ;
	assign v_1123 = (v_1130 | v_1131) ;
	assign v_1012 = (v_1128 & v_1129) ;
	assign v_612 = ((v_1125 & v_1126) & v_1127) ;
	assign v_1124 = (v_1012 & v_1123) ;
	assign v_994 = (v_158 & v_992) ;
	assign v_974 = (v_155 & v_972) ;
	assign v_950 = (v_150 & v_948) ;
	assign v_930 = (v_147 & v_928) ;
	assign v_906 = (v_142 & v_904) ;
	assign v_886 = (v_139 & v_884) ;
	assign v_862 = (v_134 & v_860) ;
	assign v_842 = (v_131 & v_840) ;
	assign v_818 = (v_126 & v_816) ;
	assign v_798 = (v_123 & v_796) ;
	assign v_774 = (v_118 & v_772) ;
	assign v_754 = (v_115 & v_752) ;
	assign v_730 = (v_110 & v_728) ;
	assign v_710 = (v_107 & v_708) ;
	assign v_686 = (v_102 & v_684) ;
	assign v_666 = (v_99 & v_664) ;
	assign v_642 = (v_94 & v_640) ;
	assign v_622 = (v_91 & v_620) ;
	assign v_594 = (v_78 & v_592) ;
	assign v_574 = (v_75 & v_572) ;
	assign v_550 = (v_70 & v_548) ;
	assign v_530 = (v_67 & v_528) ;
	assign v_506 = (v_62 & v_504) ;
	assign v_486 = (v_59 & v_484) ;
	assign v_462 = (v_54 & v_460) ;
	assign v_442 = (v_51 & v_440) ;
	assign v_418 = (v_46 & v_416) ;
	assign v_398 = (v_43 & v_396) ;
	assign v_374 = (v_38 & v_372) ;
	assign v_354 = (v_35 & v_352) ;
	assign v_330 = (v_30 & v_328) ;
	assign v_310 = (v_27 & v_308) ;
	assign v_286 = (v_22 & v_284) ;
	assign v_266 = (v_19 & v_264) ;
	assign v_242 = (v_14 & v_240) ;
	assign v_222 = (v_11 & v_220) ;
	assign v_198 = (v_6 & v_196) ;
	assign v_178 = (v_3 & v_176) ;
	assign x_1 = (v_1124 | ~v_612) ;
	assign v_995 = v_994 ;
	assign v_975 = v_974 ;
	assign v_951 = v_950 ;
	assign v_931 = v_930 ;
	assign v_907 = v_906 ;
	assign v_887 = v_886 ;
	assign v_863 = v_862 ;
	assign v_843 = v_842 ;
	assign v_819 = v_818 ;
	assign v_799 = v_798 ;
	assign v_775 = v_774 ;
	assign v_755 = v_754 ;
	assign v_731 = v_730 ;
	assign v_711 = v_710 ;
	assign v_687 = v_686 ;
	assign v_667 = v_666 ;
	assign v_643 = v_642 ;
	assign v_623 = v_622 ;
	assign v_595 = v_594 ;
	assign v_575 = v_574 ;
	assign v_551 = v_550 ;
	assign v_531 = v_530 ;
	assign v_507 = v_506 ;
	assign v_487 = v_486 ;
	assign v_463 = v_462 ;
	assign v_443 = v_442 ;
	assign v_419 = v_418 ;
	assign v_399 = v_398 ;
	assign v_375 = v_374 ;
	assign v_355 = v_354 ;
	assign v_331 = v_330 ;
	assign v_311 = v_310 ;
	assign v_287 = v_286 ;
	assign v_267 = v_266 ;
	assign v_243 = v_242 ;
	assign v_223 = v_222 ;
	assign v_199 = v_198 ;
	assign v_179 = v_178 ;
	assign o_1 = x_1 ;
endmodule
