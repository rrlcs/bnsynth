module formula(i_0,i_1,i_2,i_3,i_4,i_5,i_6, i_7,i_8,i_9,i_10,i_11,i_12,i_13,i_14,i_15, out);
	input i_0 ,i_1 ,i_2 ,i_3,i_4,i_5,i_6, i_7,i_8,i_9,i_10,i_11,i_12,i_13,i_14,i_15;
	output out;
	assign out = ((((((((((((((((i_0 ^ i_1) ^ i_2) ^ i_3) ^ i_4) ^ i_5) ^ i_6) ^ i_7) ^ i_8) ^ i_9) ^ i_10) ^ i_11) ^ i_12) ^ i_13) ^ i_14) ^ i_15)) & (~i_0 | i_15) & (~i_1 | i_14) & (~i_2 | i_13) & (~i_3 | i_12);
endmodule
