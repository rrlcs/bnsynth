// Benchmark "SKOLEMFORMULA" written by ABC on Mon May 16 20:30:33 2022

module SKOLEMFORMULA ( 
    i0,
    i1  );
  input  i0;
  output i1;
  assign i1 = 1'b1;
endmodule


