module dec (count[0] , count[1] , count[2] , count[3] , count[4] , count[5] ,count[6] , count[7] , i1[0] , i1[1] , i1[2] , i1[3] , i1[4] , i1[5] , i1[6] , i1[7] , i1[8] , i1[9] , i1[10] , i1[11] , i1[12] , i1[13] , i1[14] , i1[15] , i1[16] , i1[17] , i1[18] , i1[19] , i1[20] , i1[21] , i1[22] , i1[23] , i1[24] , i1[25] , i1[26] , i1[27] , i1[28] , i1[29] , i1[30] , i1[31] , i1[32] , i1[33] , i1[34] , i1[35] , i1[36] , i1[37] , i1[38] , i1[39] , i1[40] , i1[41] , i1[42] , i1[43] , i1[44] , i1[45] , i1[46] , i1[47] , i1[48] , i1[49] , i1[50] , i1[51] , i1[52] , i1[53] , i1[54] , i1[55] , i1[56] , i1[57] , i1[58] , i1[59] , i1[60] , i1[61] , i1[62] , i1[63] , i1[64] , i1[65] , i1[66] , i1[67] , i1[68] , i1[69] , i1[70] , i1[71] , i1[72] , i1[73] , i1[74] , i1[75] , i1[76] , i1[77] , i1[78] , i1[79] , i1[80] , i1[81] , i1[82] , i1[83] , i1[84] , i1[85] , i1[86] , i1[87] , i1[88] , i1[89] , i1[90] , i1[91] , i1[92] , i1[93] , i1[94] , i1[95] , i1[96] , i1[97] , i1[98] , i1[99] , i1[100] , i1[101] , i1[102] , i1[103] , i1[104] , i1[105] , i1[106] , i1[107] , i1[108] , i1[109] , i1[110] , i1[111] , i1[112] , i1[113] , i1[114] , i1[115] , i1[116] , i1[117] , i1[118] , i1[119] , i1[120] , i1[121] , i1[122] , i1[123] , i1[124] , i1[125] , i1[126] , i1[127] , i2[0] , i2[1] , i2[2] , i2[3] , i2[4] , i2[5] , i2[6] , i2[7] , i2[8] , i2[9] , i2[10] , i2[11] , i2[12] , i2[13] , i2[14] , i2[15] , i2[16] , i2[17] , i2[18] , i2[19] , i2[20] , i2[21] , i2[22] , i2[23] , i2[24] , i2[25] , i2[26] , i2[27] , i2[28] , i2[29] , i2[30] , i2[31] , i2[32] , i2[33] , i2[34] , i2[35] , i2[36] , i2[37] , i2[38] , i2[39] , i2[40] , i2[41] , i2[42] , i2[43] , i2[44] , i2[45] , i2[46] , i2[47] , i2[48] , i2[49] , i2[50] , i2[51] , i2[52] , i2[53] , i2[54] , i2[55] , i2[56] , i2[57] , i2[58] , i2[59] , i2[60] , i2[61] , i2[62] , i2[63] , i2[64] , i2[65] , i2[66] , i2[67] , i2[68] , i2[69] , i2[70] , i2[71] , i2[72] , i2[73] , i2[74] , i2[75] , i2[76] , i2[77] , i2[78] , i2[79] , i2[80] , i2[81] , i2[82] , i2[83] , i2[84] , i2[85] , i2[86] , i2[87] , i2[88] , i2[89] , i2[90] , i2[91] , i2[92] , i2[93] , i2[94] , i2[95] , i2[96] , i2[97] , i2[98] , i2[99] , i2[100] , i2[101] , i2[102] , i2[103] , i2[104] , i2[105] , i2[106] , i2[107] , i2[108] , i2[109] , i2[110] , i2[111] , i2[112] , i2[113] , i2[114] , i2[115] , i2[116] , i2[117] , i2[118] , i2[119] , i2[120] , i2[121] , i2[122] , i2[123] , i2[124] , i2[125] , i2[126] , i2[127]);
  input  count[0] , count[1] , count[2] , count[3] , count[4] , count[5] , count[6] , count[7], i1[0] , i1[1] , i1[2] , i1[3] , i1[4] , i1[5] , i1[6] , i1[7] , i1[8] , i1[9] , i1[10] , i1[11] , i1[12] , i1[13] , i1[14] , i1[15] , i1[16] , i1[17] , i1[18] , i1[19] , i1[20] , i1[21] , i1[22] , i1[23] , i1[24] , i1[25] , i1[26] , i1[27] , i1[28] , i1[29] , i1[30] , i1[31] , i1[32] , i1[33] , i1[34] , i1[35] , i1[36] , i1[37] , i1[38] , i1[39] , i1[40] , i1[41] , i1[42] , i1[43] , i1[44] , i1[45] , i1[46] , i1[47] , i1[48] , i1[49] , i1[50] , i1[51] , i1[52] , i1[53] , i1[54] , i1[55] , i1[56] , i1[57] , i1[58] , i1[59] , i1[60] , i1[61] , i1[62] , i1[63] , i1[64] , i1[65] , i1[66] , i1[67] , i1[68] , i1[69] , i1[70] , i1[71] , i1[72] , i1[73] , i1[74] , i1[75] , i1[76] , i1[77] , i1[78] , i1[79] , i1[80] , i1[81] , i1[82] , i1[83] , i1[84] , i1[85] , i1[86] , i1[87] , i1[88] , i1[89] , i1[90] , i1[91] , i1[92] , i1[93] , i1[94] , i1[95] , i1[96] , i1[97] , i1[98] , i1[99] , i1[100] , i1[101] , i1[102] , i1[103] , i1[104] , i1[105] , i1[106] , i1[107] , i1[108] , i1[109] , i1[110] , i1[111] , i1[112] , i1[113] , i1[114] , i1[115] , i1[116] , i1[117] , i1[118] , i1[119] , i1[120] , i1[121] , i1[122] , i1[123] , i1[124] , i1[125] , i1[126] , i1[127] , i2[0] , i2[1] , i2[2] , i2[3] , i2[4] , i2[5] , i2[6] , i2[7] , i2[8] , i2[9] , i2[10] , i2[11] , i2[12] , i2[13] , i2[14] , i2[15] , i2[16] , i2[17] , i2[18] , i2[19] , i2[20] , i2[21] , i2[22] , i2[23] , i2[24] , i2[25] , i2[26] , i2[27] , i2[28] , i2[29] , i2[30] , i2[31] , i2[32] , i2[33] , i2[34] , i2[35] , i2[36] , i2[37] , i2[38] , i2[39] , i2[40] , i2[41] , i2[42] , i2[43] , i2[44] , i2[45] , i2[46] , i2[47] , i2[48] , i2[49] , i2[50] , i2[51] , i2[52] , i2[53] , i2[54] , i2[55] , i2[56] , i2[57] , i2[58] , i2[59] , i2[60] , i2[61] , i2[62] , i2[63] , i2[64] , i2[65] , i2[66] , i2[67] , i2[68] , i2[69] , i2[70] , i2[71] , i2[72] , i2[73] , i2[74] , i2[75] , i2[76] , i2[77] , i2[78] , i2[79] , i2[80] , i2[81] , i2[82] , i2[83] , i2[84] , i2[85] , i2[86] , i2[87] , i2[88] , i2[89] , i2[90] , i2[91] , i2[92] , i2[93] , i2[94] , i2[95] , i2[96] , i2[97] , i2[98] , i2[99] , i2[100] , i2[101] , i2[102] , i2[103] , i2[104] , i2[105] , i2[106] , i2[107] , i2[108] , i2[109] , i2[110] , i2[111] , i2[112] , i2[113] , i2[114] , i2[115] , i2[116] , i2[117] , i2[118] , i2[119] , i2[120] , i2[121] , i2[122] , i2[123] , i2[124] , i2[125] , i2[126] , i2[127] ;
  output out;
  wire n265, n266, n267, n268, n269, n270, n272, n273, n275, n276, n278,
    n280, n281, n283, n284, n286, n288, n290, n291, n293, n295, n296, n298,
    n300, n302, n304, n306, n308, n309, n326, n327, n344, n345, n362, n363,
    n380, n397, n414, n431, n432, n449, n466, n483, n500, n501, n518, n535,
    n552, selectp1[0] , selectp1[1] , selectp1[2] , selectp1[3] ,
    selectp1[4] , selectp1[5] , selectp1[6] , selectp1[7] ,
    selectp1[8] , selectp1[9] , selectp1[10] , selectp1[11] ,
    selectp1[12] , selectp1[13] , selectp1[14] , selectp1[15] ,
    selectp1[16] , selectp1[17] , selectp1[18] , selectp1[19] ,
    selectp1[20] , selectp1[21] , selectp1[22] , selectp1[23] ,
    selectp1[24] , selectp1[25] , selectp1[26] , selectp1[27] ,
    selectp1[28] , selectp1[29] , selectp1[30] , selectp1[31] ,
    selectp1[32] , selectp1[33] , selectp1[34] , selectp1[35] ,
    selectp1[36] , selectp1[37] , selectp1[38] , selectp1[39] ,
    selectp1[40] , selectp1[41] , selectp1[42] , selectp1[43] ,
    selectp1[44] , selectp1[45] , selectp1[46] , selectp1[47] ,
    selectp1[48] , selectp1[49] , selectp1[50] , selectp1[51] ,
    selectp1[52] , selectp1[53] , selectp1[54] , selectp1[55] ,
    selectp1[56] , selectp1[57] , selectp1[58] , selectp1[59] ,
    selectp1[60] , selectp1[61] , selectp1[62] , selectp1[63] ,
    selectp1[64] , selectp1[65] , selectp1[66] , selectp1[67] ,
    selectp1[68] , selectp1[69] , selectp1[70] , selectp1[71] ,
    selectp1[72] , selectp1[73] , selectp1[74] , selectp1[75] ,
    selectp1[76] , selectp1[77] , selectp1[78] , selectp1[79] ,
    selectp1[80] , selectp1[81] , selectp1[82] , selectp1[83] ,
    selectp1[84] , selectp1[85] , selectp1[86] , selectp1[87] ,
    selectp1[88] , selectp1[89] , selectp1[90] , selectp1[91] ,
    selectp1[92] , selectp1[93] , selectp1[94] , selectp1[95] ,
    selectp1[96] , selectp1[97] , selectp1[98] , selectp1[99] ,
    selectp1[100] , selectp1[101] , selectp1[102] , selectp1[103] ,
    selectp1[104] , selectp1[105] , selectp1[106] , selectp1[107] ,
    selectp1[108] , selectp1[109] , selectp1[110] , selectp1[111] ,
    selectp1[112] , selectp1[113] , selectp1[114] , selectp1[115] ,
    selectp1[116] , selectp1[117] , selectp1[118] , selectp1[119] ,
    selectp1[120] , selectp1[121] , selectp1[122] , selectp1[123] ,
    selectp1[124] , selectp1[125] , selectp1[126] , selectp1[127] ,
    selectp2[0] , selectp2[1] , selectp2[2] , selectp2[3] ,
    selectp2[4] , selectp2[5] , selectp2[6] , selectp2[7] ,
    selectp2[8] , selectp2[9] , selectp2[10] , selectp2[11] ,
    selectp2[12] , selectp2[13] , selectp2[14] , selectp2[15] ,
    selectp2[16] , selectp2[17] , selectp2[18] , selectp2[19] ,
    selectp2[20] , selectp2[21] , selectp2[22] , selectp2[23] ,
    selectp2[24] , selectp2[25] , selectp2[26] , selectp2[27] ,
    selectp2[28] , selectp2[29] , selectp2[30] , selectp2[31] ,
    selectp2[32] , selectp2[33] , selectp2[34] , selectp2[35] ,
    selectp2[36] , selectp2[37] , selectp2[38] , selectp2[39] ,
    selectp2[40] , selectp2[41] , selectp2[42] , selectp2[43] ,
    selectp2[44] , selectp2[45] , selectp2[46] , selectp2[47] ,
    selectp2[48] , selectp2[49] , selectp2[50] , selectp2[51] ,
    selectp2[52] , selectp2[53] , selectp2[54] , selectp2[55] ,
    selectp2[56] , selectp2[57] , selectp2[58] , selectp2[59] ,
    selectp2[60] , selectp2[61] , selectp2[62] , selectp2[63] ,
    selectp2[64] , selectp2[65] , selectp2[66] , selectp2[67] ,
    selectp2[68] , selectp2[69] , selectp2[70] , selectp2[71] ,
    selectp2[72] , selectp2[73] , selectp2[74] , selectp2[75] ,
    selectp2[76] , selectp2[77] , selectp2[78] , selectp2[79] ,
    selectp2[80] , selectp2[81] , selectp2[82] , selectp2[83] ,
    selectp2[84] , selectp2[85] , selectp2[86] , selectp2[87] ,
    selectp2[88] , selectp2[89] , selectp2[90] , selectp2[91] ,
    selectp2[92] , selectp2[93] , selectp2[94] , selectp2[95] ,
    selectp2[96] , selectp2[97] , selectp2[98] , selectp2[99] ,
    selectp2[100] , selectp2[101] , selectp2[102] , selectp2[103] ,
    selectp2[104] , selectp2[105] , selectp2[106] , selectp2[107] ,
    selectp2[108] , selectp2[109] , selectp2[110] , selectp2[111] ,
    selectp2[112] , selectp2[113] , selectp2[114] , selectp2[115] ,
    selectp2[116] , selectp2[117] , selectp2[118] , selectp2[119] ,
    selectp2[120] , selectp2[121] , selectp2[122] , selectp2[123] ,
    selectp2[124] , selectp2[125] , selectp2[126] , selectp2[127] , selectp1_1;
  assign n265 = ~count[4]  & ~count[5] ;
  assign n266 = ~count[6]  & count[7] ;
  assign n267 = n265 & n266;
  assign n268 = ~count[0]  & ~count[2] ;
  assign n269 = ~count[1]  & ~count[3] ;
  assign n270 = n268 & n269;
  assign selectp1[0]  = n267 & n270;
  assign n272 = count[0]  & ~count[2] ;
  assign n273 = n269 & n272;
  assign selectp1[1]  = n267 & n273;
  assign n275 = count[1]  & ~count[3] ;
  assign n276 = n268 & n275;
  assign selectp1[2]  = n267 & n276;
  assign n278 = n272 & n275;
  assign selectp1[3]  = n267 & n278;
  assign n280 = ~count[0]  & count[2] ;
  assign n281 = n269 & n280;
  assign selectp1[4]  = n267 & n281;
  assign n283 = count[0]  & count[2] ;
  assign n284 = n269 & n283;
  assign selectp1[5]  = n267 & n284;
  assign n286 = n275 & n280;
  assign selectp1[6]  = n267 & n286;
  assign n288 = n275 & n283;
  assign selectp1[7]  = n267 & n288;
  assign n290 = ~count[1]  & count[3] ;
  assign n291 = n268 & n290;
  assign selectp1[8]  = n267 & n291;
  assign n293 = n272 & n290;
  assign selectp1[9]  = n267 & n293;
  assign n295 = count[1]  & count[3] ;
  assign n296 = n268 & n295;
  assign selectp1[10]  = n267 & n296;
  assign n298 = n272 & n295;
  assign selectp1[11]  = n267 & n298;
  assign n300 = n280 & n290;
  assign selectp1[12]  = n267 & n300;
  assign n302 = n283 & n290;
  assign selectp1[13]  = n267 & n302;
  assign n304 = n280 & n295;
  assign selectp1[14]  = n267 & n304;
  assign n306 = n283 & n295;
  assign selectp1[15]  = n267 & n306;
  assign n308 = count[4]  & ~count[5] ;
  assign n309 = n266 & n308;
  assign selectp1[16]  = n270 & n309;
  assign selectp1[17]  = n273 & n309;
  assign selectp1[18]  = n276 & n309;
  assign selectp1[19]  = n278 & n309;
  assign selectp1[20]  = n281 & n309;
  assign selectp1[21]  = n284 & n309;
  assign selectp1[22]  = n286 & n309;
  assign selectp1[23]  = n288 & n309;
  assign selectp1[24]  = n291 & n309;
  assign selectp1[25]  = n293 & n309;
  assign selectp1[26]  = n296 & n309;
  assign selectp1[27]  = n298 & n309;
  assign selectp1[28]  = n300 & n309;
  assign selectp1[29]  = n302 & n309;
  assign selectp1[30]  = n304 & n309;
  assign selectp1[31]  = n306 & n309;
  assign n326 = ~count[4]  & count[5] ;
  assign n327 = n266 & n326;
  assign selectp1[32]  = n270 & n327;
  assign selectp1[33]  = n273 & n327;
  assign selectp1[34]  = n276 & n327;
  assign selectp1[35]  = n278 & n327;
  assign selectp1[36]  = n281 & n327;
  assign selectp1[37]  = n284 & n327;
  assign selectp1[38]  = n286 & n327;
  assign selectp1[39]  = n288 & n327;
  assign selectp1[40]  = n291 & n327;
  assign selectp1[41]  = n293 & n327;
  assign selectp1[42]  = n296 & n327;
  assign selectp1[43]  = n298 & n327;
  assign selectp1[44]  = n300 & n327;
  assign selectp1[45]  = n302 & n327;
  assign selectp1[46]  = n304 & n327;
  assign selectp1[47]  = n306 & n327;
  assign n344 = count[4]  & count[5] ;
  assign n345 = n266 & n344;
  assign selectp1[48]  = n270 & n345;
  assign selectp1[49]  = n273 & n345;
  assign selectp1[50]  = n276 & n345;
  assign selectp1[51]  = n278 & n345;
  assign selectp1[52]  = n281 & n345;
  assign selectp1[53]  = n284 & n345;
  assign selectp1[54]  = n286 & n345;
  assign selectp1[55]  = n288 & n345;
  assign selectp1[56]  = n291 & n345;
  assign selectp1[57]  = n293 & n345;
  assign selectp1[58]  = n296 & n345;
  assign selectp1[59]  = n298 & n345;
  assign selectp1[60]  = n300 & n345;
  assign selectp1[61]  = n302 & n345;
  assign selectp1[62]  = n304 & n345;
  assign selectp1[63]  = n306 & n345;
  assign n362 = count[6]  & count[7] ;
  assign n363 = n265 & n362;
  assign selectp1[64]  = n270 & n363;
  assign selectp1[65]  = n273 & n363;
  assign selectp1[66]  = n276 & n363;
  assign selectp1[67]  = n278 & n363;
  assign selectp1[68]  = n281 & n363;
  assign selectp1[69]  = n284 & n363;
  assign selectp1[70]  = n286 & n363;
  assign selectp1[71]  = n288 & n363;
  assign selectp1[72]  = n291 & n363;
  assign selectp1[73]  = n293 & n363;
  assign selectp1[74]  = n296 & n363;
  assign selectp1[75]  = n298 & n363;
  assign selectp1[76]  = n300 & n363;
  assign selectp1[77]  = n302 & n363;
  assign selectp1[78]  = n304 & n363;
  assign selectp1[79]  = n306 & n363;
  assign n380 = n308 & n362;
  assign selectp1[80]  = n270 & n380;
  assign selectp1[81]  = n273 & n380;
  assign selectp1[82]  = n276 & n380;
  assign selectp1[83]  = n278 & n380;
  assign selectp1[84]  = n281 & n380;
  assign selectp1[85]  = n284 & n380;
  assign selectp1[86]  = n286 & n380;
  assign selectp1[87]  = n288 & n380;
  assign selectp1[88]  = n291 & n380;
  assign selectp1[89]  = n293 & n380;
  assign selectp1[90]  = n296 & n380;
  assign selectp1[91]  = n298 & n380;
  assign selectp1[92]  = n300 & n380;
  assign selectp1[93]  = n302 & n380;
  assign selectp1[94]  = n304 & n380;
  assign selectp1[95]  = n306 & n380;
  assign n397 = n326 & n362;
  assign selectp1[96]  = n270 & n397;
  assign selectp1[97]  = n273 & n397;
  assign selectp1[98]  = n276 & n397;
  assign selectp1[99]  = n278 & n397;
  assign selectp1[100]  = n281 & n397;
  assign selectp1[101]  = n284 & n397;
  assign selectp1[102]  = n286 & n397;
  assign selectp1[103]  = n288 & n397;
  assign selectp1[104]  = n291 & n397;
  assign selectp1[105]  = n293 & n397;
  assign selectp1[106]  = n296 & n397;
  assign selectp1[107]  = n298 & n397;
  assign selectp1[108]  = n300 & n397;
  assign selectp1[109]  = n302 & n397;
  assign selectp1[110]  = n304 & n397;
  assign selectp1[111]  = n306 & n397;
  assign n414 = n344 & n362;
  assign selectp1[112]  = n270 & n414;
  assign selectp1[113]  = n273 & n414;
  assign selectp1[114]  = n276 & n414;
  assign selectp1[115]  = n278 & n414;
  assign selectp1[116]  = n281 & n414;
  assign selectp1[117]  = n284 & n414;
  assign selectp1[118]  = n286 & n414;
  assign selectp1[119]  = n288 & n414;
  assign selectp1[120]  = n291 & n414;
  assign selectp1[121]  = n293 & n414;
  assign selectp1[122]  = n296 & n414;
  assign selectp1[123]  = n298 & n414;
  assign selectp1[124]  = n300 & n414;
  assign selectp1[125]  = n302 & n414;
  assign selectp1[126]  = n304 & n414;
  assign selectp1[127]  = n306 & n414;
  assign n431 = ~count[6]  & ~count[7] ;
  assign n432 = n265 & n431;
  assign selectp2[0]  = n270 & n432;
  assign selectp2[1]  = n273 & n432;
  assign selectp2[2]  = n276 & n432;
  assign selectp2[3]  = n278 & n432;
  assign selectp2[4]  = n281 & n432;
  assign selectp2[5]  = n284 & n432;
  assign selectp2[6]  = n286 & n432;
  assign selectp2[7]  = n288 & n432;
  assign selectp2[8]  = n291 & n432;
  assign selectp2[9]  = n293 & n432;
  assign selectp2[10]  = n296 & n432;
  assign selectp2[11]  = n298 & n432;
  assign selectp2[12]  = n300 & n432;
  assign selectp2[13]  = n302 & n432;
  assign selectp2[14]  = n304 & n432;
  assign selectp2[15]  = n306 & n432;
  assign n449 = n308 & n431;
  assign selectp2[16]  = n270 & n449;
  assign selectp2[17]  = n273 & n449;
  assign selectp2[18]  = n276 & n449;
  assign selectp2[19]  = n278 & n449;
  assign selectp2[20]  = n281 & n449;
  assign selectp2[21]  = n284 & n449;
  assign selectp2[22]  = n286 & n449;
  assign selectp2[23]  = n288 & n449;
  assign selectp2[24]  = n291 & n449;
  assign selectp2[25]  = n293 & n449;
  assign selectp2[26]  = n296 & n449;
  assign selectp2[27]  = n298 & n449;
  assign selectp2[28]  = n300 & n449;
  assign selectp2[29]  = n302 & n449;
  assign selectp2[30]  = n304 & n449;
  assign selectp2[31]  = n306 & n449;
  assign n466 = n326 & n431;
  assign selectp2[32]  = n270 & n466;
  assign selectp2[33]  = n273 & n466;
  assign selectp2[34]  = n276 & n466;
  assign selectp2[35]  = n278 & n466;
  assign selectp2[36]  = n281 & n466;
  assign selectp2[37]  = n284 & n466;
  assign selectp2[38]  = n286 & n466;
  assign selectp2[39]  = n288 & n466;
  assign selectp2[40]  = n291 & n466;
  assign selectp2[41]  = n293 & n466;
  assign selectp2[42]  = n296 & n466;
  assign selectp2[43]  = n298 & n466;
  assign selectp2[44]  = n300 & n466;
  assign selectp2[45]  = n302 & n466;
  assign selectp2[46]  = n304 & n466;
  assign selectp2[47]  = n306 & n466;
  assign n483 = n344 & n431;
  assign selectp2[48]  = n270 & n483;
  assign selectp2[49]  = n273 & n483;
  assign selectp2[50]  = n276 & n483;
  assign selectp2[51]  = n278 & n483;
  assign selectp2[52]  = n281 & n483;
  assign selectp2[53]  = n284 & n483;
  assign selectp2[54]  = n286 & n483;
  assign selectp2[55]  = n288 & n483;
  assign selectp2[56]  = n291 & n483;
  assign selectp2[57]  = n293 & n483;
  assign selectp2[58]  = n296 & n483;
  assign selectp2[59]  = n298 & n483;
  assign selectp2[60]  = n300 & n483;
  assign selectp2[61]  = n302 & n483;
  assign selectp2[62]  = n304 & n483;
  assign selectp2[63]  = n306 & n483;
  assign n500 = count[6]  & ~count[7] ;
  assign n501 = n265 & n500;
  assign selectp2[64]  = n270 & n501;
  assign selectp2[65]  = n273 & n501;
  assign selectp2[66]  = n276 & n501;
  assign selectp2[67]  = n278 & n501;
  assign selectp2[68]  = n281 & n501;
  assign selectp2[69]  = n284 & n501;
  assign selectp2[70]  = n286 & n501;
  assign selectp2[71]  = n288 & n501;
  assign selectp2[72]  = n291 & n501;
  assign selectp2[73]  = n293 & n501;
  assign selectp2[74]  = n296 & n501;
  assign selectp2[75]  = n298 & n501;
  assign selectp2[76]  = n300 & n501;
  assign selectp2[77]  = n302 & n501;
  assign selectp2[78]  = n304 & n501;
  assign selectp2[79]  = n306 & n501;
  assign n518 = n308 & n500;
  assign selectp2[80]  = n270 & n518;
  assign selectp2[81]  = n273 & n518;
  assign selectp2[82]  = n276 & n518;
  assign selectp2[83]  = n278 & n518;
  assign selectp2[84]  = n281 & n518;
  assign selectp2[85]  = n284 & n518;
  assign selectp2[86]  = n286 & n518;
  assign selectp2[87]  = n288 & n518;
  assign selectp2[88]  = n291 & n518;
  assign selectp2[89]  = n293 & n518;
  assign selectp2[90]  = n296 & n518;
  assign selectp2[91]  = n298 & n518;
  assign selectp2[92]  = n300 & n518;
  assign selectp2[93]  = n302 & n518;
  assign selectp2[94]  = n304 & n518;
  assign selectp2[95]  = n306 & n518;
  assign n535 = n326 & n500;
  assign selectp2[96]  = n270 & n535;
  assign selectp2[97]  = n273 & n535;
  assign selectp2[98]  = n276 & n535;
  assign selectp2[99]  = n278 & n535;
  assign selectp2[100]  = n281 & n535;
  assign selectp2[101]  = n284 & n535;
  assign selectp2[102]  = n286 & n535;
  assign selectp2[103]  = n288 & n535;
  assign selectp2[104]  = n291 & n535;
  assign selectp2[105]  = n293 & n535;
  assign selectp2[106]  = n296 & n535;
  assign selectp2[107]  = n298 & n535;
  assign selectp2[108]  = n300 & n535;
  assign selectp2[109]  = n302 & n535;
  assign selectp2[110]  = n304 & n535;
  assign selectp2[111]  = n306 & n535;
  assign n552 = n344 & n500;
  assign selectp2[112]  = n270 & n552;
  assign selectp2[113]  = n273 & n552;
  assign selectp2[114]  = n276 & n552;
  assign selectp2[115]  = n278 & n552;
  assign selectp2[116]  = n281 & n552;
  assign selectp2[117]  = n284 & n552;
  assign selectp2[118]  = n286 & n552;
  assign selectp2[119]  = n288 & n552;
  assign selectp2[120]  = n291 & n552;
  assign selectp2[121]  = n293 & n552;
  assign selectp2[122]  = n296 & n552;
  assign selectp2[123]  = n298 & n552;
  assign selectp2[124]  = n300 & n552;
  assign selectp2[125]  = n302 & n552;
  assign selectp2[126]  = n304 & n552;
  assign selectp2[127]  = n306 & n552;

  assign selectp1_1 = i1[0];
  assign out = ~(selectp1[0] ^ selectp1_1);
endmodule

