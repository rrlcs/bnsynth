// skolem function for order file variables
// Generated using findDep.cpp 
module sortnetsort10.AE.stepl.004 (v_56, v_57, v_58, v_59, v_60, v_61, v_62, v_63, v_64, v_65, v_66, v_67, v_68, v_69, v_70, v_71, v_72, v_73, v_74, v_75, v_76, v_77, v_78, v_79, v_80, v_81, v_82, v_83, v_84, v_85, v_86, v_87, v_88, v_89, v_90, v_91, v_92, v_93, v_94, v_95, v_96, v_97, v_98, v_99, v_100, v_101, v_102, v_103, v_104, v_105, v_106, v_107, v_108, v_109, v_110, v_111, v_112, v_113, v_114, v_115, v_116, v_117, v_118, v_119, v_120, v_121, v_122, v_123, v_124, v_125, v_126, v_127, v_128, v_129, v_130, v_131, v_132, v_133, v_134, v_135, v_136, v_137, v_138, v_139, v_140, v_141, v_142, v_143, v_144, v_145, v_146, v_147, v_148, v_149, v_150, v_151, v_152, v_153, v_154, v_155, v_156, v_157, v_158, v_159, v_160, v_161, v_162, v_163, v_164, v_165, v_166, v_167, v_168, v_169, v_170, v_171, v_172, v_173, v_174, v_175, v_176, v_177, v_178, v_179, v_180, v_181, v_182, v_183, v_184, v_185, v_186, v_187, v_188, v_189, v_190, v_191, v_192, v_193, v_194, v_195, v_196, v_197, v_198, v_199, v_200, v_201, v_202, v_203, v_204, v_205, v_206, v_207, v_208, v_209, v_210, v_211, v_212, v_213, v_214, v_215, v_216, v_217, v_218, v_219, v_220, v_221, v_222, v_223, v_224, v_225, v_226, v_227, v_228, v_229, v_230, v_231, v_232, v_233, v_234, v_235, v_236, v_237, v_238, v_239, v_240, v_241, v_242, v_243, v_244, v_245, v_246, v_247, v_248, v_249, v_250, v_251, v_252, v_253, v_254, v_255, v_256, v_257, v_258, v_259, v_260, v_261, v_262, v_263, v_264, v_265, v_266, v_267, v_268, v_269, v_270, v_271, v_272, v_273, v_274, v_275, v_276, v_277, v_278, v_279, v_280, v_281, v_282, v_283, v_284, v_285, v_286, v_287, v_288, v_289, v_290, v_291, v_292, v_293, v_294, v_295, v_296, v_297, v_298, v_299, v_300, v_301, v_302, v_303, v_304, v_305, v_306, v_307, v_308, v_309, v_310, v_311, v_312, v_313, v_314, v_315, v_316, v_317, v_318, v_319, v_320, v_321, v_322, v_323, v_324, v_325, v_326, v_327, v_328, v_329, v_330, v_331, v_332, v_333, v_334, v_335, v_336, v_337, v_338, v_339, v_340, v_341, v_342, v_343, v_344, v_345, v_346, v_347, v_348, v_349, v_350, v_351, v_352, v_353, v_354, v_355, v_356, v_357, v_358, v_359, v_360, v_361, v_362, v_363, v_364, v_365, v_366, v_367, v_368, v_369, v_370, v_371, v_372, v_373, v_374, v_375, v_376, v_377, v_378, v_379, v_3400, v_3401, v_3402, v_3403, v_3404, v_3405, v_3406, v_3407, v_3408, v_3409, v_3410, v_3411, v_3412, v_3413, v_3414, v_3415, v_3416, v_3417, v_3418, v_3419, v_3420, v_3421, v_3422, v_3423, v_3424, v_3425, v_3426, v_3427, v_3428, v_3429, v_3430, v_3431, v_3432, v_3433, v_3434, v_3435, v_3436, v_3437, v_3438, v_3439, v_3440, v_3441, v_3442, v_3443, v_3444, v_3445, v_3446, v_3447, v_3448, v_3449, v_3450, v_3451, v_3452, v_3453, v_3454, v_3455, v_3456, v_3457, v_3458, v_3459, v_3460, v_3461, v_3462, v_3463, v_3464, v_3465, v_3466, v_3467, v_3468, v_3469, v_3470, v_3471, v_3472, v_3473, v_3474, v_3475, v_3476, v_3477, v_3478, v_3479, v_3480, v_3481, v_3482, v_3483, v_3484, v_3485, v_3486, v_3487, v_3488, v_3489, v_3490, v_3491, v_3492, v_3493, v_3494, v_3495, v_3496, v_3497, v_3498, v_3499, v_3500, v_3501, v_3502, v_3503, v_3504, v_3505, v_3506, v_3507, v_3508, v_3509, v_3510, v_3511, v_3512, v_3513, v_3514, v_3515, v_3516, v_3517, v_3518, v_3519, v_3520, v_3521, v_3522, v_3523, v_3524, v_3525, v_3526, v_3527, v_3528, v_3529, v_3530, v_3531, v_3532, v_3533, v_3534, v_3535, v_3536, v_3537, v_3538, v_3539, v_3540, v_3541, v_3542, v_3543, v_3634, v_3635, v_3636, v_3637, v_3638, v_3639, v_3640, v_3641, v_3642, v_3643, v_3644, v_3645, v_3646, v_3647, v_3648, v_3649, v_3650, v_3651, v_3652, v_3653, v_3654, v_3655, v_3656, v_3657, v_3658, v_3659, v_3660, v_3661, v_3662, v_3663, v_3664, v_3665, v_3666, v_3667, v_3668, v_3669, v_3670, v_3671, v_3672, v_3673, v_3674, v_3675, v_3676, v_3677, v_3678, v_3679, v_3680, v_3681, v_3682, v_3683, v_3684, v_3685, v_3686, v_3687, v_3688, v_3689, v_3690, v_3691, v_3692, v_3693, v_3694, v_3695, v_3696, v_3697, v_3698, v_3699, v_3700, v_3701, v_3702, v_3703, v_3704, v_3705, v_3706, v_3707, v_3708, v_3709, v_3710, v_3711, v_3712, v_3713, v_3714, v_3715, v_3716, v_3717, v_3718, v_3719, v_3720, v_3721, v_3722, v_3723, v_3724, v_3725, v_3726, v_3727, v_3728, v_3729, v_3730, v_3731, v_3732, v_3733, v_3734, v_3735, v_3736, v_3737, v_3738, v_3739, v_3740, v_3741, v_3742, v_3743, v_3744, v_3745, v_3746, v_3747, v_3748, v_3749, v_3750, v_3751, v_3752, v_3753, v_3754, v_3755, v_3756, v_3757, v_3758, v_3759, v_3760, v_3761, v_3762, v_3763, v_3764, v_3765, v_3766, v_3767, v_3768, v_3769, v_3770, v_3771, v_3772, v_3773, v_3774, v_3775, v_3776, v_3777, v_3868, v_3869, v_3870, v_3871, v_3872, v_3873, v_3874, v_3875, v_3876, v_3877, v_3878, v_3879, v_3880, v_3881, v_3882, v_3883, v_3884, v_3885, v_3886, v_3887, v_3888, v_3889, v_3890, v_3891, v_3892, v_3893, v_3894, v_3895, v_3896, v_3897, v_3898, v_3899, v_3900, v_3901, v_3902, v_3903, v_3904, v_3905, v_3906, v_3907, v_3908, v_3909, v_3910, v_3911, v_3912, v_3913, v_3914, v_3915, v_3916, v_3917, v_3918, v_3919, v_3920, v_3921, v_3922, v_3923, v_3924, v_3925, v_3926, v_3927, v_3928, v_3929, v_3930, v_3931, v_3932, v_3933, v_3934, v_3935, v_3936, v_3937, v_3938, v_3939, v_3940, v_3941, v_3942, v_3943, v_3944, v_3945, v_3946, v_3947, v_3948, v_3949, v_3950, v_3951, v_3952, v_3953, v_3954, v_3955, v_3956, v_3957, v_3958, v_3959, v_3960, v_3961, v_3962, v_3963, v_3964, v_3965, v_3966, v_3967, v_3968, v_3969, v_3970, v_3971, v_3972, v_3973, v_3974, v_3975, v_3976, v_3977, v_3978, v_3979, v_3980, v_3981, v_3982, v_3983, v_3984, v_3985, v_3986, v_3987, v_3988, v_3989, v_3990, v_3991, v_3992, v_3993, v_3994, v_3995, v_3996, v_3997, v_3998, v_3999, v_4000, v_4001, v_4002, v_4003, v_4004, v_4005, v_4006, v_4007, v_4008, v_4009, v_4010, v_4011, v_1, v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_12, v_13, v_14, v_15, v_16, v_17, v_18, v_19, v_20, v_21, v_22, v_23, v_24, v_25, v_26, v_27, v_28, v_29, v_30, v_31, v_32, v_33, v_34, v_35, v_36, v_37, v_38, v_39, v_40, v_41, v_42, v_43, v_44, v_45, v_46, v_47, v_48, v_49, v_50, v_51, v_52, v_53, v_54, v_55, v_380, v_381, v_382, v_383, v_384, v_385, v_386, v_387, v_388, v_389, v_390, v_391, v_392, v_393, v_394, v_395, v_396, v_397, v_398, v_399, v_400, v_401, v_402, v_403, v_404, v_405, v_406, v_407, v_408, v_409, v_410, v_411, v_412, v_413, v_414, v_415, v_416, v_417, v_418, v_419, v_420, v_421, v_422, v_423, v_424, v_425, v_426, v_427, v_428, v_429, v_430, v_431, v_432, v_433, v_434, v_435, v_436, v_437, v_438, v_439, v_440, v_441, v_442, v_443, v_444, v_445, v_446, v_447, v_448, v_449, v_450, v_451, v_452, v_453, v_454, v_455, v_456, v_457, v_458, v_459, v_460, v_461, v_462, v_463, v_464, v_465, v_466, v_467, v_468, v_469, v_470, v_471, v_472, v_473, v_474, v_475, v_476, v_477, v_478, v_479, v_480, v_481, v_482, v_483, v_484, v_485, v_486, v_487, v_488, v_489, v_490, v_491, v_492, v_493, v_494, v_495, v_496, v_497, v_498, v_499, v_500, v_501, v_502, v_503, v_504, v_505, v_506, v_507, v_508, v_509, v_510, v_511, v_512, v_513, v_514, v_515, v_516, v_517, v_518, v_519, v_520, v_521, v_522, v_523, v_524, v_525, v_526, v_527, v_528, v_529, v_530, v_531, v_532, v_533, v_534, v_535, v_536, v_537, v_538, v_539, v_540, v_541, v_542, v_543, v_544, v_545, v_546, v_547, v_548, v_549, v_550, v_551, v_552, v_553, v_554, v_555, v_556, v_557, v_558, v_559, v_560, v_561, v_562, v_563, v_564, v_565, v_566, v_567, v_568, v_569, v_570, v_571, v_572, v_573, v_574, v_575, v_576, v_577, v_578, v_579, v_580, v_581, v_582, v_583, v_584, v_585, v_586, v_587, v_588, v_589, v_590, v_591, v_592, v_593, v_594, v_595, v_596, v_597, v_598, v_599, v_600, v_601, v_602, v_603, v_604, v_605, v_606, v_607, v_608, v_609, v_610, v_611, v_612, v_613, v_614, v_615, v_616, v_617, v_618, v_619, v_620, v_621, v_622, v_623, v_624, v_625, v_626, v_627, v_628, v_629, v_630, v_631, v_632, v_633, v_634, v_635, v_636, v_637, v_638, v_639, v_640, v_641, v_642, v_643, v_644, v_645, v_646, v_647, v_648, v_649, v_650, v_651, v_652, v_653, v_654, v_655, v_656, v_657, v_658, v_659, v_705, v_706, v_707, v_708, v_709, v_710, v_711, v_712, v_713, v_714, v_715, v_716, v_717, v_718, v_719, v_720, v_721, v_722, v_723, v_724, v_725, v_726, v_727, v_728, v_729, v_730, v_731, v_732, v_733, v_734, v_735, v_736, v_737, v_738, v_739, v_740, v_741, v_742, v_743, v_744, v_745, v_746, v_747, v_748, v_749, v_750, v_751, v_752, v_753, v_754, v_755, v_756, v_757, v_758, v_759, v_760, v_761, v_762, v_763, v_764, v_765, v_766, v_767, v_768, v_769, v_770, v_771, v_772, v_773, v_774, v_775, v_776, v_777, v_778, v_779, v_780, v_781, v_782, v_783, v_784, v_785, v_786, v_787, v_788, v_789, v_790, v_791, v_792, v_793, v_794, v_795, v_796, v_797, v_798, v_799, v_800, v_801, v_802, v_803, v_804, v_805, v_806, v_807, v_808, v_809, v_810, v_811, v_812, v_813, v_814, v_815, v_816, v_817, v_818, v_819, v_820, v_821, v_822, v_823, v_824, v_825, v_826, v_827, v_828, v_829, v_830, v_831, v_832, v_833, v_834, v_835, v_836, v_837, v_838, v_839, v_840, v_841, v_842, v_843, v_844, v_845, v_846, v_847, v_848, v_849, v_850, v_851, v_852, v_853, v_854, v_855, v_856, v_857, v_858, v_859, v_860, v_861, v_862, v_863, v_864, v_865, v_866, v_867, v_868, v_869, v_870, v_871, v_872, v_873, v_874, v_875, v_876, v_877, v_878, v_879, v_880, v_881, v_882, v_883, v_884, v_885, v_931, v_932, v_933, v_934, v_935, v_936, v_937, v_938, v_939, v_940, v_941, v_942, v_943, v_944, v_945, v_946, v_947, v_948, v_949, v_950, v_951, v_952, v_953, v_954, v_955, v_956, v_957, v_958, v_959, v_960, v_961, v_962, v_963, v_964, v_965, v_966, v_967, v_968, v_969, v_970, v_971, v_972, v_973, v_974, v_975, v_976, v_977, v_978, v_979, v_980, v_981, v_982, v_983, v_984, v_985, v_986, v_987, v_988, v_989, v_990, v_991, v_992, v_993, v_994, v_995, v_996, v_997, v_998, v_999, v_1000, v_1001, v_1002, v_1003, v_1004, v_1005, v_1006, v_1007, v_1008, v_1009, v_1010, v_1011, v_1012, v_1013, v_1014, v_1015, v_1016, v_1017, v_1018, v_1019, v_1020, v_1021, v_1022, v_1023, v_1024, v_1025, v_1026, v_1027, v_1028, v_1029, v_1030, v_1031, v_1032, v_1033, v_1034, v_1035, v_1036, v_1037, v_1038, v_1039, v_1040, v_1041, v_1042, v_1043, v_1044, v_1045, v_1046, v_1047, v_1048, v_1049, v_1050, v_1051, v_1052, v_1053, v_1054, v_1055, v_1056, v_1057, v_1058, v_1059, v_1060, v_1061, v_1062, v_1063, v_1064, v_1065, v_1066, v_1067, v_1068, v_1069, v_1070, v_1071, v_1072, v_1073, v_1074, v_1075, v_1076, v_1077, v_1078, v_1079, v_1080, v_1081, v_1082, v_1083, v_1084, v_1085, v_1086, v_1087, v_1088, v_1089, v_1090, v_1091, v_1092, v_1093, v_1094, v_1095, v_1096, v_1097, v_1098, v_1099, v_1100, v_1101, v_1102, v_1103, v_1104, v_1105, v_1106, v_1107, v_1108, v_1109, v_1110, v_1111, v_1157, v_1158, v_1159, v_1160, v_1161, v_1162, v_1163, v_1164, v_1165, v_1166, v_1167, v_1168, v_1169, v_1170, v_1171, v_1172, v_1173, v_1174, v_1175, v_1176, v_1177, v_1178, v_1179, v_1180, v_1181, v_1182, v_1183, v_1184, v_1185, v_1186, v_1187, v_1188, v_1189, v_1190, v_1191, v_1192, v_1193, v_1194, v_1195, v_1196, v_1197, v_1198, v_1199, v_1200, v_1201, v_1202, v_1203, v_1204, v_1205, v_1206, v_1207, v_1208, v_1209, v_1210, v_1211, v_1212, v_1213, v_1214, v_1215, v_1216, v_1217, v_1218, v_1219, v_1220, v_1221, v_1222, v_1223, v_1224, v_1225, v_1226, v_1227, v_1228, v_1229, v_1230, v_1231, v_1232, v_1233, v_1234, v_1235, v_1236, v_1237, v_1238, v_1239, v_1240, v_1241, v_1242, v_1243, v_1244, v_1245, v_1246, v_1247, v_1248, v_1249, v_1250, v_1251, v_1252, v_1253, v_1254, v_1255, v_1256, v_1257, v_1258, v_1259, v_1260, v_1261, v_1262, v_1263, v_1264, v_1265, v_1266, v_1267, v_1268, v_1269, v_1270, v_1271, v_1272, v_1273, v_1274, v_1275, v_1276, v_1277, v_1278, v_1279, v_1280, v_1281, v_1282, v_1283, v_1284, v_1285, v_1286, v_1287, v_1288, v_1289, v_1290, v_1291, v_1292, v_1293, v_1294, v_1295, v_1296, v_1297, v_1298, v_1299, v_1300, v_1301, v_1302, v_1303, v_1304, v_1305, v_1306, v_1307, v_1308, v_1309, v_1310, v_1311, v_1312, v_1313, v_1314, v_1315, v_1316, v_1317, v_1318, v_1319, v_1320, v_1321, v_1322, v_1323, v_1324, v_1325, v_1326, v_1327, v_1328, v_1329, v_1330, v_1331, v_1332, v_1333, v_1334, v_1335, v_1336, v_1337, v_1383, v_1384, v_1385, v_1386, v_1387, v_1388, v_1389, v_1390, v_1391, v_1392, v_1393, v_1394, v_1395, v_1396, v_1397, v_1398, v_1399, v_1400, v_1401, v_1402, v_1403, v_1404, v_1405, v_1406, v_1407, v_1408, v_1409, v_1410, v_1411, v_1412, v_1413, v_1414, v_1415, v_1416, v_1417, v_1418, v_1419, v_1420, v_1421, v_1422, v_1423, v_1424, v_1425, v_1426, v_1427, v_1428, v_1429, v_1430, v_1431, v_1432, v_1433, v_1434, v_1435, v_1436, v_1437, v_1438, v_1439, v_1440, v_1441, v_1442, v_1443, v_1444, v_1445, v_1446, v_1447, v_1448, v_1449, v_1450, v_1451, v_1452, v_1453, v_1454, v_1455, v_1456, v_1457, v_1458, v_1459, v_1460, v_1461, v_1462, v_1463, v_1464, v_1465, v_1466, v_1467, v_1468, v_1469, v_1470, v_1471, v_1472, v_1473, v_1474, v_1475, v_1476, v_1477, v_1478, v_1479, v_1480, v_1481, v_1482, v_1483, v_1484, v_1485, v_1486, v_1487, v_1488, v_1489, v_1490, v_1491, v_1492, v_1493, v_1494, v_1495, v_1496, v_1497, v_1498, v_1499, v_1500, v_1501, v_1502, v_1503, v_1504, v_1505, v_1506, v_1507, v_1508, v_1509, v_1510, v_1511, v_1512, v_1513, v_1514, v_1515, v_1516, v_1517, v_1518, v_1519, v_1520, v_1521, v_1522, v_1523, v_1524, v_1525, v_1526, v_1527, v_1528, v_1529, v_1530, v_1531, v_1532, v_1533, v_1534, v_1535, v_1536, v_1537, v_1538, v_1539, v_1540, v_1541, v_1542, v_1543, v_1544, v_1545, v_1546, v_1547, v_1548, v_1549, v_1550, v_1551, v_1552, v_1553, v_1554, v_1555, v_1556, v_1557, v_1558, v_1559, v_1560, v_1561, v_1562, v_1563, v_1564, v_1565, v_1566, v_1567, v_1568, v_1569, v_1570, v_1571, v_1572, v_1573, v_1574, v_1575, v_1576, v_1577, v_1578, v_1579, v_1580, v_1581, v_1582, v_1583, v_1584, v_1585, v_1586, v_1587, v_1588, v_1589, v_1590, v_1591, v_1592, v_1593, v_1594, v_1595, v_1596, v_1597, v_1598, v_1599, v_1600, v_1601, v_1602, v_1603, v_1604, v_1605, v_1606, v_1607, v_1608, v_1609, v_1610, v_1611, v_1612, v_1613, v_1614, v_1615, v_1616, v_1617, v_1618, v_1619, v_1620, v_1621, v_1622, v_1623, v_1624, v_1625, v_1626, v_1627, v_1628, v_1629, v_1630, v_1631, v_1632, v_1633, v_1634, v_1635, v_1636, v_1637, v_1638, v_1639, v_1640, v_1641, v_1642, v_1643, v_1644, v_1645, v_1646, v_1647, v_1648, v_1649, v_1650, v_1651, v_1652, v_1653, v_1654, v_1655, v_1656, v_1657, v_1658, v_1659, v_1660, v_1661, v_1662, v_1663, v_1664, v_1665, v_1666, v_1667, v_1668, v_1669, v_1670, v_1671, v_1672, v_1673, v_1674, v_1675, v_1676, v_1677, v_1678, v_1679, v_1680, v_1681, v_1682, v_1683, v_1684, v_1685, v_1686, v_1687, v_1688, v_1689, v_1690, v_1691, v_1692, v_1693, v_1694, v_1695, v_1696, v_1697, v_1698, v_1699, v_1700, v_1701, v_1702, v_1703, v_1704, v_1705, v_1706, v_1707, v_1708, v_1709, v_1710, v_1711, v_1712, v_1713, v_1714, v_1715, v_1716, v_1717, v_1718, v_1719, v_1720, v_1721, v_1722, v_1723, v_1724, v_1725, v_1726, v_1727, v_1728, v_1729, v_1730, v_1731, v_1732, v_1733, v_1734, v_1735, v_1736, v_1737, v_1738, v_1739, v_1740, v_1741, v_1742, v_1743, v_1744, v_1745, v_1746, v_1747, v_1748, v_1749, v_1750, v_1751, v_1752, v_1753, v_1754, v_1755, v_1756, v_1757, v_1758, v_1759, v_1760, v_1761, v_1762, v_1763, v_1764, v_1765, v_1766, v_1767, v_1768, v_1769, v_1770, v_1771, v_1772, v_1773, v_1774, v_1775, v_1776, v_1777, v_1778, v_1779, v_1780, v_1781, v_1782, v_1783, v_1784, v_1785, v_1786, v_1787, v_1788, v_1789, v_1790, v_1791, v_1792, v_1793, v_1794, v_1795, v_1796, v_1797, v_1798, v_1799, v_1800, v_1801, v_1802, v_1803, v_1804, v_1805, v_1806, v_1807, v_1808, v_1809, v_1810, v_1811, v_1812, v_1813, v_1814, v_1815, v_1816, v_1817, v_1818, v_1819, v_1820, v_1821, v_1822, v_1823, v_1824, v_1825, v_1826, v_1827, v_1828, v_1829, v_1830, v_1831, v_1832, v_1833, v_1834, v_1835, v_1836, v_1837, v_1838, v_1839, v_1840, v_1841, v_1842, v_1843, v_1844, v_1845, v_1846, v_1847, v_1848, v_1849, v_1850, v_1851, v_1852, v_1853, v_1854, v_1855, v_1856, v_1857, v_1858, v_1859, v_1860, v_1861, v_1862, v_1863, v_1864, v_1865, v_1866, v_1867, v_1868, v_1869, v_1870, v_1871, v_1872, v_1873, v_1874, v_1875, v_1876, v_1877, v_1878, v_1879, v_1880, v_1881, v_1882, v_1883, v_1884, v_1885, v_1886, v_1887, v_1888, v_1889, v_1890, v_1891, v_1892, v_1893, v_1894, v_1895, v_1896, v_1897, v_1898, v_1899, v_1900, v_1901, v_1902, v_1903, v_1904, v_1905, v_1906, v_1907, v_1908, v_1909, v_1910, v_1911, v_1912, v_1913, v_1914, v_1915, v_1916, v_1917, v_1918, v_1919, v_1920, v_1921, v_1922, v_1923, v_1924, v_1925, v_1926, v_1927, v_1928, v_1929, v_1930, v_1931, v_1932, v_1933, v_1934, v_1935, v_1936, v_1937, v_1938, v_1939, v_1940, v_1941, v_1942, v_1943, v_1944, v_1945, v_1946, v_1947, v_1948, v_1949, v_1950, v_1951, v_1952, v_1953, v_1954, v_1955, v_1956, v_1957, v_1958, v_1959, v_1960, v_1961, v_1962, v_1963, v_1964, v_1965, v_1966, v_1967, v_1968, v_1969, v_1970, v_1971, v_1972, v_1973, v_1974, v_1975, v_1976, v_1977, v_1978, v_1979, v_1980, v_1981, v_1982, v_1983, v_1984, v_1985, v_1986, v_1987, v_1988, v_1989, v_1990, v_1991, v_1992, v_1993, v_1994, v_1995, v_1996, v_1997, v_1998, v_1999, v_2000, v_2001, v_2002, v_2003, v_2004, v_2005, v_2006, v_2007, v_2008, v_2009, v_2010, v_2011, v_2012, v_2013, v_2014, v_2015, v_2016, v_2017, v_2018, v_2019, v_2020, v_2021, v_2022, v_2023, v_2024, v_2025, v_2026, v_2027, v_2028, v_2029, v_2030, v_2031, v_2032, v_2033, v_2034, v_2035, v_2036, v_2037, v_2038, v_2039, v_2040, v_2041, v_2042, v_2043, v_2044, v_2045, v_2046, v_2047, v_2048, v_2049, v_2050, v_2051, v_2052, v_2053, v_2054, v_2055, v_2056, v_2057, v_2058, v_2059, v_2060, v_2061, v_2062, v_2063, v_2064, v_2065, v_2066, v_2067, v_2068, v_2069, v_2070, v_2071, v_2072, v_2073, v_2074, v_2075, v_2076, v_2077, v_2078, v_2079, v_2080, v_2081, v_2082, v_2083, v_2084, v_2085, v_2086, v_2087, v_2088, v_2089, v_2090, v_2091, v_2092, v_2093, v_2094, v_2095, v_2096, v_2097, v_2098, v_2099, v_2100, v_2101, v_2102, v_2103, v_2104, v_2105, v_2106, v_2107, v_2108, v_2109, v_2110, v_2111, v_2112, v_2113, v_2114, v_2115, v_2116, v_2117, v_2118, v_2119, v_2120, v_2121, v_2122, v_2123, v_2124, v_2125, v_2126, v_2127, v_2128, v_2129, v_2130, v_2131, v_2132, v_2133, v_2134, v_2135, v_2136, v_2137, v_2138, v_2139, v_2140, v_2141, v_2142, v_2143, v_2144, v_2145, v_2146, v_2147, v_2148, v_2149, v_2150, v_2151, v_2152, v_2153, v_2154, v_2155, v_2156, v_2157, v_2158, v_2159, v_2160, v_2161, v_2162, v_2163, v_2164, v_2165, v_2166, v_2167, v_2168, v_2169, v_2170, v_2171, v_2172, v_2173, v_2174, v_2175, v_2176, v_2177, v_2178, v_2179, v_2180, v_2181, v_2182, v_2183, v_2184, v_2185, v_2186, v_2187, v_2188, v_2189, v_2190, v_2191, v_2192, v_2193, v_2194, v_2195, v_2196, v_2197, v_2198, v_2199, v_2200, v_2201, v_2202, v_2203, v_2204, v_2205, v_2206, v_2207, v_2208, v_2209, v_2210, v_2211, v_2212, v_2213, v_2214, v_2215, v_2216, v_2217, v_2218, v_2219, v_2220, v_2221, v_2222, v_2223, v_2224, v_2225, v_2226, v_2227, v_2228, v_2229, v_2230, v_2231, v_2232, v_2233, v_2234, v_2235, v_2236, v_2237, v_2238, v_2239, v_2240, v_2241, v_2242, v_2243, v_2244, v_2245, v_2246, v_2247, v_2248, v_2249, v_2250, v_2251, v_2252, v_2253, v_2254, v_2255, v_2256, v_2257, v_2258, v_2259, v_2260, v_2261, v_2262, v_2263, v_2264, v_2265, v_2266, v_2267, v_2268, v_2269, v_2270, v_2271, v_2272, v_2273, v_2274, v_2275, v_2276, v_2277, v_2278, v_2279, v_2280, v_2281, v_2282, v_2283, v_2284, v_2285, v_2286, v_2287, v_2288, v_2289, v_2290, v_2291, v_2292, v_2293, v_2294, v_2295, v_2296, v_2297, v_2298, v_2299, v_2300, v_2301, v_2302, v_2303, v_2304, v_2305, v_2306, v_2307, v_2308, v_2309, v_2310, v_2311, v_2312, v_2313, v_2314, v_2315, v_2316, v_2317, v_2318, v_2319, v_2320, v_2321, v_2322, v_2323, v_2324, v_2325, v_2326, v_2327, v_2328, v_2329, v_2330, v_2331, v_2332, v_2333, v_2334, v_2335, v_2336, v_2337, v_2338, v_2339, v_2340, v_2341, v_2342, v_2343, v_2344, v_2345, v_2346, v_2347, v_2348, v_2349, v_2350, v_2351, v_2352, v_2353, v_2354, v_2355, v_2356, v_2357, v_2358, v_2359, v_2360, v_2361, v_2362, v_2363, v_2364, v_2365, v_2366, v_2367, v_2368, v_2369, v_2370, v_2371, v_2372, v_2373, v_2374, v_2375, v_2376, v_2377, v_2378, v_2379, v_2380, v_2381, v_2382, v_2383, v_2384, v_2385, v_2386, v_2387, v_2388, v_2389, v_2390, v_2391, v_2392, v_2393, v_2394, v_2395, v_2396, v_2397, v_2398, v_2399, v_2400, v_2401, v_2402, v_2403, v_2404, v_2405, v_2406, v_2407, v_2408, v_2409, v_2410, v_2411, v_2412, v_2413, v_2414, v_2415, v_2416, v_2417, v_2418, v_2419, v_2420, v_2421, v_2422, v_2423, v_2424, v_2425, v_2426, v_2427, v_2428, v_2429, v_2430, v_2431, v_2432, v_2433, v_2434, v_2435, v_2436, v_2437, v_2438, v_2439, v_2440, v_2441, v_2442, v_2443, v_2444, v_2445, v_2446, v_2447, v_2448, v_2449, v_2450, v_2451, v_2452, v_2453, v_2454, v_2455, v_2456, v_2457, v_2458, v_2459, v_2460, v_2461, v_2462, v_2463, v_2464, v_2465, v_2466, v_2467, v_2468, v_2469, v_2470, v_2471, v_2472, v_2473, v_2474, v_2475, v_2476, v_2477, v_2478, v_2479, v_2480, v_2481, v_2482, v_2483, v_2484, v_2485, v_2486, v_2487, v_2488, v_2489, v_2490, v_2491, v_2492, v_2493, v_2494, v_2495, v_2496, v_2497, v_2498, v_2499, v_2500, v_2501, v_2502, v_2503, v_2504, v_2505, v_2506, v_2507, v_2508, v_2509, v_2510, v_2511, v_2512, v_2513, v_2514, v_2515, v_2516, v_2517, v_2518, v_2519, v_2520, v_2521, v_2522, v_2523, v_2524, v_2525, v_2526, v_2527, v_2528, v_2529, v_2530, v_2531, v_2532, v_2533, v_2534, v_2535, v_2536, v_2537, v_2538, v_2539, v_2540, v_2541, v_2542, v_2543, v_2544, v_2545, v_2546, v_2547, v_2548, v_2549, v_2550, v_2551, v_2552, v_2553, v_2554, v_2555, v_2556, v_2557, v_2558, v_2559, v_2560, v_2561, v_2562, v_2563, v_2564, v_2565, v_2566, v_2567, v_2568, v_2569, v_2570, v_2571, v_2572, v_2573, v_2574, v_2575, v_2576, v_2577, v_2578, v_2579, v_2580, v_2581, v_2582, v_2583, v_2584, v_2585, v_2586, v_2587, v_2588, v_2589, v_2590, v_2591, v_2592, v_2593, v_2594, v_2595, v_2596, v_2597, v_2598, v_2599, v_2600, v_2601, v_2602, v_2603, v_2604, v_2605, v_2606, v_2607, v_2608, v_2609, v_2610, v_2611, v_2612, v_2613, v_2614, v_2615, v_2616, v_2617, v_2618, v_2619, v_2620, v_2621, v_2622, v_2623, v_2624, v_2625, v_2626, v_2627, v_2628, v_2629, v_2630, v_2631, v_2632, v_2633, v_2634, v_2635, v_2636, v_2637, v_2638, v_2639, v_2640, v_2641, v_2642, v_2643, v_2644, v_2645, v_2646, v_2647, v_2648, v_2649, v_2650, v_2651, v_2652, v_2653, v_2654, v_2655, v_2656, v_2657, v_2658, v_2659, v_2660, v_2661, v_2662, v_2663, v_2664, v_2665, v_2666, v_2667, v_2668, v_2669, v_2670, v_2671, v_2672, v_2673, v_2674, v_2675, v_2676, v_2677, v_2678, v_2679, v_2680, v_2681, v_2682, v_2683, v_2684, v_2685, v_2686, v_2687, v_2688, v_2689, v_2690, v_2691, v_2692, v_2693, v_2694, v_2695, v_2696, v_2697, v_2698, v_2699, v_2700, v_2701, v_2702, v_2703, v_2704, v_2705, v_2706, v_2707, v_2708, v_2709, v_2710, v_2711, v_2712, v_2713, v_2714, v_2715, v_2716, v_2717, v_2718, v_2719, v_2720, v_2721, v_2722, v_2723, v_2724, v_2725, v_2726, v_2727, v_2728, v_2729, v_2730, v_2731, v_2732, v_2733, v_2734, v_2735, v_2736, v_2737, v_2738, v_2739, v_2740, v_2741, v_2742, v_2743, v_2744, v_2745, v_2746, v_2747, v_2748, v_2749, v_2750, v_2751, v_2752, v_2753, v_2754, v_2755, v_2756, v_2757, v_2758, v_2759, v_2760, v_2761, v_2762, v_2763, v_2764, v_2765, v_2766, v_2767, v_2768, v_2769, v_2770, v_2771, v_2772, v_2773, v_2774, v_2775, v_2776, v_2777, v_2778, v_2779, v_2780, v_2781, v_2782, v_2783, v_2784, v_2785, v_2786, v_2787, v_2788, v_2789, v_2790, v_2791, v_2792, v_2793, v_2794, v_2795, v_2796, v_2797, v_2798, v_2799, v_2800, v_2801, v_2802, v_2803, v_2804, v_2805, v_2806, v_2807, v_2808, v_2809, v_2810, v_2811, v_2812, v_2813, v_2814, v_2815, v_2816, v_2817, v_2818, v_2819, v_2820, v_2821, v_2822, v_2823, v_2824, v_2825, v_2826, v_2827, v_2828, v_2829, v_2830, v_2831, v_2832, v_2833, v_2834, v_2835, v_2836, v_2837, v_2838, v_2839, v_2840, v_2841, v_2842, v_2843, v_2844, v_2845, v_2846, v_2847, v_2848, v_2849, v_2850, v_2851, v_2852, v_2853, v_2854, v_2855, v_2856, v_2857, v_2858, v_2859, v_2860, v_2861, v_2862, v_2863, v_2864, v_2865, v_2866, v_2867, v_2868, v_2869, v_2870, v_2871, v_2872, v_2873, v_2874, v_2875, v_2876, v_2877, v_2878, v_2879, v_2880, v_2881, v_2882, v_2883, v_2884, v_2885, v_2886, v_2887, v_2888, v_2889, v_2890, v_2891, v_2892, v_2893, v_2894, v_2895, v_2896, v_2897, v_2898, v_2899, v_2900, v_2901, v_2902, v_2903, v_2904, v_2905, v_2906, v_2907, v_2908, v_2909, v_2910, v_2911, v_2912, v_2913, v_2914, v_2915, v_2916, v_2917, v_2918, v_2919, v_2920, v_2921, v_2922, v_2923, v_2924, v_2925, v_2926, v_2927, v_2928, v_2929, v_2930, v_2931, v_2932, v_2933, v_2934, v_2935, v_2936, v_2937, v_2938, v_2939, v_2940, v_2941, v_2942, v_2943, v_2944, v_2945, v_2946, v_2947, v_2948, v_2949, v_2950, v_2951, v_2952, v_2953, v_2954, v_2955, v_2956, v_2957, v_2958, v_2959, v_2960, v_2961, v_2962, v_2963, v_2964, v_2965, v_2966, v_2967, v_2968, v_2969, v_2970, v_2971, v_2972, v_2973, v_2974, v_2975, v_2976, v_2977, v_2978, v_2979, v_2980, v_2981, v_2982, v_2983, v_2984, v_2985, v_2986, v_2987, v_2988, v_2989, v_2990, v_2991, v_2992, v_2993, v_2994, v_2995, v_2996, v_2997, v_2998, v_2999, v_3000, v_3001, v_3002, v_3003, v_3004, v_3005, v_3006, v_3007, v_3008, v_3009, v_3010, v_3011, v_3012, v_3013, v_3014, v_3015, v_3016, v_3017, v_3018, v_3019, v_3020, v_3021, v_3022, v_3023, v_3024, v_3025, v_3026, v_3027, v_3028, v_3029, v_3030, v_3031, v_3032, v_3033, v_3034, v_3035, v_3036, v_3037, v_3038, v_3039, v_3040, v_3041, v_3042, v_3043, v_3044, v_3045, v_3046, v_3047, v_3048, v_3049, v_3050, v_3051, v_3052, v_3053, v_3054, v_3055, v_3056, v_3057, v_3058, v_3059, v_3060, v_3061, v_3062, v_3063, v_3064, v_3065, v_3066, v_3067, v_3068, v_3069, v_3070, v_3071, v_3072, v_3073, v_3074, v_3075, v_3076, v_3077, v_3078, v_3079, v_3080, v_3081, v_3082, v_3083, v_3084, v_3085, v_3086, v_3087, v_3088, v_3089, v_3090, v_3091, v_3092, v_3093, v_3094, v_3095, v_3096, v_3097, v_3098, v_3099, v_3100, v_3101, v_3102, v_3103, v_3104, v_3105, v_3106, v_3107, v_3108, v_3109, v_3110, v_3111, v_3112, v_3113, v_3114, v_3115, v_3116, v_3117, v_3118, v_3119, v_3120, v_3121, v_3122, v_3123, v_3124, v_3125, v_3126, v_3127, v_3128, v_3129, v_3130, v_3131, v_3132, v_3133, v_3134, v_3135, v_3136, v_3137, v_3138, v_3139, v_3140, v_3141, v_3142, v_3143, v_3144, v_3145, v_3146, v_3147, v_3148, v_3149, v_3150, v_3151, v_3152, v_3153, v_3154, v_3155, v_3156, v_3157, v_3158, v_3159, v_3160, v_3161, v_3162, v_3163, v_3164, v_3165, v_3166, v_3167, v_3168, v_3169, v_3170, v_3171, v_3172, v_3173, v_3174, v_3175, v_3176, v_3177, v_3178, v_3179, v_3180, v_3181, v_3182, v_3183, v_3184, v_3185, v_3186, v_3187, v_3188, v_3189, v_3190, v_3191, v_3192, v_3193, v_3194, v_3195, v_3196, v_3197, v_3198, v_3199, v_3200, v_3201, v_3202, v_3203, v_3204, v_3205, v_3206, v_3207, v_3208, v_3209, v_3210, v_3211, v_3212, v_3213, v_3214, v_3215, v_3216, v_3217, v_3218, v_3219, v_3220, v_3221, v_3222, v_3223, v_3224, v_3225, v_3226, v_3227, v_3228, v_3229, v_3230, v_3231, v_3232, v_3233, v_3234, v_3235, v_3236, v_3237, v_3238, v_3239, v_3240, v_3241, v_3242, v_3243, v_3244, v_3245, v_3246, v_3247, v_3248, v_3249, v_3250, v_3251, v_3252, v_3253, v_3254, v_3255, v_3256, v_3257, v_3258, v_3259, v_3260, v_3261, v_3262, v_3263, v_3264, v_3265, v_3266, v_3267, v_3268, v_3269, v_3270, v_3271, v_3272, v_3273, v_3274, v_3275, v_3276, v_3277, v_3278, v_3279, v_3280, v_3281, v_3282, v_3283, v_3284, v_3285, v_3286, v_3287, v_3288, v_3289, v_3290, v_3291, v_3292, v_3293, v_3294, v_3295, v_3296, v_3297, v_3298, v_3299, v_3300, v_3301, v_3302, v_3303, v_3304, v_3305, v_3306, v_3307, v_3308, v_3309, v_3310, v_3311, v_3312, v_3313, v_3314, v_3315, v_3316, v_3317, v_3318, v_3319, v_3320, v_3321, v_3322, v_3323, v_3324, v_3325, v_3326, v_3327, v_3328, v_3329, v_3330, v_3331, v_3332, v_3333, v_3334, v_3335, v_3336, v_3337, v_3338, v_3339, v_3340, v_3341, v_3342, v_3343, v_3344, v_3345, v_3346, v_3347, v_3348, v_3349, v_3350, v_3351, v_3352, v_3353, v_3354, v_3355, v_3356, v_3357, v_3358, v_3359, v_3360, v_3361, v_3362, v_3363, v_3364, v_3365, v_3366, v_3367, v_3368, v_3369, v_3370, v_3371, v_3372, v_3373, v_3374, v_3375, v_3376, v_3377, v_3378, v_3379, v_3380, v_3381, v_3382, v_3383, v_3384, v_3385, v_3386, v_3387, v_3388, v_3389, v_3390, v_3391, v_3392, v_3393, v_3394, v_3395, v_3396, v_3397, v_3398, v_3399, v_3544, v_3545, v_3546, v_3547, v_3548, v_3549, v_3550, v_3551, v_3552, v_3553, v_3554, v_3555, v_3556, v_3557, v_3558, v_3559, v_3560, v_3561, v_3562, v_3563, v_3564, v_3565, v_3566, v_3567, v_3568, v_3569, v_3570, v_3571, v_3572, v_3573, v_3574, v_3575, v_3576, v_3577, v_3578, v_3579, v_3580, v_3581, v_3582, v_3583, v_3584, v_3585, v_3586, v_3587, v_3588, v_3589, v_3590, v_3591, v_3592, v_3593, v_3594, v_3595, v_3596, v_3597, v_3598, v_3599, v_3600, v_3601, v_3602, v_3603, v_3604, v_3605, v_3606, v_3607, v_3608, v_3609, v_3610, v_3611, v_3612, v_3613, v_3614, v_3615, v_3616, v_3617, v_3618, v_3619, v_3620, v_3621, v_3622, v_3623, v_3624, v_3625, v_3626, v_3627, v_3628, v_3629, v_3630, v_3631, v_3632, v_3633, v_3778, v_3779, v_3780, v_3781, v_3782, v_3783, v_3784, v_3785, v_3786, v_3787, v_3788, v_3789, v_3790, v_3791, v_3792, v_3793, v_3794, v_3795, v_3796, v_3797, v_3798, v_3799, v_3800, v_3801, v_3802, v_3803, v_3804, v_3805, v_3806, v_3807, v_3808, v_3809, v_3810, v_3811, v_3812, v_3813, v_3814, v_3815, v_3816, v_3817, v_3818, v_3819, v_3820, v_3821, v_3822, v_3823, v_3824, v_3825, v_3826, v_3827, v_3828, v_3829, v_3830, v_3831, v_3832, v_3833, v_3834, v_3835, v_3836, v_3837, v_3838, v_3839, v_3840, v_3841, v_3842, v_3843, v_3844, v_3845, v_3846, v_3847, v_3848, v_3849, v_3850, v_3851, v_3852, v_3853, v_3854, v_3855, v_3856, v_3857, v_3858, v_3859, v_3860, v_3861, v_3862, v_3863, v_3864, v_3865, v_3866, v_3867, v_4012, v_4013, v_4014, v_4015, v_4016, v_4017, v_4018, v_4019, v_4020, v_4021, v_4022, v_4023, v_4024, v_4025, v_4026, v_4027, v_4028, v_4029, v_4030, v_4031, v_4032, v_4033, v_4034, v_4035, v_4036, v_4037, v_4038, v_4039, v_4040, v_4041, v_4042, v_4043, v_4044, v_4045, v_4046, v_4047, v_4048, v_4049, v_4050, v_4051, v_4052, v_4053, v_4054, v_4055, v_4056, v_4057, v_4058, v_4059, v_4060, v_4061, v_4062, v_4063, v_4064, v_4065, v_4066, v_4067, v_4068, v_4069, v_4070, v_4071, v_4072, v_4073, v_4074, v_4075, v_4076, v_4077, v_4078, v_4079, v_4080, v_4081, v_4082, v_4083, v_4084, v_4085, v_4086, v_4087, v_4088, v_4089, v_4090, v_4091, v_4092, v_4093, v_4094, v_4095, v_4096, v_4097, v_4098, v_4099, v_4100, v_4101, o_1);
input v_56;
input v_57;
input v_58;
input v_59;
input v_60;
input v_61;
input v_62;
input v_63;
input v_64;
input v_65;
input v_66;
input v_67;
input v_68;
input v_69;
input v_70;
input v_71;
input v_72;
input v_73;
input v_74;
input v_75;
input v_76;
input v_77;
input v_78;
input v_79;
input v_80;
input v_81;
input v_82;
input v_83;
input v_84;
input v_85;
input v_86;
input v_87;
input v_88;
input v_89;
input v_90;
input v_91;
input v_92;
input v_93;
input v_94;
input v_95;
input v_96;
input v_97;
input v_98;
input v_99;
input v_100;
input v_101;
input v_102;
input v_103;
input v_104;
input v_105;
input v_106;
input v_107;
input v_108;
input v_109;
input v_110;
input v_111;
input v_112;
input v_113;
input v_114;
input v_115;
input v_116;
input v_117;
input v_118;
input v_119;
input v_120;
input v_121;
input v_122;
input v_123;
input v_124;
input v_125;
input v_126;
input v_127;
input v_128;
input v_129;
input v_130;
input v_131;
input v_132;
input v_133;
input v_134;
input v_135;
input v_136;
input v_137;
input v_138;
input v_139;
input v_140;
input v_141;
input v_142;
input v_143;
input v_144;
input v_145;
input v_146;
input v_147;
input v_148;
input v_149;
input v_150;
input v_151;
input v_152;
input v_153;
input v_154;
input v_155;
input v_156;
input v_157;
input v_158;
input v_159;
input v_160;
input v_161;
input v_162;
input v_163;
input v_164;
input v_165;
input v_166;
input v_167;
input v_168;
input v_169;
input v_170;
input v_171;
input v_172;
input v_173;
input v_174;
input v_175;
input v_176;
input v_177;
input v_178;
input v_179;
input v_180;
input v_181;
input v_182;
input v_183;
input v_184;
input v_185;
input v_186;
input v_187;
input v_188;
input v_189;
input v_190;
input v_191;
input v_192;
input v_193;
input v_194;
input v_195;
input v_196;
input v_197;
input v_198;
input v_199;
input v_200;
input v_201;
input v_202;
input v_203;
input v_204;
input v_205;
input v_206;
input v_207;
input v_208;
input v_209;
input v_210;
input v_211;
input v_212;
input v_213;
input v_214;
input v_215;
input v_216;
input v_217;
input v_218;
input v_219;
input v_220;
input v_221;
input v_222;
input v_223;
input v_224;
input v_225;
input v_226;
input v_227;
input v_228;
input v_229;
input v_230;
input v_231;
input v_232;
input v_233;
input v_234;
input v_235;
input v_236;
input v_237;
input v_238;
input v_239;
input v_240;
input v_241;
input v_242;
input v_243;
input v_244;
input v_245;
input v_246;
input v_247;
input v_248;
input v_249;
input v_250;
input v_251;
input v_252;
input v_253;
input v_254;
input v_255;
input v_256;
input v_257;
input v_258;
input v_259;
input v_260;
input v_261;
input v_262;
input v_263;
input v_264;
input v_265;
input v_266;
input v_267;
input v_268;
input v_269;
input v_270;
input v_271;
input v_272;
input v_273;
input v_274;
input v_275;
input v_276;
input v_277;
input v_278;
input v_279;
input v_280;
input v_281;
input v_282;
input v_283;
input v_284;
input v_285;
input v_286;
input v_287;
input v_288;
input v_289;
input v_290;
input v_291;
input v_292;
input v_293;
input v_294;
input v_295;
input v_296;
input v_297;
input v_298;
input v_299;
input v_300;
input v_301;
input v_302;
input v_303;
input v_304;
input v_305;
input v_306;
input v_307;
input v_308;
input v_309;
input v_310;
input v_311;
input v_312;
input v_313;
input v_314;
input v_315;
input v_316;
input v_317;
input v_318;
input v_319;
input v_320;
input v_321;
input v_322;
input v_323;
input v_324;
input v_325;
input v_326;
input v_327;
input v_328;
input v_329;
input v_330;
input v_331;
input v_332;
input v_333;
input v_334;
input v_335;
input v_336;
input v_337;
input v_338;
input v_339;
input v_340;
input v_341;
input v_342;
input v_343;
input v_344;
input v_345;
input v_346;
input v_347;
input v_348;
input v_349;
input v_350;
input v_351;
input v_352;
input v_353;
input v_354;
input v_355;
input v_356;
input v_357;
input v_358;
input v_359;
input v_360;
input v_361;
input v_362;
input v_363;
input v_364;
input v_365;
input v_366;
input v_367;
input v_368;
input v_369;
input v_370;
input v_371;
input v_372;
input v_373;
input v_374;
input v_375;
input v_376;
input v_377;
input v_378;
input v_379;
input v_3400;
input v_3401;
input v_3402;
input v_3403;
input v_3404;
input v_3405;
input v_3406;
input v_3407;
input v_3408;
input v_3409;
input v_3410;
input v_3411;
input v_3412;
input v_3413;
input v_3414;
input v_3415;
input v_3416;
input v_3417;
input v_3418;
input v_3419;
input v_3420;
input v_3421;
input v_3422;
input v_3423;
input v_3424;
input v_3425;
input v_3426;
input v_3427;
input v_3428;
input v_3429;
input v_3430;
input v_3431;
input v_3432;
input v_3433;
input v_3434;
input v_3435;
input v_3436;
input v_3437;
input v_3438;
input v_3439;
input v_3440;
input v_3441;
input v_3442;
input v_3443;
input v_3444;
input v_3445;
input v_3446;
input v_3447;
input v_3448;
input v_3449;
input v_3450;
input v_3451;
input v_3452;
input v_3453;
input v_3454;
input v_3455;
input v_3456;
input v_3457;
input v_3458;
input v_3459;
input v_3460;
input v_3461;
input v_3462;
input v_3463;
input v_3464;
input v_3465;
input v_3466;
input v_3467;
input v_3468;
input v_3469;
input v_3470;
input v_3471;
input v_3472;
input v_3473;
input v_3474;
input v_3475;
input v_3476;
input v_3477;
input v_3478;
input v_3479;
input v_3480;
input v_3481;
input v_3482;
input v_3483;
input v_3484;
input v_3485;
input v_3486;
input v_3487;
input v_3488;
input v_3489;
input v_3490;
input v_3491;
input v_3492;
input v_3493;
input v_3494;
input v_3495;
input v_3496;
input v_3497;
input v_3498;
input v_3499;
input v_3500;
input v_3501;
input v_3502;
input v_3503;
input v_3504;
input v_3505;
input v_3506;
input v_3507;
input v_3508;
input v_3509;
input v_3510;
input v_3511;
input v_3512;
input v_3513;
input v_3514;
input v_3515;
input v_3516;
input v_3517;
input v_3518;
input v_3519;
input v_3520;
input v_3521;
input v_3522;
input v_3523;
input v_3524;
input v_3525;
input v_3526;
input v_3527;
input v_3528;
input v_3529;
input v_3530;
input v_3531;
input v_3532;
input v_3533;
input v_3534;
input v_3535;
input v_3536;
input v_3537;
input v_3538;
input v_3539;
input v_3540;
input v_3541;
input v_3542;
input v_3543;
input v_3634;
input v_3635;
input v_3636;
input v_3637;
input v_3638;
input v_3639;
input v_3640;
input v_3641;
input v_3642;
input v_3643;
input v_3644;
input v_3645;
input v_3646;
input v_3647;
input v_3648;
input v_3649;
input v_3650;
input v_3651;
input v_3652;
input v_3653;
input v_3654;
input v_3655;
input v_3656;
input v_3657;
input v_3658;
input v_3659;
input v_3660;
input v_3661;
input v_3662;
input v_3663;
input v_3664;
input v_3665;
input v_3666;
input v_3667;
input v_3668;
input v_3669;
input v_3670;
input v_3671;
input v_3672;
input v_3673;
input v_3674;
input v_3675;
input v_3676;
input v_3677;
input v_3678;
input v_3679;
input v_3680;
input v_3681;
input v_3682;
input v_3683;
input v_3684;
input v_3685;
input v_3686;
input v_3687;
input v_3688;
input v_3689;
input v_3690;
input v_3691;
input v_3692;
input v_3693;
input v_3694;
input v_3695;
input v_3696;
input v_3697;
input v_3698;
input v_3699;
input v_3700;
input v_3701;
input v_3702;
input v_3703;
input v_3704;
input v_3705;
input v_3706;
input v_3707;
input v_3708;
input v_3709;
input v_3710;
input v_3711;
input v_3712;
input v_3713;
input v_3714;
input v_3715;
input v_3716;
input v_3717;
input v_3718;
input v_3719;
input v_3720;
input v_3721;
input v_3722;
input v_3723;
input v_3724;
input v_3725;
input v_3726;
input v_3727;
input v_3728;
input v_3729;
input v_3730;
input v_3731;
input v_3732;
input v_3733;
input v_3734;
input v_3735;
input v_3736;
input v_3737;
input v_3738;
input v_3739;
input v_3740;
input v_3741;
input v_3742;
input v_3743;
input v_3744;
input v_3745;
input v_3746;
input v_3747;
input v_3748;
input v_3749;
input v_3750;
input v_3751;
input v_3752;
input v_3753;
input v_3754;
input v_3755;
input v_3756;
input v_3757;
input v_3758;
input v_3759;
input v_3760;
input v_3761;
input v_3762;
input v_3763;
input v_3764;
input v_3765;
input v_3766;
input v_3767;
input v_3768;
input v_3769;
input v_3770;
input v_3771;
input v_3772;
input v_3773;
input v_3774;
input v_3775;
input v_3776;
input v_3777;
input v_3868;
input v_3869;
input v_3870;
input v_3871;
input v_3872;
input v_3873;
input v_3874;
input v_3875;
input v_3876;
input v_3877;
input v_3878;
input v_3879;
input v_3880;
input v_3881;
input v_3882;
input v_3883;
input v_3884;
input v_3885;
input v_3886;
input v_3887;
input v_3888;
input v_3889;
input v_3890;
input v_3891;
input v_3892;
input v_3893;
input v_3894;
input v_3895;
input v_3896;
input v_3897;
input v_3898;
input v_3899;
input v_3900;
input v_3901;
input v_3902;
input v_3903;
input v_3904;
input v_3905;
input v_3906;
input v_3907;
input v_3908;
input v_3909;
input v_3910;
input v_3911;
input v_3912;
input v_3913;
input v_3914;
input v_3915;
input v_3916;
input v_3917;
input v_3918;
input v_3919;
input v_3920;
input v_3921;
input v_3922;
input v_3923;
input v_3924;
input v_3925;
input v_3926;
input v_3927;
input v_3928;
input v_3929;
input v_3930;
input v_3931;
input v_3932;
input v_3933;
input v_3934;
input v_3935;
input v_3936;
input v_3937;
input v_3938;
input v_3939;
input v_3940;
input v_3941;
input v_3942;
input v_3943;
input v_3944;
input v_3945;
input v_3946;
input v_3947;
input v_3948;
input v_3949;
input v_3950;
input v_3951;
input v_3952;
input v_3953;
input v_3954;
input v_3955;
input v_3956;
input v_3957;
input v_3958;
input v_3959;
input v_3960;
input v_3961;
input v_3962;
input v_3963;
input v_3964;
input v_3965;
input v_3966;
input v_3967;
input v_3968;
input v_3969;
input v_3970;
input v_3971;
input v_3972;
input v_3973;
input v_3974;
input v_3975;
input v_3976;
input v_3977;
input v_3978;
input v_3979;
input v_3980;
input v_3981;
input v_3982;
input v_3983;
input v_3984;
input v_3985;
input v_3986;
input v_3987;
input v_3988;
input v_3989;
input v_3990;
input v_3991;
input v_3992;
input v_3993;
input v_3994;
input v_3995;
input v_3996;
input v_3997;
input v_3998;
input v_3999;
input v_4000;
input v_4001;
input v_4002;
input v_4003;
input v_4004;
input v_4005;
input v_4006;
input v_4007;
input v_4008;
input v_4009;
input v_4010;
input v_4011;
input v_1;
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_13;
input v_14;
input v_15;
input v_16;
input v_17;
input v_18;
input v_19;
input v_20;
input v_21;
input v_22;
input v_23;
input v_24;
input v_25;
input v_26;
input v_27;
input v_28;
input v_29;
input v_30;
input v_31;
input v_32;
input v_33;
input v_34;
input v_35;
input v_36;
input v_37;
input v_38;
input v_39;
input v_40;
input v_41;
input v_42;
input v_43;
input v_44;
input v_45;
input v_46;
input v_47;
input v_48;
input v_49;
input v_50;
input v_51;
input v_52;
input v_53;
input v_54;
input v_55;
input v_380;
input v_381;
input v_382;
input v_383;
input v_384;
input v_385;
input v_386;
input v_387;
input v_388;
input v_389;
input v_390;
input v_391;
input v_392;
input v_393;
input v_394;
input v_395;
input v_396;
input v_397;
input v_398;
input v_399;
input v_400;
input v_401;
input v_402;
input v_403;
input v_404;
input v_405;
input v_406;
input v_407;
input v_408;
input v_409;
input v_410;
input v_411;
input v_412;
input v_413;
input v_414;
input v_415;
input v_416;
input v_417;
input v_418;
input v_419;
input v_420;
input v_421;
input v_422;
input v_423;
input v_424;
input v_425;
input v_426;
input v_427;
input v_428;
input v_429;
input v_430;
input v_431;
input v_432;
input v_433;
input v_434;
input v_435;
input v_436;
input v_437;
input v_438;
input v_439;
input v_440;
input v_441;
input v_442;
input v_443;
input v_444;
input v_445;
input v_446;
input v_447;
input v_448;
input v_449;
input v_450;
input v_451;
input v_452;
input v_453;
input v_454;
input v_455;
input v_456;
input v_457;
input v_458;
input v_459;
input v_460;
input v_461;
input v_462;
input v_463;
input v_464;
input v_465;
input v_466;
input v_467;
input v_468;
input v_469;
input v_470;
input v_471;
input v_472;
input v_473;
input v_474;
input v_475;
input v_476;
input v_477;
input v_478;
input v_479;
input v_480;
input v_481;
input v_482;
input v_483;
input v_484;
input v_485;
input v_486;
input v_487;
input v_488;
input v_489;
input v_490;
input v_491;
input v_492;
input v_493;
input v_494;
input v_495;
input v_496;
input v_497;
input v_498;
input v_499;
input v_500;
input v_501;
input v_502;
input v_503;
input v_504;
input v_505;
input v_506;
input v_507;
input v_508;
input v_509;
input v_510;
input v_511;
input v_512;
input v_513;
input v_514;
input v_515;
input v_516;
input v_517;
input v_518;
input v_519;
input v_520;
input v_521;
input v_522;
input v_523;
input v_524;
input v_525;
input v_526;
input v_527;
input v_528;
input v_529;
input v_530;
input v_531;
input v_532;
input v_533;
input v_534;
input v_535;
input v_536;
input v_537;
input v_538;
input v_539;
input v_540;
input v_541;
input v_542;
input v_543;
input v_544;
input v_545;
input v_546;
input v_547;
input v_548;
input v_549;
input v_550;
input v_551;
input v_552;
input v_553;
input v_554;
input v_555;
input v_556;
input v_557;
input v_558;
input v_559;
input v_560;
input v_561;
input v_562;
input v_563;
input v_564;
input v_565;
input v_566;
input v_567;
input v_568;
input v_569;
input v_570;
input v_571;
input v_572;
input v_573;
input v_574;
input v_575;
input v_576;
input v_577;
input v_578;
input v_579;
input v_580;
input v_581;
input v_582;
input v_583;
input v_584;
input v_585;
input v_586;
input v_587;
input v_588;
input v_589;
input v_590;
input v_591;
input v_592;
input v_593;
input v_594;
input v_595;
input v_596;
input v_597;
input v_598;
input v_599;
input v_600;
input v_601;
input v_602;
input v_603;
input v_604;
input v_605;
input v_606;
input v_607;
input v_608;
input v_609;
input v_610;
input v_611;
input v_612;
input v_613;
input v_614;
input v_615;
input v_616;
input v_617;
input v_618;
input v_619;
input v_620;
input v_621;
input v_622;
input v_623;
input v_624;
input v_625;
input v_626;
input v_627;
input v_628;
input v_629;
input v_630;
input v_631;
input v_632;
input v_633;
input v_634;
input v_635;
input v_636;
input v_637;
input v_638;
input v_639;
input v_640;
input v_641;
input v_642;
input v_643;
input v_644;
input v_645;
input v_646;
input v_647;
input v_648;
input v_649;
input v_650;
input v_651;
input v_652;
input v_653;
input v_654;
input v_655;
input v_656;
input v_657;
input v_658;
input v_659;
input v_705;
input v_706;
input v_707;
input v_708;
input v_709;
input v_710;
input v_711;
input v_712;
input v_713;
input v_714;
input v_715;
input v_716;
input v_717;
input v_718;
input v_719;
input v_720;
input v_721;
input v_722;
input v_723;
input v_724;
input v_725;
input v_726;
input v_727;
input v_728;
input v_729;
input v_730;
input v_731;
input v_732;
input v_733;
input v_734;
input v_735;
input v_736;
input v_737;
input v_738;
input v_739;
input v_740;
input v_741;
input v_742;
input v_743;
input v_744;
input v_745;
input v_746;
input v_747;
input v_748;
input v_749;
input v_750;
input v_751;
input v_752;
input v_753;
input v_754;
input v_755;
input v_756;
input v_757;
input v_758;
input v_759;
input v_760;
input v_761;
input v_762;
input v_763;
input v_764;
input v_765;
input v_766;
input v_767;
input v_768;
input v_769;
input v_770;
input v_771;
input v_772;
input v_773;
input v_774;
input v_775;
input v_776;
input v_777;
input v_778;
input v_779;
input v_780;
input v_781;
input v_782;
input v_783;
input v_784;
input v_785;
input v_786;
input v_787;
input v_788;
input v_789;
input v_790;
input v_791;
input v_792;
input v_793;
input v_794;
input v_795;
input v_796;
input v_797;
input v_798;
input v_799;
input v_800;
input v_801;
input v_802;
input v_803;
input v_804;
input v_805;
input v_806;
input v_807;
input v_808;
input v_809;
input v_810;
input v_811;
input v_812;
input v_813;
input v_814;
input v_815;
input v_816;
input v_817;
input v_818;
input v_819;
input v_820;
input v_821;
input v_822;
input v_823;
input v_824;
input v_825;
input v_826;
input v_827;
input v_828;
input v_829;
input v_830;
input v_831;
input v_832;
input v_833;
input v_834;
input v_835;
input v_836;
input v_837;
input v_838;
input v_839;
input v_840;
input v_841;
input v_842;
input v_843;
input v_844;
input v_845;
input v_846;
input v_847;
input v_848;
input v_849;
input v_850;
input v_851;
input v_852;
input v_853;
input v_854;
input v_855;
input v_856;
input v_857;
input v_858;
input v_859;
input v_860;
input v_861;
input v_862;
input v_863;
input v_864;
input v_865;
input v_866;
input v_867;
input v_868;
input v_869;
input v_870;
input v_871;
input v_872;
input v_873;
input v_874;
input v_875;
input v_876;
input v_877;
input v_878;
input v_879;
input v_880;
input v_881;
input v_882;
input v_883;
input v_884;
input v_885;
input v_931;
input v_932;
input v_933;
input v_934;
input v_935;
input v_936;
input v_937;
input v_938;
input v_939;
input v_940;
input v_941;
input v_942;
input v_943;
input v_944;
input v_945;
input v_946;
input v_947;
input v_948;
input v_949;
input v_950;
input v_951;
input v_952;
input v_953;
input v_954;
input v_955;
input v_956;
input v_957;
input v_958;
input v_959;
input v_960;
input v_961;
input v_962;
input v_963;
input v_964;
input v_965;
input v_966;
input v_967;
input v_968;
input v_969;
input v_970;
input v_971;
input v_972;
input v_973;
input v_974;
input v_975;
input v_976;
input v_977;
input v_978;
input v_979;
input v_980;
input v_981;
input v_982;
input v_983;
input v_984;
input v_985;
input v_986;
input v_987;
input v_988;
input v_989;
input v_990;
input v_991;
input v_992;
input v_993;
input v_994;
input v_995;
input v_996;
input v_997;
input v_998;
input v_999;
input v_1000;
input v_1001;
input v_1002;
input v_1003;
input v_1004;
input v_1005;
input v_1006;
input v_1007;
input v_1008;
input v_1009;
input v_1010;
input v_1011;
input v_1012;
input v_1013;
input v_1014;
input v_1015;
input v_1016;
input v_1017;
input v_1018;
input v_1019;
input v_1020;
input v_1021;
input v_1022;
input v_1023;
input v_1024;
input v_1025;
input v_1026;
input v_1027;
input v_1028;
input v_1029;
input v_1030;
input v_1031;
input v_1032;
input v_1033;
input v_1034;
input v_1035;
input v_1036;
input v_1037;
input v_1038;
input v_1039;
input v_1040;
input v_1041;
input v_1042;
input v_1043;
input v_1044;
input v_1045;
input v_1046;
input v_1047;
input v_1048;
input v_1049;
input v_1050;
input v_1051;
input v_1052;
input v_1053;
input v_1054;
input v_1055;
input v_1056;
input v_1057;
input v_1058;
input v_1059;
input v_1060;
input v_1061;
input v_1062;
input v_1063;
input v_1064;
input v_1065;
input v_1066;
input v_1067;
input v_1068;
input v_1069;
input v_1070;
input v_1071;
input v_1072;
input v_1073;
input v_1074;
input v_1075;
input v_1076;
input v_1077;
input v_1078;
input v_1079;
input v_1080;
input v_1081;
input v_1082;
input v_1083;
input v_1084;
input v_1085;
input v_1086;
input v_1087;
input v_1088;
input v_1089;
input v_1090;
input v_1091;
input v_1092;
input v_1093;
input v_1094;
input v_1095;
input v_1096;
input v_1097;
input v_1098;
input v_1099;
input v_1100;
input v_1101;
input v_1102;
input v_1103;
input v_1104;
input v_1105;
input v_1106;
input v_1107;
input v_1108;
input v_1109;
input v_1110;
input v_1111;
input v_1157;
input v_1158;
input v_1159;
input v_1160;
input v_1161;
input v_1162;
input v_1163;
input v_1164;
input v_1165;
input v_1166;
input v_1167;
input v_1168;
input v_1169;
input v_1170;
input v_1171;
input v_1172;
input v_1173;
input v_1174;
input v_1175;
input v_1176;
input v_1177;
input v_1178;
input v_1179;
input v_1180;
input v_1181;
input v_1182;
input v_1183;
input v_1184;
input v_1185;
input v_1186;
input v_1187;
input v_1188;
input v_1189;
input v_1190;
input v_1191;
input v_1192;
input v_1193;
input v_1194;
input v_1195;
input v_1196;
input v_1197;
input v_1198;
input v_1199;
input v_1200;
input v_1201;
input v_1202;
input v_1203;
input v_1204;
input v_1205;
input v_1206;
input v_1207;
input v_1208;
input v_1209;
input v_1210;
input v_1211;
input v_1212;
input v_1213;
input v_1214;
input v_1215;
input v_1216;
input v_1217;
input v_1218;
input v_1219;
input v_1220;
input v_1221;
input v_1222;
input v_1223;
input v_1224;
input v_1225;
input v_1226;
input v_1227;
input v_1228;
input v_1229;
input v_1230;
input v_1231;
input v_1232;
input v_1233;
input v_1234;
input v_1235;
input v_1236;
input v_1237;
input v_1238;
input v_1239;
input v_1240;
input v_1241;
input v_1242;
input v_1243;
input v_1244;
input v_1245;
input v_1246;
input v_1247;
input v_1248;
input v_1249;
input v_1250;
input v_1251;
input v_1252;
input v_1253;
input v_1254;
input v_1255;
input v_1256;
input v_1257;
input v_1258;
input v_1259;
input v_1260;
input v_1261;
input v_1262;
input v_1263;
input v_1264;
input v_1265;
input v_1266;
input v_1267;
input v_1268;
input v_1269;
input v_1270;
input v_1271;
input v_1272;
input v_1273;
input v_1274;
input v_1275;
input v_1276;
input v_1277;
input v_1278;
input v_1279;
input v_1280;
input v_1281;
input v_1282;
input v_1283;
input v_1284;
input v_1285;
input v_1286;
input v_1287;
input v_1288;
input v_1289;
input v_1290;
input v_1291;
input v_1292;
input v_1293;
input v_1294;
input v_1295;
input v_1296;
input v_1297;
input v_1298;
input v_1299;
input v_1300;
input v_1301;
input v_1302;
input v_1303;
input v_1304;
input v_1305;
input v_1306;
input v_1307;
input v_1308;
input v_1309;
input v_1310;
input v_1311;
input v_1312;
input v_1313;
input v_1314;
input v_1315;
input v_1316;
input v_1317;
input v_1318;
input v_1319;
input v_1320;
input v_1321;
input v_1322;
input v_1323;
input v_1324;
input v_1325;
input v_1326;
input v_1327;
input v_1328;
input v_1329;
input v_1330;
input v_1331;
input v_1332;
input v_1333;
input v_1334;
input v_1335;
input v_1336;
input v_1337;
input v_1383;
input v_1384;
input v_1385;
input v_1386;
input v_1387;
input v_1388;
input v_1389;
input v_1390;
input v_1391;
input v_1392;
input v_1393;
input v_1394;
input v_1395;
input v_1396;
input v_1397;
input v_1398;
input v_1399;
input v_1400;
input v_1401;
input v_1402;
input v_1403;
input v_1404;
input v_1405;
input v_1406;
input v_1407;
input v_1408;
input v_1409;
input v_1410;
input v_1411;
input v_1412;
input v_1413;
input v_1414;
input v_1415;
input v_1416;
input v_1417;
input v_1418;
input v_1419;
input v_1420;
input v_1421;
input v_1422;
input v_1423;
input v_1424;
input v_1425;
input v_1426;
input v_1427;
input v_1428;
input v_1429;
input v_1430;
input v_1431;
input v_1432;
input v_1433;
input v_1434;
input v_1435;
input v_1436;
input v_1437;
input v_1438;
input v_1439;
input v_1440;
input v_1441;
input v_1442;
input v_1443;
input v_1444;
input v_1445;
input v_1446;
input v_1447;
input v_1448;
input v_1449;
input v_1450;
input v_1451;
input v_1452;
input v_1453;
input v_1454;
input v_1455;
input v_1456;
input v_1457;
input v_1458;
input v_1459;
input v_1460;
input v_1461;
input v_1462;
input v_1463;
input v_1464;
input v_1465;
input v_1466;
input v_1467;
input v_1468;
input v_1469;
input v_1470;
input v_1471;
input v_1472;
input v_1473;
input v_1474;
input v_1475;
input v_1476;
input v_1477;
input v_1478;
input v_1479;
input v_1480;
input v_1481;
input v_1482;
input v_1483;
input v_1484;
input v_1485;
input v_1486;
input v_1487;
input v_1488;
input v_1489;
input v_1490;
input v_1491;
input v_1492;
input v_1493;
input v_1494;
input v_1495;
input v_1496;
input v_1497;
input v_1498;
input v_1499;
input v_1500;
input v_1501;
input v_1502;
input v_1503;
input v_1504;
input v_1505;
input v_1506;
input v_1507;
input v_1508;
input v_1509;
input v_1510;
input v_1511;
input v_1512;
input v_1513;
input v_1514;
input v_1515;
input v_1516;
input v_1517;
input v_1518;
input v_1519;
input v_1520;
input v_1521;
input v_1522;
input v_1523;
input v_1524;
input v_1525;
input v_1526;
input v_1527;
input v_1528;
input v_1529;
input v_1530;
input v_1531;
input v_1532;
input v_1533;
input v_1534;
input v_1535;
input v_1536;
input v_1537;
input v_1538;
input v_1539;
input v_1540;
input v_1541;
input v_1542;
input v_1543;
input v_1544;
input v_1545;
input v_1546;
input v_1547;
input v_1548;
input v_1549;
input v_1550;
input v_1551;
input v_1552;
input v_1553;
input v_1554;
input v_1555;
input v_1556;
input v_1557;
input v_1558;
input v_1559;
input v_1560;
input v_1561;
input v_1562;
input v_1563;
input v_1564;
input v_1565;
input v_1566;
input v_1567;
input v_1568;
input v_1569;
input v_1570;
input v_1571;
input v_1572;
input v_1573;
input v_1574;
input v_1575;
input v_1576;
input v_1577;
input v_1578;
input v_1579;
input v_1580;
input v_1581;
input v_1582;
input v_1583;
input v_1584;
input v_1585;
input v_1586;
input v_1587;
input v_1588;
input v_1589;
input v_1590;
input v_1591;
input v_1592;
input v_1593;
input v_1594;
input v_1595;
input v_1596;
input v_1597;
input v_1598;
input v_1599;
input v_1600;
input v_1601;
input v_1602;
input v_1603;
input v_1604;
input v_1605;
input v_1606;
input v_1607;
input v_1608;
input v_1609;
input v_1610;
input v_1611;
input v_1612;
input v_1613;
input v_1614;
input v_1615;
input v_1616;
input v_1617;
input v_1618;
input v_1619;
input v_1620;
input v_1621;
input v_1622;
input v_1623;
input v_1624;
input v_1625;
input v_1626;
input v_1627;
input v_1628;
input v_1629;
input v_1630;
input v_1631;
input v_1632;
input v_1633;
input v_1634;
input v_1635;
input v_1636;
input v_1637;
input v_1638;
input v_1639;
input v_1640;
input v_1641;
input v_1642;
input v_1643;
input v_1644;
input v_1645;
input v_1646;
input v_1647;
input v_1648;
input v_1649;
input v_1650;
input v_1651;
input v_1652;
input v_1653;
input v_1654;
input v_1655;
input v_1656;
input v_1657;
input v_1658;
input v_1659;
input v_1660;
input v_1661;
input v_1662;
input v_1663;
input v_1664;
input v_1665;
input v_1666;
input v_1667;
input v_1668;
input v_1669;
input v_1670;
input v_1671;
input v_1672;
input v_1673;
input v_1674;
input v_1675;
input v_1676;
input v_1677;
input v_1678;
input v_1679;
input v_1680;
input v_1681;
input v_1682;
input v_1683;
input v_1684;
input v_1685;
input v_1686;
input v_1687;
input v_1688;
input v_1689;
input v_1690;
input v_1691;
input v_1692;
input v_1693;
input v_1694;
input v_1695;
input v_1696;
input v_1697;
input v_1698;
input v_1699;
input v_1700;
input v_1701;
input v_1702;
input v_1703;
input v_1704;
input v_1705;
input v_1706;
input v_1707;
input v_1708;
input v_1709;
input v_1710;
input v_1711;
input v_1712;
input v_1713;
input v_1714;
input v_1715;
input v_1716;
input v_1717;
input v_1718;
input v_1719;
input v_1720;
input v_1721;
input v_1722;
input v_1723;
input v_1724;
input v_1725;
input v_1726;
input v_1727;
input v_1728;
input v_1729;
input v_1730;
input v_1731;
input v_1732;
input v_1733;
input v_1734;
input v_1735;
input v_1736;
input v_1737;
input v_1738;
input v_1739;
input v_1740;
input v_1741;
input v_1742;
input v_1743;
input v_1744;
input v_1745;
input v_1746;
input v_1747;
input v_1748;
input v_1749;
input v_1750;
input v_1751;
input v_1752;
input v_1753;
input v_1754;
input v_1755;
input v_1756;
input v_1757;
input v_1758;
input v_1759;
input v_1760;
input v_1761;
input v_1762;
input v_1763;
input v_1764;
input v_1765;
input v_1766;
input v_1767;
input v_1768;
input v_1769;
input v_1770;
input v_1771;
input v_1772;
input v_1773;
input v_1774;
input v_1775;
input v_1776;
input v_1777;
input v_1778;
input v_1779;
input v_1780;
input v_1781;
input v_1782;
input v_1783;
input v_1784;
input v_1785;
input v_1786;
input v_1787;
input v_1788;
input v_1789;
input v_1790;
input v_1791;
input v_1792;
input v_1793;
input v_1794;
input v_1795;
input v_1796;
input v_1797;
input v_1798;
input v_1799;
input v_1800;
input v_1801;
input v_1802;
input v_1803;
input v_1804;
input v_1805;
input v_1806;
input v_1807;
input v_1808;
input v_1809;
input v_1810;
input v_1811;
input v_1812;
input v_1813;
input v_1814;
input v_1815;
input v_1816;
input v_1817;
input v_1818;
input v_1819;
input v_1820;
input v_1821;
input v_1822;
input v_1823;
input v_1824;
input v_1825;
input v_1826;
input v_1827;
input v_1828;
input v_1829;
input v_1830;
input v_1831;
input v_1832;
input v_1833;
input v_1834;
input v_1835;
input v_1836;
input v_1837;
input v_1838;
input v_1839;
input v_1840;
input v_1841;
input v_1842;
input v_1843;
input v_1844;
input v_1845;
input v_1846;
input v_1847;
input v_1848;
input v_1849;
input v_1850;
input v_1851;
input v_1852;
input v_1853;
input v_1854;
input v_1855;
input v_1856;
input v_1857;
input v_1858;
input v_1859;
input v_1860;
input v_1861;
input v_1862;
input v_1863;
input v_1864;
input v_1865;
input v_1866;
input v_1867;
input v_1868;
input v_1869;
input v_1870;
input v_1871;
input v_1872;
input v_1873;
input v_1874;
input v_1875;
input v_1876;
input v_1877;
input v_1878;
input v_1879;
input v_1880;
input v_1881;
input v_1882;
input v_1883;
input v_1884;
input v_1885;
input v_1886;
input v_1887;
input v_1888;
input v_1889;
input v_1890;
input v_1891;
input v_1892;
input v_1893;
input v_1894;
input v_1895;
input v_1896;
input v_1897;
input v_1898;
input v_1899;
input v_1900;
input v_1901;
input v_1902;
input v_1903;
input v_1904;
input v_1905;
input v_1906;
input v_1907;
input v_1908;
input v_1909;
input v_1910;
input v_1911;
input v_1912;
input v_1913;
input v_1914;
input v_1915;
input v_1916;
input v_1917;
input v_1918;
input v_1919;
input v_1920;
input v_1921;
input v_1922;
input v_1923;
input v_1924;
input v_1925;
input v_1926;
input v_1927;
input v_1928;
input v_1929;
input v_1930;
input v_1931;
input v_1932;
input v_1933;
input v_1934;
input v_1935;
input v_1936;
input v_1937;
input v_1938;
input v_1939;
input v_1940;
input v_1941;
input v_1942;
input v_1943;
input v_1944;
input v_1945;
input v_1946;
input v_1947;
input v_1948;
input v_1949;
input v_1950;
input v_1951;
input v_1952;
input v_1953;
input v_1954;
input v_1955;
input v_1956;
input v_1957;
input v_1958;
input v_1959;
input v_1960;
input v_1961;
input v_1962;
input v_1963;
input v_1964;
input v_1965;
input v_1966;
input v_1967;
input v_1968;
input v_1969;
input v_1970;
input v_1971;
input v_1972;
input v_1973;
input v_1974;
input v_1975;
input v_1976;
input v_1977;
input v_1978;
input v_1979;
input v_1980;
input v_1981;
input v_1982;
input v_1983;
input v_1984;
input v_1985;
input v_1986;
input v_1987;
input v_1988;
input v_1989;
input v_1990;
input v_1991;
input v_1992;
input v_1993;
input v_1994;
input v_1995;
input v_1996;
input v_1997;
input v_1998;
input v_1999;
input v_2000;
input v_2001;
input v_2002;
input v_2003;
input v_2004;
input v_2005;
input v_2006;
input v_2007;
input v_2008;
input v_2009;
input v_2010;
input v_2011;
input v_2012;
input v_2013;
input v_2014;
input v_2015;
input v_2016;
input v_2017;
input v_2018;
input v_2019;
input v_2020;
input v_2021;
input v_2022;
input v_2023;
input v_2024;
input v_2025;
input v_2026;
input v_2027;
input v_2028;
input v_2029;
input v_2030;
input v_2031;
input v_2032;
input v_2033;
input v_2034;
input v_2035;
input v_2036;
input v_2037;
input v_2038;
input v_2039;
input v_2040;
input v_2041;
input v_2042;
input v_2043;
input v_2044;
input v_2045;
input v_2046;
input v_2047;
input v_2048;
input v_2049;
input v_2050;
input v_2051;
input v_2052;
input v_2053;
input v_2054;
input v_2055;
input v_2056;
input v_2057;
input v_2058;
input v_2059;
input v_2060;
input v_2061;
input v_2062;
input v_2063;
input v_2064;
input v_2065;
input v_2066;
input v_2067;
input v_2068;
input v_2069;
input v_2070;
input v_2071;
input v_2072;
input v_2073;
input v_2074;
input v_2075;
input v_2076;
input v_2077;
input v_2078;
input v_2079;
input v_2080;
input v_2081;
input v_2082;
input v_2083;
input v_2084;
input v_2085;
input v_2086;
input v_2087;
input v_2088;
input v_2089;
input v_2090;
input v_2091;
input v_2092;
input v_2093;
input v_2094;
input v_2095;
input v_2096;
input v_2097;
input v_2098;
input v_2099;
input v_2100;
input v_2101;
input v_2102;
input v_2103;
input v_2104;
input v_2105;
input v_2106;
input v_2107;
input v_2108;
input v_2109;
input v_2110;
input v_2111;
input v_2112;
input v_2113;
input v_2114;
input v_2115;
input v_2116;
input v_2117;
input v_2118;
input v_2119;
input v_2120;
input v_2121;
input v_2122;
input v_2123;
input v_2124;
input v_2125;
input v_2126;
input v_2127;
input v_2128;
input v_2129;
input v_2130;
input v_2131;
input v_2132;
input v_2133;
input v_2134;
input v_2135;
input v_2136;
input v_2137;
input v_2138;
input v_2139;
input v_2140;
input v_2141;
input v_2142;
input v_2143;
input v_2144;
input v_2145;
input v_2146;
input v_2147;
input v_2148;
input v_2149;
input v_2150;
input v_2151;
input v_2152;
input v_2153;
input v_2154;
input v_2155;
input v_2156;
input v_2157;
input v_2158;
input v_2159;
input v_2160;
input v_2161;
input v_2162;
input v_2163;
input v_2164;
input v_2165;
input v_2166;
input v_2167;
input v_2168;
input v_2169;
input v_2170;
input v_2171;
input v_2172;
input v_2173;
input v_2174;
input v_2175;
input v_2176;
input v_2177;
input v_2178;
input v_2179;
input v_2180;
input v_2181;
input v_2182;
input v_2183;
input v_2184;
input v_2185;
input v_2186;
input v_2187;
input v_2188;
input v_2189;
input v_2190;
input v_2191;
input v_2192;
input v_2193;
input v_2194;
input v_2195;
input v_2196;
input v_2197;
input v_2198;
input v_2199;
input v_2200;
input v_2201;
input v_2202;
input v_2203;
input v_2204;
input v_2205;
input v_2206;
input v_2207;
input v_2208;
input v_2209;
input v_2210;
input v_2211;
input v_2212;
input v_2213;
input v_2214;
input v_2215;
input v_2216;
input v_2217;
input v_2218;
input v_2219;
input v_2220;
input v_2221;
input v_2222;
input v_2223;
input v_2224;
input v_2225;
input v_2226;
input v_2227;
input v_2228;
input v_2229;
input v_2230;
input v_2231;
input v_2232;
input v_2233;
input v_2234;
input v_2235;
input v_2236;
input v_2237;
input v_2238;
input v_2239;
input v_2240;
input v_2241;
input v_2242;
input v_2243;
input v_2244;
input v_2245;
input v_2246;
input v_2247;
input v_2248;
input v_2249;
input v_2250;
input v_2251;
input v_2252;
input v_2253;
input v_2254;
input v_2255;
input v_2256;
input v_2257;
input v_2258;
input v_2259;
input v_2260;
input v_2261;
input v_2262;
input v_2263;
input v_2264;
input v_2265;
input v_2266;
input v_2267;
input v_2268;
input v_2269;
input v_2270;
input v_2271;
input v_2272;
input v_2273;
input v_2274;
input v_2275;
input v_2276;
input v_2277;
input v_2278;
input v_2279;
input v_2280;
input v_2281;
input v_2282;
input v_2283;
input v_2284;
input v_2285;
input v_2286;
input v_2287;
input v_2288;
input v_2289;
input v_2290;
input v_2291;
input v_2292;
input v_2293;
input v_2294;
input v_2295;
input v_2296;
input v_2297;
input v_2298;
input v_2299;
input v_2300;
input v_2301;
input v_2302;
input v_2303;
input v_2304;
input v_2305;
input v_2306;
input v_2307;
input v_2308;
input v_2309;
input v_2310;
input v_2311;
input v_2312;
input v_2313;
input v_2314;
input v_2315;
input v_2316;
input v_2317;
input v_2318;
input v_2319;
input v_2320;
input v_2321;
input v_2322;
input v_2323;
input v_2324;
input v_2325;
input v_2326;
input v_2327;
input v_2328;
input v_2329;
input v_2330;
input v_2331;
input v_2332;
input v_2333;
input v_2334;
input v_2335;
input v_2336;
input v_2337;
input v_2338;
input v_2339;
input v_2340;
input v_2341;
input v_2342;
input v_2343;
input v_2344;
input v_2345;
input v_2346;
input v_2347;
input v_2348;
input v_2349;
input v_2350;
input v_2351;
input v_2352;
input v_2353;
input v_2354;
input v_2355;
input v_2356;
input v_2357;
input v_2358;
input v_2359;
input v_2360;
input v_2361;
input v_2362;
input v_2363;
input v_2364;
input v_2365;
input v_2366;
input v_2367;
input v_2368;
input v_2369;
input v_2370;
input v_2371;
input v_2372;
input v_2373;
input v_2374;
input v_2375;
input v_2376;
input v_2377;
input v_2378;
input v_2379;
input v_2380;
input v_2381;
input v_2382;
input v_2383;
input v_2384;
input v_2385;
input v_2386;
input v_2387;
input v_2388;
input v_2389;
input v_2390;
input v_2391;
input v_2392;
input v_2393;
input v_2394;
input v_2395;
input v_2396;
input v_2397;
input v_2398;
input v_2399;
input v_2400;
input v_2401;
input v_2402;
input v_2403;
input v_2404;
input v_2405;
input v_2406;
input v_2407;
input v_2408;
input v_2409;
input v_2410;
input v_2411;
input v_2412;
input v_2413;
input v_2414;
input v_2415;
input v_2416;
input v_2417;
input v_2418;
input v_2419;
input v_2420;
input v_2421;
input v_2422;
input v_2423;
input v_2424;
input v_2425;
input v_2426;
input v_2427;
input v_2428;
input v_2429;
input v_2430;
input v_2431;
input v_2432;
input v_2433;
input v_2434;
input v_2435;
input v_2436;
input v_2437;
input v_2438;
input v_2439;
input v_2440;
input v_2441;
input v_2442;
input v_2443;
input v_2444;
input v_2445;
input v_2446;
input v_2447;
input v_2448;
input v_2449;
input v_2450;
input v_2451;
input v_2452;
input v_2453;
input v_2454;
input v_2455;
input v_2456;
input v_2457;
input v_2458;
input v_2459;
input v_2460;
input v_2461;
input v_2462;
input v_2463;
input v_2464;
input v_2465;
input v_2466;
input v_2467;
input v_2468;
input v_2469;
input v_2470;
input v_2471;
input v_2472;
input v_2473;
input v_2474;
input v_2475;
input v_2476;
input v_2477;
input v_2478;
input v_2479;
input v_2480;
input v_2481;
input v_2482;
input v_2483;
input v_2484;
input v_2485;
input v_2486;
input v_2487;
input v_2488;
input v_2489;
input v_2490;
input v_2491;
input v_2492;
input v_2493;
input v_2494;
input v_2495;
input v_2496;
input v_2497;
input v_2498;
input v_2499;
input v_2500;
input v_2501;
input v_2502;
input v_2503;
input v_2504;
input v_2505;
input v_2506;
input v_2507;
input v_2508;
input v_2509;
input v_2510;
input v_2511;
input v_2512;
input v_2513;
input v_2514;
input v_2515;
input v_2516;
input v_2517;
input v_2518;
input v_2519;
input v_2520;
input v_2521;
input v_2522;
input v_2523;
input v_2524;
input v_2525;
input v_2526;
input v_2527;
input v_2528;
input v_2529;
input v_2530;
input v_2531;
input v_2532;
input v_2533;
input v_2534;
input v_2535;
input v_2536;
input v_2537;
input v_2538;
input v_2539;
input v_2540;
input v_2541;
input v_2542;
input v_2543;
input v_2544;
input v_2545;
input v_2546;
input v_2547;
input v_2548;
input v_2549;
input v_2550;
input v_2551;
input v_2552;
input v_2553;
input v_2554;
input v_2555;
input v_2556;
input v_2557;
input v_2558;
input v_2559;
input v_2560;
input v_2561;
input v_2562;
input v_2563;
input v_2564;
input v_2565;
input v_2566;
input v_2567;
input v_2568;
input v_2569;
input v_2570;
input v_2571;
input v_2572;
input v_2573;
input v_2574;
input v_2575;
input v_2576;
input v_2577;
input v_2578;
input v_2579;
input v_2580;
input v_2581;
input v_2582;
input v_2583;
input v_2584;
input v_2585;
input v_2586;
input v_2587;
input v_2588;
input v_2589;
input v_2590;
input v_2591;
input v_2592;
input v_2593;
input v_2594;
input v_2595;
input v_2596;
input v_2597;
input v_2598;
input v_2599;
input v_2600;
input v_2601;
input v_2602;
input v_2603;
input v_2604;
input v_2605;
input v_2606;
input v_2607;
input v_2608;
input v_2609;
input v_2610;
input v_2611;
input v_2612;
input v_2613;
input v_2614;
input v_2615;
input v_2616;
input v_2617;
input v_2618;
input v_2619;
input v_2620;
input v_2621;
input v_2622;
input v_2623;
input v_2624;
input v_2625;
input v_2626;
input v_2627;
input v_2628;
input v_2629;
input v_2630;
input v_2631;
input v_2632;
input v_2633;
input v_2634;
input v_2635;
input v_2636;
input v_2637;
input v_2638;
input v_2639;
input v_2640;
input v_2641;
input v_2642;
input v_2643;
input v_2644;
input v_2645;
input v_2646;
input v_2647;
input v_2648;
input v_2649;
input v_2650;
input v_2651;
input v_2652;
input v_2653;
input v_2654;
input v_2655;
input v_2656;
input v_2657;
input v_2658;
input v_2659;
input v_2660;
input v_2661;
input v_2662;
input v_2663;
input v_2664;
input v_2665;
input v_2666;
input v_2667;
input v_2668;
input v_2669;
input v_2670;
input v_2671;
input v_2672;
input v_2673;
input v_2674;
input v_2675;
input v_2676;
input v_2677;
input v_2678;
input v_2679;
input v_2680;
input v_2681;
input v_2682;
input v_2683;
input v_2684;
input v_2685;
input v_2686;
input v_2687;
input v_2688;
input v_2689;
input v_2690;
input v_2691;
input v_2692;
input v_2693;
input v_2694;
input v_2695;
input v_2696;
input v_2697;
input v_2698;
input v_2699;
input v_2700;
input v_2701;
input v_2702;
input v_2703;
input v_2704;
input v_2705;
input v_2706;
input v_2707;
input v_2708;
input v_2709;
input v_2710;
input v_2711;
input v_2712;
input v_2713;
input v_2714;
input v_2715;
input v_2716;
input v_2717;
input v_2718;
input v_2719;
input v_2720;
input v_2721;
input v_2722;
input v_2723;
input v_2724;
input v_2725;
input v_2726;
input v_2727;
input v_2728;
input v_2729;
input v_2730;
input v_2731;
input v_2732;
input v_2733;
input v_2734;
input v_2735;
input v_2736;
input v_2737;
input v_2738;
input v_2739;
input v_2740;
input v_2741;
input v_2742;
input v_2743;
input v_2744;
input v_2745;
input v_2746;
input v_2747;
input v_2748;
input v_2749;
input v_2750;
input v_2751;
input v_2752;
input v_2753;
input v_2754;
input v_2755;
input v_2756;
input v_2757;
input v_2758;
input v_2759;
input v_2760;
input v_2761;
input v_2762;
input v_2763;
input v_2764;
input v_2765;
input v_2766;
input v_2767;
input v_2768;
input v_2769;
input v_2770;
input v_2771;
input v_2772;
input v_2773;
input v_2774;
input v_2775;
input v_2776;
input v_2777;
input v_2778;
input v_2779;
input v_2780;
input v_2781;
input v_2782;
input v_2783;
input v_2784;
input v_2785;
input v_2786;
input v_2787;
input v_2788;
input v_2789;
input v_2790;
input v_2791;
input v_2792;
input v_2793;
input v_2794;
input v_2795;
input v_2796;
input v_2797;
input v_2798;
input v_2799;
input v_2800;
input v_2801;
input v_2802;
input v_2803;
input v_2804;
input v_2805;
input v_2806;
input v_2807;
input v_2808;
input v_2809;
input v_2810;
input v_2811;
input v_2812;
input v_2813;
input v_2814;
input v_2815;
input v_2816;
input v_2817;
input v_2818;
input v_2819;
input v_2820;
input v_2821;
input v_2822;
input v_2823;
input v_2824;
input v_2825;
input v_2826;
input v_2827;
input v_2828;
input v_2829;
input v_2830;
input v_2831;
input v_2832;
input v_2833;
input v_2834;
input v_2835;
input v_2836;
input v_2837;
input v_2838;
input v_2839;
input v_2840;
input v_2841;
input v_2842;
input v_2843;
input v_2844;
input v_2845;
input v_2846;
input v_2847;
input v_2848;
input v_2849;
input v_2850;
input v_2851;
input v_2852;
input v_2853;
input v_2854;
input v_2855;
input v_2856;
input v_2857;
input v_2858;
input v_2859;
input v_2860;
input v_2861;
input v_2862;
input v_2863;
input v_2864;
input v_2865;
input v_2866;
input v_2867;
input v_2868;
input v_2869;
input v_2870;
input v_2871;
input v_2872;
input v_2873;
input v_2874;
input v_2875;
input v_2876;
input v_2877;
input v_2878;
input v_2879;
input v_2880;
input v_2881;
input v_2882;
input v_2883;
input v_2884;
input v_2885;
input v_2886;
input v_2887;
input v_2888;
input v_2889;
input v_2890;
input v_2891;
input v_2892;
input v_2893;
input v_2894;
input v_2895;
input v_2896;
input v_2897;
input v_2898;
input v_2899;
input v_2900;
input v_2901;
input v_2902;
input v_2903;
input v_2904;
input v_2905;
input v_2906;
input v_2907;
input v_2908;
input v_2909;
input v_2910;
input v_2911;
input v_2912;
input v_2913;
input v_2914;
input v_2915;
input v_2916;
input v_2917;
input v_2918;
input v_2919;
input v_2920;
input v_2921;
input v_2922;
input v_2923;
input v_2924;
input v_2925;
input v_2926;
input v_2927;
input v_2928;
input v_2929;
input v_2930;
input v_2931;
input v_2932;
input v_2933;
input v_2934;
input v_2935;
input v_2936;
input v_2937;
input v_2938;
input v_2939;
input v_2940;
input v_2941;
input v_2942;
input v_2943;
input v_2944;
input v_2945;
input v_2946;
input v_2947;
input v_2948;
input v_2949;
input v_2950;
input v_2951;
input v_2952;
input v_2953;
input v_2954;
input v_2955;
input v_2956;
input v_2957;
input v_2958;
input v_2959;
input v_2960;
input v_2961;
input v_2962;
input v_2963;
input v_2964;
input v_2965;
input v_2966;
input v_2967;
input v_2968;
input v_2969;
input v_2970;
input v_2971;
input v_2972;
input v_2973;
input v_2974;
input v_2975;
input v_2976;
input v_2977;
input v_2978;
input v_2979;
input v_2980;
input v_2981;
input v_2982;
input v_2983;
input v_2984;
input v_2985;
input v_2986;
input v_2987;
input v_2988;
input v_2989;
input v_2990;
input v_2991;
input v_2992;
input v_2993;
input v_2994;
input v_2995;
input v_2996;
input v_2997;
input v_2998;
input v_2999;
input v_3000;
input v_3001;
input v_3002;
input v_3003;
input v_3004;
input v_3005;
input v_3006;
input v_3007;
input v_3008;
input v_3009;
input v_3010;
input v_3011;
input v_3012;
input v_3013;
input v_3014;
input v_3015;
input v_3016;
input v_3017;
input v_3018;
input v_3019;
input v_3020;
input v_3021;
input v_3022;
input v_3023;
input v_3024;
input v_3025;
input v_3026;
input v_3027;
input v_3028;
input v_3029;
input v_3030;
input v_3031;
input v_3032;
input v_3033;
input v_3034;
input v_3035;
input v_3036;
input v_3037;
input v_3038;
input v_3039;
input v_3040;
input v_3041;
input v_3042;
input v_3043;
input v_3044;
input v_3045;
input v_3046;
input v_3047;
input v_3048;
input v_3049;
input v_3050;
input v_3051;
input v_3052;
input v_3053;
input v_3054;
input v_3055;
input v_3056;
input v_3057;
input v_3058;
input v_3059;
input v_3060;
input v_3061;
input v_3062;
input v_3063;
input v_3064;
input v_3065;
input v_3066;
input v_3067;
input v_3068;
input v_3069;
input v_3070;
input v_3071;
input v_3072;
input v_3073;
input v_3074;
input v_3075;
input v_3076;
input v_3077;
input v_3078;
input v_3079;
input v_3080;
input v_3081;
input v_3082;
input v_3083;
input v_3084;
input v_3085;
input v_3086;
input v_3087;
input v_3088;
input v_3089;
input v_3090;
input v_3091;
input v_3092;
input v_3093;
input v_3094;
input v_3095;
input v_3096;
input v_3097;
input v_3098;
input v_3099;
input v_3100;
input v_3101;
input v_3102;
input v_3103;
input v_3104;
input v_3105;
input v_3106;
input v_3107;
input v_3108;
input v_3109;
input v_3110;
input v_3111;
input v_3112;
input v_3113;
input v_3114;
input v_3115;
input v_3116;
input v_3117;
input v_3118;
input v_3119;
input v_3120;
input v_3121;
input v_3122;
input v_3123;
input v_3124;
input v_3125;
input v_3126;
input v_3127;
input v_3128;
input v_3129;
input v_3130;
input v_3131;
input v_3132;
input v_3133;
input v_3134;
input v_3135;
input v_3136;
input v_3137;
input v_3138;
input v_3139;
input v_3140;
input v_3141;
input v_3142;
input v_3143;
input v_3144;
input v_3145;
input v_3146;
input v_3147;
input v_3148;
input v_3149;
input v_3150;
input v_3151;
input v_3152;
input v_3153;
input v_3154;
input v_3155;
input v_3156;
input v_3157;
input v_3158;
input v_3159;
input v_3160;
input v_3161;
input v_3162;
input v_3163;
input v_3164;
input v_3165;
input v_3166;
input v_3167;
input v_3168;
input v_3169;
input v_3170;
input v_3171;
input v_3172;
input v_3173;
input v_3174;
input v_3175;
input v_3176;
input v_3177;
input v_3178;
input v_3179;
input v_3180;
input v_3181;
input v_3182;
input v_3183;
input v_3184;
input v_3185;
input v_3186;
input v_3187;
input v_3188;
input v_3189;
input v_3190;
input v_3191;
input v_3192;
input v_3193;
input v_3194;
input v_3195;
input v_3196;
input v_3197;
input v_3198;
input v_3199;
input v_3200;
input v_3201;
input v_3202;
input v_3203;
input v_3204;
input v_3205;
input v_3206;
input v_3207;
input v_3208;
input v_3209;
input v_3210;
input v_3211;
input v_3212;
input v_3213;
input v_3214;
input v_3215;
input v_3216;
input v_3217;
input v_3218;
input v_3219;
input v_3220;
input v_3221;
input v_3222;
input v_3223;
input v_3224;
input v_3225;
input v_3226;
input v_3227;
input v_3228;
input v_3229;
input v_3230;
input v_3231;
input v_3232;
input v_3233;
input v_3234;
input v_3235;
input v_3236;
input v_3237;
input v_3238;
input v_3239;
input v_3240;
input v_3241;
input v_3242;
input v_3243;
input v_3244;
input v_3245;
input v_3246;
input v_3247;
input v_3248;
input v_3249;
input v_3250;
input v_3251;
input v_3252;
input v_3253;
input v_3254;
input v_3255;
input v_3256;
input v_3257;
input v_3258;
input v_3259;
input v_3260;
input v_3261;
input v_3262;
input v_3263;
input v_3264;
input v_3265;
input v_3266;
input v_3267;
input v_3268;
input v_3269;
input v_3270;
input v_3271;
input v_3272;
input v_3273;
input v_3274;
input v_3275;
input v_3276;
input v_3277;
input v_3278;
input v_3279;
input v_3280;
input v_3281;
input v_3282;
input v_3283;
input v_3284;
input v_3285;
input v_3286;
input v_3287;
input v_3288;
input v_3289;
input v_3290;
input v_3291;
input v_3292;
input v_3293;
input v_3294;
input v_3295;
input v_3296;
input v_3297;
input v_3298;
input v_3299;
input v_3300;
input v_3301;
input v_3302;
input v_3303;
input v_3304;
input v_3305;
input v_3306;
input v_3307;
input v_3308;
input v_3309;
input v_3310;
input v_3311;
input v_3312;
input v_3313;
input v_3314;
input v_3315;
input v_3316;
input v_3317;
input v_3318;
input v_3319;
input v_3320;
input v_3321;
input v_3322;
input v_3323;
input v_3324;
input v_3325;
input v_3326;
input v_3327;
input v_3328;
input v_3329;
input v_3330;
input v_3331;
input v_3332;
input v_3333;
input v_3334;
input v_3335;
input v_3336;
input v_3337;
input v_3338;
input v_3339;
input v_3340;
input v_3341;
input v_3342;
input v_3343;
input v_3344;
input v_3345;
input v_3346;
input v_3347;
input v_3348;
input v_3349;
input v_3350;
input v_3351;
input v_3352;
input v_3353;
input v_3354;
input v_3355;
input v_3356;
input v_3357;
input v_3358;
input v_3359;
input v_3360;
input v_3361;
input v_3362;
input v_3363;
input v_3364;
input v_3365;
input v_3366;
input v_3367;
input v_3368;
input v_3369;
input v_3370;
input v_3371;
input v_3372;
input v_3373;
input v_3374;
input v_3375;
input v_3376;
input v_3377;
input v_3378;
input v_3379;
input v_3380;
input v_3381;
input v_3382;
input v_3383;
input v_3384;
input v_3385;
input v_3386;
input v_3387;
input v_3388;
input v_3389;
input v_3390;
input v_3391;
input v_3392;
input v_3393;
input v_3394;
input v_3395;
input v_3396;
input v_3397;
input v_3398;
input v_3399;
input v_3544;
input v_3545;
input v_3546;
input v_3547;
input v_3548;
input v_3549;
input v_3550;
input v_3551;
input v_3552;
input v_3553;
input v_3554;
input v_3555;
input v_3556;
input v_3557;
input v_3558;
input v_3559;
input v_3560;
input v_3561;
input v_3562;
input v_3563;
input v_3564;
input v_3565;
input v_3566;
input v_3567;
input v_3568;
input v_3569;
input v_3570;
input v_3571;
input v_3572;
input v_3573;
input v_3574;
input v_3575;
input v_3576;
input v_3577;
input v_3578;
input v_3579;
input v_3580;
input v_3581;
input v_3582;
input v_3583;
input v_3584;
input v_3585;
input v_3586;
input v_3587;
input v_3588;
input v_3589;
input v_3590;
input v_3591;
input v_3592;
input v_3593;
input v_3594;
input v_3595;
input v_3596;
input v_3597;
input v_3598;
input v_3599;
input v_3600;
input v_3601;
input v_3602;
input v_3603;
input v_3604;
input v_3605;
input v_3606;
input v_3607;
input v_3608;
input v_3609;
input v_3610;
input v_3611;
input v_3612;
input v_3613;
input v_3614;
input v_3615;
input v_3616;
input v_3617;
input v_3618;
input v_3619;
input v_3620;
input v_3621;
input v_3622;
input v_3623;
input v_3624;
input v_3625;
input v_3626;
input v_3627;
input v_3628;
input v_3629;
input v_3630;
input v_3631;
input v_3632;
input v_3633;
input v_3778;
input v_3779;
input v_3780;
input v_3781;
input v_3782;
input v_3783;
input v_3784;
input v_3785;
input v_3786;
input v_3787;
input v_3788;
input v_3789;
input v_3790;
input v_3791;
input v_3792;
input v_3793;
input v_3794;
input v_3795;
input v_3796;
input v_3797;
input v_3798;
input v_3799;
input v_3800;
input v_3801;
input v_3802;
input v_3803;
input v_3804;
input v_3805;
input v_3806;
input v_3807;
input v_3808;
input v_3809;
input v_3810;
input v_3811;
input v_3812;
input v_3813;
input v_3814;
input v_3815;
input v_3816;
input v_3817;
input v_3818;
input v_3819;
input v_3820;
input v_3821;
input v_3822;
input v_3823;
input v_3824;
input v_3825;
input v_3826;
input v_3827;
input v_3828;
input v_3829;
input v_3830;
input v_3831;
input v_3832;
input v_3833;
input v_3834;
input v_3835;
input v_3836;
input v_3837;
input v_3838;
input v_3839;
input v_3840;
input v_3841;
input v_3842;
input v_3843;
input v_3844;
input v_3845;
input v_3846;
input v_3847;
input v_3848;
input v_3849;
input v_3850;
input v_3851;
input v_3852;
input v_3853;
input v_3854;
input v_3855;
input v_3856;
input v_3857;
input v_3858;
input v_3859;
input v_3860;
input v_3861;
input v_3862;
input v_3863;
input v_3864;
input v_3865;
input v_3866;
input v_3867;
input v_4012;
input v_4013;
input v_4014;
input v_4015;
input v_4016;
input v_4017;
input v_4018;
input v_4019;
input v_4020;
input v_4021;
input v_4022;
input v_4023;
input v_4024;
input v_4025;
input v_4026;
input v_4027;
input v_4028;
input v_4029;
input v_4030;
input v_4031;
input v_4032;
input v_4033;
input v_4034;
input v_4035;
input v_4036;
input v_4037;
input v_4038;
input v_4039;
input v_4040;
input v_4041;
input v_4042;
input v_4043;
input v_4044;
input v_4045;
input v_4046;
input v_4047;
input v_4048;
input v_4049;
input v_4050;
input v_4051;
input v_4052;
input v_4053;
input v_4054;
input v_4055;
input v_4056;
input v_4057;
input v_4058;
input v_4059;
input v_4060;
input v_4061;
input v_4062;
input v_4063;
input v_4064;
input v_4065;
input v_4066;
input v_4067;
input v_4068;
input v_4069;
input v_4070;
input v_4071;
input v_4072;
input v_4073;
input v_4074;
input v_4075;
input v_4076;
input v_4077;
input v_4078;
input v_4079;
input v_4080;
input v_4081;
input v_4082;
input v_4083;
input v_4084;
input v_4085;
input v_4086;
input v_4087;
input v_4088;
input v_4089;
input v_4090;
input v_4091;
input v_4092;
input v_4093;
input v_4094;
input v_4095;
input v_4096;
input v_4097;
input v_4098;
input v_4099;
input v_4100;
input v_4101;
output o_1;
wire v_660;
wire v_661;
wire v_662;
wire v_663;
wire v_664;
wire v_665;
wire v_666;
wire v_667;
wire v_668;
wire v_669;
wire v_670;
wire v_671;
wire v_672;
wire v_673;
wire v_674;
wire v_675;
wire v_676;
wire v_677;
wire v_678;
wire v_679;
wire v_680;
wire v_681;
wire v_682;
wire v_683;
wire v_684;
wire v_685;
wire v_686;
wire v_687;
wire v_688;
wire v_689;
wire v_690;
wire v_691;
wire v_692;
wire v_693;
wire v_694;
wire v_695;
wire v_696;
wire v_697;
wire v_698;
wire v_699;
wire v_700;
wire v_701;
wire v_702;
wire v_703;
wire v_704;
wire v_886;
wire v_887;
wire v_888;
wire v_889;
wire v_890;
wire v_891;
wire v_892;
wire v_893;
wire v_894;
wire v_895;
wire v_896;
wire v_897;
wire v_898;
wire v_899;
wire v_900;
wire v_901;
wire v_902;
wire v_903;
wire v_904;
wire v_905;
wire v_906;
wire v_907;
wire v_908;
wire v_909;
wire v_910;
wire v_911;
wire v_912;
wire v_913;
wire v_914;
wire v_915;
wire v_916;
wire v_917;
wire v_918;
wire v_919;
wire v_920;
wire v_921;
wire v_922;
wire v_923;
wire v_924;
wire v_925;
wire v_926;
wire v_927;
wire v_928;
wire v_929;
wire v_930;
wire v_1112;
wire v_1113;
wire v_1114;
wire v_1115;
wire v_1116;
wire v_1117;
wire v_1118;
wire v_1119;
wire v_1120;
wire v_1121;
wire v_1122;
wire v_1123;
wire v_1124;
wire v_1125;
wire v_1126;
wire v_1127;
wire v_1128;
wire v_1129;
wire v_1130;
wire v_1131;
wire v_1132;
wire v_1133;
wire v_1134;
wire v_1135;
wire v_1136;
wire v_1137;
wire v_1138;
wire v_1139;
wire v_1140;
wire v_1141;
wire v_1142;
wire v_1143;
wire v_1144;
wire v_1145;
wire v_1146;
wire v_1147;
wire v_1148;
wire v_1149;
wire v_1150;
wire v_1151;
wire v_1152;
wire v_1153;
wire v_1154;
wire v_1155;
wire v_1156;
wire v_1338;
wire v_1339;
wire v_1340;
wire v_1341;
wire v_1342;
wire v_1343;
wire v_1344;
wire v_1345;
wire v_1346;
wire v_1347;
wire v_1348;
wire v_1349;
wire v_1350;
wire v_1351;
wire v_1352;
wire v_1353;
wire v_1354;
wire v_1355;
wire v_1356;
wire v_1357;
wire v_1358;
wire v_1359;
wire v_1360;
wire v_1361;
wire v_1362;
wire v_1363;
wire v_1364;
wire v_1365;
wire v_1366;
wire v_1367;
wire v_1368;
wire v_1369;
wire v_1370;
wire v_1371;
wire v_1372;
wire v_1373;
wire v_1374;
wire v_1375;
wire v_1376;
wire v_1377;
wire v_1378;
wire v_1379;
wire v_1380;
wire v_1381;
wire v_1382;
wire x_1;
wire x_2;
wire x_3;
wire x_4;
wire x_5;
wire x_6;
wire x_7;
wire x_8;
wire x_9;
wire x_10;
wire x_11;
wire x_12;
wire x_13;
wire x_14;
wire x_15;
wire x_16;
wire x_17;
wire x_18;
wire x_19;
wire x_20;
wire x_21;
wire x_22;
wire x_23;
wire x_24;
wire x_25;
wire x_26;
wire x_27;
wire x_28;
wire x_29;
wire x_30;
wire x_31;
wire x_32;
wire x_33;
wire x_34;
wire x_35;
wire x_36;
wire x_37;
wire x_38;
wire x_39;
wire x_40;
wire x_41;
wire x_42;
wire x_43;
wire x_44;
wire x_45;
wire x_46;
wire x_47;
wire x_48;
wire x_49;
wire x_50;
wire x_51;
wire x_52;
wire x_53;
wire x_54;
wire x_55;
wire x_56;
wire x_57;
wire x_58;
wire x_59;
wire x_60;
wire x_61;
wire x_62;
wire x_63;
wire x_64;
wire x_65;
wire x_66;
wire x_67;
wire x_68;
wire x_69;
wire x_70;
wire x_71;
wire x_72;
wire x_73;
wire x_74;
wire x_75;
wire x_76;
wire x_77;
wire x_78;
wire x_79;
wire x_80;
wire x_81;
wire x_82;
wire x_83;
wire x_84;
wire x_85;
wire x_86;
wire x_87;
wire x_88;
wire x_89;
wire x_90;
wire x_91;
wire x_92;
wire x_93;
wire x_94;
wire x_95;
wire x_96;
wire x_97;
wire x_98;
wire x_99;
wire x_100;
wire x_101;
wire x_102;
wire x_103;
wire x_104;
wire x_105;
wire x_106;
wire x_107;
wire x_108;
wire x_109;
wire x_110;
wire x_111;
wire x_112;
wire x_113;
wire x_114;
wire x_115;
wire x_116;
wire x_117;
wire x_118;
wire x_119;
wire x_120;
wire x_121;
wire x_122;
wire x_123;
wire x_124;
wire x_125;
wire x_126;
wire x_127;
wire x_128;
wire x_129;
wire x_130;
wire x_131;
wire x_132;
wire x_133;
wire x_134;
wire x_135;
wire x_136;
wire x_137;
wire x_138;
wire x_139;
wire x_140;
wire x_141;
wire x_142;
wire x_143;
wire x_144;
wire x_145;
wire x_146;
wire x_147;
wire x_148;
wire x_149;
wire x_150;
wire x_151;
wire x_152;
wire x_153;
wire x_154;
wire x_155;
wire x_156;
wire x_157;
wire x_158;
wire x_159;
wire x_160;
wire x_161;
wire x_162;
wire x_163;
wire x_164;
wire x_165;
wire x_166;
wire x_167;
wire x_168;
wire x_169;
wire x_170;
wire x_171;
wire x_172;
wire x_173;
wire x_174;
wire x_175;
wire x_176;
wire x_177;
wire x_178;
wire x_179;
wire x_180;
wire x_181;
wire x_182;
wire x_183;
wire x_184;
wire x_185;
wire x_186;
wire x_187;
wire x_188;
wire x_189;
wire x_190;
wire x_191;
wire x_192;
wire x_193;
wire x_194;
wire x_195;
wire x_196;
wire x_197;
wire x_198;
wire x_199;
wire x_200;
wire x_201;
wire x_202;
wire x_203;
wire x_204;
wire x_205;
wire x_206;
wire x_207;
wire x_208;
wire x_209;
wire x_210;
wire x_211;
wire x_212;
wire x_213;
wire x_214;
wire x_215;
wire x_216;
wire x_217;
wire x_218;
wire x_219;
wire x_220;
wire x_221;
wire x_222;
wire x_223;
wire x_224;
wire x_225;
wire x_226;
wire x_227;
wire x_228;
wire x_229;
wire x_230;
wire x_231;
wire x_232;
wire x_233;
wire x_234;
wire x_235;
wire x_236;
wire x_237;
wire x_238;
wire x_239;
wire x_240;
wire x_241;
wire x_242;
wire x_243;
wire x_244;
wire x_245;
wire x_246;
wire x_247;
wire x_248;
wire x_249;
wire x_250;
wire x_251;
wire x_252;
wire x_253;
wire x_254;
wire x_255;
wire x_256;
wire x_257;
wire x_258;
wire x_259;
wire x_260;
wire x_261;
wire x_262;
wire x_263;
wire x_264;
wire x_265;
wire x_266;
wire x_267;
wire x_268;
wire x_269;
wire x_270;
wire x_271;
wire x_272;
wire x_273;
wire x_274;
wire x_275;
wire x_276;
wire x_277;
wire x_278;
wire x_279;
wire x_280;
wire x_281;
wire x_282;
wire x_283;
wire x_284;
wire x_285;
wire x_286;
wire x_287;
wire x_288;
wire x_289;
wire x_290;
wire x_291;
wire x_292;
wire x_293;
wire x_294;
wire x_295;
wire x_296;
wire x_297;
wire x_298;
wire x_299;
wire x_300;
wire x_301;
wire x_302;
wire x_303;
wire x_304;
wire x_305;
wire x_306;
wire x_307;
wire x_308;
wire x_309;
wire x_310;
wire x_311;
wire x_312;
wire x_313;
wire x_314;
wire x_315;
wire x_316;
wire x_317;
wire x_318;
wire x_319;
wire x_320;
wire x_321;
wire x_322;
wire x_323;
wire x_324;
wire x_325;
wire x_326;
wire x_327;
wire x_328;
wire x_329;
wire x_330;
wire x_331;
wire x_332;
wire x_333;
wire x_334;
wire x_335;
wire x_336;
wire x_337;
wire x_338;
wire x_339;
wire x_340;
wire x_341;
wire x_342;
wire x_343;
wire x_344;
wire x_345;
wire x_346;
wire x_347;
wire x_348;
wire x_349;
wire x_350;
wire x_351;
wire x_352;
wire x_353;
wire x_354;
wire x_355;
wire x_356;
wire x_357;
wire x_358;
wire x_359;
wire x_360;
wire x_361;
wire x_362;
wire x_363;
wire x_364;
wire x_365;
wire x_366;
wire x_367;
wire x_368;
wire x_369;
wire x_370;
wire x_371;
wire x_372;
wire x_373;
wire x_374;
wire x_375;
wire x_376;
wire x_377;
wire x_378;
wire x_379;
wire x_380;
wire x_381;
wire x_382;
wire x_383;
wire x_384;
wire x_385;
wire x_386;
wire x_387;
wire x_388;
wire x_389;
wire x_390;
wire x_391;
wire x_392;
wire x_393;
wire x_394;
wire x_395;
wire x_396;
wire x_397;
wire x_398;
wire x_399;
wire x_400;
wire x_401;
wire x_402;
wire x_403;
wire x_404;
wire x_405;
wire x_406;
wire x_407;
wire x_408;
wire x_409;
wire x_410;
wire x_411;
wire x_412;
wire x_413;
wire x_414;
wire x_415;
wire x_416;
wire x_417;
wire x_418;
wire x_419;
wire x_420;
wire x_421;
wire x_422;
wire x_423;
wire x_424;
wire x_425;
wire x_426;
wire x_427;
wire x_428;
wire x_429;
wire x_430;
wire x_431;
wire x_432;
wire x_433;
wire x_434;
wire x_435;
wire x_436;
wire x_437;
wire x_438;
wire x_439;
wire x_440;
wire x_441;
wire x_442;
wire x_443;
wire x_444;
wire x_445;
wire x_446;
wire x_447;
wire x_448;
wire x_449;
wire x_450;
wire x_451;
wire x_452;
wire x_453;
wire x_454;
wire x_455;
wire x_456;
wire x_457;
wire x_458;
wire x_459;
wire x_460;
wire x_461;
wire x_462;
wire x_463;
wire x_464;
wire x_465;
wire x_466;
wire x_467;
wire x_468;
wire x_469;
wire x_470;
wire x_471;
wire x_472;
wire x_473;
wire x_474;
wire x_475;
wire x_476;
wire x_477;
wire x_478;
wire x_479;
wire x_480;
wire x_481;
wire x_482;
wire x_483;
wire x_484;
wire x_485;
wire x_486;
wire x_487;
wire x_488;
wire x_489;
wire x_490;
wire x_491;
wire x_492;
wire x_493;
wire x_494;
wire x_495;
wire x_496;
wire x_497;
wire x_498;
wire x_499;
wire x_500;
wire x_501;
wire x_502;
wire x_503;
wire x_504;
wire x_505;
wire x_506;
wire x_507;
wire x_508;
wire x_509;
wire x_510;
wire x_511;
wire x_512;
wire x_513;
wire x_514;
wire x_515;
wire x_516;
wire x_517;
wire x_518;
wire x_519;
wire x_520;
wire x_521;
wire x_522;
wire x_523;
wire x_524;
wire x_525;
wire x_526;
wire x_527;
wire x_528;
wire x_529;
wire x_530;
wire x_531;
wire x_532;
wire x_533;
wire x_534;
wire x_535;
wire x_536;
wire x_537;
wire x_538;
wire x_539;
wire x_540;
wire x_541;
wire x_542;
wire x_543;
wire x_544;
wire x_545;
wire x_546;
wire x_547;
wire x_548;
wire x_549;
wire x_550;
wire x_551;
wire x_552;
wire x_553;
wire x_554;
wire x_555;
wire x_556;
wire x_557;
wire x_558;
wire x_559;
wire x_560;
wire x_561;
wire x_562;
wire x_563;
wire x_564;
wire x_565;
wire x_566;
wire x_567;
wire x_568;
wire x_569;
wire x_570;
wire x_571;
wire x_572;
wire x_573;
wire x_574;
wire x_575;
wire x_576;
wire x_577;
wire x_578;
wire x_579;
wire x_580;
wire x_581;
wire x_582;
wire x_583;
wire x_584;
wire x_585;
wire x_586;
wire x_587;
wire x_588;
wire x_589;
wire x_590;
wire x_591;
wire x_592;
wire x_593;
wire x_594;
wire x_595;
wire x_596;
wire x_597;
wire x_598;
wire x_599;
wire x_600;
wire x_601;
wire x_602;
wire x_603;
wire x_604;
wire x_605;
wire x_606;
wire x_607;
wire x_608;
wire x_609;
wire x_610;
wire x_611;
wire x_612;
wire x_613;
wire x_614;
wire x_615;
wire x_616;
wire x_617;
wire x_618;
wire x_619;
wire x_620;
wire x_621;
wire x_622;
wire x_623;
wire x_624;
wire x_625;
wire x_626;
wire x_627;
wire x_628;
wire x_629;
wire x_630;
wire x_631;
wire x_632;
wire x_633;
wire x_634;
wire x_635;
wire x_636;
wire x_637;
wire x_638;
wire x_639;
wire x_640;
wire x_641;
wire x_642;
wire x_643;
wire x_644;
wire x_645;
wire x_646;
wire x_647;
wire x_648;
wire x_649;
wire x_650;
wire x_651;
wire x_652;
wire x_653;
wire x_654;
wire x_655;
wire x_656;
wire x_657;
wire x_658;
wire x_659;
wire x_660;
wire x_661;
wire x_662;
wire x_663;
wire x_664;
wire x_665;
wire x_666;
wire x_667;
wire x_668;
wire x_669;
wire x_670;
wire x_671;
wire x_672;
wire x_673;
wire x_674;
wire x_675;
wire x_676;
wire x_677;
wire x_678;
wire x_679;
wire x_680;
wire x_681;
wire x_682;
wire x_683;
wire x_684;
wire x_685;
wire x_686;
wire x_687;
wire x_688;
wire x_689;
wire x_690;
wire x_691;
wire x_692;
wire x_693;
wire x_694;
wire x_695;
wire x_696;
wire x_697;
wire x_698;
wire x_699;
wire x_700;
wire x_701;
wire x_702;
wire x_703;
wire x_704;
wire x_705;
wire x_706;
wire x_707;
wire x_708;
wire x_709;
wire x_710;
wire x_711;
wire x_712;
wire x_713;
wire x_714;
wire x_715;
wire x_716;
wire x_717;
wire x_718;
wire x_719;
wire x_720;
wire x_721;
wire x_722;
wire x_723;
wire x_724;
wire x_725;
wire x_726;
wire x_727;
wire x_728;
wire x_729;
wire x_730;
wire x_731;
wire x_732;
wire x_733;
wire x_734;
wire x_735;
wire x_736;
wire x_737;
wire x_738;
wire x_739;
wire x_740;
wire x_741;
wire x_742;
wire x_743;
wire x_744;
wire x_745;
wire x_746;
wire x_747;
wire x_748;
wire x_749;
wire x_750;
wire x_751;
wire x_752;
wire x_753;
wire x_754;
wire x_755;
wire x_756;
wire x_757;
wire x_758;
wire x_759;
wire x_760;
wire x_761;
wire x_762;
wire x_763;
wire x_764;
wire x_765;
wire x_766;
wire x_767;
wire x_768;
wire x_769;
wire x_770;
wire x_771;
wire x_772;
wire x_773;
wire x_774;
wire x_775;
wire x_776;
wire x_777;
wire x_778;
wire x_779;
wire x_780;
wire x_781;
wire x_782;
wire x_783;
wire x_784;
wire x_785;
wire x_786;
wire x_787;
wire x_788;
wire x_789;
wire x_790;
wire x_791;
wire x_792;
wire x_793;
wire x_794;
wire x_795;
wire x_796;
wire x_797;
wire x_798;
wire x_799;
wire x_800;
wire x_801;
wire x_802;
wire x_803;
wire x_804;
wire x_805;
wire x_806;
wire x_807;
wire x_808;
wire x_809;
wire x_810;
wire x_811;
wire x_812;
wire x_813;
wire x_814;
wire x_815;
wire x_816;
wire x_817;
wire x_818;
wire x_819;
wire x_820;
wire x_821;
wire x_822;
wire x_823;
wire x_824;
wire x_825;
wire x_826;
wire x_827;
wire x_828;
wire x_829;
wire x_830;
wire x_831;
wire x_832;
wire x_833;
wire x_834;
wire x_835;
wire x_836;
wire x_837;
wire x_838;
wire x_839;
wire x_840;
wire x_841;
wire x_842;
wire x_843;
wire x_844;
wire x_845;
wire x_846;
wire x_847;
wire x_848;
wire x_849;
wire x_850;
wire x_851;
wire x_852;
wire x_853;
wire x_854;
wire x_855;
wire x_856;
wire x_857;
wire x_858;
wire x_859;
wire x_860;
wire x_861;
wire x_862;
wire x_863;
wire x_864;
wire x_865;
wire x_866;
wire x_867;
wire x_868;
wire x_869;
wire x_870;
wire x_871;
wire x_872;
wire x_873;
wire x_874;
wire x_875;
wire x_876;
wire x_877;
wire x_878;
wire x_879;
wire x_880;
wire x_881;
wire x_882;
wire x_883;
wire x_884;
wire x_885;
wire x_886;
wire x_887;
wire x_888;
wire x_889;
wire x_890;
wire x_891;
wire x_892;
wire x_893;
wire x_894;
wire x_895;
wire x_896;
wire x_897;
wire x_898;
wire x_899;
wire x_900;
wire x_901;
wire x_902;
wire x_903;
wire x_904;
wire x_905;
wire x_906;
wire x_907;
wire x_908;
wire x_909;
wire x_910;
wire x_911;
wire x_912;
wire x_913;
wire x_914;
wire x_915;
wire x_916;
wire x_917;
wire x_918;
wire x_919;
wire x_920;
wire x_921;
wire x_922;
wire x_923;
wire x_924;
wire x_925;
wire x_926;
wire x_927;
wire x_928;
wire x_929;
wire x_930;
wire x_931;
wire x_932;
wire x_933;
wire x_934;
wire x_935;
wire x_936;
wire x_937;
wire x_938;
wire x_939;
wire x_940;
wire x_941;
wire x_942;
wire x_943;
wire x_944;
wire x_945;
wire x_946;
wire x_947;
wire x_948;
wire x_949;
wire x_950;
wire x_951;
wire x_952;
wire x_953;
wire x_954;
wire x_955;
wire x_956;
wire x_957;
wire x_958;
wire x_959;
wire x_960;
wire x_961;
wire x_962;
wire x_963;
wire x_964;
wire x_965;
wire x_966;
wire x_967;
wire x_968;
wire x_969;
wire x_970;
wire x_971;
wire x_972;
wire x_973;
wire x_974;
wire x_975;
wire x_976;
wire x_977;
wire x_978;
wire x_979;
wire x_980;
wire x_981;
wire x_982;
wire x_983;
wire x_984;
wire x_985;
wire x_986;
wire x_987;
wire x_988;
wire x_989;
wire x_990;
wire x_991;
wire x_992;
wire x_993;
wire x_994;
wire x_995;
wire x_996;
wire x_997;
wire x_998;
wire x_999;
wire x_1000;
wire x_1001;
wire x_1002;
wire x_1003;
wire x_1004;
wire x_1005;
wire x_1006;
wire x_1007;
wire x_1008;
wire x_1009;
wire x_1010;
wire x_1011;
wire x_1012;
wire x_1013;
wire x_1014;
wire x_1015;
wire x_1016;
wire x_1017;
wire x_1018;
wire x_1019;
wire x_1020;
wire x_1021;
wire x_1022;
wire x_1023;
wire x_1024;
wire x_1025;
wire x_1026;
wire x_1027;
wire x_1028;
wire x_1029;
wire x_1030;
wire x_1031;
wire x_1032;
wire x_1033;
wire x_1034;
wire x_1035;
wire x_1036;
wire x_1037;
wire x_1038;
wire x_1039;
wire x_1040;
wire x_1041;
wire x_1042;
wire x_1043;
wire x_1044;
wire x_1045;
wire x_1046;
wire x_1047;
wire x_1048;
wire x_1049;
wire x_1050;
wire x_1051;
wire x_1052;
wire x_1053;
wire x_1054;
wire x_1055;
wire x_1056;
wire x_1057;
wire x_1058;
wire x_1059;
wire x_1060;
wire x_1061;
wire x_1062;
wire x_1063;
wire x_1064;
wire x_1065;
wire x_1066;
wire x_1067;
wire x_1068;
wire x_1069;
wire x_1070;
wire x_1071;
wire x_1072;
wire x_1073;
wire x_1074;
wire x_1075;
wire x_1076;
wire x_1077;
wire x_1078;
wire x_1079;
wire x_1080;
wire x_1081;
wire x_1082;
wire x_1083;
wire x_1084;
wire x_1085;
wire x_1086;
wire x_1087;
wire x_1088;
wire x_1089;
wire x_1090;
wire x_1091;
wire x_1092;
wire x_1093;
wire x_1094;
wire x_1095;
wire x_1096;
wire x_1097;
wire x_1098;
wire x_1099;
wire x_1100;
wire x_1101;
wire x_1102;
wire x_1103;
wire x_1104;
wire x_1105;
wire x_1106;
wire x_1107;
wire x_1108;
wire x_1109;
wire x_1110;
wire x_1111;
wire x_1112;
wire x_1113;
wire x_1114;
wire x_1115;
wire x_1116;
wire x_1117;
wire x_1118;
wire x_1119;
wire x_1120;
wire x_1121;
wire x_1122;
wire x_1123;
wire x_1124;
wire x_1125;
wire x_1126;
wire x_1127;
wire x_1128;
wire x_1129;
wire x_1130;
wire x_1131;
wire x_1132;
wire x_1133;
wire x_1134;
wire x_1135;
wire x_1136;
wire x_1137;
wire x_1138;
wire x_1139;
wire x_1140;
wire x_1141;
wire x_1142;
wire x_1143;
wire x_1144;
wire x_1145;
wire x_1146;
wire x_1147;
wire x_1148;
wire x_1149;
wire x_1150;
wire x_1151;
wire x_1152;
wire x_1153;
wire x_1154;
wire x_1155;
wire x_1156;
wire x_1157;
wire x_1158;
wire x_1159;
wire x_1160;
wire x_1161;
wire x_1162;
wire x_1163;
wire x_1164;
wire x_1165;
wire x_1166;
wire x_1167;
wire x_1168;
wire x_1169;
wire x_1170;
wire x_1171;
wire x_1172;
wire x_1173;
wire x_1174;
wire x_1175;
wire x_1176;
wire x_1177;
wire x_1178;
wire x_1179;
wire x_1180;
wire x_1181;
wire x_1182;
wire x_1183;
wire x_1184;
wire x_1185;
wire x_1186;
wire x_1187;
wire x_1188;
wire x_1189;
wire x_1190;
wire x_1191;
wire x_1192;
wire x_1193;
wire x_1194;
wire x_1195;
wire x_1196;
wire x_1197;
wire x_1198;
wire x_1199;
wire x_1200;
wire x_1201;
wire x_1202;
wire x_1203;
wire x_1204;
wire x_1205;
wire x_1206;
wire x_1207;
wire x_1208;
wire x_1209;
wire x_1210;
wire x_1211;
wire x_1212;
wire x_1213;
wire x_1214;
wire x_1215;
wire x_1216;
wire x_1217;
wire x_1218;
wire x_1219;
wire x_1220;
wire x_1221;
wire x_1222;
wire x_1223;
wire x_1224;
wire x_1225;
wire x_1226;
wire x_1227;
wire x_1228;
wire x_1229;
wire x_1230;
wire x_1231;
wire x_1232;
wire x_1233;
wire x_1234;
wire x_1235;
wire x_1236;
wire x_1237;
wire x_1238;
wire x_1239;
wire x_1240;
wire x_1241;
wire x_1242;
wire x_1243;
wire x_1244;
wire x_1245;
wire x_1246;
wire x_1247;
wire x_1248;
wire x_1249;
wire x_1250;
wire x_1251;
wire x_1252;
wire x_1253;
wire x_1254;
wire x_1255;
wire x_1256;
wire x_1257;
wire x_1258;
wire x_1259;
wire x_1260;
wire x_1261;
wire x_1262;
wire x_1263;
wire x_1264;
wire x_1265;
wire x_1266;
wire x_1267;
wire x_1268;
wire x_1269;
wire x_1270;
wire x_1271;
wire x_1272;
wire x_1273;
wire x_1274;
wire x_1275;
wire x_1276;
wire x_1277;
wire x_1278;
wire x_1279;
wire x_1280;
wire x_1281;
wire x_1282;
wire x_1283;
wire x_1284;
wire x_1285;
wire x_1286;
wire x_1287;
wire x_1288;
wire x_1289;
wire x_1290;
wire x_1291;
wire x_1292;
wire x_1293;
wire x_1294;
wire x_1295;
wire x_1296;
wire x_1297;
wire x_1298;
wire x_1299;
wire x_1300;
wire x_1301;
wire x_1302;
wire x_1303;
wire x_1304;
wire x_1305;
wire x_1306;
wire x_1307;
wire x_1308;
wire x_1309;
wire x_1310;
wire x_1311;
wire x_1312;
wire x_1313;
wire x_1314;
wire x_1315;
wire x_1316;
wire x_1317;
wire x_1318;
wire x_1319;
wire x_1320;
wire x_1321;
wire x_1322;
wire x_1323;
wire x_1324;
wire x_1325;
wire x_1326;
wire x_1327;
wire x_1328;
wire x_1329;
wire x_1330;
wire x_1331;
wire x_1332;
wire x_1333;
wire x_1334;
wire x_1335;
wire x_1336;
wire x_1337;
wire x_1338;
wire x_1339;
wire x_1340;
wire x_1341;
wire x_1342;
wire x_1343;
wire x_1344;
wire x_1345;
wire x_1346;
wire x_1347;
wire x_1348;
wire x_1349;
wire x_1350;
wire x_1351;
wire x_1352;
wire x_1353;
wire x_1354;
wire x_1355;
wire x_1356;
wire x_1357;
wire x_1358;
wire x_1359;
wire x_1360;
wire x_1361;
wire x_1362;
wire x_1363;
wire x_1364;
wire x_1365;
wire x_1366;
wire x_1367;
wire x_1368;
wire x_1369;
wire x_1370;
wire x_1371;
wire x_1372;
wire x_1373;
wire x_1374;
wire x_1375;
wire x_1376;
wire x_1377;
wire x_1378;
wire x_1379;
wire x_1380;
wire x_1381;
wire x_1382;
wire x_1383;
wire x_1384;
wire x_1385;
wire x_1386;
wire x_1387;
wire x_1388;
wire x_1389;
wire x_1390;
wire x_1391;
wire x_1392;
wire x_1393;
wire x_1394;
wire x_1395;
wire x_1396;
wire x_1397;
wire x_1398;
wire x_1399;
wire x_1400;
wire x_1401;
wire x_1402;
wire x_1403;
wire x_1404;
wire x_1405;
wire x_1406;
wire x_1407;
wire x_1408;
wire x_1409;
wire x_1410;
wire x_1411;
wire x_1412;
wire x_1413;
wire x_1414;
wire x_1415;
wire x_1416;
wire x_1417;
wire x_1418;
wire x_1419;
wire x_1420;
wire x_1421;
wire x_1422;
wire x_1423;
wire x_1424;
wire x_1425;
wire x_1426;
wire x_1427;
wire x_1428;
wire x_1429;
wire x_1430;
wire x_1431;
wire x_1432;
wire x_1433;
wire x_1434;
wire x_1435;
wire x_1436;
wire x_1437;
wire x_1438;
wire x_1439;
wire x_1440;
wire x_1441;
wire x_1442;
wire x_1443;
wire x_1444;
wire x_1445;
wire x_1446;
wire x_1447;
wire x_1448;
wire x_1449;
wire x_1450;
wire x_1451;
wire x_1452;
wire x_1453;
wire x_1454;
wire x_1455;
wire x_1456;
wire x_1457;
wire x_1458;
wire x_1459;
wire x_1460;
wire x_1461;
wire x_1462;
wire x_1463;
wire x_1464;
wire x_1465;
wire x_1466;
wire x_1467;
wire x_1468;
wire x_1469;
wire x_1470;
wire x_1471;
wire x_1472;
wire x_1473;
wire x_1474;
wire x_1475;
wire x_1476;
wire x_1477;
wire x_1478;
wire x_1479;
wire x_1480;
wire x_1481;
wire x_1482;
wire x_1483;
wire x_1484;
wire x_1485;
wire x_1486;
wire x_1487;
wire x_1488;
wire x_1489;
wire x_1490;
wire x_1491;
wire x_1492;
wire x_1493;
wire x_1494;
wire x_1495;
wire x_1496;
wire x_1497;
wire x_1498;
wire x_1499;
wire x_1500;
wire x_1501;
wire x_1502;
wire x_1503;
wire x_1504;
wire x_1505;
wire x_1506;
wire x_1507;
wire x_1508;
wire x_1509;
wire x_1510;
wire x_1511;
wire x_1512;
wire x_1513;
wire x_1514;
wire x_1515;
wire x_1516;
wire x_1517;
wire x_1518;
wire x_1519;
wire x_1520;
wire x_1521;
wire x_1522;
wire x_1523;
wire x_1524;
wire x_1525;
wire x_1526;
wire x_1527;
wire x_1528;
wire x_1529;
wire x_1530;
wire x_1531;
wire x_1532;
wire x_1533;
wire x_1534;
wire x_1535;
wire x_1536;
wire x_1537;
wire x_1538;
wire x_1539;
wire x_1540;
wire x_1541;
wire x_1542;
wire x_1543;
wire x_1544;
wire x_1545;
wire x_1546;
wire x_1547;
wire x_1548;
wire x_1549;
wire x_1550;
wire x_1551;
wire x_1552;
wire x_1553;
wire x_1554;
wire x_1555;
wire x_1556;
wire x_1557;
wire x_1558;
wire x_1559;
wire x_1560;
wire x_1561;
wire x_1562;
wire x_1563;
wire x_1564;
wire x_1565;
wire x_1566;
wire x_1567;
wire x_1568;
wire x_1569;
wire x_1570;
wire x_1571;
wire x_1572;
wire x_1573;
wire x_1574;
wire x_1575;
wire x_1576;
wire x_1577;
wire x_1578;
wire x_1579;
wire x_1580;
wire x_1581;
wire x_1582;
wire x_1583;
wire x_1584;
wire x_1585;
wire x_1586;
wire x_1587;
wire x_1588;
wire x_1589;
wire x_1590;
wire x_1591;
wire x_1592;
wire x_1593;
wire x_1594;
wire x_1595;
wire x_1596;
wire x_1597;
wire x_1598;
wire x_1599;
wire x_1600;
wire x_1601;
wire x_1602;
wire x_1603;
wire x_1604;
wire x_1605;
wire x_1606;
wire x_1607;
wire x_1608;
wire x_1609;
wire x_1610;
wire x_1611;
wire x_1612;
wire x_1613;
wire x_1614;
wire x_1615;
wire x_1616;
wire x_1617;
wire x_1618;
wire x_1619;
wire x_1620;
wire x_1621;
wire x_1622;
wire x_1623;
wire x_1624;
wire x_1625;
wire x_1626;
wire x_1627;
wire x_1628;
wire x_1629;
wire x_1630;
wire x_1631;
wire x_1632;
wire x_1633;
wire x_1634;
wire x_1635;
wire x_1636;
wire x_1637;
wire x_1638;
wire x_1639;
wire x_1640;
wire x_1641;
wire x_1642;
wire x_1643;
wire x_1644;
wire x_1645;
wire x_1646;
wire x_1647;
wire x_1648;
wire x_1649;
wire x_1650;
wire x_1651;
wire x_1652;
wire x_1653;
wire x_1654;
wire x_1655;
wire x_1656;
wire x_1657;
wire x_1658;
wire x_1659;
wire x_1660;
wire x_1661;
wire x_1662;
wire x_1663;
wire x_1664;
wire x_1665;
wire x_1666;
wire x_1667;
wire x_1668;
wire x_1669;
wire x_1670;
wire x_1671;
wire x_1672;
wire x_1673;
wire x_1674;
wire x_1675;
wire x_1676;
wire x_1677;
wire x_1678;
wire x_1679;
wire x_1680;
wire x_1681;
wire x_1682;
wire x_1683;
wire x_1684;
wire x_1685;
wire x_1686;
wire x_1687;
wire x_1688;
wire x_1689;
wire x_1690;
wire x_1691;
wire x_1692;
wire x_1693;
wire x_1694;
wire x_1695;
wire x_1696;
wire x_1697;
wire x_1698;
wire x_1699;
wire x_1700;
wire x_1701;
wire x_1702;
wire x_1703;
wire x_1704;
wire x_1705;
wire x_1706;
wire x_1707;
wire x_1708;
wire x_1709;
wire x_1710;
wire x_1711;
wire x_1712;
wire x_1713;
wire x_1714;
wire x_1715;
wire x_1716;
wire x_1717;
wire x_1718;
wire x_1719;
wire x_1720;
wire x_1721;
wire x_1722;
wire x_1723;
wire x_1724;
wire x_1725;
wire x_1726;
wire x_1727;
wire x_1728;
wire x_1729;
wire x_1730;
wire x_1731;
wire x_1732;
wire x_1733;
wire x_1734;
wire x_1735;
wire x_1736;
wire x_1737;
wire x_1738;
wire x_1739;
wire x_1740;
wire x_1741;
wire x_1742;
wire x_1743;
wire x_1744;
wire x_1745;
wire x_1746;
wire x_1747;
wire x_1748;
wire x_1749;
wire x_1750;
wire x_1751;
wire x_1752;
wire x_1753;
wire x_1754;
wire x_1755;
wire x_1756;
wire x_1757;
wire x_1758;
wire x_1759;
wire x_1760;
wire x_1761;
wire x_1762;
wire x_1763;
wire x_1764;
wire x_1765;
wire x_1766;
wire x_1767;
wire x_1768;
wire x_1769;
wire x_1770;
wire x_1771;
wire x_1772;
wire x_1773;
wire x_1774;
wire x_1775;
wire x_1776;
wire x_1777;
wire x_1778;
wire x_1779;
wire x_1780;
wire x_1781;
wire x_1782;
wire x_1783;
wire x_1784;
wire x_1785;
wire x_1786;
wire x_1787;
wire x_1788;
wire x_1789;
wire x_1790;
wire x_1791;
wire x_1792;
wire x_1793;
wire x_1794;
wire x_1795;
wire x_1796;
wire x_1797;
wire x_1798;
wire x_1799;
wire x_1800;
wire x_1801;
wire x_1802;
wire x_1803;
wire x_1804;
wire x_1805;
wire x_1806;
wire x_1807;
wire x_1808;
wire x_1809;
wire x_1810;
wire x_1811;
wire x_1812;
wire x_1813;
wire x_1814;
wire x_1815;
wire x_1816;
wire x_1817;
wire x_1818;
wire x_1819;
wire x_1820;
wire x_1821;
wire x_1822;
wire x_1823;
wire x_1824;
wire x_1825;
wire x_1826;
wire x_1827;
wire x_1828;
wire x_1829;
wire x_1830;
wire x_1831;
wire x_1832;
wire x_1833;
wire x_1834;
wire x_1835;
wire x_1836;
wire x_1837;
wire x_1838;
wire x_1839;
wire x_1840;
wire x_1841;
wire x_1842;
wire x_1843;
wire x_1844;
wire x_1845;
wire x_1846;
wire x_1847;
wire x_1848;
wire x_1849;
wire x_1850;
wire x_1851;
wire x_1852;
wire x_1853;
wire x_1854;
wire x_1855;
wire x_1856;
wire x_1857;
wire x_1858;
wire x_1859;
wire x_1860;
wire x_1861;
wire x_1862;
wire x_1863;
wire x_1864;
wire x_1865;
wire x_1866;
wire x_1867;
wire x_1868;
wire x_1869;
wire x_1870;
wire x_1871;
wire x_1872;
wire x_1873;
wire x_1874;
wire x_1875;
wire x_1876;
wire x_1877;
wire x_1878;
wire x_1879;
wire x_1880;
wire x_1881;
wire x_1882;
wire x_1883;
wire x_1884;
wire x_1885;
wire x_1886;
wire x_1887;
wire x_1888;
wire x_1889;
wire x_1890;
wire x_1891;
wire x_1892;
wire x_1893;
wire x_1894;
wire x_1895;
wire x_1896;
wire x_1897;
wire x_1898;
wire x_1899;
wire x_1900;
wire x_1901;
wire x_1902;
wire x_1903;
wire x_1904;
wire x_1905;
wire x_1906;
wire x_1907;
wire x_1908;
wire x_1909;
wire x_1910;
wire x_1911;
wire x_1912;
wire x_1913;
wire x_1914;
wire x_1915;
wire x_1916;
wire x_1917;
wire x_1918;
wire x_1919;
wire x_1920;
wire x_1921;
wire x_1922;
wire x_1923;
wire x_1924;
wire x_1925;
wire x_1926;
wire x_1927;
wire x_1928;
wire x_1929;
wire x_1930;
wire x_1931;
wire x_1932;
wire x_1933;
wire x_1934;
wire x_1935;
wire x_1936;
wire x_1937;
wire x_1938;
wire x_1939;
wire x_1940;
wire x_1941;
wire x_1942;
wire x_1943;
wire x_1944;
wire x_1945;
wire x_1946;
wire x_1947;
wire x_1948;
wire x_1949;
wire x_1950;
wire x_1951;
wire x_1952;
wire x_1953;
wire x_1954;
wire x_1955;
wire x_1956;
wire x_1957;
wire x_1958;
wire x_1959;
wire x_1960;
wire x_1961;
wire x_1962;
wire x_1963;
wire x_1964;
wire x_1965;
wire x_1966;
wire x_1967;
wire x_1968;
wire x_1969;
wire x_1970;
wire x_1971;
wire x_1972;
wire x_1973;
wire x_1974;
wire x_1975;
wire x_1976;
wire x_1977;
wire x_1978;
wire x_1979;
wire x_1980;
wire x_1981;
wire x_1982;
wire x_1983;
wire x_1984;
wire x_1985;
wire x_1986;
wire x_1987;
wire x_1988;
wire x_1989;
wire x_1990;
wire x_1991;
wire x_1992;
wire x_1993;
wire x_1994;
wire x_1995;
wire x_1996;
wire x_1997;
wire x_1998;
wire x_1999;
wire x_2000;
wire x_2001;
wire x_2002;
wire x_2003;
wire x_2004;
wire x_2005;
wire x_2006;
wire x_2007;
wire x_2008;
wire x_2009;
wire x_2010;
wire x_2011;
wire x_2012;
wire x_2013;
wire x_2014;
wire x_2015;
wire x_2016;
wire x_2017;
wire x_2018;
wire x_2019;
wire x_2020;
wire x_2021;
wire x_2022;
wire x_2023;
wire x_2024;
wire x_2025;
wire x_2026;
wire x_2027;
wire x_2028;
wire x_2029;
wire x_2030;
wire x_2031;
wire x_2032;
wire x_2033;
wire x_2034;
wire x_2035;
wire x_2036;
wire x_2037;
wire x_2038;
wire x_2039;
wire x_2040;
wire x_2041;
wire x_2042;
wire x_2043;
wire x_2044;
wire x_2045;
wire x_2046;
wire x_2047;
wire x_2048;
wire x_2049;
wire x_2050;
wire x_2051;
wire x_2052;
wire x_2053;
wire x_2054;
wire x_2055;
wire x_2056;
wire x_2057;
wire x_2058;
wire x_2059;
wire x_2060;
wire x_2061;
wire x_2062;
wire x_2063;
wire x_2064;
wire x_2065;
wire x_2066;
wire x_2067;
wire x_2068;
wire x_2069;
wire x_2070;
wire x_2071;
wire x_2072;
wire x_2073;
wire x_2074;
wire x_2075;
wire x_2076;
wire x_2077;
wire x_2078;
wire x_2079;
wire x_2080;
wire x_2081;
wire x_2082;
wire x_2083;
wire x_2084;
wire x_2085;
wire x_2086;
wire x_2087;
wire x_2088;
wire x_2089;
wire x_2090;
wire x_2091;
wire x_2092;
wire x_2093;
wire x_2094;
wire x_2095;
wire x_2096;
wire x_2097;
wire x_2098;
wire x_2099;
wire x_2100;
wire x_2101;
wire x_2102;
wire x_2103;
wire x_2104;
wire x_2105;
wire x_2106;
wire x_2107;
wire x_2108;
wire x_2109;
wire x_2110;
wire x_2111;
wire x_2112;
wire x_2113;
wire x_2114;
wire x_2115;
wire x_2116;
wire x_2117;
wire x_2118;
wire x_2119;
wire x_2120;
wire x_2121;
wire x_2122;
wire x_2123;
wire x_2124;
wire x_2125;
wire x_2126;
wire x_2127;
wire x_2128;
wire x_2129;
wire x_2130;
wire x_2131;
wire x_2132;
wire x_2133;
wire x_2134;
wire x_2135;
wire x_2136;
wire x_2137;
wire x_2138;
wire x_2139;
wire x_2140;
wire x_2141;
wire x_2142;
wire x_2143;
wire x_2144;
wire x_2145;
wire x_2146;
wire x_2147;
wire x_2148;
wire x_2149;
wire x_2150;
wire x_2151;
wire x_2152;
wire x_2153;
wire x_2154;
wire x_2155;
wire x_2156;
wire x_2157;
wire x_2158;
wire x_2159;
wire x_2160;
wire x_2161;
wire x_2162;
wire x_2163;
wire x_2164;
wire x_2165;
wire x_2166;
wire x_2167;
wire x_2168;
wire x_2169;
wire x_2170;
wire x_2171;
wire x_2172;
wire x_2173;
wire x_2174;
wire x_2175;
wire x_2176;
wire x_2177;
wire x_2178;
wire x_2179;
wire x_2180;
wire x_2181;
wire x_2182;
wire x_2183;
wire x_2184;
wire x_2185;
wire x_2186;
wire x_2187;
wire x_2188;
wire x_2189;
wire x_2190;
wire x_2191;
wire x_2192;
wire x_2193;
wire x_2194;
wire x_2195;
wire x_2196;
wire x_2197;
wire x_2198;
wire x_2199;
wire x_2200;
wire x_2201;
wire x_2202;
wire x_2203;
wire x_2204;
wire x_2205;
wire x_2206;
wire x_2207;
wire x_2208;
wire x_2209;
wire x_2210;
wire x_2211;
wire x_2212;
wire x_2213;
wire x_2214;
wire x_2215;
wire x_2216;
wire x_2217;
wire x_2218;
wire x_2219;
wire x_2220;
wire x_2221;
wire x_2222;
wire x_2223;
wire x_2224;
wire x_2225;
wire x_2226;
wire x_2227;
wire x_2228;
wire x_2229;
wire x_2230;
wire x_2231;
wire x_2232;
wire x_2233;
wire x_2234;
wire x_2235;
wire x_2236;
wire x_2237;
wire x_2238;
wire x_2239;
wire x_2240;
wire x_2241;
wire x_2242;
wire x_2243;
wire x_2244;
wire x_2245;
wire x_2246;
wire x_2247;
wire x_2248;
wire x_2249;
wire x_2250;
wire x_2251;
wire x_2252;
wire x_2253;
wire x_2254;
wire x_2255;
wire x_2256;
wire x_2257;
wire x_2258;
wire x_2259;
wire x_2260;
wire x_2261;
wire x_2262;
wire x_2263;
wire x_2264;
wire x_2265;
wire x_2266;
wire x_2267;
wire x_2268;
wire x_2269;
wire x_2270;
wire x_2271;
wire x_2272;
wire x_2273;
wire x_2274;
wire x_2275;
wire x_2276;
wire x_2277;
wire x_2278;
wire x_2279;
wire x_2280;
wire x_2281;
wire x_2282;
wire x_2283;
wire x_2284;
wire x_2285;
wire x_2286;
wire x_2287;
wire x_2288;
wire x_2289;
wire x_2290;
wire x_2291;
wire x_2292;
wire x_2293;
wire x_2294;
wire x_2295;
wire x_2296;
wire x_2297;
wire x_2298;
wire x_2299;
wire x_2300;
wire x_2301;
wire x_2302;
wire x_2303;
wire x_2304;
wire x_2305;
wire x_2306;
wire x_2307;
wire x_2308;
wire x_2309;
wire x_2310;
wire x_2311;
wire x_2312;
wire x_2313;
wire x_2314;
wire x_2315;
wire x_2316;
wire x_2317;
wire x_2318;
wire x_2319;
wire x_2320;
wire x_2321;
wire x_2322;
wire x_2323;
wire x_2324;
wire x_2325;
wire x_2326;
wire x_2327;
wire x_2328;
wire x_2329;
wire x_2330;
wire x_2331;
wire x_2332;
wire x_2333;
wire x_2334;
wire x_2335;
wire x_2336;
wire x_2337;
wire x_2338;
wire x_2339;
wire x_2340;
wire x_2341;
wire x_2342;
wire x_2343;
wire x_2344;
wire x_2345;
wire x_2346;
wire x_2347;
wire x_2348;
wire x_2349;
wire x_2350;
wire x_2351;
wire x_2352;
wire x_2353;
wire x_2354;
wire x_2355;
wire x_2356;
wire x_2357;
wire x_2358;
wire x_2359;
wire x_2360;
wire x_2361;
wire x_2362;
wire x_2363;
wire x_2364;
wire x_2365;
wire x_2366;
wire x_2367;
wire x_2368;
wire x_2369;
wire x_2370;
wire x_2371;
wire x_2372;
wire x_2373;
wire x_2374;
wire x_2375;
wire x_2376;
wire x_2377;
wire x_2378;
wire x_2379;
wire x_2380;
wire x_2381;
wire x_2382;
wire x_2383;
wire x_2384;
wire x_2385;
wire x_2386;
wire x_2387;
wire x_2388;
wire x_2389;
wire x_2390;
wire x_2391;
wire x_2392;
wire x_2393;
wire x_2394;
wire x_2395;
wire x_2396;
wire x_2397;
wire x_2398;
wire x_2399;
wire x_2400;
wire x_2401;
wire x_2402;
wire x_2403;
wire x_2404;
wire x_2405;
wire x_2406;
wire x_2407;
wire x_2408;
wire x_2409;
wire x_2410;
wire x_2411;
wire x_2412;
wire x_2413;
wire x_2414;
wire x_2415;
wire x_2416;
wire x_2417;
wire x_2418;
wire x_2419;
wire x_2420;
wire x_2421;
wire x_2422;
wire x_2423;
wire x_2424;
wire x_2425;
wire x_2426;
wire x_2427;
wire x_2428;
wire x_2429;
wire x_2430;
wire x_2431;
wire x_2432;
wire x_2433;
wire x_2434;
wire x_2435;
wire x_2436;
wire x_2437;
wire x_2438;
wire x_2439;
wire x_2440;
wire x_2441;
wire x_2442;
wire x_2443;
wire x_2444;
wire x_2445;
wire x_2446;
wire x_2447;
wire x_2448;
wire x_2449;
wire x_2450;
wire x_2451;
wire x_2452;
wire x_2453;
wire x_2454;
wire x_2455;
wire x_2456;
wire x_2457;
wire x_2458;
wire x_2459;
wire x_2460;
wire x_2461;
wire x_2462;
wire x_2463;
wire x_2464;
wire x_2465;
wire x_2466;
wire x_2467;
wire x_2468;
wire x_2469;
wire x_2470;
wire x_2471;
wire x_2472;
wire x_2473;
wire x_2474;
wire x_2475;
wire x_2476;
wire x_2477;
wire x_2478;
wire x_2479;
wire x_2480;
wire x_2481;
wire x_2482;
wire x_2483;
wire x_2484;
wire x_2485;
wire x_2486;
wire x_2487;
wire x_2488;
wire x_2489;
wire x_2490;
wire x_2491;
wire x_2492;
wire x_2493;
wire x_2494;
wire x_2495;
wire x_2496;
wire x_2497;
wire x_2498;
wire x_2499;
wire x_2500;
wire x_2501;
wire x_2502;
wire x_2503;
wire x_2504;
wire x_2505;
wire x_2506;
wire x_2507;
wire x_2508;
wire x_2509;
wire x_2510;
wire x_2511;
wire x_2512;
wire x_2513;
wire x_2514;
wire x_2515;
wire x_2516;
wire x_2517;
wire x_2518;
wire x_2519;
wire x_2520;
wire x_2521;
wire x_2522;
wire x_2523;
wire x_2524;
wire x_2525;
wire x_2526;
wire x_2527;
wire x_2528;
wire x_2529;
wire x_2530;
wire x_2531;
wire x_2532;
wire x_2533;
wire x_2534;
wire x_2535;
wire x_2536;
wire x_2537;
wire x_2538;
wire x_2539;
wire x_2540;
wire x_2541;
wire x_2542;
wire x_2543;
wire x_2544;
wire x_2545;
wire x_2546;
wire x_2547;
wire x_2548;
wire x_2549;
wire x_2550;
wire x_2551;
wire x_2552;
wire x_2553;
wire x_2554;
wire x_2555;
wire x_2556;
wire x_2557;
wire x_2558;
wire x_2559;
wire x_2560;
wire x_2561;
wire x_2562;
wire x_2563;
wire x_2564;
wire x_2565;
wire x_2566;
wire x_2567;
wire x_2568;
wire x_2569;
wire x_2570;
wire x_2571;
wire x_2572;
wire x_2573;
wire x_2574;
wire x_2575;
wire x_2576;
wire x_2577;
wire x_2578;
wire x_2579;
wire x_2580;
wire x_2581;
wire x_2582;
wire x_2583;
wire x_2584;
wire x_2585;
wire x_2586;
wire x_2587;
wire x_2588;
wire x_2589;
wire x_2590;
wire x_2591;
wire x_2592;
wire x_2593;
wire x_2594;
wire x_2595;
wire x_2596;
wire x_2597;
wire x_2598;
wire x_2599;
wire x_2600;
wire x_2601;
wire x_2602;
wire x_2603;
wire x_2604;
wire x_2605;
wire x_2606;
wire x_2607;
wire x_2608;
wire x_2609;
wire x_2610;
wire x_2611;
wire x_2612;
wire x_2613;
wire x_2614;
wire x_2615;
wire x_2616;
wire x_2617;
wire x_2618;
wire x_2619;
wire x_2620;
wire x_2621;
wire x_2622;
wire x_2623;
wire x_2624;
wire x_2625;
wire x_2626;
wire x_2627;
wire x_2628;
wire x_2629;
wire x_2630;
wire x_2631;
wire x_2632;
wire x_2633;
wire x_2634;
wire x_2635;
wire x_2636;
wire x_2637;
wire x_2638;
wire x_2639;
wire x_2640;
wire x_2641;
wire x_2642;
wire x_2643;
wire x_2644;
wire x_2645;
wire x_2646;
wire x_2647;
wire x_2648;
wire x_2649;
wire x_2650;
wire x_2651;
wire x_2652;
wire x_2653;
wire x_2654;
wire x_2655;
wire x_2656;
wire x_2657;
wire x_2658;
wire x_2659;
wire x_2660;
wire x_2661;
wire x_2662;
wire x_2663;
wire x_2664;
wire x_2665;
wire x_2666;
wire x_2667;
wire x_2668;
wire x_2669;
wire x_2670;
wire x_2671;
wire x_2672;
wire x_2673;
wire x_2674;
wire x_2675;
wire x_2676;
wire x_2677;
wire x_2678;
wire x_2679;
wire x_2680;
wire x_2681;
wire x_2682;
wire x_2683;
wire x_2684;
wire x_2685;
wire x_2686;
wire x_2687;
wire x_2688;
wire x_2689;
wire x_2690;
wire x_2691;
wire x_2692;
wire x_2693;
wire x_2694;
wire x_2695;
wire x_2696;
wire x_2697;
wire x_2698;
wire x_2699;
wire x_2700;
wire x_2701;
wire x_2702;
wire x_2703;
wire x_2704;
wire x_2705;
wire x_2706;
wire x_2707;
wire x_2708;
wire x_2709;
wire x_2710;
wire x_2711;
wire x_2712;
wire x_2713;
wire x_2714;
wire x_2715;
wire x_2716;
wire x_2717;
wire x_2718;
wire x_2719;
wire x_2720;
wire x_2721;
wire x_2722;
wire x_2723;
wire x_2724;
wire x_2725;
wire x_2726;
wire x_2727;
wire x_2728;
wire x_2729;
wire x_2730;
wire x_2731;
wire x_2732;
wire x_2733;
wire x_2734;
wire x_2735;
wire x_2736;
wire x_2737;
wire x_2738;
wire x_2739;
wire x_2740;
wire x_2741;
wire x_2742;
wire x_2743;
wire x_2744;
wire x_2745;
wire x_2746;
wire x_2747;
wire x_2748;
wire x_2749;
wire x_2750;
wire x_2751;
wire x_2752;
wire x_2753;
wire x_2754;
wire x_2755;
wire x_2756;
wire x_2757;
wire x_2758;
wire x_2759;
wire x_2760;
wire x_2761;
wire x_2762;
wire x_2763;
wire x_2764;
wire x_2765;
wire x_2766;
wire x_2767;
wire x_2768;
wire x_2769;
wire x_2770;
wire x_2771;
wire x_2772;
wire x_2773;
wire x_2774;
wire x_2775;
wire x_2776;
wire x_2777;
wire x_2778;
wire x_2779;
wire x_2780;
wire x_2781;
wire x_2782;
wire x_2783;
wire x_2784;
wire x_2785;
wire x_2786;
wire x_2787;
wire x_2788;
wire x_2789;
wire x_2790;
wire x_2791;
wire x_2792;
wire x_2793;
wire x_2794;
wire x_2795;
wire x_2796;
wire x_2797;
wire x_2798;
wire x_2799;
wire x_2800;
wire x_2801;
wire x_2802;
wire x_2803;
wire x_2804;
wire x_2805;
wire x_2806;
wire x_2807;
wire x_2808;
wire x_2809;
wire x_2810;
wire x_2811;
wire x_2812;
wire x_2813;
wire x_2814;
wire x_2815;
wire x_2816;
wire x_2817;
wire x_2818;
wire x_2819;
wire x_2820;
wire x_2821;
wire x_2822;
wire x_2823;
wire x_2824;
wire x_2825;
wire x_2826;
wire x_2827;
wire x_2828;
wire x_2829;
wire x_2830;
wire x_2831;
wire x_2832;
wire x_2833;
wire x_2834;
wire x_2835;
wire x_2836;
wire x_2837;
wire x_2838;
wire x_2839;
wire x_2840;
wire x_2841;
wire x_2842;
wire x_2843;
wire x_2844;
wire x_2845;
wire x_2846;
wire x_2847;
wire x_2848;
wire x_2849;
wire x_2850;
wire x_2851;
wire x_2852;
wire x_2853;
wire x_2854;
wire x_2855;
wire x_2856;
wire x_2857;
wire x_2858;
wire x_2859;
wire x_2860;
wire x_2861;
wire x_2862;
wire x_2863;
wire x_2864;
wire x_2865;
wire x_2866;
wire x_2867;
wire x_2868;
wire x_2869;
wire x_2870;
wire x_2871;
wire x_2872;
wire x_2873;
wire x_2874;
wire x_2875;
wire x_2876;
wire x_2877;
wire x_2878;
wire x_2879;
wire x_2880;
wire x_2881;
wire x_2882;
wire x_2883;
wire x_2884;
wire x_2885;
wire x_2886;
wire x_2887;
wire x_2888;
wire x_2889;
wire x_2890;
wire x_2891;
wire x_2892;
wire x_2893;
wire x_2894;
wire x_2895;
wire x_2896;
wire x_2897;
wire x_2898;
wire x_2899;
wire x_2900;
wire x_2901;
wire x_2902;
wire x_2903;
wire x_2904;
wire x_2905;
wire x_2906;
wire x_2907;
wire x_2908;
wire x_2909;
wire x_2910;
wire x_2911;
wire x_2912;
wire x_2913;
wire x_2914;
wire x_2915;
wire x_2916;
wire x_2917;
wire x_2918;
wire x_2919;
wire x_2920;
wire x_2921;
wire x_2922;
wire x_2923;
wire x_2924;
wire x_2925;
wire x_2926;
wire x_2927;
wire x_2928;
wire x_2929;
wire x_2930;
wire x_2931;
wire x_2932;
wire x_2933;
wire x_2934;
wire x_2935;
wire x_2936;
wire x_2937;
wire x_2938;
wire x_2939;
wire x_2940;
wire x_2941;
wire x_2942;
wire x_2943;
wire x_2944;
wire x_2945;
wire x_2946;
wire x_2947;
wire x_2948;
wire x_2949;
wire x_2950;
wire x_2951;
wire x_2952;
wire x_2953;
wire x_2954;
wire x_2955;
wire x_2956;
wire x_2957;
wire x_2958;
wire x_2959;
wire x_2960;
wire x_2961;
wire x_2962;
wire x_2963;
wire x_2964;
wire x_2965;
wire x_2966;
wire x_2967;
wire x_2968;
wire x_2969;
wire x_2970;
wire x_2971;
wire x_2972;
wire x_2973;
wire x_2974;
wire x_2975;
wire x_2976;
wire x_2977;
wire x_2978;
wire x_2979;
wire x_2980;
wire x_2981;
wire x_2982;
wire x_2983;
wire x_2984;
wire x_2985;
wire x_2986;
wire x_2987;
wire x_2988;
wire x_2989;
wire x_2990;
wire x_2991;
wire x_2992;
wire x_2993;
wire x_2994;
wire x_2995;
wire x_2996;
wire x_2997;
wire x_2998;
wire x_2999;
wire x_3000;
wire x_3001;
wire x_3002;
wire x_3003;
wire x_3004;
wire x_3005;
wire x_3006;
wire x_3007;
wire x_3008;
wire x_3009;
wire x_3010;
wire x_3011;
wire x_3012;
wire x_3013;
wire x_3014;
wire x_3015;
wire x_3016;
wire x_3017;
wire x_3018;
wire x_3019;
wire x_3020;
wire x_3021;
wire x_3022;
wire x_3023;
wire x_3024;
wire x_3025;
wire x_3026;
wire x_3027;
wire x_3028;
wire x_3029;
wire x_3030;
wire x_3031;
wire x_3032;
wire x_3033;
wire x_3034;
wire x_3035;
wire x_3036;
wire x_3037;
wire x_3038;
wire x_3039;
wire x_3040;
wire x_3041;
wire x_3042;
wire x_3043;
wire x_3044;
wire x_3045;
wire x_3046;
wire x_3047;
wire x_3048;
wire x_3049;
wire x_3050;
wire x_3051;
wire x_3052;
wire x_3053;
wire x_3054;
wire x_3055;
wire x_3056;
wire x_3057;
wire x_3058;
wire x_3059;
wire x_3060;
wire x_3061;
wire x_3062;
wire x_3063;
wire x_3064;
wire x_3065;
wire x_3066;
wire x_3067;
wire x_3068;
wire x_3069;
wire x_3070;
wire x_3071;
wire x_3072;
wire x_3073;
wire x_3074;
wire x_3075;
wire x_3076;
wire x_3077;
wire x_3078;
wire x_3079;
wire x_3080;
wire x_3081;
wire x_3082;
wire x_3083;
wire x_3084;
wire x_3085;
wire x_3086;
wire x_3087;
wire x_3088;
wire x_3089;
wire x_3090;
wire x_3091;
wire x_3092;
wire x_3093;
wire x_3094;
wire x_3095;
wire x_3096;
wire x_3097;
wire x_3098;
wire x_3099;
wire x_3100;
wire x_3101;
wire x_3102;
wire x_3103;
wire x_3104;
wire x_3105;
wire x_3106;
wire x_3107;
wire x_3108;
wire x_3109;
wire x_3110;
wire x_3111;
wire x_3112;
wire x_3113;
wire x_3114;
wire x_3115;
wire x_3116;
wire x_3117;
wire x_3118;
wire x_3119;
wire x_3120;
wire x_3121;
wire x_3122;
wire x_3123;
wire x_3124;
wire x_3125;
wire x_3126;
wire x_3127;
wire x_3128;
wire x_3129;
wire x_3130;
wire x_3131;
wire x_3132;
wire x_3133;
wire x_3134;
wire x_3135;
wire x_3136;
wire x_3137;
wire x_3138;
wire x_3139;
wire x_3140;
wire x_3141;
wire x_3142;
wire x_3143;
wire x_3144;
wire x_3145;
wire x_3146;
wire x_3147;
wire x_3148;
wire x_3149;
wire x_3150;
wire x_3151;
wire x_3152;
wire x_3153;
wire x_3154;
wire x_3155;
wire x_3156;
wire x_3157;
wire x_3158;
wire x_3159;
wire x_3160;
wire x_3161;
wire x_3162;
wire x_3163;
wire x_3164;
wire x_3165;
wire x_3166;
wire x_3167;
wire x_3168;
wire x_3169;
wire x_3170;
wire x_3171;
wire x_3172;
wire x_3173;
wire x_3174;
wire x_3175;
wire x_3176;
wire x_3177;
wire x_3178;
wire x_3179;
wire x_3180;
wire x_3181;
wire x_3182;
wire x_3183;
wire x_3184;
wire x_3185;
wire x_3186;
wire x_3187;
wire x_3188;
wire x_3189;
wire x_3190;
wire x_3191;
wire x_3192;
wire x_3193;
wire x_3194;
wire x_3195;
wire x_3196;
wire x_3197;
wire x_3198;
wire x_3199;
wire x_3200;
wire x_3201;
wire x_3202;
wire x_3203;
wire x_3204;
wire x_3205;
wire x_3206;
wire x_3207;
wire x_3208;
wire x_3209;
wire x_3210;
wire x_3211;
wire x_3212;
wire x_3213;
wire x_3214;
wire x_3215;
wire x_3216;
wire x_3217;
wire x_3218;
wire x_3219;
wire x_3220;
wire x_3221;
wire x_3222;
wire x_3223;
wire x_3224;
wire x_3225;
wire x_3226;
wire x_3227;
wire x_3228;
wire x_3229;
wire x_3230;
wire x_3231;
wire x_3232;
wire x_3233;
wire x_3234;
wire x_3235;
wire x_3236;
wire x_3237;
wire x_3238;
wire x_3239;
wire x_3240;
wire x_3241;
wire x_3242;
wire x_3243;
wire x_3244;
wire x_3245;
wire x_3246;
wire x_3247;
wire x_3248;
wire x_3249;
wire x_3250;
wire x_3251;
wire x_3252;
wire x_3253;
wire x_3254;
wire x_3255;
wire x_3256;
wire x_3257;
wire x_3258;
wire x_3259;
wire x_3260;
wire x_3261;
wire x_3262;
wire x_3263;
wire x_3264;
wire x_3265;
wire x_3266;
wire x_3267;
wire x_3268;
wire x_3269;
wire x_3270;
wire x_3271;
wire x_3272;
wire x_3273;
wire x_3274;
wire x_3275;
wire x_3276;
wire x_3277;
wire x_3278;
wire x_3279;
wire x_3280;
wire x_3281;
wire x_3282;
wire x_3283;
wire x_3284;
wire x_3285;
wire x_3286;
wire x_3287;
wire x_3288;
wire x_3289;
wire x_3290;
wire x_3291;
wire x_3292;
wire x_3293;
wire x_3294;
wire x_3295;
wire x_3296;
wire x_3297;
wire x_3298;
wire x_3299;
wire x_3300;
wire x_3301;
wire x_3302;
wire x_3303;
wire x_3304;
wire x_3305;
wire x_3306;
wire x_3307;
wire x_3308;
wire x_3309;
wire x_3310;
wire x_3311;
wire x_3312;
wire x_3313;
wire x_3314;
wire x_3315;
wire x_3316;
wire x_3317;
wire x_3318;
wire x_3319;
wire x_3320;
wire x_3321;
wire x_3322;
wire x_3323;
wire x_3324;
wire x_3325;
wire x_3326;
wire x_3327;
wire x_3328;
wire x_3329;
wire x_3330;
wire x_3331;
wire x_3332;
wire x_3333;
wire x_3334;
wire x_3335;
wire x_3336;
wire x_3337;
wire x_3338;
wire x_3339;
wire x_3340;
wire x_3341;
wire x_3342;
wire x_3343;
wire x_3344;
wire x_3345;
wire x_3346;
wire x_3347;
wire x_3348;
wire x_3349;
wire x_3350;
wire x_3351;
wire x_3352;
wire x_3353;
wire x_3354;
wire x_3355;
wire x_3356;
wire x_3357;
wire x_3358;
wire x_3359;
wire x_3360;
wire x_3361;
wire x_3362;
wire x_3363;
wire x_3364;
wire x_3365;
wire x_3366;
wire x_3367;
wire x_3368;
wire x_3369;
wire x_3370;
wire x_3371;
wire x_3372;
wire x_3373;
wire x_3374;
wire x_3375;
wire x_3376;
wire x_3377;
wire x_3378;
wire x_3379;
wire x_3380;
wire x_3381;
wire x_3382;
wire x_3383;
wire x_3384;
wire x_3385;
wire x_3386;
wire x_3387;
wire x_3388;
wire x_3389;
wire x_3390;
wire x_3391;
wire x_3392;
wire x_3393;
wire x_3394;
wire x_3395;
wire x_3396;
wire x_3397;
wire x_3398;
wire x_3399;
wire x_3400;
wire x_3401;
wire x_3402;
wire x_3403;
wire x_3404;
wire x_3405;
wire x_3406;
wire x_3407;
wire x_3408;
wire x_3409;
wire x_3410;
wire x_3411;
wire x_3412;
wire x_3413;
wire x_3414;
wire x_3415;
wire x_3416;
wire x_3417;
wire x_3418;
wire x_3419;
wire x_3420;
wire x_3421;
wire x_3422;
wire x_3423;
wire x_3424;
wire x_3425;
wire x_3426;
wire x_3427;
wire x_3428;
wire x_3429;
wire x_3430;
wire x_3431;
wire x_3432;
wire x_3433;
wire x_3434;
wire x_3435;
wire x_3436;
wire x_3437;
wire x_3438;
wire x_3439;
wire x_3440;
wire x_3441;
wire x_3442;
wire x_3443;
wire x_3444;
wire x_3445;
wire x_3446;
wire x_3447;
wire x_3448;
wire x_3449;
wire x_3450;
wire x_3451;
wire x_3452;
wire x_3453;
wire x_3454;
wire x_3455;
wire x_3456;
wire x_3457;
wire x_3458;
wire x_3459;
wire x_3460;
wire x_3461;
wire x_3462;
wire x_3463;
wire x_3464;
wire x_3465;
wire x_3466;
wire x_3467;
wire x_3468;
wire x_3469;
wire x_3470;
wire x_3471;
wire x_3472;
wire x_3473;
wire x_3474;
wire x_3475;
wire x_3476;
wire x_3477;
wire x_3478;
wire x_3479;
wire x_3480;
wire x_3481;
wire x_3482;
wire x_3483;
wire x_3484;
wire x_3485;
wire x_3486;
wire x_3487;
wire x_3488;
wire x_3489;
wire x_3490;
wire x_3491;
wire x_3492;
wire x_3493;
wire x_3494;
wire x_3495;
wire x_3496;
wire x_3497;
wire x_3498;
wire x_3499;
wire x_3500;
wire x_3501;
wire x_3502;
wire x_3503;
wire x_3504;
wire x_3505;
wire x_3506;
wire x_3507;
wire x_3508;
wire x_3509;
wire x_3510;
wire x_3511;
wire x_3512;
wire x_3513;
wire x_3514;
wire x_3515;
wire x_3516;
wire x_3517;
wire x_3518;
wire x_3519;
wire x_3520;
wire x_3521;
wire x_3522;
wire x_3523;
wire x_3524;
wire x_3525;
wire x_3526;
wire x_3527;
wire x_3528;
wire x_3529;
wire x_3530;
wire x_3531;
wire x_3532;
wire x_3533;
wire x_3534;
wire x_3535;
wire x_3536;
wire x_3537;
wire x_3538;
wire x_3539;
wire x_3540;
wire x_3541;
wire x_3542;
wire x_3543;
wire x_3544;
wire x_3545;
wire x_3546;
wire x_3547;
wire x_3548;
wire x_3549;
wire x_3550;
wire x_3551;
wire x_3552;
wire x_3553;
wire x_3554;
wire x_3555;
wire x_3556;
wire x_3557;
wire x_3558;
wire x_3559;
wire x_3560;
wire x_3561;
wire x_3562;
wire x_3563;
wire x_3564;
wire x_3565;
wire x_3566;
wire x_3567;
wire x_3568;
wire x_3569;
wire x_3570;
wire x_3571;
wire x_3572;
wire x_3573;
wire x_3574;
wire x_3575;
wire x_3576;
wire x_3577;
wire x_3578;
wire x_3579;
wire x_3580;
wire x_3581;
wire x_3582;
wire x_3583;
wire x_3584;
wire x_3585;
wire x_3586;
wire x_3587;
wire x_3588;
wire x_3589;
wire x_3590;
wire x_3591;
wire x_3592;
wire x_3593;
wire x_3594;
wire x_3595;
wire x_3596;
wire x_3597;
wire x_3598;
wire x_3599;
wire x_3600;
wire x_3601;
wire x_3602;
wire x_3603;
wire x_3604;
wire x_3605;
wire x_3606;
wire x_3607;
wire x_3608;
wire x_3609;
wire x_3610;
wire x_3611;
wire x_3612;
wire x_3613;
wire x_3614;
wire x_3615;
wire x_3616;
wire x_3617;
wire x_3618;
wire x_3619;
wire x_3620;
wire x_3621;
wire x_3622;
wire x_3623;
wire x_3624;
wire x_3625;
wire x_3626;
wire x_3627;
wire x_3628;
wire x_3629;
wire x_3630;
wire x_3631;
wire x_3632;
wire x_3633;
wire x_3634;
wire x_3635;
wire x_3636;
wire x_3637;
wire x_3638;
wire x_3639;
wire x_3640;
wire x_3641;
wire x_3642;
wire x_3643;
wire x_3644;
wire x_3645;
wire x_3646;
wire x_3647;
wire x_3648;
wire x_3649;
wire x_3650;
wire x_3651;
wire x_3652;
wire x_3653;
wire x_3654;
wire x_3655;
wire x_3656;
wire x_3657;
wire x_3658;
wire x_3659;
wire x_3660;
wire x_3661;
wire x_3662;
wire x_3663;
wire x_3664;
wire x_3665;
wire x_3666;
wire x_3667;
wire x_3668;
wire x_3669;
wire x_3670;
wire x_3671;
wire x_3672;
wire x_3673;
wire x_3674;
wire x_3675;
wire x_3676;
wire x_3677;
wire x_3678;
wire x_3679;
wire x_3680;
wire x_3681;
wire x_3682;
wire x_3683;
wire x_3684;
wire x_3685;
wire x_3686;
wire x_3687;
wire x_3688;
wire x_3689;
wire x_3690;
wire x_3691;
wire x_3692;
wire x_3693;
wire x_3694;
wire x_3695;
wire x_3696;
wire x_3697;
wire x_3698;
wire x_3699;
wire x_3700;
wire x_3701;
wire x_3702;
wire x_3703;
wire x_3704;
wire x_3705;
wire x_3706;
wire x_3707;
wire x_3708;
wire x_3709;
wire x_3710;
wire x_3711;
wire x_3712;
wire x_3713;
wire x_3714;
wire x_3715;
wire x_3716;
wire x_3717;
wire x_3718;
wire x_3719;
wire x_3720;
wire x_3721;
wire x_3722;
wire x_3723;
wire x_3724;
wire x_3725;
wire x_3726;
wire x_3727;
wire x_3728;
wire x_3729;
wire x_3730;
wire x_3731;
wire x_3732;
wire x_3733;
wire x_3734;
wire x_3735;
wire x_3736;
wire x_3737;
wire x_3738;
wire x_3739;
wire x_3740;
wire x_3741;
wire x_3742;
wire x_3743;
wire x_3744;
wire x_3745;
wire x_3746;
wire x_3747;
wire x_3748;
wire x_3749;
wire x_3750;
wire x_3751;
wire x_3752;
wire x_3753;
wire x_3754;
wire x_3755;
wire x_3756;
wire x_3757;
wire x_3758;
wire x_3759;
wire x_3760;
wire x_3761;
wire x_3762;
wire x_3763;
wire x_3764;
wire x_3765;
wire x_3766;
wire x_3767;
wire x_3768;
wire x_3769;
wire x_3770;
wire x_3771;
wire x_3772;
wire x_3773;
wire x_3774;
wire x_3775;
wire x_3776;
wire x_3777;
wire x_3778;
wire x_3779;
wire x_3780;
wire x_3781;
wire x_3782;
wire x_3783;
wire x_3784;
wire x_3785;
wire x_3786;
wire x_3787;
wire x_3788;
wire x_3789;
wire x_3790;
wire x_3791;
wire x_3792;
wire x_3793;
wire x_3794;
wire x_3795;
wire x_3796;
wire x_3797;
wire x_3798;
wire x_3799;
wire x_3800;
wire x_3801;
wire x_3802;
wire x_3803;
wire x_3804;
wire x_3805;
wire x_3806;
wire x_3807;
wire x_3808;
wire x_3809;
wire x_3810;
wire x_3811;
wire x_3812;
wire x_3813;
wire x_3814;
wire x_3815;
wire x_3816;
wire x_3817;
wire x_3818;
wire x_3819;
wire x_3820;
wire x_3821;
wire x_3822;
wire x_3823;
wire x_3824;
wire x_3825;
wire x_3826;
wire x_3827;
wire x_3828;
wire x_3829;
wire x_3830;
wire x_3831;
wire x_3832;
wire x_3833;
wire x_3834;
wire x_3835;
wire x_3836;
wire x_3837;
wire x_3838;
wire x_3839;
wire x_3840;
wire x_3841;
wire x_3842;
wire x_3843;
wire x_3844;
wire x_3845;
wire x_3846;
wire x_3847;
wire x_3848;
wire x_3849;
wire x_3850;
wire x_3851;
wire x_3852;
wire x_3853;
wire x_3854;
wire x_3855;
wire x_3856;
wire x_3857;
wire x_3858;
wire x_3859;
wire x_3860;
wire x_3861;
wire x_3862;
wire x_3863;
wire x_3864;
wire x_3865;
wire x_3866;
wire x_3867;
wire x_3868;
wire x_3869;
wire x_3870;
wire x_3871;
wire x_3872;
wire x_3873;
wire x_3874;
wire x_3875;
wire x_3876;
wire x_3877;
wire x_3878;
wire x_3879;
wire x_3880;
wire x_3881;
wire x_3882;
wire x_3883;
wire x_3884;
wire x_3885;
wire x_3886;
wire x_3887;
wire x_3888;
wire x_3889;
wire x_3890;
wire x_3891;
wire x_3892;
wire x_3893;
wire x_3894;
wire x_3895;
wire x_3896;
wire x_3897;
wire x_3898;
wire x_3899;
wire x_3900;
wire x_3901;
wire x_3902;
wire x_3903;
wire x_3904;
wire x_3905;
wire x_3906;
wire x_3907;
wire x_3908;
wire x_3909;
wire x_3910;
wire x_3911;
wire x_3912;
wire x_3913;
wire x_3914;
wire x_3915;
wire x_3916;
wire x_3917;
wire x_3918;
wire x_3919;
wire x_3920;
wire x_3921;
wire x_3922;
wire x_3923;
wire x_3924;
wire x_3925;
wire x_3926;
wire x_3927;
wire x_3928;
wire x_3929;
wire x_3930;
wire x_3931;
wire x_3932;
wire x_3933;
wire x_3934;
wire x_3935;
wire x_3936;
wire x_3937;
wire x_3938;
wire x_3939;
wire x_3940;
wire x_3941;
wire x_3942;
wire x_3943;
wire x_3944;
wire x_3945;
wire x_3946;
wire x_3947;
wire x_3948;
wire x_3949;
wire x_3950;
wire x_3951;
wire x_3952;
wire x_3953;
wire x_3954;
wire x_3955;
wire x_3956;
wire x_3957;
wire x_3958;
wire x_3959;
wire x_3960;
wire x_3961;
wire x_3962;
wire x_3963;
wire x_3964;
wire x_3965;
wire x_3966;
wire x_3967;
wire x_3968;
wire x_3969;
wire x_3970;
wire x_3971;
wire x_3972;
wire x_3973;
wire x_3974;
wire x_3975;
wire x_3976;
wire x_3977;
wire x_3978;
wire x_3979;
wire x_3980;
wire x_3981;
wire x_3982;
wire x_3983;
wire x_3984;
wire x_3985;
wire x_3986;
wire x_3987;
wire x_3988;
wire x_3989;
wire x_3990;
wire x_3991;
wire x_3992;
wire x_3993;
wire x_3994;
wire x_3995;
wire x_3996;
wire x_3997;
wire x_3998;
wire x_3999;
wire x_4000;
wire x_4001;
wire x_4002;
wire x_4003;
wire x_4004;
wire x_4005;
wire x_4006;
wire x_4007;
wire x_4008;
wire x_4009;
wire x_4010;
wire x_4011;
wire x_4012;
wire x_4013;
wire x_4014;
wire x_4015;
wire x_4016;
wire x_4017;
wire x_4018;
wire x_4019;
wire x_4020;
wire x_4021;
wire x_4022;
wire x_4023;
wire x_4024;
wire x_4025;
wire x_4026;
wire x_4027;
wire x_4028;
wire x_4029;
wire x_4030;
wire x_4031;
wire x_4032;
wire x_4033;
wire x_4034;
wire x_4035;
wire x_4036;
wire x_4037;
wire x_4038;
wire x_4039;
wire x_4040;
wire x_4041;
wire x_4042;
wire x_4043;
wire x_4044;
wire x_4045;
wire x_4046;
wire x_4047;
wire x_4048;
wire x_4049;
wire x_4050;
wire x_4051;
wire x_4052;
wire x_4053;
wire x_4054;
wire x_4055;
wire x_4056;
wire x_4057;
wire x_4058;
wire x_4059;
wire x_4060;
wire x_4061;
wire x_4062;
wire x_4063;
wire x_4064;
wire x_4065;
wire x_4066;
wire x_4067;
wire x_4068;
wire x_4069;
wire x_4070;
wire x_4071;
wire x_4072;
wire x_4073;
wire x_4074;
wire x_4075;
wire x_4076;
wire x_4077;
wire x_4078;
wire x_4079;
wire x_4080;
wire x_4081;
wire x_4082;
wire x_4083;
wire x_4084;
wire x_4085;
wire x_4086;
wire x_4087;
wire x_4088;
wire x_4089;
wire x_4090;
wire x_4091;
wire x_4092;
wire x_4093;
wire x_4094;
wire x_4095;
wire x_4096;
wire x_4097;
wire x_4098;
wire x_4099;
wire x_4100;
wire x_4101;
wire x_4102;
wire x_4103;
wire x_4104;
wire x_4105;
wire x_4106;
wire x_4107;
wire x_4108;
wire x_4109;
wire x_4110;
wire x_4111;
wire x_4112;
wire x_4113;
wire x_4114;
wire x_4115;
wire x_4116;
wire x_4117;
wire x_4118;
wire x_4119;
wire x_4120;
wire x_4121;
wire x_4122;
wire x_4123;
wire x_4124;
wire x_4125;
wire x_4126;
wire x_4127;
wire x_4128;
wire x_4129;
wire x_4130;
wire x_4131;
wire x_4132;
wire x_4133;
wire x_4134;
wire x_4135;
wire x_4136;
wire x_4137;
wire x_4138;
wire x_4139;
wire x_4140;
wire x_4141;
wire x_4142;
wire x_4143;
wire x_4144;
wire x_4145;
wire x_4146;
wire x_4147;
wire x_4148;
wire x_4149;
wire x_4150;
wire x_4151;
wire x_4152;
wire x_4153;
wire x_4154;
wire x_4155;
wire x_4156;
wire x_4157;
wire x_4158;
wire x_4159;
wire x_4160;
wire x_4161;
wire x_4162;
wire x_4163;
wire x_4164;
wire x_4165;
wire x_4166;
wire x_4167;
wire x_4168;
wire x_4169;
wire x_4170;
wire x_4171;
wire x_4172;
wire x_4173;
wire x_4174;
wire x_4175;
wire x_4176;
wire x_4177;
wire x_4178;
wire x_4179;
wire x_4180;
wire x_4181;
wire x_4182;
wire x_4183;
wire x_4184;
wire x_4185;
wire x_4186;
wire x_4187;
wire x_4188;
wire x_4189;
wire x_4190;
wire x_4191;
wire x_4192;
wire x_4193;
wire x_4194;
wire x_4195;
wire x_4196;
wire x_4197;
wire x_4198;
wire x_4199;
wire x_4200;
wire x_4201;
wire x_4202;
wire x_4203;
wire x_4204;
wire x_4205;
wire x_4206;
wire x_4207;
wire x_4208;
wire x_4209;
wire x_4210;
wire x_4211;
wire x_4212;
wire x_4213;
wire x_4214;
wire x_4215;
wire x_4216;
wire x_4217;
wire x_4218;
wire x_4219;
wire x_4220;
wire x_4221;
wire x_4222;
wire x_4223;
wire x_4224;
wire x_4225;
wire x_4226;
wire x_4227;
wire x_4228;
wire x_4229;
wire x_4230;
wire x_4231;
wire x_4232;
wire x_4233;
wire x_4234;
wire x_4235;
wire x_4236;
wire x_4237;
wire x_4238;
wire x_4239;
wire x_4240;
wire x_4241;
wire x_4242;
wire x_4243;
wire x_4244;
wire x_4245;
wire x_4246;
wire x_4247;
wire x_4248;
wire x_4249;
wire x_4250;
wire x_4251;
wire x_4252;
wire x_4253;
wire x_4254;
wire x_4255;
wire x_4256;
wire x_4257;
wire x_4258;
wire x_4259;
wire x_4260;
wire x_4261;
wire x_4262;
wire x_4263;
wire x_4264;
wire x_4265;
wire x_4266;
wire x_4267;
wire x_4268;
wire x_4269;
wire x_4270;
wire x_4271;
wire x_4272;
wire x_4273;
wire x_4274;
wire x_4275;
wire x_4276;
wire x_4277;
wire x_4278;
wire x_4279;
wire x_4280;
wire x_4281;
wire x_4282;
wire x_4283;
wire x_4284;
wire x_4285;
wire x_4286;
wire x_4287;
wire x_4288;
wire x_4289;
wire x_4290;
wire x_4291;
wire x_4292;
wire x_4293;
wire x_4294;
wire x_4295;
wire x_4296;
wire x_4297;
wire x_4298;
wire x_4299;
wire x_4300;
wire x_4301;
wire x_4302;
wire x_4303;
wire x_4304;
wire x_4305;
wire x_4306;
wire x_4307;
wire x_4308;
wire x_4309;
wire x_4310;
wire x_4311;
wire x_4312;
wire x_4313;
wire x_4314;
wire x_4315;
wire x_4316;
wire x_4317;
wire x_4318;
wire x_4319;
wire x_4320;
wire x_4321;
wire x_4322;
wire x_4323;
wire x_4324;
wire x_4325;
wire x_4326;
wire x_4327;
wire x_4328;
wire x_4329;
wire x_4330;
wire x_4331;
wire x_4332;
wire x_4333;
wire x_4334;
wire x_4335;
wire x_4336;
wire x_4337;
wire x_4338;
wire x_4339;
wire x_4340;
wire x_4341;
wire x_4342;
wire x_4343;
wire x_4344;
wire x_4345;
wire x_4346;
wire x_4347;
wire x_4348;
wire x_4349;
wire x_4350;
wire x_4351;
wire x_4352;
wire x_4353;
wire x_4354;
wire x_4355;
wire x_4356;
wire x_4357;
wire x_4358;
wire x_4359;
wire x_4360;
wire x_4361;
wire x_4362;
wire x_4363;
wire x_4364;
wire x_4365;
wire x_4366;
wire x_4367;
wire x_4368;
wire x_4369;
wire x_4370;
wire x_4371;
wire x_4372;
wire x_4373;
wire x_4374;
wire x_4375;
wire x_4376;
wire x_4377;
wire x_4378;
wire x_4379;
wire x_4380;
wire x_4381;
wire x_4382;
wire x_4383;
wire x_4384;
wire x_4385;
wire x_4386;
wire x_4387;
wire x_4388;
wire x_4389;
wire x_4390;
wire x_4391;
wire x_4392;
wire x_4393;
wire x_4394;
wire x_4395;
wire x_4396;
wire x_4397;
wire x_4398;
wire x_4399;
wire x_4400;
wire x_4401;
wire x_4402;
wire x_4403;
wire x_4404;
wire x_4405;
wire x_4406;
wire x_4407;
wire x_4408;
wire x_4409;
wire x_4410;
wire x_4411;
wire x_4412;
wire x_4413;
wire x_4414;
wire x_4415;
wire x_4416;
wire x_4417;
wire x_4418;
wire x_4419;
wire x_4420;
wire x_4421;
wire x_4422;
wire x_4423;
wire x_4424;
wire x_4425;
wire x_4426;
wire x_4427;
wire x_4428;
wire x_4429;
wire x_4430;
wire x_4431;
wire x_4432;
wire x_4433;
wire x_4434;
wire x_4435;
wire x_4436;
wire x_4437;
wire x_4438;
wire x_4439;
wire x_4440;
wire x_4441;
wire x_4442;
wire x_4443;
wire x_4444;
wire x_4445;
wire x_4446;
wire x_4447;
wire x_4448;
wire x_4449;
wire x_4450;
wire x_4451;
wire x_4452;
wire x_4453;
wire x_4454;
wire x_4455;
wire x_4456;
wire x_4457;
wire x_4458;
wire x_4459;
wire x_4460;
wire x_4461;
wire x_4462;
wire x_4463;
wire x_4464;
wire x_4465;
wire x_4466;
wire x_4467;
wire x_4468;
wire x_4469;
wire x_4470;
wire x_4471;
wire x_4472;
wire x_4473;
wire x_4474;
wire x_4475;
wire x_4476;
wire x_4477;
wire x_4478;
wire x_4479;
wire x_4480;
wire x_4481;
wire x_4482;
wire x_4483;
wire x_4484;
wire x_4485;
wire x_4486;
wire x_4487;
wire x_4488;
wire x_4489;
wire x_4490;
wire x_4491;
wire x_4492;
wire x_4493;
wire x_4494;
wire x_4495;
wire x_4496;
wire x_4497;
wire x_4498;
wire x_4499;
wire x_4500;
wire x_4501;
wire x_4502;
wire x_4503;
wire x_4504;
wire x_4505;
wire x_4506;
wire x_4507;
wire x_4508;
wire x_4509;
wire x_4510;
wire x_4511;
wire x_4512;
wire x_4513;
wire x_4514;
wire x_4515;
wire x_4516;
wire x_4517;
wire x_4518;
wire x_4519;
wire x_4520;
wire x_4521;
wire x_4522;
wire x_4523;
wire x_4524;
wire x_4525;
wire x_4526;
wire x_4527;
wire x_4528;
wire x_4529;
wire x_4530;
wire x_4531;
wire x_4532;
wire x_4533;
wire x_4534;
wire x_4535;
wire x_4536;
wire x_4537;
wire x_4538;
wire x_4539;
wire x_4540;
wire x_4541;
wire x_4542;
wire x_4543;
wire x_4544;
wire x_4545;
wire x_4546;
wire x_4547;
wire x_4548;
wire x_4549;
wire x_4550;
wire x_4551;
wire x_4552;
wire x_4553;
wire x_4554;
wire x_4555;
wire x_4556;
wire x_4557;
wire x_4558;
wire x_4559;
wire x_4560;
wire x_4561;
wire x_4562;
wire x_4563;
wire x_4564;
wire x_4565;
wire x_4566;
wire x_4567;
wire x_4568;
wire x_4569;
wire x_4570;
wire x_4571;
wire x_4572;
wire x_4573;
wire x_4574;
wire x_4575;
wire x_4576;
wire x_4577;
wire x_4578;
wire x_4579;
wire x_4580;
wire x_4581;
wire x_4582;
wire x_4583;
wire x_4584;
wire x_4585;
wire x_4586;
wire x_4587;
wire x_4588;
wire x_4589;
wire x_4590;
wire x_4591;
wire x_4592;
wire x_4593;
wire x_4594;
wire x_4595;
wire x_4596;
wire x_4597;
wire x_4598;
wire x_4599;
wire x_4600;
wire x_4601;
wire x_4602;
wire x_4603;
wire x_4604;
wire x_4605;
wire x_4606;
wire x_4607;
wire x_4608;
wire x_4609;
wire x_4610;
wire x_4611;
wire x_4612;
wire x_4613;
wire x_4614;
wire x_4615;
wire x_4616;
wire x_4617;
wire x_4618;
wire x_4619;
wire x_4620;
wire x_4621;
wire x_4622;
wire x_4623;
wire x_4624;
wire x_4625;
wire x_4626;
wire x_4627;
wire x_4628;
wire x_4629;
wire x_4630;
wire x_4631;
wire x_4632;
wire x_4633;
wire x_4634;
wire x_4635;
wire x_4636;
wire x_4637;
wire x_4638;
wire x_4639;
wire x_4640;
wire x_4641;
wire x_4642;
wire x_4643;
wire x_4644;
wire x_4645;
wire x_4646;
wire x_4647;
wire x_4648;
wire x_4649;
wire x_4650;
wire x_4651;
wire x_4652;
wire x_4653;
wire x_4654;
wire x_4655;
wire x_4656;
wire x_4657;
wire x_4658;
wire x_4659;
wire x_4660;
wire x_4661;
wire x_4662;
wire x_4663;
wire x_4664;
wire x_4665;
wire x_4666;
wire x_4667;
wire x_4668;
wire x_4669;
wire x_4670;
wire x_4671;
wire x_4672;
wire x_4673;
wire x_4674;
wire x_4675;
wire x_4676;
wire x_4677;
wire x_4678;
wire x_4679;
wire x_4680;
wire x_4681;
wire x_4682;
wire x_4683;
wire x_4684;
wire x_4685;
wire x_4686;
wire x_4687;
wire x_4688;
wire x_4689;
wire x_4690;
wire x_4691;
wire x_4692;
wire x_4693;
wire x_4694;
wire x_4695;
wire x_4696;
wire x_4697;
wire x_4698;
wire x_4699;
wire x_4700;
wire x_4701;
wire x_4702;
wire x_4703;
wire x_4704;
wire x_4705;
wire x_4706;
wire x_4707;
wire x_4708;
wire x_4709;
wire x_4710;
wire x_4711;
wire x_4712;
wire x_4713;
wire x_4714;
wire x_4715;
wire x_4716;
wire x_4717;
wire x_4718;
wire x_4719;
wire x_4720;
wire x_4721;
wire x_4722;
wire x_4723;
wire x_4724;
wire x_4725;
wire x_4726;
wire x_4727;
wire x_4728;
wire x_4729;
wire x_4730;
wire x_4731;
wire x_4732;
wire x_4733;
wire x_4734;
wire x_4735;
wire x_4736;
wire x_4737;
wire x_4738;
wire x_4739;
wire x_4740;
wire x_4741;
wire x_4742;
wire x_4743;
wire x_4744;
wire x_4745;
wire x_4746;
wire x_4747;
wire x_4748;
wire x_4749;
wire x_4750;
wire x_4751;
wire x_4752;
wire x_4753;
wire x_4754;
wire x_4755;
wire x_4756;
wire x_4757;
wire x_4758;
wire x_4759;
wire x_4760;
wire x_4761;
wire x_4762;
wire x_4763;
wire x_4764;
wire x_4765;
wire x_4766;
wire x_4767;
wire x_4768;
wire x_4769;
wire x_4770;
wire x_4771;
wire x_4772;
wire x_4773;
wire x_4774;
wire x_4775;
wire x_4776;
wire x_4777;
wire x_4778;
wire x_4779;
wire x_4780;
wire x_4781;
wire x_4782;
wire x_4783;
wire x_4784;
wire x_4785;
wire x_4786;
wire x_4787;
wire x_4788;
wire x_4789;
wire x_4790;
wire x_4791;
wire x_4792;
wire x_4793;
wire x_4794;
wire x_4795;
wire x_4796;
wire x_4797;
wire x_4798;
wire x_4799;
wire x_4800;
wire x_4801;
wire x_4802;
wire x_4803;
wire x_4804;
wire x_4805;
wire x_4806;
wire x_4807;
wire x_4808;
wire x_4809;
wire x_4810;
wire x_4811;
wire x_4812;
wire x_4813;
wire x_4814;
wire x_4815;
wire x_4816;
wire x_4817;
wire x_4818;
wire x_4819;
wire x_4820;
wire x_4821;
wire x_4822;
wire x_4823;
wire x_4824;
wire x_4825;
wire x_4826;
wire x_4827;
wire x_4828;
wire x_4829;
wire x_4830;
wire x_4831;
wire x_4832;
wire x_4833;
wire x_4834;
wire x_4835;
wire x_4836;
wire x_4837;
wire x_4838;
wire x_4839;
wire x_4840;
wire x_4841;
wire x_4842;
wire x_4843;
wire x_4844;
wire x_4845;
wire x_4846;
wire x_4847;
wire x_4848;
wire x_4849;
wire x_4850;
wire x_4851;
wire x_4852;
wire x_4853;
wire x_4854;
wire x_4855;
wire x_4856;
wire x_4857;
wire x_4858;
wire x_4859;
wire x_4860;
wire x_4861;
wire x_4862;
wire x_4863;
wire x_4864;
wire x_4865;
wire x_4866;
wire x_4867;
wire x_4868;
wire x_4869;
wire x_4870;
wire x_4871;
wire x_4872;
wire x_4873;
wire x_4874;
wire x_4875;
wire x_4876;
wire x_4877;
wire x_4878;
wire x_4879;
wire x_4880;
wire x_4881;
wire x_4882;
wire x_4883;
wire x_4884;
wire x_4885;
wire x_4886;
wire x_4887;
wire x_4888;
wire x_4889;
wire x_4890;
wire x_4891;
wire x_4892;
wire x_4893;
wire x_4894;
wire x_4895;
wire x_4896;
wire x_4897;
wire x_4898;
wire x_4899;
wire x_4900;
wire x_4901;
wire x_4902;
wire x_4903;
wire x_4904;
wire x_4905;
wire x_4906;
wire x_4907;
wire x_4908;
wire x_4909;
wire x_4910;
wire x_4911;
wire x_4912;
wire x_4913;
wire x_4914;
wire x_4915;
wire x_4916;
wire x_4917;
wire x_4918;
wire x_4919;
wire x_4920;
wire x_4921;
wire x_4922;
wire x_4923;
wire x_4924;
wire x_4925;
wire x_4926;
wire x_4927;
wire x_4928;
wire x_4929;
wire x_4930;
wire x_4931;
wire x_4932;
wire x_4933;
wire x_4934;
wire x_4935;
wire x_4936;
wire x_4937;
wire x_4938;
wire x_4939;
wire x_4940;
wire x_4941;
wire x_4942;
wire x_4943;
wire x_4944;
wire x_4945;
wire x_4946;
wire x_4947;
wire x_4948;
wire x_4949;
wire x_4950;
wire x_4951;
wire x_4952;
wire x_4953;
wire x_4954;
wire x_4955;
wire x_4956;
wire x_4957;
wire x_4958;
wire x_4959;
wire x_4960;
wire x_4961;
wire x_4962;
wire x_4963;
wire x_4964;
wire x_4965;
wire x_4966;
wire x_4967;
wire x_4968;
wire x_4969;
wire x_4970;
wire x_4971;
wire x_4972;
wire x_4973;
wire x_4974;
wire x_4975;
wire x_4976;
wire x_4977;
wire x_4978;
wire x_4979;
wire x_4980;
wire x_4981;
wire x_4982;
wire x_4983;
wire x_4984;
wire x_4985;
wire x_4986;
wire x_4987;
wire x_4988;
wire x_4989;
wire x_4990;
wire x_4991;
wire x_4992;
wire x_4993;
wire x_4994;
wire x_4995;
wire x_4996;
wire x_4997;
wire x_4998;
wire x_4999;
wire x_5000;
wire x_5001;
wire x_5002;
wire x_5003;
wire x_5004;
wire x_5005;
wire x_5006;
wire x_5007;
wire x_5008;
wire x_5009;
wire x_5010;
wire x_5011;
wire x_5012;
wire x_5013;
wire x_5014;
wire x_5015;
wire x_5016;
wire x_5017;
wire x_5018;
wire x_5019;
wire x_5020;
wire x_5021;
wire x_5022;
wire x_5023;
wire x_5024;
wire x_5025;
wire x_5026;
wire x_5027;
wire x_5028;
wire x_5029;
wire x_5030;
wire x_5031;
wire x_5032;
wire x_5033;
wire x_5034;
wire x_5035;
wire x_5036;
wire x_5037;
wire x_5038;
wire x_5039;
wire x_5040;
wire x_5041;
wire x_5042;
wire x_5043;
wire x_5044;
wire x_5045;
wire x_5046;
wire x_5047;
wire x_5048;
wire x_5049;
wire x_5050;
wire x_5051;
wire x_5052;
wire x_5053;
wire x_5054;
wire x_5055;
wire x_5056;
wire x_5057;
wire x_5058;
wire x_5059;
wire x_5060;
wire x_5061;
wire x_5062;
wire x_5063;
wire x_5064;
wire x_5065;
wire x_5066;
wire x_5067;
wire x_5068;
wire x_5069;
wire x_5070;
wire x_5071;
wire x_5072;
wire x_5073;
wire x_5074;
wire x_5075;
wire x_5076;
wire x_5077;
wire x_5078;
wire x_5079;
wire x_5080;
wire x_5081;
wire x_5082;
wire x_5083;
wire x_5084;
wire x_5085;
wire x_5086;
wire x_5087;
wire x_5088;
wire x_5089;
wire x_5090;
wire x_5091;
wire x_5092;
wire x_5093;
wire x_5094;
wire x_5095;
wire x_5096;
wire x_5097;
wire x_5098;
wire x_5099;
wire x_5100;
wire x_5101;
wire x_5102;
wire x_5103;
wire x_5104;
wire x_5105;
wire x_5106;
wire x_5107;
wire x_5108;
wire x_5109;
wire x_5110;
wire x_5111;
wire x_5112;
wire x_5113;
wire x_5114;
wire x_5115;
wire x_5116;
wire x_5117;
wire x_5118;
wire x_5119;
wire x_5120;
wire x_5121;
wire x_5122;
wire x_5123;
wire x_5124;
wire x_5125;
wire x_5126;
wire x_5127;
wire x_5128;
wire x_5129;
wire x_5130;
wire x_5131;
wire x_5132;
wire x_5133;
wire x_5134;
wire x_5135;
wire x_5136;
wire x_5137;
wire x_5138;
wire x_5139;
wire x_5140;
wire x_5141;
wire x_5142;
wire x_5143;
wire x_5144;
wire x_5145;
wire x_5146;
wire x_5147;
wire x_5148;
wire x_5149;
wire x_5150;
wire x_5151;
wire x_5152;
wire x_5153;
wire x_5154;
wire x_5155;
wire x_5156;
wire x_5157;
wire x_5158;
wire x_5159;
wire x_5160;
wire x_5161;
wire x_5162;
wire x_5163;
wire x_5164;
wire x_5165;
wire x_5166;
wire x_5167;
wire x_5168;
wire x_5169;
wire x_5170;
wire x_5171;
wire x_5172;
wire x_5173;
wire x_5174;
wire x_5175;
wire x_5176;
wire x_5177;
wire x_5178;
wire x_5179;
wire x_5180;
wire x_5181;
wire x_5182;
wire x_5183;
wire x_5184;
wire x_5185;
wire x_5186;
wire x_5187;
wire x_5188;
wire x_5189;
wire x_5190;
wire x_5191;
wire x_5192;
wire x_5193;
wire x_5194;
wire x_5195;
wire x_5196;
wire x_5197;
wire x_5198;
wire x_5199;
wire x_5200;
wire x_5201;
wire x_5202;
wire x_5203;
wire x_5204;
wire x_5205;
wire x_5206;
wire x_5207;
wire x_5208;
wire x_5209;
wire x_5210;
wire x_5211;
wire x_5212;
wire x_5213;
wire x_5214;
wire x_5215;
wire x_5216;
wire x_5217;
wire x_5218;
wire x_5219;
wire x_5220;
wire x_5221;
wire x_5222;
wire x_5223;
wire x_5224;
wire x_5225;
wire x_5226;
wire x_5227;
wire x_5228;
wire x_5229;
wire x_5230;
wire x_5231;
wire x_5232;
wire x_5233;
wire x_5234;
wire x_5235;
wire x_5236;
wire x_5237;
wire x_5238;
wire x_5239;
wire x_5240;
wire x_5241;
wire x_5242;
wire x_5243;
wire x_5244;
wire x_5245;
wire x_5246;
wire x_5247;
wire x_5248;
wire x_5249;
wire x_5250;
wire x_5251;
wire x_5252;
wire x_5253;
wire x_5254;
wire x_5255;
wire x_5256;
wire x_5257;
wire x_5258;
wire x_5259;
wire x_5260;
wire x_5261;
wire x_5262;
wire x_5263;
wire x_5264;
wire x_5265;
wire x_5266;
wire x_5267;
wire x_5268;
wire x_5269;
wire x_5270;
wire x_5271;
wire x_5272;
wire x_5273;
wire x_5274;
wire x_5275;
wire x_5276;
wire x_5277;
wire x_5278;
wire x_5279;
wire x_5280;
wire x_5281;
wire x_5282;
wire x_5283;
wire x_5284;
wire x_5285;
wire x_5286;
wire x_5287;
wire x_5288;
wire x_5289;
wire x_5290;
wire x_5291;
wire x_5292;
wire x_5293;
wire x_5294;
wire x_5295;
wire x_5296;
wire x_5297;
wire x_5298;
wire x_5299;
wire x_5300;
wire x_5301;
wire x_5302;
wire x_5303;
wire x_5304;
wire x_5305;
wire x_5306;
wire x_5307;
wire x_5308;
wire x_5309;
wire x_5310;
wire x_5311;
wire x_5312;
wire x_5313;
wire x_5314;
wire x_5315;
wire x_5316;
wire x_5317;
wire x_5318;
wire x_5319;
wire x_5320;
wire x_5321;
wire x_5322;
wire x_5323;
wire x_5324;
wire x_5325;
wire x_5326;
wire x_5327;
wire x_5328;
wire x_5329;
wire x_5330;
wire x_5331;
wire x_5332;
wire x_5333;
wire x_5334;
wire x_5335;
wire x_5336;
wire x_5337;
wire x_5338;
wire x_5339;
wire x_5340;
wire x_5341;
wire x_5342;
wire x_5343;
wire x_5344;
wire x_5345;
wire x_5346;
wire x_5347;
wire x_5348;
wire x_5349;
wire x_5350;
wire x_5351;
wire x_5352;
wire x_5353;
wire x_5354;
wire x_5355;
wire x_5356;
wire x_5357;
wire x_5358;
wire x_5359;
wire x_5360;
wire x_5361;
wire x_5362;
wire x_5363;
wire x_5364;
wire x_5365;
wire x_5366;
wire x_5367;
wire x_5368;
wire x_5369;
wire x_5370;
wire x_5371;
wire x_5372;
wire x_5373;
wire x_5374;
wire x_5375;
wire x_5376;
wire x_5377;
wire x_5378;
wire x_5379;
wire x_5380;
wire x_5381;
wire x_5382;
wire x_5383;
wire x_5384;
wire x_5385;
wire x_5386;
wire x_5387;
wire x_5388;
wire x_5389;
wire x_5390;
wire x_5391;
wire x_5392;
wire x_5393;
wire x_5394;
wire x_5395;
wire x_5396;
wire x_5397;
wire x_5398;
wire x_5399;
wire x_5400;
wire x_5401;
wire x_5402;
wire x_5403;
wire x_5404;
wire x_5405;
wire x_5406;
wire x_5407;
wire x_5408;
wire x_5409;
wire x_5410;
wire x_5411;
wire x_5412;
wire x_5413;
wire x_5414;
wire x_5415;
wire x_5416;
wire x_5417;
wire x_5418;
wire x_5419;
wire x_5420;
wire x_5421;
wire x_5422;
wire x_5423;
wire x_5424;
wire x_5425;
wire x_5426;
wire x_5427;
wire x_5428;
wire x_5429;
wire x_5430;
wire x_5431;
wire x_5432;
wire x_5433;
wire x_5434;
wire x_5435;
wire x_5436;
wire x_5437;
wire x_5438;
wire x_5439;
wire x_5440;
wire x_5441;
wire x_5442;
wire x_5443;
wire x_5444;
wire x_5445;
wire x_5446;
wire x_5447;
wire x_5448;
wire x_5449;
wire x_5450;
wire x_5451;
wire x_5452;
wire x_5453;
wire x_5454;
wire x_5455;
wire x_5456;
wire x_5457;
wire x_5458;
wire x_5459;
wire x_5460;
wire x_5461;
wire x_5462;
wire x_5463;
wire x_5464;
wire x_5465;
wire x_5466;
wire x_5467;
wire x_5468;
wire x_5469;
wire x_5470;
wire x_5471;
wire x_5472;
wire x_5473;
wire x_5474;
wire x_5475;
wire x_5476;
wire x_5477;
wire x_5478;
wire x_5479;
wire x_5480;
wire x_5481;
wire x_5482;
wire x_5483;
wire x_5484;
wire x_5485;
wire x_5486;
wire x_5487;
wire x_5488;
wire x_5489;
wire x_5490;
wire x_5491;
wire x_5492;
wire x_5493;
wire x_5494;
wire x_5495;
wire x_5496;
wire x_5497;
wire x_5498;
wire x_5499;
wire x_5500;
wire x_5501;
wire x_5502;
wire x_5503;
wire x_5504;
wire x_5505;
wire x_5506;
wire x_5507;
wire x_5508;
wire x_5509;
wire x_5510;
wire x_5511;
wire x_5512;
wire x_5513;
wire x_5514;
wire x_5515;
wire x_5516;
wire x_5517;
wire x_5518;
wire x_5519;
wire x_5520;
wire x_5521;
wire x_5522;
wire x_5523;
wire x_5524;
wire x_5525;
wire x_5526;
wire x_5527;
wire x_5528;
wire x_5529;
wire x_5530;
wire x_5531;
wire x_5532;
wire x_5533;
wire x_5534;
wire x_5535;
wire x_5536;
wire x_5537;
wire x_5538;
wire x_5539;
wire x_5540;
wire x_5541;
wire x_5542;
wire x_5543;
wire x_5544;
wire x_5545;
wire x_5546;
wire x_5547;
wire x_5548;
wire x_5549;
wire x_5550;
wire x_5551;
wire x_5552;
wire x_5553;
wire x_5554;
wire x_5555;
wire x_5556;
wire x_5557;
wire x_5558;
wire x_5559;
wire x_5560;
wire x_5561;
wire x_5562;
wire x_5563;
wire x_5564;
wire x_5565;
wire x_5566;
wire x_5567;
wire x_5568;
wire x_5569;
wire x_5570;
wire x_5571;
wire x_5572;
wire x_5573;
wire x_5574;
wire x_5575;
wire x_5576;
wire x_5577;
wire x_5578;
wire x_5579;
wire x_5580;
wire x_5581;
wire x_5582;
wire x_5583;
wire x_5584;
wire x_5585;
wire x_5586;
wire x_5587;
wire x_5588;
wire x_5589;
wire x_5590;
wire x_5591;
wire x_5592;
wire x_5593;
wire x_5594;
wire x_5595;
wire x_5596;
wire x_5597;
wire x_5598;
wire x_5599;
wire x_5600;
wire x_5601;
wire x_5602;
wire x_5603;
wire x_5604;
wire x_5605;
wire x_5606;
wire x_5607;
wire x_5608;
wire x_5609;
wire x_5610;
wire x_5611;
wire x_5612;
wire x_5613;
wire x_5614;
wire x_5615;
wire x_5616;
wire x_5617;
wire x_5618;
wire x_5619;
wire x_5620;
wire x_5621;
wire x_5622;
wire x_5623;
wire x_5624;
wire x_5625;
wire x_5626;
wire x_5627;
wire x_5628;
wire x_5629;
wire x_5630;
wire x_5631;
wire x_5632;
wire x_5633;
wire x_5634;
wire x_5635;
wire x_5636;
wire x_5637;
wire x_5638;
wire x_5639;
wire x_5640;
wire x_5641;
wire x_5642;
wire x_5643;
wire x_5644;
wire x_5645;
wire x_5646;
wire x_5647;
wire x_5648;
wire x_5649;
wire x_5650;
wire x_5651;
wire x_5652;
wire x_5653;
wire x_5654;
wire x_5655;
wire x_5656;
wire x_5657;
wire x_5658;
wire x_5659;
wire x_5660;
wire x_5661;
wire x_5662;
wire x_5663;
wire x_5664;
wire x_5665;
wire x_5666;
wire x_5667;
wire x_5668;
wire x_5669;
wire x_5670;
wire x_5671;
wire x_5672;
wire x_5673;
wire x_5674;
wire x_5675;
wire x_5676;
wire x_5677;
wire x_5678;
wire x_5679;
wire x_5680;
wire x_5681;
wire x_5682;
wire x_5683;
wire x_5684;
wire x_5685;
wire x_5686;
wire x_5687;
wire x_5688;
wire x_5689;
wire x_5690;
wire x_5691;
wire x_5692;
wire x_5693;
wire x_5694;
wire x_5695;
wire x_5696;
wire x_5697;
wire x_5698;
wire x_5699;
wire x_5700;
wire x_5701;
wire x_5702;
wire x_5703;
wire x_5704;
wire x_5705;
wire x_5706;
wire x_5707;
wire x_5708;
wire x_5709;
wire x_5710;
wire x_5711;
wire x_5712;
wire x_5713;
wire x_5714;
wire x_5715;
wire x_5716;
wire x_5717;
wire x_5718;
wire x_5719;
wire x_5720;
wire x_5721;
wire x_5722;
wire x_5723;
wire x_5724;
wire x_5725;
wire x_5726;
wire x_5727;
wire x_5728;
wire x_5729;
wire x_5730;
wire x_5731;
wire x_5732;
wire x_5733;
wire x_5734;
wire x_5735;
wire x_5736;
wire x_5737;
wire x_5738;
wire x_5739;
wire x_5740;
wire x_5741;
wire x_5742;
wire x_5743;
wire x_5744;
wire x_5745;
wire x_5746;
wire x_5747;
wire x_5748;
wire x_5749;
wire x_5750;
wire x_5751;
wire x_5752;
wire x_5753;
wire x_5754;
wire x_5755;
wire x_5756;
wire x_5757;
wire x_5758;
wire x_5759;
wire x_5760;
wire x_5761;
wire x_5762;
wire x_5763;
wire x_5764;
wire x_5765;
wire x_5766;
wire x_5767;
wire x_5768;
wire x_5769;
wire x_5770;
wire x_5771;
wire x_5772;
wire x_5773;
wire x_5774;
wire x_5775;
wire x_5776;
wire x_5777;
wire x_5778;
wire x_5779;
wire x_5780;
wire x_5781;
wire x_5782;
wire x_5783;
wire x_5784;
wire x_5785;
wire x_5786;
wire x_5787;
wire x_5788;
wire x_5789;
wire x_5790;
wire x_5791;
wire x_5792;
wire x_5793;
wire x_5794;
wire x_5795;
wire x_5796;
wire x_5797;
wire x_5798;
wire x_5799;
wire x_5800;
wire x_5801;
wire x_5802;
wire x_5803;
wire x_5804;
wire x_5805;
wire x_5806;
wire x_5807;
wire x_5808;
wire x_5809;
wire x_5810;
wire x_5811;
wire x_5812;
wire x_5813;
wire x_5814;
wire x_5815;
wire x_5816;
wire x_5817;
wire x_5818;
wire x_5819;
wire x_5820;
wire x_5821;
wire x_5822;
wire x_5823;
wire x_5824;
wire x_5825;
wire x_5826;
wire x_5827;
wire x_5828;
wire x_5829;
wire x_5830;
wire x_5831;
wire x_5832;
wire x_5833;
wire x_5834;
wire x_5835;
wire x_5836;
wire x_5837;
wire x_5838;
wire x_5839;
wire x_5840;
wire x_5841;
wire x_5842;
wire x_5843;
wire x_5844;
wire x_5845;
wire x_5846;
wire x_5847;
wire x_5848;
wire x_5849;
wire x_5850;
wire x_5851;
wire x_5852;
wire x_5853;
wire x_5854;
wire x_5855;
wire x_5856;
wire x_5857;
wire x_5858;
wire x_5859;
wire x_5860;
wire x_5861;
wire x_5862;
wire x_5863;
wire x_5864;
wire x_5865;
wire x_5866;
wire x_5867;
wire x_5868;
wire x_5869;
wire x_5870;
wire x_5871;
wire x_5872;
wire x_5873;
wire x_5874;
wire x_5875;
wire x_5876;
wire x_5877;
wire x_5878;
wire x_5879;
wire x_5880;
wire x_5881;
wire x_5882;
wire x_5883;
wire x_5884;
wire x_5885;
wire x_5886;
wire x_5887;
wire x_5888;
wire x_5889;
wire x_5890;
wire x_5891;
wire x_5892;
wire x_5893;
wire x_5894;
wire x_5895;
wire x_5896;
wire x_5897;
wire x_5898;
wire x_5899;
wire x_5900;
wire x_5901;
wire x_5902;
wire x_5903;
wire x_5904;
wire x_5905;
wire x_5906;
wire x_5907;
wire x_5908;
wire x_5909;
wire x_5910;
wire x_5911;
wire x_5912;
wire x_5913;
wire x_5914;
wire x_5915;
wire x_5916;
wire x_5917;
wire x_5918;
wire x_5919;
wire x_5920;
wire x_5921;
wire x_5922;
wire x_5923;
wire x_5924;
wire x_5925;
wire x_5926;
wire x_5927;
wire x_5928;
wire x_5929;
wire x_5930;
wire x_5931;
wire x_5932;
wire x_5933;
wire x_5934;
wire x_5935;
wire x_5936;
wire x_5937;
wire x_5938;
wire x_5939;
wire x_5940;
wire x_5941;
wire x_5942;
wire x_5943;
wire x_5944;
wire x_5945;
wire x_5946;
wire x_5947;
wire x_5948;
wire x_5949;
wire x_5950;
wire x_5951;
wire x_5952;
wire x_5953;
wire x_5954;
wire x_5955;
wire x_5956;
wire x_5957;
wire x_5958;
wire x_5959;
wire x_5960;
wire x_5961;
wire x_5962;
wire x_5963;
wire x_5964;
wire x_5965;
wire x_5966;
wire x_5967;
wire x_5968;
wire x_5969;
wire x_5970;
wire x_5971;
wire x_5972;
wire x_5973;
wire x_5974;
wire x_5975;
wire x_5976;
wire x_5977;
wire x_5978;
wire x_5979;
wire x_5980;
wire x_5981;
wire x_5982;
wire x_5983;
wire x_5984;
wire x_5985;
wire x_5986;
wire x_5987;
wire x_5988;
wire x_5989;
wire x_5990;
wire x_5991;
wire x_5992;
wire x_5993;
wire x_5994;
wire x_5995;
wire x_5996;
wire x_5997;
wire x_5998;
wire x_5999;
wire x_6000;
wire x_6001;
wire x_6002;
wire x_6003;
wire x_6004;
wire x_6005;
wire x_6006;
wire x_6007;
wire x_6008;
wire x_6009;
wire x_6010;
wire x_6011;
wire x_6012;
wire x_6013;
wire x_6014;
wire x_6015;
wire x_6016;
wire x_6017;
wire x_6018;
wire x_6019;
wire x_6020;
wire x_6021;
wire x_6022;
wire x_6023;
wire x_6024;
wire x_6025;
wire x_6026;
wire x_6027;
wire x_6028;
wire x_6029;
wire x_6030;
wire x_6031;
wire x_6032;
wire x_6033;
wire x_6034;
wire x_6035;
wire x_6036;
wire x_6037;
wire x_6038;
wire x_6039;
wire x_6040;
wire x_6041;
wire x_6042;
wire x_6043;
wire x_6044;
wire x_6045;
wire x_6046;
wire x_6047;
wire x_6048;
wire x_6049;
wire x_6050;
wire x_6051;
wire x_6052;
wire x_6053;
wire x_6054;
wire x_6055;
wire x_6056;
wire x_6057;
wire x_6058;
wire x_6059;
wire x_6060;
wire x_6061;
wire x_6062;
wire x_6063;
wire x_6064;
wire x_6065;
wire x_6066;
wire x_6067;
wire x_6068;
wire x_6069;
wire x_6070;
wire x_6071;
wire x_6072;
wire x_6073;
wire x_6074;
wire x_6075;
wire x_6076;
wire x_6077;
wire x_6078;
wire x_6079;
wire x_6080;
wire x_6081;
wire x_6082;
wire x_6083;
wire x_6084;
wire x_6085;
wire x_6086;
wire x_6087;
wire x_6088;
wire x_6089;
wire x_6090;
wire x_6091;
wire x_6092;
wire x_6093;
wire x_6094;
wire x_6095;
wire x_6096;
wire x_6097;
wire x_6098;
wire x_6099;
wire x_6100;
wire x_6101;
wire x_6102;
wire x_6103;
wire x_6104;
wire x_6105;
wire x_6106;
wire x_6107;
wire x_6108;
wire x_6109;
wire x_6110;
wire x_6111;
wire x_6112;
wire x_6113;
wire x_6114;
wire x_6115;
wire x_6116;
wire x_6117;
wire x_6118;
wire x_6119;
wire x_6120;
wire x_6121;
wire x_6122;
wire x_6123;
wire x_6124;
wire x_6125;
wire x_6126;
wire x_6127;
wire x_6128;
wire x_6129;
wire x_6130;
wire x_6131;
wire x_6132;
wire x_6133;
wire x_6134;
wire x_6135;
wire x_6136;
wire x_6137;
wire x_6138;
wire x_6139;
wire x_6140;
wire x_6141;
wire x_6142;
wire x_6143;
wire x_6144;
wire x_6145;
wire x_6146;
wire x_6147;
wire x_6148;
wire x_6149;
wire x_6150;
wire x_6151;
wire x_6152;
wire x_6153;
wire x_6154;
wire x_6155;
wire x_6156;
wire x_6157;
wire x_6158;
wire x_6159;
wire x_6160;
wire x_6161;
wire x_6162;
wire x_6163;
wire x_6164;
wire x_6165;
wire x_6166;
wire x_6167;
wire x_6168;
wire x_6169;
wire x_6170;
wire x_6171;
wire x_6172;
wire x_6173;
wire x_6174;
wire x_6175;
wire x_6176;
wire x_6177;
wire x_6178;
wire x_6179;
wire x_6180;
wire x_6181;
wire x_6182;
wire x_6183;
wire x_6184;
wire x_6185;
wire x_6186;
wire x_6187;
wire x_6188;
wire x_6189;
wire x_6190;
wire x_6191;
wire x_6192;
wire x_6193;
wire x_6194;
wire x_6195;
wire x_6196;
wire x_6197;
wire x_6198;
wire x_6199;
wire x_6200;
wire x_6201;
wire x_6202;
wire x_6203;
wire x_6204;
wire x_6205;
wire x_6206;
wire x_6207;
wire x_6208;
wire x_6209;
wire x_6210;
wire x_6211;
wire x_6212;
wire x_6213;
wire x_6214;
wire x_6215;
wire x_6216;
wire x_6217;
wire x_6218;
wire x_6219;
wire x_6220;
wire x_6221;
wire x_6222;
wire x_6223;
wire x_6224;
wire x_6225;
wire x_6226;
wire x_6227;
wire x_6228;
wire x_6229;
wire x_6230;
wire x_6231;
wire x_6232;
wire x_6233;
wire x_6234;
wire x_6235;
wire x_6236;
wire x_6237;
wire x_6238;
wire x_6239;
wire x_6240;
wire x_6241;
wire x_6242;
wire x_6243;
wire x_6244;
wire x_6245;
wire x_6246;
wire x_6247;
wire x_6248;
wire x_6249;
wire x_6250;
wire x_6251;
wire x_6252;
wire x_6253;
wire x_6254;
wire x_6255;
wire x_6256;
wire x_6257;
wire x_6258;
wire x_6259;
wire x_6260;
wire x_6261;
wire x_6262;
wire x_6263;
wire x_6264;
wire x_6265;
wire x_6266;
wire x_6267;
wire x_6268;
wire x_6269;
wire x_6270;
wire x_6271;
wire x_6272;
wire x_6273;
wire x_6274;
wire x_6275;
wire x_6276;
wire x_6277;
wire x_6278;
wire x_6279;
wire x_6280;
wire x_6281;
wire x_6282;
wire x_6283;
wire x_6284;
wire x_6285;
wire x_6286;
wire x_6287;
wire x_6288;
wire x_6289;
wire x_6290;
wire x_6291;
wire x_6292;
wire x_6293;
wire x_6294;
wire x_6295;
wire x_6296;
wire x_6297;
wire x_6298;
wire x_6299;
wire x_6300;
wire x_6301;
wire x_6302;
wire x_6303;
wire x_6304;
wire x_6305;
wire x_6306;
wire x_6307;
wire x_6308;
wire x_6309;
wire x_6310;
wire x_6311;
wire x_6312;
wire x_6313;
wire x_6314;
wire x_6315;
wire x_6316;
wire x_6317;
wire x_6318;
wire x_6319;
wire x_6320;
wire x_6321;
wire x_6322;
wire x_6323;
wire x_6324;
wire x_6325;
wire x_6326;
wire x_6327;
wire x_6328;
wire x_6329;
wire x_6330;
wire x_6331;
wire x_6332;
wire x_6333;
wire x_6334;
wire x_6335;
wire x_6336;
wire x_6337;
wire x_6338;
wire x_6339;
wire x_6340;
wire x_6341;
wire x_6342;
wire x_6343;
wire x_6344;
wire x_6345;
wire x_6346;
wire x_6347;
wire x_6348;
wire x_6349;
wire x_6350;
wire x_6351;
wire x_6352;
wire x_6353;
wire x_6354;
wire x_6355;
wire x_6356;
wire x_6357;
wire x_6358;
wire x_6359;
wire x_6360;
wire x_6361;
wire x_6362;
wire x_6363;
wire x_6364;
wire x_6365;
wire x_6366;
wire x_6367;
wire x_6368;
wire x_6369;
wire x_6370;
wire x_6371;
wire x_6372;
wire x_6373;
wire x_6374;
wire x_6375;
wire x_6376;
wire x_6377;
wire x_6378;
wire x_6379;
wire x_6380;
wire x_6381;
wire x_6382;
wire x_6383;
wire x_6384;
wire x_6385;
wire x_6386;
wire x_6387;
wire x_6388;
wire x_6389;
wire x_6390;
wire x_6391;
wire x_6392;
wire x_6393;
wire x_6394;
wire x_6395;
wire x_6396;
wire x_6397;
wire x_6398;
wire x_6399;
wire x_6400;
wire x_6401;
wire x_6402;
wire x_6403;
wire x_6404;
wire x_6405;
wire x_6406;
wire x_6407;
wire x_6408;
wire x_6409;
wire x_6410;
wire x_6411;
wire x_6412;
wire x_6413;
wire x_6414;
wire x_6415;
wire x_6416;
wire x_6417;
wire x_6418;
wire x_6419;
wire x_6420;
wire x_6421;
wire x_6422;
wire x_6423;
wire x_6424;
wire x_6425;
wire x_6426;
wire x_6427;
wire x_6428;
wire x_6429;
wire x_6430;
wire x_6431;
wire x_6432;
wire x_6433;
wire x_6434;
wire x_6435;
wire x_6436;
wire x_6437;
wire x_6438;
wire x_6439;
wire x_6440;
wire x_6441;
wire x_6442;
wire x_6443;
wire x_6444;
wire x_6445;
wire x_6446;
wire x_6447;
wire x_6448;
wire x_6449;
wire x_6450;
wire x_6451;
wire x_6452;
wire x_6453;
wire x_6454;
wire x_6455;
wire x_6456;
wire x_6457;
wire x_6458;
wire x_6459;
wire x_6460;
wire x_6461;
wire x_6462;
wire x_6463;
wire x_6464;
wire x_6465;
wire x_6466;
wire x_6467;
wire x_6468;
wire x_6469;
wire x_6470;
wire x_6471;
wire x_6472;
wire x_6473;
wire x_6474;
wire x_6475;
wire x_6476;
wire x_6477;
wire x_6478;
wire x_6479;
wire x_6480;
wire x_6481;
wire x_6482;
wire x_6483;
wire x_6484;
wire x_6485;
wire x_6486;
wire x_6487;
wire x_6488;
wire x_6489;
wire x_6490;
wire x_6491;
wire x_6492;
wire x_6493;
wire x_6494;
wire x_6495;
wire x_6496;
wire x_6497;
wire x_6498;
wire x_6499;
wire x_6500;
wire x_6501;
wire x_6502;
wire x_6503;
wire x_6504;
wire x_6505;
wire x_6506;
wire x_6507;
wire x_6508;
wire x_6509;
wire x_6510;
wire x_6511;
wire x_6512;
wire x_6513;
wire x_6514;
wire x_6515;
wire x_6516;
wire x_6517;
wire x_6518;
wire x_6519;
wire x_6520;
wire x_6521;
wire x_6522;
wire x_6523;
wire x_6524;
wire x_6525;
wire x_6526;
wire x_6527;
wire x_6528;
wire x_6529;
wire x_6530;
wire x_6531;
wire x_6532;
wire x_6533;
wire x_6534;
wire x_6535;
wire x_6536;
wire x_6537;
wire x_6538;
wire x_6539;
wire x_6540;
wire x_6541;
wire x_6542;
wire x_6543;
wire x_6544;
wire x_6545;
wire x_6546;
wire x_6547;
wire x_6548;
wire x_6549;
wire x_6550;
wire x_6551;
wire x_6552;
wire x_6553;
wire x_6554;
wire x_6555;
wire x_6556;
wire x_6557;
wire x_6558;
wire x_6559;
wire x_6560;
wire x_6561;
wire x_6562;
wire x_6563;
wire x_6564;
wire x_6565;
wire x_6566;
wire x_6567;
wire x_6568;
wire x_6569;
wire x_6570;
wire x_6571;
wire x_6572;
wire x_6573;
wire x_6574;
wire x_6575;
wire x_6576;
wire x_6577;
wire x_6578;
wire x_6579;
wire x_6580;
wire x_6581;
wire x_6582;
wire x_6583;
wire x_6584;
wire x_6585;
wire x_6586;
wire x_6587;
wire x_6588;
wire x_6589;
wire x_6590;
wire x_6591;
wire x_6592;
wire x_6593;
wire x_6594;
wire x_6595;
wire x_6596;
wire x_6597;
wire x_6598;
wire x_6599;
wire x_6600;
wire x_6601;
wire x_6602;
wire x_6603;
wire x_6604;
wire x_6605;
wire x_6606;
wire x_6607;
wire x_6608;
wire x_6609;
wire x_6610;
wire x_6611;
wire x_6612;
wire x_6613;
wire x_6614;
wire x_6615;
wire x_6616;
wire x_6617;
wire x_6618;
wire x_6619;
wire x_6620;
wire x_6621;
wire x_6622;
wire x_6623;
wire x_6624;
wire x_6625;
wire x_6626;
wire x_6627;
wire x_6628;
wire x_6629;
wire x_6630;
wire x_6631;
wire x_6632;
wire x_6633;
wire x_6634;
wire x_6635;
wire x_6636;
wire x_6637;
wire x_6638;
wire x_6639;
wire x_6640;
wire x_6641;
wire x_6642;
wire x_6643;
wire x_6644;
wire x_6645;
wire x_6646;
wire x_6647;
wire x_6648;
wire x_6649;
wire x_6650;
wire x_6651;
wire x_6652;
wire x_6653;
wire x_6654;
wire x_6655;
wire x_6656;
wire x_6657;
wire x_6658;
wire x_6659;
wire x_6660;
wire x_6661;
wire x_6662;
wire x_6663;
wire x_6664;
wire x_6665;
wire x_6666;
wire x_6667;
wire x_6668;
wire x_6669;
wire x_6670;
wire x_6671;
wire x_6672;
wire x_6673;
wire x_6674;
wire x_6675;
wire x_6676;
wire x_6677;
wire x_6678;
wire x_6679;
wire x_6680;
wire x_6681;
wire x_6682;
wire x_6683;
wire x_6684;
wire x_6685;
wire x_6686;
wire x_6687;
wire x_6688;
wire x_6689;
wire x_6690;
wire x_6691;
wire x_6692;
wire x_6693;
wire x_6694;
wire x_6695;
wire x_6696;
wire x_6697;
wire x_6698;
wire x_6699;
wire x_6700;
wire x_6701;
wire x_6702;
wire x_6703;
wire x_6704;
wire x_6705;
wire x_6706;
wire x_6707;
wire x_6708;
wire x_6709;
wire x_6710;
wire x_6711;
wire x_6712;
wire x_6713;
wire x_6714;
wire x_6715;
wire x_6716;
wire x_6717;
wire x_6718;
wire x_6719;
wire x_6720;
wire x_6721;
wire x_6722;
wire x_6723;
wire x_6724;
wire x_6725;
wire x_6726;
wire x_6727;
wire x_6728;
wire x_6729;
wire x_6730;
wire x_6731;
wire x_6732;
wire x_6733;
wire x_6734;
wire x_6735;
wire x_6736;
wire x_6737;
wire x_6738;
wire x_6739;
wire x_6740;
wire x_6741;
wire x_6742;
wire x_6743;
wire x_6744;
wire x_6745;
wire x_6746;
wire x_6747;
wire x_6748;
wire x_6749;
wire x_6750;
wire x_6751;
wire x_6752;
wire x_6753;
wire x_6754;
wire x_6755;
wire x_6756;
wire x_6757;
wire x_6758;
wire x_6759;
wire x_6760;
wire x_6761;
wire x_6762;
wire x_6763;
wire x_6764;
wire x_6765;
wire x_6766;
wire x_6767;
wire x_6768;
wire x_6769;
wire x_6770;
wire x_6771;
wire x_6772;
wire x_6773;
wire x_6774;
wire x_6775;
wire x_6776;
wire x_6777;
wire x_6778;
wire x_6779;
wire x_6780;
wire x_6781;
wire x_6782;
wire x_6783;
wire x_6784;
wire x_6785;
wire x_6786;
wire x_6787;
wire x_6788;
wire x_6789;
wire x_6790;
wire x_6791;
wire x_6792;
wire x_6793;
wire x_6794;
wire x_6795;
wire x_6796;
wire x_6797;
wire x_6798;
wire x_6799;
wire x_6800;
wire x_6801;
wire x_6802;
wire x_6803;
wire x_6804;
wire x_6805;
wire x_6806;
wire x_6807;
wire x_6808;
wire x_6809;
wire x_6810;
wire x_6811;
wire x_6812;
wire x_6813;
wire x_6814;
wire x_6815;
wire x_6816;
wire x_6817;
wire x_6818;
wire x_6819;
wire x_6820;
wire x_6821;
wire x_6822;
wire x_6823;
wire x_6824;
wire x_6825;
wire x_6826;
wire x_6827;
wire x_6828;
wire x_6829;
wire x_6830;
wire x_6831;
wire x_6832;
wire x_6833;
wire x_6834;
wire x_6835;
wire x_6836;
wire x_6837;
wire x_6838;
wire x_6839;
wire x_6840;
wire x_6841;
wire x_6842;
wire x_6843;
wire x_6844;
wire x_6845;
wire x_6846;
wire x_6847;
wire x_6848;
wire x_6849;
wire x_6850;
wire x_6851;
wire x_6852;
wire x_6853;
wire x_6854;
wire x_6855;
wire x_6856;
wire x_6857;
wire x_6858;
wire x_6859;
wire x_6860;
wire x_6861;
wire x_6862;
wire x_6863;
wire x_6864;
wire x_6865;
wire x_6866;
wire x_6867;
wire x_6868;
wire x_6869;
wire x_6870;
wire x_6871;
wire x_6872;
wire x_6873;
wire x_6874;
wire x_6875;
wire x_6876;
wire x_6877;
wire x_6878;
wire x_6879;
wire x_6880;
wire x_6881;
wire x_6882;
wire x_6883;
wire x_6884;
wire x_6885;
wire x_6886;
wire x_6887;
wire x_6888;
wire x_6889;
wire x_6890;
wire x_6891;
wire x_6892;
wire x_6893;
wire x_6894;
wire x_6895;
wire x_6896;
wire x_6897;
wire x_6898;
wire x_6899;
wire x_6900;
wire x_6901;
wire x_6902;
wire x_6903;
wire x_6904;
wire x_6905;
wire x_6906;
wire x_6907;
wire x_6908;
wire x_6909;
wire x_6910;
wire x_6911;
wire x_6912;
wire x_6913;
wire x_6914;
wire x_6915;
wire x_6916;
wire x_6917;
wire x_6918;
wire x_6919;
wire x_6920;
wire x_6921;
wire x_6922;
wire x_6923;
wire x_6924;
wire x_6925;
wire x_6926;
wire x_6927;
wire x_6928;
wire x_6929;
wire x_6930;
wire x_6931;
wire x_6932;
wire x_6933;
wire x_6934;
wire x_6935;
wire x_6936;
wire x_6937;
wire x_6938;
wire x_6939;
wire x_6940;
wire x_6941;
wire x_6942;
wire x_6943;
wire x_6944;
wire x_6945;
wire x_6946;
wire x_6947;
wire x_6948;
wire x_6949;
wire x_6950;
wire x_6951;
wire x_6952;
wire x_6953;
wire x_6954;
wire x_6955;
wire x_6956;
wire x_6957;
wire x_6958;
wire x_6959;
wire x_6960;
wire x_6961;
wire x_6962;
wire x_6963;
wire x_6964;
wire x_6965;
wire x_6966;
wire x_6967;
wire x_6968;
wire x_6969;
wire x_6970;
wire x_6971;
wire x_6972;
wire x_6973;
wire x_6974;
wire x_6975;
wire x_6976;
wire x_6977;
wire x_6978;
wire x_6979;
wire x_6980;
wire x_6981;
wire x_6982;
wire x_6983;
wire x_6984;
wire x_6985;
wire x_6986;
wire x_6987;
wire x_6988;
wire x_6989;
wire x_6990;
wire x_6991;
wire x_6992;
wire x_6993;
wire x_6994;
wire x_6995;
wire x_6996;
wire x_6997;
wire x_6998;
wire x_6999;
wire x_7000;
wire x_7001;
wire x_7002;
wire x_7003;
wire x_7004;
wire x_7005;
wire x_7006;
wire x_7007;
wire x_7008;
wire x_7009;
wire x_7010;
wire x_7011;
wire x_7012;
wire x_7013;
wire x_7014;
wire x_7015;
wire x_7016;
wire x_7017;
wire x_7018;
wire x_7019;
wire x_7020;
wire x_7021;
wire x_7022;
wire x_7023;
wire x_7024;
wire x_7025;
wire x_7026;
wire x_7027;
wire x_7028;
wire x_7029;
wire x_7030;
wire x_7031;
wire x_7032;
wire x_7033;
wire x_7034;
wire x_7035;
wire x_7036;
wire x_7037;
wire x_7038;
wire x_7039;
wire x_7040;
wire x_7041;
wire x_7042;
wire x_7043;
wire x_7044;
wire x_7045;
wire x_7046;
wire x_7047;
wire x_7048;
wire x_7049;
wire x_7050;
wire x_7051;
wire x_7052;
wire x_7053;
wire x_7054;
wire x_7055;
wire x_7056;
wire x_7057;
wire x_7058;
wire x_7059;
wire x_7060;
wire x_7061;
wire x_7062;
wire x_7063;
wire x_7064;
wire x_7065;
wire x_7066;
wire x_7067;
wire x_7068;
wire x_7069;
wire x_7070;
wire x_7071;
wire x_7072;
wire x_7073;
wire x_7074;
wire x_7075;
wire x_7076;
wire x_7077;
wire x_7078;
wire x_7079;
wire x_7080;
wire x_7081;
wire x_7082;
wire x_7083;
wire x_7084;
wire x_7085;
wire x_7086;
wire x_7087;
wire x_7088;
wire x_7089;
wire x_7090;
wire x_7091;
wire x_7092;
wire x_7093;
wire x_7094;
wire x_7095;
wire x_7096;
wire x_7097;
wire x_7098;
wire x_7099;
wire x_7100;
wire x_7101;
wire x_7102;
wire x_7103;
wire x_7104;
wire x_7105;
wire x_7106;
wire x_7107;
wire x_7108;
wire x_7109;
wire x_7110;
wire x_7111;
wire x_7112;
wire x_7113;
wire x_7114;
wire x_7115;
wire x_7116;
wire x_7117;
wire x_7118;
wire x_7119;
wire x_7120;
wire x_7121;
wire x_7122;
wire x_7123;
wire x_7124;
wire x_7125;
wire x_7126;
wire x_7127;
wire x_7128;
wire x_7129;
wire x_7130;
wire x_7131;
wire x_7132;
wire x_7133;
wire x_7134;
wire x_7135;
wire x_7136;
wire x_7137;
wire x_7138;
wire x_7139;
wire x_7140;
wire x_7141;
wire x_7142;
wire x_7143;
wire x_7144;
wire x_7145;
wire x_7146;
wire x_7147;
wire x_7148;
wire x_7149;
wire x_7150;
wire x_7151;
wire x_7152;
wire x_7153;
wire x_7154;
wire x_7155;
wire x_7156;
wire x_7157;
wire x_7158;
wire x_7159;
wire x_7160;
wire x_7161;
wire x_7162;
wire x_7163;
wire x_7164;
wire x_7165;
wire x_7166;
wire x_7167;
wire x_7168;
wire x_7169;
wire x_7170;
wire x_7171;
wire x_7172;
wire x_7173;
wire x_7174;
wire x_7175;
wire x_7176;
wire x_7177;
wire x_7178;
wire x_7179;
wire x_7180;
wire x_7181;
wire x_7182;
wire x_7183;
wire x_7184;
wire x_7185;
wire x_7186;
wire x_7187;
wire x_7188;
wire x_7189;
wire x_7190;
wire x_7191;
wire x_7192;
wire x_7193;
wire x_7194;
wire x_7195;
wire x_7196;
wire x_7197;
wire x_7198;
wire x_7199;
wire x_7200;
wire x_7201;
wire x_7202;
wire x_7203;
wire x_7204;
wire x_7205;
wire x_7206;
wire x_7207;
wire x_7208;
wire x_7209;
wire x_7210;
wire x_7211;
wire x_7212;
wire x_7213;
wire x_7214;
wire x_7215;
wire x_7216;
wire x_7217;
wire x_7218;
wire x_7219;
wire x_7220;
wire x_7221;
wire x_7222;
wire x_7223;
wire x_7224;
wire x_7225;
wire x_7226;
wire x_7227;
wire x_7228;
wire x_7229;
wire x_7230;
wire x_7231;
wire x_7232;
wire x_7233;
wire x_7234;
wire x_7235;
wire x_7236;
wire x_7237;
wire x_7238;
wire x_7239;
wire x_7240;
wire x_7241;
wire x_7242;
wire x_7243;
wire x_7244;
wire x_7245;
wire x_7246;
wire x_7247;
wire x_7248;
wire x_7249;
wire x_7250;
wire x_7251;
wire x_7252;
wire x_7253;
wire x_7254;
wire x_7255;
wire x_7256;
wire x_7257;
wire x_7258;
wire x_7259;
wire x_7260;
wire x_7261;
wire x_7262;
wire x_7263;
wire x_7264;
wire x_7265;
wire x_7266;
wire x_7267;
wire x_7268;
wire x_7269;
wire x_7270;
wire x_7271;
wire x_7272;
wire x_7273;
wire x_7274;
wire x_7275;
wire x_7276;
wire x_7277;
wire x_7278;
wire x_7279;
wire x_7280;
wire x_7281;
wire x_7282;
wire x_7283;
wire x_7284;
wire x_7285;
wire x_7286;
wire x_7287;
wire x_7288;
wire x_7289;
wire x_7290;
wire x_7291;
wire x_7292;
wire x_7293;
wire x_7294;
wire x_7295;
wire x_7296;
wire x_7297;
wire x_7298;
wire x_7299;
wire x_7300;
wire x_7301;
wire x_7302;
wire x_7303;
wire x_7304;
wire x_7305;
wire x_7306;
wire x_7307;
wire x_7308;
wire x_7309;
wire x_7310;
wire x_7311;
wire x_7312;
wire x_7313;
wire x_7314;
wire x_7315;
wire x_7316;
wire x_7317;
wire x_7318;
wire x_7319;
wire x_7320;
wire x_7321;
wire x_7322;
wire x_7323;
wire x_7324;
wire x_7325;
wire x_7326;
wire x_7327;
wire x_7328;
wire x_7329;
wire x_7330;
wire x_7331;
wire x_7332;
wire x_7333;
wire x_7334;
wire x_7335;
wire x_7336;
wire x_7337;
wire x_7338;
wire x_7339;
wire x_7340;
wire x_7341;
wire x_7342;
wire x_7343;
wire x_7344;
wire x_7345;
wire x_7346;
wire x_7347;
wire x_7348;
wire x_7349;
wire x_7350;
wire x_7351;
wire x_7352;
wire x_7353;
wire x_7354;
wire x_7355;
wire x_7356;
wire x_7357;
wire x_7358;
wire x_7359;
wire x_7360;
wire x_7361;
wire x_7362;
wire x_7363;
wire x_7364;
wire x_7365;
wire x_7366;
wire x_7367;
wire x_7368;
wire x_7369;
wire x_7370;
wire x_7371;
wire x_7372;
wire x_7373;
wire x_7374;
wire x_7375;
wire x_7376;
wire x_7377;
wire x_7378;
wire x_7379;
wire x_7380;
wire x_7381;
wire x_7382;
wire x_7383;
wire x_7384;
wire x_7385;
wire x_7386;
wire x_7387;
wire x_7388;
wire x_7389;
wire x_7390;
wire x_7391;
wire x_7392;
wire x_7393;
wire x_7394;
wire x_7395;
wire x_7396;
wire x_7397;
wire x_7398;
wire x_7399;
wire x_7400;
wire x_7401;
wire x_7402;
wire x_7403;
wire x_7404;
wire x_7405;
wire x_7406;
wire x_7407;
wire x_7408;
wire x_7409;
wire x_7410;
wire x_7411;
wire x_7412;
wire x_7413;
wire x_7414;
wire x_7415;
wire x_7416;
wire x_7417;
wire x_7418;
wire x_7419;
wire x_7420;
wire x_7421;
wire x_7422;
wire x_7423;
wire x_7424;
wire x_7425;
wire x_7426;
wire x_7427;
wire x_7428;
wire x_7429;
wire x_7430;
wire x_7431;
wire x_7432;
wire x_7433;
wire x_7434;
wire x_7435;
wire x_7436;
wire x_7437;
wire x_7438;
wire x_7439;
wire x_7440;
wire x_7441;
wire x_7442;
wire x_7443;
wire x_7444;
wire x_7445;
wire x_7446;
wire x_7447;
wire x_7448;
wire x_7449;
wire x_7450;
wire x_7451;
wire x_7452;
wire x_7453;
wire x_7454;
wire x_7455;
wire x_7456;
wire x_7457;
wire x_7458;
wire x_7459;
wire x_7460;
wire x_7461;
wire x_7462;
wire x_7463;
wire x_7464;
wire x_7465;
wire x_7466;
wire x_7467;
wire x_7468;
wire x_7469;
wire x_7470;
wire x_7471;
wire x_7472;
wire x_7473;
wire x_7474;
wire x_7475;
wire x_7476;
wire x_7477;
wire x_7478;
wire x_7479;
wire x_7480;
wire x_7481;
wire x_7482;
wire x_7483;
wire x_7484;
wire x_7485;
wire x_7486;
wire x_7487;
wire x_7488;
wire x_7489;
wire x_7490;
wire x_7491;
wire x_7492;
wire x_7493;
wire x_7494;
wire x_7495;
wire x_7496;
wire x_7497;
wire x_7498;
wire x_7499;
wire x_7500;
wire x_7501;
wire x_7502;
wire x_7503;
wire x_7504;
wire x_7505;
wire x_7506;
wire x_7507;
wire x_7508;
wire x_7509;
wire x_7510;
wire x_7511;
wire x_7512;
wire x_7513;
wire x_7514;
wire x_7515;
wire x_7516;
wire x_7517;
wire x_7518;
wire x_7519;
wire x_7520;
wire x_7521;
wire x_7522;
wire x_7523;
wire x_7524;
wire x_7525;
wire x_7526;
wire x_7527;
wire x_7528;
wire x_7529;
wire x_7530;
wire x_7531;
wire x_7532;
wire x_7533;
wire x_7534;
wire x_7535;
wire x_7536;
wire x_7537;
wire x_7538;
wire x_7539;
wire x_7540;
wire x_7541;
wire x_7542;
wire x_7543;
wire x_7544;
wire x_7545;
wire x_7546;
wire x_7547;
wire x_7548;
wire x_7549;
wire x_7550;
wire x_7551;
wire x_7552;
wire x_7553;
wire x_7554;
wire x_7555;
wire x_7556;
wire x_7557;
wire x_7558;
wire x_7559;
wire x_7560;
wire x_7561;
wire x_7562;
wire x_7563;
wire x_7564;
wire x_7565;
wire x_7566;
wire x_7567;
wire x_7568;
wire x_7569;
wire x_7570;
wire x_7571;
wire x_7572;
wire x_7573;
wire x_7574;
wire x_7575;
wire x_7576;
wire x_7577;
wire x_7578;
wire x_7579;
wire x_7580;
wire x_7581;
wire x_7582;
wire x_7583;
wire x_7584;
wire x_7585;
wire x_7586;
wire x_7587;
wire x_7588;
wire x_7589;
wire x_7590;
wire x_7591;
wire x_7592;
wire x_7593;
wire x_7594;
wire x_7595;
wire x_7596;
wire x_7597;
wire x_7598;
wire x_7599;
wire x_7600;
wire x_7601;
wire x_7602;
wire x_7603;
wire x_7604;
wire x_7605;
wire x_7606;
wire x_7607;
wire x_7608;
wire x_7609;
wire x_7610;
wire x_7611;
wire x_7612;
wire x_7613;
wire x_7614;
wire x_7615;
wire x_7616;
wire x_7617;
wire x_7618;
wire x_7619;
wire x_7620;
wire x_7621;
wire x_7622;
wire x_7623;
wire x_7624;
wire x_7625;
wire x_7626;
wire x_7627;
wire x_7628;
wire x_7629;
wire x_7630;
wire x_7631;
wire x_7632;
wire x_7633;
wire x_7634;
wire x_7635;
wire x_7636;
wire x_7637;
wire x_7638;
wire x_7639;
wire x_7640;
wire x_7641;
wire x_7642;
wire x_7643;
wire x_7644;
wire x_7645;
wire x_7646;
wire x_7647;
wire x_7648;
wire x_7649;
wire x_7650;
wire x_7651;
wire x_7652;
wire x_7653;
wire x_7654;
wire x_7655;
wire x_7656;
wire x_7657;
wire x_7658;
wire x_7659;
wire x_7660;
wire x_7661;
wire x_7662;
wire x_7663;
wire x_7664;
wire x_7665;
wire x_7666;
wire x_7667;
wire x_7668;
wire x_7669;
wire x_7670;
wire x_7671;
wire x_7672;
wire x_7673;
wire x_7674;
wire x_7675;
wire x_7676;
wire x_7677;
wire x_7678;
wire x_7679;
wire x_7680;
wire x_7681;
wire x_7682;
wire x_7683;
wire x_7684;
wire x_7685;
wire x_7686;
wire x_7687;
wire x_7688;
wire x_7689;
wire x_7690;
wire x_7691;
wire x_7692;
wire x_7693;
wire x_7694;
wire x_7695;
wire x_7696;
wire x_7697;
wire x_7698;
wire x_7699;
wire x_7700;
wire x_7701;
wire x_7702;
wire x_7703;
wire x_7704;
wire x_7705;
wire x_7706;
wire x_7707;
wire x_7708;
wire x_7709;
wire x_7710;
wire x_7711;
wire x_7712;
wire x_7713;
wire x_7714;
wire x_7715;
wire x_7716;
wire x_7717;
wire x_7718;
wire x_7719;
wire x_7720;
wire x_7721;
wire x_7722;
wire x_7723;
wire x_7724;
wire x_7725;
wire x_7726;
wire x_7727;
wire x_7728;
wire x_7729;
wire x_7730;
wire x_7731;
wire x_7732;
wire x_7733;
wire x_7734;
wire x_7735;
wire x_7736;
wire x_7737;
wire x_7738;
wire x_7739;
wire x_7740;
wire x_7741;
wire x_7742;
wire x_7743;
wire x_7744;
wire x_7745;
wire x_7746;
wire x_7747;
wire x_7748;
wire x_7749;
wire x_7750;
wire x_7751;
wire x_7752;
wire x_7753;
wire x_7754;
wire x_7755;
wire x_7756;
wire x_7757;
wire x_7758;
wire x_7759;
wire x_7760;
wire x_7761;
wire x_7762;
wire x_7763;
wire x_7764;
wire x_7765;
wire x_7766;
wire x_7767;
wire x_7768;
wire x_7769;
wire x_7770;
wire x_7771;
wire x_7772;
wire x_7773;
wire x_7774;
wire x_7775;
wire x_7776;
wire x_7777;
wire x_7778;
wire x_7779;
wire x_7780;
wire x_7781;
wire x_7782;
wire x_7783;
wire x_7784;
wire x_7785;
wire x_7786;
wire x_7787;
wire x_7788;
wire x_7789;
wire x_7790;
wire x_7791;
wire x_7792;
wire x_7793;
wire x_7794;
wire x_7795;
wire x_7796;
wire x_7797;
wire x_7798;
wire x_7799;
wire x_7800;
wire x_7801;
wire x_7802;
wire x_7803;
wire x_7804;
wire x_7805;
wire x_7806;
wire x_7807;
wire x_7808;
wire x_7809;
wire x_7810;
wire x_7811;
wire x_7812;
wire x_7813;
wire x_7814;
wire x_7815;
wire x_7816;
wire x_7817;
wire x_7818;
wire x_7819;
wire x_7820;
wire x_7821;
wire x_7822;
wire x_7823;
wire x_7824;
wire x_7825;
wire x_7826;
wire x_7827;
wire x_7828;
wire x_7829;
wire x_7830;
wire x_7831;
wire x_7832;
wire x_7833;
wire x_7834;
wire x_7835;
wire x_7836;
wire x_7837;
wire x_7838;
wire x_7839;
wire x_7840;
wire x_7841;
wire x_7842;
wire x_7843;
wire x_7844;
wire x_7845;
wire x_7846;
wire x_7847;
wire x_7848;
wire x_7849;
wire x_7850;
wire x_7851;
wire x_7852;
wire x_7853;
wire x_7854;
wire x_7855;
wire x_7856;
wire x_7857;
wire x_7858;
wire x_7859;
wire x_7860;
wire x_7861;
wire x_7862;
wire x_7863;
wire x_7864;
wire x_7865;
wire x_7866;
wire x_7867;
wire x_7868;
wire x_7869;
wire x_7870;
wire x_7871;
wire x_7872;
wire x_7873;
wire x_7874;
wire x_7875;
wire x_7876;
wire x_7877;
wire x_7878;
wire x_7879;
wire x_7880;
wire x_7881;
wire x_7882;
wire x_7883;
wire x_7884;
wire x_7885;
wire x_7886;
wire x_7887;
wire x_7888;
wire x_7889;
wire x_7890;
wire x_7891;
wire x_7892;
wire x_7893;
wire x_7894;
wire x_7895;
wire x_7896;
wire x_7897;
wire x_7898;
wire x_7899;
wire x_7900;
wire x_7901;
wire x_7902;
wire x_7903;
wire x_7904;
wire x_7905;
wire x_7906;
wire x_7907;
wire x_7908;
wire x_7909;
wire x_7910;
wire x_7911;
wire x_7912;
wire x_7913;
wire x_7914;
wire x_7915;
wire x_7916;
wire x_7917;
wire x_7918;
wire x_7919;
wire x_7920;
wire x_7921;
wire x_7922;
wire x_7923;
wire x_7924;
wire x_7925;
wire x_7926;
wire x_7927;
wire x_7928;
wire x_7929;
wire x_7930;
wire x_7931;
wire x_7932;
wire x_7933;
wire x_7934;
wire x_7935;
wire x_7936;
wire x_7937;
wire x_7938;
wire x_7939;
wire x_7940;
wire x_7941;
wire x_7942;
wire x_7943;
wire x_7944;
wire x_7945;
wire x_7946;
wire x_7947;
wire x_7948;
wire x_7949;
wire x_7950;
wire x_7951;
wire x_7952;
wire x_7953;
wire x_7954;
wire x_7955;
wire x_7956;
wire x_7957;
wire x_7958;
wire x_7959;
wire x_7960;
wire x_7961;
wire x_7962;
wire x_7963;
wire x_7964;
wire x_7965;
wire x_7966;
wire x_7967;
wire x_7968;
wire x_7969;
wire x_7970;
wire x_7971;
wire x_7972;
wire x_7973;
wire x_7974;
wire x_7975;
wire x_7976;
wire x_7977;
wire x_7978;
wire x_7979;
wire x_7980;
wire x_7981;
wire x_7982;
wire x_7983;
wire x_7984;
wire x_7985;
wire x_7986;
wire x_7987;
wire x_7988;
wire x_7989;
wire x_7990;
wire x_7991;
wire x_7992;
wire x_7993;
wire x_7994;
wire x_7995;
wire x_7996;
wire x_7997;
wire x_7998;
wire x_7999;
wire x_8000;
wire x_8001;
wire x_8002;
wire x_8003;
wire x_8004;
wire x_8005;
wire x_8006;
wire x_8007;
wire x_8008;
wire x_8009;
wire x_8010;
wire x_8011;
wire x_8012;
wire x_8013;
wire x_8014;
wire x_8015;
wire x_8016;
wire x_8017;
wire x_8018;
wire x_8019;
wire x_8020;
wire x_8021;
wire x_8022;
wire x_8023;
wire x_8024;
wire x_8025;
wire x_8026;
wire x_8027;
wire x_8028;
wire x_8029;
wire x_8030;
wire x_8031;
wire x_8032;
wire x_8033;
wire x_8034;
wire x_8035;
wire x_8036;
wire x_8037;
wire x_8038;
wire x_8039;
wire x_8040;
wire x_8041;
wire x_8042;
wire x_8043;
wire x_8044;
wire x_8045;
wire x_8046;
wire x_8047;
wire x_8048;
wire x_8049;
wire x_8050;
wire x_8051;
wire x_8052;
wire x_8053;
wire x_8054;
wire x_8055;
wire x_8056;
wire x_8057;
wire x_8058;
wire x_8059;
wire x_8060;
wire x_8061;
wire x_8062;
wire x_8063;
wire x_8064;
wire x_8065;
wire x_8066;
wire x_8067;
wire x_8068;
wire x_8069;
wire x_8070;
wire x_8071;
wire x_8072;
wire x_8073;
wire x_8074;
wire x_8075;
wire x_8076;
wire x_8077;
wire x_8078;
wire x_8079;
wire x_8080;
wire x_8081;
wire x_8082;
wire x_8083;
wire x_8084;
wire x_8085;
wire x_8086;
wire x_8087;
wire x_8088;
wire x_8089;
wire x_8090;
wire x_8091;
wire x_8092;
wire x_8093;
wire x_8094;
wire x_8095;
wire x_8096;
wire x_8097;
wire x_8098;
wire x_8099;
wire x_8100;
wire x_8101;
wire x_8102;
wire x_8103;
wire x_8104;
wire x_8105;
wire x_8106;
wire x_8107;
wire x_8108;
wire x_8109;
wire x_8110;
wire x_8111;
wire x_8112;
wire x_8113;
wire x_8114;
wire x_8115;
wire x_8116;
wire x_8117;
wire x_8118;
wire x_8119;
wire x_8120;
wire x_8121;
wire x_8122;
wire x_8123;
wire x_8124;
wire x_8125;
wire x_8126;
wire x_8127;
wire x_8128;
wire x_8129;
wire x_8130;
wire x_8131;
wire x_8132;
wire x_8133;
wire x_8134;
wire x_8135;
wire x_8136;
wire x_8137;
wire x_8138;
wire x_8139;
wire x_8140;
wire x_8141;
wire x_8142;
wire x_8143;
wire x_8144;
wire x_8145;
wire x_8146;
wire x_8147;
wire x_8148;
wire x_8149;
wire x_8150;
wire x_8151;
wire x_8152;
wire x_8153;
wire x_8154;
wire x_8155;
wire x_8156;
wire x_8157;
wire x_8158;
wire x_8159;
wire x_8160;
wire x_8161;
wire x_8162;
wire x_8163;
wire x_8164;
wire x_8165;
wire x_8166;
wire x_8167;
wire x_8168;
wire x_8169;
wire x_8170;
wire x_8171;
wire x_8172;
wire x_8173;
wire x_8174;
wire x_8175;
wire x_8176;
wire x_8177;
wire x_8178;
wire x_8179;
wire x_8180;
wire x_8181;
wire x_8182;
wire x_8183;
wire x_8184;
wire x_8185;
wire x_8186;
wire x_8187;
wire x_8188;
wire x_8189;
wire x_8190;
wire x_8191;
wire x_8192;
wire x_8193;
wire x_8194;
wire x_8195;
wire x_8196;
wire x_8197;
wire x_8198;
wire x_8199;
wire x_8200;
wire x_8201;
wire x_8202;
wire x_8203;
wire x_8204;
wire x_8205;
wire x_8206;
wire x_8207;
wire x_8208;
wire x_8209;
wire x_8210;
wire x_8211;
wire x_8212;
wire x_8213;
wire x_8214;
wire x_8215;
wire x_8216;
wire x_8217;
wire x_8218;
wire x_8219;
wire x_8220;
wire x_8221;
wire x_8222;
wire x_8223;
wire x_8224;
wire x_8225;
wire x_8226;
wire x_8227;
wire x_8228;
wire x_8229;
wire x_8230;
wire x_8231;
wire x_8232;
wire x_8233;
wire x_8234;
wire x_8235;
wire x_8236;
wire x_8237;
wire x_8238;
wire x_8239;
wire x_8240;
wire x_8241;
wire x_8242;
wire x_8243;
wire x_8244;
wire x_8245;
wire x_8246;
wire x_8247;
wire x_8248;
wire x_8249;
wire x_8250;
wire x_8251;
wire x_8252;
wire x_8253;
wire x_8254;
wire x_8255;
wire x_8256;
wire x_8257;
wire x_8258;
wire x_8259;
wire x_8260;
wire x_8261;
wire x_8262;
wire x_8263;
wire x_8264;
wire x_8265;
wire x_8266;
wire x_8267;
wire x_8268;
wire x_8269;
wire x_8270;
wire x_8271;
wire x_8272;
wire x_8273;
wire x_8274;
wire x_8275;
wire x_8276;
wire x_8277;
wire x_8278;
wire x_8279;
wire x_8280;
wire x_8281;
wire x_8282;
wire x_8283;
wire x_8284;
wire x_8285;
wire x_8286;
wire x_8287;
wire x_8288;
wire x_8289;
wire x_8290;
wire x_8291;
wire x_8292;
wire x_8293;
wire x_8294;
wire x_8295;
wire x_8296;
wire x_8297;
wire x_8298;
wire x_8299;
wire x_8300;
wire x_8301;
wire x_8302;
wire x_8303;
wire x_8304;
wire x_8305;
wire x_8306;
wire x_8307;
wire x_8308;
wire x_8309;
wire x_8310;
wire x_8311;
wire x_8312;
wire x_8313;
wire x_8314;
wire x_8315;
wire x_8316;
wire x_8317;
wire x_8318;
wire x_8319;
wire x_8320;
wire x_8321;
wire x_8322;
wire x_8323;
wire x_8324;
wire x_8325;
wire x_8326;
wire x_8327;
wire x_8328;
wire x_8329;
wire x_8330;
wire x_8331;
wire x_8332;
wire x_8333;
wire x_8334;
wire x_8335;
wire x_8336;
wire x_8337;
wire x_8338;
wire x_8339;
wire x_8340;
wire x_8341;
wire x_8342;
wire x_8343;
wire x_8344;
wire x_8345;
wire x_8346;
wire x_8347;
wire x_8348;
wire x_8349;
wire x_8350;
wire x_8351;
wire x_8352;
wire x_8353;
wire x_8354;
wire x_8355;
wire x_8356;
wire x_8357;
wire x_8358;
wire x_8359;
wire x_8360;
wire x_8361;
wire x_8362;
wire x_8363;
wire x_8364;
wire x_8365;
wire x_8366;
wire x_8367;
wire x_8368;
wire x_8369;
wire x_8370;
wire x_8371;
wire x_8372;
wire x_8373;
wire x_8374;
wire x_8375;
wire x_8376;
wire x_8377;
wire x_8378;
wire x_8379;
wire x_8380;
wire x_8381;
wire x_8382;
wire x_8383;
wire x_8384;
wire x_8385;
wire x_8386;
wire x_8387;
wire x_8388;
wire x_8389;
wire x_8390;
wire x_8391;
wire x_8392;
wire x_8393;
wire x_8394;
wire x_8395;
wire x_8396;
wire x_8397;
wire x_8398;
wire x_8399;
wire x_8400;
wire x_8401;
wire x_8402;
wire x_8403;
wire x_8404;
wire x_8405;
wire x_8406;
wire x_8407;
wire x_8408;
wire x_8409;
wire x_8410;
wire x_8411;
wire x_8412;
wire x_8413;
wire x_8414;
wire x_8415;
wire x_8416;
wire x_8417;
wire x_8418;
wire x_8419;
wire x_8420;
wire x_8421;
wire x_8422;
wire x_8423;
wire x_8424;
wire x_8425;
wire x_8426;
wire x_8427;
wire x_8428;
wire x_8429;
wire x_8430;
wire x_8431;
wire x_8432;
wire x_8433;
wire x_8434;
wire x_8435;
wire x_8436;
wire x_8437;
wire x_8438;
wire x_8439;
wire x_8440;
wire x_8441;
wire x_8442;
wire x_8443;
wire x_8444;
wire x_8445;
wire x_8446;
wire x_8447;
wire x_8448;
wire x_8449;
wire x_8450;
wire x_8451;
wire x_8452;
wire x_8453;
wire x_8454;
wire x_8455;
wire x_8456;
wire x_8457;
wire x_8458;
wire x_8459;
wire x_8460;
wire x_8461;
wire x_8462;
wire x_8463;
wire x_8464;
wire x_8465;
wire x_8466;
wire x_8467;
wire x_8468;
wire x_8469;
wire x_8470;
wire x_8471;
wire x_8472;
wire x_8473;
wire x_8474;
wire x_8475;
wire x_8476;
wire x_8477;
wire x_8478;
wire x_8479;
wire x_8480;
wire x_8481;
wire x_8482;
wire x_8483;
wire x_8484;
wire x_8485;
wire x_8486;
wire x_8487;
wire x_8488;
wire x_8489;
wire x_8490;
wire x_8491;
wire x_8492;
wire x_8493;
wire x_8494;
wire x_8495;
wire x_8496;
wire x_8497;
wire x_8498;
wire x_8499;
wire x_8500;
wire x_8501;
wire x_8502;
wire x_8503;
wire x_8504;
wire x_8505;
wire x_8506;
wire x_8507;
wire x_8508;
wire x_8509;
wire x_8510;
wire x_8511;
wire x_8512;
wire x_8513;
wire x_8514;
wire x_8515;
wire x_8516;
wire x_8517;
wire x_8518;
wire x_8519;
wire x_8520;
wire x_8521;
wire x_8522;
wire x_8523;
wire x_8524;
wire x_8525;
wire x_8526;
wire x_8527;
wire x_8528;
wire x_8529;
wire x_8530;
wire x_8531;
wire x_8532;
wire x_8533;
wire x_8534;
wire x_8535;
wire x_8536;
wire x_8537;
wire x_8538;
wire x_8539;
wire x_8540;
wire x_8541;
wire x_8542;
wire x_8543;
wire x_8544;
wire x_8545;
wire x_8546;
wire x_8547;
wire x_8548;
wire x_8549;
wire x_8550;
wire x_8551;
wire x_8552;
wire x_8553;
wire x_8554;
wire x_8555;
wire x_8556;
wire x_8557;
wire x_8558;
wire x_8559;
wire x_8560;
wire x_8561;
wire x_8562;
wire x_8563;
wire x_8564;
wire x_8565;
wire x_8566;
wire x_8567;
wire x_8568;
wire x_8569;
wire x_8570;
wire x_8571;
wire x_8572;
wire x_8573;
wire x_8574;
wire x_8575;
wire x_8576;
wire x_8577;
wire x_8578;
wire x_8579;
wire x_8580;
wire x_8581;
wire x_8582;
wire x_8583;
wire x_8584;
wire x_8585;
wire x_8586;
wire x_8587;
wire x_8588;
wire x_8589;
wire x_8590;
wire x_8591;
wire x_8592;
wire x_8593;
wire x_8594;
wire x_8595;
wire x_8596;
wire x_8597;
wire x_8598;
wire x_8599;
wire x_8600;
wire x_8601;
wire x_8602;
wire x_8603;
wire x_8604;
wire x_8605;
wire x_8606;
wire x_8607;
wire x_8608;
wire x_8609;
wire x_8610;
wire x_8611;
wire x_8612;
wire x_8613;
wire x_8614;
wire x_8615;
wire x_8616;
wire x_8617;
wire x_8618;
wire x_8619;
wire x_8620;
wire x_8621;
wire x_8622;
wire x_8623;
wire x_8624;
wire x_8625;
wire x_8626;
wire x_8627;
wire x_8628;
wire x_8629;
wire x_8630;
wire x_8631;
wire x_8632;
wire x_8633;
wire x_8634;
wire x_8635;
wire x_8636;
wire x_8637;
wire x_8638;
wire x_8639;
wire x_8640;
wire x_8641;
wire x_8642;
wire x_8643;
wire x_8644;
wire x_8645;
wire x_8646;
wire x_8647;
wire x_8648;
wire x_8649;
wire x_8650;
wire x_8651;
wire x_8652;
wire x_8653;
wire x_8654;
wire x_8655;
wire x_8656;
wire x_8657;
wire x_8658;
wire x_8659;
wire x_8660;
wire x_8661;
wire x_8662;
wire x_8663;
wire x_8664;
wire x_8665;
wire x_8666;
wire x_8667;
wire x_8668;
wire x_8669;
wire x_8670;
wire x_8671;
wire x_8672;
wire x_8673;
wire x_8674;
wire x_8675;
wire x_8676;
wire x_8677;
wire x_8678;
wire x_8679;
wire x_8680;
wire x_8681;
wire x_8682;
wire x_8683;
wire x_8684;
wire x_8685;
wire x_8686;
wire x_8687;
wire x_8688;
wire x_8689;
wire x_8690;
wire x_8691;
wire x_8692;
wire x_8693;
wire x_8694;
wire x_8695;
wire x_8696;
wire x_8697;
wire x_8698;
wire x_8699;
wire x_8700;
wire x_8701;
wire x_8702;
wire x_8703;
wire x_8704;
wire x_8705;
wire x_8706;
wire x_8707;
wire x_8708;
wire x_8709;
wire x_8710;
wire x_8711;
wire x_8712;
wire x_8713;
wire x_8714;
wire x_8715;
wire x_8716;
wire x_8717;
wire x_8718;
wire x_8719;
wire x_8720;
wire x_8721;
wire x_8722;
wire x_8723;
wire x_8724;
wire x_8725;
wire x_8726;
wire x_8727;
wire x_8728;
wire x_8729;
wire x_8730;
wire x_8731;
wire x_8732;
wire x_8733;
wire x_8734;
wire x_8735;
wire x_8736;
wire x_8737;
wire x_8738;
wire x_8739;
wire x_8740;
wire x_8741;
wire x_8742;
wire x_8743;
wire x_8744;
wire x_8745;
wire x_8746;
wire x_8747;
wire x_8748;
wire x_8749;
wire x_8750;
wire x_8751;
wire x_8752;
wire x_8753;
wire x_8754;
wire x_8755;
wire x_8756;
wire x_8757;
wire x_8758;
wire x_8759;
wire x_8760;
wire x_8761;
wire x_8762;
wire x_8763;
wire x_8764;
wire x_8765;
wire x_8766;
wire x_8767;
wire x_8768;
wire x_8769;
wire x_8770;
wire x_8771;
wire x_8772;
wire x_8773;
wire x_8774;
wire x_8775;
wire x_8776;
wire x_8777;
wire x_8778;
wire x_8779;
wire x_8780;
wire x_8781;
wire x_8782;
wire x_8783;
wire x_8784;
wire x_8785;
wire x_8786;
wire x_8787;
wire x_8788;
wire x_8789;
wire x_8790;
wire x_8791;
wire x_8792;
wire x_8793;
wire x_8794;
wire x_8795;
wire x_8796;
wire x_8797;
wire x_8798;
wire x_8799;
wire x_8800;
wire x_8801;
wire x_8802;
wire x_8803;
wire x_8804;
wire x_8805;
wire x_8806;
wire x_8807;
wire x_8808;
wire x_8809;
wire x_8810;
wire x_8811;
wire x_8812;
wire x_8813;
wire x_8814;
wire x_8815;
wire x_8816;
wire x_8817;
wire x_8818;
wire x_8819;
wire x_8820;
wire x_8821;
wire x_8822;
wire x_8823;
wire x_8824;
wire x_8825;
wire x_8826;
wire x_8827;
wire x_8828;
wire x_8829;
wire x_8830;
wire x_8831;
wire x_8832;
wire x_8833;
wire x_8834;
wire x_8835;
wire x_8836;
wire x_8837;
wire x_8838;
wire x_8839;
wire x_8840;
wire x_8841;
wire x_8842;
wire x_8843;
wire x_8844;
wire x_8845;
wire x_8846;
wire x_8847;
wire x_8848;
wire x_8849;
wire x_8850;
wire x_8851;
wire x_8852;
wire x_8853;
wire x_8854;
wire x_8855;
wire x_8856;
wire x_8857;
wire x_8858;
wire x_8859;
wire x_8860;
wire x_8861;
wire x_8862;
wire x_8863;
wire x_8864;
wire x_8865;
wire x_8866;
wire x_8867;
wire x_8868;
wire x_8869;
wire x_8870;
wire x_8871;
wire x_8872;
wire x_8873;
wire x_8874;
wire x_8875;
wire x_8876;
wire x_8877;
wire x_8878;
wire x_8879;
wire x_8880;
wire x_8881;
wire x_8882;
wire x_8883;
wire x_8884;
wire x_8885;
wire x_8886;
wire x_8887;
wire x_8888;
wire x_8889;
wire x_8890;
wire x_8891;
wire x_8892;
wire x_8893;
wire x_8894;
wire x_8895;
wire x_8896;
wire x_8897;
wire x_8898;
wire x_8899;
wire x_8900;
wire x_8901;
wire x_8902;
wire x_8903;
wire x_8904;
wire x_8905;
wire x_8906;
wire x_8907;
wire x_8908;
wire x_8909;
wire x_8910;
wire x_8911;
wire x_8912;
wire x_8913;
wire x_8914;
wire x_8915;
wire x_8916;
wire x_8917;
wire x_8918;
wire x_8919;
wire x_8920;
wire x_8921;
wire x_8922;
wire x_8923;
wire x_8924;
wire x_8925;
wire x_8926;
wire x_8927;
wire x_8928;
wire x_8929;
wire x_8930;
wire x_8931;
wire x_8932;
wire x_8933;
wire x_8934;
wire x_8935;
wire x_8936;
wire x_8937;
wire x_8938;
wire x_8939;
wire x_8940;
wire x_8941;
wire x_8942;
wire x_8943;
wire x_8944;
wire x_8945;
wire x_8946;
wire x_8947;
wire x_8948;
wire x_8949;
wire x_8950;
wire x_8951;
wire x_8952;
wire x_8953;
wire x_8954;
wire x_8955;
wire x_8956;
wire x_8957;
wire x_8958;
wire x_8959;
wire x_8960;
wire x_8961;
wire x_8962;
wire x_8963;
wire x_8964;
wire x_8965;
wire x_8966;
wire x_8967;
wire x_8968;
wire x_8969;
wire x_8970;
wire x_8971;
wire x_8972;
wire x_8973;
wire x_8974;
wire x_8975;
wire x_8976;
wire x_8977;
wire x_8978;
wire x_8979;
wire x_8980;
wire x_8981;
wire x_8982;
wire x_8983;
wire x_8984;
wire x_8985;
wire x_8986;
wire x_8987;
wire x_8988;
wire x_8989;
wire x_8990;
wire x_8991;
wire x_8992;
wire x_8993;
wire x_8994;
wire x_8995;
wire x_8996;
wire x_8997;
wire x_8998;
wire x_8999;
wire x_9000;
wire x_9001;
wire x_9002;
wire x_9003;
wire x_9004;
wire x_9005;
wire x_9006;
wire x_9007;
wire x_9008;
wire x_9009;
wire x_9010;
wire x_9011;
wire x_9012;
wire x_9013;
wire x_9014;
wire x_9015;
wire x_9016;
wire x_9017;
wire x_9018;
wire x_9019;
wire x_9020;
wire x_9021;
wire x_9022;
wire x_9023;
wire x_9024;
wire x_9025;
wire x_9026;
wire x_9027;
wire x_9028;
wire x_9029;
wire x_9030;
wire x_9031;
wire x_9032;
wire x_9033;
wire x_9034;
wire x_9035;
wire x_9036;
wire x_9037;
wire x_9038;
wire x_9039;
wire x_9040;
wire x_9041;
wire x_9042;
wire x_9043;
wire x_9044;
wire x_9045;
wire x_9046;
wire x_9047;
wire x_9048;
wire x_9049;
wire x_9050;
wire x_9051;
wire x_9052;
wire x_9053;
wire x_9054;
wire x_9055;
wire x_9056;
wire x_9057;
wire x_9058;
wire x_9059;
wire x_9060;
wire x_9061;
wire x_9062;
wire x_9063;
wire x_9064;
wire x_9065;
wire x_9066;
wire x_9067;
wire x_9068;
wire x_9069;
wire x_9070;
wire x_9071;
wire x_9072;
wire x_9073;
wire x_9074;
wire x_9075;
wire x_9076;
wire x_9077;
wire x_9078;
wire x_9079;
wire x_9080;
wire x_9081;
wire x_9082;
wire x_9083;
wire x_9084;
wire x_9085;
wire x_9086;
wire x_9087;
wire x_9088;
wire x_9089;
wire x_9090;
wire x_9091;
wire x_9092;
wire x_9093;
wire x_9094;
wire x_9095;
wire x_9096;
wire x_9097;
wire x_9098;
wire x_9099;
wire x_9100;
wire x_9101;
wire x_9102;
wire x_9103;
wire x_9104;
wire x_9105;
wire x_9106;
wire x_9107;
wire x_9108;
wire x_9109;
wire x_9110;
wire x_9111;
wire x_9112;
wire x_9113;
wire x_9114;
wire x_9115;
wire x_9116;
wire x_9117;
wire x_9118;
wire x_9119;
wire x_9120;
wire x_9121;
wire x_9122;
wire x_9123;
wire x_9124;
wire x_9125;
wire x_9126;
wire x_9127;
wire x_9128;
wire x_9129;
wire x_9130;
wire x_9131;
wire x_9132;
wire x_9133;
wire x_9134;
wire x_9135;
wire x_9136;
wire x_9137;
wire x_9138;
wire x_9139;
wire x_9140;
wire x_9141;
wire x_9142;
wire x_9143;
wire x_9144;
wire x_9145;
wire x_9146;
wire x_9147;
wire x_9148;
wire x_9149;
wire x_9150;
wire x_9151;
wire x_9152;
wire x_9153;
wire x_9154;
wire x_9155;
wire x_9156;
wire x_9157;
wire x_9158;
wire x_9159;
wire x_9160;
wire x_9161;
wire x_9162;
wire x_9163;
wire x_9164;
wire x_9165;
wire x_9166;
wire x_9167;
wire x_9168;
wire x_9169;
wire x_9170;
wire x_9171;
wire x_9172;
wire x_9173;
wire x_9174;
wire x_9175;
wire x_9176;
wire x_9177;
wire x_9178;
wire x_9179;
wire x_9180;
wire x_9181;
wire x_9182;
wire x_9183;
wire x_9184;
wire x_9185;
wire x_9186;
wire x_9187;
wire x_9188;
wire x_9189;
wire x_9190;
wire x_9191;
wire x_9192;
wire x_9193;
wire x_9194;
wire x_9195;
wire x_9196;
wire x_9197;
wire x_9198;
wire x_9199;
wire x_9200;
wire x_9201;
wire x_9202;
wire x_9203;
wire x_9204;
wire x_9205;
wire x_9206;
wire x_9207;
wire x_9208;
wire x_9209;
wire x_9210;
wire x_9211;
wire x_9212;
wire x_9213;
wire x_9214;
wire x_9215;
wire x_9216;
wire x_9217;
wire x_9218;
wire x_9219;
wire x_9220;
wire x_9221;
wire x_9222;
wire x_9223;
wire x_9224;
wire x_9225;
wire x_9226;
wire x_9227;
wire x_9228;
wire x_9229;
wire x_9230;
wire x_9231;
wire x_9232;
wire x_9233;
wire x_9234;
wire x_9235;
wire x_9236;
wire x_9237;
wire x_9238;
wire x_9239;
wire x_9240;
wire x_9241;
wire x_9242;
wire x_9243;
wire x_9244;
wire x_9245;
wire x_9246;
wire x_9247;
wire x_9248;
wire x_9249;
wire x_9250;
wire x_9251;
wire x_9252;
wire x_9253;
wire x_9254;
wire x_9255;
wire x_9256;
wire x_9257;
wire x_9258;
wire x_9259;
wire x_9260;
wire x_9261;
wire x_9262;
wire x_9263;
wire x_9264;
wire x_9265;
wire x_9266;
wire x_9267;
wire x_9268;
wire x_9269;
wire x_9270;
wire x_9271;
wire x_9272;
wire x_9273;
wire x_9274;
wire x_9275;
wire x_9276;
wire x_9277;
wire x_9278;
wire x_9279;
wire x_9280;
wire x_9281;
wire x_9282;
wire x_9283;
wire x_9284;
wire x_9285;
wire x_9286;
wire x_9287;
wire x_9288;
wire x_9289;
wire x_9290;
wire x_9291;
wire x_9292;
wire x_9293;
wire x_9294;
wire x_9295;
wire x_9296;
wire x_9297;
wire x_9298;
wire x_9299;
wire x_9300;
wire x_9301;
wire x_9302;
wire x_9303;
wire x_9304;
wire x_9305;
wire x_9306;
wire x_9307;
wire x_9308;
wire x_9309;
wire x_9310;
wire x_9311;
wire x_9312;
wire x_9313;
wire x_9314;
wire x_9315;
wire x_9316;
wire x_9317;
wire x_9318;
wire x_9319;
wire x_9320;
wire x_9321;
wire x_9322;
wire x_9323;
wire x_9324;
wire x_9325;
wire x_9326;
wire x_9327;
wire x_9328;
wire x_9329;
wire x_9330;
wire x_9331;
wire x_9332;
wire x_9333;
wire x_9334;
wire x_9335;
wire x_9336;
wire x_9337;
wire x_9338;
wire x_9339;
wire x_9340;
wire x_9341;
wire x_9342;
wire x_9343;
wire x_9344;
wire x_9345;
wire x_9346;
wire x_9347;
wire x_9348;
wire x_9349;
wire x_9350;
wire x_9351;
wire x_9352;
wire x_9353;
wire x_9354;
wire x_9355;
wire x_9356;
wire x_9357;
wire x_9358;
wire x_9359;
wire x_9360;
wire x_9361;
wire x_9362;
wire x_9363;
wire x_9364;
wire x_9365;
wire x_9366;
wire x_9367;
wire x_9368;
wire x_9369;
wire x_9370;
wire x_9371;
wire x_9372;
wire x_9373;
wire x_9374;
wire x_9375;
wire x_9376;
wire x_9377;
wire x_9378;
wire x_9379;
wire x_9380;
wire x_9381;
wire x_9382;
wire x_9383;
wire x_9384;
wire x_9385;
wire x_9386;
wire x_9387;
wire x_9388;
wire x_9389;
wire x_9390;
wire x_9391;
wire x_9392;
wire x_9393;
wire x_9394;
wire x_9395;
wire x_9396;
wire x_9397;
wire x_9398;
wire x_9399;
wire x_9400;
wire x_9401;
wire x_9402;
wire x_9403;
wire x_9404;
wire x_9405;
wire x_9406;
wire x_9407;
wire x_9408;
wire x_9409;
wire x_9410;
wire x_9411;
wire x_9412;
wire x_9413;
wire x_9414;
wire x_9415;
wire x_9416;
wire x_9417;
wire x_9418;
wire x_9419;
wire x_9420;
wire x_9421;
wire x_9422;
wire x_9423;
wire x_9424;
wire x_9425;
wire x_9426;
wire x_9427;
wire x_9428;
wire x_9429;
wire x_9430;
wire x_9431;
wire x_9432;
wire x_9433;
wire x_9434;
wire x_9435;
wire x_9436;
wire x_9437;
wire x_9438;
wire x_9439;
wire x_9440;
wire x_9441;
wire x_9442;
wire x_9443;
wire x_9444;
wire x_9445;
wire x_9446;
wire x_9447;
wire x_9448;
wire x_9449;
wire x_9450;
wire x_9451;
wire x_9452;
wire x_9453;
wire x_9454;
wire x_9455;
wire x_9456;
wire x_9457;
wire x_9458;
wire x_9459;
wire x_9460;
wire x_9461;
wire x_9462;
wire x_9463;
wire x_9464;
wire x_9465;
wire x_9466;
wire x_9467;
wire x_9468;
wire x_9469;
wire x_9470;
wire x_9471;
wire x_9472;
wire x_9473;
wire x_9474;
wire x_9475;
wire x_9476;
wire x_9477;
wire x_9478;
wire x_9479;
wire x_9480;
wire x_9481;
wire x_9482;
wire x_9483;
wire x_9484;
wire x_9485;
wire x_9486;
wire x_9487;
wire x_9488;
wire x_9489;
wire x_9490;
wire x_9491;
wire x_9492;
wire x_9493;
wire x_9494;
wire x_9495;
wire x_9496;
wire x_9497;
wire x_9498;
wire x_9499;
wire x_9500;
wire x_9501;
wire x_9502;
wire x_9503;
wire x_9504;
wire x_9505;
wire x_9506;
wire x_9507;
wire x_9508;
wire x_9509;
wire x_9510;
wire x_9511;
wire x_9512;
wire x_9513;
wire x_9514;
wire x_9515;
wire x_9516;
wire x_9517;
wire x_9518;
wire x_9519;
wire x_9520;
wire x_9521;
wire x_9522;
wire x_9523;
wire x_9524;
wire x_9525;
wire x_9526;
wire x_9527;
wire x_9528;
wire x_9529;
wire x_9530;
wire x_9531;
wire x_9532;
wire x_9533;
wire x_9534;
wire x_9535;
wire x_9536;
wire x_9537;
wire x_9538;
wire x_9539;
wire x_9540;
wire x_9541;
wire x_9542;
wire x_9543;
wire x_9544;
wire x_9545;
wire x_9546;
wire x_9547;
wire x_9548;
wire x_9549;
wire x_9550;
wire x_9551;
wire x_9552;
wire x_9553;
wire x_9554;
wire x_9555;
wire x_9556;
wire x_9557;
wire x_9558;
wire x_9559;
wire x_9560;
wire x_9561;
wire x_9562;
wire x_9563;
wire x_9564;
wire x_9565;
wire x_9566;
wire x_9567;
wire x_9568;
wire x_9569;
wire x_9570;
wire x_9571;
wire x_9572;
wire x_9573;
wire x_9574;
wire x_9575;
wire x_9576;
wire x_9577;
wire x_9578;
wire x_9579;
wire x_9580;
wire x_9581;
wire x_9582;
wire x_9583;
wire x_9584;
wire x_9585;
wire x_9586;
wire x_9587;
wire x_9588;
wire x_9589;
wire x_9590;
wire x_9591;
wire x_9592;
wire x_9593;
wire x_9594;
wire x_9595;
wire x_9596;
wire x_9597;
wire x_9598;
wire x_9599;
wire x_9600;
wire x_9601;
wire x_9602;
wire x_9603;
wire x_9604;
wire x_9605;
wire x_9606;
wire x_9607;
wire x_9608;
wire x_9609;
wire x_9610;
wire x_9611;
wire x_9612;
wire x_9613;
wire x_9614;
wire x_9615;
wire x_9616;
wire x_9617;
wire x_9618;
wire x_9619;
wire x_9620;
wire x_9621;
wire x_9622;
wire x_9623;
wire x_9624;
wire x_9625;
wire x_9626;
wire x_9627;
wire x_9628;
wire x_9629;
wire x_9630;
wire x_9631;
wire x_9632;
wire x_9633;
wire x_9634;
wire x_9635;
wire x_9636;
wire x_9637;
wire x_9638;
wire x_9639;
wire x_9640;
wire x_9641;
wire x_9642;
wire x_9643;
wire x_9644;
wire x_9645;
wire x_9646;
wire x_9647;
wire x_9648;
wire x_9649;
wire x_9650;
wire x_9651;
wire x_9652;
wire x_9653;
wire x_9654;
wire x_9655;
wire x_9656;
wire x_9657;
wire x_9658;
wire x_9659;
wire x_9660;
wire x_9661;
wire x_9662;
wire x_9663;
wire x_9664;
wire x_9665;
wire x_9666;
wire x_9667;
wire x_9668;
wire x_9669;
wire x_9670;
wire x_9671;
wire x_9672;
wire x_9673;
wire x_9674;
wire x_9675;
wire x_9676;
wire x_9677;
wire x_9678;
wire x_9679;
wire x_9680;
wire x_9681;
wire x_9682;
wire x_9683;
wire x_9684;
wire x_9685;
wire x_9686;
wire x_9687;
wire x_9688;
wire x_9689;
wire x_9690;
wire x_9691;
wire x_9692;
wire x_9693;
wire x_9694;
wire x_9695;
wire x_9696;
wire x_9697;
wire x_9698;
wire x_9699;
wire x_9700;
wire x_9701;
wire x_9702;
wire x_9703;
wire x_9704;
wire x_9705;
wire x_9706;
wire x_9707;
wire x_9708;
wire x_9709;
wire x_9710;
wire x_9711;
wire x_9712;
wire x_9713;
wire x_9714;
wire x_9715;
wire x_9716;
wire x_9717;
wire x_9718;
wire x_9719;
wire x_9720;
wire x_9721;
wire x_9722;
wire x_9723;
wire x_9724;
wire x_9725;
wire x_9726;
wire x_9727;
wire x_9728;
wire x_9729;
wire x_9730;
wire x_9731;
wire x_9732;
wire x_9733;
wire x_9734;
wire x_9735;
wire x_9736;
wire x_9737;
wire x_9738;
wire x_9739;
wire x_9740;
wire x_9741;
wire x_9742;
wire x_9743;
wire x_9744;
wire x_9745;
wire x_9746;
wire x_9747;
wire x_9748;
wire x_9749;
wire x_9750;
wire x_9751;
wire x_9752;
wire x_9753;
wire x_9754;
wire x_9755;
wire x_9756;
wire x_9757;
wire x_9758;
wire x_9759;
wire x_9760;
wire x_9761;
wire x_9762;
wire x_9763;
wire x_9764;
wire x_9765;
wire x_9766;
wire x_9767;
wire x_9768;
wire x_9769;
wire x_9770;
wire x_9771;
wire x_9772;
wire x_9773;
wire x_9774;
wire x_9775;
wire x_9776;
wire x_9777;
wire x_9778;
wire x_9779;
wire x_9780;
wire x_9781;
wire x_9782;
wire x_9783;
wire x_9784;
wire x_9785;
wire x_9786;
wire x_9787;
wire x_9788;
wire x_9789;
wire x_9790;
wire x_9791;
wire x_9792;
wire x_9793;
wire x_9794;
wire x_9795;
wire x_9796;
wire x_9797;
wire x_9798;
wire x_9799;
wire x_9800;
wire x_9801;
wire x_9802;
wire x_9803;
wire x_9804;
wire x_9805;
wire x_9806;
wire x_9807;
wire x_9808;
wire x_9809;
wire x_9810;
wire x_9811;
wire x_9812;
wire x_9813;
wire x_9814;
wire x_9815;
wire x_9816;
wire x_9817;
wire x_9818;
wire x_9819;
wire x_9820;
wire x_9821;
wire x_9822;
wire x_9823;
wire x_9824;
wire x_9825;
wire x_9826;
wire x_9827;
wire x_9828;
wire x_9829;
wire x_9830;
wire x_9831;
wire x_9832;
wire x_9833;
wire x_9834;
wire x_9835;
wire x_9836;
wire x_9837;
wire x_9838;
wire x_9839;
wire x_9840;
wire x_9841;
wire x_9842;
wire x_9843;
wire x_9844;
wire x_9845;
wire x_9846;
wire x_9847;
wire x_9848;
wire x_9849;
wire x_9850;
wire x_9851;
wire x_9852;
wire x_9853;
wire x_9854;
wire x_9855;
wire x_9856;
wire x_9857;
wire x_9858;
wire x_9859;
wire x_9860;
wire x_9861;
wire x_9862;
wire x_9863;
wire x_9864;
wire x_9865;
wire x_9866;
wire x_9867;
wire x_9868;
wire x_9869;
wire x_9870;
wire x_9871;
wire x_9872;
wire x_9873;
wire x_9874;
wire x_9875;
wire x_9876;
wire x_9877;
wire x_9878;
wire x_9879;
wire x_9880;
wire x_9881;
wire x_9882;
wire x_9883;
wire x_9884;
wire x_9885;
wire x_9886;
wire x_9887;
wire x_9888;
wire x_9889;
wire x_9890;
wire x_9891;
wire x_9892;
wire x_9893;
wire x_9894;
wire x_9895;
wire x_9896;
wire x_9897;
wire x_9898;
wire x_9899;
wire x_9900;
wire x_9901;
wire x_9902;
wire x_9903;
wire x_9904;
wire x_9905;
wire x_9906;
wire x_9907;
wire x_9908;
wire x_9909;
wire x_9910;
wire x_9911;
wire x_9912;
wire x_9913;
wire x_9914;
wire x_9915;
wire x_9916;
wire x_9917;
wire x_9918;
wire x_9919;
wire x_9920;
wire x_9921;
wire x_9922;
wire x_9923;
wire x_9924;
wire x_9925;
wire x_9926;
wire x_9927;
wire x_9928;
wire x_9929;
wire x_9930;
wire x_9931;
wire x_9932;
wire x_9933;
wire x_9934;
wire x_9935;
wire x_9936;
wire x_9937;
wire x_9938;
wire x_9939;
wire x_9940;
wire x_9941;
wire x_9942;
wire x_9943;
wire x_9944;
wire x_9945;
wire x_9946;
wire x_9947;
wire x_9948;
wire x_9949;
wire x_9950;
wire x_9951;
wire x_9952;
wire x_9953;
wire x_9954;
wire x_9955;
wire x_9956;
wire x_9957;
wire x_9958;
wire x_9959;
wire x_9960;
wire x_9961;
wire x_9962;
wire x_9963;
wire x_9964;
wire x_9965;
wire x_9966;
wire x_9967;
wire x_9968;
wire x_9969;
wire x_9970;
wire x_9971;
wire x_9972;
wire x_9973;
wire x_9974;
wire x_9975;
wire x_9976;
wire x_9977;
wire x_9978;
wire x_9979;
wire x_9980;
wire x_9981;
wire x_9982;
wire x_9983;
wire x_9984;
wire x_9985;
wire x_9986;
wire x_9987;
wire x_9988;
wire x_9989;
wire x_9990;
wire x_9991;
wire x_9992;
wire x_9993;
wire x_9994;
wire x_9995;
wire x_9996;
wire x_9997;
wire x_9998;
wire x_9999;
wire x_10000;
wire x_10001;
wire x_10002;
wire x_10003;
wire x_10004;
wire x_10005;
wire x_10006;
wire x_10007;
wire x_10008;
wire x_10009;
wire x_10010;
wire x_10011;
wire x_10012;
wire x_10013;
wire x_10014;
wire x_10015;
wire x_10016;
wire x_10017;
wire x_10018;
wire x_10019;
wire x_10020;
wire x_10021;
wire x_10022;
wire x_10023;
wire x_10024;
wire x_10025;
wire x_10026;
wire x_10027;
wire x_10028;
wire x_10029;
wire x_10030;
wire x_10031;
wire x_10032;
wire x_10033;
wire x_10034;
wire x_10035;
wire x_10036;
wire x_10037;
wire x_10038;
wire x_10039;
wire x_10040;
wire x_10041;
wire x_10042;
wire x_10043;
wire x_10044;
wire x_10045;
wire x_10046;
wire x_10047;
wire x_10048;
wire x_10049;
wire x_10050;
wire x_10051;
wire x_10052;
wire x_10053;
wire x_10054;
wire x_10055;
wire x_10056;
wire x_10057;
wire x_10058;
wire x_10059;
wire x_10060;
wire x_10061;
wire x_10062;
wire x_10063;
wire x_10064;
wire x_10065;
wire x_10066;
wire x_10067;
wire x_10068;
wire x_10069;
wire x_10070;
wire x_10071;
wire x_10072;
wire x_10073;
wire x_10074;
wire x_10075;
wire x_10076;
wire x_10077;
wire x_10078;
wire x_10079;
wire x_10080;
wire x_10081;
wire x_10082;
wire x_10083;
wire x_10084;
wire x_10085;
wire x_10086;
wire x_10087;
wire x_10088;
wire x_10089;
wire x_10090;
wire x_10091;
wire x_10092;
wire x_10093;
wire x_10094;
wire x_10095;
wire x_10096;
wire x_10097;
wire x_10098;
wire x_10099;
wire x_10100;
wire x_10101;
wire x_10102;
wire x_10103;
wire x_10104;
wire x_10105;
wire x_10106;
wire x_10107;
wire x_10108;
wire x_10109;
wire x_10110;
wire x_10111;
wire x_10112;
wire x_10113;
wire x_10114;
wire x_10115;
wire x_10116;
wire x_10117;
wire x_10118;
wire x_10119;
wire x_10120;
wire x_10121;
wire x_10122;
wire x_10123;
wire x_10124;
wire x_10125;
wire x_10126;
wire x_10127;
wire x_10128;
wire x_10129;
wire x_10130;
wire x_10131;
wire x_10132;
wire x_10133;
wire x_10134;
wire x_10135;
wire x_10136;
wire x_10137;
wire x_10138;
wire x_10139;
wire x_10140;
wire x_10141;
wire x_10142;
wire x_10143;
wire x_10144;
wire x_10145;
wire x_10146;
wire x_10147;
wire x_10148;
wire x_10149;
wire x_10150;
wire x_10151;
wire x_10152;
wire x_10153;
wire x_10154;
wire x_10155;
wire x_10156;
wire x_10157;
wire x_10158;
wire x_10159;
wire x_10160;
wire x_10161;
wire x_10162;
wire x_10163;
wire x_10164;
wire x_10165;
wire x_10166;
wire x_10167;
wire x_10168;
wire x_10169;
wire x_10170;
wire x_10171;
wire x_10172;
wire x_10173;
wire x_10174;
wire x_10175;
wire x_10176;
wire x_10177;
wire x_10178;
wire x_10179;
wire x_10180;
wire x_10181;
wire x_10182;
wire x_10183;
wire x_10184;
wire x_10185;
wire x_10186;
wire x_10187;
wire x_10188;
wire x_10189;
wire x_10190;
wire x_10191;
wire x_10192;
wire x_10193;
wire x_10194;
wire x_10195;
wire x_10196;
wire x_10197;
wire x_10198;
wire x_10199;
wire x_10200;
wire x_10201;
wire x_10202;
wire x_10203;
wire x_10204;
wire x_10205;
wire x_10206;
wire x_10207;
wire x_10208;
wire x_10209;
wire x_10210;
wire x_10211;
wire x_10212;
wire x_10213;
wire x_10214;
wire x_10215;
wire x_10216;
wire x_10217;
wire x_10218;
wire x_10219;
wire x_10220;
wire x_10221;
wire x_10222;
wire x_10223;
wire x_10224;
wire x_10225;
wire x_10226;
wire x_10227;
wire x_10228;
wire x_10229;
wire x_10230;
wire x_10231;
wire x_10232;
wire x_10233;
wire x_10234;
wire x_10235;
wire x_10236;
wire x_10237;
wire x_10238;
wire x_10239;
wire x_10240;
wire x_10241;
wire x_10242;
wire x_10243;
wire x_10244;
wire x_10245;
wire x_10246;
wire x_10247;
wire x_10248;
wire x_10249;
wire x_10250;
wire x_10251;
wire x_10252;
wire x_10253;
wire x_10254;
wire x_10255;
wire x_10256;
wire x_10257;
wire x_10258;
wire x_10259;
wire x_10260;
wire x_10261;
wire x_10262;
wire x_10263;
wire x_10264;
wire x_10265;
wire x_10266;
wire x_10267;
wire x_10268;
wire x_10269;
wire x_10270;
wire x_10271;
wire x_10272;
wire x_10273;
wire x_10274;
wire x_10275;
wire x_10276;
wire x_10277;
wire x_10278;
wire x_10279;
wire x_10280;
wire x_10281;
wire x_10282;
wire x_10283;
wire x_10284;
wire x_10285;
wire x_10286;
wire x_10287;
wire x_10288;
wire x_10289;
wire x_10290;
wire x_10291;
wire x_10292;
wire x_10293;
wire x_10294;
wire x_10295;
wire x_10296;
wire x_10297;
wire x_10298;
wire x_10299;
wire x_10300;
wire x_10301;
wire x_10302;
wire x_10303;
wire x_10304;
wire x_10305;
wire x_10306;
wire x_10307;
wire x_10308;
wire x_10309;
wire x_10310;
wire x_10311;
wire x_10312;
wire x_10313;
wire x_10314;
wire x_10315;
wire x_10316;
wire x_10317;
wire x_10318;
wire x_10319;
wire x_10320;
wire x_10321;
wire x_10322;
wire x_10323;
wire x_10324;
wire x_10325;
wire x_10326;
wire x_10327;
wire x_10328;
wire x_10329;
wire x_10330;
wire x_10331;
wire x_10332;
wire x_10333;
wire x_10334;
wire x_10335;
wire x_10336;
wire x_10337;
wire x_10338;
wire x_10339;
wire x_10340;
wire x_10341;
wire x_10342;
wire x_10343;
wire x_10344;
wire x_10345;
wire x_10346;
wire x_10347;
wire x_10348;
wire x_10349;
wire x_10350;
wire x_10351;
wire x_10352;
wire x_10353;
wire x_10354;
wire x_10355;
wire x_10356;
wire x_10357;
wire x_10358;
wire x_10359;
wire x_10360;
wire x_10361;
wire x_10362;
wire x_10363;
wire x_10364;
wire x_10365;
wire x_10366;
wire x_10367;
wire x_10368;
wire x_10369;
wire x_10370;
wire x_10371;
wire x_10372;
wire x_10373;
wire x_10374;
wire x_10375;
wire x_10376;
wire x_10377;
wire x_10378;
wire x_10379;
wire x_10380;
wire x_10381;
wire x_10382;
wire x_10383;
wire x_10384;
wire x_10385;
wire x_10386;
wire x_10387;
wire x_10388;
wire x_10389;
wire x_10390;
wire x_10391;
wire x_10392;
wire x_10393;
wire x_10394;
wire x_10395;
wire x_10396;
wire x_10397;
wire x_10398;
wire x_10399;
wire x_10400;
wire x_10401;
wire x_10402;
wire x_10403;
wire x_10404;
wire x_10405;
wire x_10406;
wire x_10407;
wire x_10408;
wire x_10409;
wire x_10410;
wire x_10411;
wire x_10412;
wire x_10413;
wire x_10414;
wire x_10415;
wire x_10416;
wire x_10417;
wire x_10418;
wire x_10419;
wire x_10420;
wire x_10421;
wire x_10422;
wire x_10423;
wire x_10424;
wire x_10425;
wire x_10426;
wire x_10427;
wire x_10428;
wire x_10429;
wire x_10430;
wire x_10431;
wire x_10432;
wire x_10433;
wire x_10434;
wire x_10435;
wire x_10436;
wire x_10437;
wire x_10438;
wire x_10439;
wire x_10440;
wire x_10441;
wire x_10442;
wire x_10443;
wire x_10444;
wire x_10445;
wire x_10446;
wire x_10447;
wire x_10448;
wire x_10449;
wire x_10450;
wire x_10451;
wire x_10452;
wire x_10453;
wire x_10454;
wire x_10455;
wire x_10456;
wire x_10457;
wire x_10458;
wire x_10459;
wire x_10460;
wire x_10461;
wire x_10462;
wire x_10463;
wire x_10464;
wire x_10465;
wire x_10466;
wire x_10467;
wire x_10468;
wire x_10469;
wire x_10470;
wire x_10471;
wire x_10472;
wire x_10473;
wire x_10474;
wire x_10475;
wire x_10476;
wire x_10477;
wire x_10478;
wire x_10479;
wire x_10480;
wire x_10481;
wire x_10482;
wire x_10483;
wire x_10484;
wire x_10485;
wire x_10486;
wire x_10487;
wire x_10488;
wire x_10489;
wire x_10490;
wire x_10491;
wire x_10492;
wire x_10493;
wire x_10494;
wire x_10495;
wire x_10496;
wire x_10497;
wire x_10498;
wire x_10499;
wire x_10500;
wire x_10501;
wire x_10502;
wire x_10503;
wire x_10504;
wire x_10505;
wire x_10506;
wire x_10507;
wire x_10508;
wire x_10509;
wire x_10510;
wire x_10511;
wire x_10512;
wire x_10513;
wire x_10514;
wire x_10515;
wire x_10516;
wire x_10517;
wire x_10518;
wire x_10519;
wire x_10520;
wire x_10521;
wire x_10522;
wire x_10523;
wire x_10524;
wire x_10525;
wire x_10526;
wire x_10527;
wire x_10528;
wire x_10529;
wire x_10530;
wire x_10531;
wire x_10532;
wire x_10533;
wire x_10534;
wire x_10535;
wire x_10536;
wire x_10537;
wire x_10538;
wire x_10539;
wire x_10540;
wire x_10541;
wire x_10542;
wire x_10543;
wire x_10544;
wire x_10545;
wire x_10546;
wire x_10547;
wire x_10548;
wire x_10549;
wire x_10550;
wire x_10551;
wire x_10552;
wire x_10553;
wire x_10554;
wire x_10555;
wire x_10556;
wire x_10557;
wire x_10558;
wire x_10559;
wire x_10560;
wire x_10561;
wire x_10562;
wire x_10563;
wire x_10564;
wire x_10565;
wire x_10566;
wire x_10567;
wire x_10568;
wire x_10569;
wire x_10570;
wire x_10571;
wire x_10572;
wire x_10573;
wire x_10574;
wire x_10575;
wire x_10576;
wire x_10577;
wire x_10578;
wire x_10579;
wire x_10580;
wire x_10581;
wire x_10582;
wire x_10583;
wire x_10584;
wire x_10585;
wire x_10586;
wire x_10587;
wire x_10588;
wire x_10589;
wire x_10590;
wire x_10591;
wire x_10592;
wire x_10593;
wire x_10594;
wire x_10595;
wire x_10596;
wire x_10597;
wire x_10598;
wire x_10599;
wire x_10600;
wire x_10601;
wire x_10602;
wire x_10603;
wire x_10604;
wire x_10605;
wire x_10606;
wire x_10607;
wire x_10608;
wire x_10609;
wire x_10610;
wire x_10611;
wire x_10612;
wire x_10613;
wire x_10614;
wire x_10615;
wire x_10616;
wire x_10617;
wire x_10618;
wire x_10619;
wire x_10620;
wire x_10621;
wire x_10622;
wire x_10623;
wire x_10624;
wire x_10625;
wire x_10626;
wire x_10627;
wire x_10628;
wire x_10629;
wire x_10630;
wire x_10631;
wire x_10632;
wire x_10633;
wire x_10634;
wire x_10635;
wire x_10636;
wire x_10637;
wire x_10638;
wire x_10639;
wire x_10640;
wire x_10641;
wire x_10642;
wire x_10643;
wire x_10644;
wire x_10645;
wire x_10646;
wire x_10647;
wire x_10648;
wire x_10649;
wire x_10650;
wire x_10651;
wire x_10652;
wire x_10653;
wire x_10654;
wire x_10655;
wire x_10656;
wire x_10657;
wire x_10658;
wire x_10659;
wire x_10660;
wire x_10661;
wire x_10662;
wire x_10663;
wire x_10664;
wire x_10665;
wire x_10666;
wire x_10667;
wire x_10668;
wire x_10669;
wire x_10670;
wire x_10671;
wire x_10672;
wire x_10673;
wire x_10674;
wire x_10675;
wire x_10676;
wire x_10677;
wire x_10678;
wire x_10679;
wire x_10680;
wire x_10681;
wire x_10682;
wire x_10683;
wire x_10684;
wire x_10685;
wire x_10686;
wire x_10687;
wire x_10688;
wire x_10689;
wire x_10690;
wire x_10691;
wire x_10692;
wire x_10693;
wire x_10694;
wire x_10695;
wire x_10696;
wire x_10697;
wire x_10698;
wire x_10699;
wire x_10700;
wire x_10701;
wire x_10702;
wire x_10703;
wire x_10704;
wire x_10705;
wire x_10706;
wire x_10707;
wire x_10708;
wire x_10709;
wire x_10710;
wire x_10711;
wire x_10712;
wire x_10713;
wire x_10714;
wire x_10715;
wire x_10716;
wire x_10717;
wire x_10718;
wire x_10719;
wire x_10720;
wire x_10721;
wire x_10722;
wire x_10723;
wire x_10724;
wire x_10725;
wire x_10726;
wire x_10727;
wire x_10728;
wire x_10729;
wire x_10730;
wire x_10731;
wire x_10732;
wire x_10733;
wire x_10734;
wire x_10735;
wire x_10736;
wire x_10737;
wire x_10738;
wire x_10739;
wire x_10740;
wire x_10741;
wire x_10742;
wire x_10743;
wire x_10744;
wire x_10745;
wire x_10746;
wire x_10747;
wire x_10748;
wire x_10749;
wire x_10750;
wire x_10751;
wire x_10752;
wire x_10753;
wire x_10754;
wire x_10755;
wire x_10756;
wire x_10757;
wire x_10758;
wire x_10759;
wire x_10760;
wire x_10761;
wire x_10762;
wire x_10763;
wire x_10764;
wire x_10765;
wire x_10766;
wire x_10767;
wire x_10768;
wire x_10769;
wire x_10770;
wire x_10771;
wire x_10772;
wire x_10773;
wire x_10774;
wire x_10775;
wire x_10776;
wire x_10777;
wire x_10778;
wire x_10779;
wire x_10780;
wire x_10781;
wire x_10782;
wire x_10783;
wire x_10784;
wire x_10785;
wire x_10786;
wire x_10787;
wire x_10788;
wire x_10789;
wire x_10790;
wire x_10791;
wire x_10792;
wire x_10793;
wire x_10794;
wire x_10795;
wire x_10796;
wire x_10797;
wire x_10798;
wire x_10799;
wire x_10800;
wire x_10801;
wire x_10802;
wire x_10803;
wire x_10804;
wire x_10805;
wire x_10806;
wire x_10807;
wire x_10808;
wire x_10809;
wire x_10810;
wire x_10811;
wire x_10812;
wire x_10813;
wire x_10814;
wire x_10815;
wire x_10816;
wire x_10817;
wire x_10818;
wire x_10819;
wire x_10820;
wire x_10821;
wire x_10822;
wire x_10823;
wire x_10824;
wire x_10825;
wire x_10826;
wire x_10827;
wire x_10828;
wire x_10829;
wire x_10830;
wire x_10831;
wire x_10832;
wire x_10833;
wire x_10834;
wire x_10835;
wire x_10836;
wire x_10837;
wire x_10838;
wire x_10839;
wire x_10840;
wire x_10841;
wire x_10842;
wire x_10843;
wire x_10844;
wire x_10845;
wire x_10846;
wire x_10847;
wire x_10848;
wire x_10849;
wire x_10850;
wire x_10851;
wire x_10852;
wire x_10853;
wire x_10854;
wire x_10855;
wire x_10856;
wire x_10857;
wire x_10858;
wire x_10859;
wire x_10860;
wire x_10861;
wire x_10862;
wire x_10863;
wire x_10864;
wire x_10865;
wire x_10866;
wire x_10867;
wire x_10868;
wire x_10869;
wire x_10870;
wire x_10871;
wire x_10872;
wire x_10873;
wire x_10874;
wire x_10875;
wire x_10876;
wire x_10877;
wire x_10878;
wire x_10879;
wire x_10880;
wire x_10881;
wire x_10882;
wire x_10883;
wire x_10884;
wire x_10885;
wire x_10886;
wire x_10887;
wire x_10888;
wire x_10889;
wire x_10890;
wire x_10891;
wire x_10892;
wire x_10893;
wire x_10894;
wire x_10895;
wire x_10896;
wire x_10897;
wire x_10898;
wire x_10899;
wire x_10900;
wire x_10901;
wire x_10902;
wire x_10903;
wire x_10904;
wire x_10905;
wire x_10906;
wire x_10907;
wire x_10908;
wire x_10909;
wire x_10910;
wire x_10911;
wire x_10912;
wire x_10913;
wire x_10914;
wire x_10915;
wire x_10916;
wire x_10917;
wire x_10918;
wire x_10919;
wire x_10920;
wire x_10921;
wire x_10922;
wire x_10923;
wire x_10924;
wire x_10925;
wire x_10926;
wire x_10927;
wire x_10928;
wire x_10929;
wire x_10930;
wire x_10931;
wire x_10932;
wire x_10933;
wire x_10934;
wire x_10935;
wire x_10936;
wire x_10937;
wire x_10938;
wire x_10939;
wire x_10940;
wire x_10941;
wire x_10942;
wire x_10943;
wire x_10944;
wire x_10945;
wire x_10946;
wire x_10947;
wire x_10948;
wire x_10949;
wire x_10950;
wire x_10951;
wire x_10952;
wire x_10953;
wire x_10954;
wire x_10955;
wire x_10956;
wire x_10957;
wire x_10958;
wire x_10959;
wire x_10960;
wire x_10961;
wire x_10962;
wire x_10963;
wire x_10964;
wire x_10965;
wire x_10966;
wire x_10967;
wire x_10968;
wire x_10969;
wire x_10970;
wire x_10971;
wire x_10972;
wire x_10973;
wire x_10974;
wire x_10975;
wire x_10976;
wire x_10977;
wire x_10978;
wire x_10979;
wire x_10980;
wire x_10981;
wire x_10982;
wire x_10983;
wire x_10984;
wire x_10985;
wire x_10986;
wire x_10987;
wire x_10988;
wire x_10989;
wire x_10990;
wire x_10991;
wire x_10992;
wire x_10993;
wire x_10994;
wire x_10995;
wire x_10996;
wire x_10997;
wire x_10998;
wire x_10999;
wire x_11000;
wire x_11001;
wire x_11002;
wire x_11003;
wire x_11004;
wire x_11005;
wire x_11006;
wire x_11007;
wire x_11008;
wire x_11009;
wire x_11010;
wire x_11011;
wire x_11012;
wire x_11013;
wire x_11014;
wire x_11015;
wire x_11016;
wire x_11017;
wire x_11018;
wire x_11019;
wire x_11020;
wire x_11021;
wire x_11022;
wire x_11023;
wire x_11024;
wire x_11025;
wire x_11026;
wire x_11027;
wire x_11028;
wire x_11029;
wire x_11030;
wire x_11031;
wire x_11032;
wire x_11033;
wire x_11034;
wire x_11035;
wire x_11036;
wire x_11037;
wire x_11038;
wire x_11039;
wire x_11040;
wire x_11041;
wire x_11042;
wire x_11043;
wire x_11044;
wire x_11045;
wire x_11046;
wire x_11047;
wire x_11048;
wire x_11049;
wire x_11050;
wire x_11051;
wire x_11052;
wire x_11053;
wire x_11054;
wire x_11055;
wire x_11056;
wire x_11057;
wire x_11058;
wire x_11059;
wire x_11060;
wire x_11061;
wire x_11062;
wire x_11063;
wire x_11064;
wire x_11065;
wire x_11066;
wire x_11067;
wire x_11068;
wire x_11069;
wire x_11070;
wire x_11071;
wire x_11072;
wire x_11073;
wire x_11074;
wire x_11075;
wire x_11076;
wire x_11077;
wire x_11078;
wire x_11079;
wire x_11080;
wire x_11081;
wire x_11082;
wire x_11083;
wire x_11084;
wire x_11085;
wire x_11086;
wire x_11087;
wire x_11088;
wire x_11089;
wire x_11090;
wire x_11091;
wire x_11092;
wire x_11093;
wire x_11094;
wire x_11095;
wire x_11096;
wire x_11097;
wire x_11098;
wire x_11099;
wire x_11100;
wire x_11101;
wire x_11102;
wire x_11103;
wire x_11104;
wire x_11105;
wire x_11106;
wire x_11107;
wire x_11108;
wire x_11109;
wire x_11110;
wire x_11111;
wire x_11112;
wire x_11113;
wire x_11114;
wire x_11115;
wire x_11116;
wire x_11117;
wire x_11118;
wire x_11119;
wire x_11120;
wire x_11121;
wire x_11122;
wire x_11123;
wire x_11124;
wire x_11125;
wire x_11126;
wire x_11127;
wire x_11128;
wire x_11129;
wire x_11130;
wire x_11131;
wire x_11132;
wire x_11133;
wire x_11134;
wire x_11135;
wire x_11136;
wire x_11137;
wire x_11138;
wire x_11139;
wire x_11140;
wire x_11141;
wire x_11142;
wire x_11143;
wire x_11144;
wire x_11145;
wire x_11146;
wire x_11147;
wire x_11148;
wire x_11149;
wire x_11150;
wire x_11151;
wire x_11152;
wire x_11153;
wire x_11154;
wire x_11155;
wire x_11156;
wire x_11157;
wire x_11158;
wire x_11159;
wire x_11160;
wire x_11161;
wire x_11162;
wire x_11163;
wire x_11164;
wire x_11165;
wire x_11166;
wire x_11167;
wire x_11168;
wire x_11169;
wire x_11170;
wire x_11171;
wire x_11172;
wire x_11173;
wire x_11174;
wire x_11175;
wire x_11176;
wire x_11177;
wire x_11178;
wire x_11179;
wire x_11180;
wire x_11181;
wire x_11182;
wire x_11183;
wire x_11184;
wire x_11185;
wire x_11186;
wire x_11187;
wire x_11188;
wire x_11189;
wire x_11190;
wire x_11191;
wire x_11192;
wire x_11193;
wire x_11194;
wire x_11195;
wire x_11196;
wire x_11197;
wire x_11198;
wire x_11199;
wire x_11200;
wire x_11201;
wire x_11202;
wire x_11203;
wire x_11204;
wire x_11205;
wire x_11206;
wire x_11207;
wire x_11208;
wire x_11209;
wire x_11210;
wire x_11211;
wire x_11212;
wire x_11213;
wire x_11214;
wire x_11215;
wire x_11216;
wire x_11217;
wire x_11218;
wire x_11219;
wire x_11220;
wire x_11221;
wire x_11222;
wire x_11223;
wire x_11224;
wire x_11225;
wire x_11226;
wire x_11227;
wire x_11228;
wire x_11229;
wire x_11230;
wire x_11231;
wire x_11232;
wire x_11233;
wire x_11234;
wire x_11235;
wire x_11236;
wire x_11237;
wire x_11238;
wire x_11239;
wire x_11240;
wire x_11241;
wire x_11242;
wire x_11243;
wire x_11244;
wire x_11245;
wire x_11246;
wire x_11247;
wire x_11248;
wire x_11249;
wire x_11250;
wire x_11251;
wire x_11252;
wire x_11253;
wire x_11254;
wire x_11255;
wire x_11256;
wire x_11257;
wire x_11258;
wire x_11259;
wire x_11260;
wire x_11261;
wire x_11262;
wire x_11263;
wire x_11264;
wire x_11265;
wire x_11266;
wire x_11267;
wire x_11268;
wire x_11269;
wire x_11270;
wire x_11271;
wire x_11272;
wire x_11273;
wire x_11274;
wire x_11275;
wire x_11276;
wire x_11277;
wire x_11278;
wire x_11279;
wire x_11280;
wire x_11281;
wire x_11282;
wire x_11283;
wire x_11284;
wire x_11285;
wire x_11286;
wire x_11287;
wire x_11288;
wire x_11289;
wire x_11290;
wire x_11291;
wire x_11292;
wire x_11293;
wire x_11294;
wire x_11295;
wire x_11296;
wire x_11297;
wire x_11298;
wire x_11299;
wire x_11300;
wire x_11301;
wire x_11302;
wire x_11303;
wire x_11304;
wire x_11305;
wire x_11306;
wire x_11307;
wire x_11308;
wire x_11309;
wire x_11310;
wire x_11311;
wire x_11312;
wire x_11313;
wire x_11314;
wire x_11315;
wire x_11316;
wire x_11317;
wire x_11318;
wire x_11319;
wire x_11320;
wire x_11321;
wire x_11322;
wire x_11323;
wire x_11324;
wire x_11325;
wire x_11326;
wire x_11327;
wire x_11328;
wire x_11329;
wire x_11330;
wire x_11331;
wire x_11332;
wire x_11333;
wire x_11334;
wire x_11335;
wire x_11336;
wire x_11337;
wire x_11338;
wire x_11339;
wire x_11340;
wire x_11341;
wire x_11342;
wire x_11343;
wire x_11344;
wire x_11345;
wire x_11346;
wire x_11347;
wire x_11348;
wire x_11349;
wire x_11350;
wire x_11351;
wire x_11352;
wire x_11353;
wire x_11354;
wire x_11355;
wire x_11356;
wire x_11357;
wire x_11358;
wire x_11359;
wire x_11360;
wire x_11361;
wire x_11362;
wire x_11363;
wire x_11364;
wire x_11365;
wire x_11366;
wire x_11367;
wire x_11368;
wire x_11369;
wire x_11370;
wire x_11371;
wire x_11372;
wire x_11373;
wire x_11374;
wire x_11375;
wire x_11376;
wire x_11377;
wire x_11378;
wire x_11379;
wire x_11380;
wire x_11381;
wire x_11382;
wire x_11383;
wire x_11384;
wire x_11385;
wire x_11386;
wire x_11387;
wire x_11388;
wire x_11389;
wire x_11390;
wire x_11391;
wire x_11392;
wire x_11393;
wire x_11394;
wire x_11395;
wire x_11396;
wire x_11397;
wire x_11398;
wire x_11399;
wire x_11400;
wire x_11401;
wire x_11402;
wire x_11403;
wire x_11404;
wire x_11405;
wire x_11406;
wire x_11407;
wire x_11408;
wire x_11409;
wire x_11410;
wire x_11411;
wire x_11412;
wire x_11413;
wire x_11414;
wire x_11415;
wire x_11416;
wire x_11417;
wire x_11418;
wire x_11419;
wire x_11420;
wire x_11421;
wire x_11422;
wire x_11423;
wire x_11424;
wire x_11425;
wire x_11426;
wire x_11427;
wire x_11428;
wire x_11429;
wire x_11430;
wire x_11431;
wire x_11432;
wire x_11433;
wire x_11434;
wire x_11435;
wire x_11436;
wire x_11437;
wire x_11438;
wire x_11439;
wire x_11440;
wire x_11441;
wire x_11442;
wire x_11443;
wire x_11444;
wire x_11445;
wire x_11446;
wire x_11447;
wire x_11448;
wire x_11449;
wire x_11450;
wire x_11451;
wire x_11452;
wire x_11453;
wire x_11454;
wire x_11455;
wire x_11456;
wire x_11457;
wire x_11458;
wire x_11459;
wire x_11460;
wire x_11461;
wire x_11462;
wire x_11463;
wire x_11464;
wire x_11465;
wire x_11466;
wire x_11467;
wire x_11468;
wire x_11469;
wire x_11470;
wire x_11471;
wire x_11472;
wire x_11473;
wire x_11474;
wire x_11475;
wire x_11476;
wire x_11477;
wire x_11478;
wire x_11479;
wire x_11480;
wire x_11481;
wire x_11482;
wire x_11483;
wire x_11484;
wire x_11485;
wire x_11486;
wire x_11487;
wire x_11488;
wire x_11489;
wire x_11490;
wire x_11491;
wire x_11492;
wire x_11493;
wire x_11494;
wire x_11495;
wire x_11496;
wire x_11497;
wire x_11498;
wire x_11499;
wire x_11500;
wire x_11501;
wire x_11502;
wire x_11503;
wire x_11504;
wire x_11505;
wire x_11506;
wire x_11507;
wire x_11508;
wire x_11509;
wire x_11510;
wire x_11511;
wire x_11512;
wire x_11513;
wire x_11514;
wire x_11515;
wire x_11516;
wire x_11517;
wire x_11518;
wire x_11519;
wire x_11520;
wire x_11521;
wire x_11522;
wire x_11523;
wire x_11524;
wire x_11525;
wire x_11526;
wire x_11527;
wire x_11528;
wire x_11529;
wire x_11530;
wire x_11531;
wire x_11532;
wire x_11533;
wire x_11534;
wire x_11535;
wire x_11536;
wire x_11537;
wire x_11538;
wire x_11539;
wire x_11540;
wire x_11541;
wire x_11542;
wire x_11543;
wire x_11544;
wire x_11545;
wire x_11546;
wire x_11547;
wire x_11548;
wire x_11549;
wire x_11550;
wire x_11551;
wire x_11552;
wire x_11553;
wire x_11554;
wire x_11555;
wire x_11556;
wire x_11557;
wire x_11558;
wire x_11559;
wire x_11560;
wire x_11561;
wire x_11562;
wire x_11563;
wire x_11564;
wire x_11565;
wire x_11566;
wire x_11567;
wire x_11568;
wire x_11569;
wire x_11570;
wire x_11571;
wire x_11572;
wire x_11573;
wire x_11574;
wire x_11575;
wire x_11576;
wire x_11577;
wire x_11578;
wire x_11579;
wire x_11580;
wire x_11581;
wire x_11582;
wire x_11583;
wire x_11584;
wire x_11585;
wire x_11586;
wire x_11587;
wire x_11588;
wire x_11589;
wire x_11590;
wire x_11591;
wire x_11592;
wire x_11593;
wire x_11594;
wire x_11595;
wire x_11596;
wire x_11597;
wire x_11598;
wire x_11599;
wire x_11600;
wire x_11601;
wire x_11602;
wire x_11603;
wire x_11604;
wire x_11605;
wire x_11606;
wire x_11607;
wire x_11608;
wire x_11609;
wire x_11610;
wire x_11611;
wire x_11612;
wire x_11613;
wire x_11614;
wire x_11615;
wire x_11616;
wire x_11617;
wire x_11618;
wire x_11619;
wire x_11620;
wire x_11621;
wire x_11622;
wire x_11623;
wire x_11624;
wire x_11625;
wire x_11626;
wire x_11627;
wire x_11628;
wire x_11629;
wire x_11630;
wire x_11631;
wire x_11632;
wire x_11633;
wire x_11634;
wire x_11635;
wire x_11636;
wire x_11637;
wire x_11638;
wire x_11639;
wire x_11640;
wire x_11641;
wire x_11642;
wire x_11643;
wire x_11644;
wire x_11645;
wire x_11646;
wire x_11647;
wire x_11648;
wire x_11649;
wire x_11650;
wire x_11651;
wire x_11652;
wire x_11653;
wire x_11654;
wire x_11655;
wire x_11656;
wire x_11657;
wire x_11658;
wire x_11659;
wire x_11660;
wire x_11661;
wire x_11662;
wire x_11663;
wire x_11664;
wire x_11665;
wire x_11666;
wire x_11667;
wire x_11668;
wire x_11669;
wire x_11670;
wire x_11671;
wire x_11672;
wire x_11673;
wire x_11674;
wire x_11675;
wire x_11676;
wire x_11677;
wire x_11678;
wire x_11679;
wire x_11680;
wire x_11681;
wire x_11682;
wire x_11683;
wire x_11684;
wire x_11685;
wire x_11686;
wire x_11687;
wire x_11688;
wire x_11689;
wire x_11690;
wire x_11691;
wire x_11692;
wire x_11693;
wire x_11694;
wire x_11695;
wire x_11696;
wire x_11697;
wire x_11698;
wire x_11699;
wire x_11700;
wire x_11701;
wire x_11702;
wire x_11703;
wire x_11704;
wire x_11705;
wire x_11706;
wire x_11707;
wire x_11708;
wire x_11709;
wire x_11710;
wire x_11711;
wire x_11712;
wire x_11713;
wire x_11714;
wire x_11715;
wire x_11716;
wire x_11717;
wire x_11718;
wire x_11719;
wire x_11720;
wire x_11721;
wire x_11722;
wire x_11723;
wire x_11724;
wire x_11725;
wire x_11726;
wire x_11727;
wire x_11728;
wire x_11729;
wire x_11730;
wire x_11731;
wire x_11732;
wire x_11733;
wire x_11734;
wire x_11735;
wire x_11736;
wire x_11737;
wire x_11738;
wire x_11739;
wire x_11740;
wire x_11741;
wire x_11742;
wire x_11743;
wire x_11744;
wire x_11745;
wire x_11746;
wire x_11747;
wire x_11748;
wire x_11749;
wire x_11750;
wire x_11751;
wire x_11752;
wire x_11753;
wire x_11754;
wire x_11755;
wire x_11756;
wire x_11757;
wire x_11758;
wire x_11759;
wire x_11760;
wire x_11761;
wire x_11762;
wire x_11763;
wire x_11764;
wire x_11765;
wire x_11766;
wire x_11767;
wire x_11768;
wire x_11769;
wire x_11770;
wire x_11771;
wire x_11772;
wire x_11773;
wire x_11774;
wire x_11775;
wire x_11776;
wire x_11777;
wire x_11778;
wire x_11779;
wire x_11780;
wire x_11781;
wire x_11782;
wire x_11783;
wire x_11784;
wire x_11785;
wire x_11786;
wire x_11787;
wire x_11788;
wire x_11789;
wire x_11790;
wire x_11791;
wire x_11792;
wire x_11793;
wire x_11794;
wire x_11795;
wire x_11796;
wire x_11797;
wire x_11798;
wire x_11799;
wire x_11800;
wire x_11801;
wire x_11802;
wire x_11803;
wire x_11804;
wire x_11805;
wire x_11806;
wire x_11807;
wire x_11808;
wire x_11809;
wire x_11810;
wire x_11811;
wire x_11812;
wire x_11813;
wire x_11814;
wire x_11815;
wire x_11816;
wire x_11817;
wire x_11818;
wire x_11819;
wire x_11820;
wire x_11821;
wire x_11822;
wire x_11823;
wire x_11824;
wire x_11825;
wire x_11826;
wire x_11827;
wire x_11828;
wire x_11829;
wire x_11830;
wire x_11831;
wire x_11832;
wire x_11833;
wire x_11834;
wire x_11835;
wire x_11836;
wire x_11837;
wire x_11838;
wire x_11839;
wire x_11840;
wire x_11841;
wire x_11842;
wire x_11843;
wire x_11844;
wire x_11845;
wire x_11846;
wire x_11847;
wire x_11848;
wire x_11849;
wire x_11850;
wire x_11851;
wire x_11852;
wire x_11853;
wire x_11854;
wire x_11855;
wire x_11856;
wire x_11857;
wire x_11858;
wire x_11859;
wire x_11860;
wire x_11861;
wire x_11862;
wire x_11863;
wire x_11864;
wire x_11865;
wire x_11866;
wire x_11867;
wire x_11868;
wire x_11869;
wire x_11870;
wire x_11871;
wire x_11872;
wire x_11873;
wire x_11874;
wire x_11875;
wire x_11876;
wire x_11877;
wire x_11878;
wire x_11879;
wire x_11880;
wire x_11881;
wire x_11882;
wire x_11883;
wire x_11884;
wire x_11885;
wire x_11886;
wire x_11887;
wire x_11888;
wire x_11889;
wire x_11890;
wire x_11891;
wire x_11892;
wire x_11893;
wire x_11894;
wire x_11895;
wire x_11896;
wire x_11897;
wire x_11898;
wire x_11899;
wire x_11900;
wire x_11901;
wire x_11902;
wire x_11903;
wire x_11904;
wire x_11905;
wire x_11906;
wire x_11907;
wire x_11908;
wire x_11909;
wire x_11910;
wire x_11911;
wire x_11912;
wire x_11913;
wire x_11914;
wire x_11915;
wire x_11916;
wire x_11917;
wire x_11918;
wire x_11919;
wire x_11920;
wire x_11921;
wire x_11922;
wire x_11923;
wire x_11924;
wire x_11925;
wire x_11926;
wire x_11927;
wire x_11928;
wire x_11929;
wire x_11930;
wire x_11931;
wire x_11932;
wire x_11933;
wire x_11934;
wire x_11935;
wire x_11936;
wire x_11937;
wire x_11938;
wire x_11939;
wire x_11940;
wire x_11941;
wire x_11942;
wire x_11943;
wire x_11944;
wire x_11945;
wire x_11946;
wire x_11947;
wire x_11948;
wire x_11949;
wire x_11950;
wire x_11951;
wire x_11952;
wire x_11953;
wire x_11954;
wire x_11955;
wire x_11956;
wire x_11957;
wire x_11958;
wire x_11959;
wire x_11960;
wire x_11961;
wire x_11962;
wire x_11963;
wire x_11964;
wire x_11965;
wire x_11966;
wire x_11967;
wire x_11968;
wire x_11969;
wire x_11970;
wire x_11971;
wire x_11972;
wire x_11973;
wire x_11974;
wire x_11975;
wire x_11976;
wire x_11977;
wire x_11978;
wire x_11979;
wire x_11980;
wire x_11981;
wire x_11982;
wire x_11983;
wire x_11984;
wire x_11985;
wire x_11986;
wire x_11987;
wire x_11988;
wire x_11989;
wire x_11990;
wire x_11991;
wire x_11992;
wire x_11993;
wire x_11994;
wire x_11995;
wire x_11996;
wire x_11997;
wire x_11998;
wire x_11999;
wire x_12000;
wire x_12001;
wire x_12002;
wire x_12003;
wire x_12004;
wire x_12005;
wire x_12006;
wire x_12007;
wire x_12008;
wire x_12009;
wire x_12010;
wire x_12011;
wire x_12012;
wire x_12013;
wire x_12014;
wire x_12015;
wire x_12016;
wire x_12017;
wire x_12018;
wire x_12019;
wire x_12020;
wire x_12021;
wire x_12022;
wire x_12023;
wire x_12024;
wire x_12025;
wire x_12026;
wire x_12027;
wire x_12028;
wire x_12029;
wire x_12030;
wire x_12031;
wire x_12032;
wire x_12033;
wire x_12034;
wire x_12035;
wire x_12036;
wire x_12037;
wire x_12038;
wire x_12039;
wire x_12040;
wire x_12041;
wire x_12042;
wire x_12043;
wire x_12044;
wire x_12045;
wire x_12046;
wire x_12047;
wire x_12048;
wire x_12049;
wire x_12050;
wire x_12051;
wire x_12052;
wire x_12053;
wire x_12054;
wire x_12055;
wire x_12056;
wire x_12057;
wire x_12058;
wire x_12059;
wire x_12060;
wire x_12061;
wire x_12062;
wire x_12063;
wire x_12064;
wire x_12065;
wire x_12066;
wire x_12067;
wire x_12068;
wire x_12069;
wire x_12070;
wire x_12071;
wire x_12072;
wire x_12073;
wire x_12074;
wire x_12075;
wire x_12076;
wire x_12077;
wire x_12078;
wire x_12079;
wire x_12080;
wire x_12081;
wire x_12082;
wire x_12083;
wire x_12084;
wire x_12085;
wire x_12086;
wire x_12087;
wire x_12088;
wire x_12089;
wire x_12090;
wire x_12091;
wire x_12092;
wire x_12093;
wire x_12094;
wire x_12095;
wire x_12096;
wire x_12097;
wire x_12098;
wire x_12099;
wire x_12100;
wire x_12101;
wire x_12102;
wire x_12103;
wire x_12104;
wire x_12105;
wire x_12106;
wire x_12107;
wire x_12108;
wire x_12109;
wire x_12110;
wire x_12111;
wire x_12112;
wire x_12113;
wire x_12114;
wire x_12115;
wire x_12116;
wire x_12117;
wire x_12118;
wire x_12119;
wire x_12120;
wire x_12121;
wire x_12122;
wire x_12123;
wire x_12124;
wire x_12125;
wire x_12126;
wire x_12127;
wire x_12128;
wire x_12129;
wire x_12130;
wire x_12131;
wire x_12132;
wire x_12133;
wire x_12134;
wire x_12135;
wire x_12136;
wire x_12137;
wire x_12138;
wire x_12139;
wire x_12140;
wire x_12141;
wire x_12142;
wire x_12143;
wire x_12144;
wire x_12145;
wire x_12146;
wire x_12147;
wire x_12148;
wire x_12149;
wire x_12150;
wire x_12151;
wire x_12152;
wire x_12153;
wire x_12154;
wire x_12155;
wire x_12156;
wire x_12157;
wire x_12158;
wire x_12159;
wire x_12160;
wire x_12161;
wire x_12162;
wire x_12163;
wire x_12164;
wire x_12165;
wire x_12166;
wire x_12167;
wire x_12168;
wire x_12169;
wire x_12170;
wire x_12171;
wire x_12172;
wire x_12173;
wire x_12174;
wire x_12175;
wire x_12176;
wire x_12177;
wire x_12178;
wire x_12179;
wire x_12180;
wire x_12181;
wire x_12182;
wire x_12183;
wire x_12184;
wire x_12185;
wire x_12186;
wire x_12187;
wire x_12188;
wire x_12189;
wire x_12190;
wire x_12191;
wire x_12192;
wire x_12193;
wire x_12194;
wire x_12195;
wire x_12196;
wire x_12197;
wire x_12198;
wire x_12199;
wire x_12200;
wire x_12201;
wire x_12202;
wire x_12203;
wire x_12204;
wire x_12205;
wire x_12206;
wire x_12207;
wire x_12208;
wire x_12209;
wire x_12210;
wire x_12211;
wire x_12212;
wire x_12213;
wire x_12214;
wire x_12215;
wire x_12216;
wire x_12217;
wire x_12218;
wire x_12219;
wire x_12220;
wire x_12221;
wire x_12222;
wire x_12223;
wire x_12224;
wire x_12225;
wire x_12226;
wire x_12227;
wire x_12228;
wire x_12229;
wire x_12230;
wire x_12231;
wire x_12232;
wire x_12233;
wire x_12234;
wire x_12235;
wire x_12236;
wire x_12237;
wire x_12238;
wire x_12239;
wire x_12240;
wire x_12241;
wire x_12242;
wire x_12243;
wire x_12244;
wire x_12245;
wire x_12246;
wire x_12247;
wire x_12248;
wire x_12249;
wire x_12250;
wire x_12251;
wire x_12252;
wire x_12253;
wire x_12254;
wire x_12255;
wire x_12256;
wire x_12257;
wire x_12258;
wire x_12259;
wire x_12260;
wire x_12261;
wire x_12262;
wire x_12263;
wire x_12264;
wire x_12265;
wire x_12266;
wire x_12267;
wire x_12268;
wire x_12269;
wire x_12270;
wire x_12271;
wire x_12272;
wire x_12273;
wire x_12274;
wire x_12275;
wire x_12276;
wire x_12277;
wire x_12278;
wire x_12279;
wire x_12280;
wire x_12281;
wire x_12282;
wire x_12283;
wire x_12284;
wire x_12285;
wire x_12286;
wire x_12287;
wire x_12288;
wire x_12289;
wire x_12290;
wire x_12291;
wire x_12292;
wire x_12293;
wire x_12294;
wire x_12295;
wire x_12296;
wire x_12297;
wire x_12298;
wire x_12299;
wire x_12300;
wire x_12301;
wire x_12302;
wire x_12303;
wire x_12304;
wire x_12305;
wire x_12306;
wire x_12307;
wire x_12308;
wire x_12309;
wire x_12310;
wire x_12311;
wire x_12312;
wire x_12313;
wire x_12314;
wire x_12315;
wire x_12316;
wire x_12317;
wire x_12318;
wire x_12319;
wire x_12320;
wire x_12321;
wire x_12322;
wire x_12323;
wire x_12324;
wire x_12325;
wire x_12326;
wire x_12327;
wire x_12328;
wire x_12329;
wire x_12330;
wire x_12331;
wire x_12332;
wire x_12333;
wire x_12334;
wire x_12335;
wire x_12336;
wire x_12337;
wire x_12338;
wire x_12339;
wire x_12340;
wire x_12341;
wire x_12342;
wire x_12343;
wire x_12344;
wire x_12345;
wire x_12346;
wire x_12347;
wire x_12348;
wire x_12349;
wire x_12350;
wire x_12351;
wire x_12352;
wire x_12353;
wire x_12354;
wire x_12355;
wire x_12356;
wire x_12357;
wire x_12358;
wire x_12359;
wire x_12360;
wire x_12361;
wire x_12362;
wire x_12363;
wire x_12364;
wire x_12365;
wire x_12366;
wire x_12367;
wire x_12368;
wire x_12369;
wire x_12370;
wire x_12371;
wire x_12372;
wire x_12373;
wire x_12374;
wire x_12375;
wire x_12376;
wire x_12377;
wire x_12378;
wire x_12379;
wire x_12380;
wire x_12381;
wire x_12382;
wire x_12383;
wire x_12384;
wire x_12385;
wire x_12386;
wire x_12387;
wire x_12388;
wire x_12389;
wire x_12390;
wire x_12391;
wire x_12392;
wire x_12393;
wire x_12394;
wire x_12395;
wire x_12396;
wire x_12397;
wire x_12398;
wire x_12399;
wire x_12400;
wire x_12401;
wire x_12402;
wire x_12403;
wire x_12404;
wire x_12405;
wire x_12406;
wire x_12407;
wire x_12408;
wire x_12409;
wire x_12410;
wire x_12411;
wire x_12412;
wire x_12413;
wire x_12414;
wire x_12415;
wire x_12416;
wire x_12417;
wire x_12418;
wire x_12419;
wire x_12420;
wire x_12421;
wire x_12422;
wire x_12423;
wire x_12424;
wire x_12425;
wire x_12426;
wire x_12427;
wire x_12428;
wire x_12429;
wire x_12430;
wire x_12431;
wire x_12432;
wire x_12433;
wire x_12434;
wire x_12435;
wire x_12436;
wire x_12437;
wire x_12438;
wire x_12439;
wire x_12440;
wire x_12441;
wire x_12442;
wire x_12443;
wire x_12444;
wire x_12445;
wire x_12446;
wire x_12447;
wire x_12448;
wire x_12449;
wire x_12450;
wire x_12451;
wire x_12452;
wire x_12453;
wire x_12454;
wire x_12455;
wire x_12456;
wire x_12457;
wire x_12458;
wire x_12459;
wire x_12460;
wire x_12461;
wire x_12462;
wire x_12463;
wire x_12464;
wire x_12465;
wire x_12466;
wire x_12467;
wire x_12468;
wire x_12469;
wire x_12470;
wire x_12471;
wire x_12472;
wire x_12473;
wire x_12474;
wire x_12475;
wire x_12476;
wire x_12477;
wire x_12478;
wire x_12479;
wire x_12480;
wire x_12481;
wire x_12482;
wire x_12483;
wire x_12484;
wire x_12485;
wire x_12486;
wire x_12487;
wire x_12488;
wire x_12489;
wire x_12490;
wire x_12491;
wire x_12492;
wire x_12493;
wire x_12494;
wire x_12495;
wire x_12496;
wire x_12497;
wire x_12498;
wire x_12499;
wire x_12500;
wire x_12501;
wire x_12502;
wire x_12503;
wire x_12504;
wire x_12505;
wire x_12506;
wire x_12507;
wire x_12508;
wire x_12509;
wire x_12510;
wire x_12511;
wire x_12512;
wire x_12513;
wire x_12514;
wire x_12515;
wire x_12516;
wire x_12517;
wire x_12518;
wire x_12519;
wire x_12520;
wire x_12521;
wire x_12522;
wire x_12523;
wire x_12524;
wire x_12525;
wire x_12526;
wire x_12527;
wire x_12528;
wire x_12529;
wire x_12530;
wire x_12531;
wire x_12532;
wire x_12533;
wire x_12534;
wire x_12535;
wire x_12536;
wire x_12537;
wire x_12538;
wire x_12539;
wire x_12540;
wire x_12541;
wire x_12542;
wire x_12543;
wire x_12544;
wire x_12545;
wire x_12546;
wire x_12547;
wire x_12548;
wire x_12549;
wire x_12550;
wire x_12551;
wire x_12552;
wire x_12553;
wire x_12554;
wire x_12555;
wire x_12556;
wire x_12557;
wire x_12558;
wire x_12559;
wire x_12560;
wire x_12561;
wire x_12562;
wire x_12563;
wire x_12564;
wire x_12565;
wire x_12566;
wire x_12567;
wire x_12568;
wire x_12569;
wire x_12570;
wire x_12571;
wire x_12572;
wire x_12573;
wire x_12574;
wire x_12575;
wire x_12576;
wire x_12577;
wire x_12578;
wire x_12579;
wire x_12580;
wire x_12581;
wire x_12582;
wire x_12583;
wire x_12584;
wire x_12585;
wire x_12586;
wire x_12587;
wire x_12588;
wire x_12589;
wire x_12590;
wire x_12591;
wire x_12592;
wire x_12593;
wire x_12594;
wire x_12595;
wire x_12596;
wire x_12597;
wire x_12598;
wire x_12599;
wire x_12600;
wire x_12601;
wire x_12602;
wire x_12603;
wire x_12604;
wire x_12605;
wire x_12606;
wire x_12607;
wire x_12608;
wire x_12609;
wire x_12610;
wire x_12611;
wire x_12612;
wire x_12613;
wire x_12614;
wire x_12615;
wire x_12616;
wire x_12617;
wire x_12618;
wire x_12619;
wire x_12620;
wire x_12621;
wire x_12622;
wire x_12623;
wire x_12624;
wire x_12625;
wire x_12626;
wire x_12627;
wire x_12628;
wire x_12629;
wire x_12630;
wire x_12631;
wire x_12632;
wire x_12633;
wire x_12634;
wire x_12635;
wire x_12636;
wire x_12637;
wire x_12638;
wire x_12639;
wire x_12640;
wire x_12641;
wire x_12642;
wire x_12643;
wire x_12644;
wire x_12645;
wire x_12646;
wire x_12647;
wire x_12648;
wire x_12649;
wire x_12650;
wire x_12651;
wire x_12652;
wire x_12653;
wire x_12654;
wire x_12655;
wire x_12656;
wire x_12657;
wire x_12658;
wire x_12659;
wire x_12660;
wire x_12661;
wire x_12662;
wire x_12663;
wire x_12664;
wire x_12665;
wire x_12666;
wire x_12667;
wire x_12668;
wire x_12669;
wire x_12670;
wire x_12671;
wire x_12672;
wire x_12673;
wire x_12674;
wire x_12675;
wire x_12676;
wire x_12677;
wire x_12678;
wire x_12679;
wire x_12680;
wire x_12681;
wire x_12682;
wire x_12683;
wire x_12684;
wire x_12685;
wire x_12686;
wire x_12687;
wire x_12688;
wire x_12689;
wire x_12690;
wire x_12691;
wire x_12692;
wire x_12693;
wire x_12694;
wire x_12695;
wire x_12696;
wire x_12697;
wire x_12698;
wire x_12699;
wire x_12700;
wire x_12701;
wire x_12702;
wire x_12703;
wire x_12704;
wire x_12705;
wire x_12706;
wire x_12707;
wire x_12708;
wire x_12709;
wire x_12710;
wire x_12711;
wire x_12712;
wire x_12713;
wire x_12714;
wire x_12715;
wire x_12716;
wire x_12717;
wire x_12718;
wire x_12719;
wire x_12720;
wire x_12721;
wire x_12722;
wire x_12723;
wire x_12724;
wire x_12725;
wire x_12726;
wire x_12727;
wire x_12728;
wire x_12729;
wire x_12730;
wire x_12731;
wire x_12732;
wire x_12733;
wire x_12734;
wire x_12735;
wire x_12736;
wire x_12737;
wire x_12738;
wire x_12739;
wire x_12740;
wire x_12741;
wire x_12742;
wire x_12743;
wire x_12744;
wire x_12745;
wire x_12746;
wire x_12747;
wire x_12748;
wire x_12749;
wire x_12750;
wire x_12751;
wire x_12752;
wire x_12753;
wire x_12754;
wire x_12755;
wire x_12756;
wire x_12757;
wire x_12758;
wire x_12759;
wire x_12760;
wire x_12761;
wire x_12762;
wire x_12763;
wire x_12764;
wire x_12765;
wire x_12766;
wire x_12767;
wire x_12768;
wire x_12769;
wire x_12770;
wire x_12771;
wire x_12772;
wire x_12773;
wire x_12774;
wire x_12775;
wire x_12776;
wire x_12777;
wire x_12778;
wire x_12779;
wire x_12780;
wire x_12781;
wire x_12782;
wire x_12783;
wire x_12784;
wire x_12785;
wire x_12786;
wire x_12787;
wire x_12788;
wire x_12789;
wire x_12790;
wire x_12791;
wire x_12792;
wire x_12793;
wire x_12794;
wire x_12795;
wire x_12796;
wire x_12797;
wire x_12798;
wire x_12799;
wire x_12800;
wire x_12801;
wire x_12802;
wire x_12803;
wire x_12804;
wire x_12805;
wire x_12806;
wire x_12807;
wire x_12808;
wire x_12809;
wire x_12810;
wire x_12811;
wire x_12812;
wire x_12813;
wire x_12814;
wire x_12815;
wire x_12816;
wire x_12817;
wire x_12818;
wire x_12819;
wire x_12820;
wire x_12821;
wire x_12822;
wire x_12823;
wire x_12824;
wire x_12825;
wire x_12826;
wire x_12827;
wire x_12828;
wire x_12829;
wire x_12830;
wire x_12831;
wire x_12832;
wire x_12833;
wire x_12834;
wire x_12835;
wire x_12836;
wire x_12837;
wire x_12838;
wire x_12839;
wire x_12840;
wire x_12841;
wire x_12842;
wire x_12843;
wire x_12844;
wire x_12845;
wire x_12846;
wire x_12847;
wire x_12848;
wire x_12849;
wire x_12850;
wire x_12851;
wire x_12852;
wire x_12853;
wire x_12854;
wire x_12855;
wire x_12856;
wire x_12857;
wire x_12858;
wire x_12859;
wire x_12860;
wire x_12861;
wire x_12862;
wire x_12863;
wire x_12864;
wire x_12865;
wire x_12866;
wire x_12867;
wire x_12868;
wire x_12869;
wire x_12870;
wire x_12871;
wire x_12872;
wire x_12873;
wire x_12874;
wire x_12875;
wire x_12876;
wire x_12877;
wire x_12878;
wire x_12879;
wire x_12880;
wire x_12881;
wire x_12882;
wire x_12883;
wire x_12884;
wire x_12885;
wire x_12886;
wire x_12887;
wire x_12888;
wire x_12889;
wire x_12890;
wire x_12891;
wire x_12892;
wire x_12893;
wire x_12894;
wire x_12895;
wire x_12896;
wire x_12897;
wire x_12898;
wire x_12899;
wire x_12900;
wire x_12901;
wire x_12902;
wire x_12903;
wire x_12904;
wire x_12905;
wire x_12906;
wire x_12907;
wire x_12908;
wire x_12909;
wire x_12910;
wire x_12911;
wire x_12912;
wire x_12913;
wire x_12914;
wire x_12915;
wire x_12916;
wire x_12917;
wire x_12918;
wire x_12919;
wire x_12920;
wire x_12921;
wire x_12922;
wire x_12923;
wire x_12924;
wire x_12925;
wire x_12926;
wire x_12927;
wire x_12928;
wire x_12929;
wire x_12930;
wire x_12931;
wire x_12932;
wire x_12933;
wire x_12934;
wire x_12935;
wire x_12936;
wire x_12937;
wire x_12938;
wire x_12939;
wire x_12940;
wire x_12941;
wire x_12942;
wire x_12943;
wire x_12944;
wire x_12945;
wire x_12946;
wire x_12947;
wire x_12948;
wire x_12949;
wire x_12950;
wire x_12951;
wire x_12952;
wire x_12953;
wire x_12954;
wire x_12955;
wire x_12956;
wire x_12957;
wire x_12958;
wire x_12959;
wire x_12960;
wire x_12961;
wire x_12962;
wire x_12963;
wire x_12964;
wire x_12965;
wire x_12966;
wire x_12967;
wire x_12968;
wire x_12969;
wire x_12970;
wire x_12971;
wire x_12972;
wire x_12973;
wire x_12974;
wire x_12975;
wire x_12976;
wire x_12977;
wire x_12978;
wire x_12979;
wire x_12980;
wire x_12981;
wire x_12982;
wire x_12983;
wire x_12984;
wire x_12985;
wire x_12986;
wire x_12987;
wire x_12988;
wire x_12989;
wire x_12990;
wire x_12991;
wire x_12992;
wire x_12993;
wire x_12994;
wire x_12995;
wire x_12996;
wire x_12997;
wire x_12998;
wire x_12999;
wire x_13000;
wire x_13001;
wire x_13002;
wire x_13003;
wire x_13004;
wire x_13005;
wire x_13006;
wire x_13007;
wire x_13008;
wire x_13009;
wire x_13010;
wire x_13011;
wire x_13012;
wire x_13013;
wire x_13014;
wire x_13015;
wire x_13016;
wire x_13017;
wire x_13018;
wire x_13019;
wire x_13020;
wire x_13021;
wire x_13022;
wire x_13023;
wire x_13024;
wire x_13025;
wire x_13026;
wire x_13027;
wire x_13028;
wire x_13029;
wire x_13030;
wire x_13031;
wire x_13032;
wire x_13033;
wire x_13034;
wire x_13035;
wire x_13036;
wire x_13037;
wire x_13038;
wire x_13039;
wire x_13040;
wire x_13041;
wire x_13042;
wire x_13043;
wire x_13044;
wire x_13045;
wire x_13046;
wire x_13047;
wire x_13048;
wire x_13049;
wire x_13050;
wire x_13051;
wire x_13052;
wire x_13053;
wire x_13054;
wire x_13055;
wire x_13056;
wire x_13057;
wire x_13058;
wire x_13059;
wire x_13060;
wire x_13061;
wire x_13062;
wire x_13063;
wire x_13064;
wire x_13065;
wire x_13066;
wire x_13067;
wire x_13068;
wire x_13069;
wire x_13070;
wire x_13071;
wire x_13072;
wire x_13073;
wire x_13074;
wire x_13075;
wire x_13076;
wire x_13077;
wire x_13078;
wire x_13079;
wire x_13080;
wire x_13081;
wire x_13082;
wire x_13083;
wire x_13084;
wire x_13085;
wire x_13086;
wire x_13087;
wire x_13088;
wire x_13089;
wire x_13090;
wire x_13091;
wire x_13092;
wire x_13093;
wire x_13094;
wire x_13095;
wire x_13096;
wire x_13097;
wire x_13098;
wire x_13099;
wire x_13100;
wire x_13101;
wire x_13102;
wire x_13103;
wire x_13104;
wire x_13105;
wire x_13106;
wire x_13107;
wire x_13108;
wire x_13109;
wire x_13110;
wire x_13111;
wire x_13112;
wire x_13113;
wire x_13114;
wire x_13115;
wire x_13116;
wire x_13117;
wire x_13118;
wire x_13119;
wire x_13120;
wire x_13121;
wire x_13122;
wire x_13123;
wire x_13124;
wire x_13125;
wire x_13126;
wire x_13127;
wire x_13128;
wire x_13129;
wire x_13130;
wire x_13131;
wire x_13132;
wire x_13133;
wire x_13134;
wire x_13135;
wire x_13136;
wire x_13137;
wire x_13138;
wire x_13139;
wire x_13140;
wire x_13141;
wire x_13142;
wire x_13143;
wire x_13144;
wire x_13145;
wire x_13146;
wire x_13147;
wire x_13148;
wire x_13149;
wire x_13150;
wire x_13151;
wire x_13152;
wire x_13153;
wire x_13154;
wire x_13155;
wire x_13156;
wire x_13157;
wire x_13158;
wire x_13159;
wire x_13160;
wire x_13161;
wire x_13162;
wire x_13163;
wire x_13164;
wire x_13165;
wire x_13166;
wire x_13167;
wire x_13168;
wire x_13169;
wire x_13170;
wire x_13171;
wire x_13172;
wire x_13173;
wire x_13174;
wire x_13175;
wire x_13176;
wire x_13177;
wire x_13178;
wire x_13179;
wire x_13180;
wire x_13181;
wire x_13182;
wire x_13183;
wire x_13184;
wire x_13185;
wire x_13186;
wire x_13187;
wire x_13188;
wire x_13189;
wire x_13190;
wire x_13191;
wire x_13192;
wire x_13193;
wire x_13194;
wire x_13195;
wire x_13196;
wire x_13197;
wire x_13198;
wire x_13199;
wire x_13200;
wire x_13201;
wire x_13202;
wire x_13203;
wire x_13204;
wire x_13205;
wire x_13206;
wire x_13207;
wire x_13208;
wire x_13209;
wire x_13210;
wire x_13211;
wire x_13212;
wire x_13213;
wire x_13214;
wire x_13215;
wire x_13216;
wire x_13217;
wire x_13218;
wire x_13219;
wire x_13220;
wire x_13221;
wire x_13222;
wire x_13223;
wire x_13224;
wire x_13225;
wire x_13226;
wire x_13227;
wire x_13228;
wire x_13229;
wire x_13230;
wire x_13231;
wire x_13232;
wire x_13233;
wire x_13234;
wire x_13235;
wire x_13236;
wire x_13237;
wire x_13238;
wire x_13239;
wire x_13240;
wire x_13241;
wire x_13242;
wire x_13243;
wire x_13244;
wire x_13245;
wire x_13246;
wire x_13247;
wire x_13248;
wire x_13249;
wire x_13250;
wire x_13251;
wire x_13252;
wire x_13253;
wire x_13254;
wire x_13255;
wire x_13256;
wire x_13257;
wire x_13258;
wire x_13259;
wire x_13260;
wire x_13261;
wire x_13262;
wire x_13263;
wire x_13264;
wire x_13265;
wire x_13266;
wire x_13267;
wire x_13268;
wire x_13269;
wire x_13270;
wire x_13271;
wire x_13272;
wire x_13273;
wire x_13274;
wire x_13275;
wire x_13276;
wire x_13277;
wire x_13278;
wire x_13279;
wire x_13280;
wire x_13281;
wire x_13282;
wire x_13283;
wire x_13284;
wire x_13285;
wire x_13286;
wire x_13287;
wire x_13288;
wire x_13289;
wire x_13290;
wire x_13291;
wire x_13292;
wire x_13293;
wire x_13294;
wire x_13295;
wire x_13296;
wire x_13297;
wire x_13298;
wire x_13299;
wire x_13300;
wire x_13301;
wire x_13302;
wire x_13303;
wire x_13304;
wire x_13305;
wire x_13306;
wire x_13307;
wire x_13308;
wire x_13309;
wire x_13310;
wire x_13311;
wire x_13312;
wire x_13313;
wire x_13314;
wire x_13315;
wire x_13316;
wire x_13317;
wire x_13318;
wire x_13319;
wire x_13320;
wire x_13321;
wire x_13322;
wire x_13323;
wire x_13324;
wire x_13325;
wire x_13326;
wire x_13327;
assign v_1382 = 0;
assign v_1381 = 0;
assign v_1380 = 0;
assign v_1379 = 0;
assign v_1378 = 0;
assign v_1377 = 0;
assign v_1376 = 0;
assign v_1375 = 0;
assign v_1374 = 0;
assign v_1373 = 0;
assign v_1372 = 0;
assign v_1371 = 0;
assign v_1370 = 0;
assign v_1369 = 0;
assign v_1368 = 0;
assign v_1367 = 0;
assign v_1366 = 0;
assign v_1365 = 0;
assign v_1364 = 0;
assign v_1363 = 0;
assign v_1362 = 0;
assign v_1361 = 0;
assign v_1360 = 0;
assign v_1359 = 0;
assign v_1358 = 0;
assign v_1357 = 0;
assign v_1356 = 0;
assign v_1355 = 0;
assign v_1354 = 0;
assign v_1353 = 0;
assign v_1352 = 0;
assign v_1351 = 0;
assign v_1350 = 0;
assign v_1349 = 0;
assign v_1348 = 0;
assign v_1347 = 0;
assign v_1346 = 0;
assign v_1345 = 0;
assign v_1344 = 0;
assign v_1343 = 0;
assign v_1342 = 0;
assign v_1341 = 0;
assign v_1340 = 0;
assign v_1339 = 0;
assign v_1338 = 0;
assign v_1156 = 0;
assign v_1155 = 0;
assign v_1154 = 0;
assign v_1153 = 0;
assign v_1152 = 0;
assign v_1151 = 0;
assign v_1150 = 0;
assign v_1149 = 0;
assign v_1148 = 0;
assign v_1147 = 0;
assign v_1146 = 0;
assign v_1145 = 0;
assign v_1144 = 0;
assign v_1143 = 0;
assign v_1142 = 0;
assign v_1141 = 0;
assign v_1140 = 0;
assign v_1139 = 0;
assign v_1138 = 0;
assign v_1137 = 0;
assign v_1136 = 0;
assign v_1135 = 0;
assign v_1134 = 0;
assign v_1133 = 0;
assign v_1132 = 0;
assign v_1131 = 0;
assign v_1130 = 0;
assign v_1129 = 0;
assign v_1128 = 0;
assign v_1127 = 0;
assign v_1126 = 0;
assign v_1125 = 0;
assign v_1124 = 0;
assign v_1123 = 0;
assign v_1122 = 0;
assign v_1121 = 0;
assign v_1120 = 0;
assign v_1119 = 0;
assign v_1118 = 0;
assign v_1117 = 0;
assign v_1116 = 0;
assign v_1115 = 0;
assign v_1114 = 0;
assign v_1113 = 0;
assign v_1112 = 0;
assign v_930 = 0;
assign v_929 = 0;
assign v_928 = 0;
assign v_927 = 0;
assign v_926 = 0;
assign v_925 = 0;
assign v_924 = 0;
assign v_923 = 0;
assign v_922 = 0;
assign v_921 = 0;
assign v_920 = 0;
assign v_919 = 0;
assign v_918 = 0;
assign v_917 = 0;
assign v_916 = 0;
assign v_915 = 0;
assign v_914 = 0;
assign v_913 = 0;
assign v_912 = 0;
assign v_911 = 0;
assign v_910 = 0;
assign v_909 = 0;
assign v_908 = 0;
assign v_907 = 0;
assign v_906 = 0;
assign v_905 = 0;
assign v_904 = 0;
assign v_903 = 0;
assign v_902 = 0;
assign v_901 = 0;
assign v_900 = 0;
assign v_899 = 0;
assign v_898 = 0;
assign v_897 = 0;
assign v_896 = 0;
assign v_895 = 0;
assign v_894 = 0;
assign v_893 = 0;
assign v_892 = 0;
assign v_891 = 0;
assign v_890 = 0;
assign v_889 = 0;
assign v_888 = 0;
assign v_887 = 0;
assign v_886 = 0;
assign v_704 = 0;
assign v_703 = 0;
assign v_702 = 0;
assign v_701 = 0;
assign v_700 = 0;
assign v_699 = 0;
assign v_698 = 0;
assign v_697 = 0;
assign v_696 = 0;
assign v_695 = 0;
assign v_694 = 0;
assign v_693 = 0;
assign v_692 = 0;
assign v_691 = 0;
assign v_690 = 0;
assign v_689 = 0;
assign v_688 = 0;
assign v_687 = 0;
assign v_686 = 0;
assign v_685 = 0;
assign v_684 = 0;
assign v_683 = 0;
assign v_682 = 0;
assign v_681 = 0;
assign v_680 = 0;
assign v_679 = 0;
assign v_678 = 0;
assign v_677 = 0;
assign v_676 = 0;
assign v_675 = 0;
assign v_674 = 0;
assign v_673 = 0;
assign v_672 = 0;
assign v_671 = 0;
assign v_670 = 0;
assign v_669 = 0;
assign v_668 = 0;
assign v_667 = 0;
assign v_666 = 0;
assign v_665 = 0;
assign v_664 = 0;
assign v_663 = 0;
assign v_662 = 0;
assign v_661 = 0;
assign v_660 = 0;
assign x_1 = v_1383 | v_1384 | v_1385 | v_1386 | v_1387 | v_1388 | v_1389 | v_1390 | v_1391 | v_1392 | v_1393 | v_1394 | v_1395 | v_1396 | v_1397 | v_1398 | v_1399 | v_1400 | v_1401 | v_1402 | v_1403 | v_1404 | v_1405 | v_1406 | v_1407 | v_1408 | v_1409 | v_1410 | v_1411 | v_1412 | v_1413 | v_1414 | v_1415 | v_1416 | v_1417 | v_1418 | v_1419 | v_1420 | v_1421 | v_1422 | v_1423 | v_1424 | v_1425 | v_1426 | v_1427 | v_1428 | v_1429 | v_1430 | v_1431 | v_1432 | v_1433 | v_1434 | v_1435 | v_1436 | v_1437 | v_1438 | v_1439 | v_1440 | v_1441 | v_1442 | v_1443 | v_1444 | v_1445 | v_1446 | v_1447 | v_1448 | v_1449 | v_1450 | v_1451 | v_1452 | v_1453 | v_1454 | v_1455 | v_1456 | v_1457 | v_1458 | v_1459 | v_1460 | v_1461 | v_1462 | v_1463 | v_1464 | v_1465 | v_1466 | v_1467 | v_1468 | v_1469 | v_1470 | v_1471 | v_1472 | v_1473 | v_1474 | v_1475 | v_1476 | v_1477 | v_1478 | v_1479 | v_1480 | v_1481 | v_1482 | v_1483 | v_1484 | v_1485 | v_1486 | v_1487 | v_1488 | v_1489 | v_1490 | v_1491 | v_1492 | v_1493 | v_1494 | v_1495 | v_1496 | v_1497 | v_1498 | v_1499 | v_1500 | v_1501 | v_1502 | v_1503 | v_1504 | v_1505 | v_1506 | v_1507 | v_1508 | v_1509 | v_1510 | v_1511 | v_1512 | v_1513 | v_1514 | v_1515 | v_1516 | v_1517 | v_1518 | v_1519 | v_1520 | v_1521 | v_1522 | v_1523 | v_1524 | v_1525 | v_1526 | v_1527 | v_1528 | v_1529 | v_1530 | v_1531 | v_1532 | v_1533 | v_1534 | v_1535 | v_1536 | v_1537 | v_1538 | v_1539 | v_1540 | v_1541 | v_1542 | v_1543 | v_1544 | v_1545 | v_1546 | v_1547 | v_1548 | v_1549 | v_1550 | v_1551 | v_1552 | v_1553 | v_1554 | v_1555 | v_1556 | v_1557 | v_1558 | v_1559 | v_1560 | v_1561 | v_1562 | v_1563 | v_1564 | v_1565 | v_1566 | v_1567 | v_1568 | v_1569 | v_1570 | v_1571 | v_1572 | v_1573 | v_1574 | v_1575 | v_1576 | v_1577 | v_1578 | v_1579 | v_1580 | v_1581 | v_1582 | v_1583 | v_1584 | v_1585 | v_1586 | v_1587 | v_1588 | v_1589 | v_1590 | v_1591 | v_1592 | v_1593 | v_1594 | v_1595 | v_1596 | v_1597 | v_1598 | v_1599 | v_1600 | v_1601 | v_1602 | v_1603 | v_1604 | v_1605 | v_1606 | v_1607 | v_1608 | v_1609 | v_1610 | v_1611 | v_1612 | v_1613 | v_1614 | v_1615 | v_1616 | v_1617 | v_1618 | v_1619 | v_1620 | v_1621 | v_1622 | v_1623 | v_1624 | v_1625 | v_1626 | v_1627 | v_1628 | v_1629 | v_1630 | v_1631 | v_1632 | v_1633 | v_1634 | v_1635 | v_1636 | v_1637 | v_1638 | v_1639 | v_1640 | v_1641 | v_1642 | v_1643 | v_1644 | v_1645 | v_1646 | v_1647 | v_1648 | v_1649 | v_1650 | v_1651 | v_1652 | v_1653 | v_1654 | v_1655 | v_1656 | v_1657 | v_1658 | v_1659 | v_1660 | v_1661 | v_1662 | v_1663 | v_1664 | v_1665 | v_1666 | v_1667 | v_1668 | v_1669 | v_1670 | v_1671 | v_1672 | v_1673 | v_1674 | v_1675 | v_1676 | v_1677 | v_1678 | v_1679 | v_1680 | v_1681 | v_1682 | v_1683 | v_1684 | v_1685 | v_1686 | v_1687 | v_1688 | v_1689 | v_1690 | v_1691 | v_1692 | v_1693 | v_1694 | v_1695 | v_1696 | v_1697 | v_1698 | v_1699 | v_1700 | v_1701 | v_1702 | v_1703 | v_1704 | v_1705 | v_1706 | v_1707 | v_1708 | v_1709 | v_1710 | v_1711 | v_1712 | v_1713 | v_1714 | v_1715 | v_1716 | v_1717 | v_1718 | v_1719 | v_1720 | v_1721 | v_1722 | v_1723 | v_1724 | v_1725 | v_1726 | v_1727 | v_1728 | v_1729 | v_1730 | v_1731 | v_1732 | v_1733 | v_1734 | v_1735 | v_1736 | v_1737 | v_1738 | v_1739 | v_1740 | v_1741 | v_1742 | v_1743 | v_1744 | v_1745 | v_1746 | v_1747 | v_1748 | v_1749 | v_1750 | v_1751 | v_1752 | v_1753 | v_1754 | v_1755 | v_1756 | v_1757 | v_1758 | v_1759 | v_1760 | v_1761 | v_1762 | v_1763 | v_1764 | v_1765 | v_1766 | v_1767 | v_1768 | v_1769 | v_1770 | v_1771 | v_1772 | v_1773 | v_1774 | v_1775 | v_1776 | v_1777 | v_1778 | v_1779 | v_1780 | v_1781 | v_1782 | v_1783 | v_1784 | v_1785 | v_1786 | v_1787 | v_1788 | v_1789 | v_1790 | v_1791 | v_1792 | v_1793 | v_1794 | v_1795 | v_1796 | v_1797 | v_1798 | v_1799 | v_1800 | v_1801 | v_1802 | v_1803 | v_1804 | v_1805 | v_1806 | v_1807 | v_1808 | v_1809 | v_1810 | v_1811 | v_1812 | v_1813 | v_1814 | v_1815 | v_1816 | v_1817 | v_1818 | v_1819 | v_1820 | v_1821 | v_1822 | v_1823 | v_1824 | v_1825 | v_1826 | v_1827 | v_1828 | v_1829 | v_1830 | v_1831 | v_1832 | v_1833 | v_1834 | v_1835 | v_1836 | v_1837 | v_1838 | v_1839 | v_1840 | v_1841 | v_1842 | v_1843 | v_1844 | v_1845 | v_1846 | v_1847 | v_1848 | v_1849 | v_1850 | v_1851 | v_1852 | v_1853 | v_1854 | v_1855 | v_1856 | v_1857 | v_1858 | v_1859 | v_1860 | v_1861 | v_1862 | v_1863 | v_1864 | v_1865 | v_1866 | v_1867 | v_1868 | v_1869 | v_1870 | v_1871 | v_1872 | v_1873 | v_1874 | v_1875 | v_1876 | v_1877 | v_1878 | v_1879 | v_1880 | v_1881 | v_1882 | v_1883 | v_1884 | v_1885 | v_1886 | v_1887 | v_1888 | v_1889 | v_1890 | v_1891 | v_1892 | v_1893 | v_1894 | v_1895 | v_1896 | v_1897 | v_1898 | v_1899 | v_1900 | v_1901 | v_1902 | v_1903 | v_1904 | v_1905 | v_1906 | v_1907 | v_1908 | v_1909 | v_1910 | v_1911 | v_1912 | v_1913 | v_1914 | v_1915 | v_1916 | v_1917 | v_1918 | v_1919 | v_1920 | v_1921 | v_1922 | v_1923 | v_1924 | v_1925 | v_1926 | v_1927 | v_1928 | v_1929 | v_1930 | v_1931 | v_1932 | v_1933 | v_1934 | v_1935 | v_1936 | v_1937 | v_1938 | v_1939 | v_1940 | v_1941 | v_1942 | v_1943 | v_1944 | v_1945 | v_1946 | v_1947 | v_1948 | v_1949 | v_1950 | v_1951 | v_1952 | v_1953 | v_1954 | v_1955 | v_1956 | v_1957 | v_1958 | v_1959 | v_1960 | v_1961 | v_1962 | v_1963 | v_1964 | v_1965 | v_1966 | v_1967 | v_1968 | v_1969 | v_1970 | v_1971 | v_1972 | v_1973 | v_1974 | v_1975 | v_1976 | v_1977 | v_1978 | v_1979 | v_1980 | v_1981 | v_1982 | v_1983 | v_1984 | v_1985 | v_1986 | v_1987 | v_1988 | v_1989 | v_1990 | v_1991 | v_1992 | v_1993 | v_1994 | v_1995 | v_1996 | v_1997 | v_1998 | v_1999 | v_2000 | v_2001 | v_2002 | v_2003 | v_2004 | v_2005 | v_2006 | v_2007 | v_2008 | v_2009 | v_2010 | v_2011 | v_2012 | v_2013 | v_2014 | v_2015 | v_2016 | v_2017 | v_2018 | v_2019 | v_2020 | v_2021 | v_2022 | v_2023 | v_2024 | v_2025 | v_2026 | v_2027 | v_2028 | v_2029 | v_2030 | v_2031 | v_2032 | v_2033 | v_2034 | v_2035 | v_2036 | v_2037 | v_2038 | v_2039 | v_2040 | v_2041 | v_2042 | v_2043 | v_2044 | v_2045 | v_2046 | v_2047 | v_2048 | v_2049 | v_2050 | v_2051 | v_2052 | v_2053 | v_2054 | v_2055 | v_2056 | v_2057 | v_2058 | v_2059 | v_2060 | v_2061 | v_2062 | v_2063 | v_2064 | v_2065 | v_2066 | v_2067 | v_2068 | v_2069 | v_2070 | v_2071 | v_2072 | v_2073 | v_2074 | v_2075 | v_2076 | v_2077 | v_2078 | v_2079 | v_2080 | v_2081 | v_2082 | v_2083 | v_2084 | v_2085 | v_2086 | v_2087 | v_2088 | v_2089 | v_2090 | v_2091 | v_2092 | v_2093 | v_2094 | v_2095 | v_2096 | v_2097 | v_2098 | v_2099 | v_2100 | v_2101 | v_2102 | v_2103 | v_2104 | v_2105 | v_2106 | v_2107 | v_2108 | v_2109 | v_2110 | v_2111 | v_2112 | v_2113 | v_2114 | v_2115 | v_2116 | v_2117 | v_2118 | v_2119 | v_2120 | v_2121 | v_2122 | v_2123 | v_2124 | v_2125 | v_2126 | v_2127 | v_2128 | v_2129 | v_2130 | v_2131 | v_2132 | v_2133 | v_2134 | v_2135 | v_2136 | v_2137 | v_2138 | v_2139 | v_2140 | v_2141 | v_2142 | v_2143 | v_2144 | v_2145 | v_2146 | v_2147 | v_2148 | v_2149 | v_2150 | v_2151 | v_2152 | v_2153 | v_2154 | v_2155 | v_2156 | v_2157 | v_2158 | v_2159 | v_2160 | v_2161 | v_2162 | v_2163 | v_2164 | v_2165 | v_2166 | v_2167 | v_2168 | v_2169 | v_2170 | v_2171 | v_2172 | v_2173 | v_2174 | v_2175 | v_2176 | v_2177 | v_2178 | v_2179 | v_2180 | v_2181 | v_2182 | v_2183 | v_2184 | v_2185 | v_2186 | v_2187 | v_2188 | v_2189 | v_2190 | v_2191 | v_2192 | v_2193 | v_2194 | v_2195 | v_2196 | v_2197 | v_2198 | v_2199 | v_2200 | v_2201 | v_2202 | v_2203 | v_2204 | v_2205 | v_2206 | v_2207 | v_2208 | v_2209 | v_2210 | v_2211 | v_2212 | v_2213 | v_2214 | v_2215 | v_2216 | v_2217 | v_2218 | v_2219 | v_2220 | v_2221 | v_2222 | v_2223 | v_2224 | v_2225 | v_2226 | v_2227 | v_2228 | v_2229 | v_2230 | v_2231 | v_2232 | v_2233 | v_2234 | v_2235 | v_2236 | v_2237 | v_2238 | v_2239 | v_2240 | v_2241 | v_2242 | v_2243 | v_2244 | v_2245 | v_2246 | v_2247 | v_2248 | v_2249 | v_2250 | v_2251 | v_2252 | v_2253 | v_2254 | v_2255 | v_2256 | v_2257 | v_2258 | v_2259 | v_2260 | v_2261 | v_2262 | v_2263 | v_2264 | v_2265 | v_2266 | v_2267 | v_2268 | v_2269 | v_2270 | v_2271 | v_2272 | v_2273 | v_2274 | v_2275 | v_2276 | v_2277 | v_2278 | v_2279 | v_2280 | v_2281 | v_2282 | v_2283 | v_2284 | v_2285 | v_2286 | v_2287 | v_2288 | v_2289 | v_2290 | v_2291 | v_2292 | v_2293 | v_2294 | v_2295 | v_2296 | v_2297 | v_2298 | v_2299 | v_2300 | v_2301 | v_2302 | v_2303 | v_2304 | v_2305 | v_2306 | v_2307 | v_2308 | v_2309 | v_2310 | v_2311 | v_2312 | v_2313 | v_2314 | v_2315 | v_2316 | v_2317 | v_2318 | v_2319 | v_2320 | v_2321 | v_2322 | v_2323 | v_2324 | v_2325 | v_2326 | v_2327 | v_2328 | v_2329 | v_2330 | v_2331 | v_2332 | v_2333 | v_2334 | v_2335 | v_2336 | v_2337 | v_2338 | v_2339 | v_2340 | v_2341 | v_2342 | v_2343 | v_2344 | v_2345 | v_2346 | v_2347 | v_2348 | v_2349 | v_2350 | v_2351 | v_2352 | v_2353 | v_2354 | v_2355 | v_2356 | v_2357 | v_2358 | v_2359 | v_2360 | v_2361 | v_2362 | v_2363 | v_2364 | v_2365 | v_2366 | v_2367 | v_2368 | v_2369 | v_2370 | v_2371 | v_2372 | v_2373 | v_2374 | v_2375 | v_2376 | v_2377 | v_2378 | v_2379 | v_2380 | v_2381 | v_2382 | v_2383 | v_2384 | v_2385 | v_2386 | v_2387 | v_2388 | v_2389 | v_2390 | v_2391 | v_2392 | v_2393 | v_2394 | v_2395 | v_2396 | v_2397 | v_2398 | v_2399 | v_2400 | v_2401 | v_2402 | v_2403 | v_2404 | v_2405 | v_2406 | v_2407 | v_2408 | v_2409 | v_2410 | v_2411 | v_2412 | v_2413 | v_2414 | v_2415 | v_2416 | v_2417 | v_2418 | v_2419 | v_2420 | v_2421 | v_2422 | v_2423 | v_2424 | v_2425 | v_2426 | v_2427 | v_2428 | v_2429 | v_2430 | v_2431 | v_2432 | v_2433 | v_2434 | v_2435 | v_2436 | v_2437 | v_2438 | v_2439 | v_2440 | v_2441 | v_2442 | v_2443 | v_2444 | v_2445 | v_2446 | v_2447 | v_2448 | v_2449 | v_2450 | v_2451 | v_2452 | v_2453 | v_2454 | v_2455 | v_2456 | v_2457 | v_2458 | v_2459 | v_2460 | v_2461 | v_2462 | v_2463 | v_2464 | v_2465 | v_2466 | v_2467 | v_2468 | v_2469 | v_2470 | v_2471 | v_2472 | v_2473 | v_2474 | v_2475 | v_2476 | v_2477 | v_2478 | v_2479 | v_2480 | v_2481 | v_2482 | v_2483 | v_2484 | v_2485 | v_2486 | v_2487 | v_2488 | v_2489 | v_2490 | v_2491 | v_2492 | v_2493 | v_2494 | v_2495 | v_2496 | v_2497 | v_2498 | v_2499 | v_2500 | v_2501 | v_2502 | v_2503 | v_2504 | v_2505 | v_2506 | v_2507 | v_2508 | v_2509 | v_2510 | v_2511 | v_2512 | v_2513 | v_2514 | v_2515 | v_2516 | v_2517 | v_2518 | v_2519 | v_2520 | v_2521 | v_2522 | v_2523 | v_2524 | v_2525 | v_2526 | v_2527 | v_2528 | v_2529 | v_2530 | v_2531 | v_2532 | v_2533 | v_2534 | v_2535 | v_2536 | v_2537 | v_2538 | v_2539 | v_2540 | v_2541 | v_2542 | v_2543 | v_2544 | v_2545 | v_2546 | v_2547 | v_2548 | v_2549 | v_2550 | v_2551 | v_2552 | v_2553 | v_2554 | v_2555 | v_2556 | v_2557 | v_2558 | v_2559 | v_2560 | v_2561 | v_2562 | v_2563 | v_2564 | v_2565 | v_2566 | v_2567 | v_2568 | v_2569 | v_2570 | v_2571 | v_2572 | v_2573 | v_2574 | v_2575 | v_2576 | v_2577 | v_2578 | v_2579 | v_2580 | v_2581 | v_2582 | v_2583 | v_2584 | v_2585 | v_2586 | v_2587 | v_2588 | v_2589 | v_2590 | v_2591 | v_2592 | v_2593 | v_2594 | v_2595 | v_2596 | v_2597 | v_2598 | v_2599 | v_2600 | v_2601 | v_2602 | v_2603 | v_2604 | v_2605 | v_2606 | v_2607 | v_2608 | v_2609 | v_2610 | v_2611 | v_2612 | v_2613 | v_2614 | v_2615 | v_2616 | v_2617 | v_2618 | v_2619 | v_2620 | v_2621 | v_2622 | v_2623 | v_2624 | v_2625 | v_2626 | v_2627 | v_2628 | v_2629 | v_2630 | v_2631 | v_2632 | v_2633 | v_2634 | v_2635 | v_2636 | v_2637 | v_2638 | v_2639 | v_2640 | v_2641 | v_2642 | v_2643 | v_2644 | v_2645 | v_2646 | v_2647 | v_2648 | v_2649 | v_2650 | v_2651 | v_2652 | v_2653 | v_2654 | v_2655 | v_2656 | v_2657 | v_2658 | v_2659 | v_2660 | v_2661 | v_2662 | v_2663 | v_2664 | v_2665 | v_2666 | v_2667 | v_2668 | v_2669 | v_2670 | v_2671 | v_2672 | v_2673 | v_2674 | v_2675 | v_2676 | v_2677 | v_2678 | v_2679 | v_2680 | v_2681 | v_2682 | v_2683 | v_2684 | v_2685 | v_2686 | v_2687 | v_2688 | v_2689 | v_2690 | v_2691 | v_2692 | v_2693 | v_2694 | v_2695 | v_2696 | v_2697 | v_2698 | v_2699 | v_2700 | v_2701 | v_2702 | v_2703 | v_2704 | v_2705 | v_2706 | v_2707 | v_2708 | v_2709 | v_2710 | v_2711 | v_2712 | v_2713 | v_2714 | v_2715 | v_2716 | v_2717 | v_2718 | v_2719 | v_2720 | v_2721 | v_2722 | v_2723 | v_2724 | v_2725 | v_2726 | v_2727 | v_2728 | v_2729 | v_2730 | v_2731 | v_2732 | v_2733 | v_2734 | v_2735 | v_2736 | v_2737 | v_2738 | v_2739 | v_2740 | v_2741 | v_2742 | v_2743 | v_2744 | v_2745 | v_2746 | v_2747 | v_2748 | v_2749 | v_2750 | v_2751 | v_2752 | v_2753 | v_2754 | v_2755 | v_2756 | v_2757 | v_2758 | v_2759 | v_2760 | v_2761 | v_2762 | v_2763 | v_2764 | v_2765 | v_2766 | v_2767 | v_2768 | v_2769 | v_2770 | v_2771 | v_2772 | v_2773 | v_2774 | v_2775 | v_2776 | v_2777 | v_2778 | v_2779 | v_2780 | v_2781 | v_2782 | v_2783 | v_2784 | v_2785 | v_2786 | v_2787 | v_2788 | v_2789 | v_2790 | v_2791 | v_2792 | v_2793 | v_2794 | v_2795 | v_2796 | v_2797 | v_2798 | v_2799 | v_2800 | v_2801 | v_2802 | v_2803 | v_2804 | v_2805 | v_2806 | v_2807 | v_2808 | v_2809 | v_2810 | v_2811 | v_2812 | v_2813 | v_2814 | v_2815 | v_2816 | v_2817 | v_2818 | v_2819 | v_2820 | v_2821 | v_2822 | v_2823 | v_2824 | v_2825 | v_2826 | v_2827 | v_2828 | v_2829 | v_2830 | v_2831 | v_2832 | v_2833 | v_2834 | v_2835 | v_2836 | v_2837 | v_2838 | v_2839 | v_2840 | v_2841 | v_2842 | v_2843 | v_2844 | v_2845 | v_2846 | v_2847 | v_2848 | v_2849 | v_2850 | v_2851 | v_2852 | v_2853 | v_2854 | v_2855 | v_2856 | v_2857 | v_2858 | v_2859 | v_2860 | v_2861 | v_2862 | v_2863 | v_2864 | v_2865 | v_2866 | v_2867 | v_2868 | v_2869 | v_2870 | v_2871 | v_2872 | v_2873 | v_2874 | v_2875 | v_2876 | v_2877 | v_2878 | v_2879 | v_2880 | v_2881 | v_2882 | v_2883 | v_2884 | v_2885 | v_2886 | v_2887 | v_2888 | v_2889 | v_2890 | v_2891 | v_2892 | v_2893 | v_2894 | v_2895 | v_2896 | v_2897 | v_2898 | v_2899 | v_2900 | v_2901 | v_2902 | v_2903 | v_2904 | v_2905 | v_2906 | v_2907 | v_2908 | v_2909 | v_2910 | v_2911 | v_2912 | v_2913 | v_2914 | v_2915 | v_2916 | v_2917 | v_2918 | v_2919 | v_2920 | v_2921 | v_2922 | v_2923 | v_2924 | v_2925 | v_2926 | v_2927 | v_2928 | v_2929 | v_2930 | v_2931 | v_2932 | v_2933 | v_2934 | v_2935 | v_2936 | v_2937 | v_2938 | v_2939 | v_2940 | v_2941 | v_2942 | v_2943 | v_2944 | v_2945 | v_2946 | v_2947 | v_2948 | v_2949 | v_2950 | v_2951 | v_2952 | v_2953 | v_2954 | v_2955 | v_2956 | v_2957 | v_2958 | v_2959 | v_2960 | v_2961 | v_2962 | v_2963 | v_2964 | v_2965 | v_2966 | v_2967 | v_2968 | v_2969 | v_2970 | v_2971 | v_2972 | v_2973 | v_2974 | v_2975 | v_2976 | v_2977 | v_2978 | v_2979 | v_2980 | v_2981 | v_2982 | v_2983 | v_2984 | v_2985 | v_2986 | v_2987 | v_2988 | v_2989 | v_2990 | v_2991 | v_2992 | v_2993 | v_2994 | v_2995 | v_2996 | v_2997 | v_2998 | v_2999 | v_3000 | v_3001 | v_3002 | v_3003 | v_3004 | v_3005 | v_3006 | v_3007 | v_3008 | v_3009 | v_3010 | v_3011 | v_3012 | v_3013 | v_3014 | v_3015 | v_3016 | v_3017 | v_3018 | v_3019 | v_3020 | v_3021 | v_3022 | v_3023 | v_3024 | v_3025 | v_3026 | v_3027 | v_3028 | v_3029 | v_3030 | v_3031 | v_3032 | v_3033 | v_3034 | v_3035 | v_3036 | v_3037 | v_3038 | v_3039 | v_3040 | v_3041 | v_3042 | v_3043 | v_3044 | v_3045 | v_3046 | v_3047 | v_3048 | v_3049 | v_3050 | v_3051 | v_3052 | v_3053 | v_3054 | v_3055 | v_3056 | v_3057 | v_3058 | v_3059 | v_3060 | v_3061 | v_3062 | v_3063 | v_3064 | v_3065 | v_3066 | v_3067 | v_3068 | v_3069 | v_3070 | v_3071 | v_3072 | v_3073 | v_3074 | v_3075 | v_3076 | v_3077 | v_3078 | v_3079 | v_3080 | v_3081 | v_3082 | v_3083 | v_3084 | v_3085 | v_3086 | v_3087 | v_3088 | v_3089 | v_3090 | v_3091 | v_3092 | v_3093 | v_3094 | v_3095 | v_3096 | v_3097 | v_3098 | v_3099 | v_3100 | v_3101 | v_3102 | v_3103 | v_3104 | v_3105 | v_3106 | v_3107 | v_3108 | v_3109 | v_3110 | v_3111 | v_3112 | v_3113 | v_3114 | v_3115 | v_3116 | v_3117 | v_3118 | v_3119 | v_3120 | v_3121 | v_3122 | v_3123 | v_3124 | v_3125 | v_3126 | v_3127 | v_3128 | v_3129 | v_3130 | v_3131 | v_3132 | v_3133 | v_3134 | v_3135 | v_3136 | v_3137 | v_3138 | v_3139 | v_3140 | v_3141 | v_3142 | v_3143 | v_3144 | v_3145 | v_3146 | v_3147 | v_3148 | v_3149 | v_3150 | v_3151 | v_3152 | v_3153 | v_3154 | v_3155 | v_3156 | v_3157 | v_3158 | v_3159 | v_3160 | v_3161 | v_3162 | v_3163 | v_3164 | v_3165 | v_3166 | v_3167 | v_3168 | v_3169 | v_3170 | v_3171 | v_3172 | v_3173 | v_3174 | v_3175 | v_3176 | v_3177 | v_3178 | v_3179 | v_3180 | v_3181 | v_3182 | v_3183 | v_3184 | v_3185 | v_3186 | v_3187 | v_3188 | v_3189 | v_3190 | v_3191 | v_3192 | v_3193 | v_3194 | v_3195 | v_3196 | v_3197 | v_3198 | v_3199 | v_3200 | v_3201 | v_3202 | v_3203 | v_3204 | v_3205 | v_3206 | v_3207 | v_3208 | v_3209 | v_3210 | v_3211 | v_3212 | v_3213 | v_3214 | v_3215 | v_3216 | v_3217 | v_3218 | v_3219 | v_3220 | v_3221 | v_3222 | v_3223 | v_3224 | v_3225 | v_3226 | v_3227 | v_3228 | v_3229 | v_3230 | v_3231 | v_3232 | v_3233 | v_3234 | v_3235 | v_3236 | v_3237 | v_3238 | v_3239 | v_3240 | v_3241 | v_3242 | v_3243 | v_3244 | v_3245 | v_3246 | v_3247 | v_3248 | v_3249 | v_3250 | v_3251 | v_3252 | v_3253 | v_3254 | v_3255 | v_3256 | v_3257 | v_3258 | v_3259 | v_3260 | v_3261 | v_3262 | v_3263 | v_3264 | v_3265 | v_3266 | v_3267 | v_3268 | v_3269 | v_3270 | v_3271 | v_3272 | v_3273 | v_3274 | v_3275 | v_3276 | v_3277 | v_3278 | v_3279 | v_3280 | v_3281 | v_3282 | v_3283 | v_3284 | v_3285 | v_3286 | v_3287 | v_3288 | v_3289 | v_3290 | v_3291 | v_3292 | v_3293 | v_3294 | v_3295 | v_3296 | v_3297 | v_3298 | v_3299 | v_3300 | v_3301 | v_3302 | v_3303 | v_3304 | v_3305 | v_3306 | v_3307 | v_3308 | v_3309 | v_3310 | v_3311 | v_3312 | v_3313 | v_3314 | v_3315 | v_3316 | v_3317 | v_3318 | v_3319 | v_3320 | v_3321 | v_3322 | v_3323 | v_3324 | v_3325 | v_3326 | v_3327 | v_3328 | v_3329 | v_3330 | v_3331 | v_3332 | v_3333 | v_3334 | v_3335 | v_3336 | v_3337 | v_3338 | v_3339 | v_3340 | v_3341 | v_3342 | v_3343 | v_3344 | v_3345 | v_3346 | v_3347 | v_3348 | v_3349 | v_3350 | v_3351 | v_3352 | v_3353 | v_3354 | v_3355 | v_3356 | v_3357 | v_3358 | v_3359 | v_3360 | v_3361 | v_3362 | v_3363 | v_3364 | v_3365 | v_3366 | v_3367 | v_3368 | v_3369 | v_3370 | v_3371 | v_3372 | v_3373 | v_3374 | v_3375 | v_3376 | v_3377 | v_3378 | v_3379 | v_3380 | v_3381 | v_3382 | v_3383 | v_3384 | v_3385 | v_3386 | v_3387 | v_3388 | v_3389 | v_3390 | v_3391 | v_3392 | v_3393 | v_3394 | v_3395 | v_3396 | v_3397 | v_3398 | v_3399;
assign x_2 = ~v_1383 | v_1337;
assign x_3 = ~v_1384 | v_306;
assign x_4 = ~v_1384 | ~v_307;
assign x_5 = ~v_1385 | v_64;
assign x_6 = ~v_1385 | ~v_307;
assign x_7 = ~v_1386 | v_306;
assign x_8 = ~v_1386 | v_64;
assign x_9 = ~v_1387 | v_305;
assign x_10 = ~v_1387 | ~v_306;
assign x_11 = ~v_1388 | v_63;
assign x_12 = ~v_1388 | ~v_306;
assign x_13 = ~v_1389 | v_305;
assign x_14 = ~v_1389 | v_63;
assign x_15 = ~v_1390 | v_304;
assign x_16 = ~v_1390 | ~v_305;
assign x_17 = ~v_1391 | v_62;
assign x_18 = ~v_1391 | ~v_305;
assign x_19 = ~v_1392 | v_304;
assign x_20 = ~v_1392 | v_62;
assign x_21 = ~v_1393 | v_303;
assign x_22 = ~v_1393 | ~v_304;
assign x_23 = ~v_1394 | v_61;
assign x_24 = ~v_1394 | ~v_304;
assign x_25 = ~v_1395 | v_303;
assign x_26 = ~v_1395 | v_61;
assign x_27 = ~v_1396 | v_302;
assign x_28 = ~v_1396 | ~v_303;
assign x_29 = ~v_1397 | v_60;
assign x_30 = ~v_1397 | ~v_303;
assign x_31 = ~v_1398 | v_302;
assign x_32 = ~v_1398 | v_60;
assign x_33 = ~v_1399 | v_301;
assign x_34 = ~v_1399 | ~v_302;
assign x_35 = ~v_1400 | v_59;
assign x_36 = ~v_1400 | ~v_302;
assign x_37 = ~v_1401 | v_301;
assign x_38 = ~v_1401 | v_59;
assign x_39 = ~v_1402 | v_300;
assign x_40 = ~v_1402 | ~v_301;
assign x_41 = ~v_1403 | v_58;
assign x_42 = ~v_1403 | ~v_301;
assign x_43 = ~v_1404 | v_300;
assign x_44 = ~v_1404 | v_58;
assign x_45 = ~v_1405 | v_56;
assign x_46 = ~v_1405 | ~v_300;
assign x_47 = ~v_1406 | v_57;
assign x_48 = ~v_1406 | ~v_300;
assign x_49 = ~v_1407 | v_56;
assign x_50 = ~v_1407 | v_57;
assign x_51 = ~v_1408 | v_298;
assign x_52 = ~v_1408 | ~v_299;
assign x_53 = ~v_1409 | v_72;
assign x_54 = ~v_1409 | ~v_299;
assign x_55 = ~v_1410 | v_298;
assign x_56 = ~v_1410 | v_72;
assign x_57 = ~v_1411 | v_297;
assign x_58 = ~v_1411 | ~v_298;
assign x_59 = ~v_1412 | v_71;
assign x_60 = ~v_1412 | ~v_298;
assign x_61 = ~v_1413 | v_297;
assign x_62 = ~v_1413 | v_71;
assign x_63 = ~v_1414 | v_296;
assign x_64 = ~v_1414 | ~v_297;
assign x_65 = ~v_1415 | v_70;
assign x_66 = ~v_1415 | ~v_297;
assign x_67 = ~v_1416 | v_296;
assign x_68 = ~v_1416 | v_70;
assign x_69 = ~v_1417 | v_295;
assign x_70 = ~v_1417 | ~v_296;
assign x_71 = ~v_1418 | v_69;
assign x_72 = ~v_1418 | ~v_296;
assign x_73 = ~v_1419 | v_295;
assign x_74 = ~v_1419 | v_69;
assign x_75 = ~v_1420 | v_294;
assign x_76 = ~v_1420 | ~v_295;
assign x_77 = ~v_1421 | v_68;
assign x_78 = ~v_1421 | ~v_295;
assign x_79 = ~v_1422 | v_294;
assign x_80 = ~v_1422 | v_68;
assign x_81 = ~v_1423 | v_293;
assign x_82 = ~v_1423 | ~v_294;
assign x_83 = ~v_1424 | v_67;
assign x_84 = ~v_1424 | ~v_294;
assign x_85 = ~v_1425 | v_293;
assign x_86 = ~v_1425 | v_67;
assign x_87 = ~v_1426 | v_65;
assign x_88 = ~v_1426 | ~v_293;
assign x_89 = ~v_1427 | v_66;
assign x_90 = ~v_1427 | ~v_293;
assign x_91 = ~v_1428 | v_65;
assign x_92 = ~v_1428 | v_66;
assign x_93 = ~v_1429 | v_56;
assign x_94 = ~v_1429 | v_72;
assign x_95 = ~v_1430 | v_56;
assign x_96 = ~v_1430 | v_71;
assign x_97 = ~v_1431 | v_56;
assign x_98 = ~v_1431 | v_70;
assign x_99 = ~v_1432 | v_56;
assign x_100 = ~v_1432 | v_69;
assign x_101 = ~v_1433 | v_56;
assign x_102 = ~v_1433 | v_68;
assign x_103 = ~v_1434 | v_56;
assign x_104 = ~v_1434 | v_67;
assign x_105 = ~v_1435 | v_56;
assign x_106 = ~v_1435 | v_66;
assign x_107 = ~v_1436 | v_56;
assign x_108 = ~v_1436 | v_65;
assign x_109 = ~v_1437 | v_291;
assign x_110 = ~v_1437 | ~v_292;
assign x_111 = ~v_1438 | v_79;
assign x_112 = ~v_1438 | ~v_292;
assign x_113 = ~v_1439 | v_291;
assign x_114 = ~v_1439 | v_79;
assign x_115 = ~v_1440 | v_290;
assign x_116 = ~v_1440 | ~v_291;
assign x_117 = ~v_1441 | v_78;
assign x_118 = ~v_1441 | ~v_291;
assign x_119 = ~v_1442 | v_290;
assign x_120 = ~v_1442 | v_78;
assign x_121 = ~v_1443 | v_289;
assign x_122 = ~v_1443 | ~v_290;
assign x_123 = ~v_1444 | v_77;
assign x_124 = ~v_1444 | ~v_290;
assign x_125 = ~v_1445 | v_289;
assign x_126 = ~v_1445 | v_77;
assign x_127 = ~v_1446 | v_288;
assign x_128 = ~v_1446 | ~v_289;
assign x_129 = ~v_1447 | v_76;
assign x_130 = ~v_1447 | ~v_289;
assign x_131 = ~v_1448 | v_288;
assign x_132 = ~v_1448 | v_76;
assign x_133 = ~v_1449 | v_287;
assign x_134 = ~v_1449 | ~v_288;
assign x_135 = ~v_1450 | v_75;
assign x_136 = ~v_1450 | ~v_288;
assign x_137 = ~v_1451 | v_287;
assign x_138 = ~v_1451 | v_75;
assign x_139 = ~v_1452 | v_73;
assign x_140 = ~v_1452 | ~v_287;
assign x_141 = ~v_1453 | v_74;
assign x_142 = ~v_1453 | ~v_287;
assign x_143 = ~v_1454 | v_73;
assign x_144 = ~v_1454 | v_74;
assign x_145 = ~v_1455 | v_286;
assign x_146 = ~v_1455 | v_79;
assign x_147 = ~v_1456 | v_286;
assign x_148 = ~v_1456 | v_78;
assign x_149 = ~v_1457 | v_286;
assign x_150 = ~v_1457 | v_77;
assign x_151 = ~v_1458 | v_286;
assign x_152 = ~v_1458 | v_76;
assign x_153 = ~v_1459 | v_286;
assign x_154 = ~v_1459 | v_75;
assign x_155 = ~v_1460 | v_286;
assign x_156 = ~v_1460 | v_74;
assign x_157 = ~v_1461 | v_286;
assign x_158 = ~v_1461 | v_73;
assign x_159 = ~v_1462 | v_57;
assign x_160 = ~v_1462 | ~v_286;
assign x_161 = ~v_1463 | v_65;
assign x_162 = ~v_1463 | ~v_286;
assign x_163 = ~v_1464 | v_57;
assign x_164 = ~v_1464 | v_65;
assign x_165 = ~v_1465 | v_284;
assign x_166 = ~v_1465 | ~v_285;
assign x_167 = ~v_1466 | v_85;
assign x_168 = ~v_1466 | ~v_285;
assign x_169 = ~v_1467 | v_284;
assign x_170 = ~v_1467 | v_85;
assign x_171 = ~v_1468 | v_283;
assign x_172 = ~v_1468 | ~v_284;
assign x_173 = ~v_1469 | v_84;
assign x_174 = ~v_1469 | ~v_284;
assign x_175 = ~v_1470 | v_283;
assign x_176 = ~v_1470 | v_84;
assign x_177 = ~v_1471 | v_282;
assign x_178 = ~v_1471 | ~v_283;
assign x_179 = ~v_1472 | v_83;
assign x_180 = ~v_1472 | ~v_283;
assign x_181 = ~v_1473 | v_282;
assign x_182 = ~v_1473 | v_83;
assign x_183 = ~v_1474 | v_281;
assign x_184 = ~v_1474 | ~v_282;
assign x_185 = ~v_1475 | v_82;
assign x_186 = ~v_1475 | ~v_282;
assign x_187 = ~v_1476 | v_281;
assign x_188 = ~v_1476 | v_82;
assign x_189 = ~v_1477 | v_80;
assign x_190 = ~v_1477 | ~v_281;
assign x_191 = ~v_1478 | v_81;
assign x_192 = ~v_1478 | ~v_281;
assign x_193 = ~v_1479 | v_80;
assign x_194 = ~v_1479 | v_81;
assign x_195 = ~v_1480 | v_280;
assign x_196 = ~v_1480 | v_85;
assign x_197 = ~v_1481 | v_280;
assign x_198 = ~v_1481 | v_84;
assign x_199 = ~v_1482 | v_280;
assign x_200 = ~v_1482 | v_83;
assign x_201 = ~v_1483 | v_280;
assign x_202 = ~v_1483 | v_82;
assign x_203 = ~v_1484 | v_280;
assign x_204 = ~v_1484 | v_81;
assign x_205 = ~v_1485 | v_280;
assign x_206 = ~v_1485 | v_80;
assign x_207 = ~v_1486 | v_279;
assign x_208 = ~v_1486 | ~v_280;
assign x_209 = ~v_1487 | v_73;
assign x_210 = ~v_1487 | ~v_280;
assign x_211 = ~v_1488 | v_279;
assign x_212 = ~v_1488 | v_73;
assign x_213 = ~v_1489 | v_58;
assign x_214 = ~v_1489 | ~v_279;
assign x_215 = ~v_1490 | v_66;
assign x_216 = ~v_1490 | ~v_279;
assign x_217 = ~v_1491 | v_58;
assign x_218 = ~v_1491 | v_66;
assign x_219 = ~v_1492 | v_277;
assign x_220 = ~v_1492 | ~v_278;
assign x_221 = ~v_1493 | v_90;
assign x_222 = ~v_1493 | ~v_278;
assign x_223 = ~v_1494 | v_277;
assign x_224 = ~v_1494 | v_90;
assign x_225 = ~v_1495 | v_276;
assign x_226 = ~v_1495 | ~v_277;
assign x_227 = ~v_1496 | v_89;
assign x_228 = ~v_1496 | ~v_277;
assign x_229 = ~v_1497 | v_276;
assign x_230 = ~v_1497 | v_89;
assign x_231 = ~v_1498 | v_275;
assign x_232 = ~v_1498 | ~v_276;
assign x_233 = ~v_1499 | v_88;
assign x_234 = ~v_1499 | ~v_276;
assign x_235 = ~v_1500 | v_275;
assign x_236 = ~v_1500 | v_88;
assign x_237 = ~v_1501 | v_86;
assign x_238 = ~v_1501 | ~v_275;
assign x_239 = ~v_1502 | v_87;
assign x_240 = ~v_1502 | ~v_275;
assign x_241 = ~v_1503 | v_86;
assign x_242 = ~v_1503 | v_87;
assign x_243 = ~v_1504 | v_274;
assign x_244 = ~v_1504 | v_90;
assign x_245 = ~v_1505 | v_274;
assign x_246 = ~v_1505 | v_89;
assign x_247 = ~v_1506 | v_274;
assign x_248 = ~v_1506 | v_88;
assign x_249 = ~v_1507 | v_274;
assign x_250 = ~v_1507 | v_87;
assign x_251 = ~v_1508 | v_274;
assign x_252 = ~v_1508 | v_86;
assign x_253 = ~v_1509 | v_273;
assign x_254 = ~v_1509 | ~v_274;
assign x_255 = ~v_1510 | v_80;
assign x_256 = ~v_1510 | ~v_274;
assign x_257 = ~v_1511 | v_273;
assign x_258 = ~v_1511 | v_80;
assign x_259 = ~v_1512 | v_272;
assign x_260 = ~v_1512 | ~v_273;
assign x_261 = ~v_1513 | v_74;
assign x_262 = ~v_1513 | ~v_273;
assign x_263 = ~v_1514 | v_272;
assign x_264 = ~v_1514 | v_74;
assign x_265 = ~v_1515 | v_59;
assign x_266 = ~v_1515 | ~v_272;
assign x_267 = ~v_1516 | v_67;
assign x_268 = ~v_1516 | ~v_272;
assign x_269 = ~v_1517 | v_59;
assign x_270 = ~v_1517 | v_67;
assign x_271 = ~v_1518 | v_270;
assign x_272 = ~v_1518 | ~v_271;
assign x_273 = ~v_1519 | v_94;
assign x_274 = ~v_1519 | ~v_271;
assign x_275 = ~v_1520 | v_270;
assign x_276 = ~v_1520 | v_94;
assign x_277 = ~v_1521 | v_269;
assign x_278 = ~v_1521 | ~v_270;
assign x_279 = ~v_1522 | v_93;
assign x_280 = ~v_1522 | ~v_270;
assign x_281 = ~v_1523 | v_269;
assign x_282 = ~v_1523 | v_93;
assign x_283 = ~v_1524 | v_91;
assign x_284 = ~v_1524 | ~v_269;
assign x_285 = ~v_1525 | v_92;
assign x_286 = ~v_1525 | ~v_269;
assign x_287 = ~v_1526 | v_91;
assign x_288 = ~v_1526 | v_92;
assign x_289 = ~v_1527 | v_268;
assign x_290 = ~v_1527 | v_94;
assign x_291 = ~v_1528 | v_268;
assign x_292 = ~v_1528 | v_93;
assign x_293 = ~v_1529 | v_268;
assign x_294 = ~v_1529 | v_92;
assign x_295 = ~v_1530 | v_268;
assign x_296 = ~v_1530 | v_91;
assign x_297 = ~v_1531 | v_267;
assign x_298 = ~v_1531 | ~v_268;
assign x_299 = ~v_1532 | v_86;
assign x_300 = ~v_1532 | ~v_268;
assign x_301 = ~v_1533 | v_267;
assign x_302 = ~v_1533 | v_86;
assign x_303 = ~v_1534 | v_266;
assign x_304 = ~v_1534 | ~v_267;
assign x_305 = ~v_1535 | v_81;
assign x_306 = ~v_1535 | ~v_267;
assign x_307 = ~v_1536 | v_266;
assign x_308 = ~v_1536 | v_81;
assign x_309 = ~v_1537 | v_265;
assign x_310 = ~v_1537 | ~v_266;
assign x_311 = ~v_1538 | v_75;
assign x_312 = ~v_1538 | ~v_266;
assign x_313 = ~v_1539 | v_265;
assign x_314 = ~v_1539 | v_75;
assign x_315 = ~v_1540 | v_60;
assign x_316 = ~v_1540 | ~v_265;
assign x_317 = ~v_1541 | v_68;
assign x_318 = ~v_1541 | ~v_265;
assign x_319 = ~v_1542 | v_60;
assign x_320 = ~v_1542 | v_68;
assign x_321 = ~v_1543 | v_263;
assign x_322 = ~v_1543 | ~v_264;
assign x_323 = ~v_1544 | v_97;
assign x_324 = ~v_1544 | ~v_264;
assign x_325 = ~v_1545 | v_263;
assign x_326 = ~v_1545 | v_97;
assign x_327 = ~v_1546 | v_95;
assign x_328 = ~v_1546 | ~v_263;
assign x_329 = ~v_1547 | v_96;
assign x_330 = ~v_1547 | ~v_263;
assign x_331 = ~v_1548 | v_95;
assign x_332 = ~v_1548 | v_96;
assign x_333 = ~v_1549 | v_262;
assign x_334 = ~v_1549 | v_97;
assign x_335 = ~v_1550 | v_262;
assign x_336 = ~v_1550 | v_96;
assign x_337 = ~v_1551 | v_262;
assign x_338 = ~v_1551 | v_95;
assign x_339 = ~v_1552 | v_261;
assign x_340 = ~v_1552 | ~v_262;
assign x_341 = ~v_1553 | v_91;
assign x_342 = ~v_1553 | ~v_262;
assign x_343 = ~v_1554 | v_261;
assign x_344 = ~v_1554 | v_91;
assign x_345 = ~v_1555 | v_260;
assign x_346 = ~v_1555 | ~v_261;
assign x_347 = ~v_1556 | v_87;
assign x_348 = ~v_1556 | ~v_261;
assign x_349 = ~v_1557 | v_260;
assign x_350 = ~v_1557 | v_87;
assign x_351 = ~v_1558 | v_259;
assign x_352 = ~v_1558 | ~v_260;
assign x_353 = ~v_1559 | v_82;
assign x_354 = ~v_1559 | ~v_260;
assign x_355 = ~v_1560 | v_259;
assign x_356 = ~v_1560 | v_82;
assign x_357 = ~v_1561 | v_258;
assign x_358 = ~v_1561 | ~v_259;
assign x_359 = ~v_1562 | v_76;
assign x_360 = ~v_1562 | ~v_259;
assign x_361 = ~v_1563 | v_258;
assign x_362 = ~v_1563 | v_76;
assign x_363 = ~v_1564 | v_61;
assign x_364 = ~v_1564 | ~v_258;
assign x_365 = ~v_1565 | v_69;
assign x_366 = ~v_1565 | ~v_258;
assign x_367 = ~v_1566 | v_61;
assign x_368 = ~v_1566 | v_69;
assign x_369 = ~v_1567 | v_98;
assign x_370 = ~v_1567 | ~v_257;
assign x_371 = ~v_1568 | v_99;
assign x_372 = ~v_1568 | ~v_257;
assign x_373 = ~v_1569 | v_98;
assign x_374 = ~v_1569 | v_99;
assign x_375 = ~v_1570 | v_256;
assign x_376 = ~v_1570 | v_99;
assign x_377 = ~v_1571 | v_256;
assign x_378 = ~v_1571 | v_98;
assign x_379 = ~v_1572 | v_255;
assign x_380 = ~v_1572 | ~v_256;
assign x_381 = ~v_1573 | v_95;
assign x_382 = ~v_1573 | ~v_256;
assign x_383 = ~v_1574 | v_255;
assign x_384 = ~v_1574 | v_95;
assign x_385 = ~v_1575 | v_254;
assign x_386 = ~v_1575 | ~v_255;
assign x_387 = ~v_1576 | v_92;
assign x_388 = ~v_1576 | ~v_255;
assign x_389 = ~v_1577 | v_254;
assign x_390 = ~v_1577 | v_92;
assign x_391 = ~v_1578 | v_253;
assign x_392 = ~v_1578 | ~v_254;
assign x_393 = ~v_1579 | v_88;
assign x_394 = ~v_1579 | ~v_254;
assign x_395 = ~v_1580 | v_253;
assign x_396 = ~v_1580 | v_88;
assign x_397 = ~v_1581 | v_252;
assign x_398 = ~v_1581 | ~v_253;
assign x_399 = ~v_1582 | v_83;
assign x_400 = ~v_1582 | ~v_253;
assign x_401 = ~v_1583 | v_252;
assign x_402 = ~v_1583 | v_83;
assign x_403 = ~v_1584 | v_251;
assign x_404 = ~v_1584 | ~v_252;
assign x_405 = ~v_1585 | v_77;
assign x_406 = ~v_1585 | ~v_252;
assign x_407 = ~v_1586 | v_251;
assign x_408 = ~v_1586 | v_77;
assign x_409 = ~v_1587 | v_62;
assign x_410 = ~v_1587 | ~v_251;
assign x_411 = ~v_1588 | v_70;
assign x_412 = ~v_1588 | ~v_251;
assign x_413 = ~v_1589 | v_62;
assign x_414 = ~v_1589 | v_70;
assign x_415 = ~v_1590 | v_250;
assign x_416 = ~v_1590 | v_100;
assign x_417 = ~v_1591 | v_249;
assign x_418 = ~v_1591 | ~v_250;
assign x_419 = ~v_1592 | v_98;
assign x_420 = ~v_1592 | ~v_250;
assign x_421 = ~v_1593 | v_249;
assign x_422 = ~v_1593 | v_98;
assign x_423 = ~v_1594 | v_248;
assign x_424 = ~v_1594 | ~v_249;
assign x_425 = ~v_1595 | v_96;
assign x_426 = ~v_1595 | ~v_249;
assign x_427 = ~v_1596 | v_248;
assign x_428 = ~v_1596 | v_96;
assign x_429 = ~v_1597 | v_247;
assign x_430 = ~v_1597 | ~v_248;
assign x_431 = ~v_1598 | v_93;
assign x_432 = ~v_1598 | ~v_248;
assign x_433 = ~v_1599 | v_247;
assign x_434 = ~v_1599 | v_93;
assign x_435 = ~v_1600 | v_246;
assign x_436 = ~v_1600 | ~v_247;
assign x_437 = ~v_1601 | v_89;
assign x_438 = ~v_1601 | ~v_247;
assign x_439 = ~v_1602 | v_246;
assign x_440 = ~v_1602 | v_89;
assign x_441 = ~v_1603 | v_245;
assign x_442 = ~v_1603 | ~v_246;
assign x_443 = ~v_1604 | v_84;
assign x_444 = ~v_1604 | ~v_246;
assign x_445 = ~v_1605 | v_245;
assign x_446 = ~v_1605 | v_84;
assign x_447 = ~v_1606 | v_244;
assign x_448 = ~v_1606 | ~v_245;
assign x_449 = ~v_1607 | v_78;
assign x_450 = ~v_1607 | ~v_245;
assign x_451 = ~v_1608 | v_244;
assign x_452 = ~v_1608 | v_78;
assign x_453 = ~v_1609 | v_63;
assign x_454 = ~v_1609 | ~v_244;
assign x_455 = ~v_1610 | v_71;
assign x_456 = ~v_1610 | ~v_244;
assign x_457 = ~v_1611 | v_63;
assign x_458 = ~v_1611 | v_71;
assign x_459 = ~v_1612 | v_242;
assign x_460 = ~v_1612 | ~v_243;
assign x_461 = ~v_1613 | v_100;
assign x_462 = ~v_1613 | ~v_243;
assign x_463 = ~v_1614 | v_242;
assign x_464 = ~v_1614 | v_100;
assign x_465 = ~v_1615 | v_241;
assign x_466 = ~v_1615 | ~v_242;
assign x_467 = ~v_1616 | v_99;
assign x_468 = ~v_1616 | ~v_242;
assign x_469 = ~v_1617 | v_241;
assign x_470 = ~v_1617 | v_99;
assign x_471 = ~v_1618 | v_240;
assign x_472 = ~v_1618 | ~v_241;
assign x_473 = ~v_1619 | v_97;
assign x_474 = ~v_1619 | ~v_241;
assign x_475 = ~v_1620 | v_240;
assign x_476 = ~v_1620 | v_97;
assign x_477 = ~v_1621 | v_239;
assign x_478 = ~v_1621 | ~v_240;
assign x_479 = ~v_1622 | v_94;
assign x_480 = ~v_1622 | ~v_240;
assign x_481 = ~v_1623 | v_239;
assign x_482 = ~v_1623 | v_94;
assign x_483 = ~v_1624 | v_238;
assign x_484 = ~v_1624 | ~v_239;
assign x_485 = ~v_1625 | v_90;
assign x_486 = ~v_1625 | ~v_239;
assign x_487 = ~v_1626 | v_238;
assign x_488 = ~v_1626 | v_90;
assign x_489 = ~v_1627 | v_237;
assign x_490 = ~v_1627 | ~v_238;
assign x_491 = ~v_1628 | v_85;
assign x_492 = ~v_1628 | ~v_238;
assign x_493 = ~v_1629 | v_237;
assign x_494 = ~v_1629 | v_85;
assign x_495 = ~v_1630 | v_236;
assign x_496 = ~v_1630 | ~v_237;
assign x_497 = ~v_1631 | v_79;
assign x_498 = ~v_1631 | ~v_237;
assign x_499 = ~v_1632 | v_236;
assign x_500 = ~v_1632 | v_79;
assign x_501 = ~v_1633 | v_64;
assign x_502 = ~v_1633 | ~v_236;
assign x_503 = ~v_1634 | v_72;
assign x_504 = ~v_1634 | ~v_236;
assign x_505 = ~v_1635 | v_64;
assign x_506 = ~v_1635 | v_72;
assign x_507 = ~v_1636 | v_378;
assign x_508 = ~v_1636 | ~v_379;
assign x_509 = ~v_1637 | v_56;
assign x_510 = ~v_1637 | ~v_379;
assign x_511 = ~v_1638 | v_378;
assign x_512 = ~v_1638 | v_56;
assign x_513 = ~v_1639 | v_377;
assign x_514 = ~v_1639 | ~v_378;
assign x_515 = ~v_1640 | v_57;
assign x_516 = ~v_1640 | ~v_378;
assign x_517 = ~v_1641 | v_377;
assign x_518 = ~v_1641 | v_57;
assign x_519 = ~v_1642 | v_376;
assign x_520 = ~v_1642 | ~v_377;
assign x_521 = ~v_1643 | v_58;
assign x_522 = ~v_1643 | ~v_377;
assign x_523 = ~v_1644 | v_376;
assign x_524 = ~v_1644 | v_58;
assign x_525 = ~v_1645 | v_375;
assign x_526 = ~v_1645 | ~v_376;
assign x_527 = ~v_1646 | v_59;
assign x_528 = ~v_1646 | ~v_376;
assign x_529 = ~v_1647 | v_375;
assign x_530 = ~v_1647 | v_59;
assign x_531 = ~v_1648 | v_374;
assign x_532 = ~v_1648 | ~v_375;
assign x_533 = ~v_1649 | v_60;
assign x_534 = ~v_1649 | ~v_375;
assign x_535 = ~v_1650 | v_374;
assign x_536 = ~v_1650 | v_60;
assign x_537 = ~v_1651 | v_373;
assign x_538 = ~v_1651 | ~v_374;
assign x_539 = ~v_1652 | v_61;
assign x_540 = ~v_1652 | ~v_374;
assign x_541 = ~v_1653 | v_373;
assign x_542 = ~v_1653 | v_61;
assign x_543 = ~v_1654 | v_372;
assign x_544 = ~v_1654 | ~v_373;
assign x_545 = ~v_1655 | v_62;
assign x_546 = ~v_1655 | ~v_373;
assign x_547 = ~v_1656 | v_372;
assign x_548 = ~v_1656 | v_62;
assign x_549 = ~v_1657 | v_64;
assign x_550 = ~v_1657 | ~v_372;
assign x_551 = ~v_1658 | v_63;
assign x_552 = ~v_1658 | ~v_372;
assign x_553 = ~v_1659 | v_64;
assign x_554 = ~v_1659 | v_63;
assign x_555 = ~v_1660 | v_371;
assign x_556 = ~v_1660 | v_56;
assign x_557 = ~v_1661 | v_370;
assign x_558 = ~v_1661 | ~v_371;
assign x_559 = ~v_1662 | v_65;
assign x_560 = ~v_1662 | ~v_371;
assign x_561 = ~v_1663 | v_370;
assign x_562 = ~v_1663 | v_65;
assign x_563 = ~v_1664 | v_369;
assign x_564 = ~v_1664 | ~v_370;
assign x_565 = ~v_1665 | v_66;
assign x_566 = ~v_1665 | ~v_370;
assign x_567 = ~v_1666 | v_369;
assign x_568 = ~v_1666 | v_66;
assign x_569 = ~v_1667 | v_368;
assign x_570 = ~v_1667 | ~v_369;
assign x_571 = ~v_1668 | v_67;
assign x_572 = ~v_1668 | ~v_369;
assign x_573 = ~v_1669 | v_368;
assign x_574 = ~v_1669 | v_67;
assign x_575 = ~v_1670 | v_367;
assign x_576 = ~v_1670 | ~v_368;
assign x_577 = ~v_1671 | v_68;
assign x_578 = ~v_1671 | ~v_368;
assign x_579 = ~v_1672 | v_367;
assign x_580 = ~v_1672 | v_68;
assign x_581 = ~v_1673 | v_366;
assign x_582 = ~v_1673 | ~v_367;
assign x_583 = ~v_1674 | v_69;
assign x_584 = ~v_1674 | ~v_367;
assign x_585 = ~v_1675 | v_366;
assign x_586 = ~v_1675 | v_69;
assign x_587 = ~v_1676 | v_365;
assign x_588 = ~v_1676 | ~v_366;
assign x_589 = ~v_1677 | v_70;
assign x_590 = ~v_1677 | ~v_366;
assign x_591 = ~v_1678 | v_365;
assign x_592 = ~v_1678 | v_70;
assign x_593 = ~v_1679 | v_72;
assign x_594 = ~v_1679 | ~v_365;
assign x_595 = ~v_1680 | v_71;
assign x_596 = ~v_1680 | ~v_365;
assign x_597 = ~v_1681 | v_72;
assign x_598 = ~v_1681 | v_71;
assign x_599 = ~v_1682 | v_364;
assign x_600 = ~v_1682 | v_57;
assign x_601 = ~v_1683 | v_364;
assign x_602 = ~v_1683 | v_65;
assign x_603 = ~v_1684 | v_363;
assign x_604 = ~v_1684 | ~v_364;
assign x_605 = ~v_1685 | v_73;
assign x_606 = ~v_1685 | ~v_364;
assign x_607 = ~v_1686 | v_363;
assign x_608 = ~v_1686 | v_73;
assign x_609 = ~v_1687 | v_362;
assign x_610 = ~v_1687 | ~v_363;
assign x_611 = ~v_1688 | v_74;
assign x_612 = ~v_1688 | ~v_363;
assign x_613 = ~v_1689 | v_362;
assign x_614 = ~v_1689 | v_74;
assign x_615 = ~v_1690 | v_361;
assign x_616 = ~v_1690 | ~v_362;
assign x_617 = ~v_1691 | v_75;
assign x_618 = ~v_1691 | ~v_362;
assign x_619 = ~v_1692 | v_361;
assign x_620 = ~v_1692 | v_75;
assign x_621 = ~v_1693 | v_360;
assign x_622 = ~v_1693 | ~v_361;
assign x_623 = ~v_1694 | v_76;
assign x_624 = ~v_1694 | ~v_361;
assign x_625 = ~v_1695 | v_360;
assign x_626 = ~v_1695 | v_76;
assign x_627 = ~v_1696 | v_359;
assign x_628 = ~v_1696 | ~v_360;
assign x_629 = ~v_1697 | v_77;
assign x_630 = ~v_1697 | ~v_360;
assign x_631 = ~v_1698 | v_359;
assign x_632 = ~v_1698 | v_77;
assign x_633 = ~v_1699 | v_79;
assign x_634 = ~v_1699 | ~v_359;
assign x_635 = ~v_1700 | v_78;
assign x_636 = ~v_1700 | ~v_359;
assign x_637 = ~v_1701 | v_79;
assign x_638 = ~v_1701 | v_78;
assign x_639 = ~v_1702 | v_65;
assign x_640 = ~v_1702 | ~v_358;
assign x_641 = ~v_1703 | v_57;
assign x_642 = ~v_1703 | ~v_358;
assign x_643 = ~v_1704 | v_65;
assign x_644 = ~v_1704 | v_57;
assign x_645 = ~v_1705 | v_357;
assign x_646 = ~v_1705 | v_58;
assign x_647 = ~v_1706 | v_357;
assign x_648 = ~v_1706 | v_66;
assign x_649 = ~v_1707 | v_357;
assign x_650 = ~v_1707 | v_73;
assign x_651 = ~v_1708 | v_356;
assign x_652 = ~v_1708 | ~v_357;
assign x_653 = ~v_1709 | v_80;
assign x_654 = ~v_1709 | ~v_357;
assign x_655 = ~v_1710 | v_356;
assign x_656 = ~v_1710 | v_80;
assign x_657 = ~v_1711 | v_355;
assign x_658 = ~v_1711 | ~v_356;
assign x_659 = ~v_1712 | v_81;
assign x_660 = ~v_1712 | ~v_356;
assign x_661 = ~v_1713 | v_355;
assign x_662 = ~v_1713 | v_81;
assign x_663 = ~v_1714 | v_354;
assign x_664 = ~v_1714 | ~v_355;
assign x_665 = ~v_1715 | v_82;
assign x_666 = ~v_1715 | ~v_355;
assign x_667 = ~v_1716 | v_354;
assign x_668 = ~v_1716 | v_82;
assign x_669 = ~v_1717 | v_353;
assign x_670 = ~v_1717 | ~v_354;
assign x_671 = ~v_1718 | v_83;
assign x_672 = ~v_1718 | ~v_354;
assign x_673 = ~v_1719 | v_353;
assign x_674 = ~v_1719 | v_83;
assign x_675 = ~v_1720 | v_85;
assign x_676 = ~v_1720 | ~v_353;
assign x_677 = ~v_1721 | v_84;
assign x_678 = ~v_1721 | ~v_353;
assign x_679 = ~v_1722 | v_85;
assign x_680 = ~v_1722 | v_84;
assign x_681 = ~v_1723 | v_351;
assign x_682 = ~v_1723 | ~v_352;
assign x_683 = ~v_1724 | v_58;
assign x_684 = ~v_1724 | ~v_352;
assign x_685 = ~v_1725 | v_351;
assign x_686 = ~v_1725 | v_58;
assign x_687 = ~v_1726 | v_73;
assign x_688 = ~v_1726 | ~v_351;
assign x_689 = ~v_1727 | v_66;
assign x_690 = ~v_1727 | ~v_351;
assign x_691 = ~v_1728 | v_73;
assign x_692 = ~v_1728 | v_66;
assign x_693 = ~v_1729 | v_350;
assign x_694 = ~v_1729 | v_59;
assign x_695 = ~v_1730 | v_350;
assign x_696 = ~v_1730 | v_67;
assign x_697 = ~v_1731 | v_350;
assign x_698 = ~v_1731 | v_74;
assign x_699 = ~v_1732 | v_350;
assign x_700 = ~v_1732 | v_80;
assign x_701 = ~v_1733 | v_349;
assign x_702 = ~v_1733 | ~v_350;
assign x_703 = ~v_1734 | v_86;
assign x_704 = ~v_1734 | ~v_350;
assign x_705 = ~v_1735 | v_349;
assign x_706 = ~v_1735 | v_86;
assign x_707 = ~v_1736 | v_348;
assign x_708 = ~v_1736 | ~v_349;
assign x_709 = ~v_1737 | v_87;
assign x_710 = ~v_1737 | ~v_349;
assign x_711 = ~v_1738 | v_348;
assign x_712 = ~v_1738 | v_87;
assign x_713 = ~v_1739 | v_347;
assign x_714 = ~v_1739 | ~v_348;
assign x_715 = ~v_1740 | v_88;
assign x_716 = ~v_1740 | ~v_348;
assign x_717 = ~v_1741 | v_347;
assign x_718 = ~v_1741 | v_88;
assign x_719 = ~v_1742 | v_90;
assign x_720 = ~v_1742 | ~v_347;
assign x_721 = ~v_1743 | v_89;
assign x_722 = ~v_1743 | ~v_347;
assign x_723 = ~v_1744 | v_90;
assign x_724 = ~v_1744 | v_89;
assign x_725 = ~v_1745 | v_345;
assign x_726 = ~v_1745 | ~v_346;
assign x_727 = ~v_1746 | v_59;
assign x_728 = ~v_1746 | ~v_346;
assign x_729 = ~v_1747 | v_345;
assign x_730 = ~v_1747 | v_59;
assign x_731 = ~v_1748 | v_344;
assign x_732 = ~v_1748 | ~v_345;
assign x_733 = ~v_1749 | v_67;
assign x_734 = ~v_1749 | ~v_345;
assign x_735 = ~v_1750 | v_344;
assign x_736 = ~v_1750 | v_67;
assign x_737 = ~v_1751 | v_80;
assign x_738 = ~v_1751 | ~v_344;
assign x_739 = ~v_1752 | v_74;
assign x_740 = ~v_1752 | ~v_344;
assign x_741 = ~v_1753 | v_80;
assign x_742 = ~v_1753 | v_74;
assign x_743 = ~v_1754 | v_343;
assign x_744 = ~v_1754 | v_60;
assign x_745 = ~v_1755 | v_343;
assign x_746 = ~v_1755 | v_68;
assign x_747 = ~v_1756 | v_343;
assign x_748 = ~v_1756 | v_75;
assign x_749 = ~v_1757 | v_343;
assign x_750 = ~v_1757 | v_81;
assign x_751 = ~v_1758 | v_343;
assign x_752 = ~v_1758 | v_86;
assign x_753 = ~v_1759 | v_342;
assign x_754 = ~v_1759 | ~v_343;
assign x_755 = ~v_1760 | v_91;
assign x_756 = ~v_1760 | ~v_343;
assign x_757 = ~v_1761 | v_342;
assign x_758 = ~v_1761 | v_91;
assign x_759 = ~v_1762 | v_341;
assign x_760 = ~v_1762 | ~v_342;
assign x_761 = ~v_1763 | v_92;
assign x_762 = ~v_1763 | ~v_342;
assign x_763 = ~v_1764 | v_341;
assign x_764 = ~v_1764 | v_92;
assign x_765 = ~v_1765 | v_94;
assign x_766 = ~v_1765 | ~v_341;
assign x_767 = ~v_1766 | v_93;
assign x_768 = ~v_1766 | ~v_341;
assign x_769 = ~v_1767 | v_94;
assign x_770 = ~v_1767 | v_93;
assign x_771 = ~v_1768 | v_339;
assign x_772 = ~v_1768 | ~v_340;
assign x_773 = ~v_1769 | v_60;
assign x_774 = ~v_1769 | ~v_340;
assign x_775 = ~v_1770 | v_339;
assign x_776 = ~v_1770 | v_60;
assign x_777 = ~v_1771 | v_338;
assign x_778 = ~v_1771 | ~v_339;
assign x_779 = ~v_1772 | v_68;
assign x_780 = ~v_1772 | ~v_339;
assign x_781 = ~v_1773 | v_338;
assign x_782 = ~v_1773 | v_68;
assign x_783 = ~v_1774 | v_337;
assign x_784 = ~v_1774 | ~v_338;
assign x_785 = ~v_1775 | v_75;
assign x_786 = ~v_1775 | ~v_338;
assign x_787 = ~v_1776 | v_337;
assign x_788 = ~v_1776 | v_75;
assign x_789 = ~v_1777 | v_86;
assign x_790 = ~v_1777 | ~v_337;
assign x_791 = ~v_1778 | v_81;
assign x_792 = ~v_1778 | ~v_337;
assign x_793 = ~v_1779 | v_86;
assign x_794 = ~v_1779 | v_81;
assign x_795 = ~v_1780 | v_336;
assign x_796 = ~v_1780 | v_61;
assign x_797 = ~v_1781 | v_336;
assign x_798 = ~v_1781 | v_69;
assign x_799 = ~v_1782 | v_336;
assign x_800 = ~v_1782 | v_76;
assign x_801 = ~v_1783 | v_336;
assign x_802 = ~v_1783 | v_82;
assign x_803 = ~v_1784 | v_336;
assign x_804 = ~v_1784 | v_87;
assign x_805 = ~v_1785 | v_336;
assign x_806 = ~v_1785 | v_91;
assign x_807 = ~v_1786 | v_335;
assign x_808 = ~v_1786 | ~v_336;
assign x_809 = ~v_1787 | v_95;
assign x_810 = ~v_1787 | ~v_336;
assign x_811 = ~v_1788 | v_335;
assign x_812 = ~v_1788 | v_95;
assign x_813 = ~v_1789 | v_97;
assign x_814 = ~v_1789 | ~v_335;
assign x_815 = ~v_1790 | v_96;
assign x_816 = ~v_1790 | ~v_335;
assign x_817 = ~v_1791 | v_97;
assign x_818 = ~v_1791 | v_96;
assign x_819 = ~v_1792 | v_333;
assign x_820 = ~v_1792 | ~v_334;
assign x_821 = ~v_1793 | v_61;
assign x_822 = ~v_1793 | ~v_334;
assign x_823 = ~v_1794 | v_333;
assign x_824 = ~v_1794 | v_61;
assign x_825 = ~v_1795 | v_332;
assign x_826 = ~v_1795 | ~v_333;
assign x_827 = ~v_1796 | v_69;
assign x_828 = ~v_1796 | ~v_333;
assign x_829 = ~v_1797 | v_332;
assign x_830 = ~v_1797 | v_69;
assign x_831 = ~v_1798 | v_331;
assign x_832 = ~v_1798 | ~v_332;
assign x_833 = ~v_1799 | v_76;
assign x_834 = ~v_1799 | ~v_332;
assign x_835 = ~v_1800 | v_331;
assign x_836 = ~v_1800 | v_76;
assign x_837 = ~v_1801 | v_330;
assign x_838 = ~v_1801 | ~v_331;
assign x_839 = ~v_1802 | v_82;
assign x_840 = ~v_1802 | ~v_331;
assign x_841 = ~v_1803 | v_330;
assign x_842 = ~v_1803 | v_82;
assign x_843 = ~v_1804 | v_91;
assign x_844 = ~v_1804 | ~v_330;
assign x_845 = ~v_1805 | v_87;
assign x_846 = ~v_1805 | ~v_330;
assign x_847 = ~v_1806 | v_91;
assign x_848 = ~v_1806 | v_87;
assign x_849 = ~v_1807 | v_329;
assign x_850 = ~v_1807 | v_62;
assign x_851 = ~v_1808 | v_329;
assign x_852 = ~v_1808 | v_70;
assign x_853 = ~v_1809 | v_329;
assign x_854 = ~v_1809 | v_77;
assign x_855 = ~v_1810 | v_329;
assign x_856 = ~v_1810 | v_83;
assign x_857 = ~v_1811 | v_329;
assign x_858 = ~v_1811 | v_88;
assign x_859 = ~v_1812 | v_329;
assign x_860 = ~v_1812 | v_92;
assign x_861 = ~v_1813 | v_329;
assign x_862 = ~v_1813 | v_95;
assign x_863 = ~v_1814 | v_99;
assign x_864 = ~v_1814 | ~v_329;
assign x_865 = ~v_1815 | v_98;
assign x_866 = ~v_1815 | ~v_329;
assign x_867 = ~v_1816 | v_99;
assign x_868 = ~v_1816 | v_98;
assign x_869 = ~v_1817 | v_327;
assign x_870 = ~v_1817 | ~v_328;
assign x_871 = ~v_1818 | v_62;
assign x_872 = ~v_1818 | ~v_328;
assign x_873 = ~v_1819 | v_327;
assign x_874 = ~v_1819 | v_62;
assign x_875 = ~v_1820 | v_326;
assign x_876 = ~v_1820 | ~v_327;
assign x_877 = ~v_1821 | v_70;
assign x_878 = ~v_1821 | ~v_327;
assign x_879 = ~v_1822 | v_326;
assign x_880 = ~v_1822 | v_70;
assign x_881 = ~v_1823 | v_325;
assign x_882 = ~v_1823 | ~v_326;
assign x_883 = ~v_1824 | v_77;
assign x_884 = ~v_1824 | ~v_326;
assign x_885 = ~v_1825 | v_325;
assign x_886 = ~v_1825 | v_77;
assign x_887 = ~v_1826 | v_324;
assign x_888 = ~v_1826 | ~v_325;
assign x_889 = ~v_1827 | v_83;
assign x_890 = ~v_1827 | ~v_325;
assign x_891 = ~v_1828 | v_324;
assign x_892 = ~v_1828 | v_83;
assign x_893 = ~v_1829 | v_323;
assign x_894 = ~v_1829 | ~v_324;
assign x_895 = ~v_1830 | v_88;
assign x_896 = ~v_1830 | ~v_324;
assign x_897 = ~v_1831 | v_323;
assign x_898 = ~v_1831 | v_88;
assign x_899 = ~v_1832 | v_95;
assign x_900 = ~v_1832 | ~v_323;
assign x_901 = ~v_1833 | v_92;
assign x_902 = ~v_1833 | ~v_323;
assign x_903 = ~v_1834 | v_95;
assign x_904 = ~v_1834 | v_92;
assign x_905 = ~v_1835 | v_100;
assign x_906 = ~v_1835 | v_63;
assign x_907 = ~v_1836 | v_100;
assign x_908 = ~v_1836 | v_71;
assign x_909 = ~v_1837 | v_100;
assign x_910 = ~v_1837 | v_78;
assign x_911 = ~v_1838 | v_100;
assign x_912 = ~v_1838 | v_84;
assign x_913 = ~v_1839 | v_100;
assign x_914 = ~v_1839 | v_89;
assign x_915 = ~v_1840 | v_100;
assign x_916 = ~v_1840 | v_93;
assign x_917 = ~v_1841 | v_100;
assign x_918 = ~v_1841 | v_96;
assign x_919 = ~v_1842 | v_100;
assign x_920 = ~v_1842 | v_98;
assign x_921 = ~v_1843 | v_321;
assign x_922 = ~v_1843 | ~v_322;
assign x_923 = ~v_1844 | v_63;
assign x_924 = ~v_1844 | ~v_322;
assign x_925 = ~v_1845 | v_321;
assign x_926 = ~v_1845 | v_63;
assign x_927 = ~v_1846 | v_320;
assign x_928 = ~v_1846 | ~v_321;
assign x_929 = ~v_1847 | v_71;
assign x_930 = ~v_1847 | ~v_321;
assign x_931 = ~v_1848 | v_320;
assign x_932 = ~v_1848 | v_71;
assign x_933 = ~v_1849 | v_319;
assign x_934 = ~v_1849 | ~v_320;
assign x_935 = ~v_1850 | v_78;
assign x_936 = ~v_1850 | ~v_320;
assign x_937 = ~v_1851 | v_319;
assign x_938 = ~v_1851 | v_78;
assign x_939 = ~v_1852 | v_318;
assign x_940 = ~v_1852 | ~v_319;
assign x_941 = ~v_1853 | v_84;
assign x_942 = ~v_1853 | ~v_319;
assign x_943 = ~v_1854 | v_318;
assign x_944 = ~v_1854 | v_84;
assign x_945 = ~v_1855 | v_317;
assign x_946 = ~v_1855 | ~v_318;
assign x_947 = ~v_1856 | v_89;
assign x_948 = ~v_1856 | ~v_318;
assign x_949 = ~v_1857 | v_317;
assign x_950 = ~v_1857 | v_89;
assign x_951 = ~v_1858 | v_316;
assign x_952 = ~v_1858 | ~v_317;
assign x_953 = ~v_1859 | v_93;
assign x_954 = ~v_1859 | ~v_317;
assign x_955 = ~v_1860 | v_316;
assign x_956 = ~v_1860 | v_93;
assign x_957 = ~v_1861 | v_98;
assign x_958 = ~v_1861 | ~v_316;
assign x_959 = ~v_1862 | v_96;
assign x_960 = ~v_1862 | ~v_316;
assign x_961 = ~v_1863 | v_98;
assign x_962 = ~v_1863 | v_96;
assign x_963 = ~v_1864 | v_314;
assign x_964 = ~v_1864 | ~v_315;
assign x_965 = ~v_1865 | v_64;
assign x_966 = ~v_1865 | ~v_315;
assign x_967 = ~v_1866 | v_314;
assign x_968 = ~v_1866 | v_64;
assign x_969 = ~v_1867 | v_313;
assign x_970 = ~v_1867 | ~v_314;
assign x_971 = ~v_1868 | v_72;
assign x_972 = ~v_1868 | ~v_314;
assign x_973 = ~v_1869 | v_313;
assign x_974 = ~v_1869 | v_72;
assign x_975 = ~v_1870 | v_312;
assign x_976 = ~v_1870 | ~v_313;
assign x_977 = ~v_1871 | v_79;
assign x_978 = ~v_1871 | ~v_313;
assign x_979 = ~v_1872 | v_312;
assign x_980 = ~v_1872 | v_79;
assign x_981 = ~v_1873 | v_311;
assign x_982 = ~v_1873 | ~v_312;
assign x_983 = ~v_1874 | v_85;
assign x_984 = ~v_1874 | ~v_312;
assign x_985 = ~v_1875 | v_311;
assign x_986 = ~v_1875 | v_85;
assign x_987 = ~v_1876 | v_310;
assign x_988 = ~v_1876 | ~v_311;
assign x_989 = ~v_1877 | v_90;
assign x_990 = ~v_1877 | ~v_311;
assign x_991 = ~v_1878 | v_310;
assign x_992 = ~v_1878 | v_90;
assign x_993 = ~v_1879 | v_309;
assign x_994 = ~v_1879 | ~v_310;
assign x_995 = ~v_1880 | v_94;
assign x_996 = ~v_1880 | ~v_310;
assign x_997 = ~v_1881 | v_309;
assign x_998 = ~v_1881 | v_94;
assign x_999 = ~v_1882 | v_308;
assign x_1000 = ~v_1882 | ~v_309;
assign x_1001 = ~v_1883 | v_97;
assign x_1002 = ~v_1883 | ~v_309;
assign x_1003 = ~v_1884 | v_308;
assign x_1004 = ~v_1884 | v_97;
assign x_1005 = ~v_1885 | v_100;
assign x_1006 = ~v_1885 | ~v_308;
assign x_1007 = ~v_1886 | v_99;
assign x_1008 = ~v_1886 | ~v_308;
assign x_1009 = ~v_1887 | v_100;
assign x_1010 = ~v_1887 | v_99;
assign x_1011 = ~v_1888 | v_3470;
assign x_1012 = ~v_1888 | ~v_3471;
assign x_1013 = ~v_1889 | v_109;
assign x_1014 = ~v_1889 | ~v_3471;
assign x_1015 = ~v_1890 | v_3470;
assign x_1016 = ~v_1890 | v_109;
assign x_1017 = ~v_1891 | v_3469;
assign x_1018 = ~v_1891 | ~v_3470;
assign x_1019 = ~v_1892 | v_108;
assign x_1020 = ~v_1892 | ~v_3470;
assign x_1021 = ~v_1893 | v_3469;
assign x_1022 = ~v_1893 | v_108;
assign x_1023 = ~v_1894 | v_3468;
assign x_1024 = ~v_1894 | ~v_3469;
assign x_1025 = ~v_1895 | v_107;
assign x_1026 = ~v_1895 | ~v_3469;
assign x_1027 = ~v_1896 | v_3468;
assign x_1028 = ~v_1896 | v_107;
assign x_1029 = ~v_1897 | v_3467;
assign x_1030 = ~v_1897 | ~v_3468;
assign x_1031 = ~v_1898 | v_106;
assign x_1032 = ~v_1898 | ~v_3468;
assign x_1033 = ~v_1899 | v_3467;
assign x_1034 = ~v_1899 | v_106;
assign x_1035 = ~v_1900 | v_3466;
assign x_1036 = ~v_1900 | ~v_3467;
assign x_1037 = ~v_1901 | v_105;
assign x_1038 = ~v_1901 | ~v_3467;
assign x_1039 = ~v_1902 | v_3466;
assign x_1040 = ~v_1902 | v_105;
assign x_1041 = ~v_1903 | v_3465;
assign x_1042 = ~v_1903 | ~v_3466;
assign x_1043 = ~v_1904 | v_104;
assign x_1044 = ~v_1904 | ~v_3466;
assign x_1045 = ~v_1905 | v_3465;
assign x_1046 = ~v_1905 | v_104;
assign x_1047 = ~v_1906 | v_3464;
assign x_1048 = ~v_1906 | ~v_3465;
assign x_1049 = ~v_1907 | v_103;
assign x_1050 = ~v_1907 | ~v_3465;
assign x_1051 = ~v_1908 | v_3464;
assign x_1052 = ~v_1908 | v_103;
assign x_1053 = ~v_1909 | v_101;
assign x_1054 = ~v_1909 | ~v_3464;
assign x_1055 = ~v_1910 | v_102;
assign x_1056 = ~v_1910 | ~v_3464;
assign x_1057 = ~v_1911 | v_101;
assign x_1058 = ~v_1911 | v_102;
assign x_1059 = ~v_1912 | v_3462;
assign x_1060 = ~v_1912 | ~v_3463;
assign x_1061 = ~v_1913 | v_117;
assign x_1062 = ~v_1913 | ~v_3463;
assign x_1063 = ~v_1914 | v_3462;
assign x_1064 = ~v_1914 | v_117;
assign x_1065 = ~v_1915 | v_3461;
assign x_1066 = ~v_1915 | ~v_3462;
assign x_1067 = ~v_1916 | v_116;
assign x_1068 = ~v_1916 | ~v_3462;
assign x_1069 = ~v_1917 | v_3461;
assign x_1070 = ~v_1917 | v_116;
assign x_1071 = ~v_1918 | v_3460;
assign x_1072 = ~v_1918 | ~v_3461;
assign x_1073 = ~v_1919 | v_115;
assign x_1074 = ~v_1919 | ~v_3461;
assign x_1075 = ~v_1920 | v_3460;
assign x_1076 = ~v_1920 | v_115;
assign x_1077 = ~v_1921 | v_3459;
assign x_1078 = ~v_1921 | ~v_3460;
assign x_1079 = ~v_1922 | v_114;
assign x_1080 = ~v_1922 | ~v_3460;
assign x_1081 = ~v_1923 | v_3459;
assign x_1082 = ~v_1923 | v_114;
assign x_1083 = ~v_1924 | v_3458;
assign x_1084 = ~v_1924 | ~v_3459;
assign x_1085 = ~v_1925 | v_113;
assign x_1086 = ~v_1925 | ~v_3459;
assign x_1087 = ~v_1926 | v_3458;
assign x_1088 = ~v_1926 | v_113;
assign x_1089 = ~v_1927 | v_3457;
assign x_1090 = ~v_1927 | ~v_3458;
assign x_1091 = ~v_1928 | v_112;
assign x_1092 = ~v_1928 | ~v_3458;
assign x_1093 = ~v_1929 | v_3457;
assign x_1094 = ~v_1929 | v_112;
assign x_1095 = ~v_1930 | v_110;
assign x_1096 = ~v_1930 | ~v_3457;
assign x_1097 = ~v_1931 | v_111;
assign x_1098 = ~v_1931 | ~v_3457;
assign x_1099 = ~v_1932 | v_110;
assign x_1100 = ~v_1932 | v_111;
assign x_1101 = ~v_1933 | v_101;
assign x_1102 = ~v_1933 | v_117;
assign x_1103 = ~v_1934 | v_101;
assign x_1104 = ~v_1934 | v_116;
assign x_1105 = ~v_1935 | v_101;
assign x_1106 = ~v_1935 | v_115;
assign x_1107 = ~v_1936 | v_101;
assign x_1108 = ~v_1936 | v_114;
assign x_1109 = ~v_1937 | v_101;
assign x_1110 = ~v_1937 | v_113;
assign x_1111 = ~v_1938 | v_101;
assign x_1112 = ~v_1938 | v_112;
assign x_1113 = ~v_1939 | v_101;
assign x_1114 = ~v_1939 | v_111;
assign x_1115 = ~v_1940 | v_101;
assign x_1116 = ~v_1940 | v_110;
assign x_1117 = ~v_1941 | v_3455;
assign x_1118 = ~v_1941 | ~v_3456;
assign x_1119 = ~v_1942 | v_124;
assign x_1120 = ~v_1942 | ~v_3456;
assign x_1121 = ~v_1943 | v_3455;
assign x_1122 = ~v_1943 | v_124;
assign x_1123 = ~v_1944 | v_3454;
assign x_1124 = ~v_1944 | ~v_3455;
assign x_1125 = ~v_1945 | v_123;
assign x_1126 = ~v_1945 | ~v_3455;
assign x_1127 = ~v_1946 | v_3454;
assign x_1128 = ~v_1946 | v_123;
assign x_1129 = ~v_1947 | v_3453;
assign x_1130 = ~v_1947 | ~v_3454;
assign x_1131 = ~v_1948 | v_122;
assign x_1132 = ~v_1948 | ~v_3454;
assign x_1133 = ~v_1949 | v_3453;
assign x_1134 = ~v_1949 | v_122;
assign x_1135 = ~v_1950 | v_3452;
assign x_1136 = ~v_1950 | ~v_3453;
assign x_1137 = ~v_1951 | v_121;
assign x_1138 = ~v_1951 | ~v_3453;
assign x_1139 = ~v_1952 | v_3452;
assign x_1140 = ~v_1952 | v_121;
assign x_1141 = ~v_1953 | v_3451;
assign x_1142 = ~v_1953 | ~v_3452;
assign x_1143 = ~v_1954 | v_120;
assign x_1144 = ~v_1954 | ~v_3452;
assign x_1145 = ~v_1955 | v_3451;
assign x_1146 = ~v_1955 | v_120;
assign x_1147 = ~v_1956 | v_118;
assign x_1148 = ~v_1956 | ~v_3451;
assign x_1149 = ~v_1957 | v_119;
assign x_1150 = ~v_1957 | ~v_3451;
assign x_1151 = ~v_1958 | v_118;
assign x_1152 = ~v_1958 | v_119;
assign x_1153 = ~v_1959 | v_3450;
assign x_1154 = ~v_1959 | v_124;
assign x_1155 = ~v_1960 | v_3450;
assign x_1156 = ~v_1960 | v_123;
assign x_1157 = ~v_1961 | v_3450;
assign x_1158 = ~v_1961 | v_122;
assign x_1159 = ~v_1962 | v_3450;
assign x_1160 = ~v_1962 | v_121;
assign x_1161 = ~v_1963 | v_3450;
assign x_1162 = ~v_1963 | v_120;
assign x_1163 = ~v_1964 | v_3450;
assign x_1164 = ~v_1964 | v_119;
assign x_1165 = ~v_1965 | v_3450;
assign x_1166 = ~v_1965 | v_118;
assign x_1167 = ~v_1966 | v_102;
assign x_1168 = ~v_1966 | ~v_3450;
assign x_1169 = ~v_1967 | v_110;
assign x_1170 = ~v_1967 | ~v_3450;
assign x_1171 = ~v_1968 | v_102;
assign x_1172 = ~v_1968 | v_110;
assign x_1173 = ~v_1969 | v_3448;
assign x_1174 = ~v_1969 | ~v_3449;
assign x_1175 = ~v_1970 | v_130;
assign x_1176 = ~v_1970 | ~v_3449;
assign x_1177 = ~v_1971 | v_3448;
assign x_1178 = ~v_1971 | v_130;
assign x_1179 = ~v_1972 | v_3447;
assign x_1180 = ~v_1972 | ~v_3448;
assign x_1181 = ~v_1973 | v_129;
assign x_1182 = ~v_1973 | ~v_3448;
assign x_1183 = ~v_1974 | v_3447;
assign x_1184 = ~v_1974 | v_129;
assign x_1185 = ~v_1975 | v_3446;
assign x_1186 = ~v_1975 | ~v_3447;
assign x_1187 = ~v_1976 | v_128;
assign x_1188 = ~v_1976 | ~v_3447;
assign x_1189 = ~v_1977 | v_3446;
assign x_1190 = ~v_1977 | v_128;
assign x_1191 = ~v_1978 | v_3445;
assign x_1192 = ~v_1978 | ~v_3446;
assign x_1193 = ~v_1979 | v_127;
assign x_1194 = ~v_1979 | ~v_3446;
assign x_1195 = ~v_1980 | v_3445;
assign x_1196 = ~v_1980 | v_127;
assign x_1197 = ~v_1981 | v_125;
assign x_1198 = ~v_1981 | ~v_3445;
assign x_1199 = ~v_1982 | v_126;
assign x_1200 = ~v_1982 | ~v_3445;
assign x_1201 = ~v_1983 | v_125;
assign x_1202 = ~v_1983 | v_126;
assign x_1203 = ~v_1984 | v_3444;
assign x_1204 = ~v_1984 | v_130;
assign x_1205 = ~v_1985 | v_3444;
assign x_1206 = ~v_1985 | v_129;
assign x_1207 = ~v_1986 | v_3444;
assign x_1208 = ~v_1986 | v_128;
assign x_1209 = ~v_1987 | v_3444;
assign x_1210 = ~v_1987 | v_127;
assign x_1211 = ~v_1988 | v_3444;
assign x_1212 = ~v_1988 | v_126;
assign x_1213 = ~v_1989 | v_3444;
assign x_1214 = ~v_1989 | v_125;
assign x_1215 = ~v_1990 | v_3443;
assign x_1216 = ~v_1990 | ~v_3444;
assign x_1217 = ~v_1991 | v_118;
assign x_1218 = ~v_1991 | ~v_3444;
assign x_1219 = ~v_1992 | v_3443;
assign x_1220 = ~v_1992 | v_118;
assign x_1221 = ~v_1993 | v_103;
assign x_1222 = ~v_1993 | ~v_3443;
assign x_1223 = ~v_1994 | v_111;
assign x_1224 = ~v_1994 | ~v_3443;
assign x_1225 = ~v_1995 | v_103;
assign x_1226 = ~v_1995 | v_111;
assign x_1227 = ~v_1996 | v_3441;
assign x_1228 = ~v_1996 | ~v_3442;
assign x_1229 = ~v_1997 | v_135;
assign x_1230 = ~v_1997 | ~v_3442;
assign x_1231 = ~v_1998 | v_3441;
assign x_1232 = ~v_1998 | v_135;
assign x_1233 = ~v_1999 | v_3440;
assign x_1234 = ~v_1999 | ~v_3441;
assign x_1235 = ~v_2000 | v_134;
assign x_1236 = ~v_2000 | ~v_3441;
assign x_1237 = ~v_2001 | v_3440;
assign x_1238 = ~v_2001 | v_134;
assign x_1239 = ~v_2002 | v_3439;
assign x_1240 = ~v_2002 | ~v_3440;
assign x_1241 = ~v_2003 | v_133;
assign x_1242 = ~v_2003 | ~v_3440;
assign x_1243 = ~v_2004 | v_3439;
assign x_1244 = ~v_2004 | v_133;
assign x_1245 = ~v_2005 | v_131;
assign x_1246 = ~v_2005 | ~v_3439;
assign x_1247 = ~v_2006 | v_132;
assign x_1248 = ~v_2006 | ~v_3439;
assign x_1249 = ~v_2007 | v_131;
assign x_1250 = ~v_2007 | v_132;
assign x_1251 = ~v_2008 | v_3438;
assign x_1252 = ~v_2008 | v_135;
assign x_1253 = ~v_2009 | v_3438;
assign x_1254 = ~v_2009 | v_134;
assign x_1255 = ~v_2010 | v_3438;
assign x_1256 = ~v_2010 | v_133;
assign x_1257 = ~v_2011 | v_3438;
assign x_1258 = ~v_2011 | v_132;
assign x_1259 = ~v_2012 | v_3438;
assign x_1260 = ~v_2012 | v_131;
assign x_1261 = ~v_2013 | v_3437;
assign x_1262 = ~v_2013 | ~v_3438;
assign x_1263 = ~v_2014 | v_125;
assign x_1264 = ~v_2014 | ~v_3438;
assign x_1265 = ~v_2015 | v_3437;
assign x_1266 = ~v_2015 | v_125;
assign x_1267 = ~v_2016 | v_3436;
assign x_1268 = ~v_2016 | ~v_3437;
assign x_1269 = ~v_2017 | v_119;
assign x_1270 = ~v_2017 | ~v_3437;
assign x_1271 = ~v_2018 | v_3436;
assign x_1272 = ~v_2018 | v_119;
assign x_1273 = ~v_2019 | v_104;
assign x_1274 = ~v_2019 | ~v_3436;
assign x_1275 = ~v_2020 | v_112;
assign x_1276 = ~v_2020 | ~v_3436;
assign x_1277 = ~v_2021 | v_104;
assign x_1278 = ~v_2021 | v_112;
assign x_1279 = ~v_2022 | v_3434;
assign x_1280 = ~v_2022 | ~v_3435;
assign x_1281 = ~v_2023 | v_139;
assign x_1282 = ~v_2023 | ~v_3435;
assign x_1283 = ~v_2024 | v_3434;
assign x_1284 = ~v_2024 | v_139;
assign x_1285 = ~v_2025 | v_3433;
assign x_1286 = ~v_2025 | ~v_3434;
assign x_1287 = ~v_2026 | v_138;
assign x_1288 = ~v_2026 | ~v_3434;
assign x_1289 = ~v_2027 | v_3433;
assign x_1290 = ~v_2027 | v_138;
assign x_1291 = ~v_2028 | v_136;
assign x_1292 = ~v_2028 | ~v_3433;
assign x_1293 = ~v_2029 | v_137;
assign x_1294 = ~v_2029 | ~v_3433;
assign x_1295 = ~v_2030 | v_136;
assign x_1296 = ~v_2030 | v_137;
assign x_1297 = ~v_2031 | v_3432;
assign x_1298 = ~v_2031 | v_139;
assign x_1299 = ~v_2032 | v_3432;
assign x_1300 = ~v_2032 | v_138;
assign x_1301 = ~v_2033 | v_3432;
assign x_1302 = ~v_2033 | v_137;
assign x_1303 = ~v_2034 | v_3432;
assign x_1304 = ~v_2034 | v_136;
assign x_1305 = ~v_2035 | v_3431;
assign x_1306 = ~v_2035 | ~v_3432;
assign x_1307 = ~v_2036 | v_131;
assign x_1308 = ~v_2036 | ~v_3432;
assign x_1309 = ~v_2037 | v_3431;
assign x_1310 = ~v_2037 | v_131;
assign x_1311 = ~v_2038 | v_3430;
assign x_1312 = ~v_2038 | ~v_3431;
assign x_1313 = ~v_2039 | v_126;
assign x_1314 = ~v_2039 | ~v_3431;
assign x_1315 = ~v_2040 | v_3430;
assign x_1316 = ~v_2040 | v_126;
assign x_1317 = ~v_2041 | v_3429;
assign x_1318 = ~v_2041 | ~v_3430;
assign x_1319 = ~v_2042 | v_120;
assign x_1320 = ~v_2042 | ~v_3430;
assign x_1321 = ~v_2043 | v_3429;
assign x_1322 = ~v_2043 | v_120;
assign x_1323 = ~v_2044 | v_105;
assign x_1324 = ~v_2044 | ~v_3429;
assign x_1325 = ~v_2045 | v_113;
assign x_1326 = ~v_2045 | ~v_3429;
assign x_1327 = ~v_2046 | v_105;
assign x_1328 = ~v_2046 | v_113;
assign x_1329 = ~v_2047 | v_3427;
assign x_1330 = ~v_2047 | ~v_3428;
assign x_1331 = ~v_2048 | v_142;
assign x_1332 = ~v_2048 | ~v_3428;
assign x_1333 = ~v_2049 | v_3427;
assign x_1334 = ~v_2049 | v_142;
assign x_1335 = ~v_2050 | v_140;
assign x_1336 = ~v_2050 | ~v_3427;
assign x_1337 = ~v_2051 | v_141;
assign x_1338 = ~v_2051 | ~v_3427;
assign x_1339 = ~v_2052 | v_140;
assign x_1340 = ~v_2052 | v_141;
assign x_1341 = ~v_2053 | v_3426;
assign x_1342 = ~v_2053 | v_142;
assign x_1343 = ~v_2054 | v_3426;
assign x_1344 = ~v_2054 | v_141;
assign x_1345 = ~v_2055 | v_3426;
assign x_1346 = ~v_2055 | v_140;
assign x_1347 = ~v_2056 | v_3425;
assign x_1348 = ~v_2056 | ~v_3426;
assign x_1349 = ~v_2057 | v_136;
assign x_1350 = ~v_2057 | ~v_3426;
assign x_1351 = ~v_2058 | v_3425;
assign x_1352 = ~v_2058 | v_136;
assign x_1353 = ~v_2059 | v_3424;
assign x_1354 = ~v_2059 | ~v_3425;
assign x_1355 = ~v_2060 | v_132;
assign x_1356 = ~v_2060 | ~v_3425;
assign x_1357 = ~v_2061 | v_3424;
assign x_1358 = ~v_2061 | v_132;
assign x_1359 = ~v_2062 | v_3423;
assign x_1360 = ~v_2062 | ~v_3424;
assign x_1361 = ~v_2063 | v_127;
assign x_1362 = ~v_2063 | ~v_3424;
assign x_1363 = ~v_2064 | v_3423;
assign x_1364 = ~v_2064 | v_127;
assign x_1365 = ~v_2065 | v_3422;
assign x_1366 = ~v_2065 | ~v_3423;
assign x_1367 = ~v_2066 | v_121;
assign x_1368 = ~v_2066 | ~v_3423;
assign x_1369 = ~v_2067 | v_3422;
assign x_1370 = ~v_2067 | v_121;
assign x_1371 = ~v_2068 | v_106;
assign x_1372 = ~v_2068 | ~v_3422;
assign x_1373 = ~v_2069 | v_114;
assign x_1374 = ~v_2069 | ~v_3422;
assign x_1375 = ~v_2070 | v_106;
assign x_1376 = ~v_2070 | v_114;
assign x_1377 = ~v_2071 | v_143;
assign x_1378 = ~v_2071 | ~v_3421;
assign x_1379 = ~v_2072 | v_144;
assign x_1380 = ~v_2072 | ~v_3421;
assign x_1381 = ~v_2073 | v_143;
assign x_1382 = ~v_2073 | v_144;
assign x_1383 = ~v_2074 | v_3420;
assign x_1384 = ~v_2074 | v_144;
assign x_1385 = ~v_2075 | v_3420;
assign x_1386 = ~v_2075 | v_143;
assign x_1387 = ~v_2076 | v_3419;
assign x_1388 = ~v_2076 | ~v_3420;
assign x_1389 = ~v_2077 | v_140;
assign x_1390 = ~v_2077 | ~v_3420;
assign x_1391 = ~v_2078 | v_3419;
assign x_1392 = ~v_2078 | v_140;
assign x_1393 = ~v_2079 | v_3418;
assign x_1394 = ~v_2079 | ~v_3419;
assign x_1395 = ~v_2080 | v_137;
assign x_1396 = ~v_2080 | ~v_3419;
assign x_1397 = ~v_2081 | v_3418;
assign x_1398 = ~v_2081 | v_137;
assign x_1399 = ~v_2082 | v_3417;
assign x_1400 = ~v_2082 | ~v_3418;
assign x_1401 = ~v_2083 | v_133;
assign x_1402 = ~v_2083 | ~v_3418;
assign x_1403 = ~v_2084 | v_3417;
assign x_1404 = ~v_2084 | v_133;
assign x_1405 = ~v_2085 | v_3416;
assign x_1406 = ~v_2085 | ~v_3417;
assign x_1407 = ~v_2086 | v_128;
assign x_1408 = ~v_2086 | ~v_3417;
assign x_1409 = ~v_2087 | v_3416;
assign x_1410 = ~v_2087 | v_128;
assign x_1411 = ~v_2088 | v_3415;
assign x_1412 = ~v_2088 | ~v_3416;
assign x_1413 = ~v_2089 | v_122;
assign x_1414 = ~v_2089 | ~v_3416;
assign x_1415 = ~v_2090 | v_3415;
assign x_1416 = ~v_2090 | v_122;
assign x_1417 = ~v_2091 | v_107;
assign x_1418 = ~v_2091 | ~v_3415;
assign x_1419 = ~v_2092 | v_115;
assign x_1420 = ~v_2092 | ~v_3415;
assign x_1421 = ~v_2093 | v_107;
assign x_1422 = ~v_2093 | v_115;
assign x_1423 = ~v_2094 | v_3414;
assign x_1424 = ~v_2094 | v_145;
assign x_1425 = ~v_2095 | v_3413;
assign x_1426 = ~v_2095 | ~v_3414;
assign x_1427 = ~v_2096 | v_143;
assign x_1428 = ~v_2096 | ~v_3414;
assign x_1429 = ~v_2097 | v_3413;
assign x_1430 = ~v_2097 | v_143;
assign x_1431 = ~v_2098 | v_3412;
assign x_1432 = ~v_2098 | ~v_3413;
assign x_1433 = ~v_2099 | v_141;
assign x_1434 = ~v_2099 | ~v_3413;
assign x_1435 = ~v_2100 | v_3412;
assign x_1436 = ~v_2100 | v_141;
assign x_1437 = ~v_2101 | v_3411;
assign x_1438 = ~v_2101 | ~v_3412;
assign x_1439 = ~v_2102 | v_138;
assign x_1440 = ~v_2102 | ~v_3412;
assign x_1441 = ~v_2103 | v_3411;
assign x_1442 = ~v_2103 | v_138;
assign x_1443 = ~v_2104 | v_3410;
assign x_1444 = ~v_2104 | ~v_3411;
assign x_1445 = ~v_2105 | v_134;
assign x_1446 = ~v_2105 | ~v_3411;
assign x_1447 = ~v_2106 | v_3410;
assign x_1448 = ~v_2106 | v_134;
assign x_1449 = ~v_2107 | v_3409;
assign x_1450 = ~v_2107 | ~v_3410;
assign x_1451 = ~v_2108 | v_129;
assign x_1452 = ~v_2108 | ~v_3410;
assign x_1453 = ~v_2109 | v_3409;
assign x_1454 = ~v_2109 | v_129;
assign x_1455 = ~v_2110 | v_3408;
assign x_1456 = ~v_2110 | ~v_3409;
assign x_1457 = ~v_2111 | v_123;
assign x_1458 = ~v_2111 | ~v_3409;
assign x_1459 = ~v_2112 | v_3408;
assign x_1460 = ~v_2112 | v_123;
assign x_1461 = ~v_2113 | v_108;
assign x_1462 = ~v_2113 | ~v_3408;
assign x_1463 = ~v_2114 | v_116;
assign x_1464 = ~v_2114 | ~v_3408;
assign x_1465 = ~v_2115 | v_108;
assign x_1466 = ~v_2115 | v_116;
assign x_1467 = ~v_2116 | v_3406;
assign x_1468 = ~v_2116 | ~v_3407;
assign x_1469 = ~v_2117 | v_145;
assign x_1470 = ~v_2117 | ~v_3407;
assign x_1471 = ~v_2118 | v_3406;
assign x_1472 = ~v_2118 | v_145;
assign x_1473 = ~v_2119 | v_3405;
assign x_1474 = ~v_2119 | ~v_3406;
assign x_1475 = ~v_2120 | v_144;
assign x_1476 = ~v_2120 | ~v_3406;
assign x_1477 = ~v_2121 | v_3405;
assign x_1478 = ~v_2121 | v_144;
assign x_1479 = ~v_2122 | v_3404;
assign x_1480 = ~v_2122 | ~v_3405;
assign x_1481 = ~v_2123 | v_142;
assign x_1482 = ~v_2123 | ~v_3405;
assign x_1483 = ~v_2124 | v_3404;
assign x_1484 = ~v_2124 | v_142;
assign x_1485 = ~v_2125 | v_3403;
assign x_1486 = ~v_2125 | ~v_3404;
assign x_1487 = ~v_2126 | v_139;
assign x_1488 = ~v_2126 | ~v_3404;
assign x_1489 = ~v_2127 | v_3403;
assign x_1490 = ~v_2127 | v_139;
assign x_1491 = ~v_2128 | v_3402;
assign x_1492 = ~v_2128 | ~v_3403;
assign x_1493 = ~v_2129 | v_135;
assign x_1494 = ~v_2129 | ~v_3403;
assign x_1495 = ~v_2130 | v_3402;
assign x_1496 = ~v_2130 | v_135;
assign x_1497 = ~v_2131 | v_3401;
assign x_1498 = ~v_2131 | ~v_3402;
assign x_1499 = ~v_2132 | v_130;
assign x_1500 = ~v_2132 | ~v_3402;
assign x_1501 = ~v_2133 | v_3401;
assign x_1502 = ~v_2133 | v_130;
assign x_1503 = ~v_2134 | v_3400;
assign x_1504 = ~v_2134 | ~v_3401;
assign x_1505 = ~v_2135 | v_124;
assign x_1506 = ~v_2135 | ~v_3401;
assign x_1507 = ~v_2136 | v_3400;
assign x_1508 = ~v_2136 | v_124;
assign x_1509 = ~v_2137 | v_109;
assign x_1510 = ~v_2137 | ~v_3400;
assign x_1511 = ~v_2138 | v_117;
assign x_1512 = ~v_2138 | ~v_3400;
assign x_1513 = ~v_2139 | v_109;
assign x_1514 = ~v_2139 | v_117;
assign x_1515 = ~v_2140 | v_3542;
assign x_1516 = ~v_2140 | ~v_3543;
assign x_1517 = ~v_2141 | v_101;
assign x_1518 = ~v_2141 | ~v_3543;
assign x_1519 = ~v_2142 | v_3542;
assign x_1520 = ~v_2142 | v_101;
assign x_1521 = ~v_2143 | v_3541;
assign x_1522 = ~v_2143 | ~v_3542;
assign x_1523 = ~v_2144 | v_102;
assign x_1524 = ~v_2144 | ~v_3542;
assign x_1525 = ~v_2145 | v_3541;
assign x_1526 = ~v_2145 | v_102;
assign x_1527 = ~v_2146 | v_3540;
assign x_1528 = ~v_2146 | ~v_3541;
assign x_1529 = ~v_2147 | v_103;
assign x_1530 = ~v_2147 | ~v_3541;
assign x_1531 = ~v_2148 | v_3540;
assign x_1532 = ~v_2148 | v_103;
assign x_1533 = ~v_2149 | v_3539;
assign x_1534 = ~v_2149 | ~v_3540;
assign x_1535 = ~v_2150 | v_104;
assign x_1536 = ~v_2150 | ~v_3540;
assign x_1537 = ~v_2151 | v_3539;
assign x_1538 = ~v_2151 | v_104;
assign x_1539 = ~v_2152 | v_3538;
assign x_1540 = ~v_2152 | ~v_3539;
assign x_1541 = ~v_2153 | v_105;
assign x_1542 = ~v_2153 | ~v_3539;
assign x_1543 = ~v_2154 | v_3538;
assign x_1544 = ~v_2154 | v_105;
assign x_1545 = ~v_2155 | v_3537;
assign x_1546 = ~v_2155 | ~v_3538;
assign x_1547 = ~v_2156 | v_106;
assign x_1548 = ~v_2156 | ~v_3538;
assign x_1549 = ~v_2157 | v_3537;
assign x_1550 = ~v_2157 | v_106;
assign x_1551 = ~v_2158 | v_3536;
assign x_1552 = ~v_2158 | ~v_3537;
assign x_1553 = ~v_2159 | v_107;
assign x_1554 = ~v_2159 | ~v_3537;
assign x_1555 = ~v_2160 | v_3536;
assign x_1556 = ~v_2160 | v_107;
assign x_1557 = ~v_2161 | v_109;
assign x_1558 = ~v_2161 | ~v_3536;
assign x_1559 = ~v_2162 | v_108;
assign x_1560 = ~v_2162 | ~v_3536;
assign x_1561 = ~v_2163 | v_109;
assign x_1562 = ~v_2163 | v_108;
assign x_1563 = ~v_2164 | v_3535;
assign x_1564 = ~v_2164 | v_101;
assign x_1565 = ~v_2165 | v_3534;
assign x_1566 = ~v_2165 | ~v_3535;
assign x_1567 = ~v_2166 | v_110;
assign x_1568 = ~v_2166 | ~v_3535;
assign x_1569 = ~v_2167 | v_3534;
assign x_1570 = ~v_2167 | v_110;
assign x_1571 = ~v_2168 | v_3533;
assign x_1572 = ~v_2168 | ~v_3534;
assign x_1573 = ~v_2169 | v_111;
assign x_1574 = ~v_2169 | ~v_3534;
assign x_1575 = ~v_2170 | v_3533;
assign x_1576 = ~v_2170 | v_111;
assign x_1577 = ~v_2171 | v_3532;
assign x_1578 = ~v_2171 | ~v_3533;
assign x_1579 = ~v_2172 | v_112;
assign x_1580 = ~v_2172 | ~v_3533;
assign x_1581 = ~v_2173 | v_3532;
assign x_1582 = ~v_2173 | v_112;
assign x_1583 = ~v_2174 | v_3531;
assign x_1584 = ~v_2174 | ~v_3532;
assign x_1585 = ~v_2175 | v_113;
assign x_1586 = ~v_2175 | ~v_3532;
assign x_1587 = ~v_2176 | v_3531;
assign x_1588 = ~v_2176 | v_113;
assign x_1589 = ~v_2177 | v_3530;
assign x_1590 = ~v_2177 | ~v_3531;
assign x_1591 = ~v_2178 | v_114;
assign x_1592 = ~v_2178 | ~v_3531;
assign x_1593 = ~v_2179 | v_3530;
assign x_1594 = ~v_2179 | v_114;
assign x_1595 = ~v_2180 | v_3529;
assign x_1596 = ~v_2180 | ~v_3530;
assign x_1597 = ~v_2181 | v_115;
assign x_1598 = ~v_2181 | ~v_3530;
assign x_1599 = ~v_2182 | v_3529;
assign x_1600 = ~v_2182 | v_115;
assign x_1601 = ~v_2183 | v_117;
assign x_1602 = ~v_2183 | ~v_3529;
assign x_1603 = ~v_2184 | v_116;
assign x_1604 = ~v_2184 | ~v_3529;
assign x_1605 = ~v_2185 | v_117;
assign x_1606 = ~v_2185 | v_116;
assign x_1607 = ~v_2186 | v_3528;
assign x_1608 = ~v_2186 | v_102;
assign x_1609 = ~v_2187 | v_3528;
assign x_1610 = ~v_2187 | v_110;
assign x_1611 = ~v_2188 | v_3527;
assign x_1612 = ~v_2188 | ~v_3528;
assign x_1613 = ~v_2189 | v_118;
assign x_1614 = ~v_2189 | ~v_3528;
assign x_1615 = ~v_2190 | v_3527;
assign x_1616 = ~v_2190 | v_118;
assign x_1617 = ~v_2191 | v_3526;
assign x_1618 = ~v_2191 | ~v_3527;
assign x_1619 = ~v_2192 | v_119;
assign x_1620 = ~v_2192 | ~v_3527;
assign x_1621 = ~v_2193 | v_3526;
assign x_1622 = ~v_2193 | v_119;
assign x_1623 = ~v_2194 | v_3525;
assign x_1624 = ~v_2194 | ~v_3526;
assign x_1625 = ~v_2195 | v_120;
assign x_1626 = ~v_2195 | ~v_3526;
assign x_1627 = ~v_2196 | v_3525;
assign x_1628 = ~v_2196 | v_120;
assign x_1629 = ~v_2197 | v_3524;
assign x_1630 = ~v_2197 | ~v_3525;
assign x_1631 = ~v_2198 | v_121;
assign x_1632 = ~v_2198 | ~v_3525;
assign x_1633 = ~v_2199 | v_3524;
assign x_1634 = ~v_2199 | v_121;
assign x_1635 = ~v_2200 | v_3523;
assign x_1636 = ~v_2200 | ~v_3524;
assign x_1637 = ~v_2201 | v_122;
assign x_1638 = ~v_2201 | ~v_3524;
assign x_1639 = ~v_2202 | v_3523;
assign x_1640 = ~v_2202 | v_122;
assign x_1641 = ~v_2203 | v_124;
assign x_1642 = ~v_2203 | ~v_3523;
assign x_1643 = ~v_2204 | v_123;
assign x_1644 = ~v_2204 | ~v_3523;
assign x_1645 = ~v_2205 | v_124;
assign x_1646 = ~v_2205 | v_123;
assign x_1647 = ~v_2206 | v_110;
assign x_1648 = ~v_2206 | ~v_3522;
assign x_1649 = ~v_2207 | v_102;
assign x_1650 = ~v_2207 | ~v_3522;
assign x_1651 = ~v_2208 | v_110;
assign x_1652 = ~v_2208 | v_102;
assign x_1653 = ~v_2209 | v_3521;
assign x_1654 = ~v_2209 | v_103;
assign x_1655 = ~v_2210 | v_3521;
assign x_1656 = ~v_2210 | v_111;
assign x_1657 = ~v_2211 | v_3521;
assign x_1658 = ~v_2211 | v_118;
assign x_1659 = ~v_2212 | v_3520;
assign x_1660 = ~v_2212 | ~v_3521;
assign x_1661 = ~v_2213 | v_125;
assign x_1662 = ~v_2213 | ~v_3521;
assign x_1663 = ~v_2214 | v_3520;
assign x_1664 = ~v_2214 | v_125;
assign x_1665 = ~v_2215 | v_3519;
assign x_1666 = ~v_2215 | ~v_3520;
assign x_1667 = ~v_2216 | v_126;
assign x_1668 = ~v_2216 | ~v_3520;
assign x_1669 = ~v_2217 | v_3519;
assign x_1670 = ~v_2217 | v_126;
assign x_1671 = ~v_2218 | v_3518;
assign x_1672 = ~v_2218 | ~v_3519;
assign x_1673 = ~v_2219 | v_127;
assign x_1674 = ~v_2219 | ~v_3519;
assign x_1675 = ~v_2220 | v_3518;
assign x_1676 = ~v_2220 | v_127;
assign x_1677 = ~v_2221 | v_3517;
assign x_1678 = ~v_2221 | ~v_3518;
assign x_1679 = ~v_2222 | v_128;
assign x_1680 = ~v_2222 | ~v_3518;
assign x_1681 = ~v_2223 | v_3517;
assign x_1682 = ~v_2223 | v_128;
assign x_1683 = ~v_2224 | v_130;
assign x_1684 = ~v_2224 | ~v_3517;
assign x_1685 = ~v_2225 | v_129;
assign x_1686 = ~v_2225 | ~v_3517;
assign x_1687 = ~v_2226 | v_130;
assign x_1688 = ~v_2226 | v_129;
assign x_1689 = ~v_2227 | v_3515;
assign x_1690 = ~v_2227 | ~v_3516;
assign x_1691 = ~v_2228 | v_103;
assign x_1692 = ~v_2228 | ~v_3516;
assign x_1693 = ~v_2229 | v_3515;
assign x_1694 = ~v_2229 | v_103;
assign x_1695 = ~v_2230 | v_118;
assign x_1696 = ~v_2230 | ~v_3515;
assign x_1697 = ~v_2231 | v_111;
assign x_1698 = ~v_2231 | ~v_3515;
assign x_1699 = ~v_2232 | v_118;
assign x_1700 = ~v_2232 | v_111;
assign x_1701 = ~v_2233 | v_3514;
assign x_1702 = ~v_2233 | v_104;
assign x_1703 = ~v_2234 | v_3514;
assign x_1704 = ~v_2234 | v_112;
assign x_1705 = ~v_2235 | v_3514;
assign x_1706 = ~v_2235 | v_119;
assign x_1707 = ~v_2236 | v_3514;
assign x_1708 = ~v_2236 | v_125;
assign x_1709 = ~v_2237 | v_3513;
assign x_1710 = ~v_2237 | ~v_3514;
assign x_1711 = ~v_2238 | v_131;
assign x_1712 = ~v_2238 | ~v_3514;
assign x_1713 = ~v_2239 | v_3513;
assign x_1714 = ~v_2239 | v_131;
assign x_1715 = ~v_2240 | v_3512;
assign x_1716 = ~v_2240 | ~v_3513;
assign x_1717 = ~v_2241 | v_132;
assign x_1718 = ~v_2241 | ~v_3513;
assign x_1719 = ~v_2242 | v_3512;
assign x_1720 = ~v_2242 | v_132;
assign x_1721 = ~v_2243 | v_3511;
assign x_1722 = ~v_2243 | ~v_3512;
assign x_1723 = ~v_2244 | v_133;
assign x_1724 = ~v_2244 | ~v_3512;
assign x_1725 = ~v_2245 | v_3511;
assign x_1726 = ~v_2245 | v_133;
assign x_1727 = ~v_2246 | v_135;
assign x_1728 = ~v_2246 | ~v_3511;
assign x_1729 = ~v_2247 | v_134;
assign x_1730 = ~v_2247 | ~v_3511;
assign x_1731 = ~v_2248 | v_135;
assign x_1732 = ~v_2248 | v_134;
assign x_1733 = ~v_2249 | v_3509;
assign x_1734 = ~v_2249 | ~v_3510;
assign x_1735 = ~v_2250 | v_104;
assign x_1736 = ~v_2250 | ~v_3510;
assign x_1737 = ~v_2251 | v_3509;
assign x_1738 = ~v_2251 | v_104;
assign x_1739 = ~v_2252 | v_3508;
assign x_1740 = ~v_2252 | ~v_3509;
assign x_1741 = ~v_2253 | v_112;
assign x_1742 = ~v_2253 | ~v_3509;
assign x_1743 = ~v_2254 | v_3508;
assign x_1744 = ~v_2254 | v_112;
assign x_1745 = ~v_2255 | v_125;
assign x_1746 = ~v_2255 | ~v_3508;
assign x_1747 = ~v_2256 | v_119;
assign x_1748 = ~v_2256 | ~v_3508;
assign x_1749 = ~v_2257 | v_125;
assign x_1750 = ~v_2257 | v_119;
assign x_1751 = ~v_2258 | v_3507;
assign x_1752 = ~v_2258 | v_105;
assign x_1753 = ~v_2259 | v_3507;
assign x_1754 = ~v_2259 | v_113;
assign x_1755 = ~v_2260 | v_3507;
assign x_1756 = ~v_2260 | v_120;
assign x_1757 = ~v_2261 | v_3507;
assign x_1758 = ~v_2261 | v_126;
assign x_1759 = ~v_2262 | v_3507;
assign x_1760 = ~v_2262 | v_131;
assign x_1761 = ~v_2263 | v_3506;
assign x_1762 = ~v_2263 | ~v_3507;
assign x_1763 = ~v_2264 | v_136;
assign x_1764 = ~v_2264 | ~v_3507;
assign x_1765 = ~v_2265 | v_3506;
assign x_1766 = ~v_2265 | v_136;
assign x_1767 = ~v_2266 | v_3505;
assign x_1768 = ~v_2266 | ~v_3506;
assign x_1769 = ~v_2267 | v_137;
assign x_1770 = ~v_2267 | ~v_3506;
assign x_1771 = ~v_2268 | v_3505;
assign x_1772 = ~v_2268 | v_137;
assign x_1773 = ~v_2269 | v_139;
assign x_1774 = ~v_2269 | ~v_3505;
assign x_1775 = ~v_2270 | v_138;
assign x_1776 = ~v_2270 | ~v_3505;
assign x_1777 = ~v_2271 | v_139;
assign x_1778 = ~v_2271 | v_138;
assign x_1779 = ~v_2272 | v_3503;
assign x_1780 = ~v_2272 | ~v_3504;
assign x_1781 = ~v_2273 | v_105;
assign x_1782 = ~v_2273 | ~v_3504;
assign x_1783 = ~v_2274 | v_3503;
assign x_1784 = ~v_2274 | v_105;
assign x_1785 = ~v_2275 | v_3502;
assign x_1786 = ~v_2275 | ~v_3503;
assign x_1787 = ~v_2276 | v_113;
assign x_1788 = ~v_2276 | ~v_3503;
assign x_1789 = ~v_2277 | v_3502;
assign x_1790 = ~v_2277 | v_113;
assign x_1791 = ~v_2278 | v_3501;
assign x_1792 = ~v_2278 | ~v_3502;
assign x_1793 = ~v_2279 | v_120;
assign x_1794 = ~v_2279 | ~v_3502;
assign x_1795 = ~v_2280 | v_3501;
assign x_1796 = ~v_2280 | v_120;
assign x_1797 = ~v_2281 | v_131;
assign x_1798 = ~v_2281 | ~v_3501;
assign x_1799 = ~v_2282 | v_126;
assign x_1800 = ~v_2282 | ~v_3501;
assign x_1801 = ~v_2283 | v_131;
assign x_1802 = ~v_2283 | v_126;
assign x_1803 = ~v_2284 | v_3500;
assign x_1804 = ~v_2284 | v_106;
assign x_1805 = ~v_2285 | v_3500;
assign x_1806 = ~v_2285 | v_114;
assign x_1807 = ~v_2286 | v_3500;
assign x_1808 = ~v_2286 | v_121;
assign x_1809 = ~v_2287 | v_3500;
assign x_1810 = ~v_2287 | v_127;
assign x_1811 = ~v_2288 | v_3500;
assign x_1812 = ~v_2288 | v_132;
assign x_1813 = ~v_2289 | v_3500;
assign x_1814 = ~v_2289 | v_136;
assign x_1815 = ~v_2290 | v_3499;
assign x_1816 = ~v_2290 | ~v_3500;
assign x_1817 = ~v_2291 | v_140;
assign x_1818 = ~v_2291 | ~v_3500;
assign x_1819 = ~v_2292 | v_3499;
assign x_1820 = ~v_2292 | v_140;
assign x_1821 = ~v_2293 | v_142;
assign x_1822 = ~v_2293 | ~v_3499;
assign x_1823 = ~v_2294 | v_141;
assign x_1824 = ~v_2294 | ~v_3499;
assign x_1825 = ~v_2295 | v_142;
assign x_1826 = ~v_2295 | v_141;
assign x_1827 = ~v_2296 | v_3497;
assign x_1828 = ~v_2296 | ~v_3498;
assign x_1829 = ~v_2297 | v_106;
assign x_1830 = ~v_2297 | ~v_3498;
assign x_1831 = ~v_2298 | v_3497;
assign x_1832 = ~v_2298 | v_106;
assign x_1833 = ~v_2299 | v_3496;
assign x_1834 = ~v_2299 | ~v_3497;
assign x_1835 = ~v_2300 | v_114;
assign x_1836 = ~v_2300 | ~v_3497;
assign x_1837 = ~v_2301 | v_3496;
assign x_1838 = ~v_2301 | v_114;
assign x_1839 = ~v_2302 | v_3495;
assign x_1840 = ~v_2302 | ~v_3496;
assign x_1841 = ~v_2303 | v_121;
assign x_1842 = ~v_2303 | ~v_3496;
assign x_1843 = ~v_2304 | v_3495;
assign x_1844 = ~v_2304 | v_121;
assign x_1845 = ~v_2305 | v_3494;
assign x_1846 = ~v_2305 | ~v_3495;
assign x_1847 = ~v_2306 | v_127;
assign x_1848 = ~v_2306 | ~v_3495;
assign x_1849 = ~v_2307 | v_3494;
assign x_1850 = ~v_2307 | v_127;
assign x_1851 = ~v_2308 | v_136;
assign x_1852 = ~v_2308 | ~v_3494;
assign x_1853 = ~v_2309 | v_132;
assign x_1854 = ~v_2309 | ~v_3494;
assign x_1855 = ~v_2310 | v_136;
assign x_1856 = ~v_2310 | v_132;
assign x_1857 = ~v_2311 | v_3493;
assign x_1858 = ~v_2311 | v_107;
assign x_1859 = ~v_2312 | v_3493;
assign x_1860 = ~v_2312 | v_115;
assign x_1861 = ~v_2313 | v_3493;
assign x_1862 = ~v_2313 | v_122;
assign x_1863 = ~v_2314 | v_3493;
assign x_1864 = ~v_2314 | v_128;
assign x_1865 = ~v_2315 | v_3493;
assign x_1866 = ~v_2315 | v_133;
assign x_1867 = ~v_2316 | v_3493;
assign x_1868 = ~v_2316 | v_137;
assign x_1869 = ~v_2317 | v_3493;
assign x_1870 = ~v_2317 | v_140;
assign x_1871 = ~v_2318 | v_144;
assign x_1872 = ~v_2318 | ~v_3493;
assign x_1873 = ~v_2319 | v_143;
assign x_1874 = ~v_2319 | ~v_3493;
assign x_1875 = ~v_2320 | v_144;
assign x_1876 = ~v_2320 | v_143;
assign x_1877 = ~v_2321 | v_3491;
assign x_1878 = ~v_2321 | ~v_3492;
assign x_1879 = ~v_2322 | v_107;
assign x_1880 = ~v_2322 | ~v_3492;
assign x_1881 = ~v_2323 | v_3491;
assign x_1882 = ~v_2323 | v_107;
assign x_1883 = ~v_2324 | v_3490;
assign x_1884 = ~v_2324 | ~v_3491;
assign x_1885 = ~v_2325 | v_115;
assign x_1886 = ~v_2325 | ~v_3491;
assign x_1887 = ~v_2326 | v_3490;
assign x_1888 = ~v_2326 | v_115;
assign x_1889 = ~v_2327 | v_3489;
assign x_1890 = ~v_2327 | ~v_3490;
assign x_1891 = ~v_2328 | v_122;
assign x_1892 = ~v_2328 | ~v_3490;
assign x_1893 = ~v_2329 | v_3489;
assign x_1894 = ~v_2329 | v_122;
assign x_1895 = ~v_2330 | v_3488;
assign x_1896 = ~v_2330 | ~v_3489;
assign x_1897 = ~v_2331 | v_128;
assign x_1898 = ~v_2331 | ~v_3489;
assign x_1899 = ~v_2332 | v_3488;
assign x_1900 = ~v_2332 | v_128;
assign x_1901 = ~v_2333 | v_3487;
assign x_1902 = ~v_2333 | ~v_3488;
assign x_1903 = ~v_2334 | v_133;
assign x_1904 = ~v_2334 | ~v_3488;
assign x_1905 = ~v_2335 | v_3487;
assign x_1906 = ~v_2335 | v_133;
assign x_1907 = ~v_2336 | v_140;
assign x_1908 = ~v_2336 | ~v_3487;
assign x_1909 = ~v_2337 | v_137;
assign x_1910 = ~v_2337 | ~v_3487;
assign x_1911 = ~v_2338 | v_140;
assign x_1912 = ~v_2338 | v_137;
assign x_1913 = ~v_2339 | v_145;
assign x_1914 = ~v_2339 | v_108;
assign x_1915 = ~v_2340 | v_145;
assign x_1916 = ~v_2340 | v_116;
assign x_1917 = ~v_2341 | v_145;
assign x_1918 = ~v_2341 | v_123;
assign x_1919 = ~v_2342 | v_145;
assign x_1920 = ~v_2342 | v_129;
assign x_1921 = ~v_2343 | v_145;
assign x_1922 = ~v_2343 | v_134;
assign x_1923 = ~v_2344 | v_145;
assign x_1924 = ~v_2344 | v_138;
assign x_1925 = ~v_2345 | v_145;
assign x_1926 = ~v_2345 | v_141;
assign x_1927 = ~v_2346 | v_145;
assign x_1928 = ~v_2346 | v_143;
assign x_1929 = ~v_2347 | v_3485;
assign x_1930 = ~v_2347 | ~v_3486;
assign x_1931 = ~v_2348 | v_108;
assign x_1932 = ~v_2348 | ~v_3486;
assign x_1933 = ~v_2349 | v_3485;
assign x_1934 = ~v_2349 | v_108;
assign x_1935 = ~v_2350 | v_3484;
assign x_1936 = ~v_2350 | ~v_3485;
assign x_1937 = ~v_2351 | v_116;
assign x_1938 = ~v_2351 | ~v_3485;
assign x_1939 = ~v_2352 | v_3484;
assign x_1940 = ~v_2352 | v_116;
assign x_1941 = ~v_2353 | v_3483;
assign x_1942 = ~v_2353 | ~v_3484;
assign x_1943 = ~v_2354 | v_123;
assign x_1944 = ~v_2354 | ~v_3484;
assign x_1945 = ~v_2355 | v_3483;
assign x_1946 = ~v_2355 | v_123;
assign x_1947 = ~v_2356 | v_3482;
assign x_1948 = ~v_2356 | ~v_3483;
assign x_1949 = ~v_2357 | v_129;
assign x_1950 = ~v_2357 | ~v_3483;
assign x_1951 = ~v_2358 | v_3482;
assign x_1952 = ~v_2358 | v_129;
assign x_1953 = ~v_2359 | v_3481;
assign x_1954 = ~v_2359 | ~v_3482;
assign x_1955 = ~v_2360 | v_134;
assign x_1956 = ~v_2360 | ~v_3482;
assign x_1957 = ~v_2361 | v_3481;
assign x_1958 = ~v_2361 | v_134;
assign x_1959 = ~v_2362 | v_3480;
assign x_1960 = ~v_2362 | ~v_3481;
assign x_1961 = ~v_2363 | v_138;
assign x_1962 = ~v_2363 | ~v_3481;
assign x_1963 = ~v_2364 | v_3480;
assign x_1964 = ~v_2364 | v_138;
assign x_1965 = ~v_2365 | v_143;
assign x_1966 = ~v_2365 | ~v_3480;
assign x_1967 = ~v_2366 | v_141;
assign x_1968 = ~v_2366 | ~v_3480;
assign x_1969 = ~v_2367 | v_143;
assign x_1970 = ~v_2367 | v_141;
assign x_1971 = ~v_2368 | v_3478;
assign x_1972 = ~v_2368 | ~v_3479;
assign x_1973 = ~v_2369 | v_109;
assign x_1974 = ~v_2369 | ~v_3479;
assign x_1975 = ~v_2370 | v_3478;
assign x_1976 = ~v_2370 | v_109;
assign x_1977 = ~v_2371 | v_3477;
assign x_1978 = ~v_2371 | ~v_3478;
assign x_1979 = ~v_2372 | v_117;
assign x_1980 = ~v_2372 | ~v_3478;
assign x_1981 = ~v_2373 | v_3477;
assign x_1982 = ~v_2373 | v_117;
assign x_1983 = ~v_2374 | v_3476;
assign x_1984 = ~v_2374 | ~v_3477;
assign x_1985 = ~v_2375 | v_124;
assign x_1986 = ~v_2375 | ~v_3477;
assign x_1987 = ~v_2376 | v_3476;
assign x_1988 = ~v_2376 | v_124;
assign x_1989 = ~v_2377 | v_3475;
assign x_1990 = ~v_2377 | ~v_3476;
assign x_1991 = ~v_2378 | v_130;
assign x_1992 = ~v_2378 | ~v_3476;
assign x_1993 = ~v_2379 | v_3475;
assign x_1994 = ~v_2379 | v_130;
assign x_1995 = ~v_2380 | v_3474;
assign x_1996 = ~v_2380 | ~v_3475;
assign x_1997 = ~v_2381 | v_135;
assign x_1998 = ~v_2381 | ~v_3475;
assign x_1999 = ~v_2382 | v_3474;
assign x_2000 = ~v_2382 | v_135;
assign x_2001 = ~v_2383 | v_3473;
assign x_2002 = ~v_2383 | ~v_3474;
assign x_2003 = ~v_2384 | v_139;
assign x_2004 = ~v_2384 | ~v_3474;
assign x_2005 = ~v_2385 | v_3473;
assign x_2006 = ~v_2385 | v_139;
assign x_2007 = ~v_2386 | v_3472;
assign x_2008 = ~v_2386 | ~v_3473;
assign x_2009 = ~v_2387 | v_142;
assign x_2010 = ~v_2387 | ~v_3473;
assign x_2011 = ~v_2388 | v_3472;
assign x_2012 = ~v_2388 | v_142;
assign x_2013 = ~v_2389 | v_145;
assign x_2014 = ~v_2389 | ~v_3472;
assign x_2015 = ~v_2390 | v_144;
assign x_2016 = ~v_2390 | ~v_3472;
assign x_2017 = ~v_2391 | v_145;
assign x_2018 = ~v_2391 | v_144;
assign x_2019 = ~v_2392 | v_3704;
assign x_2020 = ~v_2392 | ~v_3705;
assign x_2021 = ~v_2393 | v_154;
assign x_2022 = ~v_2393 | ~v_3705;
assign x_2023 = ~v_2394 | v_3704;
assign x_2024 = ~v_2394 | v_154;
assign x_2025 = ~v_2395 | v_3703;
assign x_2026 = ~v_2395 | ~v_3704;
assign x_2027 = ~v_2396 | v_153;
assign x_2028 = ~v_2396 | ~v_3704;
assign x_2029 = ~v_2397 | v_3703;
assign x_2030 = ~v_2397 | v_153;
assign x_2031 = ~v_2398 | v_3702;
assign x_2032 = ~v_2398 | ~v_3703;
assign x_2033 = ~v_2399 | v_152;
assign x_2034 = ~v_2399 | ~v_3703;
assign x_2035 = ~v_2400 | v_3702;
assign x_2036 = ~v_2400 | v_152;
assign x_2037 = ~v_2401 | v_3701;
assign x_2038 = ~v_2401 | ~v_3702;
assign x_2039 = ~v_2402 | v_151;
assign x_2040 = ~v_2402 | ~v_3702;
assign x_2041 = ~v_2403 | v_3701;
assign x_2042 = ~v_2403 | v_151;
assign x_2043 = ~v_2404 | v_3700;
assign x_2044 = ~v_2404 | ~v_3701;
assign x_2045 = ~v_2405 | v_150;
assign x_2046 = ~v_2405 | ~v_3701;
assign x_2047 = ~v_2406 | v_3700;
assign x_2048 = ~v_2406 | v_150;
assign x_2049 = ~v_2407 | v_3699;
assign x_2050 = ~v_2407 | ~v_3700;
assign x_2051 = ~v_2408 | v_149;
assign x_2052 = ~v_2408 | ~v_3700;
assign x_2053 = ~v_2409 | v_3699;
assign x_2054 = ~v_2409 | v_149;
assign x_2055 = ~v_2410 | v_3698;
assign x_2056 = ~v_2410 | ~v_3699;
assign x_2057 = ~v_2411 | v_148;
assign x_2058 = ~v_2411 | ~v_3699;
assign x_2059 = ~v_2412 | v_3698;
assign x_2060 = ~v_2412 | v_148;
assign x_2061 = ~v_2413 | v_146;
assign x_2062 = ~v_2413 | ~v_3698;
assign x_2063 = ~v_2414 | v_147;
assign x_2064 = ~v_2414 | ~v_3698;
assign x_2065 = ~v_2415 | v_146;
assign x_2066 = ~v_2415 | v_147;
assign x_2067 = ~v_2416 | v_3696;
assign x_2068 = ~v_2416 | ~v_3697;
assign x_2069 = ~v_2417 | v_162;
assign x_2070 = ~v_2417 | ~v_3697;
assign x_2071 = ~v_2418 | v_3696;
assign x_2072 = ~v_2418 | v_162;
assign x_2073 = ~v_2419 | v_3695;
assign x_2074 = ~v_2419 | ~v_3696;
assign x_2075 = ~v_2420 | v_161;
assign x_2076 = ~v_2420 | ~v_3696;
assign x_2077 = ~v_2421 | v_3695;
assign x_2078 = ~v_2421 | v_161;
assign x_2079 = ~v_2422 | v_3694;
assign x_2080 = ~v_2422 | ~v_3695;
assign x_2081 = ~v_2423 | v_160;
assign x_2082 = ~v_2423 | ~v_3695;
assign x_2083 = ~v_2424 | v_3694;
assign x_2084 = ~v_2424 | v_160;
assign x_2085 = ~v_2425 | v_3693;
assign x_2086 = ~v_2425 | ~v_3694;
assign x_2087 = ~v_2426 | v_159;
assign x_2088 = ~v_2426 | ~v_3694;
assign x_2089 = ~v_2427 | v_3693;
assign x_2090 = ~v_2427 | v_159;
assign x_2091 = ~v_2428 | v_3692;
assign x_2092 = ~v_2428 | ~v_3693;
assign x_2093 = ~v_2429 | v_158;
assign x_2094 = ~v_2429 | ~v_3693;
assign x_2095 = ~v_2430 | v_3692;
assign x_2096 = ~v_2430 | v_158;
assign x_2097 = ~v_2431 | v_3691;
assign x_2098 = ~v_2431 | ~v_3692;
assign x_2099 = ~v_2432 | v_157;
assign x_2100 = ~v_2432 | ~v_3692;
assign x_2101 = ~v_2433 | v_3691;
assign x_2102 = ~v_2433 | v_157;
assign x_2103 = ~v_2434 | v_155;
assign x_2104 = ~v_2434 | ~v_3691;
assign x_2105 = ~v_2435 | v_156;
assign x_2106 = ~v_2435 | ~v_3691;
assign x_2107 = ~v_2436 | v_155;
assign x_2108 = ~v_2436 | v_156;
assign x_2109 = ~v_2437 | v_146;
assign x_2110 = ~v_2437 | v_162;
assign x_2111 = ~v_2438 | v_146;
assign x_2112 = ~v_2438 | v_161;
assign x_2113 = ~v_2439 | v_146;
assign x_2114 = ~v_2439 | v_160;
assign x_2115 = ~v_2440 | v_146;
assign x_2116 = ~v_2440 | v_159;
assign x_2117 = ~v_2441 | v_146;
assign x_2118 = ~v_2441 | v_158;
assign x_2119 = ~v_2442 | v_146;
assign x_2120 = ~v_2442 | v_157;
assign x_2121 = ~v_2443 | v_146;
assign x_2122 = ~v_2443 | v_156;
assign x_2123 = ~v_2444 | v_146;
assign x_2124 = ~v_2444 | v_155;
assign x_2125 = ~v_2445 | v_3689;
assign x_2126 = ~v_2445 | ~v_3690;
assign x_2127 = ~v_2446 | v_169;
assign x_2128 = ~v_2446 | ~v_3690;
assign x_2129 = ~v_2447 | v_3689;
assign x_2130 = ~v_2447 | v_169;
assign x_2131 = ~v_2448 | v_3688;
assign x_2132 = ~v_2448 | ~v_3689;
assign x_2133 = ~v_2449 | v_168;
assign x_2134 = ~v_2449 | ~v_3689;
assign x_2135 = ~v_2450 | v_3688;
assign x_2136 = ~v_2450 | v_168;
assign x_2137 = ~v_2451 | v_3687;
assign x_2138 = ~v_2451 | ~v_3688;
assign x_2139 = ~v_2452 | v_167;
assign x_2140 = ~v_2452 | ~v_3688;
assign x_2141 = ~v_2453 | v_3687;
assign x_2142 = ~v_2453 | v_167;
assign x_2143 = ~v_2454 | v_3686;
assign x_2144 = ~v_2454 | ~v_3687;
assign x_2145 = ~v_2455 | v_166;
assign x_2146 = ~v_2455 | ~v_3687;
assign x_2147 = ~v_2456 | v_3686;
assign x_2148 = ~v_2456 | v_166;
assign x_2149 = ~v_2457 | v_3685;
assign x_2150 = ~v_2457 | ~v_3686;
assign x_2151 = ~v_2458 | v_165;
assign x_2152 = ~v_2458 | ~v_3686;
assign x_2153 = ~v_2459 | v_3685;
assign x_2154 = ~v_2459 | v_165;
assign x_2155 = ~v_2460 | v_163;
assign x_2156 = ~v_2460 | ~v_3685;
assign x_2157 = ~v_2461 | v_164;
assign x_2158 = ~v_2461 | ~v_3685;
assign x_2159 = ~v_2462 | v_163;
assign x_2160 = ~v_2462 | v_164;
assign x_2161 = ~v_2463 | v_3684;
assign x_2162 = ~v_2463 | v_169;
assign x_2163 = ~v_2464 | v_3684;
assign x_2164 = ~v_2464 | v_168;
assign x_2165 = ~v_2465 | v_3684;
assign x_2166 = ~v_2465 | v_167;
assign x_2167 = ~v_2466 | v_3684;
assign x_2168 = ~v_2466 | v_166;
assign x_2169 = ~v_2467 | v_3684;
assign x_2170 = ~v_2467 | v_165;
assign x_2171 = ~v_2468 | v_3684;
assign x_2172 = ~v_2468 | v_164;
assign x_2173 = ~v_2469 | v_3684;
assign x_2174 = ~v_2469 | v_163;
assign x_2175 = ~v_2470 | v_147;
assign x_2176 = ~v_2470 | ~v_3684;
assign x_2177 = ~v_2471 | v_155;
assign x_2178 = ~v_2471 | ~v_3684;
assign x_2179 = ~v_2472 | v_147;
assign x_2180 = ~v_2472 | v_155;
assign x_2181 = ~v_2473 | v_3682;
assign x_2182 = ~v_2473 | ~v_3683;
assign x_2183 = ~v_2474 | v_175;
assign x_2184 = ~v_2474 | ~v_3683;
assign x_2185 = ~v_2475 | v_3682;
assign x_2186 = ~v_2475 | v_175;
assign x_2187 = ~v_2476 | v_3681;
assign x_2188 = ~v_2476 | ~v_3682;
assign x_2189 = ~v_2477 | v_174;
assign x_2190 = ~v_2477 | ~v_3682;
assign x_2191 = ~v_2478 | v_3681;
assign x_2192 = ~v_2478 | v_174;
assign x_2193 = ~v_2479 | v_3680;
assign x_2194 = ~v_2479 | ~v_3681;
assign x_2195 = ~v_2480 | v_173;
assign x_2196 = ~v_2480 | ~v_3681;
assign x_2197 = ~v_2481 | v_3680;
assign x_2198 = ~v_2481 | v_173;
assign x_2199 = ~v_2482 | v_3679;
assign x_2200 = ~v_2482 | ~v_3680;
assign x_2201 = ~v_2483 | v_172;
assign x_2202 = ~v_2483 | ~v_3680;
assign x_2203 = ~v_2484 | v_3679;
assign x_2204 = ~v_2484 | v_172;
assign x_2205 = ~v_2485 | v_170;
assign x_2206 = ~v_2485 | ~v_3679;
assign x_2207 = ~v_2486 | v_171;
assign x_2208 = ~v_2486 | ~v_3679;
assign x_2209 = ~v_2487 | v_170;
assign x_2210 = ~v_2487 | v_171;
assign x_2211 = ~v_2488 | v_3678;
assign x_2212 = ~v_2488 | v_175;
assign x_2213 = ~v_2489 | v_3678;
assign x_2214 = ~v_2489 | v_174;
assign x_2215 = ~v_2490 | v_3678;
assign x_2216 = ~v_2490 | v_173;
assign x_2217 = ~v_2491 | v_3678;
assign x_2218 = ~v_2491 | v_172;
assign x_2219 = ~v_2492 | v_3678;
assign x_2220 = ~v_2492 | v_171;
assign x_2221 = ~v_2493 | v_3678;
assign x_2222 = ~v_2493 | v_170;
assign x_2223 = ~v_2494 | v_3677;
assign x_2224 = ~v_2494 | ~v_3678;
assign x_2225 = ~v_2495 | v_163;
assign x_2226 = ~v_2495 | ~v_3678;
assign x_2227 = ~v_2496 | v_3677;
assign x_2228 = ~v_2496 | v_163;
assign x_2229 = ~v_2497 | v_148;
assign x_2230 = ~v_2497 | ~v_3677;
assign x_2231 = ~v_2498 | v_156;
assign x_2232 = ~v_2498 | ~v_3677;
assign x_2233 = ~v_2499 | v_148;
assign x_2234 = ~v_2499 | v_156;
assign x_2235 = ~v_2500 | v_3675;
assign x_2236 = ~v_2500 | ~v_3676;
assign x_2237 = ~v_2501 | v_180;
assign x_2238 = ~v_2501 | ~v_3676;
assign x_2239 = ~v_2502 | v_3675;
assign x_2240 = ~v_2502 | v_180;
assign x_2241 = ~v_2503 | v_3674;
assign x_2242 = ~v_2503 | ~v_3675;
assign x_2243 = ~v_2504 | v_179;
assign x_2244 = ~v_2504 | ~v_3675;
assign x_2245 = ~v_2505 | v_3674;
assign x_2246 = ~v_2505 | v_179;
assign x_2247 = ~v_2506 | v_3673;
assign x_2248 = ~v_2506 | ~v_3674;
assign x_2249 = ~v_2507 | v_178;
assign x_2250 = ~v_2507 | ~v_3674;
assign x_2251 = ~v_2508 | v_3673;
assign x_2252 = ~v_2508 | v_178;
assign x_2253 = ~v_2509 | v_176;
assign x_2254 = ~v_2509 | ~v_3673;
assign x_2255 = ~v_2510 | v_177;
assign x_2256 = ~v_2510 | ~v_3673;
assign x_2257 = ~v_2511 | v_176;
assign x_2258 = ~v_2511 | v_177;
assign x_2259 = ~v_2512 | v_3672;
assign x_2260 = ~v_2512 | v_180;
assign x_2261 = ~v_2513 | v_3672;
assign x_2262 = ~v_2513 | v_179;
assign x_2263 = ~v_2514 | v_3672;
assign x_2264 = ~v_2514 | v_178;
assign x_2265 = ~v_2515 | v_3672;
assign x_2266 = ~v_2515 | v_177;
assign x_2267 = ~v_2516 | v_3672;
assign x_2268 = ~v_2516 | v_176;
assign x_2269 = ~v_2517 | v_3671;
assign x_2270 = ~v_2517 | ~v_3672;
assign x_2271 = ~v_2518 | v_170;
assign x_2272 = ~v_2518 | ~v_3672;
assign x_2273 = ~v_2519 | v_3671;
assign x_2274 = ~v_2519 | v_170;
assign x_2275 = ~v_2520 | v_3670;
assign x_2276 = ~v_2520 | ~v_3671;
assign x_2277 = ~v_2521 | v_164;
assign x_2278 = ~v_2521 | ~v_3671;
assign x_2279 = ~v_2522 | v_3670;
assign x_2280 = ~v_2522 | v_164;
assign x_2281 = ~v_2523 | v_149;
assign x_2282 = ~v_2523 | ~v_3670;
assign x_2283 = ~v_2524 | v_157;
assign x_2284 = ~v_2524 | ~v_3670;
assign x_2285 = ~v_2525 | v_149;
assign x_2286 = ~v_2525 | v_157;
assign x_2287 = ~v_2526 | v_3668;
assign x_2288 = ~v_2526 | ~v_3669;
assign x_2289 = ~v_2527 | v_184;
assign x_2290 = ~v_2527 | ~v_3669;
assign x_2291 = ~v_2528 | v_3668;
assign x_2292 = ~v_2528 | v_184;
assign x_2293 = ~v_2529 | v_3667;
assign x_2294 = ~v_2529 | ~v_3668;
assign x_2295 = ~v_2530 | v_183;
assign x_2296 = ~v_2530 | ~v_3668;
assign x_2297 = ~v_2531 | v_3667;
assign x_2298 = ~v_2531 | v_183;
assign x_2299 = ~v_2532 | v_181;
assign x_2300 = ~v_2532 | ~v_3667;
assign x_2301 = ~v_2533 | v_182;
assign x_2302 = ~v_2533 | ~v_3667;
assign x_2303 = ~v_2534 | v_181;
assign x_2304 = ~v_2534 | v_182;
assign x_2305 = ~v_2535 | v_3666;
assign x_2306 = ~v_2535 | v_184;
assign x_2307 = ~v_2536 | v_3666;
assign x_2308 = ~v_2536 | v_183;
assign x_2309 = ~v_2537 | v_3666;
assign x_2310 = ~v_2537 | v_182;
assign x_2311 = ~v_2538 | v_3666;
assign x_2312 = ~v_2538 | v_181;
assign x_2313 = ~v_2539 | v_3665;
assign x_2314 = ~v_2539 | ~v_3666;
assign x_2315 = ~v_2540 | v_176;
assign x_2316 = ~v_2540 | ~v_3666;
assign x_2317 = ~v_2541 | v_3665;
assign x_2318 = ~v_2541 | v_176;
assign x_2319 = ~v_2542 | v_3664;
assign x_2320 = ~v_2542 | ~v_3665;
assign x_2321 = ~v_2543 | v_171;
assign x_2322 = ~v_2543 | ~v_3665;
assign x_2323 = ~v_2544 | v_3664;
assign x_2324 = ~v_2544 | v_171;
assign x_2325 = ~v_2545 | v_3663;
assign x_2326 = ~v_2545 | ~v_3664;
assign x_2327 = ~v_2546 | v_165;
assign x_2328 = ~v_2546 | ~v_3664;
assign x_2329 = ~v_2547 | v_3663;
assign x_2330 = ~v_2547 | v_165;
assign x_2331 = ~v_2548 | v_150;
assign x_2332 = ~v_2548 | ~v_3663;
assign x_2333 = ~v_2549 | v_158;
assign x_2334 = ~v_2549 | ~v_3663;
assign x_2335 = ~v_2550 | v_150;
assign x_2336 = ~v_2550 | v_158;
assign x_2337 = ~v_2551 | v_3661;
assign x_2338 = ~v_2551 | ~v_3662;
assign x_2339 = ~v_2552 | v_187;
assign x_2340 = ~v_2552 | ~v_3662;
assign x_2341 = ~v_2553 | v_3661;
assign x_2342 = ~v_2553 | v_187;
assign x_2343 = ~v_2554 | v_185;
assign x_2344 = ~v_2554 | ~v_3661;
assign x_2345 = ~v_2555 | v_186;
assign x_2346 = ~v_2555 | ~v_3661;
assign x_2347 = ~v_2556 | v_185;
assign x_2348 = ~v_2556 | v_186;
assign x_2349 = ~v_2557 | v_3660;
assign x_2350 = ~v_2557 | v_187;
assign x_2351 = ~v_2558 | v_3660;
assign x_2352 = ~v_2558 | v_186;
assign x_2353 = ~v_2559 | v_3660;
assign x_2354 = ~v_2559 | v_185;
assign x_2355 = ~v_2560 | v_3659;
assign x_2356 = ~v_2560 | ~v_3660;
assign x_2357 = ~v_2561 | v_181;
assign x_2358 = ~v_2561 | ~v_3660;
assign x_2359 = ~v_2562 | v_3659;
assign x_2360 = ~v_2562 | v_181;
assign x_2361 = ~v_2563 | v_3658;
assign x_2362 = ~v_2563 | ~v_3659;
assign x_2363 = ~v_2564 | v_177;
assign x_2364 = ~v_2564 | ~v_3659;
assign x_2365 = ~v_2565 | v_3658;
assign x_2366 = ~v_2565 | v_177;
assign x_2367 = ~v_2566 | v_3657;
assign x_2368 = ~v_2566 | ~v_3658;
assign x_2369 = ~v_2567 | v_172;
assign x_2370 = ~v_2567 | ~v_3658;
assign x_2371 = ~v_2568 | v_3657;
assign x_2372 = ~v_2568 | v_172;
assign x_2373 = ~v_2569 | v_3656;
assign x_2374 = ~v_2569 | ~v_3657;
assign x_2375 = ~v_2570 | v_166;
assign x_2376 = ~v_2570 | ~v_3657;
assign x_2377 = ~v_2571 | v_3656;
assign x_2378 = ~v_2571 | v_166;
assign x_2379 = ~v_2572 | v_151;
assign x_2380 = ~v_2572 | ~v_3656;
assign x_2381 = ~v_2573 | v_159;
assign x_2382 = ~v_2573 | ~v_3656;
assign x_2383 = ~v_2574 | v_151;
assign x_2384 = ~v_2574 | v_159;
assign x_2385 = ~v_2575 | v_188;
assign x_2386 = ~v_2575 | ~v_3655;
assign x_2387 = ~v_2576 | v_189;
assign x_2388 = ~v_2576 | ~v_3655;
assign x_2389 = ~v_2577 | v_188;
assign x_2390 = ~v_2577 | v_189;
assign x_2391 = ~v_2578 | v_3654;
assign x_2392 = ~v_2578 | v_189;
assign x_2393 = ~v_2579 | v_3654;
assign x_2394 = ~v_2579 | v_188;
assign x_2395 = ~v_2580 | v_3653;
assign x_2396 = ~v_2580 | ~v_3654;
assign x_2397 = ~v_2581 | v_185;
assign x_2398 = ~v_2581 | ~v_3654;
assign x_2399 = ~v_2582 | v_3653;
assign x_2400 = ~v_2582 | v_185;
assign x_2401 = ~v_2583 | v_3652;
assign x_2402 = ~v_2583 | ~v_3653;
assign x_2403 = ~v_2584 | v_182;
assign x_2404 = ~v_2584 | ~v_3653;
assign x_2405 = ~v_2585 | v_3652;
assign x_2406 = ~v_2585 | v_182;
assign x_2407 = ~v_2586 | v_3651;
assign x_2408 = ~v_2586 | ~v_3652;
assign x_2409 = ~v_2587 | v_178;
assign x_2410 = ~v_2587 | ~v_3652;
assign x_2411 = ~v_2588 | v_3651;
assign x_2412 = ~v_2588 | v_178;
assign x_2413 = ~v_2589 | v_3650;
assign x_2414 = ~v_2589 | ~v_3651;
assign x_2415 = ~v_2590 | v_173;
assign x_2416 = ~v_2590 | ~v_3651;
assign x_2417 = ~v_2591 | v_3650;
assign x_2418 = ~v_2591 | v_173;
assign x_2419 = ~v_2592 | v_3649;
assign x_2420 = ~v_2592 | ~v_3650;
assign x_2421 = ~v_2593 | v_167;
assign x_2422 = ~v_2593 | ~v_3650;
assign x_2423 = ~v_2594 | v_3649;
assign x_2424 = ~v_2594 | v_167;
assign x_2425 = ~v_2595 | v_152;
assign x_2426 = ~v_2595 | ~v_3649;
assign x_2427 = ~v_2596 | v_160;
assign x_2428 = ~v_2596 | ~v_3649;
assign x_2429 = ~v_2597 | v_152;
assign x_2430 = ~v_2597 | v_160;
assign x_2431 = ~v_2598 | v_3648;
assign x_2432 = ~v_2598 | v_190;
assign x_2433 = ~v_2599 | v_3647;
assign x_2434 = ~v_2599 | ~v_3648;
assign x_2435 = ~v_2600 | v_188;
assign x_2436 = ~v_2600 | ~v_3648;
assign x_2437 = ~v_2601 | v_3647;
assign x_2438 = ~v_2601 | v_188;
assign x_2439 = ~v_2602 | v_3646;
assign x_2440 = ~v_2602 | ~v_3647;
assign x_2441 = ~v_2603 | v_186;
assign x_2442 = ~v_2603 | ~v_3647;
assign x_2443 = ~v_2604 | v_3646;
assign x_2444 = ~v_2604 | v_186;
assign x_2445 = ~v_2605 | v_3645;
assign x_2446 = ~v_2605 | ~v_3646;
assign x_2447 = ~v_2606 | v_183;
assign x_2448 = ~v_2606 | ~v_3646;
assign x_2449 = ~v_2607 | v_3645;
assign x_2450 = ~v_2607 | v_183;
assign x_2451 = ~v_2608 | v_3644;
assign x_2452 = ~v_2608 | ~v_3645;
assign x_2453 = ~v_2609 | v_179;
assign x_2454 = ~v_2609 | ~v_3645;
assign x_2455 = ~v_2610 | v_3644;
assign x_2456 = ~v_2610 | v_179;
assign x_2457 = ~v_2611 | v_3643;
assign x_2458 = ~v_2611 | ~v_3644;
assign x_2459 = ~v_2612 | v_174;
assign x_2460 = ~v_2612 | ~v_3644;
assign x_2461 = ~v_2613 | v_3643;
assign x_2462 = ~v_2613 | v_174;
assign x_2463 = ~v_2614 | v_3642;
assign x_2464 = ~v_2614 | ~v_3643;
assign x_2465 = ~v_2615 | v_168;
assign x_2466 = ~v_2615 | ~v_3643;
assign x_2467 = ~v_2616 | v_3642;
assign x_2468 = ~v_2616 | v_168;
assign x_2469 = ~v_2617 | v_153;
assign x_2470 = ~v_2617 | ~v_3642;
assign x_2471 = ~v_2618 | v_161;
assign x_2472 = ~v_2618 | ~v_3642;
assign x_2473 = ~v_2619 | v_153;
assign x_2474 = ~v_2619 | v_161;
assign x_2475 = ~v_2620 | v_3640;
assign x_2476 = ~v_2620 | ~v_3641;
assign x_2477 = ~v_2621 | v_190;
assign x_2478 = ~v_2621 | ~v_3641;
assign x_2479 = ~v_2622 | v_3640;
assign x_2480 = ~v_2622 | v_190;
assign x_2481 = ~v_2623 | v_3639;
assign x_2482 = ~v_2623 | ~v_3640;
assign x_2483 = ~v_2624 | v_189;
assign x_2484 = ~v_2624 | ~v_3640;
assign x_2485 = ~v_2625 | v_3639;
assign x_2486 = ~v_2625 | v_189;
assign x_2487 = ~v_2626 | v_3638;
assign x_2488 = ~v_2626 | ~v_3639;
assign x_2489 = ~v_2627 | v_187;
assign x_2490 = ~v_2627 | ~v_3639;
assign x_2491 = ~v_2628 | v_3638;
assign x_2492 = ~v_2628 | v_187;
assign x_2493 = ~v_2629 | v_3637;
assign x_2494 = ~v_2629 | ~v_3638;
assign x_2495 = ~v_2630 | v_184;
assign x_2496 = ~v_2630 | ~v_3638;
assign x_2497 = ~v_2631 | v_3637;
assign x_2498 = ~v_2631 | v_184;
assign x_2499 = ~v_2632 | v_3636;
assign x_2500 = ~v_2632 | ~v_3637;
assign x_2501 = ~v_2633 | v_180;
assign x_2502 = ~v_2633 | ~v_3637;
assign x_2503 = ~v_2634 | v_3636;
assign x_2504 = ~v_2634 | v_180;
assign x_2505 = ~v_2635 | v_3635;
assign x_2506 = ~v_2635 | ~v_3636;
assign x_2507 = ~v_2636 | v_175;
assign x_2508 = ~v_2636 | ~v_3636;
assign x_2509 = ~v_2637 | v_3635;
assign x_2510 = ~v_2637 | v_175;
assign x_2511 = ~v_2638 | v_3634;
assign x_2512 = ~v_2638 | ~v_3635;
assign x_2513 = ~v_2639 | v_169;
assign x_2514 = ~v_2639 | ~v_3635;
assign x_2515 = ~v_2640 | v_3634;
assign x_2516 = ~v_2640 | v_169;
assign x_2517 = ~v_2641 | v_154;
assign x_2518 = ~v_2641 | ~v_3634;
assign x_2519 = ~v_2642 | v_162;
assign x_2520 = ~v_2642 | ~v_3634;
assign x_2521 = ~v_2643 | v_154;
assign x_2522 = ~v_2643 | v_162;
assign x_2523 = ~v_2644 | v_3776;
assign x_2524 = ~v_2644 | ~v_3777;
assign x_2525 = ~v_2645 | v_146;
assign x_2526 = ~v_2645 | ~v_3777;
assign x_2527 = ~v_2646 | v_3776;
assign x_2528 = ~v_2646 | v_146;
assign x_2529 = ~v_2647 | v_3775;
assign x_2530 = ~v_2647 | ~v_3776;
assign x_2531 = ~v_2648 | v_147;
assign x_2532 = ~v_2648 | ~v_3776;
assign x_2533 = ~v_2649 | v_3775;
assign x_2534 = ~v_2649 | v_147;
assign x_2535 = ~v_2650 | v_3774;
assign x_2536 = ~v_2650 | ~v_3775;
assign x_2537 = ~v_2651 | v_148;
assign x_2538 = ~v_2651 | ~v_3775;
assign x_2539 = ~v_2652 | v_3774;
assign x_2540 = ~v_2652 | v_148;
assign x_2541 = ~v_2653 | v_3773;
assign x_2542 = ~v_2653 | ~v_3774;
assign x_2543 = ~v_2654 | v_149;
assign x_2544 = ~v_2654 | ~v_3774;
assign x_2545 = ~v_2655 | v_3773;
assign x_2546 = ~v_2655 | v_149;
assign x_2547 = ~v_2656 | v_3772;
assign x_2548 = ~v_2656 | ~v_3773;
assign x_2549 = ~v_2657 | v_150;
assign x_2550 = ~v_2657 | ~v_3773;
assign x_2551 = ~v_2658 | v_3772;
assign x_2552 = ~v_2658 | v_150;
assign x_2553 = ~v_2659 | v_3771;
assign x_2554 = ~v_2659 | ~v_3772;
assign x_2555 = ~v_2660 | v_151;
assign x_2556 = ~v_2660 | ~v_3772;
assign x_2557 = ~v_2661 | v_3771;
assign x_2558 = ~v_2661 | v_151;
assign x_2559 = ~v_2662 | v_3770;
assign x_2560 = ~v_2662 | ~v_3771;
assign x_2561 = ~v_2663 | v_152;
assign x_2562 = ~v_2663 | ~v_3771;
assign x_2563 = ~v_2664 | v_3770;
assign x_2564 = ~v_2664 | v_152;
assign x_2565 = ~v_2665 | v_154;
assign x_2566 = ~v_2665 | ~v_3770;
assign x_2567 = ~v_2666 | v_153;
assign x_2568 = ~v_2666 | ~v_3770;
assign x_2569 = ~v_2667 | v_154;
assign x_2570 = ~v_2667 | v_153;
assign x_2571 = ~v_2668 | v_3769;
assign x_2572 = ~v_2668 | v_146;
assign x_2573 = ~v_2669 | v_3768;
assign x_2574 = ~v_2669 | ~v_3769;
assign x_2575 = ~v_2670 | v_155;
assign x_2576 = ~v_2670 | ~v_3769;
assign x_2577 = ~v_2671 | v_3768;
assign x_2578 = ~v_2671 | v_155;
assign x_2579 = ~v_2672 | v_3767;
assign x_2580 = ~v_2672 | ~v_3768;
assign x_2581 = ~v_2673 | v_156;
assign x_2582 = ~v_2673 | ~v_3768;
assign x_2583 = ~v_2674 | v_3767;
assign x_2584 = ~v_2674 | v_156;
assign x_2585 = ~v_2675 | v_3766;
assign x_2586 = ~v_2675 | ~v_3767;
assign x_2587 = ~v_2676 | v_157;
assign x_2588 = ~v_2676 | ~v_3767;
assign x_2589 = ~v_2677 | v_3766;
assign x_2590 = ~v_2677 | v_157;
assign x_2591 = ~v_2678 | v_3765;
assign x_2592 = ~v_2678 | ~v_3766;
assign x_2593 = ~v_2679 | v_158;
assign x_2594 = ~v_2679 | ~v_3766;
assign x_2595 = ~v_2680 | v_3765;
assign x_2596 = ~v_2680 | v_158;
assign x_2597 = ~v_2681 | v_3764;
assign x_2598 = ~v_2681 | ~v_3765;
assign x_2599 = ~v_2682 | v_159;
assign x_2600 = ~v_2682 | ~v_3765;
assign x_2601 = ~v_2683 | v_3764;
assign x_2602 = ~v_2683 | v_159;
assign x_2603 = ~v_2684 | v_3763;
assign x_2604 = ~v_2684 | ~v_3764;
assign x_2605 = ~v_2685 | v_160;
assign x_2606 = ~v_2685 | ~v_3764;
assign x_2607 = ~v_2686 | v_3763;
assign x_2608 = ~v_2686 | v_160;
assign x_2609 = ~v_2687 | v_162;
assign x_2610 = ~v_2687 | ~v_3763;
assign x_2611 = ~v_2688 | v_161;
assign x_2612 = ~v_2688 | ~v_3763;
assign x_2613 = ~v_2689 | v_162;
assign x_2614 = ~v_2689 | v_161;
assign x_2615 = ~v_2690 | v_3762;
assign x_2616 = ~v_2690 | v_147;
assign x_2617 = ~v_2691 | v_3762;
assign x_2618 = ~v_2691 | v_155;
assign x_2619 = ~v_2692 | v_3761;
assign x_2620 = ~v_2692 | ~v_3762;
assign x_2621 = ~v_2693 | v_163;
assign x_2622 = ~v_2693 | ~v_3762;
assign x_2623 = ~v_2694 | v_3761;
assign x_2624 = ~v_2694 | v_163;
assign x_2625 = ~v_2695 | v_3760;
assign x_2626 = ~v_2695 | ~v_3761;
assign x_2627 = ~v_2696 | v_164;
assign x_2628 = ~v_2696 | ~v_3761;
assign x_2629 = ~v_2697 | v_3760;
assign x_2630 = ~v_2697 | v_164;
assign x_2631 = ~v_2698 | v_3759;
assign x_2632 = ~v_2698 | ~v_3760;
assign x_2633 = ~v_2699 | v_165;
assign x_2634 = ~v_2699 | ~v_3760;
assign x_2635 = ~v_2700 | v_3759;
assign x_2636 = ~v_2700 | v_165;
assign x_2637 = ~v_2701 | v_3758;
assign x_2638 = ~v_2701 | ~v_3759;
assign x_2639 = ~v_2702 | v_166;
assign x_2640 = ~v_2702 | ~v_3759;
assign x_2641 = ~v_2703 | v_3758;
assign x_2642 = ~v_2703 | v_166;
assign x_2643 = ~v_2704 | v_3757;
assign x_2644 = ~v_2704 | ~v_3758;
assign x_2645 = ~v_2705 | v_167;
assign x_2646 = ~v_2705 | ~v_3758;
assign x_2647 = ~v_2706 | v_3757;
assign x_2648 = ~v_2706 | v_167;
assign x_2649 = ~v_2707 | v_169;
assign x_2650 = ~v_2707 | ~v_3757;
assign x_2651 = ~v_2708 | v_168;
assign x_2652 = ~v_2708 | ~v_3757;
assign x_2653 = ~v_2709 | v_169;
assign x_2654 = ~v_2709 | v_168;
assign x_2655 = ~v_2710 | v_155;
assign x_2656 = ~v_2710 | ~v_3756;
assign x_2657 = ~v_2711 | v_147;
assign x_2658 = ~v_2711 | ~v_3756;
assign x_2659 = ~v_2712 | v_155;
assign x_2660 = ~v_2712 | v_147;
assign x_2661 = ~v_2713 | v_3755;
assign x_2662 = ~v_2713 | v_148;
assign x_2663 = ~v_2714 | v_3755;
assign x_2664 = ~v_2714 | v_156;
assign x_2665 = ~v_2715 | v_3755;
assign x_2666 = ~v_2715 | v_163;
assign x_2667 = ~v_2716 | v_3754;
assign x_2668 = ~v_2716 | ~v_3755;
assign x_2669 = ~v_2717 | v_170;
assign x_2670 = ~v_2717 | ~v_3755;
assign x_2671 = ~v_2718 | v_3754;
assign x_2672 = ~v_2718 | v_170;
assign x_2673 = ~v_2719 | v_3753;
assign x_2674 = ~v_2719 | ~v_3754;
assign x_2675 = ~v_2720 | v_171;
assign x_2676 = ~v_2720 | ~v_3754;
assign x_2677 = ~v_2721 | v_3753;
assign x_2678 = ~v_2721 | v_171;
assign x_2679 = ~v_2722 | v_3752;
assign x_2680 = ~v_2722 | ~v_3753;
assign x_2681 = ~v_2723 | v_172;
assign x_2682 = ~v_2723 | ~v_3753;
assign x_2683 = ~v_2724 | v_3752;
assign x_2684 = ~v_2724 | v_172;
assign x_2685 = ~v_2725 | v_3751;
assign x_2686 = ~v_2725 | ~v_3752;
assign x_2687 = ~v_2726 | v_173;
assign x_2688 = ~v_2726 | ~v_3752;
assign x_2689 = ~v_2727 | v_3751;
assign x_2690 = ~v_2727 | v_173;
assign x_2691 = ~v_2728 | v_175;
assign x_2692 = ~v_2728 | ~v_3751;
assign x_2693 = ~v_2729 | v_174;
assign x_2694 = ~v_2729 | ~v_3751;
assign x_2695 = ~v_2730 | v_175;
assign x_2696 = ~v_2730 | v_174;
assign x_2697 = ~v_2731 | v_3749;
assign x_2698 = ~v_2731 | ~v_3750;
assign x_2699 = ~v_2732 | v_148;
assign x_2700 = ~v_2732 | ~v_3750;
assign x_2701 = ~v_2733 | v_3749;
assign x_2702 = ~v_2733 | v_148;
assign x_2703 = ~v_2734 | v_163;
assign x_2704 = ~v_2734 | ~v_3749;
assign x_2705 = ~v_2735 | v_156;
assign x_2706 = ~v_2735 | ~v_3749;
assign x_2707 = ~v_2736 | v_163;
assign x_2708 = ~v_2736 | v_156;
assign x_2709 = ~v_2737 | v_3748;
assign x_2710 = ~v_2737 | v_149;
assign x_2711 = ~v_2738 | v_3748;
assign x_2712 = ~v_2738 | v_157;
assign x_2713 = ~v_2739 | v_3748;
assign x_2714 = ~v_2739 | v_164;
assign x_2715 = ~v_2740 | v_3748;
assign x_2716 = ~v_2740 | v_170;
assign x_2717 = ~v_2741 | v_3747;
assign x_2718 = ~v_2741 | ~v_3748;
assign x_2719 = ~v_2742 | v_176;
assign x_2720 = ~v_2742 | ~v_3748;
assign x_2721 = ~v_2743 | v_3747;
assign x_2722 = ~v_2743 | v_176;
assign x_2723 = ~v_2744 | v_3746;
assign x_2724 = ~v_2744 | ~v_3747;
assign x_2725 = ~v_2745 | v_177;
assign x_2726 = ~v_2745 | ~v_3747;
assign x_2727 = ~v_2746 | v_3746;
assign x_2728 = ~v_2746 | v_177;
assign x_2729 = ~v_2747 | v_3745;
assign x_2730 = ~v_2747 | ~v_3746;
assign x_2731 = ~v_2748 | v_178;
assign x_2732 = ~v_2748 | ~v_3746;
assign x_2733 = ~v_2749 | v_3745;
assign x_2734 = ~v_2749 | v_178;
assign x_2735 = ~v_2750 | v_180;
assign x_2736 = ~v_2750 | ~v_3745;
assign x_2737 = ~v_2751 | v_179;
assign x_2738 = ~v_2751 | ~v_3745;
assign x_2739 = ~v_2752 | v_180;
assign x_2740 = ~v_2752 | v_179;
assign x_2741 = ~v_2753 | v_3743;
assign x_2742 = ~v_2753 | ~v_3744;
assign x_2743 = ~v_2754 | v_149;
assign x_2744 = ~v_2754 | ~v_3744;
assign x_2745 = ~v_2755 | v_3743;
assign x_2746 = ~v_2755 | v_149;
assign x_2747 = ~v_2756 | v_3742;
assign x_2748 = ~v_2756 | ~v_3743;
assign x_2749 = ~v_2757 | v_157;
assign x_2750 = ~v_2757 | ~v_3743;
assign x_2751 = ~v_2758 | v_3742;
assign x_2752 = ~v_2758 | v_157;
assign x_2753 = ~v_2759 | v_170;
assign x_2754 = ~v_2759 | ~v_3742;
assign x_2755 = ~v_2760 | v_164;
assign x_2756 = ~v_2760 | ~v_3742;
assign x_2757 = ~v_2761 | v_170;
assign x_2758 = ~v_2761 | v_164;
assign x_2759 = ~v_2762 | v_3741;
assign x_2760 = ~v_2762 | v_150;
assign x_2761 = ~v_2763 | v_3741;
assign x_2762 = ~v_2763 | v_158;
assign x_2763 = ~v_2764 | v_3741;
assign x_2764 = ~v_2764 | v_165;
assign x_2765 = ~v_2765 | v_3741;
assign x_2766 = ~v_2765 | v_171;
assign x_2767 = ~v_2766 | v_3741;
assign x_2768 = ~v_2766 | v_176;
assign x_2769 = ~v_2767 | v_3740;
assign x_2770 = ~v_2767 | ~v_3741;
assign x_2771 = ~v_2768 | v_181;
assign x_2772 = ~v_2768 | ~v_3741;
assign x_2773 = ~v_2769 | v_3740;
assign x_2774 = ~v_2769 | v_181;
assign x_2775 = ~v_2770 | v_3739;
assign x_2776 = ~v_2770 | ~v_3740;
assign x_2777 = ~v_2771 | v_182;
assign x_2778 = ~v_2771 | ~v_3740;
assign x_2779 = ~v_2772 | v_3739;
assign x_2780 = ~v_2772 | v_182;
assign x_2781 = ~v_2773 | v_184;
assign x_2782 = ~v_2773 | ~v_3739;
assign x_2783 = ~v_2774 | v_183;
assign x_2784 = ~v_2774 | ~v_3739;
assign x_2785 = ~v_2775 | v_184;
assign x_2786 = ~v_2775 | v_183;
assign x_2787 = ~v_2776 | v_3737;
assign x_2788 = ~v_2776 | ~v_3738;
assign x_2789 = ~v_2777 | v_150;
assign x_2790 = ~v_2777 | ~v_3738;
assign x_2791 = ~v_2778 | v_3737;
assign x_2792 = ~v_2778 | v_150;
assign x_2793 = ~v_2779 | v_3736;
assign x_2794 = ~v_2779 | ~v_3737;
assign x_2795 = ~v_2780 | v_158;
assign x_2796 = ~v_2780 | ~v_3737;
assign x_2797 = ~v_2781 | v_3736;
assign x_2798 = ~v_2781 | v_158;
assign x_2799 = ~v_2782 | v_3735;
assign x_2800 = ~v_2782 | ~v_3736;
assign x_2801 = ~v_2783 | v_165;
assign x_2802 = ~v_2783 | ~v_3736;
assign x_2803 = ~v_2784 | v_3735;
assign x_2804 = ~v_2784 | v_165;
assign x_2805 = ~v_2785 | v_176;
assign x_2806 = ~v_2785 | ~v_3735;
assign x_2807 = ~v_2786 | v_171;
assign x_2808 = ~v_2786 | ~v_3735;
assign x_2809 = ~v_2787 | v_176;
assign x_2810 = ~v_2787 | v_171;
assign x_2811 = ~v_2788 | v_3734;
assign x_2812 = ~v_2788 | v_151;
assign x_2813 = ~v_2789 | v_3734;
assign x_2814 = ~v_2789 | v_159;
assign x_2815 = ~v_2790 | v_3734;
assign x_2816 = ~v_2790 | v_166;
assign x_2817 = ~v_2791 | v_3734;
assign x_2818 = ~v_2791 | v_172;
assign x_2819 = ~v_2792 | v_3734;
assign x_2820 = ~v_2792 | v_177;
assign x_2821 = ~v_2793 | v_3734;
assign x_2822 = ~v_2793 | v_181;
assign x_2823 = ~v_2794 | v_3733;
assign x_2824 = ~v_2794 | ~v_3734;
assign x_2825 = ~v_2795 | v_185;
assign x_2826 = ~v_2795 | ~v_3734;
assign x_2827 = ~v_2796 | v_3733;
assign x_2828 = ~v_2796 | v_185;
assign x_2829 = ~v_2797 | v_187;
assign x_2830 = ~v_2797 | ~v_3733;
assign x_2831 = ~v_2798 | v_186;
assign x_2832 = ~v_2798 | ~v_3733;
assign x_2833 = ~v_2799 | v_187;
assign x_2834 = ~v_2799 | v_186;
assign x_2835 = ~v_2800 | v_3731;
assign x_2836 = ~v_2800 | ~v_3732;
assign x_2837 = ~v_2801 | v_151;
assign x_2838 = ~v_2801 | ~v_3732;
assign x_2839 = ~v_2802 | v_3731;
assign x_2840 = ~v_2802 | v_151;
assign x_2841 = ~v_2803 | v_3730;
assign x_2842 = ~v_2803 | ~v_3731;
assign x_2843 = ~v_2804 | v_159;
assign x_2844 = ~v_2804 | ~v_3731;
assign x_2845 = ~v_2805 | v_3730;
assign x_2846 = ~v_2805 | v_159;
assign x_2847 = ~v_2806 | v_3729;
assign x_2848 = ~v_2806 | ~v_3730;
assign x_2849 = ~v_2807 | v_166;
assign x_2850 = ~v_2807 | ~v_3730;
assign x_2851 = ~v_2808 | v_3729;
assign x_2852 = ~v_2808 | v_166;
assign x_2853 = ~v_2809 | v_3728;
assign x_2854 = ~v_2809 | ~v_3729;
assign x_2855 = ~v_2810 | v_172;
assign x_2856 = ~v_2810 | ~v_3729;
assign x_2857 = ~v_2811 | v_3728;
assign x_2858 = ~v_2811 | v_172;
assign x_2859 = ~v_2812 | v_181;
assign x_2860 = ~v_2812 | ~v_3728;
assign x_2861 = ~v_2813 | v_177;
assign x_2862 = ~v_2813 | ~v_3728;
assign x_2863 = ~v_2814 | v_181;
assign x_2864 = ~v_2814 | v_177;
assign x_2865 = ~v_2815 | v_3727;
assign x_2866 = ~v_2815 | v_152;
assign x_2867 = ~v_2816 | v_3727;
assign x_2868 = ~v_2816 | v_160;
assign x_2869 = ~v_2817 | v_3727;
assign x_2870 = ~v_2817 | v_167;
assign x_2871 = ~v_2818 | v_3727;
assign x_2872 = ~v_2818 | v_173;
assign x_2873 = ~v_2819 | v_3727;
assign x_2874 = ~v_2819 | v_178;
assign x_2875 = ~v_2820 | v_3727;
assign x_2876 = ~v_2820 | v_182;
assign x_2877 = ~v_2821 | v_3727;
assign x_2878 = ~v_2821 | v_185;
assign x_2879 = ~v_2822 | v_189;
assign x_2880 = ~v_2822 | ~v_3727;
assign x_2881 = ~v_2823 | v_188;
assign x_2882 = ~v_2823 | ~v_3727;
assign x_2883 = ~v_2824 | v_189;
assign x_2884 = ~v_2824 | v_188;
assign x_2885 = ~v_2825 | v_3725;
assign x_2886 = ~v_2825 | ~v_3726;
assign x_2887 = ~v_2826 | v_152;
assign x_2888 = ~v_2826 | ~v_3726;
assign x_2889 = ~v_2827 | v_3725;
assign x_2890 = ~v_2827 | v_152;
assign x_2891 = ~v_2828 | v_3724;
assign x_2892 = ~v_2828 | ~v_3725;
assign x_2893 = ~v_2829 | v_160;
assign x_2894 = ~v_2829 | ~v_3725;
assign x_2895 = ~v_2830 | v_3724;
assign x_2896 = ~v_2830 | v_160;
assign x_2897 = ~v_2831 | v_3723;
assign x_2898 = ~v_2831 | ~v_3724;
assign x_2899 = ~v_2832 | v_167;
assign x_2900 = ~v_2832 | ~v_3724;
assign x_2901 = ~v_2833 | v_3723;
assign x_2902 = ~v_2833 | v_167;
assign x_2903 = ~v_2834 | v_3722;
assign x_2904 = ~v_2834 | ~v_3723;
assign x_2905 = ~v_2835 | v_173;
assign x_2906 = ~v_2835 | ~v_3723;
assign x_2907 = ~v_2836 | v_3722;
assign x_2908 = ~v_2836 | v_173;
assign x_2909 = ~v_2837 | v_3721;
assign x_2910 = ~v_2837 | ~v_3722;
assign x_2911 = ~v_2838 | v_178;
assign x_2912 = ~v_2838 | ~v_3722;
assign x_2913 = ~v_2839 | v_3721;
assign x_2914 = ~v_2839 | v_178;
assign x_2915 = ~v_2840 | v_185;
assign x_2916 = ~v_2840 | ~v_3721;
assign x_2917 = ~v_2841 | v_182;
assign x_2918 = ~v_2841 | ~v_3721;
assign x_2919 = ~v_2842 | v_185;
assign x_2920 = ~v_2842 | v_182;
assign x_2921 = ~v_2843 | v_190;
assign x_2922 = ~v_2843 | v_153;
assign x_2923 = ~v_2844 | v_190;
assign x_2924 = ~v_2844 | v_161;
assign x_2925 = ~v_2845 | v_190;
assign x_2926 = ~v_2845 | v_168;
assign x_2927 = ~v_2846 | v_190;
assign x_2928 = ~v_2846 | v_174;
assign x_2929 = ~v_2847 | v_190;
assign x_2930 = ~v_2847 | v_179;
assign x_2931 = ~v_2848 | v_190;
assign x_2932 = ~v_2848 | v_183;
assign x_2933 = ~v_2849 | v_190;
assign x_2934 = ~v_2849 | v_186;
assign x_2935 = ~v_2850 | v_190;
assign x_2936 = ~v_2850 | v_188;
assign x_2937 = ~v_2851 | v_3719;
assign x_2938 = ~v_2851 | ~v_3720;
assign x_2939 = ~v_2852 | v_153;
assign x_2940 = ~v_2852 | ~v_3720;
assign x_2941 = ~v_2853 | v_3719;
assign x_2942 = ~v_2853 | v_153;
assign x_2943 = ~v_2854 | v_3718;
assign x_2944 = ~v_2854 | ~v_3719;
assign x_2945 = ~v_2855 | v_161;
assign x_2946 = ~v_2855 | ~v_3719;
assign x_2947 = ~v_2856 | v_3718;
assign x_2948 = ~v_2856 | v_161;
assign x_2949 = ~v_2857 | v_3717;
assign x_2950 = ~v_2857 | ~v_3718;
assign x_2951 = ~v_2858 | v_168;
assign x_2952 = ~v_2858 | ~v_3718;
assign x_2953 = ~v_2859 | v_3717;
assign x_2954 = ~v_2859 | v_168;
assign x_2955 = ~v_2860 | v_3716;
assign x_2956 = ~v_2860 | ~v_3717;
assign x_2957 = ~v_2861 | v_174;
assign x_2958 = ~v_2861 | ~v_3717;
assign x_2959 = ~v_2862 | v_3716;
assign x_2960 = ~v_2862 | v_174;
assign x_2961 = ~v_2863 | v_3715;
assign x_2962 = ~v_2863 | ~v_3716;
assign x_2963 = ~v_2864 | v_179;
assign x_2964 = ~v_2864 | ~v_3716;
assign x_2965 = ~v_2865 | v_3715;
assign x_2966 = ~v_2865 | v_179;
assign x_2967 = ~v_2866 | v_3714;
assign x_2968 = ~v_2866 | ~v_3715;
assign x_2969 = ~v_2867 | v_183;
assign x_2970 = ~v_2867 | ~v_3715;
assign x_2971 = ~v_2868 | v_3714;
assign x_2972 = ~v_2868 | v_183;
assign x_2973 = ~v_2869 | v_188;
assign x_2974 = ~v_2869 | ~v_3714;
assign x_2975 = ~v_2870 | v_186;
assign x_2976 = ~v_2870 | ~v_3714;
assign x_2977 = ~v_2871 | v_188;
assign x_2978 = ~v_2871 | v_186;
assign x_2979 = ~v_2872 | v_3712;
assign x_2980 = ~v_2872 | ~v_3713;
assign x_2981 = ~v_2873 | v_154;
assign x_2982 = ~v_2873 | ~v_3713;
assign x_2983 = ~v_2874 | v_3712;
assign x_2984 = ~v_2874 | v_154;
assign x_2985 = ~v_2875 | v_3711;
assign x_2986 = ~v_2875 | ~v_3712;
assign x_2987 = ~v_2876 | v_162;
assign x_2988 = ~v_2876 | ~v_3712;
assign x_2989 = ~v_2877 | v_3711;
assign x_2990 = ~v_2877 | v_162;
assign x_2991 = ~v_2878 | v_3710;
assign x_2992 = ~v_2878 | ~v_3711;
assign x_2993 = ~v_2879 | v_169;
assign x_2994 = ~v_2879 | ~v_3711;
assign x_2995 = ~v_2880 | v_3710;
assign x_2996 = ~v_2880 | v_169;
assign x_2997 = ~v_2881 | v_3709;
assign x_2998 = ~v_2881 | ~v_3710;
assign x_2999 = ~v_2882 | v_175;
assign x_3000 = ~v_2882 | ~v_3710;
assign x_3001 = ~v_2883 | v_3709;
assign x_3002 = ~v_2883 | v_175;
assign x_3003 = ~v_2884 | v_3708;
assign x_3004 = ~v_2884 | ~v_3709;
assign x_3005 = ~v_2885 | v_180;
assign x_3006 = ~v_2885 | ~v_3709;
assign x_3007 = ~v_2886 | v_3708;
assign x_3008 = ~v_2886 | v_180;
assign x_3009 = ~v_2887 | v_3707;
assign x_3010 = ~v_2887 | ~v_3708;
assign x_3011 = ~v_2888 | v_184;
assign x_3012 = ~v_2888 | ~v_3708;
assign x_3013 = ~v_2889 | v_3707;
assign x_3014 = ~v_2889 | v_184;
assign x_3015 = ~v_2890 | v_3706;
assign x_3016 = ~v_2890 | ~v_3707;
assign x_3017 = ~v_2891 | v_187;
assign x_3018 = ~v_2891 | ~v_3707;
assign x_3019 = ~v_2892 | v_3706;
assign x_3020 = ~v_2892 | v_187;
assign x_3021 = ~v_2893 | v_190;
assign x_3022 = ~v_2893 | ~v_3706;
assign x_3023 = ~v_2894 | v_189;
assign x_3024 = ~v_2894 | ~v_3706;
assign x_3025 = ~v_2895 | v_190;
assign x_3026 = ~v_2895 | v_189;
assign x_3027 = ~v_2896 | v_3938;
assign x_3028 = ~v_2896 | ~v_3939;
assign x_3029 = ~v_2897 | v_199;
assign x_3030 = ~v_2897 | ~v_3939;
assign x_3031 = ~v_2898 | v_3938;
assign x_3032 = ~v_2898 | v_199;
assign x_3033 = ~v_2899 | v_3937;
assign x_3034 = ~v_2899 | ~v_3938;
assign x_3035 = ~v_2900 | v_198;
assign x_3036 = ~v_2900 | ~v_3938;
assign x_3037 = ~v_2901 | v_3937;
assign x_3038 = ~v_2901 | v_198;
assign x_3039 = ~v_2902 | v_3936;
assign x_3040 = ~v_2902 | ~v_3937;
assign x_3041 = ~v_2903 | v_197;
assign x_3042 = ~v_2903 | ~v_3937;
assign x_3043 = ~v_2904 | v_3936;
assign x_3044 = ~v_2904 | v_197;
assign x_3045 = ~v_2905 | v_3935;
assign x_3046 = ~v_2905 | ~v_3936;
assign x_3047 = ~v_2906 | v_196;
assign x_3048 = ~v_2906 | ~v_3936;
assign x_3049 = ~v_2907 | v_3935;
assign x_3050 = ~v_2907 | v_196;
assign x_3051 = ~v_2908 | v_3934;
assign x_3052 = ~v_2908 | ~v_3935;
assign x_3053 = ~v_2909 | v_195;
assign x_3054 = ~v_2909 | ~v_3935;
assign x_3055 = ~v_2910 | v_3934;
assign x_3056 = ~v_2910 | v_195;
assign x_3057 = ~v_2911 | v_3933;
assign x_3058 = ~v_2911 | ~v_3934;
assign x_3059 = ~v_2912 | v_194;
assign x_3060 = ~v_2912 | ~v_3934;
assign x_3061 = ~v_2913 | v_3933;
assign x_3062 = ~v_2913 | v_194;
assign x_3063 = ~v_2914 | v_3932;
assign x_3064 = ~v_2914 | ~v_3933;
assign x_3065 = ~v_2915 | v_193;
assign x_3066 = ~v_2915 | ~v_3933;
assign x_3067 = ~v_2916 | v_3932;
assign x_3068 = ~v_2916 | v_193;
assign x_3069 = ~v_2917 | v_191;
assign x_3070 = ~v_2917 | ~v_3932;
assign x_3071 = ~v_2918 | v_192;
assign x_3072 = ~v_2918 | ~v_3932;
assign x_3073 = ~v_2919 | v_191;
assign x_3074 = ~v_2919 | v_192;
assign x_3075 = ~v_2920 | v_3930;
assign x_3076 = ~v_2920 | ~v_3931;
assign x_3077 = ~v_2921 | v_207;
assign x_3078 = ~v_2921 | ~v_3931;
assign x_3079 = ~v_2922 | v_3930;
assign x_3080 = ~v_2922 | v_207;
assign x_3081 = ~v_2923 | v_3929;
assign x_3082 = ~v_2923 | ~v_3930;
assign x_3083 = ~v_2924 | v_206;
assign x_3084 = ~v_2924 | ~v_3930;
assign x_3085 = ~v_2925 | v_3929;
assign x_3086 = ~v_2925 | v_206;
assign x_3087 = ~v_2926 | v_3928;
assign x_3088 = ~v_2926 | ~v_3929;
assign x_3089 = ~v_2927 | v_205;
assign x_3090 = ~v_2927 | ~v_3929;
assign x_3091 = ~v_2928 | v_3928;
assign x_3092 = ~v_2928 | v_205;
assign x_3093 = ~v_2929 | v_3927;
assign x_3094 = ~v_2929 | ~v_3928;
assign x_3095 = ~v_2930 | v_204;
assign x_3096 = ~v_2930 | ~v_3928;
assign x_3097 = ~v_2931 | v_3927;
assign x_3098 = ~v_2931 | v_204;
assign x_3099 = ~v_2932 | v_3926;
assign x_3100 = ~v_2932 | ~v_3927;
assign x_3101 = ~v_2933 | v_203;
assign x_3102 = ~v_2933 | ~v_3927;
assign x_3103 = ~v_2934 | v_3926;
assign x_3104 = ~v_2934 | v_203;
assign x_3105 = ~v_2935 | v_3925;
assign x_3106 = ~v_2935 | ~v_3926;
assign x_3107 = ~v_2936 | v_202;
assign x_3108 = ~v_2936 | ~v_3926;
assign x_3109 = ~v_2937 | v_3925;
assign x_3110 = ~v_2937 | v_202;
assign x_3111 = ~v_2938 | v_200;
assign x_3112 = ~v_2938 | ~v_3925;
assign x_3113 = ~v_2939 | v_201;
assign x_3114 = ~v_2939 | ~v_3925;
assign x_3115 = ~v_2940 | v_200;
assign x_3116 = ~v_2940 | v_201;
assign x_3117 = ~v_2941 | v_191;
assign x_3118 = ~v_2941 | v_207;
assign x_3119 = ~v_2942 | v_191;
assign x_3120 = ~v_2942 | v_206;
assign x_3121 = ~v_2943 | v_191;
assign x_3122 = ~v_2943 | v_205;
assign x_3123 = ~v_2944 | v_191;
assign x_3124 = ~v_2944 | v_204;
assign x_3125 = ~v_2945 | v_191;
assign x_3126 = ~v_2945 | v_203;
assign x_3127 = ~v_2946 | v_191;
assign x_3128 = ~v_2946 | v_202;
assign x_3129 = ~v_2947 | v_191;
assign x_3130 = ~v_2947 | v_201;
assign x_3131 = ~v_2948 | v_191;
assign x_3132 = ~v_2948 | v_200;
assign x_3133 = ~v_2949 | v_3923;
assign x_3134 = ~v_2949 | ~v_3924;
assign x_3135 = ~v_2950 | v_214;
assign x_3136 = ~v_2950 | ~v_3924;
assign x_3137 = ~v_2951 | v_3923;
assign x_3138 = ~v_2951 | v_214;
assign x_3139 = ~v_2952 | v_3922;
assign x_3140 = ~v_2952 | ~v_3923;
assign x_3141 = ~v_2953 | v_213;
assign x_3142 = ~v_2953 | ~v_3923;
assign x_3143 = ~v_2954 | v_3922;
assign x_3144 = ~v_2954 | v_213;
assign x_3145 = ~v_2955 | v_3921;
assign x_3146 = ~v_2955 | ~v_3922;
assign x_3147 = ~v_2956 | v_212;
assign x_3148 = ~v_2956 | ~v_3922;
assign x_3149 = ~v_2957 | v_3921;
assign x_3150 = ~v_2957 | v_212;
assign x_3151 = ~v_2958 | v_3920;
assign x_3152 = ~v_2958 | ~v_3921;
assign x_3153 = ~v_2959 | v_211;
assign x_3154 = ~v_2959 | ~v_3921;
assign x_3155 = ~v_2960 | v_3920;
assign x_3156 = ~v_2960 | v_211;
assign x_3157 = ~v_2961 | v_3919;
assign x_3158 = ~v_2961 | ~v_3920;
assign x_3159 = ~v_2962 | v_210;
assign x_3160 = ~v_2962 | ~v_3920;
assign x_3161 = ~v_2963 | v_3919;
assign x_3162 = ~v_2963 | v_210;
assign x_3163 = ~v_2964 | v_208;
assign x_3164 = ~v_2964 | ~v_3919;
assign x_3165 = ~v_2965 | v_209;
assign x_3166 = ~v_2965 | ~v_3919;
assign x_3167 = ~v_2966 | v_208;
assign x_3168 = ~v_2966 | v_209;
assign x_3169 = ~v_2967 | v_3918;
assign x_3170 = ~v_2967 | v_214;
assign x_3171 = ~v_2968 | v_3918;
assign x_3172 = ~v_2968 | v_213;
assign x_3173 = ~v_2969 | v_3918;
assign x_3174 = ~v_2969 | v_212;
assign x_3175 = ~v_2970 | v_3918;
assign x_3176 = ~v_2970 | v_211;
assign x_3177 = ~v_2971 | v_3918;
assign x_3178 = ~v_2971 | v_210;
assign x_3179 = ~v_2972 | v_3918;
assign x_3180 = ~v_2972 | v_209;
assign x_3181 = ~v_2973 | v_3918;
assign x_3182 = ~v_2973 | v_208;
assign x_3183 = ~v_2974 | v_192;
assign x_3184 = ~v_2974 | ~v_3918;
assign x_3185 = ~v_2975 | v_200;
assign x_3186 = ~v_2975 | ~v_3918;
assign x_3187 = ~v_2976 | v_192;
assign x_3188 = ~v_2976 | v_200;
assign x_3189 = ~v_2977 | v_3916;
assign x_3190 = ~v_2977 | ~v_3917;
assign x_3191 = ~v_2978 | v_220;
assign x_3192 = ~v_2978 | ~v_3917;
assign x_3193 = ~v_2979 | v_3916;
assign x_3194 = ~v_2979 | v_220;
assign x_3195 = ~v_2980 | v_3915;
assign x_3196 = ~v_2980 | ~v_3916;
assign x_3197 = ~v_2981 | v_219;
assign x_3198 = ~v_2981 | ~v_3916;
assign x_3199 = ~v_2982 | v_3915;
assign x_3200 = ~v_2982 | v_219;
assign x_3201 = ~v_2983 | v_3914;
assign x_3202 = ~v_2983 | ~v_3915;
assign x_3203 = ~v_2984 | v_218;
assign x_3204 = ~v_2984 | ~v_3915;
assign x_3205 = ~v_2985 | v_3914;
assign x_3206 = ~v_2985 | v_218;
assign x_3207 = ~v_2986 | v_3913;
assign x_3208 = ~v_2986 | ~v_3914;
assign x_3209 = ~v_2987 | v_217;
assign x_3210 = ~v_2987 | ~v_3914;
assign x_3211 = ~v_2988 | v_3913;
assign x_3212 = ~v_2988 | v_217;
assign x_3213 = ~v_2989 | v_215;
assign x_3214 = ~v_2989 | ~v_3913;
assign x_3215 = ~v_2990 | v_216;
assign x_3216 = ~v_2990 | ~v_3913;
assign x_3217 = ~v_2991 | v_215;
assign x_3218 = ~v_2991 | v_216;
assign x_3219 = ~v_2992 | v_3912;
assign x_3220 = ~v_2992 | v_220;
assign x_3221 = ~v_2993 | v_3912;
assign x_3222 = ~v_2993 | v_219;
assign x_3223 = ~v_2994 | v_3912;
assign x_3224 = ~v_2994 | v_218;
assign x_3225 = ~v_2995 | v_3912;
assign x_3226 = ~v_2995 | v_217;
assign x_3227 = ~v_2996 | v_3912;
assign x_3228 = ~v_2996 | v_216;
assign x_3229 = ~v_2997 | v_3912;
assign x_3230 = ~v_2997 | v_215;
assign x_3231 = ~v_2998 | v_3911;
assign x_3232 = ~v_2998 | ~v_3912;
assign x_3233 = ~v_2999 | v_208;
assign x_3234 = ~v_2999 | ~v_3912;
assign x_3235 = ~v_3000 | v_3911;
assign x_3236 = ~v_3000 | v_208;
assign x_3237 = ~v_3001 | v_193;
assign x_3238 = ~v_3001 | ~v_3911;
assign x_3239 = ~v_3002 | v_201;
assign x_3240 = ~v_3002 | ~v_3911;
assign x_3241 = ~v_3003 | v_193;
assign x_3242 = ~v_3003 | v_201;
assign x_3243 = ~v_3004 | v_3909;
assign x_3244 = ~v_3004 | ~v_3910;
assign x_3245 = ~v_3005 | v_225;
assign x_3246 = ~v_3005 | ~v_3910;
assign x_3247 = ~v_3006 | v_3909;
assign x_3248 = ~v_3006 | v_225;
assign x_3249 = ~v_3007 | v_3908;
assign x_3250 = ~v_3007 | ~v_3909;
assign x_3251 = ~v_3008 | v_224;
assign x_3252 = ~v_3008 | ~v_3909;
assign x_3253 = ~v_3009 | v_3908;
assign x_3254 = ~v_3009 | v_224;
assign x_3255 = ~v_3010 | v_3907;
assign x_3256 = ~v_3010 | ~v_3908;
assign x_3257 = ~v_3011 | v_223;
assign x_3258 = ~v_3011 | ~v_3908;
assign x_3259 = ~v_3012 | v_3907;
assign x_3260 = ~v_3012 | v_223;
assign x_3261 = ~v_3013 | v_221;
assign x_3262 = ~v_3013 | ~v_3907;
assign x_3263 = ~v_3014 | v_222;
assign x_3264 = ~v_3014 | ~v_3907;
assign x_3265 = ~v_3015 | v_221;
assign x_3266 = ~v_3015 | v_222;
assign x_3267 = ~v_3016 | v_3906;
assign x_3268 = ~v_3016 | v_225;
assign x_3269 = ~v_3017 | v_3906;
assign x_3270 = ~v_3017 | v_224;
assign x_3271 = ~v_3018 | v_3906;
assign x_3272 = ~v_3018 | v_223;
assign x_3273 = ~v_3019 | v_3906;
assign x_3274 = ~v_3019 | v_222;
assign x_3275 = ~v_3020 | v_3906;
assign x_3276 = ~v_3020 | v_221;
assign x_3277 = ~v_3021 | v_3905;
assign x_3278 = ~v_3021 | ~v_3906;
assign x_3279 = ~v_3022 | v_215;
assign x_3280 = ~v_3022 | ~v_3906;
assign x_3281 = ~v_3023 | v_3905;
assign x_3282 = ~v_3023 | v_215;
assign x_3283 = ~v_3024 | v_3904;
assign x_3284 = ~v_3024 | ~v_3905;
assign x_3285 = ~v_3025 | v_209;
assign x_3286 = ~v_3025 | ~v_3905;
assign x_3287 = ~v_3026 | v_3904;
assign x_3288 = ~v_3026 | v_209;
assign x_3289 = ~v_3027 | v_194;
assign x_3290 = ~v_3027 | ~v_3904;
assign x_3291 = ~v_3028 | v_202;
assign x_3292 = ~v_3028 | ~v_3904;
assign x_3293 = ~v_3029 | v_194;
assign x_3294 = ~v_3029 | v_202;
assign x_3295 = ~v_3030 | v_3902;
assign x_3296 = ~v_3030 | ~v_3903;
assign x_3297 = ~v_3031 | v_229;
assign x_3298 = ~v_3031 | ~v_3903;
assign x_3299 = ~v_3032 | v_3902;
assign x_3300 = ~v_3032 | v_229;
assign x_3301 = ~v_3033 | v_3901;
assign x_3302 = ~v_3033 | ~v_3902;
assign x_3303 = ~v_3034 | v_228;
assign x_3304 = ~v_3034 | ~v_3902;
assign x_3305 = ~v_3035 | v_3901;
assign x_3306 = ~v_3035 | v_228;
assign x_3307 = ~v_3036 | v_226;
assign x_3308 = ~v_3036 | ~v_3901;
assign x_3309 = ~v_3037 | v_227;
assign x_3310 = ~v_3037 | ~v_3901;
assign x_3311 = ~v_3038 | v_226;
assign x_3312 = ~v_3038 | v_227;
assign x_3313 = ~v_3039 | v_3900;
assign x_3314 = ~v_3039 | v_229;
assign x_3315 = ~v_3040 | v_3900;
assign x_3316 = ~v_3040 | v_228;
assign x_3317 = ~v_3041 | v_3900;
assign x_3318 = ~v_3041 | v_227;
assign x_3319 = ~v_3042 | v_3900;
assign x_3320 = ~v_3042 | v_226;
assign x_3321 = ~v_3043 | v_3899;
assign x_3322 = ~v_3043 | ~v_3900;
assign x_3323 = ~v_3044 | v_221;
assign x_3324 = ~v_3044 | ~v_3900;
assign x_3325 = ~v_3045 | v_3899;
assign x_3326 = ~v_3045 | v_221;
assign x_3327 = ~v_3046 | v_3898;
assign x_3328 = ~v_3046 | ~v_3899;
assign x_3329 = ~v_3047 | v_216;
assign x_3330 = ~v_3047 | ~v_3899;
assign x_3331 = ~v_3048 | v_3898;
assign x_3332 = ~v_3048 | v_216;
assign x_3333 = ~v_3049 | v_3897;
assign x_3334 = ~v_3049 | ~v_3898;
assign x_3335 = ~v_3050 | v_210;
assign x_3336 = ~v_3050 | ~v_3898;
assign x_3337 = ~v_3051 | v_3897;
assign x_3338 = ~v_3051 | v_210;
assign x_3339 = ~v_3052 | v_195;
assign x_3340 = ~v_3052 | ~v_3897;
assign x_3341 = ~v_3053 | v_203;
assign x_3342 = ~v_3053 | ~v_3897;
assign x_3343 = ~v_3054 | v_195;
assign x_3344 = ~v_3054 | v_203;
assign x_3345 = ~v_3055 | v_3895;
assign x_3346 = ~v_3055 | ~v_3896;
assign x_3347 = ~v_3056 | v_232;
assign x_3348 = ~v_3056 | ~v_3896;
assign x_3349 = ~v_3057 | v_3895;
assign x_3350 = ~v_3057 | v_232;
assign x_3351 = ~v_3058 | v_230;
assign x_3352 = ~v_3058 | ~v_3895;
assign x_3353 = ~v_3059 | v_231;
assign x_3354 = ~v_3059 | ~v_3895;
assign x_3355 = ~v_3060 | v_230;
assign x_3356 = ~v_3060 | v_231;
assign x_3357 = ~v_3061 | v_3894;
assign x_3358 = ~v_3061 | v_232;
assign x_3359 = ~v_3062 | v_3894;
assign x_3360 = ~v_3062 | v_231;
assign x_3361 = ~v_3063 | v_3894;
assign x_3362 = ~v_3063 | v_230;
assign x_3363 = ~v_3064 | v_3893;
assign x_3364 = ~v_3064 | ~v_3894;
assign x_3365 = ~v_3065 | v_226;
assign x_3366 = ~v_3065 | ~v_3894;
assign x_3367 = ~v_3066 | v_3893;
assign x_3368 = ~v_3066 | v_226;
assign x_3369 = ~v_3067 | v_3892;
assign x_3370 = ~v_3067 | ~v_3893;
assign x_3371 = ~v_3068 | v_222;
assign x_3372 = ~v_3068 | ~v_3893;
assign x_3373 = ~v_3069 | v_3892;
assign x_3374 = ~v_3069 | v_222;
assign x_3375 = ~v_3070 | v_3891;
assign x_3376 = ~v_3070 | ~v_3892;
assign x_3377 = ~v_3071 | v_217;
assign x_3378 = ~v_3071 | ~v_3892;
assign x_3379 = ~v_3072 | v_3891;
assign x_3380 = ~v_3072 | v_217;
assign x_3381 = ~v_3073 | v_3890;
assign x_3382 = ~v_3073 | ~v_3891;
assign x_3383 = ~v_3074 | v_211;
assign x_3384 = ~v_3074 | ~v_3891;
assign x_3385 = ~v_3075 | v_3890;
assign x_3386 = ~v_3075 | v_211;
assign x_3387 = ~v_3076 | v_196;
assign x_3388 = ~v_3076 | ~v_3890;
assign x_3389 = ~v_3077 | v_204;
assign x_3390 = ~v_3077 | ~v_3890;
assign x_3391 = ~v_3078 | v_196;
assign x_3392 = ~v_3078 | v_204;
assign x_3393 = ~v_3079 | v_233;
assign x_3394 = ~v_3079 | ~v_3889;
assign x_3395 = ~v_3080 | v_234;
assign x_3396 = ~v_3080 | ~v_3889;
assign x_3397 = ~v_3081 | v_233;
assign x_3398 = ~v_3081 | v_234;
assign x_3399 = ~v_3082 | v_3888;
assign x_3400 = ~v_3082 | v_234;
assign x_3401 = ~v_3083 | v_3888;
assign x_3402 = ~v_3083 | v_233;
assign x_3403 = ~v_3084 | v_3887;
assign x_3404 = ~v_3084 | ~v_3888;
assign x_3405 = ~v_3085 | v_230;
assign x_3406 = ~v_3085 | ~v_3888;
assign x_3407 = ~v_3086 | v_3887;
assign x_3408 = ~v_3086 | v_230;
assign x_3409 = ~v_3087 | v_3886;
assign x_3410 = ~v_3087 | ~v_3887;
assign x_3411 = ~v_3088 | v_227;
assign x_3412 = ~v_3088 | ~v_3887;
assign x_3413 = ~v_3089 | v_3886;
assign x_3414 = ~v_3089 | v_227;
assign x_3415 = ~v_3090 | v_3885;
assign x_3416 = ~v_3090 | ~v_3886;
assign x_3417 = ~v_3091 | v_223;
assign x_3418 = ~v_3091 | ~v_3886;
assign x_3419 = ~v_3092 | v_3885;
assign x_3420 = ~v_3092 | v_223;
assign x_3421 = ~v_3093 | v_3884;
assign x_3422 = ~v_3093 | ~v_3885;
assign x_3423 = ~v_3094 | v_218;
assign x_3424 = ~v_3094 | ~v_3885;
assign x_3425 = ~v_3095 | v_3884;
assign x_3426 = ~v_3095 | v_218;
assign x_3427 = ~v_3096 | v_3883;
assign x_3428 = ~v_3096 | ~v_3884;
assign x_3429 = ~v_3097 | v_212;
assign x_3430 = ~v_3097 | ~v_3884;
assign x_3431 = ~v_3098 | v_3883;
assign x_3432 = ~v_3098 | v_212;
assign x_3433 = ~v_3099 | v_197;
assign x_3434 = ~v_3099 | ~v_3883;
assign x_3435 = ~v_3100 | v_205;
assign x_3436 = ~v_3100 | ~v_3883;
assign x_3437 = ~v_3101 | v_197;
assign x_3438 = ~v_3101 | v_205;
assign x_3439 = ~v_3102 | v_3882;
assign x_3440 = ~v_3102 | v_235;
assign x_3441 = ~v_3103 | v_3881;
assign x_3442 = ~v_3103 | ~v_3882;
assign x_3443 = ~v_3104 | v_233;
assign x_3444 = ~v_3104 | ~v_3882;
assign x_3445 = ~v_3105 | v_3881;
assign x_3446 = ~v_3105 | v_233;
assign x_3447 = ~v_3106 | v_3880;
assign x_3448 = ~v_3106 | ~v_3881;
assign x_3449 = ~v_3107 | v_231;
assign x_3450 = ~v_3107 | ~v_3881;
assign x_3451 = ~v_3108 | v_3880;
assign x_3452 = ~v_3108 | v_231;
assign x_3453 = ~v_3109 | v_3879;
assign x_3454 = ~v_3109 | ~v_3880;
assign x_3455 = ~v_3110 | v_228;
assign x_3456 = ~v_3110 | ~v_3880;
assign x_3457 = ~v_3111 | v_3879;
assign x_3458 = ~v_3111 | v_228;
assign x_3459 = ~v_3112 | v_3878;
assign x_3460 = ~v_3112 | ~v_3879;
assign x_3461 = ~v_3113 | v_224;
assign x_3462 = ~v_3113 | ~v_3879;
assign x_3463 = ~v_3114 | v_3878;
assign x_3464 = ~v_3114 | v_224;
assign x_3465 = ~v_3115 | v_3877;
assign x_3466 = ~v_3115 | ~v_3878;
assign x_3467 = ~v_3116 | v_219;
assign x_3468 = ~v_3116 | ~v_3878;
assign x_3469 = ~v_3117 | v_3877;
assign x_3470 = ~v_3117 | v_219;
assign x_3471 = ~v_3118 | v_3876;
assign x_3472 = ~v_3118 | ~v_3877;
assign x_3473 = ~v_3119 | v_213;
assign x_3474 = ~v_3119 | ~v_3877;
assign x_3475 = ~v_3120 | v_3876;
assign x_3476 = ~v_3120 | v_213;
assign x_3477 = ~v_3121 | v_198;
assign x_3478 = ~v_3121 | ~v_3876;
assign x_3479 = ~v_3122 | v_206;
assign x_3480 = ~v_3122 | ~v_3876;
assign x_3481 = ~v_3123 | v_198;
assign x_3482 = ~v_3123 | v_206;
assign x_3483 = ~v_3124 | v_3874;
assign x_3484 = ~v_3124 | ~v_3875;
assign x_3485 = ~v_3125 | v_235;
assign x_3486 = ~v_3125 | ~v_3875;
assign x_3487 = ~v_3126 | v_3874;
assign x_3488 = ~v_3126 | v_235;
assign x_3489 = ~v_3127 | v_3873;
assign x_3490 = ~v_3127 | ~v_3874;
assign x_3491 = ~v_3128 | v_234;
assign x_3492 = ~v_3128 | ~v_3874;
assign x_3493 = ~v_3129 | v_3873;
assign x_3494 = ~v_3129 | v_234;
assign x_3495 = ~v_3130 | v_3872;
assign x_3496 = ~v_3130 | ~v_3873;
assign x_3497 = ~v_3131 | v_232;
assign x_3498 = ~v_3131 | ~v_3873;
assign x_3499 = ~v_3132 | v_3872;
assign x_3500 = ~v_3132 | v_232;
assign x_3501 = ~v_3133 | v_3871;
assign x_3502 = ~v_3133 | ~v_3872;
assign x_3503 = ~v_3134 | v_229;
assign x_3504 = ~v_3134 | ~v_3872;
assign x_3505 = ~v_3135 | v_3871;
assign x_3506 = ~v_3135 | v_229;
assign x_3507 = ~v_3136 | v_3870;
assign x_3508 = ~v_3136 | ~v_3871;
assign x_3509 = ~v_3137 | v_225;
assign x_3510 = ~v_3137 | ~v_3871;
assign x_3511 = ~v_3138 | v_3870;
assign x_3512 = ~v_3138 | v_225;
assign x_3513 = ~v_3139 | v_3869;
assign x_3514 = ~v_3139 | ~v_3870;
assign x_3515 = ~v_3140 | v_220;
assign x_3516 = ~v_3140 | ~v_3870;
assign x_3517 = ~v_3141 | v_3869;
assign x_3518 = ~v_3141 | v_220;
assign x_3519 = ~v_3142 | v_3868;
assign x_3520 = ~v_3142 | ~v_3869;
assign x_3521 = ~v_3143 | v_214;
assign x_3522 = ~v_3143 | ~v_3869;
assign x_3523 = ~v_3144 | v_3868;
assign x_3524 = ~v_3144 | v_214;
assign x_3525 = ~v_3145 | v_199;
assign x_3526 = ~v_3145 | ~v_3868;
assign x_3527 = ~v_3146 | v_207;
assign x_3528 = ~v_3146 | ~v_3868;
assign x_3529 = ~v_3147 | v_199;
assign x_3530 = ~v_3147 | v_207;
assign x_3531 = ~v_3148 | v_4010;
assign x_3532 = ~v_3148 | ~v_4011;
assign x_3533 = ~v_3149 | v_191;
assign x_3534 = ~v_3149 | ~v_4011;
assign x_3535 = ~v_3150 | v_4010;
assign x_3536 = ~v_3150 | v_191;
assign x_3537 = ~v_3151 | v_4009;
assign x_3538 = ~v_3151 | ~v_4010;
assign x_3539 = ~v_3152 | v_192;
assign x_3540 = ~v_3152 | ~v_4010;
assign x_3541 = ~v_3153 | v_4009;
assign x_3542 = ~v_3153 | v_192;
assign x_3543 = ~v_3154 | v_4008;
assign x_3544 = ~v_3154 | ~v_4009;
assign x_3545 = ~v_3155 | v_193;
assign x_3546 = ~v_3155 | ~v_4009;
assign x_3547 = ~v_3156 | v_4008;
assign x_3548 = ~v_3156 | v_193;
assign x_3549 = ~v_3157 | v_4007;
assign x_3550 = ~v_3157 | ~v_4008;
assign x_3551 = ~v_3158 | v_194;
assign x_3552 = ~v_3158 | ~v_4008;
assign x_3553 = ~v_3159 | v_4007;
assign x_3554 = ~v_3159 | v_194;
assign x_3555 = ~v_3160 | v_4006;
assign x_3556 = ~v_3160 | ~v_4007;
assign x_3557 = ~v_3161 | v_195;
assign x_3558 = ~v_3161 | ~v_4007;
assign x_3559 = ~v_3162 | v_4006;
assign x_3560 = ~v_3162 | v_195;
assign x_3561 = ~v_3163 | v_4005;
assign x_3562 = ~v_3163 | ~v_4006;
assign x_3563 = ~v_3164 | v_196;
assign x_3564 = ~v_3164 | ~v_4006;
assign x_3565 = ~v_3165 | v_4005;
assign x_3566 = ~v_3165 | v_196;
assign x_3567 = ~v_3166 | v_4004;
assign x_3568 = ~v_3166 | ~v_4005;
assign x_3569 = ~v_3167 | v_197;
assign x_3570 = ~v_3167 | ~v_4005;
assign x_3571 = ~v_3168 | v_4004;
assign x_3572 = ~v_3168 | v_197;
assign x_3573 = ~v_3169 | v_199;
assign x_3574 = ~v_3169 | ~v_4004;
assign x_3575 = ~v_3170 | v_198;
assign x_3576 = ~v_3170 | ~v_4004;
assign x_3577 = ~v_3171 | v_199;
assign x_3578 = ~v_3171 | v_198;
assign x_3579 = ~v_3172 | v_4003;
assign x_3580 = ~v_3172 | v_191;
assign x_3581 = ~v_3173 | v_4002;
assign x_3582 = ~v_3173 | ~v_4003;
assign x_3583 = ~v_3174 | v_200;
assign x_3584 = ~v_3174 | ~v_4003;
assign x_3585 = ~v_3175 | v_4002;
assign x_3586 = ~v_3175 | v_200;
assign x_3587 = ~v_3176 | v_4001;
assign x_3588 = ~v_3176 | ~v_4002;
assign x_3589 = ~v_3177 | v_201;
assign x_3590 = ~v_3177 | ~v_4002;
assign x_3591 = ~v_3178 | v_4001;
assign x_3592 = ~v_3178 | v_201;
assign x_3593 = ~v_3179 | v_4000;
assign x_3594 = ~v_3179 | ~v_4001;
assign x_3595 = ~v_3180 | v_202;
assign x_3596 = ~v_3180 | ~v_4001;
assign x_3597 = ~v_3181 | v_4000;
assign x_3598 = ~v_3181 | v_202;
assign x_3599 = ~v_3182 | v_3999;
assign x_3600 = ~v_3182 | ~v_4000;
assign x_3601 = ~v_3183 | v_203;
assign x_3602 = ~v_3183 | ~v_4000;
assign x_3603 = ~v_3184 | v_3999;
assign x_3604 = ~v_3184 | v_203;
assign x_3605 = ~v_3185 | v_3998;
assign x_3606 = ~v_3185 | ~v_3999;
assign x_3607 = ~v_3186 | v_204;
assign x_3608 = ~v_3186 | ~v_3999;
assign x_3609 = ~v_3187 | v_3998;
assign x_3610 = ~v_3187 | v_204;
assign x_3611 = ~v_3188 | v_3997;
assign x_3612 = ~v_3188 | ~v_3998;
assign x_3613 = ~v_3189 | v_205;
assign x_3614 = ~v_3189 | ~v_3998;
assign x_3615 = ~v_3190 | v_3997;
assign x_3616 = ~v_3190 | v_205;
assign x_3617 = ~v_3191 | v_207;
assign x_3618 = ~v_3191 | ~v_3997;
assign x_3619 = ~v_3192 | v_206;
assign x_3620 = ~v_3192 | ~v_3997;
assign x_3621 = ~v_3193 | v_207;
assign x_3622 = ~v_3193 | v_206;
assign x_3623 = ~v_3194 | v_3996;
assign x_3624 = ~v_3194 | v_192;
assign x_3625 = ~v_3195 | v_3996;
assign x_3626 = ~v_3195 | v_200;
assign x_3627 = ~v_3196 | v_3995;
assign x_3628 = ~v_3196 | ~v_3996;
assign x_3629 = ~v_3197 | v_208;
assign x_3630 = ~v_3197 | ~v_3996;
assign x_3631 = ~v_3198 | v_3995;
assign x_3632 = ~v_3198 | v_208;
assign x_3633 = ~v_3199 | v_3994;
assign x_3634 = ~v_3199 | ~v_3995;
assign x_3635 = ~v_3200 | v_209;
assign x_3636 = ~v_3200 | ~v_3995;
assign x_3637 = ~v_3201 | v_3994;
assign x_3638 = ~v_3201 | v_209;
assign x_3639 = ~v_3202 | v_3993;
assign x_3640 = ~v_3202 | ~v_3994;
assign x_3641 = ~v_3203 | v_210;
assign x_3642 = ~v_3203 | ~v_3994;
assign x_3643 = ~v_3204 | v_3993;
assign x_3644 = ~v_3204 | v_210;
assign x_3645 = ~v_3205 | v_3992;
assign x_3646 = ~v_3205 | ~v_3993;
assign x_3647 = ~v_3206 | v_211;
assign x_3648 = ~v_3206 | ~v_3993;
assign x_3649 = ~v_3207 | v_3992;
assign x_3650 = ~v_3207 | v_211;
assign x_3651 = ~v_3208 | v_3991;
assign x_3652 = ~v_3208 | ~v_3992;
assign x_3653 = ~v_3209 | v_212;
assign x_3654 = ~v_3209 | ~v_3992;
assign x_3655 = ~v_3210 | v_3991;
assign x_3656 = ~v_3210 | v_212;
assign x_3657 = ~v_3211 | v_214;
assign x_3658 = ~v_3211 | ~v_3991;
assign x_3659 = ~v_3212 | v_213;
assign x_3660 = ~v_3212 | ~v_3991;
assign x_3661 = ~v_3213 | v_214;
assign x_3662 = ~v_3213 | v_213;
assign x_3663 = ~v_3214 | v_200;
assign x_3664 = ~v_3214 | ~v_3990;
assign x_3665 = ~v_3215 | v_192;
assign x_3666 = ~v_3215 | ~v_3990;
assign x_3667 = ~v_3216 | v_200;
assign x_3668 = ~v_3216 | v_192;
assign x_3669 = ~v_3217 | v_3989;
assign x_3670 = ~v_3217 | v_193;
assign x_3671 = ~v_3218 | v_3989;
assign x_3672 = ~v_3218 | v_201;
assign x_3673 = ~v_3219 | v_3989;
assign x_3674 = ~v_3219 | v_208;
assign x_3675 = ~v_3220 | v_3988;
assign x_3676 = ~v_3220 | ~v_3989;
assign x_3677 = ~v_3221 | v_215;
assign x_3678 = ~v_3221 | ~v_3989;
assign x_3679 = ~v_3222 | v_3988;
assign x_3680 = ~v_3222 | v_215;
assign x_3681 = ~v_3223 | v_3987;
assign x_3682 = ~v_3223 | ~v_3988;
assign x_3683 = ~v_3224 | v_216;
assign x_3684 = ~v_3224 | ~v_3988;
assign x_3685 = ~v_3225 | v_3987;
assign x_3686 = ~v_3225 | v_216;
assign x_3687 = ~v_3226 | v_3986;
assign x_3688 = ~v_3226 | ~v_3987;
assign x_3689 = ~v_3227 | v_217;
assign x_3690 = ~v_3227 | ~v_3987;
assign x_3691 = ~v_3228 | v_3986;
assign x_3692 = ~v_3228 | v_217;
assign x_3693 = ~v_3229 | v_3985;
assign x_3694 = ~v_3229 | ~v_3986;
assign x_3695 = ~v_3230 | v_218;
assign x_3696 = ~v_3230 | ~v_3986;
assign x_3697 = ~v_3231 | v_3985;
assign x_3698 = ~v_3231 | v_218;
assign x_3699 = ~v_3232 | v_220;
assign x_3700 = ~v_3232 | ~v_3985;
assign x_3701 = ~v_3233 | v_219;
assign x_3702 = ~v_3233 | ~v_3985;
assign x_3703 = ~v_3234 | v_220;
assign x_3704 = ~v_3234 | v_219;
assign x_3705 = ~v_3235 | v_3983;
assign x_3706 = ~v_3235 | ~v_3984;
assign x_3707 = ~v_3236 | v_193;
assign x_3708 = ~v_3236 | ~v_3984;
assign x_3709 = ~v_3237 | v_3983;
assign x_3710 = ~v_3237 | v_193;
assign x_3711 = ~v_3238 | v_208;
assign x_3712 = ~v_3238 | ~v_3983;
assign x_3713 = ~v_3239 | v_201;
assign x_3714 = ~v_3239 | ~v_3983;
assign x_3715 = ~v_3240 | v_208;
assign x_3716 = ~v_3240 | v_201;
assign x_3717 = ~v_3241 | v_3982;
assign x_3718 = ~v_3241 | v_194;
assign x_3719 = ~v_3242 | v_3982;
assign x_3720 = ~v_3242 | v_202;
assign x_3721 = ~v_3243 | v_3982;
assign x_3722 = ~v_3243 | v_209;
assign x_3723 = ~v_3244 | v_3982;
assign x_3724 = ~v_3244 | v_215;
assign x_3725 = ~v_3245 | v_3981;
assign x_3726 = ~v_3245 | ~v_3982;
assign x_3727 = ~v_3246 | v_221;
assign x_3728 = ~v_3246 | ~v_3982;
assign x_3729 = ~v_3247 | v_3981;
assign x_3730 = ~v_3247 | v_221;
assign x_3731 = ~v_3248 | v_3980;
assign x_3732 = ~v_3248 | ~v_3981;
assign x_3733 = ~v_3249 | v_222;
assign x_3734 = ~v_3249 | ~v_3981;
assign x_3735 = ~v_3250 | v_3980;
assign x_3736 = ~v_3250 | v_222;
assign x_3737 = ~v_3251 | v_3979;
assign x_3738 = ~v_3251 | ~v_3980;
assign x_3739 = ~v_3252 | v_223;
assign x_3740 = ~v_3252 | ~v_3980;
assign x_3741 = ~v_3253 | v_3979;
assign x_3742 = ~v_3253 | v_223;
assign x_3743 = ~v_3254 | v_225;
assign x_3744 = ~v_3254 | ~v_3979;
assign x_3745 = ~v_3255 | v_224;
assign x_3746 = ~v_3255 | ~v_3979;
assign x_3747 = ~v_3256 | v_225;
assign x_3748 = ~v_3256 | v_224;
assign x_3749 = ~v_3257 | v_3977;
assign x_3750 = ~v_3257 | ~v_3978;
assign x_3751 = ~v_3258 | v_194;
assign x_3752 = ~v_3258 | ~v_3978;
assign x_3753 = ~v_3259 | v_3977;
assign x_3754 = ~v_3259 | v_194;
assign x_3755 = ~v_3260 | v_3976;
assign x_3756 = ~v_3260 | ~v_3977;
assign x_3757 = ~v_3261 | v_202;
assign x_3758 = ~v_3261 | ~v_3977;
assign x_3759 = ~v_3262 | v_3976;
assign x_3760 = ~v_3262 | v_202;
assign x_3761 = ~v_3263 | v_215;
assign x_3762 = ~v_3263 | ~v_3976;
assign x_3763 = ~v_3264 | v_209;
assign x_3764 = ~v_3264 | ~v_3976;
assign x_3765 = ~v_3265 | v_215;
assign x_3766 = ~v_3265 | v_209;
assign x_3767 = ~v_3266 | v_3975;
assign x_3768 = ~v_3266 | v_195;
assign x_3769 = ~v_3267 | v_3975;
assign x_3770 = ~v_3267 | v_203;
assign x_3771 = ~v_3268 | v_3975;
assign x_3772 = ~v_3268 | v_210;
assign x_3773 = ~v_3269 | v_3975;
assign x_3774 = ~v_3269 | v_216;
assign x_3775 = ~v_3270 | v_3975;
assign x_3776 = ~v_3270 | v_221;
assign x_3777 = ~v_3271 | v_3974;
assign x_3778 = ~v_3271 | ~v_3975;
assign x_3779 = ~v_3272 | v_226;
assign x_3780 = ~v_3272 | ~v_3975;
assign x_3781 = ~v_3273 | v_3974;
assign x_3782 = ~v_3273 | v_226;
assign x_3783 = ~v_3274 | v_3973;
assign x_3784 = ~v_3274 | ~v_3974;
assign x_3785 = ~v_3275 | v_227;
assign x_3786 = ~v_3275 | ~v_3974;
assign x_3787 = ~v_3276 | v_3973;
assign x_3788 = ~v_3276 | v_227;
assign x_3789 = ~v_3277 | v_229;
assign x_3790 = ~v_3277 | ~v_3973;
assign x_3791 = ~v_3278 | v_228;
assign x_3792 = ~v_3278 | ~v_3973;
assign x_3793 = ~v_3279 | v_229;
assign x_3794 = ~v_3279 | v_228;
assign x_3795 = ~v_3280 | v_3971;
assign x_3796 = ~v_3280 | ~v_3972;
assign x_3797 = ~v_3281 | v_195;
assign x_3798 = ~v_3281 | ~v_3972;
assign x_3799 = ~v_3282 | v_3971;
assign x_3800 = ~v_3282 | v_195;
assign x_3801 = ~v_3283 | v_3970;
assign x_3802 = ~v_3283 | ~v_3971;
assign x_3803 = ~v_3284 | v_203;
assign x_3804 = ~v_3284 | ~v_3971;
assign x_3805 = ~v_3285 | v_3970;
assign x_3806 = ~v_3285 | v_203;
assign x_3807 = ~v_3286 | v_3969;
assign x_3808 = ~v_3286 | ~v_3970;
assign x_3809 = ~v_3287 | v_210;
assign x_3810 = ~v_3287 | ~v_3970;
assign x_3811 = ~v_3288 | v_3969;
assign x_3812 = ~v_3288 | v_210;
assign x_3813 = ~v_3289 | v_221;
assign x_3814 = ~v_3289 | ~v_3969;
assign x_3815 = ~v_3290 | v_216;
assign x_3816 = ~v_3290 | ~v_3969;
assign x_3817 = ~v_3291 | v_221;
assign x_3818 = ~v_3291 | v_216;
assign x_3819 = ~v_3292 | v_3968;
assign x_3820 = ~v_3292 | v_196;
assign x_3821 = ~v_3293 | v_3968;
assign x_3822 = ~v_3293 | v_204;
assign x_3823 = ~v_3294 | v_3968;
assign x_3824 = ~v_3294 | v_211;
assign x_3825 = ~v_3295 | v_3968;
assign x_3826 = ~v_3295 | v_217;
assign x_3827 = ~v_3296 | v_3968;
assign x_3828 = ~v_3296 | v_222;
assign x_3829 = ~v_3297 | v_3968;
assign x_3830 = ~v_3297 | v_226;
assign x_3831 = ~v_3298 | v_3967;
assign x_3832 = ~v_3298 | ~v_3968;
assign x_3833 = ~v_3299 | v_230;
assign x_3834 = ~v_3299 | ~v_3968;
assign x_3835 = ~v_3300 | v_3967;
assign x_3836 = ~v_3300 | v_230;
assign x_3837 = ~v_3301 | v_232;
assign x_3838 = ~v_3301 | ~v_3967;
assign x_3839 = ~v_3302 | v_231;
assign x_3840 = ~v_3302 | ~v_3967;
assign x_3841 = ~v_3303 | v_232;
assign x_3842 = ~v_3303 | v_231;
assign x_3843 = ~v_3304 | v_3965;
assign x_3844 = ~v_3304 | ~v_3966;
assign x_3845 = ~v_3305 | v_196;
assign x_3846 = ~v_3305 | ~v_3966;
assign x_3847 = ~v_3306 | v_3965;
assign x_3848 = ~v_3306 | v_196;
assign x_3849 = ~v_3307 | v_3964;
assign x_3850 = ~v_3307 | ~v_3965;
assign x_3851 = ~v_3308 | v_204;
assign x_3852 = ~v_3308 | ~v_3965;
assign x_3853 = ~v_3309 | v_3964;
assign x_3854 = ~v_3309 | v_204;
assign x_3855 = ~v_3310 | v_3963;
assign x_3856 = ~v_3310 | ~v_3964;
assign x_3857 = ~v_3311 | v_211;
assign x_3858 = ~v_3311 | ~v_3964;
assign x_3859 = ~v_3312 | v_3963;
assign x_3860 = ~v_3312 | v_211;
assign x_3861 = ~v_3313 | v_3962;
assign x_3862 = ~v_3313 | ~v_3963;
assign x_3863 = ~v_3314 | v_217;
assign x_3864 = ~v_3314 | ~v_3963;
assign x_3865 = ~v_3315 | v_3962;
assign x_3866 = ~v_3315 | v_217;
assign x_3867 = ~v_3316 | v_226;
assign x_3868 = ~v_3316 | ~v_3962;
assign x_3869 = ~v_3317 | v_222;
assign x_3870 = ~v_3317 | ~v_3962;
assign x_3871 = ~v_3318 | v_226;
assign x_3872 = ~v_3318 | v_222;
assign x_3873 = ~v_3319 | v_3961;
assign x_3874 = ~v_3319 | v_197;
assign x_3875 = ~v_3320 | v_3961;
assign x_3876 = ~v_3320 | v_205;
assign x_3877 = ~v_3321 | v_3961;
assign x_3878 = ~v_3321 | v_212;
assign x_3879 = ~v_3322 | v_3961;
assign x_3880 = ~v_3322 | v_218;
assign x_3881 = ~v_3323 | v_3961;
assign x_3882 = ~v_3323 | v_223;
assign x_3883 = ~v_3324 | v_3961;
assign x_3884 = ~v_3324 | v_227;
assign x_3885 = ~v_3325 | v_3961;
assign x_3886 = ~v_3325 | v_230;
assign x_3887 = ~v_3326 | v_234;
assign x_3888 = ~v_3326 | ~v_3961;
assign x_3889 = ~v_3327 | v_233;
assign x_3890 = ~v_3327 | ~v_3961;
assign x_3891 = ~v_3328 | v_234;
assign x_3892 = ~v_3328 | v_233;
assign x_3893 = ~v_3329 | v_3959;
assign x_3894 = ~v_3329 | ~v_3960;
assign x_3895 = ~v_3330 | v_197;
assign x_3896 = ~v_3330 | ~v_3960;
assign x_3897 = ~v_3331 | v_3959;
assign x_3898 = ~v_3331 | v_197;
assign x_3899 = ~v_3332 | v_3958;
assign x_3900 = ~v_3332 | ~v_3959;
assign x_3901 = ~v_3333 | v_205;
assign x_3902 = ~v_3333 | ~v_3959;
assign x_3903 = ~v_3334 | v_3958;
assign x_3904 = ~v_3334 | v_205;
assign x_3905 = ~v_3335 | v_3957;
assign x_3906 = ~v_3335 | ~v_3958;
assign x_3907 = ~v_3336 | v_212;
assign x_3908 = ~v_3336 | ~v_3958;
assign x_3909 = ~v_3337 | v_3957;
assign x_3910 = ~v_3337 | v_212;
assign x_3911 = ~v_3338 | v_3956;
assign x_3912 = ~v_3338 | ~v_3957;
assign x_3913 = ~v_3339 | v_218;
assign x_3914 = ~v_3339 | ~v_3957;
assign x_3915 = ~v_3340 | v_3956;
assign x_3916 = ~v_3340 | v_218;
assign x_3917 = ~v_3341 | v_3955;
assign x_3918 = ~v_3341 | ~v_3956;
assign x_3919 = ~v_3342 | v_223;
assign x_3920 = ~v_3342 | ~v_3956;
assign x_3921 = ~v_3343 | v_3955;
assign x_3922 = ~v_3343 | v_223;
assign x_3923 = ~v_3344 | v_230;
assign x_3924 = ~v_3344 | ~v_3955;
assign x_3925 = ~v_3345 | v_227;
assign x_3926 = ~v_3345 | ~v_3955;
assign x_3927 = ~v_3346 | v_230;
assign x_3928 = ~v_3346 | v_227;
assign x_3929 = ~v_3347 | v_235;
assign x_3930 = ~v_3347 | v_198;
assign x_3931 = ~v_3348 | v_235;
assign x_3932 = ~v_3348 | v_206;
assign x_3933 = ~v_3349 | v_235;
assign x_3934 = ~v_3349 | v_213;
assign x_3935 = ~v_3350 | v_235;
assign x_3936 = ~v_3350 | v_219;
assign x_3937 = ~v_3351 | v_235;
assign x_3938 = ~v_3351 | v_224;
assign x_3939 = ~v_3352 | v_235;
assign x_3940 = ~v_3352 | v_228;
assign x_3941 = ~v_3353 | v_235;
assign x_3942 = ~v_3353 | v_231;
assign x_3943 = ~v_3354 | v_235;
assign x_3944 = ~v_3354 | v_233;
assign x_3945 = ~v_3355 | v_3953;
assign x_3946 = ~v_3355 | ~v_3954;
assign x_3947 = ~v_3356 | v_198;
assign x_3948 = ~v_3356 | ~v_3954;
assign x_3949 = ~v_3357 | v_3953;
assign x_3950 = ~v_3357 | v_198;
assign x_3951 = ~v_3358 | v_3952;
assign x_3952 = ~v_3358 | ~v_3953;
assign x_3953 = ~v_3359 | v_206;
assign x_3954 = ~v_3359 | ~v_3953;
assign x_3955 = ~v_3360 | v_3952;
assign x_3956 = ~v_3360 | v_206;
assign x_3957 = ~v_3361 | v_3951;
assign x_3958 = ~v_3361 | ~v_3952;
assign x_3959 = ~v_3362 | v_213;
assign x_3960 = ~v_3362 | ~v_3952;
assign x_3961 = ~v_3363 | v_3951;
assign x_3962 = ~v_3363 | v_213;
assign x_3963 = ~v_3364 | v_3950;
assign x_3964 = ~v_3364 | ~v_3951;
assign x_3965 = ~v_3365 | v_219;
assign x_3966 = ~v_3365 | ~v_3951;
assign x_3967 = ~v_3366 | v_3950;
assign x_3968 = ~v_3366 | v_219;
assign x_3969 = ~v_3367 | v_3949;
assign x_3970 = ~v_3367 | ~v_3950;
assign x_3971 = ~v_3368 | v_224;
assign x_3972 = ~v_3368 | ~v_3950;
assign x_3973 = ~v_3369 | v_3949;
assign x_3974 = ~v_3369 | v_224;
assign x_3975 = ~v_3370 | v_3948;
assign x_3976 = ~v_3370 | ~v_3949;
assign x_3977 = ~v_3371 | v_228;
assign x_3978 = ~v_3371 | ~v_3949;
assign x_3979 = ~v_3372 | v_3948;
assign x_3980 = ~v_3372 | v_228;
assign x_3981 = ~v_3373 | v_233;
assign x_3982 = ~v_3373 | ~v_3948;
assign x_3983 = ~v_3374 | v_231;
assign x_3984 = ~v_3374 | ~v_3948;
assign x_3985 = ~v_3375 | v_233;
assign x_3986 = ~v_3375 | v_231;
assign x_3987 = ~v_3376 | v_3946;
assign x_3988 = ~v_3376 | ~v_3947;
assign x_3989 = ~v_3377 | v_199;
assign x_3990 = ~v_3377 | ~v_3947;
assign x_3991 = ~v_3378 | v_3946;
assign x_3992 = ~v_3378 | v_199;
assign x_3993 = ~v_3379 | v_3945;
assign x_3994 = ~v_3379 | ~v_3946;
assign x_3995 = ~v_3380 | v_207;
assign x_3996 = ~v_3380 | ~v_3946;
assign x_3997 = ~v_3381 | v_3945;
assign x_3998 = ~v_3381 | v_207;
assign x_3999 = ~v_3382 | v_3944;
assign x_4000 = ~v_3382 | ~v_3945;
assign x_4001 = ~v_3383 | v_214;
assign x_4002 = ~v_3383 | ~v_3945;
assign x_4003 = ~v_3384 | v_3944;
assign x_4004 = ~v_3384 | v_214;
assign x_4005 = ~v_3385 | v_3943;
assign x_4006 = ~v_3385 | ~v_3944;
assign x_4007 = ~v_3386 | v_220;
assign x_4008 = ~v_3386 | ~v_3944;
assign x_4009 = ~v_3387 | v_3943;
assign x_4010 = ~v_3387 | v_220;
assign x_4011 = ~v_3388 | v_3942;
assign x_4012 = ~v_3388 | ~v_3943;
assign x_4013 = ~v_3389 | v_225;
assign x_4014 = ~v_3389 | ~v_3943;
assign x_4015 = ~v_3390 | v_3942;
assign x_4016 = ~v_3390 | v_225;
assign x_4017 = ~v_3391 | v_3941;
assign x_4018 = ~v_3391 | ~v_3942;
assign x_4019 = ~v_3392 | v_229;
assign x_4020 = ~v_3392 | ~v_3942;
assign x_4021 = ~v_3393 | v_3941;
assign x_4022 = ~v_3393 | v_229;
assign x_4023 = ~v_3394 | v_3940;
assign x_4024 = ~v_3394 | ~v_3941;
assign x_4025 = ~v_3395 | v_232;
assign x_4026 = ~v_3395 | ~v_3941;
assign x_4027 = ~v_3396 | v_3940;
assign x_4028 = ~v_3396 | v_232;
assign x_4029 = ~v_3397 | v_235;
assign x_4030 = ~v_3397 | ~v_3940;
assign x_4031 = ~v_3398 | v_234;
assign x_4032 = ~v_3398 | ~v_3940;
assign x_4033 = ~v_3399 | v_235;
assign x_4034 = ~v_3399 | v_234;
assign x_4035 = ~v_1337 | v_1 | ~v_12;
assign x_4036 = ~v_1337 | ~v_1 | v_12 | v_388 | v_387 | v_386 | v_385 | v_384 | v_383 | v_382 | v_381 | v_380;
assign x_4037 = ~v_1337 | ~v_388 | v_1336;
assign x_4038 = ~v_1337 | ~v_56 | ~v_1 | v_2 | v_388;
assign x_4039 = ~v_1337 | ~v_387 | v_1335;
assign x_4040 = ~v_1337 | ~v_57 | ~v_1 | v_3 | v_387;
assign x_4041 = ~v_1337 | ~v_386 | v_1334;
assign x_4042 = ~v_1337 | ~v_58 | ~v_1 | v_4 | v_386;
assign x_4043 = ~v_1337 | ~v_385 | v_1333;
assign x_4044 = ~v_1337 | ~v_59 | ~v_1 | v_5 | v_385;
assign x_4045 = ~v_1337 | ~v_384 | v_1332;
assign x_4046 = ~v_1337 | ~v_60 | ~v_1 | v_6 | v_384;
assign x_4047 = ~v_1337 | ~v_383 | v_1331;
assign x_4048 = ~v_1337 | ~v_61 | ~v_1 | v_7 | v_383;
assign x_4049 = ~v_1337 | ~v_382 | v_1330;
assign x_4050 = ~v_1337 | ~v_62 | ~v_1 | v_8 | v_382;
assign x_4051 = ~v_1337 | ~v_381 | v_1329;
assign x_4052 = ~v_1337 | ~v_63 | ~v_1 | v_9 | v_381;
assign x_4053 = ~v_1337 | ~v_380 | v_1328;
assign x_4054 = ~v_1337 | ~v_64 | ~v_1 | v_10 | v_380;
assign x_4055 = ~v_1337 | v_2 | ~v_13 | v_389;
assign x_4056 = ~v_1337 | ~v_2 | v_13 | v_397 | v_396 | v_395 | v_394 | v_393 | v_392 | v_391 | v_390;
assign x_4057 = ~v_1337 | ~v_389 | v_1327;
assign x_4058 = ~v_1337 | ~v_56 | ~v_1 | v_2 | v_389;
assign x_4059 = ~v_1337 | ~v_397 | v_1326;
assign x_4060 = ~v_1337 | ~v_65 | ~v_2 | v_3 | v_397;
assign x_4061 = ~v_1337 | ~v_396 | v_1325;
assign x_4062 = ~v_1337 | ~v_66 | ~v_2 | v_4 | v_396;
assign x_4063 = ~v_1337 | ~v_395 | v_1324;
assign x_4064 = ~v_1337 | ~v_67 | ~v_2 | v_5 | v_395;
assign x_4065 = ~v_1337 | ~v_394 | v_1323;
assign x_4066 = ~v_1337 | ~v_68 | ~v_2 | v_6 | v_394;
assign x_4067 = ~v_1337 | ~v_393 | v_1322;
assign x_4068 = ~v_1337 | ~v_69 | ~v_2 | v_7 | v_393;
assign x_4069 = ~v_1337 | ~v_392 | v_1321;
assign x_4070 = ~v_1337 | ~v_70 | ~v_2 | v_8 | v_392;
assign x_4071 = ~v_1337 | ~v_391 | v_1320;
assign x_4072 = ~v_1337 | ~v_71 | ~v_2 | v_9 | v_391;
assign x_4073 = ~v_1337 | ~v_390 | v_1319;
assign x_4074 = ~v_1337 | ~v_72 | ~v_2 | v_10 | v_390;
assign x_4075 = ~v_1337 | v_3 | ~v_14 | v_399 | v_398;
assign x_4076 = ~v_1337 | ~v_3 | v_14 | v_406 | v_405 | v_404 | v_403 | v_402 | v_401 | v_400;
assign x_4077 = ~v_1337 | ~v_399 | v_1318;
assign x_4078 = ~v_1337 | ~v_57 | ~v_1 | v_3 | v_399;
assign x_4079 = ~v_1337 | ~v_398 | v_1317;
assign x_4080 = ~v_1337 | ~v_65 | ~v_2 | v_3 | v_398;
assign x_4081 = ~v_1337 | ~v_406 | v_1316;
assign x_4082 = ~v_1337 | ~v_73 | ~v_3 | v_4 | v_406;
assign x_4083 = ~v_1337 | ~v_405 | v_1315;
assign x_4084 = ~v_1337 | ~v_74 | ~v_3 | v_5 | v_405;
assign x_4085 = ~v_1337 | ~v_404 | v_1314;
assign x_4086 = ~v_1337 | ~v_75 | ~v_3 | v_6 | v_404;
assign x_4087 = ~v_1337 | ~v_403 | v_1313;
assign x_4088 = ~v_1337 | ~v_76 | ~v_3 | v_7 | v_403;
assign x_4089 = ~v_1337 | ~v_402 | v_1312;
assign x_4090 = ~v_1337 | ~v_77 | ~v_3 | v_8 | v_402;
assign x_4091 = ~v_1337 | ~v_401 | v_1311;
assign x_4092 = ~v_1337 | ~v_78 | ~v_3 | v_9 | v_401;
assign x_4093 = ~v_1337 | ~v_400 | v_1310;
assign x_4094 = ~v_1337 | ~v_79 | ~v_3 | v_10 | v_400;
assign x_4095 = ~v_1337 | v_4 | ~v_15 | v_409 | v_408 | v_407;
assign x_4096 = ~v_1337 | ~v_4 | v_15 | v_415 | v_414 | v_413 | v_412 | v_411 | v_410;
assign x_4097 = ~v_1337 | ~v_409 | v_1309;
assign x_4098 = ~v_1337 | ~v_58 | ~v_1 | v_4 | v_409;
assign x_4099 = ~v_1337 | ~v_408 | v_1308;
assign x_4100 = ~v_1337 | ~v_66 | ~v_2 | v_4 | v_408;
assign x_4101 = ~v_1337 | ~v_407 | v_1307;
assign x_4102 = ~v_1337 | ~v_73 | ~v_3 | v_4 | v_407;
assign x_4103 = ~v_1337 | ~v_415 | v_1306;
assign x_4104 = ~v_1337 | ~v_80 | ~v_4 | v_5 | v_415;
assign x_4105 = ~v_1337 | ~v_414 | v_1305;
assign x_4106 = ~v_1337 | ~v_81 | ~v_4 | v_6 | v_414;
assign x_4107 = ~v_1337 | ~v_413 | v_1304;
assign x_4108 = ~v_1337 | ~v_82 | ~v_4 | v_7 | v_413;
assign x_4109 = ~v_1337 | ~v_412 | v_1303;
assign x_4110 = ~v_1337 | ~v_83 | ~v_4 | v_8 | v_412;
assign x_4111 = ~v_1337 | ~v_411 | v_1302;
assign x_4112 = ~v_1337 | ~v_84 | ~v_4 | v_9 | v_411;
assign x_4113 = ~v_1337 | ~v_410 | v_1301;
assign x_4114 = ~v_1337 | ~v_85 | ~v_4 | v_10 | v_410;
assign x_4115 = ~v_1337 | v_5 | ~v_16 | v_419 | v_418 | v_417 | v_416;
assign x_4116 = ~v_1337 | ~v_5 | v_16 | v_424 | v_423 | v_422 | v_421 | v_420;
assign x_4117 = ~v_1337 | ~v_419 | v_1300;
assign x_4118 = ~v_1337 | ~v_59 | ~v_1 | v_5 | v_419;
assign x_4119 = ~v_1337 | ~v_418 | v_1299;
assign x_4120 = ~v_1337 | ~v_67 | ~v_2 | v_5 | v_418;
assign x_4121 = ~v_1337 | ~v_417 | v_1298;
assign x_4122 = ~v_1337 | ~v_74 | ~v_3 | v_5 | v_417;
assign x_4123 = ~v_1337 | ~v_416 | v_1297;
assign x_4124 = ~v_1337 | ~v_80 | ~v_4 | v_5 | v_416;
assign x_4125 = ~v_1337 | ~v_424 | v_1296;
assign x_4126 = ~v_1337 | ~v_86 | ~v_5 | v_6 | v_424;
assign x_4127 = ~v_1337 | ~v_423 | v_1295;
assign x_4128 = ~v_1337 | ~v_87 | ~v_5 | v_7 | v_423;
assign x_4129 = ~v_1337 | ~v_422 | v_1294;
assign x_4130 = ~v_1337 | ~v_88 | ~v_5 | v_8 | v_422;
assign x_4131 = ~v_1337 | ~v_421 | v_1293;
assign x_4132 = ~v_1337 | ~v_89 | ~v_5 | v_9 | v_421;
assign x_4133 = ~v_1337 | ~v_420 | v_1292;
assign x_4134 = ~v_1337 | ~v_90 | ~v_5 | v_10 | v_420;
assign x_4135 = ~v_1337 | v_6 | ~v_17 | v_429 | v_428 | v_427 | v_426 | v_425;
assign x_4136 = ~v_1337 | ~v_6 | v_17 | v_433 | v_432 | v_431 | v_430;
assign x_4137 = ~v_1337 | ~v_429 | v_1291;
assign x_4138 = ~v_1337 | ~v_60 | ~v_1 | v_6 | v_429;
assign x_4139 = ~v_1337 | ~v_428 | v_1290;
assign x_4140 = ~v_1337 | ~v_68 | ~v_2 | v_6 | v_428;
assign x_4141 = ~v_1337 | ~v_427 | v_1289;
assign x_4142 = ~v_1337 | ~v_75 | ~v_3 | v_6 | v_427;
assign x_4143 = ~v_1337 | ~v_426 | v_1288;
assign x_4144 = ~v_1337 | ~v_81 | ~v_4 | v_6 | v_426;
assign x_4145 = ~v_1337 | ~v_425 | v_1287;
assign x_4146 = ~v_1337 | ~v_86 | ~v_5 | v_6 | v_425;
assign x_4147 = ~v_1337 | ~v_433 | v_1286;
assign x_4148 = ~v_1337 | ~v_91 | ~v_6 | v_7 | v_433;
assign x_4149 = ~v_1337 | ~v_432 | v_1285;
assign x_4150 = ~v_1337 | ~v_92 | ~v_6 | v_8 | v_432;
assign x_4151 = ~v_1337 | ~v_431 | v_1284;
assign x_4152 = ~v_1337 | ~v_93 | ~v_6 | v_9 | v_431;
assign x_4153 = ~v_1337 | ~v_430 | v_1283;
assign x_4154 = ~v_1337 | ~v_94 | ~v_6 | v_10 | v_430;
assign x_4155 = ~v_1337 | v_7 | ~v_18 | v_439 | v_438 | v_437 | v_436 | v_435 | v_434;
assign x_4156 = ~v_1337 | ~v_7 | v_18 | v_442 | v_441 | v_440;
assign x_4157 = ~v_1337 | ~v_439 | v_1282;
assign x_4158 = ~v_1337 | ~v_61 | ~v_1 | v_7 | v_439;
assign x_4159 = ~v_1337 | ~v_438 | v_1281;
assign x_4160 = ~v_1337 | ~v_69 | ~v_2 | v_7 | v_438;
assign x_4161 = ~v_1337 | ~v_437 | v_1280;
assign x_4162 = ~v_1337 | ~v_76 | ~v_3 | v_7 | v_437;
assign x_4163 = ~v_1337 | ~v_436 | v_1279;
assign x_4164 = ~v_1337 | ~v_82 | ~v_4 | v_7 | v_436;
assign x_4165 = ~v_1337 | ~v_435 | v_1278;
assign x_4166 = ~v_1337 | ~v_87 | ~v_5 | v_7 | v_435;
assign x_4167 = ~v_1337 | ~v_434 | v_1277;
assign x_4168 = ~v_1337 | ~v_91 | ~v_6 | v_7 | v_434;
assign x_4169 = ~v_1337 | ~v_442 | v_1276;
assign x_4170 = ~v_1337 | ~v_95 | ~v_7 | v_8 | v_442;
assign x_4171 = ~v_1337 | ~v_441 | v_1275;
assign x_4172 = ~v_1337 | ~v_96 | ~v_7 | v_9 | v_441;
assign x_4173 = ~v_1337 | ~v_440 | v_1274;
assign x_4174 = ~v_1337 | ~v_97 | ~v_7 | v_10 | v_440;
assign x_4175 = ~v_1337 | v_8 | ~v_19 | v_449 | v_448 | v_447 | v_446 | v_445 | v_444 | v_443;
assign x_4176 = ~v_1337 | ~v_8 | v_19 | v_451 | v_450;
assign x_4177 = ~v_1337 | ~v_449 | v_1273;
assign x_4178 = ~v_1337 | ~v_62 | ~v_1 | v_8 | v_449;
assign x_4179 = ~v_1337 | ~v_448 | v_1272;
assign x_4180 = ~v_1337 | ~v_70 | ~v_2 | v_8 | v_448;
assign x_4181 = ~v_1337 | ~v_447 | v_1271;
assign x_4182 = ~v_1337 | ~v_77 | ~v_3 | v_8 | v_447;
assign x_4183 = ~v_1337 | ~v_446 | v_1270;
assign x_4184 = ~v_1337 | ~v_83 | ~v_4 | v_8 | v_446;
assign x_4185 = ~v_1337 | ~v_445 | v_1269;
assign x_4186 = ~v_1337 | ~v_88 | ~v_5 | v_8 | v_445;
assign x_4187 = ~v_1337 | ~v_444 | v_1268;
assign x_4188 = ~v_1337 | ~v_92 | ~v_6 | v_8 | v_444;
assign x_4189 = ~v_1337 | ~v_443 | v_1267;
assign x_4190 = ~v_1337 | ~v_95 | ~v_7 | v_8 | v_443;
assign x_4191 = ~v_1337 | ~v_451 | v_1266;
assign x_4192 = ~v_1337 | ~v_98 | ~v_8 | v_9 | v_451;
assign x_4193 = ~v_1337 | ~v_450 | v_1265;
assign x_4194 = ~v_1337 | ~v_99 | ~v_8 | v_10 | v_450;
assign x_4195 = ~v_1337 | v_9 | ~v_20 | v_459 | v_458 | v_457 | v_456 | v_455 | v_454 | v_453 | v_452;
assign x_4196 = ~v_1337 | ~v_9 | v_20 | v_460;
assign x_4197 = ~v_1337 | ~v_459 | v_1264;
assign x_4198 = ~v_1337 | ~v_63 | ~v_1 | v_9 | v_459;
assign x_4199 = ~v_1337 | ~v_458 | v_1263;
assign x_4200 = ~v_1337 | ~v_71 | ~v_2 | v_9 | v_458;
assign x_4201 = ~v_1337 | ~v_457 | v_1262;
assign x_4202 = ~v_1337 | ~v_78 | ~v_3 | v_9 | v_457;
assign x_4203 = ~v_1337 | ~v_456 | v_1261;
assign x_4204 = ~v_1337 | ~v_84 | ~v_4 | v_9 | v_456;
assign x_4205 = ~v_1337 | ~v_455 | v_1260;
assign x_4206 = ~v_1337 | ~v_89 | ~v_5 | v_9 | v_455;
assign x_4207 = ~v_1337 | ~v_454 | v_1259;
assign x_4208 = ~v_1337 | ~v_93 | ~v_6 | v_9 | v_454;
assign x_4209 = ~v_1337 | ~v_453 | v_1258;
assign x_4210 = ~v_1337 | ~v_96 | ~v_7 | v_9 | v_453;
assign x_4211 = ~v_1337 | ~v_452 | v_1257;
assign x_4212 = ~v_1337 | ~v_98 | ~v_8 | v_9 | v_452;
assign x_4213 = ~v_1337 | ~v_460 | v_1256;
assign x_4214 = ~v_1337 | ~v_100 | ~v_9 | v_10 | v_460;
assign x_4215 = ~v_1337 | v_10 | ~v_21 | v_469 | v_468 | v_467 | v_466 | v_465 | v_464 | v_463 | v_462 | v_461;
assign x_4216 = ~v_1337 | ~v_10 | v_21;
assign x_4217 = ~v_1337 | ~v_469 | v_1255;
assign x_4218 = ~v_1337 | ~v_64 | ~v_1 | v_10 | v_469;
assign x_4219 = ~v_1337 | ~v_468 | v_1254;
assign x_4220 = ~v_1337 | ~v_72 | ~v_2 | v_10 | v_468;
assign x_4221 = ~v_1337 | ~v_467 | v_1253;
assign x_4222 = ~v_1337 | ~v_79 | ~v_3 | v_10 | v_467;
assign x_4223 = ~v_1337 | ~v_466 | v_1252;
assign x_4224 = ~v_1337 | ~v_85 | ~v_4 | v_10 | v_466;
assign x_4225 = ~v_1337 | ~v_465 | v_1251;
assign x_4226 = ~v_1337 | ~v_90 | ~v_5 | v_10 | v_465;
assign x_4227 = ~v_1337 | ~v_464 | v_1250;
assign x_4228 = ~v_1337 | ~v_94 | ~v_6 | v_10 | v_464;
assign x_4229 = ~v_1337 | ~v_463 | v_1249;
assign x_4230 = ~v_1337 | ~v_97 | ~v_7 | v_10 | v_463;
assign x_4231 = ~v_1337 | ~v_462 | v_1248;
assign x_4232 = ~v_1337 | ~v_99 | ~v_8 | v_10 | v_462;
assign x_4233 = ~v_1337 | ~v_461 | v_1247;
assign x_4234 = ~v_1337 | ~v_100 | ~v_9 | v_10 | v_461;
assign x_4235 = ~v_1337 | v_11 | ~v_22;
assign x_4236 = ~v_1337 | ~v_11 | v_22;
assign x_4237 = ~v_1337 | v_1245 | v_1246;
assign x_4238 = ~v_1337 | v_1243 | v_1244;
assign x_4239 = ~v_1337 | v_1241 | v_1242;
assign x_4240 = ~v_1337 | v_1239 | v_1240;
assign x_4241 = ~v_1337 | v_1237 | v_1238;
assign x_4242 = ~v_1337 | v_1235 | v_1236;
assign x_4243 = ~v_1337 | v_1233 | v_1234;
assign x_4244 = ~v_1337 | v_1231 | v_1232;
assign x_4245 = ~v_1337 | v_1229 | v_1230;
assign x_4246 = ~v_1337 | v_1227 | v_1228;
assign x_4247 = ~v_1337 | v_1225 | v_1226;
assign x_4248 = ~v_1337 | v_1223 | v_1224;
assign x_4249 = ~v_1337 | v_1221 | v_1222;
assign x_4250 = ~v_1337 | v_1219 | v_1220;
assign x_4251 = ~v_1337 | v_1217 | v_1218;
assign x_4252 = ~v_1337 | v_1215 | v_1216;
assign x_4253 = ~v_1337 | v_1213 | v_1214;
assign x_4254 = ~v_1337 | v_1211 | v_1212;
assign x_4255 = ~v_1337 | v_1209 | v_1210;
assign x_4256 = ~v_1337 | v_1207 | v_1208;
assign x_4257 = ~v_1337 | v_1205 | v_1206;
assign x_4258 = ~v_1337 | v_1203 | v_1204;
assign x_4259 = ~v_1337 | v_1201 | v_1202;
assign x_4260 = ~v_1337 | v_1199 | v_1200;
assign x_4261 = ~v_1337 | v_1197 | v_1198;
assign x_4262 = ~v_1337 | v_1195 | v_1196;
assign x_4263 = ~v_1337 | v_1193 | v_1194;
assign x_4264 = ~v_1337 | v_1191 | v_1192;
assign x_4265 = ~v_1337 | v_1189 | v_1190;
assign x_4266 = ~v_1337 | v_1187 | v_1188;
assign x_4267 = ~v_1337 | v_1185 | v_1186;
assign x_4268 = ~v_1337 | v_1183 | v_1184;
assign x_4269 = ~v_1337 | v_1181 | v_1182;
assign x_4270 = ~v_1337 | v_1179 | v_1180;
assign x_4271 = ~v_1337 | v_1177 | v_1178;
assign x_4272 = ~v_1337 | v_1175 | v_1176;
assign x_4273 = ~v_1337 | v_1173 | v_1174;
assign x_4274 = ~v_1337 | v_1171 | v_1172;
assign x_4275 = ~v_1337 | v_1169 | v_1170;
assign x_4276 = ~v_1337 | v_1167 | v_1168;
assign x_4277 = ~v_1337 | v_1165 | v_1166;
assign x_4278 = ~v_1337 | v_1163 | v_1164;
assign x_4279 = ~v_1337 | v_1161 | v_1162;
assign x_4280 = ~v_1337 | v_1159 | v_1160;
assign x_4281 = ~v_1337 | v_1157 | v_1158;
assign x_4282 = ~v_1337 | v_1111;
assign x_4283 = ~v_1336 | v_56;
assign x_4284 = ~v_1336 | v_1;
assign x_4285 = ~v_1336 | ~v_2;
assign x_4286 = ~v_1335 | v_57;
assign x_4287 = ~v_1335 | v_1;
assign x_4288 = ~v_1335 | ~v_3;
assign x_4289 = ~v_1334 | v_58;
assign x_4290 = ~v_1334 | v_1;
assign x_4291 = ~v_1334 | ~v_4;
assign x_4292 = ~v_1333 | v_59;
assign x_4293 = ~v_1333 | v_1;
assign x_4294 = ~v_1333 | ~v_5;
assign x_4295 = ~v_1332 | v_60;
assign x_4296 = ~v_1332 | v_1;
assign x_4297 = ~v_1332 | ~v_6;
assign x_4298 = ~v_1331 | v_61;
assign x_4299 = ~v_1331 | v_1;
assign x_4300 = ~v_1331 | ~v_7;
assign x_4301 = ~v_1330 | v_62;
assign x_4302 = ~v_1330 | v_1;
assign x_4303 = ~v_1330 | ~v_8;
assign x_4304 = ~v_1329 | v_63;
assign x_4305 = ~v_1329 | v_1;
assign x_4306 = ~v_1329 | ~v_9;
assign x_4307 = ~v_1328 | v_64;
assign x_4308 = ~v_1328 | v_1;
assign x_4309 = ~v_1328 | ~v_10;
assign x_4310 = ~v_1327 | v_56;
assign x_4311 = ~v_1327 | v_1;
assign x_4312 = ~v_1327 | ~v_2;
assign x_4313 = ~v_1326 | v_65;
assign x_4314 = ~v_1326 | v_2;
assign x_4315 = ~v_1326 | ~v_3;
assign x_4316 = ~v_1325 | v_66;
assign x_4317 = ~v_1325 | v_2;
assign x_4318 = ~v_1325 | ~v_4;
assign x_4319 = ~v_1324 | v_67;
assign x_4320 = ~v_1324 | v_2;
assign x_4321 = ~v_1324 | ~v_5;
assign x_4322 = ~v_1323 | v_68;
assign x_4323 = ~v_1323 | v_2;
assign x_4324 = ~v_1323 | ~v_6;
assign x_4325 = ~v_1322 | v_69;
assign x_4326 = ~v_1322 | v_2;
assign x_4327 = ~v_1322 | ~v_7;
assign x_4328 = ~v_1321 | v_70;
assign x_4329 = ~v_1321 | v_2;
assign x_4330 = ~v_1321 | ~v_8;
assign x_4331 = ~v_1320 | v_71;
assign x_4332 = ~v_1320 | v_2;
assign x_4333 = ~v_1320 | ~v_9;
assign x_4334 = ~v_1319 | v_72;
assign x_4335 = ~v_1319 | v_2;
assign x_4336 = ~v_1319 | ~v_10;
assign x_4337 = ~v_1318 | v_57;
assign x_4338 = ~v_1318 | v_1;
assign x_4339 = ~v_1318 | ~v_3;
assign x_4340 = ~v_1317 | v_65;
assign x_4341 = ~v_1317 | v_2;
assign x_4342 = ~v_1317 | ~v_3;
assign x_4343 = ~v_1316 | v_73;
assign x_4344 = ~v_1316 | v_3;
assign x_4345 = ~v_1316 | ~v_4;
assign x_4346 = ~v_1315 | v_74;
assign x_4347 = ~v_1315 | v_3;
assign x_4348 = ~v_1315 | ~v_5;
assign x_4349 = ~v_1314 | v_75;
assign x_4350 = ~v_1314 | v_3;
assign x_4351 = ~v_1314 | ~v_6;
assign x_4352 = ~v_1313 | v_76;
assign x_4353 = ~v_1313 | v_3;
assign x_4354 = ~v_1313 | ~v_7;
assign x_4355 = ~v_1312 | v_77;
assign x_4356 = ~v_1312 | v_3;
assign x_4357 = ~v_1312 | ~v_8;
assign x_4358 = ~v_1311 | v_78;
assign x_4359 = ~v_1311 | v_3;
assign x_4360 = ~v_1311 | ~v_9;
assign x_4361 = ~v_1310 | v_79;
assign x_4362 = ~v_1310 | v_3;
assign x_4363 = ~v_1310 | ~v_10;
assign x_4364 = ~v_1309 | v_58;
assign x_4365 = ~v_1309 | v_1;
assign x_4366 = ~v_1309 | ~v_4;
assign x_4367 = ~v_1308 | v_66;
assign x_4368 = ~v_1308 | v_2;
assign x_4369 = ~v_1308 | ~v_4;
assign x_4370 = ~v_1307 | v_73;
assign x_4371 = ~v_1307 | v_3;
assign x_4372 = ~v_1307 | ~v_4;
assign x_4373 = ~v_1306 | v_80;
assign x_4374 = ~v_1306 | v_4;
assign x_4375 = ~v_1306 | ~v_5;
assign x_4376 = ~v_1305 | v_81;
assign x_4377 = ~v_1305 | v_4;
assign x_4378 = ~v_1305 | ~v_6;
assign x_4379 = ~v_1304 | v_82;
assign x_4380 = ~v_1304 | v_4;
assign x_4381 = ~v_1304 | ~v_7;
assign x_4382 = ~v_1303 | v_83;
assign x_4383 = ~v_1303 | v_4;
assign x_4384 = ~v_1303 | ~v_8;
assign x_4385 = ~v_1302 | v_84;
assign x_4386 = ~v_1302 | v_4;
assign x_4387 = ~v_1302 | ~v_9;
assign x_4388 = ~v_1301 | v_85;
assign x_4389 = ~v_1301 | v_4;
assign x_4390 = ~v_1301 | ~v_10;
assign x_4391 = ~v_1300 | v_59;
assign x_4392 = ~v_1300 | v_1;
assign x_4393 = ~v_1300 | ~v_5;
assign x_4394 = ~v_1299 | v_67;
assign x_4395 = ~v_1299 | v_2;
assign x_4396 = ~v_1299 | ~v_5;
assign x_4397 = ~v_1298 | v_74;
assign x_4398 = ~v_1298 | v_3;
assign x_4399 = ~v_1298 | ~v_5;
assign x_4400 = ~v_1297 | v_80;
assign x_4401 = ~v_1297 | v_4;
assign x_4402 = ~v_1297 | ~v_5;
assign x_4403 = ~v_1296 | v_86;
assign x_4404 = ~v_1296 | v_5;
assign x_4405 = ~v_1296 | ~v_6;
assign x_4406 = ~v_1295 | v_87;
assign x_4407 = ~v_1295 | v_5;
assign x_4408 = ~v_1295 | ~v_7;
assign x_4409 = ~v_1294 | v_88;
assign x_4410 = ~v_1294 | v_5;
assign x_4411 = ~v_1294 | ~v_8;
assign x_4412 = ~v_1293 | v_89;
assign x_4413 = ~v_1293 | v_5;
assign x_4414 = ~v_1293 | ~v_9;
assign x_4415 = ~v_1292 | v_90;
assign x_4416 = ~v_1292 | v_5;
assign x_4417 = ~v_1292 | ~v_10;
assign x_4418 = ~v_1291 | v_60;
assign x_4419 = ~v_1291 | v_1;
assign x_4420 = ~v_1291 | ~v_6;
assign x_4421 = ~v_1290 | v_68;
assign x_4422 = ~v_1290 | v_2;
assign x_4423 = ~v_1290 | ~v_6;
assign x_4424 = ~v_1289 | v_75;
assign x_4425 = ~v_1289 | v_3;
assign x_4426 = ~v_1289 | ~v_6;
assign x_4427 = ~v_1288 | v_81;
assign x_4428 = ~v_1288 | v_4;
assign x_4429 = ~v_1288 | ~v_6;
assign x_4430 = ~v_1287 | v_86;
assign x_4431 = ~v_1287 | v_5;
assign x_4432 = ~v_1287 | ~v_6;
assign x_4433 = ~v_1286 | v_91;
assign x_4434 = ~v_1286 | v_6;
assign x_4435 = ~v_1286 | ~v_7;
assign x_4436 = ~v_1285 | v_92;
assign x_4437 = ~v_1285 | v_6;
assign x_4438 = ~v_1285 | ~v_8;
assign x_4439 = ~v_1284 | v_93;
assign x_4440 = ~v_1284 | v_6;
assign x_4441 = ~v_1284 | ~v_9;
assign x_4442 = ~v_1283 | v_94;
assign x_4443 = ~v_1283 | v_6;
assign x_4444 = ~v_1283 | ~v_10;
assign x_4445 = ~v_1282 | v_61;
assign x_4446 = ~v_1282 | v_1;
assign x_4447 = ~v_1282 | ~v_7;
assign x_4448 = ~v_1281 | v_69;
assign x_4449 = ~v_1281 | v_2;
assign x_4450 = ~v_1281 | ~v_7;
assign x_4451 = ~v_1280 | v_76;
assign x_4452 = ~v_1280 | v_3;
assign x_4453 = ~v_1280 | ~v_7;
assign x_4454 = ~v_1279 | v_82;
assign x_4455 = ~v_1279 | v_4;
assign x_4456 = ~v_1279 | ~v_7;
assign x_4457 = ~v_1278 | v_87;
assign x_4458 = ~v_1278 | v_5;
assign x_4459 = ~v_1278 | ~v_7;
assign x_4460 = ~v_1277 | v_91;
assign x_4461 = ~v_1277 | v_6;
assign x_4462 = ~v_1277 | ~v_7;
assign x_4463 = ~v_1276 | v_95;
assign x_4464 = ~v_1276 | v_7;
assign x_4465 = ~v_1276 | ~v_8;
assign x_4466 = ~v_1275 | v_96;
assign x_4467 = ~v_1275 | v_7;
assign x_4468 = ~v_1275 | ~v_9;
assign x_4469 = ~v_1274 | v_97;
assign x_4470 = ~v_1274 | v_7;
assign x_4471 = ~v_1274 | ~v_10;
assign x_4472 = ~v_1273 | v_62;
assign x_4473 = ~v_1273 | v_1;
assign x_4474 = ~v_1273 | ~v_8;
assign x_4475 = ~v_1272 | v_70;
assign x_4476 = ~v_1272 | v_2;
assign x_4477 = ~v_1272 | ~v_8;
assign x_4478 = ~v_1271 | v_77;
assign x_4479 = ~v_1271 | v_3;
assign x_4480 = ~v_1271 | ~v_8;
assign x_4481 = ~v_1270 | v_83;
assign x_4482 = ~v_1270 | v_4;
assign x_4483 = ~v_1270 | ~v_8;
assign x_4484 = ~v_1269 | v_88;
assign x_4485 = ~v_1269 | v_5;
assign x_4486 = ~v_1269 | ~v_8;
assign x_4487 = ~v_1268 | v_92;
assign x_4488 = ~v_1268 | v_6;
assign x_4489 = ~v_1268 | ~v_8;
assign x_4490 = ~v_1267 | v_95;
assign x_4491 = ~v_1267 | v_7;
assign x_4492 = ~v_1267 | ~v_8;
assign x_4493 = ~v_1266 | v_98;
assign x_4494 = ~v_1266 | v_8;
assign x_4495 = ~v_1266 | ~v_9;
assign x_4496 = ~v_1265 | v_99;
assign x_4497 = ~v_1265 | v_8;
assign x_4498 = ~v_1265 | ~v_10;
assign x_4499 = ~v_1264 | v_63;
assign x_4500 = ~v_1264 | v_1;
assign x_4501 = ~v_1264 | ~v_9;
assign x_4502 = ~v_1263 | v_71;
assign x_4503 = ~v_1263 | v_2;
assign x_4504 = ~v_1263 | ~v_9;
assign x_4505 = ~v_1262 | v_78;
assign x_4506 = ~v_1262 | v_3;
assign x_4507 = ~v_1262 | ~v_9;
assign x_4508 = ~v_1261 | v_84;
assign x_4509 = ~v_1261 | v_4;
assign x_4510 = ~v_1261 | ~v_9;
assign x_4511 = ~v_1260 | v_89;
assign x_4512 = ~v_1260 | v_5;
assign x_4513 = ~v_1260 | ~v_9;
assign x_4514 = ~v_1259 | v_93;
assign x_4515 = ~v_1259 | v_6;
assign x_4516 = ~v_1259 | ~v_9;
assign x_4517 = ~v_1258 | v_96;
assign x_4518 = ~v_1258 | v_7;
assign x_4519 = ~v_1258 | ~v_9;
assign x_4520 = ~v_1257 | v_98;
assign x_4521 = ~v_1257 | v_8;
assign x_4522 = ~v_1257 | ~v_9;
assign x_4523 = ~v_1256 | v_100;
assign x_4524 = ~v_1256 | v_9;
assign x_4525 = ~v_1256 | ~v_10;
assign x_4526 = ~v_1255 | v_64;
assign x_4527 = ~v_1255 | v_1;
assign x_4528 = ~v_1255 | ~v_10;
assign x_4529 = ~v_1254 | v_72;
assign x_4530 = ~v_1254 | v_2;
assign x_4531 = ~v_1254 | ~v_10;
assign x_4532 = ~v_1253 | v_79;
assign x_4533 = ~v_1253 | v_3;
assign x_4534 = ~v_1253 | ~v_10;
assign x_4535 = ~v_1252 | v_85;
assign x_4536 = ~v_1252 | v_4;
assign x_4537 = ~v_1252 | ~v_10;
assign x_4538 = ~v_1251 | v_90;
assign x_4539 = ~v_1251 | v_5;
assign x_4540 = ~v_1251 | ~v_10;
assign x_4541 = ~v_1250 | v_94;
assign x_4542 = ~v_1250 | v_6;
assign x_4543 = ~v_1250 | ~v_10;
assign x_4544 = ~v_1249 | v_97;
assign x_4545 = ~v_1249 | v_7;
assign x_4546 = ~v_1249 | ~v_10;
assign x_4547 = ~v_1248 | v_99;
assign x_4548 = ~v_1248 | v_8;
assign x_4549 = ~v_1248 | ~v_10;
assign x_4550 = ~v_1247 | v_100;
assign x_4551 = ~v_1247 | v_9;
assign x_4552 = ~v_1247 | ~v_10;
assign x_4553 = ~v_1245 | ~v_56 | ~v_1 | v_2;
assign x_4554 = ~v_1246 | ~v_12;
assign x_4555 = ~v_1246 | v_13;
assign x_4556 = ~v_1243 | ~v_57 | ~v_1 | v_3;
assign x_4557 = ~v_1244 | ~v_12;
assign x_4558 = ~v_1244 | v_14;
assign x_4559 = ~v_1241 | ~v_58 | ~v_1 | v_4;
assign x_4560 = ~v_1242 | ~v_12;
assign x_4561 = ~v_1242 | v_15;
assign x_4562 = ~v_1239 | ~v_59 | ~v_1 | v_5;
assign x_4563 = ~v_1240 | ~v_12;
assign x_4564 = ~v_1240 | v_16;
assign x_4565 = ~v_1237 | ~v_60 | ~v_1 | v_6;
assign x_4566 = ~v_1238 | ~v_12;
assign x_4567 = ~v_1238 | v_17;
assign x_4568 = ~v_1235 | ~v_61 | ~v_1 | v_7;
assign x_4569 = ~v_1236 | ~v_12;
assign x_4570 = ~v_1236 | v_18;
assign x_4571 = ~v_1233 | ~v_62 | ~v_1 | v_8;
assign x_4572 = ~v_1234 | ~v_12;
assign x_4573 = ~v_1234 | v_19;
assign x_4574 = ~v_1231 | ~v_63 | ~v_1 | v_9;
assign x_4575 = ~v_1232 | ~v_12;
assign x_4576 = ~v_1232 | v_20;
assign x_4577 = ~v_1229 | ~v_64 | ~v_1 | v_10;
assign x_4578 = ~v_1230 | ~v_12;
assign x_4579 = ~v_1230 | v_21;
assign x_4580 = ~v_1227 | ~v_65 | ~v_2 | v_3;
assign x_4581 = ~v_1228 | ~v_13;
assign x_4582 = ~v_1228 | v_14;
assign x_4583 = ~v_1225 | ~v_66 | ~v_2 | v_4;
assign x_4584 = ~v_1226 | ~v_13;
assign x_4585 = ~v_1226 | v_15;
assign x_4586 = ~v_1223 | ~v_67 | ~v_2 | v_5;
assign x_4587 = ~v_1224 | ~v_13;
assign x_4588 = ~v_1224 | v_16;
assign x_4589 = ~v_1221 | ~v_68 | ~v_2 | v_6;
assign x_4590 = ~v_1222 | ~v_13;
assign x_4591 = ~v_1222 | v_17;
assign x_4592 = ~v_1219 | ~v_69 | ~v_2 | v_7;
assign x_4593 = ~v_1220 | ~v_13;
assign x_4594 = ~v_1220 | v_18;
assign x_4595 = ~v_1217 | ~v_70 | ~v_2 | v_8;
assign x_4596 = ~v_1218 | ~v_13;
assign x_4597 = ~v_1218 | v_19;
assign x_4598 = ~v_1215 | ~v_71 | ~v_2 | v_9;
assign x_4599 = ~v_1216 | ~v_13;
assign x_4600 = ~v_1216 | v_20;
assign x_4601 = ~v_1213 | ~v_72 | ~v_2 | v_10;
assign x_4602 = ~v_1214 | ~v_13;
assign x_4603 = ~v_1214 | v_21;
assign x_4604 = ~v_1211 | ~v_73 | ~v_3 | v_4;
assign x_4605 = ~v_1212 | ~v_14;
assign x_4606 = ~v_1212 | v_15;
assign x_4607 = ~v_1209 | ~v_74 | ~v_3 | v_5;
assign x_4608 = ~v_1210 | ~v_14;
assign x_4609 = ~v_1210 | v_16;
assign x_4610 = ~v_1207 | ~v_75 | ~v_3 | v_6;
assign x_4611 = ~v_1208 | ~v_14;
assign x_4612 = ~v_1208 | v_17;
assign x_4613 = ~v_1205 | ~v_76 | ~v_3 | v_7;
assign x_4614 = ~v_1206 | ~v_14;
assign x_4615 = ~v_1206 | v_18;
assign x_4616 = ~v_1203 | ~v_77 | ~v_3 | v_8;
assign x_4617 = ~v_1204 | ~v_14;
assign x_4618 = ~v_1204 | v_19;
assign x_4619 = ~v_1201 | ~v_78 | ~v_3 | v_9;
assign x_4620 = ~v_1202 | ~v_14;
assign x_4621 = ~v_1202 | v_20;
assign x_4622 = ~v_1199 | ~v_79 | ~v_3 | v_10;
assign x_4623 = ~v_1200 | ~v_14;
assign x_4624 = ~v_1200 | v_21;
assign x_4625 = ~v_1197 | ~v_80 | ~v_4 | v_5;
assign x_4626 = ~v_1198 | ~v_15;
assign x_4627 = ~v_1198 | v_16;
assign x_4628 = ~v_1195 | ~v_81 | ~v_4 | v_6;
assign x_4629 = ~v_1196 | ~v_15;
assign x_4630 = ~v_1196 | v_17;
assign x_4631 = ~v_1193 | ~v_82 | ~v_4 | v_7;
assign x_4632 = ~v_1194 | ~v_15;
assign x_4633 = ~v_1194 | v_18;
assign x_4634 = ~v_1191 | ~v_83 | ~v_4 | v_8;
assign x_4635 = ~v_1192 | ~v_15;
assign x_4636 = ~v_1192 | v_19;
assign x_4637 = ~v_1189 | ~v_84 | ~v_4 | v_9;
assign x_4638 = ~v_1190 | ~v_15;
assign x_4639 = ~v_1190 | v_20;
assign x_4640 = ~v_1187 | ~v_85 | ~v_4 | v_10;
assign x_4641 = ~v_1188 | ~v_15;
assign x_4642 = ~v_1188 | v_21;
assign x_4643 = ~v_1185 | ~v_86 | ~v_5 | v_6;
assign x_4644 = ~v_1186 | ~v_16;
assign x_4645 = ~v_1186 | v_17;
assign x_4646 = ~v_1183 | ~v_87 | ~v_5 | v_7;
assign x_4647 = ~v_1184 | ~v_16;
assign x_4648 = ~v_1184 | v_18;
assign x_4649 = ~v_1181 | ~v_88 | ~v_5 | v_8;
assign x_4650 = ~v_1182 | ~v_16;
assign x_4651 = ~v_1182 | v_19;
assign x_4652 = ~v_1179 | ~v_89 | ~v_5 | v_9;
assign x_4653 = ~v_1180 | ~v_16;
assign x_4654 = ~v_1180 | v_20;
assign x_4655 = ~v_1177 | ~v_90 | ~v_5 | v_10;
assign x_4656 = ~v_1178 | ~v_16;
assign x_4657 = ~v_1178 | v_21;
assign x_4658 = ~v_1175 | ~v_91 | ~v_6 | v_7;
assign x_4659 = ~v_1176 | ~v_17;
assign x_4660 = ~v_1176 | v_18;
assign x_4661 = ~v_1173 | ~v_92 | ~v_6 | v_8;
assign x_4662 = ~v_1174 | ~v_17;
assign x_4663 = ~v_1174 | v_19;
assign x_4664 = ~v_1171 | ~v_93 | ~v_6 | v_9;
assign x_4665 = ~v_1172 | ~v_17;
assign x_4666 = ~v_1172 | v_20;
assign x_4667 = ~v_1169 | ~v_94 | ~v_6 | v_10;
assign x_4668 = ~v_1170 | ~v_17;
assign x_4669 = ~v_1170 | v_21;
assign x_4670 = ~v_1167 | ~v_95 | ~v_7 | v_8;
assign x_4671 = ~v_1168 | ~v_18;
assign x_4672 = ~v_1168 | v_19;
assign x_4673 = ~v_1165 | ~v_96 | ~v_7 | v_9;
assign x_4674 = ~v_1166 | ~v_18;
assign x_4675 = ~v_1166 | v_20;
assign x_4676 = ~v_1163 | ~v_97 | ~v_7 | v_10;
assign x_4677 = ~v_1164 | ~v_18;
assign x_4678 = ~v_1164 | v_21;
assign x_4679 = ~v_1161 | ~v_98 | ~v_8 | v_9;
assign x_4680 = ~v_1162 | ~v_19;
assign x_4681 = ~v_1162 | v_20;
assign x_4682 = ~v_1159 | ~v_99 | ~v_8 | v_10;
assign x_4683 = ~v_1160 | ~v_19;
assign x_4684 = ~v_1160 | v_21;
assign x_4685 = ~v_1157 | ~v_100 | ~v_9 | v_10;
assign x_4686 = ~v_1158 | ~v_20;
assign x_4687 = ~v_1158 | v_21;
assign x_4688 = ~v_1111 | v_12 | ~v_23;
assign x_4689 = ~v_1111 | ~v_12 | v_23 | v_3552 | v_3551 | v_3550 | v_3549 | v_3548 | v_3547 | v_3546 | v_3545 | v_3544;
assign x_4690 = ~v_1111 | ~v_3552 | v_1110;
assign x_4691 = ~v_1111 | ~v_101 | ~v_12 | v_13 | v_3552;
assign x_4692 = ~v_1111 | ~v_3551 | v_1109;
assign x_4693 = ~v_1111 | ~v_102 | ~v_12 | v_14 | v_3551;
assign x_4694 = ~v_1111 | ~v_3550 | v_1108;
assign x_4695 = ~v_1111 | ~v_103 | ~v_12 | v_15 | v_3550;
assign x_4696 = ~v_1111 | ~v_3549 | v_1107;
assign x_4697 = ~v_1111 | ~v_104 | ~v_12 | v_16 | v_3549;
assign x_4698 = ~v_1111 | ~v_3548 | v_1106;
assign x_4699 = ~v_1111 | ~v_105 | ~v_12 | v_17 | v_3548;
assign x_4700 = ~v_1111 | ~v_3547 | v_1105;
assign x_4701 = ~v_1111 | ~v_106 | ~v_12 | v_18 | v_3547;
assign x_4702 = ~v_1111 | ~v_3546 | v_1104;
assign x_4703 = ~v_1111 | ~v_107 | ~v_12 | v_19 | v_3546;
assign x_4704 = ~v_1111 | ~v_3545 | v_1103;
assign x_4705 = ~v_1111 | ~v_108 | ~v_12 | v_20 | v_3545;
assign x_4706 = ~v_1111 | ~v_3544 | v_1102;
assign x_4707 = ~v_1111 | ~v_109 | ~v_12 | v_21 | v_3544;
assign x_4708 = ~v_1111 | v_13 | ~v_24 | v_3553;
assign x_4709 = ~v_1111 | ~v_13 | v_24 | v_3561 | v_3560 | v_3559 | v_3558 | v_3557 | v_3556 | v_3555 | v_3554;
assign x_4710 = ~v_1111 | ~v_3553 | v_1101;
assign x_4711 = ~v_1111 | ~v_101 | ~v_12 | v_13 | v_3553;
assign x_4712 = ~v_1111 | ~v_3561 | v_1100;
assign x_4713 = ~v_1111 | ~v_110 | ~v_13 | v_14 | v_3561;
assign x_4714 = ~v_1111 | ~v_3560 | v_1099;
assign x_4715 = ~v_1111 | ~v_111 | ~v_13 | v_15 | v_3560;
assign x_4716 = ~v_1111 | ~v_3559 | v_1098;
assign x_4717 = ~v_1111 | ~v_112 | ~v_13 | v_16 | v_3559;
assign x_4718 = ~v_1111 | ~v_3558 | v_1097;
assign x_4719 = ~v_1111 | ~v_113 | ~v_13 | v_17 | v_3558;
assign x_4720 = ~v_1111 | ~v_3557 | v_1096;
assign x_4721 = ~v_1111 | ~v_114 | ~v_13 | v_18 | v_3557;
assign x_4722 = ~v_1111 | ~v_3556 | v_1095;
assign x_4723 = ~v_1111 | ~v_115 | ~v_13 | v_19 | v_3556;
assign x_4724 = ~v_1111 | ~v_3555 | v_1094;
assign x_4725 = ~v_1111 | ~v_116 | ~v_13 | v_20 | v_3555;
assign x_4726 = ~v_1111 | ~v_3554 | v_1093;
assign x_4727 = ~v_1111 | ~v_117 | ~v_13 | v_21 | v_3554;
assign x_4728 = ~v_1111 | v_14 | ~v_25 | v_3563 | v_3562;
assign x_4729 = ~v_1111 | ~v_14 | v_25 | v_3570 | v_3569 | v_3568 | v_3567 | v_3566 | v_3565 | v_3564;
assign x_4730 = ~v_1111 | ~v_3563 | v_1092;
assign x_4731 = ~v_1111 | ~v_102 | ~v_12 | v_14 | v_3563;
assign x_4732 = ~v_1111 | ~v_3562 | v_1091;
assign x_4733 = ~v_1111 | ~v_110 | ~v_13 | v_14 | v_3562;
assign x_4734 = ~v_1111 | ~v_3570 | v_1090;
assign x_4735 = ~v_1111 | ~v_118 | ~v_14 | v_15 | v_3570;
assign x_4736 = ~v_1111 | ~v_3569 | v_1089;
assign x_4737 = ~v_1111 | ~v_119 | ~v_14 | v_16 | v_3569;
assign x_4738 = ~v_1111 | ~v_3568 | v_1088;
assign x_4739 = ~v_1111 | ~v_120 | ~v_14 | v_17 | v_3568;
assign x_4740 = ~v_1111 | ~v_3567 | v_1087;
assign x_4741 = ~v_1111 | ~v_121 | ~v_14 | v_18 | v_3567;
assign x_4742 = ~v_1111 | ~v_3566 | v_1086;
assign x_4743 = ~v_1111 | ~v_122 | ~v_14 | v_19 | v_3566;
assign x_4744 = ~v_1111 | ~v_3565 | v_1085;
assign x_4745 = ~v_1111 | ~v_123 | ~v_14 | v_20 | v_3565;
assign x_4746 = ~v_1111 | ~v_3564 | v_1084;
assign x_4747 = ~v_1111 | ~v_124 | ~v_14 | v_21 | v_3564;
assign x_4748 = ~v_1111 | v_15 | ~v_26 | v_3573 | v_3572 | v_3571;
assign x_4749 = ~v_1111 | ~v_15 | v_26 | v_3579 | v_3578 | v_3577 | v_3576 | v_3575 | v_3574;
assign x_4750 = ~v_1111 | ~v_3573 | v_1083;
assign x_4751 = ~v_1111 | ~v_103 | ~v_12 | v_15 | v_3573;
assign x_4752 = ~v_1111 | ~v_3572 | v_1082;
assign x_4753 = ~v_1111 | ~v_111 | ~v_13 | v_15 | v_3572;
assign x_4754 = ~v_1111 | ~v_3571 | v_1081;
assign x_4755 = ~v_1111 | ~v_118 | ~v_14 | v_15 | v_3571;
assign x_4756 = ~v_1111 | ~v_3579 | v_1080;
assign x_4757 = ~v_1111 | ~v_125 | ~v_15 | v_16 | v_3579;
assign x_4758 = ~v_1111 | ~v_3578 | v_1079;
assign x_4759 = ~v_1111 | ~v_126 | ~v_15 | v_17 | v_3578;
assign x_4760 = ~v_1111 | ~v_3577 | v_1078;
assign x_4761 = ~v_1111 | ~v_127 | ~v_15 | v_18 | v_3577;
assign x_4762 = ~v_1111 | ~v_3576 | v_1077;
assign x_4763 = ~v_1111 | ~v_128 | ~v_15 | v_19 | v_3576;
assign x_4764 = ~v_1111 | ~v_3575 | v_1076;
assign x_4765 = ~v_1111 | ~v_129 | ~v_15 | v_20 | v_3575;
assign x_4766 = ~v_1111 | ~v_3574 | v_1075;
assign x_4767 = ~v_1111 | ~v_130 | ~v_15 | v_21 | v_3574;
assign x_4768 = ~v_1111 | v_16 | ~v_27 | v_3583 | v_3582 | v_3581 | v_3580;
assign x_4769 = ~v_1111 | ~v_16 | v_27 | v_3588 | v_3587 | v_3586 | v_3585 | v_3584;
assign x_4770 = ~v_1111 | ~v_3583 | v_1074;
assign x_4771 = ~v_1111 | ~v_104 | ~v_12 | v_16 | v_3583;
assign x_4772 = ~v_1111 | ~v_3582 | v_1073;
assign x_4773 = ~v_1111 | ~v_112 | ~v_13 | v_16 | v_3582;
assign x_4774 = ~v_1111 | ~v_3581 | v_1072;
assign x_4775 = ~v_1111 | ~v_119 | ~v_14 | v_16 | v_3581;
assign x_4776 = ~v_1111 | ~v_3580 | v_1071;
assign x_4777 = ~v_1111 | ~v_125 | ~v_15 | v_16 | v_3580;
assign x_4778 = ~v_1111 | ~v_3588 | v_1070;
assign x_4779 = ~v_1111 | ~v_131 | ~v_16 | v_17 | v_3588;
assign x_4780 = ~v_1111 | ~v_3587 | v_1069;
assign x_4781 = ~v_1111 | ~v_132 | ~v_16 | v_18 | v_3587;
assign x_4782 = ~v_1111 | ~v_3586 | v_1068;
assign x_4783 = ~v_1111 | ~v_133 | ~v_16 | v_19 | v_3586;
assign x_4784 = ~v_1111 | ~v_3585 | v_1067;
assign x_4785 = ~v_1111 | ~v_134 | ~v_16 | v_20 | v_3585;
assign x_4786 = ~v_1111 | ~v_3584 | v_1066;
assign x_4787 = ~v_1111 | ~v_135 | ~v_16 | v_21 | v_3584;
assign x_4788 = ~v_1111 | v_17 | ~v_28 | v_3593 | v_3592 | v_3591 | v_3590 | v_3589;
assign x_4789 = ~v_1111 | ~v_17 | v_28 | v_3597 | v_3596 | v_3595 | v_3594;
assign x_4790 = ~v_1111 | ~v_3593 | v_1065;
assign x_4791 = ~v_1111 | ~v_105 | ~v_12 | v_17 | v_3593;
assign x_4792 = ~v_1111 | ~v_3592 | v_1064;
assign x_4793 = ~v_1111 | ~v_113 | ~v_13 | v_17 | v_3592;
assign x_4794 = ~v_1111 | ~v_3591 | v_1063;
assign x_4795 = ~v_1111 | ~v_120 | ~v_14 | v_17 | v_3591;
assign x_4796 = ~v_1111 | ~v_3590 | v_1062;
assign x_4797 = ~v_1111 | ~v_126 | ~v_15 | v_17 | v_3590;
assign x_4798 = ~v_1111 | ~v_3589 | v_1061;
assign x_4799 = ~v_1111 | ~v_131 | ~v_16 | v_17 | v_3589;
assign x_4800 = ~v_1111 | ~v_3597 | v_1060;
assign x_4801 = ~v_1111 | ~v_136 | ~v_17 | v_18 | v_3597;
assign x_4802 = ~v_1111 | ~v_3596 | v_1059;
assign x_4803 = ~v_1111 | ~v_137 | ~v_17 | v_19 | v_3596;
assign x_4804 = ~v_1111 | ~v_3595 | v_1058;
assign x_4805 = ~v_1111 | ~v_138 | ~v_17 | v_20 | v_3595;
assign x_4806 = ~v_1111 | ~v_3594 | v_1057;
assign x_4807 = ~v_1111 | ~v_139 | ~v_17 | v_21 | v_3594;
assign x_4808 = ~v_1111 | v_18 | ~v_29 | v_3603 | v_3602 | v_3601 | v_3600 | v_3599 | v_3598;
assign x_4809 = ~v_1111 | ~v_18 | v_29 | v_3606 | v_3605 | v_3604;
assign x_4810 = ~v_1111 | ~v_3603 | v_1056;
assign x_4811 = ~v_1111 | ~v_106 | ~v_12 | v_18 | v_3603;
assign x_4812 = ~v_1111 | ~v_3602 | v_1055;
assign x_4813 = ~v_1111 | ~v_114 | ~v_13 | v_18 | v_3602;
assign x_4814 = ~v_1111 | ~v_3601 | v_1054;
assign x_4815 = ~v_1111 | ~v_121 | ~v_14 | v_18 | v_3601;
assign x_4816 = ~v_1111 | ~v_3600 | v_1053;
assign x_4817 = ~v_1111 | ~v_127 | ~v_15 | v_18 | v_3600;
assign x_4818 = ~v_1111 | ~v_3599 | v_1052;
assign x_4819 = ~v_1111 | ~v_132 | ~v_16 | v_18 | v_3599;
assign x_4820 = ~v_1111 | ~v_3598 | v_1051;
assign x_4821 = ~v_1111 | ~v_136 | ~v_17 | v_18 | v_3598;
assign x_4822 = ~v_1111 | ~v_3606 | v_1050;
assign x_4823 = ~v_1111 | ~v_140 | ~v_18 | v_19 | v_3606;
assign x_4824 = ~v_1111 | ~v_3605 | v_1049;
assign x_4825 = ~v_1111 | ~v_141 | ~v_18 | v_20 | v_3605;
assign x_4826 = ~v_1111 | ~v_3604 | v_1048;
assign x_4827 = ~v_1111 | ~v_142 | ~v_18 | v_21 | v_3604;
assign x_4828 = ~v_1111 | v_19 | ~v_30 | v_3613 | v_3612 | v_3611 | v_3610 | v_3609 | v_3608 | v_3607;
assign x_4829 = ~v_1111 | ~v_19 | v_30 | v_3615 | v_3614;
assign x_4830 = ~v_1111 | ~v_3613 | v_1047;
assign x_4831 = ~v_1111 | ~v_107 | ~v_12 | v_19 | v_3613;
assign x_4832 = ~v_1111 | ~v_3612 | v_1046;
assign x_4833 = ~v_1111 | ~v_115 | ~v_13 | v_19 | v_3612;
assign x_4834 = ~v_1111 | ~v_3611 | v_1045;
assign x_4835 = ~v_1111 | ~v_122 | ~v_14 | v_19 | v_3611;
assign x_4836 = ~v_1111 | ~v_3610 | v_1044;
assign x_4837 = ~v_1111 | ~v_128 | ~v_15 | v_19 | v_3610;
assign x_4838 = ~v_1111 | ~v_3609 | v_1043;
assign x_4839 = ~v_1111 | ~v_133 | ~v_16 | v_19 | v_3609;
assign x_4840 = ~v_1111 | ~v_3608 | v_1042;
assign x_4841 = ~v_1111 | ~v_137 | ~v_17 | v_19 | v_3608;
assign x_4842 = ~v_1111 | ~v_3607 | v_1041;
assign x_4843 = ~v_1111 | ~v_140 | ~v_18 | v_19 | v_3607;
assign x_4844 = ~v_1111 | ~v_3615 | v_1040;
assign x_4845 = ~v_1111 | ~v_143 | ~v_19 | v_20 | v_3615;
assign x_4846 = ~v_1111 | ~v_3614 | v_1039;
assign x_4847 = ~v_1111 | ~v_144 | ~v_19 | v_21 | v_3614;
assign x_4848 = ~v_1111 | v_20 | ~v_31 | v_3623 | v_3622 | v_3621 | v_3620 | v_3619 | v_3618 | v_3617 | v_3616;
assign x_4849 = ~v_1111 | ~v_20 | v_31 | v_3624;
assign x_4850 = ~v_1111 | ~v_3623 | v_1038;
assign x_4851 = ~v_1111 | ~v_108 | ~v_12 | v_20 | v_3623;
assign x_4852 = ~v_1111 | ~v_3622 | v_1037;
assign x_4853 = ~v_1111 | ~v_116 | ~v_13 | v_20 | v_3622;
assign x_4854 = ~v_1111 | ~v_3621 | v_1036;
assign x_4855 = ~v_1111 | ~v_123 | ~v_14 | v_20 | v_3621;
assign x_4856 = ~v_1111 | ~v_3620 | v_1035;
assign x_4857 = ~v_1111 | ~v_129 | ~v_15 | v_20 | v_3620;
assign x_4858 = ~v_1111 | ~v_3619 | v_1034;
assign x_4859 = ~v_1111 | ~v_134 | ~v_16 | v_20 | v_3619;
assign x_4860 = ~v_1111 | ~v_3618 | v_1033;
assign x_4861 = ~v_1111 | ~v_138 | ~v_17 | v_20 | v_3618;
assign x_4862 = ~v_1111 | ~v_3617 | v_1032;
assign x_4863 = ~v_1111 | ~v_141 | ~v_18 | v_20 | v_3617;
assign x_4864 = ~v_1111 | ~v_3616 | v_1031;
assign x_4865 = ~v_1111 | ~v_143 | ~v_19 | v_20 | v_3616;
assign x_4866 = ~v_1111 | ~v_3624 | v_1030;
assign x_4867 = ~v_1111 | ~v_145 | ~v_20 | v_21 | v_3624;
assign x_4868 = ~v_1111 | v_21 | ~v_32 | v_3633 | v_3632 | v_3631 | v_3630 | v_3629 | v_3628 | v_3627 | v_3626 | v_3625;
assign x_4869 = ~v_1111 | ~v_21 | v_32;
assign x_4870 = ~v_1111 | ~v_3633 | v_1029;
assign x_4871 = ~v_1111 | ~v_109 | ~v_12 | v_21 | v_3633;
assign x_4872 = ~v_1111 | ~v_3632 | v_1028;
assign x_4873 = ~v_1111 | ~v_117 | ~v_13 | v_21 | v_3632;
assign x_4874 = ~v_1111 | ~v_3631 | v_1027;
assign x_4875 = ~v_1111 | ~v_124 | ~v_14 | v_21 | v_3631;
assign x_4876 = ~v_1111 | ~v_3630 | v_1026;
assign x_4877 = ~v_1111 | ~v_130 | ~v_15 | v_21 | v_3630;
assign x_4878 = ~v_1111 | ~v_3629 | v_1025;
assign x_4879 = ~v_1111 | ~v_135 | ~v_16 | v_21 | v_3629;
assign x_4880 = ~v_1111 | ~v_3628 | v_1024;
assign x_4881 = ~v_1111 | ~v_139 | ~v_17 | v_21 | v_3628;
assign x_4882 = ~v_1111 | ~v_3627 | v_1023;
assign x_4883 = ~v_1111 | ~v_142 | ~v_18 | v_21 | v_3627;
assign x_4884 = ~v_1111 | ~v_3626 | v_1022;
assign x_4885 = ~v_1111 | ~v_144 | ~v_19 | v_21 | v_3626;
assign x_4886 = ~v_1111 | ~v_3625 | v_1021;
assign x_4887 = ~v_1111 | ~v_145 | ~v_20 | v_21 | v_3625;
assign x_4888 = ~v_1111 | v_22 | ~v_33;
assign x_4889 = ~v_1111 | ~v_22 | v_33;
assign x_4890 = ~v_1111 | v_1019 | v_1020;
assign x_4891 = ~v_1111 | v_1017 | v_1018;
assign x_4892 = ~v_1111 | v_1015 | v_1016;
assign x_4893 = ~v_1111 | v_1013 | v_1014;
assign x_4894 = ~v_1111 | v_1011 | v_1012;
assign x_4895 = ~v_1111 | v_1009 | v_1010;
assign x_4896 = ~v_1111 | v_1007 | v_1008;
assign x_4897 = ~v_1111 | v_1005 | v_1006;
assign x_4898 = ~v_1111 | v_1003 | v_1004;
assign x_4899 = ~v_1111 | v_1001 | v_1002;
assign x_4900 = ~v_1111 | v_999 | v_1000;
assign x_4901 = ~v_1111 | v_997 | v_998;
assign x_4902 = ~v_1111 | v_995 | v_996;
assign x_4903 = ~v_1111 | v_993 | v_994;
assign x_4904 = ~v_1111 | v_991 | v_992;
assign x_4905 = ~v_1111 | v_989 | v_990;
assign x_4906 = ~v_1111 | v_987 | v_988;
assign x_4907 = ~v_1111 | v_985 | v_986;
assign x_4908 = ~v_1111 | v_983 | v_984;
assign x_4909 = ~v_1111 | v_981 | v_982;
assign x_4910 = ~v_1111 | v_979 | v_980;
assign x_4911 = ~v_1111 | v_977 | v_978;
assign x_4912 = ~v_1111 | v_975 | v_976;
assign x_4913 = ~v_1111 | v_973 | v_974;
assign x_4914 = ~v_1111 | v_971 | v_972;
assign x_4915 = ~v_1111 | v_969 | v_970;
assign x_4916 = ~v_1111 | v_967 | v_968;
assign x_4917 = ~v_1111 | v_965 | v_966;
assign x_4918 = ~v_1111 | v_963 | v_964;
assign x_4919 = ~v_1111 | v_961 | v_962;
assign x_4920 = ~v_1111 | v_959 | v_960;
assign x_4921 = ~v_1111 | v_957 | v_958;
assign x_4922 = ~v_1111 | v_955 | v_956;
assign x_4923 = ~v_1111 | v_953 | v_954;
assign x_4924 = ~v_1111 | v_951 | v_952;
assign x_4925 = ~v_1111 | v_949 | v_950;
assign x_4926 = ~v_1111 | v_947 | v_948;
assign x_4927 = ~v_1111 | v_945 | v_946;
assign x_4928 = ~v_1111 | v_943 | v_944;
assign x_4929 = ~v_1111 | v_941 | v_942;
assign x_4930 = ~v_1111 | v_939 | v_940;
assign x_4931 = ~v_1111 | v_937 | v_938;
assign x_4932 = ~v_1111 | v_935 | v_936;
assign x_4933 = ~v_1111 | v_933 | v_934;
assign x_4934 = ~v_1111 | v_931 | v_932;
assign x_4935 = ~v_1111 | v_885;
assign x_4936 = ~v_1110 | v_101;
assign x_4937 = ~v_1110 | v_12;
assign x_4938 = ~v_1110 | ~v_13;
assign x_4939 = ~v_1109 | v_102;
assign x_4940 = ~v_1109 | v_12;
assign x_4941 = ~v_1109 | ~v_14;
assign x_4942 = ~v_1108 | v_103;
assign x_4943 = ~v_1108 | v_12;
assign x_4944 = ~v_1108 | ~v_15;
assign x_4945 = ~v_1107 | v_104;
assign x_4946 = ~v_1107 | v_12;
assign x_4947 = ~v_1107 | ~v_16;
assign x_4948 = ~v_1106 | v_105;
assign x_4949 = ~v_1106 | v_12;
assign x_4950 = ~v_1106 | ~v_17;
assign x_4951 = ~v_1105 | v_106;
assign x_4952 = ~v_1105 | v_12;
assign x_4953 = ~v_1105 | ~v_18;
assign x_4954 = ~v_1104 | v_107;
assign x_4955 = ~v_1104 | v_12;
assign x_4956 = ~v_1104 | ~v_19;
assign x_4957 = ~v_1103 | v_108;
assign x_4958 = ~v_1103 | v_12;
assign x_4959 = ~v_1103 | ~v_20;
assign x_4960 = ~v_1102 | v_109;
assign x_4961 = ~v_1102 | v_12;
assign x_4962 = ~v_1102 | ~v_21;
assign x_4963 = ~v_1101 | v_101;
assign x_4964 = ~v_1101 | v_12;
assign x_4965 = ~v_1101 | ~v_13;
assign x_4966 = ~v_1100 | v_110;
assign x_4967 = ~v_1100 | v_13;
assign x_4968 = ~v_1100 | ~v_14;
assign x_4969 = ~v_1099 | v_111;
assign x_4970 = ~v_1099 | v_13;
assign x_4971 = ~v_1099 | ~v_15;
assign x_4972 = ~v_1098 | v_112;
assign x_4973 = ~v_1098 | v_13;
assign x_4974 = ~v_1098 | ~v_16;
assign x_4975 = ~v_1097 | v_113;
assign x_4976 = ~v_1097 | v_13;
assign x_4977 = ~v_1097 | ~v_17;
assign x_4978 = ~v_1096 | v_114;
assign x_4979 = ~v_1096 | v_13;
assign x_4980 = ~v_1096 | ~v_18;
assign x_4981 = ~v_1095 | v_115;
assign x_4982 = ~v_1095 | v_13;
assign x_4983 = ~v_1095 | ~v_19;
assign x_4984 = ~v_1094 | v_116;
assign x_4985 = ~v_1094 | v_13;
assign x_4986 = ~v_1094 | ~v_20;
assign x_4987 = ~v_1093 | v_117;
assign x_4988 = ~v_1093 | v_13;
assign x_4989 = ~v_1093 | ~v_21;
assign x_4990 = ~v_1092 | v_102;
assign x_4991 = ~v_1092 | v_12;
assign x_4992 = ~v_1092 | ~v_14;
assign x_4993 = ~v_1091 | v_110;
assign x_4994 = ~v_1091 | v_13;
assign x_4995 = ~v_1091 | ~v_14;
assign x_4996 = ~v_1090 | v_118;
assign x_4997 = ~v_1090 | v_14;
assign x_4998 = ~v_1090 | ~v_15;
assign x_4999 = ~v_1089 | v_119;
assign x_5000 = ~v_1089 | v_14;
assign x_5001 = ~v_1089 | ~v_16;
assign x_5002 = ~v_1088 | v_120;
assign x_5003 = ~v_1088 | v_14;
assign x_5004 = ~v_1088 | ~v_17;
assign x_5005 = ~v_1087 | v_121;
assign x_5006 = ~v_1087 | v_14;
assign x_5007 = ~v_1087 | ~v_18;
assign x_5008 = ~v_1086 | v_122;
assign x_5009 = ~v_1086 | v_14;
assign x_5010 = ~v_1086 | ~v_19;
assign x_5011 = ~v_1085 | v_123;
assign x_5012 = ~v_1085 | v_14;
assign x_5013 = ~v_1085 | ~v_20;
assign x_5014 = ~v_1084 | v_124;
assign x_5015 = ~v_1084 | v_14;
assign x_5016 = ~v_1084 | ~v_21;
assign x_5017 = ~v_1083 | v_103;
assign x_5018 = ~v_1083 | v_12;
assign x_5019 = ~v_1083 | ~v_15;
assign x_5020 = ~v_1082 | v_111;
assign x_5021 = ~v_1082 | v_13;
assign x_5022 = ~v_1082 | ~v_15;
assign x_5023 = ~v_1081 | v_118;
assign x_5024 = ~v_1081 | v_14;
assign x_5025 = ~v_1081 | ~v_15;
assign x_5026 = ~v_1080 | v_125;
assign x_5027 = ~v_1080 | v_15;
assign x_5028 = ~v_1080 | ~v_16;
assign x_5029 = ~v_1079 | v_126;
assign x_5030 = ~v_1079 | v_15;
assign x_5031 = ~v_1079 | ~v_17;
assign x_5032 = ~v_1078 | v_127;
assign x_5033 = ~v_1078 | v_15;
assign x_5034 = ~v_1078 | ~v_18;
assign x_5035 = ~v_1077 | v_128;
assign x_5036 = ~v_1077 | v_15;
assign x_5037 = ~v_1077 | ~v_19;
assign x_5038 = ~v_1076 | v_129;
assign x_5039 = ~v_1076 | v_15;
assign x_5040 = ~v_1076 | ~v_20;
assign x_5041 = ~v_1075 | v_130;
assign x_5042 = ~v_1075 | v_15;
assign x_5043 = ~v_1075 | ~v_21;
assign x_5044 = ~v_1074 | v_104;
assign x_5045 = ~v_1074 | v_12;
assign x_5046 = ~v_1074 | ~v_16;
assign x_5047 = ~v_1073 | v_112;
assign x_5048 = ~v_1073 | v_13;
assign x_5049 = ~v_1073 | ~v_16;
assign x_5050 = ~v_1072 | v_119;
assign x_5051 = ~v_1072 | v_14;
assign x_5052 = ~v_1072 | ~v_16;
assign x_5053 = ~v_1071 | v_125;
assign x_5054 = ~v_1071 | v_15;
assign x_5055 = ~v_1071 | ~v_16;
assign x_5056 = ~v_1070 | v_131;
assign x_5057 = ~v_1070 | v_16;
assign x_5058 = ~v_1070 | ~v_17;
assign x_5059 = ~v_1069 | v_132;
assign x_5060 = ~v_1069 | v_16;
assign x_5061 = ~v_1069 | ~v_18;
assign x_5062 = ~v_1068 | v_133;
assign x_5063 = ~v_1068 | v_16;
assign x_5064 = ~v_1068 | ~v_19;
assign x_5065 = ~v_1067 | v_134;
assign x_5066 = ~v_1067 | v_16;
assign x_5067 = ~v_1067 | ~v_20;
assign x_5068 = ~v_1066 | v_135;
assign x_5069 = ~v_1066 | v_16;
assign x_5070 = ~v_1066 | ~v_21;
assign x_5071 = ~v_1065 | v_105;
assign x_5072 = ~v_1065 | v_12;
assign x_5073 = ~v_1065 | ~v_17;
assign x_5074 = ~v_1064 | v_113;
assign x_5075 = ~v_1064 | v_13;
assign x_5076 = ~v_1064 | ~v_17;
assign x_5077 = ~v_1063 | v_120;
assign x_5078 = ~v_1063 | v_14;
assign x_5079 = ~v_1063 | ~v_17;
assign x_5080 = ~v_1062 | v_126;
assign x_5081 = ~v_1062 | v_15;
assign x_5082 = ~v_1062 | ~v_17;
assign x_5083 = ~v_1061 | v_131;
assign x_5084 = ~v_1061 | v_16;
assign x_5085 = ~v_1061 | ~v_17;
assign x_5086 = ~v_1060 | v_136;
assign x_5087 = ~v_1060 | v_17;
assign x_5088 = ~v_1060 | ~v_18;
assign x_5089 = ~v_1059 | v_137;
assign x_5090 = ~v_1059 | v_17;
assign x_5091 = ~v_1059 | ~v_19;
assign x_5092 = ~v_1058 | v_138;
assign x_5093 = ~v_1058 | v_17;
assign x_5094 = ~v_1058 | ~v_20;
assign x_5095 = ~v_1057 | v_139;
assign x_5096 = ~v_1057 | v_17;
assign x_5097 = ~v_1057 | ~v_21;
assign x_5098 = ~v_1056 | v_106;
assign x_5099 = ~v_1056 | v_12;
assign x_5100 = ~v_1056 | ~v_18;
assign x_5101 = ~v_1055 | v_114;
assign x_5102 = ~v_1055 | v_13;
assign x_5103 = ~v_1055 | ~v_18;
assign x_5104 = ~v_1054 | v_121;
assign x_5105 = ~v_1054 | v_14;
assign x_5106 = ~v_1054 | ~v_18;
assign x_5107 = ~v_1053 | v_127;
assign x_5108 = ~v_1053 | v_15;
assign x_5109 = ~v_1053 | ~v_18;
assign x_5110 = ~v_1052 | v_132;
assign x_5111 = ~v_1052 | v_16;
assign x_5112 = ~v_1052 | ~v_18;
assign x_5113 = ~v_1051 | v_136;
assign x_5114 = ~v_1051 | v_17;
assign x_5115 = ~v_1051 | ~v_18;
assign x_5116 = ~v_1050 | v_140;
assign x_5117 = ~v_1050 | v_18;
assign x_5118 = ~v_1050 | ~v_19;
assign x_5119 = ~v_1049 | v_141;
assign x_5120 = ~v_1049 | v_18;
assign x_5121 = ~v_1049 | ~v_20;
assign x_5122 = ~v_1048 | v_142;
assign x_5123 = ~v_1048 | v_18;
assign x_5124 = ~v_1048 | ~v_21;
assign x_5125 = ~v_1047 | v_107;
assign x_5126 = ~v_1047 | v_12;
assign x_5127 = ~v_1047 | ~v_19;
assign x_5128 = ~v_1046 | v_115;
assign x_5129 = ~v_1046 | v_13;
assign x_5130 = ~v_1046 | ~v_19;
assign x_5131 = ~v_1045 | v_122;
assign x_5132 = ~v_1045 | v_14;
assign x_5133 = ~v_1045 | ~v_19;
assign x_5134 = ~v_1044 | v_128;
assign x_5135 = ~v_1044 | v_15;
assign x_5136 = ~v_1044 | ~v_19;
assign x_5137 = ~v_1043 | v_133;
assign x_5138 = ~v_1043 | v_16;
assign x_5139 = ~v_1043 | ~v_19;
assign x_5140 = ~v_1042 | v_137;
assign x_5141 = ~v_1042 | v_17;
assign x_5142 = ~v_1042 | ~v_19;
assign x_5143 = ~v_1041 | v_140;
assign x_5144 = ~v_1041 | v_18;
assign x_5145 = ~v_1041 | ~v_19;
assign x_5146 = ~v_1040 | v_143;
assign x_5147 = ~v_1040 | v_19;
assign x_5148 = ~v_1040 | ~v_20;
assign x_5149 = ~v_1039 | v_144;
assign x_5150 = ~v_1039 | v_19;
assign x_5151 = ~v_1039 | ~v_21;
assign x_5152 = ~v_1038 | v_108;
assign x_5153 = ~v_1038 | v_12;
assign x_5154 = ~v_1038 | ~v_20;
assign x_5155 = ~v_1037 | v_116;
assign x_5156 = ~v_1037 | v_13;
assign x_5157 = ~v_1037 | ~v_20;
assign x_5158 = ~v_1036 | v_123;
assign x_5159 = ~v_1036 | v_14;
assign x_5160 = ~v_1036 | ~v_20;
assign x_5161 = ~v_1035 | v_129;
assign x_5162 = ~v_1035 | v_15;
assign x_5163 = ~v_1035 | ~v_20;
assign x_5164 = ~v_1034 | v_134;
assign x_5165 = ~v_1034 | v_16;
assign x_5166 = ~v_1034 | ~v_20;
assign x_5167 = ~v_1033 | v_138;
assign x_5168 = ~v_1033 | v_17;
assign x_5169 = ~v_1033 | ~v_20;
assign x_5170 = ~v_1032 | v_141;
assign x_5171 = ~v_1032 | v_18;
assign x_5172 = ~v_1032 | ~v_20;
assign x_5173 = ~v_1031 | v_143;
assign x_5174 = ~v_1031 | v_19;
assign x_5175 = ~v_1031 | ~v_20;
assign x_5176 = ~v_1030 | v_145;
assign x_5177 = ~v_1030 | v_20;
assign x_5178 = ~v_1030 | ~v_21;
assign x_5179 = ~v_1029 | v_109;
assign x_5180 = ~v_1029 | v_12;
assign x_5181 = ~v_1029 | ~v_21;
assign x_5182 = ~v_1028 | v_117;
assign x_5183 = ~v_1028 | v_13;
assign x_5184 = ~v_1028 | ~v_21;
assign x_5185 = ~v_1027 | v_124;
assign x_5186 = ~v_1027 | v_14;
assign x_5187 = ~v_1027 | ~v_21;
assign x_5188 = ~v_1026 | v_130;
assign x_5189 = ~v_1026 | v_15;
assign x_5190 = ~v_1026 | ~v_21;
assign x_5191 = ~v_1025 | v_135;
assign x_5192 = ~v_1025 | v_16;
assign x_5193 = ~v_1025 | ~v_21;
assign x_5194 = ~v_1024 | v_139;
assign x_5195 = ~v_1024 | v_17;
assign x_5196 = ~v_1024 | ~v_21;
assign x_5197 = ~v_1023 | v_142;
assign x_5198 = ~v_1023 | v_18;
assign x_5199 = ~v_1023 | ~v_21;
assign x_5200 = ~v_1022 | v_144;
assign x_5201 = ~v_1022 | v_19;
assign x_5202 = ~v_1022 | ~v_21;
assign x_5203 = ~v_1021 | v_145;
assign x_5204 = ~v_1021 | v_20;
assign x_5205 = ~v_1021 | ~v_21;
assign x_5206 = ~v_1019 | ~v_101 | ~v_12 | v_13;
assign x_5207 = ~v_1020 | ~v_23;
assign x_5208 = ~v_1020 | v_24;
assign x_5209 = ~v_1017 | ~v_102 | ~v_12 | v_14;
assign x_5210 = ~v_1018 | ~v_23;
assign x_5211 = ~v_1018 | v_25;
assign x_5212 = ~v_1015 | ~v_103 | ~v_12 | v_15;
assign x_5213 = ~v_1016 | ~v_23;
assign x_5214 = ~v_1016 | v_26;
assign x_5215 = ~v_1013 | ~v_104 | ~v_12 | v_16;
assign x_5216 = ~v_1014 | ~v_23;
assign x_5217 = ~v_1014 | v_27;
assign x_5218 = ~v_1011 | ~v_105 | ~v_12 | v_17;
assign x_5219 = ~v_1012 | ~v_23;
assign x_5220 = ~v_1012 | v_28;
assign x_5221 = ~v_1009 | ~v_106 | ~v_12 | v_18;
assign x_5222 = ~v_1010 | ~v_23;
assign x_5223 = ~v_1010 | v_29;
assign x_5224 = ~v_1007 | ~v_107 | ~v_12 | v_19;
assign x_5225 = ~v_1008 | ~v_23;
assign x_5226 = ~v_1008 | v_30;
assign x_5227 = ~v_1005 | ~v_108 | ~v_12 | v_20;
assign x_5228 = ~v_1006 | ~v_23;
assign x_5229 = ~v_1006 | v_31;
assign x_5230 = ~v_1003 | ~v_109 | ~v_12 | v_21;
assign x_5231 = ~v_1004 | ~v_23;
assign x_5232 = ~v_1004 | v_32;
assign x_5233 = ~v_1001 | ~v_110 | ~v_13 | v_14;
assign x_5234 = ~v_1002 | ~v_24;
assign x_5235 = ~v_1002 | v_25;
assign x_5236 = ~v_999 | ~v_111 | ~v_13 | v_15;
assign x_5237 = ~v_1000 | ~v_24;
assign x_5238 = ~v_1000 | v_26;
assign x_5239 = ~v_997 | ~v_112 | ~v_13 | v_16;
assign x_5240 = ~v_998 | ~v_24;
assign x_5241 = ~v_998 | v_27;
assign x_5242 = ~v_995 | ~v_113 | ~v_13 | v_17;
assign x_5243 = ~v_996 | ~v_24;
assign x_5244 = ~v_996 | v_28;
assign x_5245 = ~v_993 | ~v_114 | ~v_13 | v_18;
assign x_5246 = ~v_994 | ~v_24;
assign x_5247 = ~v_994 | v_29;
assign x_5248 = ~v_991 | ~v_115 | ~v_13 | v_19;
assign x_5249 = ~v_992 | ~v_24;
assign x_5250 = ~v_992 | v_30;
assign x_5251 = ~v_989 | ~v_116 | ~v_13 | v_20;
assign x_5252 = ~v_990 | ~v_24;
assign x_5253 = ~v_990 | v_31;
assign x_5254 = ~v_987 | ~v_117 | ~v_13 | v_21;
assign x_5255 = ~v_988 | ~v_24;
assign x_5256 = ~v_988 | v_32;
assign x_5257 = ~v_985 | ~v_118 | ~v_14 | v_15;
assign x_5258 = ~v_986 | ~v_25;
assign x_5259 = ~v_986 | v_26;
assign x_5260 = ~v_983 | ~v_119 | ~v_14 | v_16;
assign x_5261 = ~v_984 | ~v_25;
assign x_5262 = ~v_984 | v_27;
assign x_5263 = ~v_981 | ~v_120 | ~v_14 | v_17;
assign x_5264 = ~v_982 | ~v_25;
assign x_5265 = ~v_982 | v_28;
assign x_5266 = ~v_979 | ~v_121 | ~v_14 | v_18;
assign x_5267 = ~v_980 | ~v_25;
assign x_5268 = ~v_980 | v_29;
assign x_5269 = ~v_977 | ~v_122 | ~v_14 | v_19;
assign x_5270 = ~v_978 | ~v_25;
assign x_5271 = ~v_978 | v_30;
assign x_5272 = ~v_975 | ~v_123 | ~v_14 | v_20;
assign x_5273 = ~v_976 | ~v_25;
assign x_5274 = ~v_976 | v_31;
assign x_5275 = ~v_973 | ~v_124 | ~v_14 | v_21;
assign x_5276 = ~v_974 | ~v_25;
assign x_5277 = ~v_974 | v_32;
assign x_5278 = ~v_971 | ~v_125 | ~v_15 | v_16;
assign x_5279 = ~v_972 | ~v_26;
assign x_5280 = ~v_972 | v_27;
assign x_5281 = ~v_969 | ~v_126 | ~v_15 | v_17;
assign x_5282 = ~v_970 | ~v_26;
assign x_5283 = ~v_970 | v_28;
assign x_5284 = ~v_967 | ~v_127 | ~v_15 | v_18;
assign x_5285 = ~v_968 | ~v_26;
assign x_5286 = ~v_968 | v_29;
assign x_5287 = ~v_965 | ~v_128 | ~v_15 | v_19;
assign x_5288 = ~v_966 | ~v_26;
assign x_5289 = ~v_966 | v_30;
assign x_5290 = ~v_963 | ~v_129 | ~v_15 | v_20;
assign x_5291 = ~v_964 | ~v_26;
assign x_5292 = ~v_964 | v_31;
assign x_5293 = ~v_961 | ~v_130 | ~v_15 | v_21;
assign x_5294 = ~v_962 | ~v_26;
assign x_5295 = ~v_962 | v_32;
assign x_5296 = ~v_959 | ~v_131 | ~v_16 | v_17;
assign x_5297 = ~v_960 | ~v_27;
assign x_5298 = ~v_960 | v_28;
assign x_5299 = ~v_957 | ~v_132 | ~v_16 | v_18;
assign x_5300 = ~v_958 | ~v_27;
assign x_5301 = ~v_958 | v_29;
assign x_5302 = ~v_955 | ~v_133 | ~v_16 | v_19;
assign x_5303 = ~v_956 | ~v_27;
assign x_5304 = ~v_956 | v_30;
assign x_5305 = ~v_953 | ~v_134 | ~v_16 | v_20;
assign x_5306 = ~v_954 | ~v_27;
assign x_5307 = ~v_954 | v_31;
assign x_5308 = ~v_951 | ~v_135 | ~v_16 | v_21;
assign x_5309 = ~v_952 | ~v_27;
assign x_5310 = ~v_952 | v_32;
assign x_5311 = ~v_949 | ~v_136 | ~v_17 | v_18;
assign x_5312 = ~v_950 | ~v_28;
assign x_5313 = ~v_950 | v_29;
assign x_5314 = ~v_947 | ~v_137 | ~v_17 | v_19;
assign x_5315 = ~v_948 | ~v_28;
assign x_5316 = ~v_948 | v_30;
assign x_5317 = ~v_945 | ~v_138 | ~v_17 | v_20;
assign x_5318 = ~v_946 | ~v_28;
assign x_5319 = ~v_946 | v_31;
assign x_5320 = ~v_943 | ~v_139 | ~v_17 | v_21;
assign x_5321 = ~v_944 | ~v_28;
assign x_5322 = ~v_944 | v_32;
assign x_5323 = ~v_941 | ~v_140 | ~v_18 | v_19;
assign x_5324 = ~v_942 | ~v_29;
assign x_5325 = ~v_942 | v_30;
assign x_5326 = ~v_939 | ~v_141 | ~v_18 | v_20;
assign x_5327 = ~v_940 | ~v_29;
assign x_5328 = ~v_940 | v_31;
assign x_5329 = ~v_937 | ~v_142 | ~v_18 | v_21;
assign x_5330 = ~v_938 | ~v_29;
assign x_5331 = ~v_938 | v_32;
assign x_5332 = ~v_935 | ~v_143 | ~v_19 | v_20;
assign x_5333 = ~v_936 | ~v_30;
assign x_5334 = ~v_936 | v_31;
assign x_5335 = ~v_933 | ~v_144 | ~v_19 | v_21;
assign x_5336 = ~v_934 | ~v_30;
assign x_5337 = ~v_934 | v_32;
assign x_5338 = ~v_931 | ~v_145 | ~v_20 | v_21;
assign x_5339 = ~v_932 | ~v_31;
assign x_5340 = ~v_932 | v_32;
assign x_5341 = ~v_885 | v_23 | ~v_34;
assign x_5342 = ~v_885 | ~v_23 | v_34 | v_3786 | v_3785 | v_3784 | v_3783 | v_3782 | v_3781 | v_3780 | v_3779 | v_3778;
assign x_5343 = ~v_885 | ~v_3786 | v_884;
assign x_5344 = ~v_885 | ~v_146 | ~v_23 | v_24 | v_3786;
assign x_5345 = ~v_885 | ~v_3785 | v_883;
assign x_5346 = ~v_885 | ~v_147 | ~v_23 | v_25 | v_3785;
assign x_5347 = ~v_885 | ~v_3784 | v_882;
assign x_5348 = ~v_885 | ~v_148 | ~v_23 | v_26 | v_3784;
assign x_5349 = ~v_885 | ~v_3783 | v_881;
assign x_5350 = ~v_885 | ~v_149 | ~v_23 | v_27 | v_3783;
assign x_5351 = ~v_885 | ~v_3782 | v_880;
assign x_5352 = ~v_885 | ~v_150 | ~v_23 | v_28 | v_3782;
assign x_5353 = ~v_885 | ~v_3781 | v_879;
assign x_5354 = ~v_885 | ~v_151 | ~v_23 | v_29 | v_3781;
assign x_5355 = ~v_885 | ~v_3780 | v_878;
assign x_5356 = ~v_885 | ~v_152 | ~v_23 | v_30 | v_3780;
assign x_5357 = ~v_885 | ~v_3779 | v_877;
assign x_5358 = ~v_885 | ~v_153 | ~v_23 | v_31 | v_3779;
assign x_5359 = ~v_885 | ~v_3778 | v_876;
assign x_5360 = ~v_885 | ~v_154 | ~v_23 | v_32 | v_3778;
assign x_5361 = ~v_885 | v_24 | ~v_35 | v_3787;
assign x_5362 = ~v_885 | ~v_24 | v_35 | v_3795 | v_3794 | v_3793 | v_3792 | v_3791 | v_3790 | v_3789 | v_3788;
assign x_5363 = ~v_885 | ~v_3787 | v_875;
assign x_5364 = ~v_885 | ~v_146 | ~v_23 | v_24 | v_3787;
assign x_5365 = ~v_885 | ~v_3795 | v_874;
assign x_5366 = ~v_885 | ~v_155 | ~v_24 | v_25 | v_3795;
assign x_5367 = ~v_885 | ~v_3794 | v_873;
assign x_5368 = ~v_885 | ~v_156 | ~v_24 | v_26 | v_3794;
assign x_5369 = ~v_885 | ~v_3793 | v_872;
assign x_5370 = ~v_885 | ~v_157 | ~v_24 | v_27 | v_3793;
assign x_5371 = ~v_885 | ~v_3792 | v_871;
assign x_5372 = ~v_885 | ~v_158 | ~v_24 | v_28 | v_3792;
assign x_5373 = ~v_885 | ~v_3791 | v_870;
assign x_5374 = ~v_885 | ~v_159 | ~v_24 | v_29 | v_3791;
assign x_5375 = ~v_885 | ~v_3790 | v_869;
assign x_5376 = ~v_885 | ~v_160 | ~v_24 | v_30 | v_3790;
assign x_5377 = ~v_885 | ~v_3789 | v_868;
assign x_5378 = ~v_885 | ~v_161 | ~v_24 | v_31 | v_3789;
assign x_5379 = ~v_885 | ~v_3788 | v_867;
assign x_5380 = ~v_885 | ~v_162 | ~v_24 | v_32 | v_3788;
assign x_5381 = ~v_885 | v_25 | ~v_36 | v_3797 | v_3796;
assign x_5382 = ~v_885 | ~v_25 | v_36 | v_3804 | v_3803 | v_3802 | v_3801 | v_3800 | v_3799 | v_3798;
assign x_5383 = ~v_885 | ~v_3797 | v_866;
assign x_5384 = ~v_885 | ~v_147 | ~v_23 | v_25 | v_3797;
assign x_5385 = ~v_885 | ~v_3796 | v_865;
assign x_5386 = ~v_885 | ~v_155 | ~v_24 | v_25 | v_3796;
assign x_5387 = ~v_885 | ~v_3804 | v_864;
assign x_5388 = ~v_885 | ~v_163 | ~v_25 | v_26 | v_3804;
assign x_5389 = ~v_885 | ~v_3803 | v_863;
assign x_5390 = ~v_885 | ~v_164 | ~v_25 | v_27 | v_3803;
assign x_5391 = ~v_885 | ~v_3802 | v_862;
assign x_5392 = ~v_885 | ~v_165 | ~v_25 | v_28 | v_3802;
assign x_5393 = ~v_885 | ~v_3801 | v_861;
assign x_5394 = ~v_885 | ~v_166 | ~v_25 | v_29 | v_3801;
assign x_5395 = ~v_885 | ~v_3800 | v_860;
assign x_5396 = ~v_885 | ~v_167 | ~v_25 | v_30 | v_3800;
assign x_5397 = ~v_885 | ~v_3799 | v_859;
assign x_5398 = ~v_885 | ~v_168 | ~v_25 | v_31 | v_3799;
assign x_5399 = ~v_885 | ~v_3798 | v_858;
assign x_5400 = ~v_885 | ~v_169 | ~v_25 | v_32 | v_3798;
assign x_5401 = ~v_885 | v_26 | ~v_37 | v_3807 | v_3806 | v_3805;
assign x_5402 = ~v_885 | ~v_26 | v_37 | v_3813 | v_3812 | v_3811 | v_3810 | v_3809 | v_3808;
assign x_5403 = ~v_885 | ~v_3807 | v_857;
assign x_5404 = ~v_885 | ~v_148 | ~v_23 | v_26 | v_3807;
assign x_5405 = ~v_885 | ~v_3806 | v_856;
assign x_5406 = ~v_885 | ~v_156 | ~v_24 | v_26 | v_3806;
assign x_5407 = ~v_885 | ~v_3805 | v_855;
assign x_5408 = ~v_885 | ~v_163 | ~v_25 | v_26 | v_3805;
assign x_5409 = ~v_885 | ~v_3813 | v_854;
assign x_5410 = ~v_885 | ~v_170 | ~v_26 | v_27 | v_3813;
assign x_5411 = ~v_885 | ~v_3812 | v_853;
assign x_5412 = ~v_885 | ~v_171 | ~v_26 | v_28 | v_3812;
assign x_5413 = ~v_885 | ~v_3811 | v_852;
assign x_5414 = ~v_885 | ~v_172 | ~v_26 | v_29 | v_3811;
assign x_5415 = ~v_885 | ~v_3810 | v_851;
assign x_5416 = ~v_885 | ~v_173 | ~v_26 | v_30 | v_3810;
assign x_5417 = ~v_885 | ~v_3809 | v_850;
assign x_5418 = ~v_885 | ~v_174 | ~v_26 | v_31 | v_3809;
assign x_5419 = ~v_885 | ~v_3808 | v_849;
assign x_5420 = ~v_885 | ~v_175 | ~v_26 | v_32 | v_3808;
assign x_5421 = ~v_885 | v_27 | ~v_38 | v_3817 | v_3816 | v_3815 | v_3814;
assign x_5422 = ~v_885 | ~v_27 | v_38 | v_3822 | v_3821 | v_3820 | v_3819 | v_3818;
assign x_5423 = ~v_885 | ~v_3817 | v_848;
assign x_5424 = ~v_885 | ~v_149 | ~v_23 | v_27 | v_3817;
assign x_5425 = ~v_885 | ~v_3816 | v_847;
assign x_5426 = ~v_885 | ~v_157 | ~v_24 | v_27 | v_3816;
assign x_5427 = ~v_885 | ~v_3815 | v_846;
assign x_5428 = ~v_885 | ~v_164 | ~v_25 | v_27 | v_3815;
assign x_5429 = ~v_885 | ~v_3814 | v_845;
assign x_5430 = ~v_885 | ~v_170 | ~v_26 | v_27 | v_3814;
assign x_5431 = ~v_885 | ~v_3822 | v_844;
assign x_5432 = ~v_885 | ~v_176 | ~v_27 | v_28 | v_3822;
assign x_5433 = ~v_885 | ~v_3821 | v_843;
assign x_5434 = ~v_885 | ~v_177 | ~v_27 | v_29 | v_3821;
assign x_5435 = ~v_885 | ~v_3820 | v_842;
assign x_5436 = ~v_885 | ~v_178 | ~v_27 | v_30 | v_3820;
assign x_5437 = ~v_885 | ~v_3819 | v_841;
assign x_5438 = ~v_885 | ~v_179 | ~v_27 | v_31 | v_3819;
assign x_5439 = ~v_885 | ~v_3818 | v_840;
assign x_5440 = ~v_885 | ~v_180 | ~v_27 | v_32 | v_3818;
assign x_5441 = ~v_885 | v_28 | ~v_39 | v_3827 | v_3826 | v_3825 | v_3824 | v_3823;
assign x_5442 = ~v_885 | ~v_28 | v_39 | v_3831 | v_3830 | v_3829 | v_3828;
assign x_5443 = ~v_885 | ~v_3827 | v_839;
assign x_5444 = ~v_885 | ~v_150 | ~v_23 | v_28 | v_3827;
assign x_5445 = ~v_885 | ~v_3826 | v_838;
assign x_5446 = ~v_885 | ~v_158 | ~v_24 | v_28 | v_3826;
assign x_5447 = ~v_885 | ~v_3825 | v_837;
assign x_5448 = ~v_885 | ~v_165 | ~v_25 | v_28 | v_3825;
assign x_5449 = ~v_885 | ~v_3824 | v_836;
assign x_5450 = ~v_885 | ~v_171 | ~v_26 | v_28 | v_3824;
assign x_5451 = ~v_885 | ~v_3823 | v_835;
assign x_5452 = ~v_885 | ~v_176 | ~v_27 | v_28 | v_3823;
assign x_5453 = ~v_885 | ~v_3831 | v_834;
assign x_5454 = ~v_885 | ~v_181 | ~v_28 | v_29 | v_3831;
assign x_5455 = ~v_885 | ~v_3830 | v_833;
assign x_5456 = ~v_885 | ~v_182 | ~v_28 | v_30 | v_3830;
assign x_5457 = ~v_885 | ~v_3829 | v_832;
assign x_5458 = ~v_885 | ~v_183 | ~v_28 | v_31 | v_3829;
assign x_5459 = ~v_885 | ~v_3828 | v_831;
assign x_5460 = ~v_885 | ~v_184 | ~v_28 | v_32 | v_3828;
assign x_5461 = ~v_885 | v_29 | ~v_40 | v_3837 | v_3836 | v_3835 | v_3834 | v_3833 | v_3832;
assign x_5462 = ~v_885 | ~v_29 | v_40 | v_3840 | v_3839 | v_3838;
assign x_5463 = ~v_885 | ~v_3837 | v_830;
assign x_5464 = ~v_885 | ~v_151 | ~v_23 | v_29 | v_3837;
assign x_5465 = ~v_885 | ~v_3836 | v_829;
assign x_5466 = ~v_885 | ~v_159 | ~v_24 | v_29 | v_3836;
assign x_5467 = ~v_885 | ~v_3835 | v_828;
assign x_5468 = ~v_885 | ~v_166 | ~v_25 | v_29 | v_3835;
assign x_5469 = ~v_885 | ~v_3834 | v_827;
assign x_5470 = ~v_885 | ~v_172 | ~v_26 | v_29 | v_3834;
assign x_5471 = ~v_885 | ~v_3833 | v_826;
assign x_5472 = ~v_885 | ~v_177 | ~v_27 | v_29 | v_3833;
assign x_5473 = ~v_885 | ~v_3832 | v_825;
assign x_5474 = ~v_885 | ~v_181 | ~v_28 | v_29 | v_3832;
assign x_5475 = ~v_885 | ~v_3840 | v_824;
assign x_5476 = ~v_885 | ~v_185 | ~v_29 | v_30 | v_3840;
assign x_5477 = ~v_885 | ~v_3839 | v_823;
assign x_5478 = ~v_885 | ~v_186 | ~v_29 | v_31 | v_3839;
assign x_5479 = ~v_885 | ~v_3838 | v_822;
assign x_5480 = ~v_885 | ~v_187 | ~v_29 | v_32 | v_3838;
assign x_5481 = ~v_885 | v_30 | ~v_41 | v_3847 | v_3846 | v_3845 | v_3844 | v_3843 | v_3842 | v_3841;
assign x_5482 = ~v_885 | ~v_30 | v_41 | v_3849 | v_3848;
assign x_5483 = ~v_885 | ~v_3847 | v_821;
assign x_5484 = ~v_885 | ~v_152 | ~v_23 | v_30 | v_3847;
assign x_5485 = ~v_885 | ~v_3846 | v_820;
assign x_5486 = ~v_885 | ~v_160 | ~v_24 | v_30 | v_3846;
assign x_5487 = ~v_885 | ~v_3845 | v_819;
assign x_5488 = ~v_885 | ~v_167 | ~v_25 | v_30 | v_3845;
assign x_5489 = ~v_885 | ~v_3844 | v_818;
assign x_5490 = ~v_885 | ~v_173 | ~v_26 | v_30 | v_3844;
assign x_5491 = ~v_885 | ~v_3843 | v_817;
assign x_5492 = ~v_885 | ~v_178 | ~v_27 | v_30 | v_3843;
assign x_5493 = ~v_885 | ~v_3842 | v_816;
assign x_5494 = ~v_885 | ~v_182 | ~v_28 | v_30 | v_3842;
assign x_5495 = ~v_885 | ~v_3841 | v_815;
assign x_5496 = ~v_885 | ~v_185 | ~v_29 | v_30 | v_3841;
assign x_5497 = ~v_885 | ~v_3849 | v_814;
assign x_5498 = ~v_885 | ~v_188 | ~v_30 | v_31 | v_3849;
assign x_5499 = ~v_885 | ~v_3848 | v_813;
assign x_5500 = ~v_885 | ~v_189 | ~v_30 | v_32 | v_3848;
assign x_5501 = ~v_885 | v_31 | ~v_42 | v_3857 | v_3856 | v_3855 | v_3854 | v_3853 | v_3852 | v_3851 | v_3850;
assign x_5502 = ~v_885 | ~v_31 | v_42 | v_3858;
assign x_5503 = ~v_885 | ~v_3857 | v_812;
assign x_5504 = ~v_885 | ~v_153 | ~v_23 | v_31 | v_3857;
assign x_5505 = ~v_885 | ~v_3856 | v_811;
assign x_5506 = ~v_885 | ~v_161 | ~v_24 | v_31 | v_3856;
assign x_5507 = ~v_885 | ~v_3855 | v_810;
assign x_5508 = ~v_885 | ~v_168 | ~v_25 | v_31 | v_3855;
assign x_5509 = ~v_885 | ~v_3854 | v_809;
assign x_5510 = ~v_885 | ~v_174 | ~v_26 | v_31 | v_3854;
assign x_5511 = ~v_885 | ~v_3853 | v_808;
assign x_5512 = ~v_885 | ~v_179 | ~v_27 | v_31 | v_3853;
assign x_5513 = ~v_885 | ~v_3852 | v_807;
assign x_5514 = ~v_885 | ~v_183 | ~v_28 | v_31 | v_3852;
assign x_5515 = ~v_885 | ~v_3851 | v_806;
assign x_5516 = ~v_885 | ~v_186 | ~v_29 | v_31 | v_3851;
assign x_5517 = ~v_885 | ~v_3850 | v_805;
assign x_5518 = ~v_885 | ~v_188 | ~v_30 | v_31 | v_3850;
assign x_5519 = ~v_885 | ~v_3858 | v_804;
assign x_5520 = ~v_885 | ~v_190 | ~v_31 | v_32 | v_3858;
assign x_5521 = ~v_885 | v_32 | ~v_43 | v_3867 | v_3866 | v_3865 | v_3864 | v_3863 | v_3862 | v_3861 | v_3860 | v_3859;
assign x_5522 = ~v_885 | ~v_32 | v_43;
assign x_5523 = ~v_885 | ~v_3867 | v_803;
assign x_5524 = ~v_885 | ~v_154 | ~v_23 | v_32 | v_3867;
assign x_5525 = ~v_885 | ~v_3866 | v_802;
assign x_5526 = ~v_885 | ~v_162 | ~v_24 | v_32 | v_3866;
assign x_5527 = ~v_885 | ~v_3865 | v_801;
assign x_5528 = ~v_885 | ~v_169 | ~v_25 | v_32 | v_3865;
assign x_5529 = ~v_885 | ~v_3864 | v_800;
assign x_5530 = ~v_885 | ~v_175 | ~v_26 | v_32 | v_3864;
assign x_5531 = ~v_885 | ~v_3863 | v_799;
assign x_5532 = ~v_885 | ~v_180 | ~v_27 | v_32 | v_3863;
assign x_5533 = ~v_885 | ~v_3862 | v_798;
assign x_5534 = ~v_885 | ~v_184 | ~v_28 | v_32 | v_3862;
assign x_5535 = ~v_885 | ~v_3861 | v_797;
assign x_5536 = ~v_885 | ~v_187 | ~v_29 | v_32 | v_3861;
assign x_5537 = ~v_885 | ~v_3860 | v_796;
assign x_5538 = ~v_885 | ~v_189 | ~v_30 | v_32 | v_3860;
assign x_5539 = ~v_885 | ~v_3859 | v_795;
assign x_5540 = ~v_885 | ~v_190 | ~v_31 | v_32 | v_3859;
assign x_5541 = ~v_885 | v_33 | ~v_44;
assign x_5542 = ~v_885 | ~v_33 | v_44;
assign x_5543 = ~v_885 | v_793 | v_794;
assign x_5544 = ~v_885 | v_791 | v_792;
assign x_5545 = ~v_885 | v_789 | v_790;
assign x_5546 = ~v_885 | v_787 | v_788;
assign x_5547 = ~v_885 | v_785 | v_786;
assign x_5548 = ~v_885 | v_783 | v_784;
assign x_5549 = ~v_885 | v_781 | v_782;
assign x_5550 = ~v_885 | v_779 | v_780;
assign x_5551 = ~v_885 | v_777 | v_778;
assign x_5552 = ~v_885 | v_775 | v_776;
assign x_5553 = ~v_885 | v_773 | v_774;
assign x_5554 = ~v_885 | v_771 | v_772;
assign x_5555 = ~v_885 | v_769 | v_770;
assign x_5556 = ~v_885 | v_767 | v_768;
assign x_5557 = ~v_885 | v_765 | v_766;
assign x_5558 = ~v_885 | v_763 | v_764;
assign x_5559 = ~v_885 | v_761 | v_762;
assign x_5560 = ~v_885 | v_759 | v_760;
assign x_5561 = ~v_885 | v_757 | v_758;
assign x_5562 = ~v_885 | v_755 | v_756;
assign x_5563 = ~v_885 | v_753 | v_754;
assign x_5564 = ~v_885 | v_751 | v_752;
assign x_5565 = ~v_885 | v_749 | v_750;
assign x_5566 = ~v_885 | v_747 | v_748;
assign x_5567 = ~v_885 | v_745 | v_746;
assign x_5568 = ~v_885 | v_743 | v_744;
assign x_5569 = ~v_885 | v_741 | v_742;
assign x_5570 = ~v_885 | v_739 | v_740;
assign x_5571 = ~v_885 | v_737 | v_738;
assign x_5572 = ~v_885 | v_735 | v_736;
assign x_5573 = ~v_885 | v_733 | v_734;
assign x_5574 = ~v_885 | v_731 | v_732;
assign x_5575 = ~v_885 | v_729 | v_730;
assign x_5576 = ~v_885 | v_727 | v_728;
assign x_5577 = ~v_885 | v_725 | v_726;
assign x_5578 = ~v_885 | v_723 | v_724;
assign x_5579 = ~v_885 | v_721 | v_722;
assign x_5580 = ~v_885 | v_719 | v_720;
assign x_5581 = ~v_885 | v_717 | v_718;
assign x_5582 = ~v_885 | v_715 | v_716;
assign x_5583 = ~v_885 | v_713 | v_714;
assign x_5584 = ~v_885 | v_711 | v_712;
assign x_5585 = ~v_885 | v_709 | v_710;
assign x_5586 = ~v_885 | v_707 | v_708;
assign x_5587 = ~v_885 | v_705 | v_706;
assign x_5588 = ~v_885 | v_659;
assign x_5589 = ~v_884 | v_146;
assign x_5590 = ~v_884 | v_23;
assign x_5591 = ~v_884 | ~v_24;
assign x_5592 = ~v_883 | v_147;
assign x_5593 = ~v_883 | v_23;
assign x_5594 = ~v_883 | ~v_25;
assign x_5595 = ~v_882 | v_148;
assign x_5596 = ~v_882 | v_23;
assign x_5597 = ~v_882 | ~v_26;
assign x_5598 = ~v_881 | v_149;
assign x_5599 = ~v_881 | v_23;
assign x_5600 = ~v_881 | ~v_27;
assign x_5601 = ~v_880 | v_150;
assign x_5602 = ~v_880 | v_23;
assign x_5603 = ~v_880 | ~v_28;
assign x_5604 = ~v_879 | v_151;
assign x_5605 = ~v_879 | v_23;
assign x_5606 = ~v_879 | ~v_29;
assign x_5607 = ~v_878 | v_152;
assign x_5608 = ~v_878 | v_23;
assign x_5609 = ~v_878 | ~v_30;
assign x_5610 = ~v_877 | v_153;
assign x_5611 = ~v_877 | v_23;
assign x_5612 = ~v_877 | ~v_31;
assign x_5613 = ~v_876 | v_154;
assign x_5614 = ~v_876 | v_23;
assign x_5615 = ~v_876 | ~v_32;
assign x_5616 = ~v_875 | v_146;
assign x_5617 = ~v_875 | v_23;
assign x_5618 = ~v_875 | ~v_24;
assign x_5619 = ~v_874 | v_155;
assign x_5620 = ~v_874 | v_24;
assign x_5621 = ~v_874 | ~v_25;
assign x_5622 = ~v_873 | v_156;
assign x_5623 = ~v_873 | v_24;
assign x_5624 = ~v_873 | ~v_26;
assign x_5625 = ~v_872 | v_157;
assign x_5626 = ~v_872 | v_24;
assign x_5627 = ~v_872 | ~v_27;
assign x_5628 = ~v_871 | v_158;
assign x_5629 = ~v_871 | v_24;
assign x_5630 = ~v_871 | ~v_28;
assign x_5631 = ~v_870 | v_159;
assign x_5632 = ~v_870 | v_24;
assign x_5633 = ~v_870 | ~v_29;
assign x_5634 = ~v_869 | v_160;
assign x_5635 = ~v_869 | v_24;
assign x_5636 = ~v_869 | ~v_30;
assign x_5637 = ~v_868 | v_161;
assign x_5638 = ~v_868 | v_24;
assign x_5639 = ~v_868 | ~v_31;
assign x_5640 = ~v_867 | v_162;
assign x_5641 = ~v_867 | v_24;
assign x_5642 = ~v_867 | ~v_32;
assign x_5643 = ~v_866 | v_147;
assign x_5644 = ~v_866 | v_23;
assign x_5645 = ~v_866 | ~v_25;
assign x_5646 = ~v_865 | v_155;
assign x_5647 = ~v_865 | v_24;
assign x_5648 = ~v_865 | ~v_25;
assign x_5649 = ~v_864 | v_163;
assign x_5650 = ~v_864 | v_25;
assign x_5651 = ~v_864 | ~v_26;
assign x_5652 = ~v_863 | v_164;
assign x_5653 = ~v_863 | v_25;
assign x_5654 = ~v_863 | ~v_27;
assign x_5655 = ~v_862 | v_165;
assign x_5656 = ~v_862 | v_25;
assign x_5657 = ~v_862 | ~v_28;
assign x_5658 = ~v_861 | v_166;
assign x_5659 = ~v_861 | v_25;
assign x_5660 = ~v_861 | ~v_29;
assign x_5661 = ~v_860 | v_167;
assign x_5662 = ~v_860 | v_25;
assign x_5663 = ~v_860 | ~v_30;
assign x_5664 = ~v_859 | v_168;
assign x_5665 = ~v_859 | v_25;
assign x_5666 = ~v_859 | ~v_31;
assign x_5667 = ~v_858 | v_169;
assign x_5668 = ~v_858 | v_25;
assign x_5669 = ~v_858 | ~v_32;
assign x_5670 = ~v_857 | v_148;
assign x_5671 = ~v_857 | v_23;
assign x_5672 = ~v_857 | ~v_26;
assign x_5673 = ~v_856 | v_156;
assign x_5674 = ~v_856 | v_24;
assign x_5675 = ~v_856 | ~v_26;
assign x_5676 = ~v_855 | v_163;
assign x_5677 = ~v_855 | v_25;
assign x_5678 = ~v_855 | ~v_26;
assign x_5679 = ~v_854 | v_170;
assign x_5680 = ~v_854 | v_26;
assign x_5681 = ~v_854 | ~v_27;
assign x_5682 = ~v_853 | v_171;
assign x_5683 = ~v_853 | v_26;
assign x_5684 = ~v_853 | ~v_28;
assign x_5685 = ~v_852 | v_172;
assign x_5686 = ~v_852 | v_26;
assign x_5687 = ~v_852 | ~v_29;
assign x_5688 = ~v_851 | v_173;
assign x_5689 = ~v_851 | v_26;
assign x_5690 = ~v_851 | ~v_30;
assign x_5691 = ~v_850 | v_174;
assign x_5692 = ~v_850 | v_26;
assign x_5693 = ~v_850 | ~v_31;
assign x_5694 = ~v_849 | v_175;
assign x_5695 = ~v_849 | v_26;
assign x_5696 = ~v_849 | ~v_32;
assign x_5697 = ~v_848 | v_149;
assign x_5698 = ~v_848 | v_23;
assign x_5699 = ~v_848 | ~v_27;
assign x_5700 = ~v_847 | v_157;
assign x_5701 = ~v_847 | v_24;
assign x_5702 = ~v_847 | ~v_27;
assign x_5703 = ~v_846 | v_164;
assign x_5704 = ~v_846 | v_25;
assign x_5705 = ~v_846 | ~v_27;
assign x_5706 = ~v_845 | v_170;
assign x_5707 = ~v_845 | v_26;
assign x_5708 = ~v_845 | ~v_27;
assign x_5709 = ~v_844 | v_176;
assign x_5710 = ~v_844 | v_27;
assign x_5711 = ~v_844 | ~v_28;
assign x_5712 = ~v_843 | v_177;
assign x_5713 = ~v_843 | v_27;
assign x_5714 = ~v_843 | ~v_29;
assign x_5715 = ~v_842 | v_178;
assign x_5716 = ~v_842 | v_27;
assign x_5717 = ~v_842 | ~v_30;
assign x_5718 = ~v_841 | v_179;
assign x_5719 = ~v_841 | v_27;
assign x_5720 = ~v_841 | ~v_31;
assign x_5721 = ~v_840 | v_180;
assign x_5722 = ~v_840 | v_27;
assign x_5723 = ~v_840 | ~v_32;
assign x_5724 = ~v_839 | v_150;
assign x_5725 = ~v_839 | v_23;
assign x_5726 = ~v_839 | ~v_28;
assign x_5727 = ~v_838 | v_158;
assign x_5728 = ~v_838 | v_24;
assign x_5729 = ~v_838 | ~v_28;
assign x_5730 = ~v_837 | v_165;
assign x_5731 = ~v_837 | v_25;
assign x_5732 = ~v_837 | ~v_28;
assign x_5733 = ~v_836 | v_171;
assign x_5734 = ~v_836 | v_26;
assign x_5735 = ~v_836 | ~v_28;
assign x_5736 = ~v_835 | v_176;
assign x_5737 = ~v_835 | v_27;
assign x_5738 = ~v_835 | ~v_28;
assign x_5739 = ~v_834 | v_181;
assign x_5740 = ~v_834 | v_28;
assign x_5741 = ~v_834 | ~v_29;
assign x_5742 = ~v_833 | v_182;
assign x_5743 = ~v_833 | v_28;
assign x_5744 = ~v_833 | ~v_30;
assign x_5745 = ~v_832 | v_183;
assign x_5746 = ~v_832 | v_28;
assign x_5747 = ~v_832 | ~v_31;
assign x_5748 = ~v_831 | v_184;
assign x_5749 = ~v_831 | v_28;
assign x_5750 = ~v_831 | ~v_32;
assign x_5751 = ~v_830 | v_151;
assign x_5752 = ~v_830 | v_23;
assign x_5753 = ~v_830 | ~v_29;
assign x_5754 = ~v_829 | v_159;
assign x_5755 = ~v_829 | v_24;
assign x_5756 = ~v_829 | ~v_29;
assign x_5757 = ~v_828 | v_166;
assign x_5758 = ~v_828 | v_25;
assign x_5759 = ~v_828 | ~v_29;
assign x_5760 = ~v_827 | v_172;
assign x_5761 = ~v_827 | v_26;
assign x_5762 = ~v_827 | ~v_29;
assign x_5763 = ~v_826 | v_177;
assign x_5764 = ~v_826 | v_27;
assign x_5765 = ~v_826 | ~v_29;
assign x_5766 = ~v_825 | v_181;
assign x_5767 = ~v_825 | v_28;
assign x_5768 = ~v_825 | ~v_29;
assign x_5769 = ~v_824 | v_185;
assign x_5770 = ~v_824 | v_29;
assign x_5771 = ~v_824 | ~v_30;
assign x_5772 = ~v_823 | v_186;
assign x_5773 = ~v_823 | v_29;
assign x_5774 = ~v_823 | ~v_31;
assign x_5775 = ~v_822 | v_187;
assign x_5776 = ~v_822 | v_29;
assign x_5777 = ~v_822 | ~v_32;
assign x_5778 = ~v_821 | v_152;
assign x_5779 = ~v_821 | v_23;
assign x_5780 = ~v_821 | ~v_30;
assign x_5781 = ~v_820 | v_160;
assign x_5782 = ~v_820 | v_24;
assign x_5783 = ~v_820 | ~v_30;
assign x_5784 = ~v_819 | v_167;
assign x_5785 = ~v_819 | v_25;
assign x_5786 = ~v_819 | ~v_30;
assign x_5787 = ~v_818 | v_173;
assign x_5788 = ~v_818 | v_26;
assign x_5789 = ~v_818 | ~v_30;
assign x_5790 = ~v_817 | v_178;
assign x_5791 = ~v_817 | v_27;
assign x_5792 = ~v_817 | ~v_30;
assign x_5793 = ~v_816 | v_182;
assign x_5794 = ~v_816 | v_28;
assign x_5795 = ~v_816 | ~v_30;
assign x_5796 = ~v_815 | v_185;
assign x_5797 = ~v_815 | v_29;
assign x_5798 = ~v_815 | ~v_30;
assign x_5799 = ~v_814 | v_188;
assign x_5800 = ~v_814 | v_30;
assign x_5801 = ~v_814 | ~v_31;
assign x_5802 = ~v_813 | v_189;
assign x_5803 = ~v_813 | v_30;
assign x_5804 = ~v_813 | ~v_32;
assign x_5805 = ~v_812 | v_153;
assign x_5806 = ~v_812 | v_23;
assign x_5807 = ~v_812 | ~v_31;
assign x_5808 = ~v_811 | v_161;
assign x_5809 = ~v_811 | v_24;
assign x_5810 = ~v_811 | ~v_31;
assign x_5811 = ~v_810 | v_168;
assign x_5812 = ~v_810 | v_25;
assign x_5813 = ~v_810 | ~v_31;
assign x_5814 = ~v_809 | v_174;
assign x_5815 = ~v_809 | v_26;
assign x_5816 = ~v_809 | ~v_31;
assign x_5817 = ~v_808 | v_179;
assign x_5818 = ~v_808 | v_27;
assign x_5819 = ~v_808 | ~v_31;
assign x_5820 = ~v_807 | v_183;
assign x_5821 = ~v_807 | v_28;
assign x_5822 = ~v_807 | ~v_31;
assign x_5823 = ~v_806 | v_186;
assign x_5824 = ~v_806 | v_29;
assign x_5825 = ~v_806 | ~v_31;
assign x_5826 = ~v_805 | v_188;
assign x_5827 = ~v_805 | v_30;
assign x_5828 = ~v_805 | ~v_31;
assign x_5829 = ~v_804 | v_190;
assign x_5830 = ~v_804 | v_31;
assign x_5831 = ~v_804 | ~v_32;
assign x_5832 = ~v_803 | v_154;
assign x_5833 = ~v_803 | v_23;
assign x_5834 = ~v_803 | ~v_32;
assign x_5835 = ~v_802 | v_162;
assign x_5836 = ~v_802 | v_24;
assign x_5837 = ~v_802 | ~v_32;
assign x_5838 = ~v_801 | v_169;
assign x_5839 = ~v_801 | v_25;
assign x_5840 = ~v_801 | ~v_32;
assign x_5841 = ~v_800 | v_175;
assign x_5842 = ~v_800 | v_26;
assign x_5843 = ~v_800 | ~v_32;
assign x_5844 = ~v_799 | v_180;
assign x_5845 = ~v_799 | v_27;
assign x_5846 = ~v_799 | ~v_32;
assign x_5847 = ~v_798 | v_184;
assign x_5848 = ~v_798 | v_28;
assign x_5849 = ~v_798 | ~v_32;
assign x_5850 = ~v_797 | v_187;
assign x_5851 = ~v_797 | v_29;
assign x_5852 = ~v_797 | ~v_32;
assign x_5853 = ~v_796 | v_189;
assign x_5854 = ~v_796 | v_30;
assign x_5855 = ~v_796 | ~v_32;
assign x_5856 = ~v_795 | v_190;
assign x_5857 = ~v_795 | v_31;
assign x_5858 = ~v_795 | ~v_32;
assign x_5859 = ~v_793 | ~v_146 | ~v_23 | v_24;
assign x_5860 = ~v_794 | ~v_34;
assign x_5861 = ~v_794 | v_35;
assign x_5862 = ~v_791 | ~v_147 | ~v_23 | v_25;
assign x_5863 = ~v_792 | ~v_34;
assign x_5864 = ~v_792 | v_36;
assign x_5865 = ~v_789 | ~v_148 | ~v_23 | v_26;
assign x_5866 = ~v_790 | ~v_34;
assign x_5867 = ~v_790 | v_37;
assign x_5868 = ~v_787 | ~v_149 | ~v_23 | v_27;
assign x_5869 = ~v_788 | ~v_34;
assign x_5870 = ~v_788 | v_38;
assign x_5871 = ~v_785 | ~v_150 | ~v_23 | v_28;
assign x_5872 = ~v_786 | ~v_34;
assign x_5873 = ~v_786 | v_39;
assign x_5874 = ~v_783 | ~v_151 | ~v_23 | v_29;
assign x_5875 = ~v_784 | ~v_34;
assign x_5876 = ~v_784 | v_40;
assign x_5877 = ~v_781 | ~v_152 | ~v_23 | v_30;
assign x_5878 = ~v_782 | ~v_34;
assign x_5879 = ~v_782 | v_41;
assign x_5880 = ~v_779 | ~v_153 | ~v_23 | v_31;
assign x_5881 = ~v_780 | ~v_34;
assign x_5882 = ~v_780 | v_42;
assign x_5883 = ~v_777 | ~v_154 | ~v_23 | v_32;
assign x_5884 = ~v_778 | ~v_34;
assign x_5885 = ~v_778 | v_43;
assign x_5886 = ~v_775 | ~v_155 | ~v_24 | v_25;
assign x_5887 = ~v_776 | ~v_35;
assign x_5888 = ~v_776 | v_36;
assign x_5889 = ~v_773 | ~v_156 | ~v_24 | v_26;
assign x_5890 = ~v_774 | ~v_35;
assign x_5891 = ~v_774 | v_37;
assign x_5892 = ~v_771 | ~v_157 | ~v_24 | v_27;
assign x_5893 = ~v_772 | ~v_35;
assign x_5894 = ~v_772 | v_38;
assign x_5895 = ~v_769 | ~v_158 | ~v_24 | v_28;
assign x_5896 = ~v_770 | ~v_35;
assign x_5897 = ~v_770 | v_39;
assign x_5898 = ~v_767 | ~v_159 | ~v_24 | v_29;
assign x_5899 = ~v_768 | ~v_35;
assign x_5900 = ~v_768 | v_40;
assign x_5901 = ~v_765 | ~v_160 | ~v_24 | v_30;
assign x_5902 = ~v_766 | ~v_35;
assign x_5903 = ~v_766 | v_41;
assign x_5904 = ~v_763 | ~v_161 | ~v_24 | v_31;
assign x_5905 = ~v_764 | ~v_35;
assign x_5906 = ~v_764 | v_42;
assign x_5907 = ~v_761 | ~v_162 | ~v_24 | v_32;
assign x_5908 = ~v_762 | ~v_35;
assign x_5909 = ~v_762 | v_43;
assign x_5910 = ~v_759 | ~v_163 | ~v_25 | v_26;
assign x_5911 = ~v_760 | ~v_36;
assign x_5912 = ~v_760 | v_37;
assign x_5913 = ~v_757 | ~v_164 | ~v_25 | v_27;
assign x_5914 = ~v_758 | ~v_36;
assign x_5915 = ~v_758 | v_38;
assign x_5916 = ~v_755 | ~v_165 | ~v_25 | v_28;
assign x_5917 = ~v_756 | ~v_36;
assign x_5918 = ~v_756 | v_39;
assign x_5919 = ~v_753 | ~v_166 | ~v_25 | v_29;
assign x_5920 = ~v_754 | ~v_36;
assign x_5921 = ~v_754 | v_40;
assign x_5922 = ~v_751 | ~v_167 | ~v_25 | v_30;
assign x_5923 = ~v_752 | ~v_36;
assign x_5924 = ~v_752 | v_41;
assign x_5925 = ~v_749 | ~v_168 | ~v_25 | v_31;
assign x_5926 = ~v_750 | ~v_36;
assign x_5927 = ~v_750 | v_42;
assign x_5928 = ~v_747 | ~v_169 | ~v_25 | v_32;
assign x_5929 = ~v_748 | ~v_36;
assign x_5930 = ~v_748 | v_43;
assign x_5931 = ~v_745 | ~v_170 | ~v_26 | v_27;
assign x_5932 = ~v_746 | ~v_37;
assign x_5933 = ~v_746 | v_38;
assign x_5934 = ~v_743 | ~v_171 | ~v_26 | v_28;
assign x_5935 = ~v_744 | ~v_37;
assign x_5936 = ~v_744 | v_39;
assign x_5937 = ~v_741 | ~v_172 | ~v_26 | v_29;
assign x_5938 = ~v_742 | ~v_37;
assign x_5939 = ~v_742 | v_40;
assign x_5940 = ~v_739 | ~v_173 | ~v_26 | v_30;
assign x_5941 = ~v_740 | ~v_37;
assign x_5942 = ~v_740 | v_41;
assign x_5943 = ~v_737 | ~v_174 | ~v_26 | v_31;
assign x_5944 = ~v_738 | ~v_37;
assign x_5945 = ~v_738 | v_42;
assign x_5946 = ~v_735 | ~v_175 | ~v_26 | v_32;
assign x_5947 = ~v_736 | ~v_37;
assign x_5948 = ~v_736 | v_43;
assign x_5949 = ~v_733 | ~v_176 | ~v_27 | v_28;
assign x_5950 = ~v_734 | ~v_38;
assign x_5951 = ~v_734 | v_39;
assign x_5952 = ~v_731 | ~v_177 | ~v_27 | v_29;
assign x_5953 = ~v_732 | ~v_38;
assign x_5954 = ~v_732 | v_40;
assign x_5955 = ~v_729 | ~v_178 | ~v_27 | v_30;
assign x_5956 = ~v_730 | ~v_38;
assign x_5957 = ~v_730 | v_41;
assign x_5958 = ~v_727 | ~v_179 | ~v_27 | v_31;
assign x_5959 = ~v_728 | ~v_38;
assign x_5960 = ~v_728 | v_42;
assign x_5961 = ~v_725 | ~v_180 | ~v_27 | v_32;
assign x_5962 = ~v_726 | ~v_38;
assign x_5963 = ~v_726 | v_43;
assign x_5964 = ~v_723 | ~v_181 | ~v_28 | v_29;
assign x_5965 = ~v_724 | ~v_39;
assign x_5966 = ~v_724 | v_40;
assign x_5967 = ~v_721 | ~v_182 | ~v_28 | v_30;
assign x_5968 = ~v_722 | ~v_39;
assign x_5969 = ~v_722 | v_41;
assign x_5970 = ~v_719 | ~v_183 | ~v_28 | v_31;
assign x_5971 = ~v_720 | ~v_39;
assign x_5972 = ~v_720 | v_42;
assign x_5973 = ~v_717 | ~v_184 | ~v_28 | v_32;
assign x_5974 = ~v_718 | ~v_39;
assign x_5975 = ~v_718 | v_43;
assign x_5976 = ~v_715 | ~v_185 | ~v_29 | v_30;
assign x_5977 = ~v_716 | ~v_40;
assign x_5978 = ~v_716 | v_41;
assign x_5979 = ~v_713 | ~v_186 | ~v_29 | v_31;
assign x_5980 = ~v_714 | ~v_40;
assign x_5981 = ~v_714 | v_42;
assign x_5982 = ~v_711 | ~v_187 | ~v_29 | v_32;
assign x_5983 = ~v_712 | ~v_40;
assign x_5984 = ~v_712 | v_43;
assign x_5985 = ~v_709 | ~v_188 | ~v_30 | v_31;
assign x_5986 = ~v_710 | ~v_41;
assign x_5987 = ~v_710 | v_42;
assign x_5988 = ~v_707 | ~v_189 | ~v_30 | v_32;
assign x_5989 = ~v_708 | ~v_41;
assign x_5990 = ~v_708 | v_43;
assign x_5991 = ~v_705 | ~v_190 | ~v_31 | v_32;
assign x_5992 = ~v_706 | ~v_42;
assign x_5993 = ~v_706 | v_43;
assign x_5994 = ~v_659 | v_34 | ~v_45;
assign x_5995 = ~v_659 | ~v_34 | v_45 | v_4020 | v_4019 | v_4018 | v_4017 | v_4016 | v_4015 | v_4014 | v_4013 | v_4012;
assign x_5996 = ~v_659 | ~v_4020 | v_658;
assign x_5997 = ~v_659 | ~v_191 | ~v_34 | v_35 | v_4020;
assign x_5998 = ~v_659 | ~v_4019 | v_657;
assign x_5999 = ~v_659 | ~v_192 | ~v_34 | v_36 | v_4019;
assign x_6000 = ~v_659 | ~v_4018 | v_656;
assign x_6001 = ~v_659 | ~v_193 | ~v_34 | v_37 | v_4018;
assign x_6002 = ~v_659 | ~v_4017 | v_655;
assign x_6003 = ~v_659 | ~v_194 | ~v_34 | v_38 | v_4017;
assign x_6004 = ~v_659 | ~v_4016 | v_654;
assign x_6005 = ~v_659 | ~v_195 | ~v_34 | v_39 | v_4016;
assign x_6006 = ~v_659 | ~v_4015 | v_653;
assign x_6007 = ~v_659 | ~v_196 | ~v_34 | v_40 | v_4015;
assign x_6008 = ~v_659 | ~v_4014 | v_652;
assign x_6009 = ~v_659 | ~v_197 | ~v_34 | v_41 | v_4014;
assign x_6010 = ~v_659 | ~v_4013 | v_651;
assign x_6011 = ~v_659 | ~v_198 | ~v_34 | v_42 | v_4013;
assign x_6012 = ~v_659 | ~v_4012 | v_650;
assign x_6013 = ~v_659 | ~v_199 | ~v_34 | v_43 | v_4012;
assign x_6014 = ~v_659 | v_35 | ~v_46 | v_4021;
assign x_6015 = ~v_659 | ~v_35 | v_46 | v_4029 | v_4028 | v_4027 | v_4026 | v_4025 | v_4024 | v_4023 | v_4022;
assign x_6016 = ~v_659 | ~v_4021 | v_649;
assign x_6017 = ~v_659 | ~v_191 | ~v_34 | v_35 | v_4021;
assign x_6018 = ~v_659 | ~v_4029 | v_648;
assign x_6019 = ~v_659 | ~v_200 | ~v_35 | v_36 | v_4029;
assign x_6020 = ~v_659 | ~v_4028 | v_647;
assign x_6021 = ~v_659 | ~v_201 | ~v_35 | v_37 | v_4028;
assign x_6022 = ~v_659 | ~v_4027 | v_646;
assign x_6023 = ~v_659 | ~v_202 | ~v_35 | v_38 | v_4027;
assign x_6024 = ~v_659 | ~v_4026 | v_645;
assign x_6025 = ~v_659 | ~v_203 | ~v_35 | v_39 | v_4026;
assign x_6026 = ~v_659 | ~v_4025 | v_644;
assign x_6027 = ~v_659 | ~v_204 | ~v_35 | v_40 | v_4025;
assign x_6028 = ~v_659 | ~v_4024 | v_643;
assign x_6029 = ~v_659 | ~v_205 | ~v_35 | v_41 | v_4024;
assign x_6030 = ~v_659 | ~v_4023 | v_642;
assign x_6031 = ~v_659 | ~v_206 | ~v_35 | v_42 | v_4023;
assign x_6032 = ~v_659 | ~v_4022 | v_641;
assign x_6033 = ~v_659 | ~v_207 | ~v_35 | v_43 | v_4022;
assign x_6034 = ~v_659 | v_36 | ~v_47 | v_4031 | v_4030;
assign x_6035 = ~v_659 | ~v_36 | v_47 | v_4038 | v_4037 | v_4036 | v_4035 | v_4034 | v_4033 | v_4032;
assign x_6036 = ~v_659 | ~v_4031 | v_640;
assign x_6037 = ~v_659 | ~v_192 | ~v_34 | v_36 | v_4031;
assign x_6038 = ~v_659 | ~v_4030 | v_639;
assign x_6039 = ~v_659 | ~v_200 | ~v_35 | v_36 | v_4030;
assign x_6040 = ~v_659 | ~v_4038 | v_638;
assign x_6041 = ~v_659 | ~v_208 | ~v_36 | v_37 | v_4038;
assign x_6042 = ~v_659 | ~v_4037 | v_637;
assign x_6043 = ~v_659 | ~v_209 | ~v_36 | v_38 | v_4037;
assign x_6044 = ~v_659 | ~v_4036 | v_636;
assign x_6045 = ~v_659 | ~v_210 | ~v_36 | v_39 | v_4036;
assign x_6046 = ~v_659 | ~v_4035 | v_635;
assign x_6047 = ~v_659 | ~v_211 | ~v_36 | v_40 | v_4035;
assign x_6048 = ~v_659 | ~v_4034 | v_634;
assign x_6049 = ~v_659 | ~v_212 | ~v_36 | v_41 | v_4034;
assign x_6050 = ~v_659 | ~v_4033 | v_633;
assign x_6051 = ~v_659 | ~v_213 | ~v_36 | v_42 | v_4033;
assign x_6052 = ~v_659 | ~v_4032 | v_632;
assign x_6053 = ~v_659 | ~v_214 | ~v_36 | v_43 | v_4032;
assign x_6054 = ~v_659 | v_37 | ~v_48 | v_4041 | v_4040 | v_4039;
assign x_6055 = ~v_659 | ~v_37 | v_48 | v_4047 | v_4046 | v_4045 | v_4044 | v_4043 | v_4042;
assign x_6056 = ~v_659 | ~v_4041 | v_631;
assign x_6057 = ~v_659 | ~v_193 | ~v_34 | v_37 | v_4041;
assign x_6058 = ~v_659 | ~v_4040 | v_630;
assign x_6059 = ~v_659 | ~v_201 | ~v_35 | v_37 | v_4040;
assign x_6060 = ~v_659 | ~v_4039 | v_629;
assign x_6061 = ~v_659 | ~v_208 | ~v_36 | v_37 | v_4039;
assign x_6062 = ~v_659 | ~v_4047 | v_628;
assign x_6063 = ~v_659 | ~v_215 | ~v_37 | v_38 | v_4047;
assign x_6064 = ~v_659 | ~v_4046 | v_627;
assign x_6065 = ~v_659 | ~v_216 | ~v_37 | v_39 | v_4046;
assign x_6066 = ~v_659 | ~v_4045 | v_626;
assign x_6067 = ~v_659 | ~v_217 | ~v_37 | v_40 | v_4045;
assign x_6068 = ~v_659 | ~v_4044 | v_625;
assign x_6069 = ~v_659 | ~v_218 | ~v_37 | v_41 | v_4044;
assign x_6070 = ~v_659 | ~v_4043 | v_624;
assign x_6071 = ~v_659 | ~v_219 | ~v_37 | v_42 | v_4043;
assign x_6072 = ~v_659 | ~v_4042 | v_623;
assign x_6073 = ~v_659 | ~v_220 | ~v_37 | v_43 | v_4042;
assign x_6074 = ~v_659 | v_38 | ~v_49 | v_4051 | v_4050 | v_4049 | v_4048;
assign x_6075 = ~v_659 | ~v_38 | v_49 | v_4056 | v_4055 | v_4054 | v_4053 | v_4052;
assign x_6076 = ~v_659 | ~v_4051 | v_622;
assign x_6077 = ~v_659 | ~v_194 | ~v_34 | v_38 | v_4051;
assign x_6078 = ~v_659 | ~v_4050 | v_621;
assign x_6079 = ~v_659 | ~v_202 | ~v_35 | v_38 | v_4050;
assign x_6080 = ~v_659 | ~v_4049 | v_620;
assign x_6081 = ~v_659 | ~v_209 | ~v_36 | v_38 | v_4049;
assign x_6082 = ~v_659 | ~v_4048 | v_619;
assign x_6083 = ~v_659 | ~v_215 | ~v_37 | v_38 | v_4048;
assign x_6084 = ~v_659 | ~v_4056 | v_618;
assign x_6085 = ~v_659 | ~v_221 | ~v_38 | v_39 | v_4056;
assign x_6086 = ~v_659 | ~v_4055 | v_617;
assign x_6087 = ~v_659 | ~v_222 | ~v_38 | v_40 | v_4055;
assign x_6088 = ~v_659 | ~v_4054 | v_616;
assign x_6089 = ~v_659 | ~v_223 | ~v_38 | v_41 | v_4054;
assign x_6090 = ~v_659 | ~v_4053 | v_615;
assign x_6091 = ~v_659 | ~v_224 | ~v_38 | v_42 | v_4053;
assign x_6092 = ~v_659 | ~v_4052 | v_614;
assign x_6093 = ~v_659 | ~v_225 | ~v_38 | v_43 | v_4052;
assign x_6094 = ~v_659 | v_39 | ~v_50 | v_4061 | v_4060 | v_4059 | v_4058 | v_4057;
assign x_6095 = ~v_659 | ~v_39 | v_50 | v_4065 | v_4064 | v_4063 | v_4062;
assign x_6096 = ~v_659 | ~v_4061 | v_613;
assign x_6097 = ~v_659 | ~v_195 | ~v_34 | v_39 | v_4061;
assign x_6098 = ~v_659 | ~v_4060 | v_612;
assign x_6099 = ~v_659 | ~v_203 | ~v_35 | v_39 | v_4060;
assign x_6100 = ~v_659 | ~v_4059 | v_611;
assign x_6101 = ~v_659 | ~v_210 | ~v_36 | v_39 | v_4059;
assign x_6102 = ~v_659 | ~v_4058 | v_610;
assign x_6103 = ~v_659 | ~v_216 | ~v_37 | v_39 | v_4058;
assign x_6104 = ~v_659 | ~v_4057 | v_609;
assign x_6105 = ~v_659 | ~v_221 | ~v_38 | v_39 | v_4057;
assign x_6106 = ~v_659 | ~v_4065 | v_608;
assign x_6107 = ~v_659 | ~v_226 | ~v_39 | v_40 | v_4065;
assign x_6108 = ~v_659 | ~v_4064 | v_607;
assign x_6109 = ~v_659 | ~v_227 | ~v_39 | v_41 | v_4064;
assign x_6110 = ~v_659 | ~v_4063 | v_606;
assign x_6111 = ~v_659 | ~v_228 | ~v_39 | v_42 | v_4063;
assign x_6112 = ~v_659 | ~v_4062 | v_605;
assign x_6113 = ~v_659 | ~v_229 | ~v_39 | v_43 | v_4062;
assign x_6114 = ~v_659 | v_40 | ~v_51 | v_4071 | v_4070 | v_4069 | v_4068 | v_4067 | v_4066;
assign x_6115 = ~v_659 | ~v_40 | v_51 | v_4074 | v_4073 | v_4072;
assign x_6116 = ~v_659 | ~v_4071 | v_604;
assign x_6117 = ~v_659 | ~v_196 | ~v_34 | v_40 | v_4071;
assign x_6118 = ~v_659 | ~v_4070 | v_603;
assign x_6119 = ~v_659 | ~v_204 | ~v_35 | v_40 | v_4070;
assign x_6120 = ~v_659 | ~v_4069 | v_602;
assign x_6121 = ~v_659 | ~v_211 | ~v_36 | v_40 | v_4069;
assign x_6122 = ~v_659 | ~v_4068 | v_601;
assign x_6123 = ~v_659 | ~v_217 | ~v_37 | v_40 | v_4068;
assign x_6124 = ~v_659 | ~v_4067 | v_600;
assign x_6125 = ~v_659 | ~v_222 | ~v_38 | v_40 | v_4067;
assign x_6126 = ~v_659 | ~v_4066 | v_599;
assign x_6127 = ~v_659 | ~v_226 | ~v_39 | v_40 | v_4066;
assign x_6128 = ~v_659 | ~v_4074 | v_598;
assign x_6129 = ~v_659 | ~v_230 | ~v_40 | v_41 | v_4074;
assign x_6130 = ~v_659 | ~v_4073 | v_597;
assign x_6131 = ~v_659 | ~v_231 | ~v_40 | v_42 | v_4073;
assign x_6132 = ~v_659 | ~v_4072 | v_596;
assign x_6133 = ~v_659 | ~v_232 | ~v_40 | v_43 | v_4072;
assign x_6134 = ~v_659 | v_41 | ~v_52 | v_4081 | v_4080 | v_4079 | v_4078 | v_4077 | v_4076 | v_4075;
assign x_6135 = ~v_659 | ~v_41 | v_52 | v_4083 | v_4082;
assign x_6136 = ~v_659 | ~v_4081 | v_595;
assign x_6137 = ~v_659 | ~v_197 | ~v_34 | v_41 | v_4081;
assign x_6138 = ~v_659 | ~v_4080 | v_594;
assign x_6139 = ~v_659 | ~v_205 | ~v_35 | v_41 | v_4080;
assign x_6140 = ~v_659 | ~v_4079 | v_593;
assign x_6141 = ~v_659 | ~v_212 | ~v_36 | v_41 | v_4079;
assign x_6142 = ~v_659 | ~v_4078 | v_592;
assign x_6143 = ~v_659 | ~v_218 | ~v_37 | v_41 | v_4078;
assign x_6144 = ~v_659 | ~v_4077 | v_591;
assign x_6145 = ~v_659 | ~v_223 | ~v_38 | v_41 | v_4077;
assign x_6146 = ~v_659 | ~v_4076 | v_590;
assign x_6147 = ~v_659 | ~v_227 | ~v_39 | v_41 | v_4076;
assign x_6148 = ~v_659 | ~v_4075 | v_589;
assign x_6149 = ~v_659 | ~v_230 | ~v_40 | v_41 | v_4075;
assign x_6150 = ~v_659 | ~v_4083 | v_588;
assign x_6151 = ~v_659 | ~v_233 | ~v_41 | v_42 | v_4083;
assign x_6152 = ~v_659 | ~v_4082 | v_587;
assign x_6153 = ~v_659 | ~v_234 | ~v_41 | v_43 | v_4082;
assign x_6154 = ~v_659 | v_42 | ~v_53 | v_4091 | v_4090 | v_4089 | v_4088 | v_4087 | v_4086 | v_4085 | v_4084;
assign x_6155 = ~v_659 | ~v_42 | v_53 | v_4092;
assign x_6156 = ~v_659 | ~v_4091 | v_586;
assign x_6157 = ~v_659 | ~v_198 | ~v_34 | v_42 | v_4091;
assign x_6158 = ~v_659 | ~v_4090 | v_585;
assign x_6159 = ~v_659 | ~v_206 | ~v_35 | v_42 | v_4090;
assign x_6160 = ~v_659 | ~v_4089 | v_584;
assign x_6161 = ~v_659 | ~v_213 | ~v_36 | v_42 | v_4089;
assign x_6162 = ~v_659 | ~v_4088 | v_583;
assign x_6163 = ~v_659 | ~v_219 | ~v_37 | v_42 | v_4088;
assign x_6164 = ~v_659 | ~v_4087 | v_582;
assign x_6165 = ~v_659 | ~v_224 | ~v_38 | v_42 | v_4087;
assign x_6166 = ~v_659 | ~v_4086 | v_581;
assign x_6167 = ~v_659 | ~v_228 | ~v_39 | v_42 | v_4086;
assign x_6168 = ~v_659 | ~v_4085 | v_580;
assign x_6169 = ~v_659 | ~v_231 | ~v_40 | v_42 | v_4085;
assign x_6170 = ~v_659 | ~v_4084 | v_579;
assign x_6171 = ~v_659 | ~v_233 | ~v_41 | v_42 | v_4084;
assign x_6172 = ~v_659 | ~v_4092 | v_578;
assign x_6173 = ~v_659 | ~v_235 | ~v_42 | v_43 | v_4092;
assign x_6174 = ~v_659 | v_43 | ~v_54 | v_4101 | v_4100 | v_4099 | v_4098 | v_4097 | v_4096 | v_4095 | v_4094 | v_4093;
assign x_6175 = ~v_659 | ~v_43 | v_54;
assign x_6176 = ~v_659 | ~v_4101 | v_577;
assign x_6177 = ~v_659 | ~v_199 | ~v_34 | v_43 | v_4101;
assign x_6178 = ~v_659 | ~v_4100 | v_576;
assign x_6179 = ~v_659 | ~v_207 | ~v_35 | v_43 | v_4100;
assign x_6180 = ~v_659 | ~v_4099 | v_575;
assign x_6181 = ~v_659 | ~v_214 | ~v_36 | v_43 | v_4099;
assign x_6182 = ~v_659 | ~v_4098 | v_574;
assign x_6183 = ~v_659 | ~v_220 | ~v_37 | v_43 | v_4098;
assign x_6184 = ~v_659 | ~v_4097 | v_573;
assign x_6185 = ~v_659 | ~v_225 | ~v_38 | v_43 | v_4097;
assign x_6186 = ~v_659 | ~v_4096 | v_572;
assign x_6187 = ~v_659 | ~v_229 | ~v_39 | v_43 | v_4096;
assign x_6188 = ~v_659 | ~v_4095 | v_571;
assign x_6189 = ~v_659 | ~v_232 | ~v_40 | v_43 | v_4095;
assign x_6190 = ~v_659 | ~v_4094 | v_570;
assign x_6191 = ~v_659 | ~v_234 | ~v_41 | v_43 | v_4094;
assign x_6192 = ~v_659 | ~v_4093 | v_569;
assign x_6193 = ~v_659 | ~v_235 | ~v_42 | v_43 | v_4093;
assign x_6194 = ~v_659 | v_44 | ~v_55;
assign x_6195 = ~v_659 | ~v_44 | v_55;
assign x_6196 = ~v_659 | v_567 | v_568;
assign x_6197 = ~v_659 | v_565 | v_566;
assign x_6198 = ~v_659 | v_563 | v_564;
assign x_6199 = ~v_659 | v_561 | v_562;
assign x_6200 = ~v_659 | v_559 | v_560;
assign x_6201 = ~v_659 | v_557 | v_558;
assign x_6202 = ~v_659 | v_555 | v_556;
assign x_6203 = ~v_659 | v_553 | v_554;
assign x_6204 = ~v_659 | v_551 | v_552;
assign x_6205 = ~v_659 | v_549 | v_550;
assign x_6206 = ~v_659 | v_547 | v_548;
assign x_6207 = ~v_659 | v_545 | v_546;
assign x_6208 = ~v_659 | v_543 | v_544;
assign x_6209 = ~v_659 | v_541 | v_542;
assign x_6210 = ~v_659 | v_539 | v_540;
assign x_6211 = ~v_659 | v_537 | v_538;
assign x_6212 = ~v_659 | v_535 | v_536;
assign x_6213 = ~v_659 | v_533 | v_534;
assign x_6214 = ~v_659 | v_531 | v_532;
assign x_6215 = ~v_659 | v_529 | v_530;
assign x_6216 = ~v_659 | v_527 | v_528;
assign x_6217 = ~v_659 | v_525 | v_526;
assign x_6218 = ~v_659 | v_523 | v_524;
assign x_6219 = ~v_659 | v_521 | v_522;
assign x_6220 = ~v_659 | v_519 | v_520;
assign x_6221 = ~v_659 | v_517 | v_518;
assign x_6222 = ~v_659 | v_515 | v_516;
assign x_6223 = ~v_659 | v_513 | v_514;
assign x_6224 = ~v_659 | v_511 | v_512;
assign x_6225 = ~v_659 | v_509 | v_510;
assign x_6226 = ~v_659 | v_507 | v_508;
assign x_6227 = ~v_659 | v_505 | v_506;
assign x_6228 = ~v_659 | v_503 | v_504;
assign x_6229 = ~v_659 | v_501 | v_502;
assign x_6230 = ~v_659 | v_499 | v_500;
assign x_6231 = ~v_659 | v_497 | v_498;
assign x_6232 = ~v_659 | v_495 | v_496;
assign x_6233 = ~v_659 | v_493 | v_494;
assign x_6234 = ~v_659 | v_491 | v_492;
assign x_6235 = ~v_659 | v_489 | v_490;
assign x_6236 = ~v_659 | v_487 | v_488;
assign x_6237 = ~v_659 | v_485 | v_486;
assign x_6238 = ~v_659 | v_483 | v_484;
assign x_6239 = ~v_659 | v_481 | v_482;
assign x_6240 = ~v_659 | v_479 | v_480;
assign x_6241 = ~v_659 | v_470 | v_471 | v_472 | v_473 | v_474 | v_475 | v_476 | v_477 | v_478;
assign x_6242 = ~v_658 | v_191;
assign x_6243 = ~v_658 | v_34;
assign x_6244 = ~v_658 | ~v_35;
assign x_6245 = ~v_657 | v_192;
assign x_6246 = ~v_657 | v_34;
assign x_6247 = ~v_657 | ~v_36;
assign x_6248 = ~v_656 | v_193;
assign x_6249 = ~v_656 | v_34;
assign x_6250 = ~v_656 | ~v_37;
assign x_6251 = ~v_655 | v_194;
assign x_6252 = ~v_655 | v_34;
assign x_6253 = ~v_655 | ~v_38;
assign x_6254 = ~v_654 | v_195;
assign x_6255 = ~v_654 | v_34;
assign x_6256 = ~v_654 | ~v_39;
assign x_6257 = ~v_653 | v_196;
assign x_6258 = ~v_653 | v_34;
assign x_6259 = ~v_653 | ~v_40;
assign x_6260 = ~v_652 | v_197;
assign x_6261 = ~v_652 | v_34;
assign x_6262 = ~v_652 | ~v_41;
assign x_6263 = ~v_651 | v_198;
assign x_6264 = ~v_651 | v_34;
assign x_6265 = ~v_651 | ~v_42;
assign x_6266 = ~v_650 | v_199;
assign x_6267 = ~v_650 | v_34;
assign x_6268 = ~v_650 | ~v_43;
assign x_6269 = ~v_649 | v_191;
assign x_6270 = ~v_649 | v_34;
assign x_6271 = ~v_649 | ~v_35;
assign x_6272 = ~v_648 | v_200;
assign x_6273 = ~v_648 | v_35;
assign x_6274 = ~v_648 | ~v_36;
assign x_6275 = ~v_647 | v_201;
assign x_6276 = ~v_647 | v_35;
assign x_6277 = ~v_647 | ~v_37;
assign x_6278 = ~v_646 | v_202;
assign x_6279 = ~v_646 | v_35;
assign x_6280 = ~v_646 | ~v_38;
assign x_6281 = ~v_645 | v_203;
assign x_6282 = ~v_645 | v_35;
assign x_6283 = ~v_645 | ~v_39;
assign x_6284 = ~v_644 | v_204;
assign x_6285 = ~v_644 | v_35;
assign x_6286 = ~v_644 | ~v_40;
assign x_6287 = ~v_643 | v_205;
assign x_6288 = ~v_643 | v_35;
assign x_6289 = ~v_643 | ~v_41;
assign x_6290 = ~v_642 | v_206;
assign x_6291 = ~v_642 | v_35;
assign x_6292 = ~v_642 | ~v_42;
assign x_6293 = ~v_641 | v_207;
assign x_6294 = ~v_641 | v_35;
assign x_6295 = ~v_641 | ~v_43;
assign x_6296 = ~v_640 | v_192;
assign x_6297 = ~v_640 | v_34;
assign x_6298 = ~v_640 | ~v_36;
assign x_6299 = ~v_639 | v_200;
assign x_6300 = ~v_639 | v_35;
assign x_6301 = ~v_639 | ~v_36;
assign x_6302 = ~v_638 | v_208;
assign x_6303 = ~v_638 | v_36;
assign x_6304 = ~v_638 | ~v_37;
assign x_6305 = ~v_637 | v_209;
assign x_6306 = ~v_637 | v_36;
assign x_6307 = ~v_637 | ~v_38;
assign x_6308 = ~v_636 | v_210;
assign x_6309 = ~v_636 | v_36;
assign x_6310 = ~v_636 | ~v_39;
assign x_6311 = ~v_635 | v_211;
assign x_6312 = ~v_635 | v_36;
assign x_6313 = ~v_635 | ~v_40;
assign x_6314 = ~v_634 | v_212;
assign x_6315 = ~v_634 | v_36;
assign x_6316 = ~v_634 | ~v_41;
assign x_6317 = ~v_633 | v_213;
assign x_6318 = ~v_633 | v_36;
assign x_6319 = ~v_633 | ~v_42;
assign x_6320 = ~v_632 | v_214;
assign x_6321 = ~v_632 | v_36;
assign x_6322 = ~v_632 | ~v_43;
assign x_6323 = ~v_631 | v_193;
assign x_6324 = ~v_631 | v_34;
assign x_6325 = ~v_631 | ~v_37;
assign x_6326 = ~v_630 | v_201;
assign x_6327 = ~v_630 | v_35;
assign x_6328 = ~v_630 | ~v_37;
assign x_6329 = ~v_629 | v_208;
assign x_6330 = ~v_629 | v_36;
assign x_6331 = ~v_629 | ~v_37;
assign x_6332 = ~v_628 | v_215;
assign x_6333 = ~v_628 | v_37;
assign x_6334 = ~v_628 | ~v_38;
assign x_6335 = ~v_627 | v_216;
assign x_6336 = ~v_627 | v_37;
assign x_6337 = ~v_627 | ~v_39;
assign x_6338 = ~v_626 | v_217;
assign x_6339 = ~v_626 | v_37;
assign x_6340 = ~v_626 | ~v_40;
assign x_6341 = ~v_625 | v_218;
assign x_6342 = ~v_625 | v_37;
assign x_6343 = ~v_625 | ~v_41;
assign x_6344 = ~v_624 | v_219;
assign x_6345 = ~v_624 | v_37;
assign x_6346 = ~v_624 | ~v_42;
assign x_6347 = ~v_623 | v_220;
assign x_6348 = ~v_623 | v_37;
assign x_6349 = ~v_623 | ~v_43;
assign x_6350 = ~v_622 | v_194;
assign x_6351 = ~v_622 | v_34;
assign x_6352 = ~v_622 | ~v_38;
assign x_6353 = ~v_621 | v_202;
assign x_6354 = ~v_621 | v_35;
assign x_6355 = ~v_621 | ~v_38;
assign x_6356 = ~v_620 | v_209;
assign x_6357 = ~v_620 | v_36;
assign x_6358 = ~v_620 | ~v_38;
assign x_6359 = ~v_619 | v_215;
assign x_6360 = ~v_619 | v_37;
assign x_6361 = ~v_619 | ~v_38;
assign x_6362 = ~v_618 | v_221;
assign x_6363 = ~v_618 | v_38;
assign x_6364 = ~v_618 | ~v_39;
assign x_6365 = ~v_617 | v_222;
assign x_6366 = ~v_617 | v_38;
assign x_6367 = ~v_617 | ~v_40;
assign x_6368 = ~v_616 | v_223;
assign x_6369 = ~v_616 | v_38;
assign x_6370 = ~v_616 | ~v_41;
assign x_6371 = ~v_615 | v_224;
assign x_6372 = ~v_615 | v_38;
assign x_6373 = ~v_615 | ~v_42;
assign x_6374 = ~v_614 | v_225;
assign x_6375 = ~v_614 | v_38;
assign x_6376 = ~v_614 | ~v_43;
assign x_6377 = ~v_613 | v_195;
assign x_6378 = ~v_613 | v_34;
assign x_6379 = ~v_613 | ~v_39;
assign x_6380 = ~v_612 | v_203;
assign x_6381 = ~v_612 | v_35;
assign x_6382 = ~v_612 | ~v_39;
assign x_6383 = ~v_611 | v_210;
assign x_6384 = ~v_611 | v_36;
assign x_6385 = ~v_611 | ~v_39;
assign x_6386 = ~v_610 | v_216;
assign x_6387 = ~v_610 | v_37;
assign x_6388 = ~v_610 | ~v_39;
assign x_6389 = ~v_609 | v_221;
assign x_6390 = ~v_609 | v_38;
assign x_6391 = ~v_609 | ~v_39;
assign x_6392 = ~v_608 | v_226;
assign x_6393 = ~v_608 | v_39;
assign x_6394 = ~v_608 | ~v_40;
assign x_6395 = ~v_607 | v_227;
assign x_6396 = ~v_607 | v_39;
assign x_6397 = ~v_607 | ~v_41;
assign x_6398 = ~v_606 | v_228;
assign x_6399 = ~v_606 | v_39;
assign x_6400 = ~v_606 | ~v_42;
assign x_6401 = ~v_605 | v_229;
assign x_6402 = ~v_605 | v_39;
assign x_6403 = ~v_605 | ~v_43;
assign x_6404 = ~v_604 | v_196;
assign x_6405 = ~v_604 | v_34;
assign x_6406 = ~v_604 | ~v_40;
assign x_6407 = ~v_603 | v_204;
assign x_6408 = ~v_603 | v_35;
assign x_6409 = ~v_603 | ~v_40;
assign x_6410 = ~v_602 | v_211;
assign x_6411 = ~v_602 | v_36;
assign x_6412 = ~v_602 | ~v_40;
assign x_6413 = ~v_601 | v_217;
assign x_6414 = ~v_601 | v_37;
assign x_6415 = ~v_601 | ~v_40;
assign x_6416 = ~v_600 | v_222;
assign x_6417 = ~v_600 | v_38;
assign x_6418 = ~v_600 | ~v_40;
assign x_6419 = ~v_599 | v_226;
assign x_6420 = ~v_599 | v_39;
assign x_6421 = ~v_599 | ~v_40;
assign x_6422 = ~v_598 | v_230;
assign x_6423 = ~v_598 | v_40;
assign x_6424 = ~v_598 | ~v_41;
assign x_6425 = ~v_597 | v_231;
assign x_6426 = ~v_597 | v_40;
assign x_6427 = ~v_597 | ~v_42;
assign x_6428 = ~v_596 | v_232;
assign x_6429 = ~v_596 | v_40;
assign x_6430 = ~v_596 | ~v_43;
assign x_6431 = ~v_595 | v_197;
assign x_6432 = ~v_595 | v_34;
assign x_6433 = ~v_595 | ~v_41;
assign x_6434 = ~v_594 | v_205;
assign x_6435 = ~v_594 | v_35;
assign x_6436 = ~v_594 | ~v_41;
assign x_6437 = ~v_593 | v_212;
assign x_6438 = ~v_593 | v_36;
assign x_6439 = ~v_593 | ~v_41;
assign x_6440 = ~v_592 | v_218;
assign x_6441 = ~v_592 | v_37;
assign x_6442 = ~v_592 | ~v_41;
assign x_6443 = ~v_591 | v_223;
assign x_6444 = ~v_591 | v_38;
assign x_6445 = ~v_591 | ~v_41;
assign x_6446 = ~v_590 | v_227;
assign x_6447 = ~v_590 | v_39;
assign x_6448 = ~v_590 | ~v_41;
assign x_6449 = ~v_589 | v_230;
assign x_6450 = ~v_589 | v_40;
assign x_6451 = ~v_589 | ~v_41;
assign x_6452 = ~v_588 | v_233;
assign x_6453 = ~v_588 | v_41;
assign x_6454 = ~v_588 | ~v_42;
assign x_6455 = ~v_587 | v_234;
assign x_6456 = ~v_587 | v_41;
assign x_6457 = ~v_587 | ~v_43;
assign x_6458 = ~v_586 | v_198;
assign x_6459 = ~v_586 | v_34;
assign x_6460 = ~v_586 | ~v_42;
assign x_6461 = ~v_585 | v_206;
assign x_6462 = ~v_585 | v_35;
assign x_6463 = ~v_585 | ~v_42;
assign x_6464 = ~v_584 | v_213;
assign x_6465 = ~v_584 | v_36;
assign x_6466 = ~v_584 | ~v_42;
assign x_6467 = ~v_583 | v_219;
assign x_6468 = ~v_583 | v_37;
assign x_6469 = ~v_583 | ~v_42;
assign x_6470 = ~v_582 | v_224;
assign x_6471 = ~v_582 | v_38;
assign x_6472 = ~v_582 | ~v_42;
assign x_6473 = ~v_581 | v_228;
assign x_6474 = ~v_581 | v_39;
assign x_6475 = ~v_581 | ~v_42;
assign x_6476 = ~v_580 | v_231;
assign x_6477 = ~v_580 | v_40;
assign x_6478 = ~v_580 | ~v_42;
assign x_6479 = ~v_579 | v_233;
assign x_6480 = ~v_579 | v_41;
assign x_6481 = ~v_579 | ~v_42;
assign x_6482 = ~v_578 | v_235;
assign x_6483 = ~v_578 | v_42;
assign x_6484 = ~v_578 | ~v_43;
assign x_6485 = ~v_577 | v_199;
assign x_6486 = ~v_577 | v_34;
assign x_6487 = ~v_577 | ~v_43;
assign x_6488 = ~v_576 | v_207;
assign x_6489 = ~v_576 | v_35;
assign x_6490 = ~v_576 | ~v_43;
assign x_6491 = ~v_575 | v_214;
assign x_6492 = ~v_575 | v_36;
assign x_6493 = ~v_575 | ~v_43;
assign x_6494 = ~v_574 | v_220;
assign x_6495 = ~v_574 | v_37;
assign x_6496 = ~v_574 | ~v_43;
assign x_6497 = ~v_573 | v_225;
assign x_6498 = ~v_573 | v_38;
assign x_6499 = ~v_573 | ~v_43;
assign x_6500 = ~v_572 | v_229;
assign x_6501 = ~v_572 | v_39;
assign x_6502 = ~v_572 | ~v_43;
assign x_6503 = ~v_571 | v_232;
assign x_6504 = ~v_571 | v_40;
assign x_6505 = ~v_571 | ~v_43;
assign x_6506 = ~v_570 | v_234;
assign x_6507 = ~v_570 | v_41;
assign x_6508 = ~v_570 | ~v_43;
assign x_6509 = ~v_569 | v_235;
assign x_6510 = ~v_569 | v_42;
assign x_6511 = ~v_569 | ~v_43;
assign x_6512 = ~v_567 | ~v_191 | ~v_34 | v_35;
assign x_6513 = ~v_568 | ~v_45;
assign x_6514 = ~v_568 | v_46;
assign x_6515 = ~v_565 | ~v_192 | ~v_34 | v_36;
assign x_6516 = ~v_566 | ~v_45;
assign x_6517 = ~v_566 | v_47;
assign x_6518 = ~v_563 | ~v_193 | ~v_34 | v_37;
assign x_6519 = ~v_564 | ~v_45;
assign x_6520 = ~v_564 | v_48;
assign x_6521 = ~v_561 | ~v_194 | ~v_34 | v_38;
assign x_6522 = ~v_562 | ~v_45;
assign x_6523 = ~v_562 | v_49;
assign x_6524 = ~v_559 | ~v_195 | ~v_34 | v_39;
assign x_6525 = ~v_560 | ~v_45;
assign x_6526 = ~v_560 | v_50;
assign x_6527 = ~v_557 | ~v_196 | ~v_34 | v_40;
assign x_6528 = ~v_558 | ~v_45;
assign x_6529 = ~v_558 | v_51;
assign x_6530 = ~v_555 | ~v_197 | ~v_34 | v_41;
assign x_6531 = ~v_556 | ~v_45;
assign x_6532 = ~v_556 | v_52;
assign x_6533 = ~v_553 | ~v_198 | ~v_34 | v_42;
assign x_6534 = ~v_554 | ~v_45;
assign x_6535 = ~v_554 | v_53;
assign x_6536 = ~v_551 | ~v_199 | ~v_34 | v_43;
assign x_6537 = ~v_552 | ~v_45;
assign x_6538 = ~v_552 | v_54;
assign x_6539 = ~v_549 | ~v_200 | ~v_35 | v_36;
assign x_6540 = ~v_550 | ~v_46;
assign x_6541 = ~v_550 | v_47;
assign x_6542 = ~v_547 | ~v_201 | ~v_35 | v_37;
assign x_6543 = ~v_548 | ~v_46;
assign x_6544 = ~v_548 | v_48;
assign x_6545 = ~v_545 | ~v_202 | ~v_35 | v_38;
assign x_6546 = ~v_546 | ~v_46;
assign x_6547 = ~v_546 | v_49;
assign x_6548 = ~v_543 | ~v_203 | ~v_35 | v_39;
assign x_6549 = ~v_544 | ~v_46;
assign x_6550 = ~v_544 | v_50;
assign x_6551 = ~v_541 | ~v_204 | ~v_35 | v_40;
assign x_6552 = ~v_542 | ~v_46;
assign x_6553 = ~v_542 | v_51;
assign x_6554 = ~v_539 | ~v_205 | ~v_35 | v_41;
assign x_6555 = ~v_540 | ~v_46;
assign x_6556 = ~v_540 | v_52;
assign x_6557 = ~v_537 | ~v_206 | ~v_35 | v_42;
assign x_6558 = ~v_538 | ~v_46;
assign x_6559 = ~v_538 | v_53;
assign x_6560 = ~v_535 | ~v_207 | ~v_35 | v_43;
assign x_6561 = ~v_536 | ~v_46;
assign x_6562 = ~v_536 | v_54;
assign x_6563 = ~v_533 | ~v_208 | ~v_36 | v_37;
assign x_6564 = ~v_534 | ~v_47;
assign x_6565 = ~v_534 | v_48;
assign x_6566 = ~v_531 | ~v_209 | ~v_36 | v_38;
assign x_6567 = ~v_532 | ~v_47;
assign x_6568 = ~v_532 | v_49;
assign x_6569 = ~v_529 | ~v_210 | ~v_36 | v_39;
assign x_6570 = ~v_530 | ~v_47;
assign x_6571 = ~v_530 | v_50;
assign x_6572 = ~v_527 | ~v_211 | ~v_36 | v_40;
assign x_6573 = ~v_528 | ~v_47;
assign x_6574 = ~v_528 | v_51;
assign x_6575 = ~v_525 | ~v_212 | ~v_36 | v_41;
assign x_6576 = ~v_526 | ~v_47;
assign x_6577 = ~v_526 | v_52;
assign x_6578 = ~v_523 | ~v_213 | ~v_36 | v_42;
assign x_6579 = ~v_524 | ~v_47;
assign x_6580 = ~v_524 | v_53;
assign x_6581 = ~v_521 | ~v_214 | ~v_36 | v_43;
assign x_6582 = ~v_522 | ~v_47;
assign x_6583 = ~v_522 | v_54;
assign x_6584 = ~v_519 | ~v_215 | ~v_37 | v_38;
assign x_6585 = ~v_520 | ~v_48;
assign x_6586 = ~v_520 | v_49;
assign x_6587 = ~v_517 | ~v_216 | ~v_37 | v_39;
assign x_6588 = ~v_518 | ~v_48;
assign x_6589 = ~v_518 | v_50;
assign x_6590 = ~v_515 | ~v_217 | ~v_37 | v_40;
assign x_6591 = ~v_516 | ~v_48;
assign x_6592 = ~v_516 | v_51;
assign x_6593 = ~v_513 | ~v_218 | ~v_37 | v_41;
assign x_6594 = ~v_514 | ~v_48;
assign x_6595 = ~v_514 | v_52;
assign x_6596 = ~v_511 | ~v_219 | ~v_37 | v_42;
assign x_6597 = ~v_512 | ~v_48;
assign x_6598 = ~v_512 | v_53;
assign x_6599 = ~v_509 | ~v_220 | ~v_37 | v_43;
assign x_6600 = ~v_510 | ~v_48;
assign x_6601 = ~v_510 | v_54;
assign x_6602 = ~v_507 | ~v_221 | ~v_38 | v_39;
assign x_6603 = ~v_508 | ~v_49;
assign x_6604 = ~v_508 | v_50;
assign x_6605 = ~v_505 | ~v_222 | ~v_38 | v_40;
assign x_6606 = ~v_506 | ~v_49;
assign x_6607 = ~v_506 | v_51;
assign x_6608 = ~v_503 | ~v_223 | ~v_38 | v_41;
assign x_6609 = ~v_504 | ~v_49;
assign x_6610 = ~v_504 | v_52;
assign x_6611 = ~v_501 | ~v_224 | ~v_38 | v_42;
assign x_6612 = ~v_502 | ~v_49;
assign x_6613 = ~v_502 | v_53;
assign x_6614 = ~v_499 | ~v_225 | ~v_38 | v_43;
assign x_6615 = ~v_500 | ~v_49;
assign x_6616 = ~v_500 | v_54;
assign x_6617 = ~v_497 | ~v_226 | ~v_39 | v_40;
assign x_6618 = ~v_498 | ~v_50;
assign x_6619 = ~v_498 | v_51;
assign x_6620 = ~v_495 | ~v_227 | ~v_39 | v_41;
assign x_6621 = ~v_496 | ~v_50;
assign x_6622 = ~v_496 | v_52;
assign x_6623 = ~v_493 | ~v_228 | ~v_39 | v_42;
assign x_6624 = ~v_494 | ~v_50;
assign x_6625 = ~v_494 | v_53;
assign x_6626 = ~v_491 | ~v_229 | ~v_39 | v_43;
assign x_6627 = ~v_492 | ~v_50;
assign x_6628 = ~v_492 | v_54;
assign x_6629 = ~v_489 | ~v_230 | ~v_40 | v_41;
assign x_6630 = ~v_490 | ~v_51;
assign x_6631 = ~v_490 | v_52;
assign x_6632 = ~v_487 | ~v_231 | ~v_40 | v_42;
assign x_6633 = ~v_488 | ~v_51;
assign x_6634 = ~v_488 | v_53;
assign x_6635 = ~v_485 | ~v_232 | ~v_40 | v_43;
assign x_6636 = ~v_486 | ~v_51;
assign x_6637 = ~v_486 | v_54;
assign x_6638 = ~v_483 | ~v_233 | ~v_41 | v_42;
assign x_6639 = ~v_484 | ~v_52;
assign x_6640 = ~v_484 | v_53;
assign x_6641 = ~v_481 | ~v_234 | ~v_41 | v_43;
assign x_6642 = ~v_482 | ~v_52;
assign x_6643 = ~v_482 | v_54;
assign x_6644 = ~v_479 | ~v_235 | ~v_42 | v_43;
assign x_6645 = ~v_480 | ~v_53;
assign x_6646 = ~v_480 | v_54;
assign x_6647 = ~v_470 | v_45;
assign x_6648 = ~v_470 | ~v_46;
assign x_6649 = ~v_471 | v_46;
assign x_6650 = ~v_471 | ~v_47;
assign x_6651 = ~v_472 | v_47;
assign x_6652 = ~v_472 | ~v_48;
assign x_6653 = ~v_473 | v_48;
assign x_6654 = ~v_473 | ~v_49;
assign x_6655 = ~v_474 | v_49;
assign x_6656 = ~v_474 | ~v_50;
assign x_6657 = ~v_475 | v_50;
assign x_6658 = ~v_475 | ~v_51;
assign x_6659 = ~v_476 | v_51;
assign x_6660 = ~v_476 | ~v_52;
assign x_6661 = ~v_477 | v_52;
assign x_6662 = ~v_477 | ~v_53;
assign x_6663 = ~v_478 | v_53;
assign x_6664 = ~v_478 | ~v_54;
assign x_6665 = x_2 & x_3;
assign x_6666 = x_1 & x_6665;
assign x_6667 = x_5 & x_6;
assign x_6668 = x_4 & x_6667;
assign x_6669 = x_6666 & x_6668;
assign x_6670 = x_8 & x_9;
assign x_6671 = x_7 & x_6670;
assign x_6672 = x_10 & x_11;
assign x_6673 = x_12 & x_13;
assign x_6674 = x_6672 & x_6673;
assign x_6675 = x_6671 & x_6674;
assign x_6676 = x_6669 & x_6675;
assign x_6677 = x_15 & x_16;
assign x_6678 = x_14 & x_6677;
assign x_6679 = x_18 & x_19;
assign x_6680 = x_17 & x_6679;
assign x_6681 = x_6678 & x_6680;
assign x_6682 = x_21 & x_22;
assign x_6683 = x_20 & x_6682;
assign x_6684 = x_23 & x_24;
assign x_6685 = x_25 & x_26;
assign x_6686 = x_6684 & x_6685;
assign x_6687 = x_6683 & x_6686;
assign x_6688 = x_6681 & x_6687;
assign x_6689 = x_6676 & x_6688;
assign x_6690 = x_28 & x_29;
assign x_6691 = x_27 & x_6690;
assign x_6692 = x_31 & x_32;
assign x_6693 = x_30 & x_6692;
assign x_6694 = x_6691 & x_6693;
assign x_6695 = x_34 & x_35;
assign x_6696 = x_33 & x_6695;
assign x_6697 = x_36 & x_37;
assign x_6698 = x_38 & x_39;
assign x_6699 = x_6697 & x_6698;
assign x_6700 = x_6696 & x_6699;
assign x_6701 = x_6694 & x_6700;
assign x_6702 = x_41 & x_42;
assign x_6703 = x_40 & x_6702;
assign x_6704 = x_44 & x_45;
assign x_6705 = x_43 & x_6704;
assign x_6706 = x_6703 & x_6705;
assign x_6707 = x_47 & x_48;
assign x_6708 = x_46 & x_6707;
assign x_6709 = x_49 & x_50;
assign x_6710 = x_51 & x_52;
assign x_6711 = x_6709 & x_6710;
assign x_6712 = x_6708 & x_6711;
assign x_6713 = x_6706 & x_6712;
assign x_6714 = x_6701 & x_6713;
assign x_6715 = x_6689 & x_6714;
assign x_6716 = x_54 & x_55;
assign x_6717 = x_53 & x_6716;
assign x_6718 = x_57 & x_58;
assign x_6719 = x_56 & x_6718;
assign x_6720 = x_6717 & x_6719;
assign x_6721 = x_60 & x_61;
assign x_6722 = x_59 & x_6721;
assign x_6723 = x_62 & x_63;
assign x_6724 = x_64 & x_65;
assign x_6725 = x_6723 & x_6724;
assign x_6726 = x_6722 & x_6725;
assign x_6727 = x_6720 & x_6726;
assign x_6728 = x_67 & x_68;
assign x_6729 = x_66 & x_6728;
assign x_6730 = x_70 & x_71;
assign x_6731 = x_69 & x_6730;
assign x_6732 = x_6729 & x_6731;
assign x_6733 = x_73 & x_74;
assign x_6734 = x_72 & x_6733;
assign x_6735 = x_75 & x_76;
assign x_6736 = x_77 & x_78;
assign x_6737 = x_6735 & x_6736;
assign x_6738 = x_6734 & x_6737;
assign x_6739 = x_6732 & x_6738;
assign x_6740 = x_6727 & x_6739;
assign x_6741 = x_80 & x_81;
assign x_6742 = x_79 & x_6741;
assign x_6743 = x_83 & x_84;
assign x_6744 = x_82 & x_6743;
assign x_6745 = x_6742 & x_6744;
assign x_6746 = x_86 & x_87;
assign x_6747 = x_85 & x_6746;
assign x_6748 = x_88 & x_89;
assign x_6749 = x_90 & x_91;
assign x_6750 = x_6748 & x_6749;
assign x_6751 = x_6747 & x_6750;
assign x_6752 = x_6745 & x_6751;
assign x_6753 = x_93 & x_94;
assign x_6754 = x_92 & x_6753;
assign x_6755 = x_96 & x_97;
assign x_6756 = x_95 & x_6755;
assign x_6757 = x_6754 & x_6756;
assign x_6758 = x_99 & x_100;
assign x_6759 = x_98 & x_6758;
assign x_6760 = x_101 & x_102;
assign x_6761 = x_103 & x_104;
assign x_6762 = x_6760 & x_6761;
assign x_6763 = x_6759 & x_6762;
assign x_6764 = x_6757 & x_6763;
assign x_6765 = x_6752 & x_6764;
assign x_6766 = x_6740 & x_6765;
assign x_6767 = x_6715 & x_6766;
assign x_6768 = x_106 & x_107;
assign x_6769 = x_105 & x_6768;
assign x_6770 = x_109 & x_110;
assign x_6771 = x_108 & x_6770;
assign x_6772 = x_6769 & x_6771;
assign x_6773 = x_112 & x_113;
assign x_6774 = x_111 & x_6773;
assign x_6775 = x_114 & x_115;
assign x_6776 = x_116 & x_117;
assign x_6777 = x_6775 & x_6776;
assign x_6778 = x_6774 & x_6777;
assign x_6779 = x_6772 & x_6778;
assign x_6780 = x_119 & x_120;
assign x_6781 = x_118 & x_6780;
assign x_6782 = x_122 & x_123;
assign x_6783 = x_121 & x_6782;
assign x_6784 = x_6781 & x_6783;
assign x_6785 = x_125 & x_126;
assign x_6786 = x_124 & x_6785;
assign x_6787 = x_127 & x_128;
assign x_6788 = x_129 & x_130;
assign x_6789 = x_6787 & x_6788;
assign x_6790 = x_6786 & x_6789;
assign x_6791 = x_6784 & x_6790;
assign x_6792 = x_6779 & x_6791;
assign x_6793 = x_132 & x_133;
assign x_6794 = x_131 & x_6793;
assign x_6795 = x_135 & x_136;
assign x_6796 = x_134 & x_6795;
assign x_6797 = x_6794 & x_6796;
assign x_6798 = x_138 & x_139;
assign x_6799 = x_137 & x_6798;
assign x_6800 = x_140 & x_141;
assign x_6801 = x_142 & x_143;
assign x_6802 = x_6800 & x_6801;
assign x_6803 = x_6799 & x_6802;
assign x_6804 = x_6797 & x_6803;
assign x_6805 = x_145 & x_146;
assign x_6806 = x_144 & x_6805;
assign x_6807 = x_148 & x_149;
assign x_6808 = x_147 & x_6807;
assign x_6809 = x_6806 & x_6808;
assign x_6810 = x_151 & x_152;
assign x_6811 = x_150 & x_6810;
assign x_6812 = x_153 & x_154;
assign x_6813 = x_155 & x_156;
assign x_6814 = x_6812 & x_6813;
assign x_6815 = x_6811 & x_6814;
assign x_6816 = x_6809 & x_6815;
assign x_6817 = x_6804 & x_6816;
assign x_6818 = x_6792 & x_6817;
assign x_6819 = x_158 & x_159;
assign x_6820 = x_157 & x_6819;
assign x_6821 = x_161 & x_162;
assign x_6822 = x_160 & x_6821;
assign x_6823 = x_6820 & x_6822;
assign x_6824 = x_164 & x_165;
assign x_6825 = x_163 & x_6824;
assign x_6826 = x_166 & x_167;
assign x_6827 = x_168 & x_169;
assign x_6828 = x_6826 & x_6827;
assign x_6829 = x_6825 & x_6828;
assign x_6830 = x_6823 & x_6829;
assign x_6831 = x_171 & x_172;
assign x_6832 = x_170 & x_6831;
assign x_6833 = x_174 & x_175;
assign x_6834 = x_173 & x_6833;
assign x_6835 = x_6832 & x_6834;
assign x_6836 = x_177 & x_178;
assign x_6837 = x_176 & x_6836;
assign x_6838 = x_179 & x_180;
assign x_6839 = x_181 & x_182;
assign x_6840 = x_6838 & x_6839;
assign x_6841 = x_6837 & x_6840;
assign x_6842 = x_6835 & x_6841;
assign x_6843 = x_6830 & x_6842;
assign x_6844 = x_184 & x_185;
assign x_6845 = x_183 & x_6844;
assign x_6846 = x_187 & x_188;
assign x_6847 = x_186 & x_6846;
assign x_6848 = x_6845 & x_6847;
assign x_6849 = x_190 & x_191;
assign x_6850 = x_189 & x_6849;
assign x_6851 = x_192 & x_193;
assign x_6852 = x_194 & x_195;
assign x_6853 = x_6851 & x_6852;
assign x_6854 = x_6850 & x_6853;
assign x_6855 = x_6848 & x_6854;
assign x_6856 = x_197 & x_198;
assign x_6857 = x_196 & x_6856;
assign x_6858 = x_200 & x_201;
assign x_6859 = x_199 & x_6858;
assign x_6860 = x_6857 & x_6859;
assign x_6861 = x_203 & x_204;
assign x_6862 = x_202 & x_6861;
assign x_6863 = x_205 & x_206;
assign x_6864 = x_207 & x_208;
assign x_6865 = x_6863 & x_6864;
assign x_6866 = x_6862 & x_6865;
assign x_6867 = x_6860 & x_6866;
assign x_6868 = x_6855 & x_6867;
assign x_6869 = x_6843 & x_6868;
assign x_6870 = x_6818 & x_6869;
assign x_6871 = x_6767 & x_6870;
assign x_6872 = x_210 & x_211;
assign x_6873 = x_209 & x_6872;
assign x_6874 = x_213 & x_214;
assign x_6875 = x_212 & x_6874;
assign x_6876 = x_6873 & x_6875;
assign x_6877 = x_216 & x_217;
assign x_6878 = x_215 & x_6877;
assign x_6879 = x_218 & x_219;
assign x_6880 = x_220 & x_221;
assign x_6881 = x_6879 & x_6880;
assign x_6882 = x_6878 & x_6881;
assign x_6883 = x_6876 & x_6882;
assign x_6884 = x_223 & x_224;
assign x_6885 = x_222 & x_6884;
assign x_6886 = x_226 & x_227;
assign x_6887 = x_225 & x_6886;
assign x_6888 = x_6885 & x_6887;
assign x_6889 = x_229 & x_230;
assign x_6890 = x_228 & x_6889;
assign x_6891 = x_231 & x_232;
assign x_6892 = x_233 & x_234;
assign x_6893 = x_6891 & x_6892;
assign x_6894 = x_6890 & x_6893;
assign x_6895 = x_6888 & x_6894;
assign x_6896 = x_6883 & x_6895;
assign x_6897 = x_236 & x_237;
assign x_6898 = x_235 & x_6897;
assign x_6899 = x_239 & x_240;
assign x_6900 = x_238 & x_6899;
assign x_6901 = x_6898 & x_6900;
assign x_6902 = x_242 & x_243;
assign x_6903 = x_241 & x_6902;
assign x_6904 = x_244 & x_245;
assign x_6905 = x_246 & x_247;
assign x_6906 = x_6904 & x_6905;
assign x_6907 = x_6903 & x_6906;
assign x_6908 = x_6901 & x_6907;
assign x_6909 = x_249 & x_250;
assign x_6910 = x_248 & x_6909;
assign x_6911 = x_252 & x_253;
assign x_6912 = x_251 & x_6911;
assign x_6913 = x_6910 & x_6912;
assign x_6914 = x_255 & x_256;
assign x_6915 = x_254 & x_6914;
assign x_6916 = x_257 & x_258;
assign x_6917 = x_259 & x_260;
assign x_6918 = x_6916 & x_6917;
assign x_6919 = x_6915 & x_6918;
assign x_6920 = x_6913 & x_6919;
assign x_6921 = x_6908 & x_6920;
assign x_6922 = x_6896 & x_6921;
assign x_6923 = x_262 & x_263;
assign x_6924 = x_261 & x_6923;
assign x_6925 = x_265 & x_266;
assign x_6926 = x_264 & x_6925;
assign x_6927 = x_6924 & x_6926;
assign x_6928 = x_268 & x_269;
assign x_6929 = x_267 & x_6928;
assign x_6930 = x_270 & x_271;
assign x_6931 = x_272 & x_273;
assign x_6932 = x_6930 & x_6931;
assign x_6933 = x_6929 & x_6932;
assign x_6934 = x_6927 & x_6933;
assign x_6935 = x_275 & x_276;
assign x_6936 = x_274 & x_6935;
assign x_6937 = x_278 & x_279;
assign x_6938 = x_277 & x_6937;
assign x_6939 = x_6936 & x_6938;
assign x_6940 = x_281 & x_282;
assign x_6941 = x_280 & x_6940;
assign x_6942 = x_283 & x_284;
assign x_6943 = x_285 & x_286;
assign x_6944 = x_6942 & x_6943;
assign x_6945 = x_6941 & x_6944;
assign x_6946 = x_6939 & x_6945;
assign x_6947 = x_6934 & x_6946;
assign x_6948 = x_288 & x_289;
assign x_6949 = x_287 & x_6948;
assign x_6950 = x_291 & x_292;
assign x_6951 = x_290 & x_6950;
assign x_6952 = x_6949 & x_6951;
assign x_6953 = x_294 & x_295;
assign x_6954 = x_293 & x_6953;
assign x_6955 = x_296 & x_297;
assign x_6956 = x_298 & x_299;
assign x_6957 = x_6955 & x_6956;
assign x_6958 = x_6954 & x_6957;
assign x_6959 = x_6952 & x_6958;
assign x_6960 = x_301 & x_302;
assign x_6961 = x_300 & x_6960;
assign x_6962 = x_304 & x_305;
assign x_6963 = x_303 & x_6962;
assign x_6964 = x_6961 & x_6963;
assign x_6965 = x_307 & x_308;
assign x_6966 = x_306 & x_6965;
assign x_6967 = x_309 & x_310;
assign x_6968 = x_311 & x_312;
assign x_6969 = x_6967 & x_6968;
assign x_6970 = x_6966 & x_6969;
assign x_6971 = x_6964 & x_6970;
assign x_6972 = x_6959 & x_6971;
assign x_6973 = x_6947 & x_6972;
assign x_6974 = x_6922 & x_6973;
assign x_6975 = x_314 & x_315;
assign x_6976 = x_313 & x_6975;
assign x_6977 = x_317 & x_318;
assign x_6978 = x_316 & x_6977;
assign x_6979 = x_6976 & x_6978;
assign x_6980 = x_320 & x_321;
assign x_6981 = x_319 & x_6980;
assign x_6982 = x_322 & x_323;
assign x_6983 = x_324 & x_325;
assign x_6984 = x_6982 & x_6983;
assign x_6985 = x_6981 & x_6984;
assign x_6986 = x_6979 & x_6985;
assign x_6987 = x_327 & x_328;
assign x_6988 = x_326 & x_6987;
assign x_6989 = x_330 & x_331;
assign x_6990 = x_329 & x_6989;
assign x_6991 = x_6988 & x_6990;
assign x_6992 = x_333 & x_334;
assign x_6993 = x_332 & x_6992;
assign x_6994 = x_335 & x_336;
assign x_6995 = x_337 & x_338;
assign x_6996 = x_6994 & x_6995;
assign x_6997 = x_6993 & x_6996;
assign x_6998 = x_6991 & x_6997;
assign x_6999 = x_6986 & x_6998;
assign x_7000 = x_340 & x_341;
assign x_7001 = x_339 & x_7000;
assign x_7002 = x_343 & x_344;
assign x_7003 = x_342 & x_7002;
assign x_7004 = x_7001 & x_7003;
assign x_7005 = x_346 & x_347;
assign x_7006 = x_345 & x_7005;
assign x_7007 = x_348 & x_349;
assign x_7008 = x_350 & x_351;
assign x_7009 = x_7007 & x_7008;
assign x_7010 = x_7006 & x_7009;
assign x_7011 = x_7004 & x_7010;
assign x_7012 = x_353 & x_354;
assign x_7013 = x_352 & x_7012;
assign x_7014 = x_356 & x_357;
assign x_7015 = x_355 & x_7014;
assign x_7016 = x_7013 & x_7015;
assign x_7017 = x_359 & x_360;
assign x_7018 = x_358 & x_7017;
assign x_7019 = x_361 & x_362;
assign x_7020 = x_363 & x_364;
assign x_7021 = x_7019 & x_7020;
assign x_7022 = x_7018 & x_7021;
assign x_7023 = x_7016 & x_7022;
assign x_7024 = x_7011 & x_7023;
assign x_7025 = x_6999 & x_7024;
assign x_7026 = x_366 & x_367;
assign x_7027 = x_365 & x_7026;
assign x_7028 = x_369 & x_370;
assign x_7029 = x_368 & x_7028;
assign x_7030 = x_7027 & x_7029;
assign x_7031 = x_372 & x_373;
assign x_7032 = x_371 & x_7031;
assign x_7033 = x_374 & x_375;
assign x_7034 = x_376 & x_377;
assign x_7035 = x_7033 & x_7034;
assign x_7036 = x_7032 & x_7035;
assign x_7037 = x_7030 & x_7036;
assign x_7038 = x_379 & x_380;
assign x_7039 = x_378 & x_7038;
assign x_7040 = x_382 & x_383;
assign x_7041 = x_381 & x_7040;
assign x_7042 = x_7039 & x_7041;
assign x_7043 = x_385 & x_386;
assign x_7044 = x_384 & x_7043;
assign x_7045 = x_387 & x_388;
assign x_7046 = x_389 & x_390;
assign x_7047 = x_7045 & x_7046;
assign x_7048 = x_7044 & x_7047;
assign x_7049 = x_7042 & x_7048;
assign x_7050 = x_7037 & x_7049;
assign x_7051 = x_392 & x_393;
assign x_7052 = x_391 & x_7051;
assign x_7053 = x_395 & x_396;
assign x_7054 = x_394 & x_7053;
assign x_7055 = x_7052 & x_7054;
assign x_7056 = x_398 & x_399;
assign x_7057 = x_397 & x_7056;
assign x_7058 = x_400 & x_401;
assign x_7059 = x_402 & x_403;
assign x_7060 = x_7058 & x_7059;
assign x_7061 = x_7057 & x_7060;
assign x_7062 = x_7055 & x_7061;
assign x_7063 = x_405 & x_406;
assign x_7064 = x_404 & x_7063;
assign x_7065 = x_408 & x_409;
assign x_7066 = x_407 & x_7065;
assign x_7067 = x_7064 & x_7066;
assign x_7068 = x_411 & x_412;
assign x_7069 = x_410 & x_7068;
assign x_7070 = x_413 & x_414;
assign x_7071 = x_415 & x_416;
assign x_7072 = x_7070 & x_7071;
assign x_7073 = x_7069 & x_7072;
assign x_7074 = x_7067 & x_7073;
assign x_7075 = x_7062 & x_7074;
assign x_7076 = x_7050 & x_7075;
assign x_7077 = x_7025 & x_7076;
assign x_7078 = x_6974 & x_7077;
assign x_7079 = x_6871 & x_7078;
assign x_7080 = x_418 & x_419;
assign x_7081 = x_417 & x_7080;
assign x_7082 = x_421 & x_422;
assign x_7083 = x_420 & x_7082;
assign x_7084 = x_7081 & x_7083;
assign x_7085 = x_424 & x_425;
assign x_7086 = x_423 & x_7085;
assign x_7087 = x_426 & x_427;
assign x_7088 = x_428 & x_429;
assign x_7089 = x_7087 & x_7088;
assign x_7090 = x_7086 & x_7089;
assign x_7091 = x_7084 & x_7090;
assign x_7092 = x_431 & x_432;
assign x_7093 = x_430 & x_7092;
assign x_7094 = x_434 & x_435;
assign x_7095 = x_433 & x_7094;
assign x_7096 = x_7093 & x_7095;
assign x_7097 = x_437 & x_438;
assign x_7098 = x_436 & x_7097;
assign x_7099 = x_439 & x_440;
assign x_7100 = x_441 & x_442;
assign x_7101 = x_7099 & x_7100;
assign x_7102 = x_7098 & x_7101;
assign x_7103 = x_7096 & x_7102;
assign x_7104 = x_7091 & x_7103;
assign x_7105 = x_444 & x_445;
assign x_7106 = x_443 & x_7105;
assign x_7107 = x_447 & x_448;
assign x_7108 = x_446 & x_7107;
assign x_7109 = x_7106 & x_7108;
assign x_7110 = x_450 & x_451;
assign x_7111 = x_449 & x_7110;
assign x_7112 = x_452 & x_453;
assign x_7113 = x_454 & x_455;
assign x_7114 = x_7112 & x_7113;
assign x_7115 = x_7111 & x_7114;
assign x_7116 = x_7109 & x_7115;
assign x_7117 = x_457 & x_458;
assign x_7118 = x_456 & x_7117;
assign x_7119 = x_460 & x_461;
assign x_7120 = x_459 & x_7119;
assign x_7121 = x_7118 & x_7120;
assign x_7122 = x_463 & x_464;
assign x_7123 = x_462 & x_7122;
assign x_7124 = x_465 & x_466;
assign x_7125 = x_467 & x_468;
assign x_7126 = x_7124 & x_7125;
assign x_7127 = x_7123 & x_7126;
assign x_7128 = x_7121 & x_7127;
assign x_7129 = x_7116 & x_7128;
assign x_7130 = x_7104 & x_7129;
assign x_7131 = x_470 & x_471;
assign x_7132 = x_469 & x_7131;
assign x_7133 = x_473 & x_474;
assign x_7134 = x_472 & x_7133;
assign x_7135 = x_7132 & x_7134;
assign x_7136 = x_476 & x_477;
assign x_7137 = x_475 & x_7136;
assign x_7138 = x_478 & x_479;
assign x_7139 = x_480 & x_481;
assign x_7140 = x_7138 & x_7139;
assign x_7141 = x_7137 & x_7140;
assign x_7142 = x_7135 & x_7141;
assign x_7143 = x_483 & x_484;
assign x_7144 = x_482 & x_7143;
assign x_7145 = x_486 & x_487;
assign x_7146 = x_485 & x_7145;
assign x_7147 = x_7144 & x_7146;
assign x_7148 = x_489 & x_490;
assign x_7149 = x_488 & x_7148;
assign x_7150 = x_491 & x_492;
assign x_7151 = x_493 & x_494;
assign x_7152 = x_7150 & x_7151;
assign x_7153 = x_7149 & x_7152;
assign x_7154 = x_7147 & x_7153;
assign x_7155 = x_7142 & x_7154;
assign x_7156 = x_496 & x_497;
assign x_7157 = x_495 & x_7156;
assign x_7158 = x_499 & x_500;
assign x_7159 = x_498 & x_7158;
assign x_7160 = x_7157 & x_7159;
assign x_7161 = x_502 & x_503;
assign x_7162 = x_501 & x_7161;
assign x_7163 = x_504 & x_505;
assign x_7164 = x_506 & x_507;
assign x_7165 = x_7163 & x_7164;
assign x_7166 = x_7162 & x_7165;
assign x_7167 = x_7160 & x_7166;
assign x_7168 = x_509 & x_510;
assign x_7169 = x_508 & x_7168;
assign x_7170 = x_512 & x_513;
assign x_7171 = x_511 & x_7170;
assign x_7172 = x_7169 & x_7171;
assign x_7173 = x_515 & x_516;
assign x_7174 = x_514 & x_7173;
assign x_7175 = x_517 & x_518;
assign x_7176 = x_519 & x_520;
assign x_7177 = x_7175 & x_7176;
assign x_7178 = x_7174 & x_7177;
assign x_7179 = x_7172 & x_7178;
assign x_7180 = x_7167 & x_7179;
assign x_7181 = x_7155 & x_7180;
assign x_7182 = x_7130 & x_7181;
assign x_7183 = x_522 & x_523;
assign x_7184 = x_521 & x_7183;
assign x_7185 = x_525 & x_526;
assign x_7186 = x_524 & x_7185;
assign x_7187 = x_7184 & x_7186;
assign x_7188 = x_528 & x_529;
assign x_7189 = x_527 & x_7188;
assign x_7190 = x_530 & x_531;
assign x_7191 = x_532 & x_533;
assign x_7192 = x_7190 & x_7191;
assign x_7193 = x_7189 & x_7192;
assign x_7194 = x_7187 & x_7193;
assign x_7195 = x_535 & x_536;
assign x_7196 = x_534 & x_7195;
assign x_7197 = x_538 & x_539;
assign x_7198 = x_537 & x_7197;
assign x_7199 = x_7196 & x_7198;
assign x_7200 = x_541 & x_542;
assign x_7201 = x_540 & x_7200;
assign x_7202 = x_543 & x_544;
assign x_7203 = x_545 & x_546;
assign x_7204 = x_7202 & x_7203;
assign x_7205 = x_7201 & x_7204;
assign x_7206 = x_7199 & x_7205;
assign x_7207 = x_7194 & x_7206;
assign x_7208 = x_548 & x_549;
assign x_7209 = x_547 & x_7208;
assign x_7210 = x_551 & x_552;
assign x_7211 = x_550 & x_7210;
assign x_7212 = x_7209 & x_7211;
assign x_7213 = x_554 & x_555;
assign x_7214 = x_553 & x_7213;
assign x_7215 = x_556 & x_557;
assign x_7216 = x_558 & x_559;
assign x_7217 = x_7215 & x_7216;
assign x_7218 = x_7214 & x_7217;
assign x_7219 = x_7212 & x_7218;
assign x_7220 = x_561 & x_562;
assign x_7221 = x_560 & x_7220;
assign x_7222 = x_564 & x_565;
assign x_7223 = x_563 & x_7222;
assign x_7224 = x_7221 & x_7223;
assign x_7225 = x_567 & x_568;
assign x_7226 = x_566 & x_7225;
assign x_7227 = x_569 & x_570;
assign x_7228 = x_571 & x_572;
assign x_7229 = x_7227 & x_7228;
assign x_7230 = x_7226 & x_7229;
assign x_7231 = x_7224 & x_7230;
assign x_7232 = x_7219 & x_7231;
assign x_7233 = x_7207 & x_7232;
assign x_7234 = x_574 & x_575;
assign x_7235 = x_573 & x_7234;
assign x_7236 = x_577 & x_578;
assign x_7237 = x_576 & x_7236;
assign x_7238 = x_7235 & x_7237;
assign x_7239 = x_580 & x_581;
assign x_7240 = x_579 & x_7239;
assign x_7241 = x_582 & x_583;
assign x_7242 = x_584 & x_585;
assign x_7243 = x_7241 & x_7242;
assign x_7244 = x_7240 & x_7243;
assign x_7245 = x_7238 & x_7244;
assign x_7246 = x_587 & x_588;
assign x_7247 = x_586 & x_7246;
assign x_7248 = x_590 & x_591;
assign x_7249 = x_589 & x_7248;
assign x_7250 = x_7247 & x_7249;
assign x_7251 = x_593 & x_594;
assign x_7252 = x_592 & x_7251;
assign x_7253 = x_595 & x_596;
assign x_7254 = x_597 & x_598;
assign x_7255 = x_7253 & x_7254;
assign x_7256 = x_7252 & x_7255;
assign x_7257 = x_7250 & x_7256;
assign x_7258 = x_7245 & x_7257;
assign x_7259 = x_600 & x_601;
assign x_7260 = x_599 & x_7259;
assign x_7261 = x_603 & x_604;
assign x_7262 = x_602 & x_7261;
assign x_7263 = x_7260 & x_7262;
assign x_7264 = x_606 & x_607;
assign x_7265 = x_605 & x_7264;
assign x_7266 = x_608 & x_609;
assign x_7267 = x_610 & x_611;
assign x_7268 = x_7266 & x_7267;
assign x_7269 = x_7265 & x_7268;
assign x_7270 = x_7263 & x_7269;
assign x_7271 = x_613 & x_614;
assign x_7272 = x_612 & x_7271;
assign x_7273 = x_616 & x_617;
assign x_7274 = x_615 & x_7273;
assign x_7275 = x_7272 & x_7274;
assign x_7276 = x_619 & x_620;
assign x_7277 = x_618 & x_7276;
assign x_7278 = x_621 & x_622;
assign x_7279 = x_623 & x_624;
assign x_7280 = x_7278 & x_7279;
assign x_7281 = x_7277 & x_7280;
assign x_7282 = x_7275 & x_7281;
assign x_7283 = x_7270 & x_7282;
assign x_7284 = x_7258 & x_7283;
assign x_7285 = x_7233 & x_7284;
assign x_7286 = x_7182 & x_7285;
assign x_7287 = x_626 & x_627;
assign x_7288 = x_625 & x_7287;
assign x_7289 = x_629 & x_630;
assign x_7290 = x_628 & x_7289;
assign x_7291 = x_7288 & x_7290;
assign x_7292 = x_632 & x_633;
assign x_7293 = x_631 & x_7292;
assign x_7294 = x_634 & x_635;
assign x_7295 = x_636 & x_637;
assign x_7296 = x_7294 & x_7295;
assign x_7297 = x_7293 & x_7296;
assign x_7298 = x_7291 & x_7297;
assign x_7299 = x_639 & x_640;
assign x_7300 = x_638 & x_7299;
assign x_7301 = x_642 & x_643;
assign x_7302 = x_641 & x_7301;
assign x_7303 = x_7300 & x_7302;
assign x_7304 = x_645 & x_646;
assign x_7305 = x_644 & x_7304;
assign x_7306 = x_647 & x_648;
assign x_7307 = x_649 & x_650;
assign x_7308 = x_7306 & x_7307;
assign x_7309 = x_7305 & x_7308;
assign x_7310 = x_7303 & x_7309;
assign x_7311 = x_7298 & x_7310;
assign x_7312 = x_652 & x_653;
assign x_7313 = x_651 & x_7312;
assign x_7314 = x_655 & x_656;
assign x_7315 = x_654 & x_7314;
assign x_7316 = x_7313 & x_7315;
assign x_7317 = x_658 & x_659;
assign x_7318 = x_657 & x_7317;
assign x_7319 = x_660 & x_661;
assign x_7320 = x_662 & x_663;
assign x_7321 = x_7319 & x_7320;
assign x_7322 = x_7318 & x_7321;
assign x_7323 = x_7316 & x_7322;
assign x_7324 = x_665 & x_666;
assign x_7325 = x_664 & x_7324;
assign x_7326 = x_668 & x_669;
assign x_7327 = x_667 & x_7326;
assign x_7328 = x_7325 & x_7327;
assign x_7329 = x_671 & x_672;
assign x_7330 = x_670 & x_7329;
assign x_7331 = x_673 & x_674;
assign x_7332 = x_675 & x_676;
assign x_7333 = x_7331 & x_7332;
assign x_7334 = x_7330 & x_7333;
assign x_7335 = x_7328 & x_7334;
assign x_7336 = x_7323 & x_7335;
assign x_7337 = x_7311 & x_7336;
assign x_7338 = x_678 & x_679;
assign x_7339 = x_677 & x_7338;
assign x_7340 = x_681 & x_682;
assign x_7341 = x_680 & x_7340;
assign x_7342 = x_7339 & x_7341;
assign x_7343 = x_684 & x_685;
assign x_7344 = x_683 & x_7343;
assign x_7345 = x_686 & x_687;
assign x_7346 = x_688 & x_689;
assign x_7347 = x_7345 & x_7346;
assign x_7348 = x_7344 & x_7347;
assign x_7349 = x_7342 & x_7348;
assign x_7350 = x_691 & x_692;
assign x_7351 = x_690 & x_7350;
assign x_7352 = x_694 & x_695;
assign x_7353 = x_693 & x_7352;
assign x_7354 = x_7351 & x_7353;
assign x_7355 = x_697 & x_698;
assign x_7356 = x_696 & x_7355;
assign x_7357 = x_699 & x_700;
assign x_7358 = x_701 & x_702;
assign x_7359 = x_7357 & x_7358;
assign x_7360 = x_7356 & x_7359;
assign x_7361 = x_7354 & x_7360;
assign x_7362 = x_7349 & x_7361;
assign x_7363 = x_704 & x_705;
assign x_7364 = x_703 & x_7363;
assign x_7365 = x_707 & x_708;
assign x_7366 = x_706 & x_7365;
assign x_7367 = x_7364 & x_7366;
assign x_7368 = x_710 & x_711;
assign x_7369 = x_709 & x_7368;
assign x_7370 = x_712 & x_713;
assign x_7371 = x_714 & x_715;
assign x_7372 = x_7370 & x_7371;
assign x_7373 = x_7369 & x_7372;
assign x_7374 = x_7367 & x_7373;
assign x_7375 = x_717 & x_718;
assign x_7376 = x_716 & x_7375;
assign x_7377 = x_720 & x_721;
assign x_7378 = x_719 & x_7377;
assign x_7379 = x_7376 & x_7378;
assign x_7380 = x_723 & x_724;
assign x_7381 = x_722 & x_7380;
assign x_7382 = x_725 & x_726;
assign x_7383 = x_727 & x_728;
assign x_7384 = x_7382 & x_7383;
assign x_7385 = x_7381 & x_7384;
assign x_7386 = x_7379 & x_7385;
assign x_7387 = x_7374 & x_7386;
assign x_7388 = x_7362 & x_7387;
assign x_7389 = x_7337 & x_7388;
assign x_7390 = x_730 & x_731;
assign x_7391 = x_729 & x_7390;
assign x_7392 = x_733 & x_734;
assign x_7393 = x_732 & x_7392;
assign x_7394 = x_7391 & x_7393;
assign x_7395 = x_736 & x_737;
assign x_7396 = x_735 & x_7395;
assign x_7397 = x_738 & x_739;
assign x_7398 = x_740 & x_741;
assign x_7399 = x_7397 & x_7398;
assign x_7400 = x_7396 & x_7399;
assign x_7401 = x_7394 & x_7400;
assign x_7402 = x_743 & x_744;
assign x_7403 = x_742 & x_7402;
assign x_7404 = x_746 & x_747;
assign x_7405 = x_745 & x_7404;
assign x_7406 = x_7403 & x_7405;
assign x_7407 = x_749 & x_750;
assign x_7408 = x_748 & x_7407;
assign x_7409 = x_751 & x_752;
assign x_7410 = x_753 & x_754;
assign x_7411 = x_7409 & x_7410;
assign x_7412 = x_7408 & x_7411;
assign x_7413 = x_7406 & x_7412;
assign x_7414 = x_7401 & x_7413;
assign x_7415 = x_756 & x_757;
assign x_7416 = x_755 & x_7415;
assign x_7417 = x_759 & x_760;
assign x_7418 = x_758 & x_7417;
assign x_7419 = x_7416 & x_7418;
assign x_7420 = x_762 & x_763;
assign x_7421 = x_761 & x_7420;
assign x_7422 = x_764 & x_765;
assign x_7423 = x_766 & x_767;
assign x_7424 = x_7422 & x_7423;
assign x_7425 = x_7421 & x_7424;
assign x_7426 = x_7419 & x_7425;
assign x_7427 = x_769 & x_770;
assign x_7428 = x_768 & x_7427;
assign x_7429 = x_772 & x_773;
assign x_7430 = x_771 & x_7429;
assign x_7431 = x_7428 & x_7430;
assign x_7432 = x_775 & x_776;
assign x_7433 = x_774 & x_7432;
assign x_7434 = x_777 & x_778;
assign x_7435 = x_779 & x_780;
assign x_7436 = x_7434 & x_7435;
assign x_7437 = x_7433 & x_7436;
assign x_7438 = x_7431 & x_7437;
assign x_7439 = x_7426 & x_7438;
assign x_7440 = x_7414 & x_7439;
assign x_7441 = x_782 & x_783;
assign x_7442 = x_781 & x_7441;
assign x_7443 = x_785 & x_786;
assign x_7444 = x_784 & x_7443;
assign x_7445 = x_7442 & x_7444;
assign x_7446 = x_788 & x_789;
assign x_7447 = x_787 & x_7446;
assign x_7448 = x_790 & x_791;
assign x_7449 = x_792 & x_793;
assign x_7450 = x_7448 & x_7449;
assign x_7451 = x_7447 & x_7450;
assign x_7452 = x_7445 & x_7451;
assign x_7453 = x_795 & x_796;
assign x_7454 = x_794 & x_7453;
assign x_7455 = x_798 & x_799;
assign x_7456 = x_797 & x_7455;
assign x_7457 = x_7454 & x_7456;
assign x_7458 = x_801 & x_802;
assign x_7459 = x_800 & x_7458;
assign x_7460 = x_803 & x_804;
assign x_7461 = x_805 & x_806;
assign x_7462 = x_7460 & x_7461;
assign x_7463 = x_7459 & x_7462;
assign x_7464 = x_7457 & x_7463;
assign x_7465 = x_7452 & x_7464;
assign x_7466 = x_808 & x_809;
assign x_7467 = x_807 & x_7466;
assign x_7468 = x_811 & x_812;
assign x_7469 = x_810 & x_7468;
assign x_7470 = x_7467 & x_7469;
assign x_7471 = x_814 & x_815;
assign x_7472 = x_813 & x_7471;
assign x_7473 = x_816 & x_817;
assign x_7474 = x_818 & x_819;
assign x_7475 = x_7473 & x_7474;
assign x_7476 = x_7472 & x_7475;
assign x_7477 = x_7470 & x_7476;
assign x_7478 = x_821 & x_822;
assign x_7479 = x_820 & x_7478;
assign x_7480 = x_823 & x_824;
assign x_7481 = x_825 & x_826;
assign x_7482 = x_7480 & x_7481;
assign x_7483 = x_7479 & x_7482;
assign x_7484 = x_828 & x_829;
assign x_7485 = x_827 & x_7484;
assign x_7486 = x_830 & x_831;
assign x_7487 = x_832 & x_833;
assign x_7488 = x_7486 & x_7487;
assign x_7489 = x_7485 & x_7488;
assign x_7490 = x_7483 & x_7489;
assign x_7491 = x_7477 & x_7490;
assign x_7492 = x_7465 & x_7491;
assign x_7493 = x_7440 & x_7492;
assign x_7494 = x_7389 & x_7493;
assign x_7495 = x_7286 & x_7494;
assign x_7496 = x_7079 & x_7495;
assign x_7497 = x_835 & x_836;
assign x_7498 = x_834 & x_7497;
assign x_7499 = x_838 & x_839;
assign x_7500 = x_837 & x_7499;
assign x_7501 = x_7498 & x_7500;
assign x_7502 = x_841 & x_842;
assign x_7503 = x_840 & x_7502;
assign x_7504 = x_843 & x_844;
assign x_7505 = x_845 & x_846;
assign x_7506 = x_7504 & x_7505;
assign x_7507 = x_7503 & x_7506;
assign x_7508 = x_7501 & x_7507;
assign x_7509 = x_848 & x_849;
assign x_7510 = x_847 & x_7509;
assign x_7511 = x_851 & x_852;
assign x_7512 = x_850 & x_7511;
assign x_7513 = x_7510 & x_7512;
assign x_7514 = x_854 & x_855;
assign x_7515 = x_853 & x_7514;
assign x_7516 = x_856 & x_857;
assign x_7517 = x_858 & x_859;
assign x_7518 = x_7516 & x_7517;
assign x_7519 = x_7515 & x_7518;
assign x_7520 = x_7513 & x_7519;
assign x_7521 = x_7508 & x_7520;
assign x_7522 = x_861 & x_862;
assign x_7523 = x_860 & x_7522;
assign x_7524 = x_864 & x_865;
assign x_7525 = x_863 & x_7524;
assign x_7526 = x_7523 & x_7525;
assign x_7527 = x_867 & x_868;
assign x_7528 = x_866 & x_7527;
assign x_7529 = x_869 & x_870;
assign x_7530 = x_871 & x_872;
assign x_7531 = x_7529 & x_7530;
assign x_7532 = x_7528 & x_7531;
assign x_7533 = x_7526 & x_7532;
assign x_7534 = x_874 & x_875;
assign x_7535 = x_873 & x_7534;
assign x_7536 = x_877 & x_878;
assign x_7537 = x_876 & x_7536;
assign x_7538 = x_7535 & x_7537;
assign x_7539 = x_880 & x_881;
assign x_7540 = x_879 & x_7539;
assign x_7541 = x_882 & x_883;
assign x_7542 = x_884 & x_885;
assign x_7543 = x_7541 & x_7542;
assign x_7544 = x_7540 & x_7543;
assign x_7545 = x_7538 & x_7544;
assign x_7546 = x_7533 & x_7545;
assign x_7547 = x_7521 & x_7546;
assign x_7548 = x_887 & x_888;
assign x_7549 = x_886 & x_7548;
assign x_7550 = x_890 & x_891;
assign x_7551 = x_889 & x_7550;
assign x_7552 = x_7549 & x_7551;
assign x_7553 = x_893 & x_894;
assign x_7554 = x_892 & x_7553;
assign x_7555 = x_895 & x_896;
assign x_7556 = x_897 & x_898;
assign x_7557 = x_7555 & x_7556;
assign x_7558 = x_7554 & x_7557;
assign x_7559 = x_7552 & x_7558;
assign x_7560 = x_900 & x_901;
assign x_7561 = x_899 & x_7560;
assign x_7562 = x_903 & x_904;
assign x_7563 = x_902 & x_7562;
assign x_7564 = x_7561 & x_7563;
assign x_7565 = x_906 & x_907;
assign x_7566 = x_905 & x_7565;
assign x_7567 = x_908 & x_909;
assign x_7568 = x_910 & x_911;
assign x_7569 = x_7567 & x_7568;
assign x_7570 = x_7566 & x_7569;
assign x_7571 = x_7564 & x_7570;
assign x_7572 = x_7559 & x_7571;
assign x_7573 = x_913 & x_914;
assign x_7574 = x_912 & x_7573;
assign x_7575 = x_916 & x_917;
assign x_7576 = x_915 & x_7575;
assign x_7577 = x_7574 & x_7576;
assign x_7578 = x_919 & x_920;
assign x_7579 = x_918 & x_7578;
assign x_7580 = x_921 & x_922;
assign x_7581 = x_923 & x_924;
assign x_7582 = x_7580 & x_7581;
assign x_7583 = x_7579 & x_7582;
assign x_7584 = x_7577 & x_7583;
assign x_7585 = x_926 & x_927;
assign x_7586 = x_925 & x_7585;
assign x_7587 = x_929 & x_930;
assign x_7588 = x_928 & x_7587;
assign x_7589 = x_7586 & x_7588;
assign x_7590 = x_932 & x_933;
assign x_7591 = x_931 & x_7590;
assign x_7592 = x_934 & x_935;
assign x_7593 = x_936 & x_937;
assign x_7594 = x_7592 & x_7593;
assign x_7595 = x_7591 & x_7594;
assign x_7596 = x_7589 & x_7595;
assign x_7597 = x_7584 & x_7596;
assign x_7598 = x_7572 & x_7597;
assign x_7599 = x_7547 & x_7598;
assign x_7600 = x_939 & x_940;
assign x_7601 = x_938 & x_7600;
assign x_7602 = x_942 & x_943;
assign x_7603 = x_941 & x_7602;
assign x_7604 = x_7601 & x_7603;
assign x_7605 = x_945 & x_946;
assign x_7606 = x_944 & x_7605;
assign x_7607 = x_947 & x_948;
assign x_7608 = x_949 & x_950;
assign x_7609 = x_7607 & x_7608;
assign x_7610 = x_7606 & x_7609;
assign x_7611 = x_7604 & x_7610;
assign x_7612 = x_952 & x_953;
assign x_7613 = x_951 & x_7612;
assign x_7614 = x_955 & x_956;
assign x_7615 = x_954 & x_7614;
assign x_7616 = x_7613 & x_7615;
assign x_7617 = x_958 & x_959;
assign x_7618 = x_957 & x_7617;
assign x_7619 = x_960 & x_961;
assign x_7620 = x_962 & x_963;
assign x_7621 = x_7619 & x_7620;
assign x_7622 = x_7618 & x_7621;
assign x_7623 = x_7616 & x_7622;
assign x_7624 = x_7611 & x_7623;
assign x_7625 = x_965 & x_966;
assign x_7626 = x_964 & x_7625;
assign x_7627 = x_968 & x_969;
assign x_7628 = x_967 & x_7627;
assign x_7629 = x_7626 & x_7628;
assign x_7630 = x_971 & x_972;
assign x_7631 = x_970 & x_7630;
assign x_7632 = x_973 & x_974;
assign x_7633 = x_975 & x_976;
assign x_7634 = x_7632 & x_7633;
assign x_7635 = x_7631 & x_7634;
assign x_7636 = x_7629 & x_7635;
assign x_7637 = x_978 & x_979;
assign x_7638 = x_977 & x_7637;
assign x_7639 = x_981 & x_982;
assign x_7640 = x_980 & x_7639;
assign x_7641 = x_7638 & x_7640;
assign x_7642 = x_984 & x_985;
assign x_7643 = x_983 & x_7642;
assign x_7644 = x_986 & x_987;
assign x_7645 = x_988 & x_989;
assign x_7646 = x_7644 & x_7645;
assign x_7647 = x_7643 & x_7646;
assign x_7648 = x_7641 & x_7647;
assign x_7649 = x_7636 & x_7648;
assign x_7650 = x_7624 & x_7649;
assign x_7651 = x_991 & x_992;
assign x_7652 = x_990 & x_7651;
assign x_7653 = x_994 & x_995;
assign x_7654 = x_993 & x_7653;
assign x_7655 = x_7652 & x_7654;
assign x_7656 = x_997 & x_998;
assign x_7657 = x_996 & x_7656;
assign x_7658 = x_999 & x_1000;
assign x_7659 = x_1001 & x_1002;
assign x_7660 = x_7658 & x_7659;
assign x_7661 = x_7657 & x_7660;
assign x_7662 = x_7655 & x_7661;
assign x_7663 = x_1004 & x_1005;
assign x_7664 = x_1003 & x_7663;
assign x_7665 = x_1007 & x_1008;
assign x_7666 = x_1006 & x_7665;
assign x_7667 = x_7664 & x_7666;
assign x_7668 = x_1010 & x_1011;
assign x_7669 = x_1009 & x_7668;
assign x_7670 = x_1012 & x_1013;
assign x_7671 = x_1014 & x_1015;
assign x_7672 = x_7670 & x_7671;
assign x_7673 = x_7669 & x_7672;
assign x_7674 = x_7667 & x_7673;
assign x_7675 = x_7662 & x_7674;
assign x_7676 = x_1017 & x_1018;
assign x_7677 = x_1016 & x_7676;
assign x_7678 = x_1020 & x_1021;
assign x_7679 = x_1019 & x_7678;
assign x_7680 = x_7677 & x_7679;
assign x_7681 = x_1023 & x_1024;
assign x_7682 = x_1022 & x_7681;
assign x_7683 = x_1025 & x_1026;
assign x_7684 = x_1027 & x_1028;
assign x_7685 = x_7683 & x_7684;
assign x_7686 = x_7682 & x_7685;
assign x_7687 = x_7680 & x_7686;
assign x_7688 = x_1030 & x_1031;
assign x_7689 = x_1029 & x_7688;
assign x_7690 = x_1033 & x_1034;
assign x_7691 = x_1032 & x_7690;
assign x_7692 = x_7689 & x_7691;
assign x_7693 = x_1036 & x_1037;
assign x_7694 = x_1035 & x_7693;
assign x_7695 = x_1038 & x_1039;
assign x_7696 = x_1040 & x_1041;
assign x_7697 = x_7695 & x_7696;
assign x_7698 = x_7694 & x_7697;
assign x_7699 = x_7692 & x_7698;
assign x_7700 = x_7687 & x_7699;
assign x_7701 = x_7675 & x_7700;
assign x_7702 = x_7650 & x_7701;
assign x_7703 = x_7599 & x_7702;
assign x_7704 = x_1043 & x_1044;
assign x_7705 = x_1042 & x_7704;
assign x_7706 = x_1046 & x_1047;
assign x_7707 = x_1045 & x_7706;
assign x_7708 = x_7705 & x_7707;
assign x_7709 = x_1049 & x_1050;
assign x_7710 = x_1048 & x_7709;
assign x_7711 = x_1051 & x_1052;
assign x_7712 = x_1053 & x_1054;
assign x_7713 = x_7711 & x_7712;
assign x_7714 = x_7710 & x_7713;
assign x_7715 = x_7708 & x_7714;
assign x_7716 = x_1056 & x_1057;
assign x_7717 = x_1055 & x_7716;
assign x_7718 = x_1059 & x_1060;
assign x_7719 = x_1058 & x_7718;
assign x_7720 = x_7717 & x_7719;
assign x_7721 = x_1062 & x_1063;
assign x_7722 = x_1061 & x_7721;
assign x_7723 = x_1064 & x_1065;
assign x_7724 = x_1066 & x_1067;
assign x_7725 = x_7723 & x_7724;
assign x_7726 = x_7722 & x_7725;
assign x_7727 = x_7720 & x_7726;
assign x_7728 = x_7715 & x_7727;
assign x_7729 = x_1069 & x_1070;
assign x_7730 = x_1068 & x_7729;
assign x_7731 = x_1072 & x_1073;
assign x_7732 = x_1071 & x_7731;
assign x_7733 = x_7730 & x_7732;
assign x_7734 = x_1075 & x_1076;
assign x_7735 = x_1074 & x_7734;
assign x_7736 = x_1077 & x_1078;
assign x_7737 = x_1079 & x_1080;
assign x_7738 = x_7736 & x_7737;
assign x_7739 = x_7735 & x_7738;
assign x_7740 = x_7733 & x_7739;
assign x_7741 = x_1082 & x_1083;
assign x_7742 = x_1081 & x_7741;
assign x_7743 = x_1085 & x_1086;
assign x_7744 = x_1084 & x_7743;
assign x_7745 = x_7742 & x_7744;
assign x_7746 = x_1088 & x_1089;
assign x_7747 = x_1087 & x_7746;
assign x_7748 = x_1090 & x_1091;
assign x_7749 = x_1092 & x_1093;
assign x_7750 = x_7748 & x_7749;
assign x_7751 = x_7747 & x_7750;
assign x_7752 = x_7745 & x_7751;
assign x_7753 = x_7740 & x_7752;
assign x_7754 = x_7728 & x_7753;
assign x_7755 = x_1095 & x_1096;
assign x_7756 = x_1094 & x_7755;
assign x_7757 = x_1098 & x_1099;
assign x_7758 = x_1097 & x_7757;
assign x_7759 = x_7756 & x_7758;
assign x_7760 = x_1101 & x_1102;
assign x_7761 = x_1100 & x_7760;
assign x_7762 = x_1103 & x_1104;
assign x_7763 = x_1105 & x_1106;
assign x_7764 = x_7762 & x_7763;
assign x_7765 = x_7761 & x_7764;
assign x_7766 = x_7759 & x_7765;
assign x_7767 = x_1108 & x_1109;
assign x_7768 = x_1107 & x_7767;
assign x_7769 = x_1111 & x_1112;
assign x_7770 = x_1110 & x_7769;
assign x_7771 = x_7768 & x_7770;
assign x_7772 = x_1114 & x_1115;
assign x_7773 = x_1113 & x_7772;
assign x_7774 = x_1116 & x_1117;
assign x_7775 = x_1118 & x_1119;
assign x_7776 = x_7774 & x_7775;
assign x_7777 = x_7773 & x_7776;
assign x_7778 = x_7771 & x_7777;
assign x_7779 = x_7766 & x_7778;
assign x_7780 = x_1121 & x_1122;
assign x_7781 = x_1120 & x_7780;
assign x_7782 = x_1124 & x_1125;
assign x_7783 = x_1123 & x_7782;
assign x_7784 = x_7781 & x_7783;
assign x_7785 = x_1127 & x_1128;
assign x_7786 = x_1126 & x_7785;
assign x_7787 = x_1129 & x_1130;
assign x_7788 = x_1131 & x_1132;
assign x_7789 = x_7787 & x_7788;
assign x_7790 = x_7786 & x_7789;
assign x_7791 = x_7784 & x_7790;
assign x_7792 = x_1134 & x_1135;
assign x_7793 = x_1133 & x_7792;
assign x_7794 = x_1137 & x_1138;
assign x_7795 = x_1136 & x_7794;
assign x_7796 = x_7793 & x_7795;
assign x_7797 = x_1140 & x_1141;
assign x_7798 = x_1139 & x_7797;
assign x_7799 = x_1142 & x_1143;
assign x_7800 = x_1144 & x_1145;
assign x_7801 = x_7799 & x_7800;
assign x_7802 = x_7798 & x_7801;
assign x_7803 = x_7796 & x_7802;
assign x_7804 = x_7791 & x_7803;
assign x_7805 = x_7779 & x_7804;
assign x_7806 = x_7754 & x_7805;
assign x_7807 = x_1147 & x_1148;
assign x_7808 = x_1146 & x_7807;
assign x_7809 = x_1150 & x_1151;
assign x_7810 = x_1149 & x_7809;
assign x_7811 = x_7808 & x_7810;
assign x_7812 = x_1153 & x_1154;
assign x_7813 = x_1152 & x_7812;
assign x_7814 = x_1155 & x_1156;
assign x_7815 = x_1157 & x_1158;
assign x_7816 = x_7814 & x_7815;
assign x_7817 = x_7813 & x_7816;
assign x_7818 = x_7811 & x_7817;
assign x_7819 = x_1160 & x_1161;
assign x_7820 = x_1159 & x_7819;
assign x_7821 = x_1163 & x_1164;
assign x_7822 = x_1162 & x_7821;
assign x_7823 = x_7820 & x_7822;
assign x_7824 = x_1166 & x_1167;
assign x_7825 = x_1165 & x_7824;
assign x_7826 = x_1168 & x_1169;
assign x_7827 = x_1170 & x_1171;
assign x_7828 = x_7826 & x_7827;
assign x_7829 = x_7825 & x_7828;
assign x_7830 = x_7823 & x_7829;
assign x_7831 = x_7818 & x_7830;
assign x_7832 = x_1173 & x_1174;
assign x_7833 = x_1172 & x_7832;
assign x_7834 = x_1176 & x_1177;
assign x_7835 = x_1175 & x_7834;
assign x_7836 = x_7833 & x_7835;
assign x_7837 = x_1179 & x_1180;
assign x_7838 = x_1178 & x_7837;
assign x_7839 = x_1181 & x_1182;
assign x_7840 = x_1183 & x_1184;
assign x_7841 = x_7839 & x_7840;
assign x_7842 = x_7838 & x_7841;
assign x_7843 = x_7836 & x_7842;
assign x_7844 = x_1186 & x_1187;
assign x_7845 = x_1185 & x_7844;
assign x_7846 = x_1189 & x_1190;
assign x_7847 = x_1188 & x_7846;
assign x_7848 = x_7845 & x_7847;
assign x_7849 = x_1192 & x_1193;
assign x_7850 = x_1191 & x_7849;
assign x_7851 = x_1194 & x_1195;
assign x_7852 = x_1196 & x_1197;
assign x_7853 = x_7851 & x_7852;
assign x_7854 = x_7850 & x_7853;
assign x_7855 = x_7848 & x_7854;
assign x_7856 = x_7843 & x_7855;
assign x_7857 = x_7831 & x_7856;
assign x_7858 = x_1199 & x_1200;
assign x_7859 = x_1198 & x_7858;
assign x_7860 = x_1202 & x_1203;
assign x_7861 = x_1201 & x_7860;
assign x_7862 = x_7859 & x_7861;
assign x_7863 = x_1205 & x_1206;
assign x_7864 = x_1204 & x_7863;
assign x_7865 = x_1207 & x_1208;
assign x_7866 = x_1209 & x_1210;
assign x_7867 = x_7865 & x_7866;
assign x_7868 = x_7864 & x_7867;
assign x_7869 = x_7862 & x_7868;
assign x_7870 = x_1212 & x_1213;
assign x_7871 = x_1211 & x_7870;
assign x_7872 = x_1215 & x_1216;
assign x_7873 = x_1214 & x_7872;
assign x_7874 = x_7871 & x_7873;
assign x_7875 = x_1218 & x_1219;
assign x_7876 = x_1217 & x_7875;
assign x_7877 = x_1220 & x_1221;
assign x_7878 = x_1222 & x_1223;
assign x_7879 = x_7877 & x_7878;
assign x_7880 = x_7876 & x_7879;
assign x_7881 = x_7874 & x_7880;
assign x_7882 = x_7869 & x_7881;
assign x_7883 = x_1225 & x_1226;
assign x_7884 = x_1224 & x_7883;
assign x_7885 = x_1228 & x_1229;
assign x_7886 = x_1227 & x_7885;
assign x_7887 = x_7884 & x_7886;
assign x_7888 = x_1231 & x_1232;
assign x_7889 = x_1230 & x_7888;
assign x_7890 = x_1233 & x_1234;
assign x_7891 = x_1235 & x_1236;
assign x_7892 = x_7890 & x_7891;
assign x_7893 = x_7889 & x_7892;
assign x_7894 = x_7887 & x_7893;
assign x_7895 = x_1238 & x_1239;
assign x_7896 = x_1237 & x_7895;
assign x_7897 = x_1241 & x_1242;
assign x_7898 = x_1240 & x_7897;
assign x_7899 = x_7896 & x_7898;
assign x_7900 = x_1244 & x_1245;
assign x_7901 = x_1243 & x_7900;
assign x_7902 = x_1246 & x_1247;
assign x_7903 = x_1248 & x_1249;
assign x_7904 = x_7902 & x_7903;
assign x_7905 = x_7901 & x_7904;
assign x_7906 = x_7899 & x_7905;
assign x_7907 = x_7894 & x_7906;
assign x_7908 = x_7882 & x_7907;
assign x_7909 = x_7857 & x_7908;
assign x_7910 = x_7806 & x_7909;
assign x_7911 = x_7703 & x_7910;
assign x_7912 = x_1251 & x_1252;
assign x_7913 = x_1250 & x_7912;
assign x_7914 = x_1254 & x_1255;
assign x_7915 = x_1253 & x_7914;
assign x_7916 = x_7913 & x_7915;
assign x_7917 = x_1257 & x_1258;
assign x_7918 = x_1256 & x_7917;
assign x_7919 = x_1259 & x_1260;
assign x_7920 = x_1261 & x_1262;
assign x_7921 = x_7919 & x_7920;
assign x_7922 = x_7918 & x_7921;
assign x_7923 = x_7916 & x_7922;
assign x_7924 = x_1264 & x_1265;
assign x_7925 = x_1263 & x_7924;
assign x_7926 = x_1267 & x_1268;
assign x_7927 = x_1266 & x_7926;
assign x_7928 = x_7925 & x_7927;
assign x_7929 = x_1270 & x_1271;
assign x_7930 = x_1269 & x_7929;
assign x_7931 = x_1272 & x_1273;
assign x_7932 = x_1274 & x_1275;
assign x_7933 = x_7931 & x_7932;
assign x_7934 = x_7930 & x_7933;
assign x_7935 = x_7928 & x_7934;
assign x_7936 = x_7923 & x_7935;
assign x_7937 = x_1277 & x_1278;
assign x_7938 = x_1276 & x_7937;
assign x_7939 = x_1280 & x_1281;
assign x_7940 = x_1279 & x_7939;
assign x_7941 = x_7938 & x_7940;
assign x_7942 = x_1283 & x_1284;
assign x_7943 = x_1282 & x_7942;
assign x_7944 = x_1285 & x_1286;
assign x_7945 = x_1287 & x_1288;
assign x_7946 = x_7944 & x_7945;
assign x_7947 = x_7943 & x_7946;
assign x_7948 = x_7941 & x_7947;
assign x_7949 = x_1290 & x_1291;
assign x_7950 = x_1289 & x_7949;
assign x_7951 = x_1293 & x_1294;
assign x_7952 = x_1292 & x_7951;
assign x_7953 = x_7950 & x_7952;
assign x_7954 = x_1296 & x_1297;
assign x_7955 = x_1295 & x_7954;
assign x_7956 = x_1298 & x_1299;
assign x_7957 = x_1300 & x_1301;
assign x_7958 = x_7956 & x_7957;
assign x_7959 = x_7955 & x_7958;
assign x_7960 = x_7953 & x_7959;
assign x_7961 = x_7948 & x_7960;
assign x_7962 = x_7936 & x_7961;
assign x_7963 = x_1303 & x_1304;
assign x_7964 = x_1302 & x_7963;
assign x_7965 = x_1306 & x_1307;
assign x_7966 = x_1305 & x_7965;
assign x_7967 = x_7964 & x_7966;
assign x_7968 = x_1309 & x_1310;
assign x_7969 = x_1308 & x_7968;
assign x_7970 = x_1311 & x_1312;
assign x_7971 = x_1313 & x_1314;
assign x_7972 = x_7970 & x_7971;
assign x_7973 = x_7969 & x_7972;
assign x_7974 = x_7967 & x_7973;
assign x_7975 = x_1316 & x_1317;
assign x_7976 = x_1315 & x_7975;
assign x_7977 = x_1319 & x_1320;
assign x_7978 = x_1318 & x_7977;
assign x_7979 = x_7976 & x_7978;
assign x_7980 = x_1322 & x_1323;
assign x_7981 = x_1321 & x_7980;
assign x_7982 = x_1324 & x_1325;
assign x_7983 = x_1326 & x_1327;
assign x_7984 = x_7982 & x_7983;
assign x_7985 = x_7981 & x_7984;
assign x_7986 = x_7979 & x_7985;
assign x_7987 = x_7974 & x_7986;
assign x_7988 = x_1329 & x_1330;
assign x_7989 = x_1328 & x_7988;
assign x_7990 = x_1332 & x_1333;
assign x_7991 = x_1331 & x_7990;
assign x_7992 = x_7989 & x_7991;
assign x_7993 = x_1335 & x_1336;
assign x_7994 = x_1334 & x_7993;
assign x_7995 = x_1337 & x_1338;
assign x_7996 = x_1339 & x_1340;
assign x_7997 = x_7995 & x_7996;
assign x_7998 = x_7994 & x_7997;
assign x_7999 = x_7992 & x_7998;
assign x_8000 = x_1342 & x_1343;
assign x_8001 = x_1341 & x_8000;
assign x_8002 = x_1345 & x_1346;
assign x_8003 = x_1344 & x_8002;
assign x_8004 = x_8001 & x_8003;
assign x_8005 = x_1348 & x_1349;
assign x_8006 = x_1347 & x_8005;
assign x_8007 = x_1350 & x_1351;
assign x_8008 = x_1352 & x_1353;
assign x_8009 = x_8007 & x_8008;
assign x_8010 = x_8006 & x_8009;
assign x_8011 = x_8004 & x_8010;
assign x_8012 = x_7999 & x_8011;
assign x_8013 = x_7987 & x_8012;
assign x_8014 = x_7962 & x_8013;
assign x_8015 = x_1355 & x_1356;
assign x_8016 = x_1354 & x_8015;
assign x_8017 = x_1358 & x_1359;
assign x_8018 = x_1357 & x_8017;
assign x_8019 = x_8016 & x_8018;
assign x_8020 = x_1361 & x_1362;
assign x_8021 = x_1360 & x_8020;
assign x_8022 = x_1363 & x_1364;
assign x_8023 = x_1365 & x_1366;
assign x_8024 = x_8022 & x_8023;
assign x_8025 = x_8021 & x_8024;
assign x_8026 = x_8019 & x_8025;
assign x_8027 = x_1368 & x_1369;
assign x_8028 = x_1367 & x_8027;
assign x_8029 = x_1371 & x_1372;
assign x_8030 = x_1370 & x_8029;
assign x_8031 = x_8028 & x_8030;
assign x_8032 = x_1374 & x_1375;
assign x_8033 = x_1373 & x_8032;
assign x_8034 = x_1376 & x_1377;
assign x_8035 = x_1378 & x_1379;
assign x_8036 = x_8034 & x_8035;
assign x_8037 = x_8033 & x_8036;
assign x_8038 = x_8031 & x_8037;
assign x_8039 = x_8026 & x_8038;
assign x_8040 = x_1381 & x_1382;
assign x_8041 = x_1380 & x_8040;
assign x_8042 = x_1384 & x_1385;
assign x_8043 = x_1383 & x_8042;
assign x_8044 = x_8041 & x_8043;
assign x_8045 = x_1387 & x_1388;
assign x_8046 = x_1386 & x_8045;
assign x_8047 = x_1389 & x_1390;
assign x_8048 = x_1391 & x_1392;
assign x_8049 = x_8047 & x_8048;
assign x_8050 = x_8046 & x_8049;
assign x_8051 = x_8044 & x_8050;
assign x_8052 = x_1394 & x_1395;
assign x_8053 = x_1393 & x_8052;
assign x_8054 = x_1397 & x_1398;
assign x_8055 = x_1396 & x_8054;
assign x_8056 = x_8053 & x_8055;
assign x_8057 = x_1400 & x_1401;
assign x_8058 = x_1399 & x_8057;
assign x_8059 = x_1402 & x_1403;
assign x_8060 = x_1404 & x_1405;
assign x_8061 = x_8059 & x_8060;
assign x_8062 = x_8058 & x_8061;
assign x_8063 = x_8056 & x_8062;
assign x_8064 = x_8051 & x_8063;
assign x_8065 = x_8039 & x_8064;
assign x_8066 = x_1407 & x_1408;
assign x_8067 = x_1406 & x_8066;
assign x_8068 = x_1410 & x_1411;
assign x_8069 = x_1409 & x_8068;
assign x_8070 = x_8067 & x_8069;
assign x_8071 = x_1413 & x_1414;
assign x_8072 = x_1412 & x_8071;
assign x_8073 = x_1415 & x_1416;
assign x_8074 = x_1417 & x_1418;
assign x_8075 = x_8073 & x_8074;
assign x_8076 = x_8072 & x_8075;
assign x_8077 = x_8070 & x_8076;
assign x_8078 = x_1420 & x_1421;
assign x_8079 = x_1419 & x_8078;
assign x_8080 = x_1423 & x_1424;
assign x_8081 = x_1422 & x_8080;
assign x_8082 = x_8079 & x_8081;
assign x_8083 = x_1426 & x_1427;
assign x_8084 = x_1425 & x_8083;
assign x_8085 = x_1428 & x_1429;
assign x_8086 = x_1430 & x_1431;
assign x_8087 = x_8085 & x_8086;
assign x_8088 = x_8084 & x_8087;
assign x_8089 = x_8082 & x_8088;
assign x_8090 = x_8077 & x_8089;
assign x_8091 = x_1433 & x_1434;
assign x_8092 = x_1432 & x_8091;
assign x_8093 = x_1436 & x_1437;
assign x_8094 = x_1435 & x_8093;
assign x_8095 = x_8092 & x_8094;
assign x_8096 = x_1439 & x_1440;
assign x_8097 = x_1438 & x_8096;
assign x_8098 = x_1441 & x_1442;
assign x_8099 = x_1443 & x_1444;
assign x_8100 = x_8098 & x_8099;
assign x_8101 = x_8097 & x_8100;
assign x_8102 = x_8095 & x_8101;
assign x_8103 = x_1446 & x_1447;
assign x_8104 = x_1445 & x_8103;
assign x_8105 = x_1449 & x_1450;
assign x_8106 = x_1448 & x_8105;
assign x_8107 = x_8104 & x_8106;
assign x_8108 = x_1452 & x_1453;
assign x_8109 = x_1451 & x_8108;
assign x_8110 = x_1454 & x_1455;
assign x_8111 = x_1456 & x_1457;
assign x_8112 = x_8110 & x_8111;
assign x_8113 = x_8109 & x_8112;
assign x_8114 = x_8107 & x_8113;
assign x_8115 = x_8102 & x_8114;
assign x_8116 = x_8090 & x_8115;
assign x_8117 = x_8065 & x_8116;
assign x_8118 = x_8014 & x_8117;
assign x_8119 = x_1459 & x_1460;
assign x_8120 = x_1458 & x_8119;
assign x_8121 = x_1462 & x_1463;
assign x_8122 = x_1461 & x_8121;
assign x_8123 = x_8120 & x_8122;
assign x_8124 = x_1465 & x_1466;
assign x_8125 = x_1464 & x_8124;
assign x_8126 = x_1467 & x_1468;
assign x_8127 = x_1469 & x_1470;
assign x_8128 = x_8126 & x_8127;
assign x_8129 = x_8125 & x_8128;
assign x_8130 = x_8123 & x_8129;
assign x_8131 = x_1472 & x_1473;
assign x_8132 = x_1471 & x_8131;
assign x_8133 = x_1475 & x_1476;
assign x_8134 = x_1474 & x_8133;
assign x_8135 = x_8132 & x_8134;
assign x_8136 = x_1478 & x_1479;
assign x_8137 = x_1477 & x_8136;
assign x_8138 = x_1480 & x_1481;
assign x_8139 = x_1482 & x_1483;
assign x_8140 = x_8138 & x_8139;
assign x_8141 = x_8137 & x_8140;
assign x_8142 = x_8135 & x_8141;
assign x_8143 = x_8130 & x_8142;
assign x_8144 = x_1485 & x_1486;
assign x_8145 = x_1484 & x_8144;
assign x_8146 = x_1488 & x_1489;
assign x_8147 = x_1487 & x_8146;
assign x_8148 = x_8145 & x_8147;
assign x_8149 = x_1491 & x_1492;
assign x_8150 = x_1490 & x_8149;
assign x_8151 = x_1493 & x_1494;
assign x_8152 = x_1495 & x_1496;
assign x_8153 = x_8151 & x_8152;
assign x_8154 = x_8150 & x_8153;
assign x_8155 = x_8148 & x_8154;
assign x_8156 = x_1498 & x_1499;
assign x_8157 = x_1497 & x_8156;
assign x_8158 = x_1501 & x_1502;
assign x_8159 = x_1500 & x_8158;
assign x_8160 = x_8157 & x_8159;
assign x_8161 = x_1504 & x_1505;
assign x_8162 = x_1503 & x_8161;
assign x_8163 = x_1506 & x_1507;
assign x_8164 = x_1508 & x_1509;
assign x_8165 = x_8163 & x_8164;
assign x_8166 = x_8162 & x_8165;
assign x_8167 = x_8160 & x_8166;
assign x_8168 = x_8155 & x_8167;
assign x_8169 = x_8143 & x_8168;
assign x_8170 = x_1511 & x_1512;
assign x_8171 = x_1510 & x_8170;
assign x_8172 = x_1514 & x_1515;
assign x_8173 = x_1513 & x_8172;
assign x_8174 = x_8171 & x_8173;
assign x_8175 = x_1517 & x_1518;
assign x_8176 = x_1516 & x_8175;
assign x_8177 = x_1519 & x_1520;
assign x_8178 = x_1521 & x_1522;
assign x_8179 = x_8177 & x_8178;
assign x_8180 = x_8176 & x_8179;
assign x_8181 = x_8174 & x_8180;
assign x_8182 = x_1524 & x_1525;
assign x_8183 = x_1523 & x_8182;
assign x_8184 = x_1527 & x_1528;
assign x_8185 = x_1526 & x_8184;
assign x_8186 = x_8183 & x_8185;
assign x_8187 = x_1530 & x_1531;
assign x_8188 = x_1529 & x_8187;
assign x_8189 = x_1532 & x_1533;
assign x_8190 = x_1534 & x_1535;
assign x_8191 = x_8189 & x_8190;
assign x_8192 = x_8188 & x_8191;
assign x_8193 = x_8186 & x_8192;
assign x_8194 = x_8181 & x_8193;
assign x_8195 = x_1537 & x_1538;
assign x_8196 = x_1536 & x_8195;
assign x_8197 = x_1540 & x_1541;
assign x_8198 = x_1539 & x_8197;
assign x_8199 = x_8196 & x_8198;
assign x_8200 = x_1543 & x_1544;
assign x_8201 = x_1542 & x_8200;
assign x_8202 = x_1545 & x_1546;
assign x_8203 = x_1547 & x_1548;
assign x_8204 = x_8202 & x_8203;
assign x_8205 = x_8201 & x_8204;
assign x_8206 = x_8199 & x_8205;
assign x_8207 = x_1550 & x_1551;
assign x_8208 = x_1549 & x_8207;
assign x_8209 = x_1553 & x_1554;
assign x_8210 = x_1552 & x_8209;
assign x_8211 = x_8208 & x_8210;
assign x_8212 = x_1556 & x_1557;
assign x_8213 = x_1555 & x_8212;
assign x_8214 = x_1558 & x_1559;
assign x_8215 = x_1560 & x_1561;
assign x_8216 = x_8214 & x_8215;
assign x_8217 = x_8213 & x_8216;
assign x_8218 = x_8211 & x_8217;
assign x_8219 = x_8206 & x_8218;
assign x_8220 = x_8194 & x_8219;
assign x_8221 = x_8169 & x_8220;
assign x_8222 = x_1563 & x_1564;
assign x_8223 = x_1562 & x_8222;
assign x_8224 = x_1566 & x_1567;
assign x_8225 = x_1565 & x_8224;
assign x_8226 = x_8223 & x_8225;
assign x_8227 = x_1569 & x_1570;
assign x_8228 = x_1568 & x_8227;
assign x_8229 = x_1571 & x_1572;
assign x_8230 = x_1573 & x_1574;
assign x_8231 = x_8229 & x_8230;
assign x_8232 = x_8228 & x_8231;
assign x_8233 = x_8226 & x_8232;
assign x_8234 = x_1576 & x_1577;
assign x_8235 = x_1575 & x_8234;
assign x_8236 = x_1579 & x_1580;
assign x_8237 = x_1578 & x_8236;
assign x_8238 = x_8235 & x_8237;
assign x_8239 = x_1582 & x_1583;
assign x_8240 = x_1581 & x_8239;
assign x_8241 = x_1584 & x_1585;
assign x_8242 = x_1586 & x_1587;
assign x_8243 = x_8241 & x_8242;
assign x_8244 = x_8240 & x_8243;
assign x_8245 = x_8238 & x_8244;
assign x_8246 = x_8233 & x_8245;
assign x_8247 = x_1589 & x_1590;
assign x_8248 = x_1588 & x_8247;
assign x_8249 = x_1592 & x_1593;
assign x_8250 = x_1591 & x_8249;
assign x_8251 = x_8248 & x_8250;
assign x_8252 = x_1595 & x_1596;
assign x_8253 = x_1594 & x_8252;
assign x_8254 = x_1597 & x_1598;
assign x_8255 = x_1599 & x_1600;
assign x_8256 = x_8254 & x_8255;
assign x_8257 = x_8253 & x_8256;
assign x_8258 = x_8251 & x_8257;
assign x_8259 = x_1602 & x_1603;
assign x_8260 = x_1601 & x_8259;
assign x_8261 = x_1605 & x_1606;
assign x_8262 = x_1604 & x_8261;
assign x_8263 = x_8260 & x_8262;
assign x_8264 = x_1608 & x_1609;
assign x_8265 = x_1607 & x_8264;
assign x_8266 = x_1610 & x_1611;
assign x_8267 = x_1612 & x_1613;
assign x_8268 = x_8266 & x_8267;
assign x_8269 = x_8265 & x_8268;
assign x_8270 = x_8263 & x_8269;
assign x_8271 = x_8258 & x_8270;
assign x_8272 = x_8246 & x_8271;
assign x_8273 = x_1615 & x_1616;
assign x_8274 = x_1614 & x_8273;
assign x_8275 = x_1618 & x_1619;
assign x_8276 = x_1617 & x_8275;
assign x_8277 = x_8274 & x_8276;
assign x_8278 = x_1621 & x_1622;
assign x_8279 = x_1620 & x_8278;
assign x_8280 = x_1623 & x_1624;
assign x_8281 = x_1625 & x_1626;
assign x_8282 = x_8280 & x_8281;
assign x_8283 = x_8279 & x_8282;
assign x_8284 = x_8277 & x_8283;
assign x_8285 = x_1628 & x_1629;
assign x_8286 = x_1627 & x_8285;
assign x_8287 = x_1631 & x_1632;
assign x_8288 = x_1630 & x_8287;
assign x_8289 = x_8286 & x_8288;
assign x_8290 = x_1634 & x_1635;
assign x_8291 = x_1633 & x_8290;
assign x_8292 = x_1636 & x_1637;
assign x_8293 = x_1638 & x_1639;
assign x_8294 = x_8292 & x_8293;
assign x_8295 = x_8291 & x_8294;
assign x_8296 = x_8289 & x_8295;
assign x_8297 = x_8284 & x_8296;
assign x_8298 = x_1641 & x_1642;
assign x_8299 = x_1640 & x_8298;
assign x_8300 = x_1644 & x_1645;
assign x_8301 = x_1643 & x_8300;
assign x_8302 = x_8299 & x_8301;
assign x_8303 = x_1647 & x_1648;
assign x_8304 = x_1646 & x_8303;
assign x_8305 = x_1649 & x_1650;
assign x_8306 = x_1651 & x_1652;
assign x_8307 = x_8305 & x_8306;
assign x_8308 = x_8304 & x_8307;
assign x_8309 = x_8302 & x_8308;
assign x_8310 = x_1654 & x_1655;
assign x_8311 = x_1653 & x_8310;
assign x_8312 = x_1656 & x_1657;
assign x_8313 = x_1658 & x_1659;
assign x_8314 = x_8312 & x_8313;
assign x_8315 = x_8311 & x_8314;
assign x_8316 = x_1661 & x_1662;
assign x_8317 = x_1660 & x_8316;
assign x_8318 = x_1663 & x_1664;
assign x_8319 = x_1665 & x_1666;
assign x_8320 = x_8318 & x_8319;
assign x_8321 = x_8317 & x_8320;
assign x_8322 = x_8315 & x_8321;
assign x_8323 = x_8309 & x_8322;
assign x_8324 = x_8297 & x_8323;
assign x_8325 = x_8272 & x_8324;
assign x_8326 = x_8221 & x_8325;
assign x_8327 = x_8118 & x_8326;
assign x_8328 = x_7911 & x_8327;
assign x_8329 = x_7496 & x_8328;
assign x_8330 = x_1668 & x_1669;
assign x_8331 = x_1667 & x_8330;
assign x_8332 = x_1671 & x_1672;
assign x_8333 = x_1670 & x_8332;
assign x_8334 = x_8331 & x_8333;
assign x_8335 = x_1674 & x_1675;
assign x_8336 = x_1673 & x_8335;
assign x_8337 = x_1676 & x_1677;
assign x_8338 = x_1678 & x_1679;
assign x_8339 = x_8337 & x_8338;
assign x_8340 = x_8336 & x_8339;
assign x_8341 = x_8334 & x_8340;
assign x_8342 = x_1681 & x_1682;
assign x_8343 = x_1680 & x_8342;
assign x_8344 = x_1684 & x_1685;
assign x_8345 = x_1683 & x_8344;
assign x_8346 = x_8343 & x_8345;
assign x_8347 = x_1687 & x_1688;
assign x_8348 = x_1686 & x_8347;
assign x_8349 = x_1689 & x_1690;
assign x_8350 = x_1691 & x_1692;
assign x_8351 = x_8349 & x_8350;
assign x_8352 = x_8348 & x_8351;
assign x_8353 = x_8346 & x_8352;
assign x_8354 = x_8341 & x_8353;
assign x_8355 = x_1694 & x_1695;
assign x_8356 = x_1693 & x_8355;
assign x_8357 = x_1697 & x_1698;
assign x_8358 = x_1696 & x_8357;
assign x_8359 = x_8356 & x_8358;
assign x_8360 = x_1700 & x_1701;
assign x_8361 = x_1699 & x_8360;
assign x_8362 = x_1702 & x_1703;
assign x_8363 = x_1704 & x_1705;
assign x_8364 = x_8362 & x_8363;
assign x_8365 = x_8361 & x_8364;
assign x_8366 = x_8359 & x_8365;
assign x_8367 = x_1707 & x_1708;
assign x_8368 = x_1706 & x_8367;
assign x_8369 = x_1710 & x_1711;
assign x_8370 = x_1709 & x_8369;
assign x_8371 = x_8368 & x_8370;
assign x_8372 = x_1713 & x_1714;
assign x_8373 = x_1712 & x_8372;
assign x_8374 = x_1715 & x_1716;
assign x_8375 = x_1717 & x_1718;
assign x_8376 = x_8374 & x_8375;
assign x_8377 = x_8373 & x_8376;
assign x_8378 = x_8371 & x_8377;
assign x_8379 = x_8366 & x_8378;
assign x_8380 = x_8354 & x_8379;
assign x_8381 = x_1720 & x_1721;
assign x_8382 = x_1719 & x_8381;
assign x_8383 = x_1723 & x_1724;
assign x_8384 = x_1722 & x_8383;
assign x_8385 = x_8382 & x_8384;
assign x_8386 = x_1726 & x_1727;
assign x_8387 = x_1725 & x_8386;
assign x_8388 = x_1728 & x_1729;
assign x_8389 = x_1730 & x_1731;
assign x_8390 = x_8388 & x_8389;
assign x_8391 = x_8387 & x_8390;
assign x_8392 = x_8385 & x_8391;
assign x_8393 = x_1733 & x_1734;
assign x_8394 = x_1732 & x_8393;
assign x_8395 = x_1736 & x_1737;
assign x_8396 = x_1735 & x_8395;
assign x_8397 = x_8394 & x_8396;
assign x_8398 = x_1739 & x_1740;
assign x_8399 = x_1738 & x_8398;
assign x_8400 = x_1741 & x_1742;
assign x_8401 = x_1743 & x_1744;
assign x_8402 = x_8400 & x_8401;
assign x_8403 = x_8399 & x_8402;
assign x_8404 = x_8397 & x_8403;
assign x_8405 = x_8392 & x_8404;
assign x_8406 = x_1746 & x_1747;
assign x_8407 = x_1745 & x_8406;
assign x_8408 = x_1749 & x_1750;
assign x_8409 = x_1748 & x_8408;
assign x_8410 = x_8407 & x_8409;
assign x_8411 = x_1752 & x_1753;
assign x_8412 = x_1751 & x_8411;
assign x_8413 = x_1754 & x_1755;
assign x_8414 = x_1756 & x_1757;
assign x_8415 = x_8413 & x_8414;
assign x_8416 = x_8412 & x_8415;
assign x_8417 = x_8410 & x_8416;
assign x_8418 = x_1759 & x_1760;
assign x_8419 = x_1758 & x_8418;
assign x_8420 = x_1762 & x_1763;
assign x_8421 = x_1761 & x_8420;
assign x_8422 = x_8419 & x_8421;
assign x_8423 = x_1765 & x_1766;
assign x_8424 = x_1764 & x_8423;
assign x_8425 = x_1767 & x_1768;
assign x_8426 = x_1769 & x_1770;
assign x_8427 = x_8425 & x_8426;
assign x_8428 = x_8424 & x_8427;
assign x_8429 = x_8422 & x_8428;
assign x_8430 = x_8417 & x_8429;
assign x_8431 = x_8405 & x_8430;
assign x_8432 = x_8380 & x_8431;
assign x_8433 = x_1772 & x_1773;
assign x_8434 = x_1771 & x_8433;
assign x_8435 = x_1775 & x_1776;
assign x_8436 = x_1774 & x_8435;
assign x_8437 = x_8434 & x_8436;
assign x_8438 = x_1778 & x_1779;
assign x_8439 = x_1777 & x_8438;
assign x_8440 = x_1780 & x_1781;
assign x_8441 = x_1782 & x_1783;
assign x_8442 = x_8440 & x_8441;
assign x_8443 = x_8439 & x_8442;
assign x_8444 = x_8437 & x_8443;
assign x_8445 = x_1785 & x_1786;
assign x_8446 = x_1784 & x_8445;
assign x_8447 = x_1788 & x_1789;
assign x_8448 = x_1787 & x_8447;
assign x_8449 = x_8446 & x_8448;
assign x_8450 = x_1791 & x_1792;
assign x_8451 = x_1790 & x_8450;
assign x_8452 = x_1793 & x_1794;
assign x_8453 = x_1795 & x_1796;
assign x_8454 = x_8452 & x_8453;
assign x_8455 = x_8451 & x_8454;
assign x_8456 = x_8449 & x_8455;
assign x_8457 = x_8444 & x_8456;
assign x_8458 = x_1798 & x_1799;
assign x_8459 = x_1797 & x_8458;
assign x_8460 = x_1801 & x_1802;
assign x_8461 = x_1800 & x_8460;
assign x_8462 = x_8459 & x_8461;
assign x_8463 = x_1804 & x_1805;
assign x_8464 = x_1803 & x_8463;
assign x_8465 = x_1806 & x_1807;
assign x_8466 = x_1808 & x_1809;
assign x_8467 = x_8465 & x_8466;
assign x_8468 = x_8464 & x_8467;
assign x_8469 = x_8462 & x_8468;
assign x_8470 = x_1811 & x_1812;
assign x_8471 = x_1810 & x_8470;
assign x_8472 = x_1814 & x_1815;
assign x_8473 = x_1813 & x_8472;
assign x_8474 = x_8471 & x_8473;
assign x_8475 = x_1817 & x_1818;
assign x_8476 = x_1816 & x_8475;
assign x_8477 = x_1819 & x_1820;
assign x_8478 = x_1821 & x_1822;
assign x_8479 = x_8477 & x_8478;
assign x_8480 = x_8476 & x_8479;
assign x_8481 = x_8474 & x_8480;
assign x_8482 = x_8469 & x_8481;
assign x_8483 = x_8457 & x_8482;
assign x_8484 = x_1824 & x_1825;
assign x_8485 = x_1823 & x_8484;
assign x_8486 = x_1827 & x_1828;
assign x_8487 = x_1826 & x_8486;
assign x_8488 = x_8485 & x_8487;
assign x_8489 = x_1830 & x_1831;
assign x_8490 = x_1829 & x_8489;
assign x_8491 = x_1832 & x_1833;
assign x_8492 = x_1834 & x_1835;
assign x_8493 = x_8491 & x_8492;
assign x_8494 = x_8490 & x_8493;
assign x_8495 = x_8488 & x_8494;
assign x_8496 = x_1837 & x_1838;
assign x_8497 = x_1836 & x_8496;
assign x_8498 = x_1840 & x_1841;
assign x_8499 = x_1839 & x_8498;
assign x_8500 = x_8497 & x_8499;
assign x_8501 = x_1843 & x_1844;
assign x_8502 = x_1842 & x_8501;
assign x_8503 = x_1845 & x_1846;
assign x_8504 = x_1847 & x_1848;
assign x_8505 = x_8503 & x_8504;
assign x_8506 = x_8502 & x_8505;
assign x_8507 = x_8500 & x_8506;
assign x_8508 = x_8495 & x_8507;
assign x_8509 = x_1850 & x_1851;
assign x_8510 = x_1849 & x_8509;
assign x_8511 = x_1853 & x_1854;
assign x_8512 = x_1852 & x_8511;
assign x_8513 = x_8510 & x_8512;
assign x_8514 = x_1856 & x_1857;
assign x_8515 = x_1855 & x_8514;
assign x_8516 = x_1858 & x_1859;
assign x_8517 = x_1860 & x_1861;
assign x_8518 = x_8516 & x_8517;
assign x_8519 = x_8515 & x_8518;
assign x_8520 = x_8513 & x_8519;
assign x_8521 = x_1863 & x_1864;
assign x_8522 = x_1862 & x_8521;
assign x_8523 = x_1866 & x_1867;
assign x_8524 = x_1865 & x_8523;
assign x_8525 = x_8522 & x_8524;
assign x_8526 = x_1869 & x_1870;
assign x_8527 = x_1868 & x_8526;
assign x_8528 = x_1871 & x_1872;
assign x_8529 = x_1873 & x_1874;
assign x_8530 = x_8528 & x_8529;
assign x_8531 = x_8527 & x_8530;
assign x_8532 = x_8525 & x_8531;
assign x_8533 = x_8520 & x_8532;
assign x_8534 = x_8508 & x_8533;
assign x_8535 = x_8483 & x_8534;
assign x_8536 = x_8432 & x_8535;
assign x_8537 = x_1876 & x_1877;
assign x_8538 = x_1875 & x_8537;
assign x_8539 = x_1879 & x_1880;
assign x_8540 = x_1878 & x_8539;
assign x_8541 = x_8538 & x_8540;
assign x_8542 = x_1882 & x_1883;
assign x_8543 = x_1881 & x_8542;
assign x_8544 = x_1884 & x_1885;
assign x_8545 = x_1886 & x_1887;
assign x_8546 = x_8544 & x_8545;
assign x_8547 = x_8543 & x_8546;
assign x_8548 = x_8541 & x_8547;
assign x_8549 = x_1889 & x_1890;
assign x_8550 = x_1888 & x_8549;
assign x_8551 = x_1892 & x_1893;
assign x_8552 = x_1891 & x_8551;
assign x_8553 = x_8550 & x_8552;
assign x_8554 = x_1895 & x_1896;
assign x_8555 = x_1894 & x_8554;
assign x_8556 = x_1897 & x_1898;
assign x_8557 = x_1899 & x_1900;
assign x_8558 = x_8556 & x_8557;
assign x_8559 = x_8555 & x_8558;
assign x_8560 = x_8553 & x_8559;
assign x_8561 = x_8548 & x_8560;
assign x_8562 = x_1902 & x_1903;
assign x_8563 = x_1901 & x_8562;
assign x_8564 = x_1905 & x_1906;
assign x_8565 = x_1904 & x_8564;
assign x_8566 = x_8563 & x_8565;
assign x_8567 = x_1908 & x_1909;
assign x_8568 = x_1907 & x_8567;
assign x_8569 = x_1910 & x_1911;
assign x_8570 = x_1912 & x_1913;
assign x_8571 = x_8569 & x_8570;
assign x_8572 = x_8568 & x_8571;
assign x_8573 = x_8566 & x_8572;
assign x_8574 = x_1915 & x_1916;
assign x_8575 = x_1914 & x_8574;
assign x_8576 = x_1918 & x_1919;
assign x_8577 = x_1917 & x_8576;
assign x_8578 = x_8575 & x_8577;
assign x_8579 = x_1921 & x_1922;
assign x_8580 = x_1920 & x_8579;
assign x_8581 = x_1923 & x_1924;
assign x_8582 = x_1925 & x_1926;
assign x_8583 = x_8581 & x_8582;
assign x_8584 = x_8580 & x_8583;
assign x_8585 = x_8578 & x_8584;
assign x_8586 = x_8573 & x_8585;
assign x_8587 = x_8561 & x_8586;
assign x_8588 = x_1928 & x_1929;
assign x_8589 = x_1927 & x_8588;
assign x_8590 = x_1931 & x_1932;
assign x_8591 = x_1930 & x_8590;
assign x_8592 = x_8589 & x_8591;
assign x_8593 = x_1934 & x_1935;
assign x_8594 = x_1933 & x_8593;
assign x_8595 = x_1936 & x_1937;
assign x_8596 = x_1938 & x_1939;
assign x_8597 = x_8595 & x_8596;
assign x_8598 = x_8594 & x_8597;
assign x_8599 = x_8592 & x_8598;
assign x_8600 = x_1941 & x_1942;
assign x_8601 = x_1940 & x_8600;
assign x_8602 = x_1944 & x_1945;
assign x_8603 = x_1943 & x_8602;
assign x_8604 = x_8601 & x_8603;
assign x_8605 = x_1947 & x_1948;
assign x_8606 = x_1946 & x_8605;
assign x_8607 = x_1949 & x_1950;
assign x_8608 = x_1951 & x_1952;
assign x_8609 = x_8607 & x_8608;
assign x_8610 = x_8606 & x_8609;
assign x_8611 = x_8604 & x_8610;
assign x_8612 = x_8599 & x_8611;
assign x_8613 = x_1954 & x_1955;
assign x_8614 = x_1953 & x_8613;
assign x_8615 = x_1957 & x_1958;
assign x_8616 = x_1956 & x_8615;
assign x_8617 = x_8614 & x_8616;
assign x_8618 = x_1960 & x_1961;
assign x_8619 = x_1959 & x_8618;
assign x_8620 = x_1962 & x_1963;
assign x_8621 = x_1964 & x_1965;
assign x_8622 = x_8620 & x_8621;
assign x_8623 = x_8619 & x_8622;
assign x_8624 = x_8617 & x_8623;
assign x_8625 = x_1967 & x_1968;
assign x_8626 = x_1966 & x_8625;
assign x_8627 = x_1970 & x_1971;
assign x_8628 = x_1969 & x_8627;
assign x_8629 = x_8626 & x_8628;
assign x_8630 = x_1973 & x_1974;
assign x_8631 = x_1972 & x_8630;
assign x_8632 = x_1975 & x_1976;
assign x_8633 = x_1977 & x_1978;
assign x_8634 = x_8632 & x_8633;
assign x_8635 = x_8631 & x_8634;
assign x_8636 = x_8629 & x_8635;
assign x_8637 = x_8624 & x_8636;
assign x_8638 = x_8612 & x_8637;
assign x_8639 = x_8587 & x_8638;
assign x_8640 = x_1980 & x_1981;
assign x_8641 = x_1979 & x_8640;
assign x_8642 = x_1983 & x_1984;
assign x_8643 = x_1982 & x_8642;
assign x_8644 = x_8641 & x_8643;
assign x_8645 = x_1986 & x_1987;
assign x_8646 = x_1985 & x_8645;
assign x_8647 = x_1988 & x_1989;
assign x_8648 = x_1990 & x_1991;
assign x_8649 = x_8647 & x_8648;
assign x_8650 = x_8646 & x_8649;
assign x_8651 = x_8644 & x_8650;
assign x_8652 = x_1993 & x_1994;
assign x_8653 = x_1992 & x_8652;
assign x_8654 = x_1996 & x_1997;
assign x_8655 = x_1995 & x_8654;
assign x_8656 = x_8653 & x_8655;
assign x_8657 = x_1999 & x_2000;
assign x_8658 = x_1998 & x_8657;
assign x_8659 = x_2001 & x_2002;
assign x_8660 = x_2003 & x_2004;
assign x_8661 = x_8659 & x_8660;
assign x_8662 = x_8658 & x_8661;
assign x_8663 = x_8656 & x_8662;
assign x_8664 = x_8651 & x_8663;
assign x_8665 = x_2006 & x_2007;
assign x_8666 = x_2005 & x_8665;
assign x_8667 = x_2009 & x_2010;
assign x_8668 = x_2008 & x_8667;
assign x_8669 = x_8666 & x_8668;
assign x_8670 = x_2012 & x_2013;
assign x_8671 = x_2011 & x_8670;
assign x_8672 = x_2014 & x_2015;
assign x_8673 = x_2016 & x_2017;
assign x_8674 = x_8672 & x_8673;
assign x_8675 = x_8671 & x_8674;
assign x_8676 = x_8669 & x_8675;
assign x_8677 = x_2019 & x_2020;
assign x_8678 = x_2018 & x_8677;
assign x_8679 = x_2022 & x_2023;
assign x_8680 = x_2021 & x_8679;
assign x_8681 = x_8678 & x_8680;
assign x_8682 = x_2025 & x_2026;
assign x_8683 = x_2024 & x_8682;
assign x_8684 = x_2027 & x_2028;
assign x_8685 = x_2029 & x_2030;
assign x_8686 = x_8684 & x_8685;
assign x_8687 = x_8683 & x_8686;
assign x_8688 = x_8681 & x_8687;
assign x_8689 = x_8676 & x_8688;
assign x_8690 = x_8664 & x_8689;
assign x_8691 = x_2032 & x_2033;
assign x_8692 = x_2031 & x_8691;
assign x_8693 = x_2035 & x_2036;
assign x_8694 = x_2034 & x_8693;
assign x_8695 = x_8692 & x_8694;
assign x_8696 = x_2038 & x_2039;
assign x_8697 = x_2037 & x_8696;
assign x_8698 = x_2040 & x_2041;
assign x_8699 = x_2042 & x_2043;
assign x_8700 = x_8698 & x_8699;
assign x_8701 = x_8697 & x_8700;
assign x_8702 = x_8695 & x_8701;
assign x_8703 = x_2045 & x_2046;
assign x_8704 = x_2044 & x_8703;
assign x_8705 = x_2048 & x_2049;
assign x_8706 = x_2047 & x_8705;
assign x_8707 = x_8704 & x_8706;
assign x_8708 = x_2051 & x_2052;
assign x_8709 = x_2050 & x_8708;
assign x_8710 = x_2053 & x_2054;
assign x_8711 = x_2055 & x_2056;
assign x_8712 = x_8710 & x_8711;
assign x_8713 = x_8709 & x_8712;
assign x_8714 = x_8707 & x_8713;
assign x_8715 = x_8702 & x_8714;
assign x_8716 = x_2058 & x_2059;
assign x_8717 = x_2057 & x_8716;
assign x_8718 = x_2061 & x_2062;
assign x_8719 = x_2060 & x_8718;
assign x_8720 = x_8717 & x_8719;
assign x_8721 = x_2064 & x_2065;
assign x_8722 = x_2063 & x_8721;
assign x_8723 = x_2066 & x_2067;
assign x_8724 = x_2068 & x_2069;
assign x_8725 = x_8723 & x_8724;
assign x_8726 = x_8722 & x_8725;
assign x_8727 = x_8720 & x_8726;
assign x_8728 = x_2071 & x_2072;
assign x_8729 = x_2070 & x_8728;
assign x_8730 = x_2074 & x_2075;
assign x_8731 = x_2073 & x_8730;
assign x_8732 = x_8729 & x_8731;
assign x_8733 = x_2077 & x_2078;
assign x_8734 = x_2076 & x_8733;
assign x_8735 = x_2079 & x_2080;
assign x_8736 = x_2081 & x_2082;
assign x_8737 = x_8735 & x_8736;
assign x_8738 = x_8734 & x_8737;
assign x_8739 = x_8732 & x_8738;
assign x_8740 = x_8727 & x_8739;
assign x_8741 = x_8715 & x_8740;
assign x_8742 = x_8690 & x_8741;
assign x_8743 = x_8639 & x_8742;
assign x_8744 = x_8536 & x_8743;
assign x_8745 = x_2084 & x_2085;
assign x_8746 = x_2083 & x_8745;
assign x_8747 = x_2087 & x_2088;
assign x_8748 = x_2086 & x_8747;
assign x_8749 = x_8746 & x_8748;
assign x_8750 = x_2090 & x_2091;
assign x_8751 = x_2089 & x_8750;
assign x_8752 = x_2092 & x_2093;
assign x_8753 = x_2094 & x_2095;
assign x_8754 = x_8752 & x_8753;
assign x_8755 = x_8751 & x_8754;
assign x_8756 = x_8749 & x_8755;
assign x_8757 = x_2097 & x_2098;
assign x_8758 = x_2096 & x_8757;
assign x_8759 = x_2100 & x_2101;
assign x_8760 = x_2099 & x_8759;
assign x_8761 = x_8758 & x_8760;
assign x_8762 = x_2103 & x_2104;
assign x_8763 = x_2102 & x_8762;
assign x_8764 = x_2105 & x_2106;
assign x_8765 = x_2107 & x_2108;
assign x_8766 = x_8764 & x_8765;
assign x_8767 = x_8763 & x_8766;
assign x_8768 = x_8761 & x_8767;
assign x_8769 = x_8756 & x_8768;
assign x_8770 = x_2110 & x_2111;
assign x_8771 = x_2109 & x_8770;
assign x_8772 = x_2113 & x_2114;
assign x_8773 = x_2112 & x_8772;
assign x_8774 = x_8771 & x_8773;
assign x_8775 = x_2116 & x_2117;
assign x_8776 = x_2115 & x_8775;
assign x_8777 = x_2118 & x_2119;
assign x_8778 = x_2120 & x_2121;
assign x_8779 = x_8777 & x_8778;
assign x_8780 = x_8776 & x_8779;
assign x_8781 = x_8774 & x_8780;
assign x_8782 = x_2123 & x_2124;
assign x_8783 = x_2122 & x_8782;
assign x_8784 = x_2126 & x_2127;
assign x_8785 = x_2125 & x_8784;
assign x_8786 = x_8783 & x_8785;
assign x_8787 = x_2129 & x_2130;
assign x_8788 = x_2128 & x_8787;
assign x_8789 = x_2131 & x_2132;
assign x_8790 = x_2133 & x_2134;
assign x_8791 = x_8789 & x_8790;
assign x_8792 = x_8788 & x_8791;
assign x_8793 = x_8786 & x_8792;
assign x_8794 = x_8781 & x_8793;
assign x_8795 = x_8769 & x_8794;
assign x_8796 = x_2136 & x_2137;
assign x_8797 = x_2135 & x_8796;
assign x_8798 = x_2139 & x_2140;
assign x_8799 = x_2138 & x_8798;
assign x_8800 = x_8797 & x_8799;
assign x_8801 = x_2142 & x_2143;
assign x_8802 = x_2141 & x_8801;
assign x_8803 = x_2144 & x_2145;
assign x_8804 = x_2146 & x_2147;
assign x_8805 = x_8803 & x_8804;
assign x_8806 = x_8802 & x_8805;
assign x_8807 = x_8800 & x_8806;
assign x_8808 = x_2149 & x_2150;
assign x_8809 = x_2148 & x_8808;
assign x_8810 = x_2152 & x_2153;
assign x_8811 = x_2151 & x_8810;
assign x_8812 = x_8809 & x_8811;
assign x_8813 = x_2155 & x_2156;
assign x_8814 = x_2154 & x_8813;
assign x_8815 = x_2157 & x_2158;
assign x_8816 = x_2159 & x_2160;
assign x_8817 = x_8815 & x_8816;
assign x_8818 = x_8814 & x_8817;
assign x_8819 = x_8812 & x_8818;
assign x_8820 = x_8807 & x_8819;
assign x_8821 = x_2162 & x_2163;
assign x_8822 = x_2161 & x_8821;
assign x_8823 = x_2165 & x_2166;
assign x_8824 = x_2164 & x_8823;
assign x_8825 = x_8822 & x_8824;
assign x_8826 = x_2168 & x_2169;
assign x_8827 = x_2167 & x_8826;
assign x_8828 = x_2170 & x_2171;
assign x_8829 = x_2172 & x_2173;
assign x_8830 = x_8828 & x_8829;
assign x_8831 = x_8827 & x_8830;
assign x_8832 = x_8825 & x_8831;
assign x_8833 = x_2175 & x_2176;
assign x_8834 = x_2174 & x_8833;
assign x_8835 = x_2178 & x_2179;
assign x_8836 = x_2177 & x_8835;
assign x_8837 = x_8834 & x_8836;
assign x_8838 = x_2181 & x_2182;
assign x_8839 = x_2180 & x_8838;
assign x_8840 = x_2183 & x_2184;
assign x_8841 = x_2185 & x_2186;
assign x_8842 = x_8840 & x_8841;
assign x_8843 = x_8839 & x_8842;
assign x_8844 = x_8837 & x_8843;
assign x_8845 = x_8832 & x_8844;
assign x_8846 = x_8820 & x_8845;
assign x_8847 = x_8795 & x_8846;
assign x_8848 = x_2188 & x_2189;
assign x_8849 = x_2187 & x_8848;
assign x_8850 = x_2191 & x_2192;
assign x_8851 = x_2190 & x_8850;
assign x_8852 = x_8849 & x_8851;
assign x_8853 = x_2194 & x_2195;
assign x_8854 = x_2193 & x_8853;
assign x_8855 = x_2196 & x_2197;
assign x_8856 = x_2198 & x_2199;
assign x_8857 = x_8855 & x_8856;
assign x_8858 = x_8854 & x_8857;
assign x_8859 = x_8852 & x_8858;
assign x_8860 = x_2201 & x_2202;
assign x_8861 = x_2200 & x_8860;
assign x_8862 = x_2204 & x_2205;
assign x_8863 = x_2203 & x_8862;
assign x_8864 = x_8861 & x_8863;
assign x_8865 = x_2207 & x_2208;
assign x_8866 = x_2206 & x_8865;
assign x_8867 = x_2209 & x_2210;
assign x_8868 = x_2211 & x_2212;
assign x_8869 = x_8867 & x_8868;
assign x_8870 = x_8866 & x_8869;
assign x_8871 = x_8864 & x_8870;
assign x_8872 = x_8859 & x_8871;
assign x_8873 = x_2214 & x_2215;
assign x_8874 = x_2213 & x_8873;
assign x_8875 = x_2217 & x_2218;
assign x_8876 = x_2216 & x_8875;
assign x_8877 = x_8874 & x_8876;
assign x_8878 = x_2220 & x_2221;
assign x_8879 = x_2219 & x_8878;
assign x_8880 = x_2222 & x_2223;
assign x_8881 = x_2224 & x_2225;
assign x_8882 = x_8880 & x_8881;
assign x_8883 = x_8879 & x_8882;
assign x_8884 = x_8877 & x_8883;
assign x_8885 = x_2227 & x_2228;
assign x_8886 = x_2226 & x_8885;
assign x_8887 = x_2230 & x_2231;
assign x_8888 = x_2229 & x_8887;
assign x_8889 = x_8886 & x_8888;
assign x_8890 = x_2233 & x_2234;
assign x_8891 = x_2232 & x_8890;
assign x_8892 = x_2235 & x_2236;
assign x_8893 = x_2237 & x_2238;
assign x_8894 = x_8892 & x_8893;
assign x_8895 = x_8891 & x_8894;
assign x_8896 = x_8889 & x_8895;
assign x_8897 = x_8884 & x_8896;
assign x_8898 = x_8872 & x_8897;
assign x_8899 = x_2240 & x_2241;
assign x_8900 = x_2239 & x_8899;
assign x_8901 = x_2243 & x_2244;
assign x_8902 = x_2242 & x_8901;
assign x_8903 = x_8900 & x_8902;
assign x_8904 = x_2246 & x_2247;
assign x_8905 = x_2245 & x_8904;
assign x_8906 = x_2248 & x_2249;
assign x_8907 = x_2250 & x_2251;
assign x_8908 = x_8906 & x_8907;
assign x_8909 = x_8905 & x_8908;
assign x_8910 = x_8903 & x_8909;
assign x_8911 = x_2253 & x_2254;
assign x_8912 = x_2252 & x_8911;
assign x_8913 = x_2256 & x_2257;
assign x_8914 = x_2255 & x_8913;
assign x_8915 = x_8912 & x_8914;
assign x_8916 = x_2259 & x_2260;
assign x_8917 = x_2258 & x_8916;
assign x_8918 = x_2261 & x_2262;
assign x_8919 = x_2263 & x_2264;
assign x_8920 = x_8918 & x_8919;
assign x_8921 = x_8917 & x_8920;
assign x_8922 = x_8915 & x_8921;
assign x_8923 = x_8910 & x_8922;
assign x_8924 = x_2266 & x_2267;
assign x_8925 = x_2265 & x_8924;
assign x_8926 = x_2269 & x_2270;
assign x_8927 = x_2268 & x_8926;
assign x_8928 = x_8925 & x_8927;
assign x_8929 = x_2272 & x_2273;
assign x_8930 = x_2271 & x_8929;
assign x_8931 = x_2274 & x_2275;
assign x_8932 = x_2276 & x_2277;
assign x_8933 = x_8931 & x_8932;
assign x_8934 = x_8930 & x_8933;
assign x_8935 = x_8928 & x_8934;
assign x_8936 = x_2279 & x_2280;
assign x_8937 = x_2278 & x_8936;
assign x_8938 = x_2282 & x_2283;
assign x_8939 = x_2281 & x_8938;
assign x_8940 = x_8937 & x_8939;
assign x_8941 = x_2285 & x_2286;
assign x_8942 = x_2284 & x_8941;
assign x_8943 = x_2287 & x_2288;
assign x_8944 = x_2289 & x_2290;
assign x_8945 = x_8943 & x_8944;
assign x_8946 = x_8942 & x_8945;
assign x_8947 = x_8940 & x_8946;
assign x_8948 = x_8935 & x_8947;
assign x_8949 = x_8923 & x_8948;
assign x_8950 = x_8898 & x_8949;
assign x_8951 = x_8847 & x_8950;
assign x_8952 = x_2292 & x_2293;
assign x_8953 = x_2291 & x_8952;
assign x_8954 = x_2295 & x_2296;
assign x_8955 = x_2294 & x_8954;
assign x_8956 = x_8953 & x_8955;
assign x_8957 = x_2298 & x_2299;
assign x_8958 = x_2297 & x_8957;
assign x_8959 = x_2300 & x_2301;
assign x_8960 = x_2302 & x_2303;
assign x_8961 = x_8959 & x_8960;
assign x_8962 = x_8958 & x_8961;
assign x_8963 = x_8956 & x_8962;
assign x_8964 = x_2305 & x_2306;
assign x_8965 = x_2304 & x_8964;
assign x_8966 = x_2308 & x_2309;
assign x_8967 = x_2307 & x_8966;
assign x_8968 = x_8965 & x_8967;
assign x_8969 = x_2311 & x_2312;
assign x_8970 = x_2310 & x_8969;
assign x_8971 = x_2313 & x_2314;
assign x_8972 = x_2315 & x_2316;
assign x_8973 = x_8971 & x_8972;
assign x_8974 = x_8970 & x_8973;
assign x_8975 = x_8968 & x_8974;
assign x_8976 = x_8963 & x_8975;
assign x_8977 = x_2318 & x_2319;
assign x_8978 = x_2317 & x_8977;
assign x_8979 = x_2321 & x_2322;
assign x_8980 = x_2320 & x_8979;
assign x_8981 = x_8978 & x_8980;
assign x_8982 = x_2324 & x_2325;
assign x_8983 = x_2323 & x_8982;
assign x_8984 = x_2326 & x_2327;
assign x_8985 = x_2328 & x_2329;
assign x_8986 = x_8984 & x_8985;
assign x_8987 = x_8983 & x_8986;
assign x_8988 = x_8981 & x_8987;
assign x_8989 = x_2331 & x_2332;
assign x_8990 = x_2330 & x_8989;
assign x_8991 = x_2334 & x_2335;
assign x_8992 = x_2333 & x_8991;
assign x_8993 = x_8990 & x_8992;
assign x_8994 = x_2337 & x_2338;
assign x_8995 = x_2336 & x_8994;
assign x_8996 = x_2339 & x_2340;
assign x_8997 = x_2341 & x_2342;
assign x_8998 = x_8996 & x_8997;
assign x_8999 = x_8995 & x_8998;
assign x_9000 = x_8993 & x_8999;
assign x_9001 = x_8988 & x_9000;
assign x_9002 = x_8976 & x_9001;
assign x_9003 = x_2344 & x_2345;
assign x_9004 = x_2343 & x_9003;
assign x_9005 = x_2347 & x_2348;
assign x_9006 = x_2346 & x_9005;
assign x_9007 = x_9004 & x_9006;
assign x_9008 = x_2350 & x_2351;
assign x_9009 = x_2349 & x_9008;
assign x_9010 = x_2352 & x_2353;
assign x_9011 = x_2354 & x_2355;
assign x_9012 = x_9010 & x_9011;
assign x_9013 = x_9009 & x_9012;
assign x_9014 = x_9007 & x_9013;
assign x_9015 = x_2357 & x_2358;
assign x_9016 = x_2356 & x_9015;
assign x_9017 = x_2360 & x_2361;
assign x_9018 = x_2359 & x_9017;
assign x_9019 = x_9016 & x_9018;
assign x_9020 = x_2363 & x_2364;
assign x_9021 = x_2362 & x_9020;
assign x_9022 = x_2365 & x_2366;
assign x_9023 = x_2367 & x_2368;
assign x_9024 = x_9022 & x_9023;
assign x_9025 = x_9021 & x_9024;
assign x_9026 = x_9019 & x_9025;
assign x_9027 = x_9014 & x_9026;
assign x_9028 = x_2370 & x_2371;
assign x_9029 = x_2369 & x_9028;
assign x_9030 = x_2373 & x_2374;
assign x_9031 = x_2372 & x_9030;
assign x_9032 = x_9029 & x_9031;
assign x_9033 = x_2376 & x_2377;
assign x_9034 = x_2375 & x_9033;
assign x_9035 = x_2378 & x_2379;
assign x_9036 = x_2380 & x_2381;
assign x_9037 = x_9035 & x_9036;
assign x_9038 = x_9034 & x_9037;
assign x_9039 = x_9032 & x_9038;
assign x_9040 = x_2383 & x_2384;
assign x_9041 = x_2382 & x_9040;
assign x_9042 = x_2386 & x_2387;
assign x_9043 = x_2385 & x_9042;
assign x_9044 = x_9041 & x_9043;
assign x_9045 = x_2389 & x_2390;
assign x_9046 = x_2388 & x_9045;
assign x_9047 = x_2391 & x_2392;
assign x_9048 = x_2393 & x_2394;
assign x_9049 = x_9047 & x_9048;
assign x_9050 = x_9046 & x_9049;
assign x_9051 = x_9044 & x_9050;
assign x_9052 = x_9039 & x_9051;
assign x_9053 = x_9027 & x_9052;
assign x_9054 = x_9002 & x_9053;
assign x_9055 = x_2396 & x_2397;
assign x_9056 = x_2395 & x_9055;
assign x_9057 = x_2399 & x_2400;
assign x_9058 = x_2398 & x_9057;
assign x_9059 = x_9056 & x_9058;
assign x_9060 = x_2402 & x_2403;
assign x_9061 = x_2401 & x_9060;
assign x_9062 = x_2404 & x_2405;
assign x_9063 = x_2406 & x_2407;
assign x_9064 = x_9062 & x_9063;
assign x_9065 = x_9061 & x_9064;
assign x_9066 = x_9059 & x_9065;
assign x_9067 = x_2409 & x_2410;
assign x_9068 = x_2408 & x_9067;
assign x_9069 = x_2412 & x_2413;
assign x_9070 = x_2411 & x_9069;
assign x_9071 = x_9068 & x_9070;
assign x_9072 = x_2415 & x_2416;
assign x_9073 = x_2414 & x_9072;
assign x_9074 = x_2417 & x_2418;
assign x_9075 = x_2419 & x_2420;
assign x_9076 = x_9074 & x_9075;
assign x_9077 = x_9073 & x_9076;
assign x_9078 = x_9071 & x_9077;
assign x_9079 = x_9066 & x_9078;
assign x_9080 = x_2422 & x_2423;
assign x_9081 = x_2421 & x_9080;
assign x_9082 = x_2425 & x_2426;
assign x_9083 = x_2424 & x_9082;
assign x_9084 = x_9081 & x_9083;
assign x_9085 = x_2428 & x_2429;
assign x_9086 = x_2427 & x_9085;
assign x_9087 = x_2430 & x_2431;
assign x_9088 = x_2432 & x_2433;
assign x_9089 = x_9087 & x_9088;
assign x_9090 = x_9086 & x_9089;
assign x_9091 = x_9084 & x_9090;
assign x_9092 = x_2435 & x_2436;
assign x_9093 = x_2434 & x_9092;
assign x_9094 = x_2438 & x_2439;
assign x_9095 = x_2437 & x_9094;
assign x_9096 = x_9093 & x_9095;
assign x_9097 = x_2441 & x_2442;
assign x_9098 = x_2440 & x_9097;
assign x_9099 = x_2443 & x_2444;
assign x_9100 = x_2445 & x_2446;
assign x_9101 = x_9099 & x_9100;
assign x_9102 = x_9098 & x_9101;
assign x_9103 = x_9096 & x_9102;
assign x_9104 = x_9091 & x_9103;
assign x_9105 = x_9079 & x_9104;
assign x_9106 = x_2448 & x_2449;
assign x_9107 = x_2447 & x_9106;
assign x_9108 = x_2451 & x_2452;
assign x_9109 = x_2450 & x_9108;
assign x_9110 = x_9107 & x_9109;
assign x_9111 = x_2454 & x_2455;
assign x_9112 = x_2453 & x_9111;
assign x_9113 = x_2456 & x_2457;
assign x_9114 = x_2458 & x_2459;
assign x_9115 = x_9113 & x_9114;
assign x_9116 = x_9112 & x_9115;
assign x_9117 = x_9110 & x_9116;
assign x_9118 = x_2461 & x_2462;
assign x_9119 = x_2460 & x_9118;
assign x_9120 = x_2464 & x_2465;
assign x_9121 = x_2463 & x_9120;
assign x_9122 = x_9119 & x_9121;
assign x_9123 = x_2467 & x_2468;
assign x_9124 = x_2466 & x_9123;
assign x_9125 = x_2469 & x_2470;
assign x_9126 = x_2471 & x_2472;
assign x_9127 = x_9125 & x_9126;
assign x_9128 = x_9124 & x_9127;
assign x_9129 = x_9122 & x_9128;
assign x_9130 = x_9117 & x_9129;
assign x_9131 = x_2474 & x_2475;
assign x_9132 = x_2473 & x_9131;
assign x_9133 = x_2477 & x_2478;
assign x_9134 = x_2476 & x_9133;
assign x_9135 = x_9132 & x_9134;
assign x_9136 = x_2480 & x_2481;
assign x_9137 = x_2479 & x_9136;
assign x_9138 = x_2482 & x_2483;
assign x_9139 = x_2484 & x_2485;
assign x_9140 = x_9138 & x_9139;
assign x_9141 = x_9137 & x_9140;
assign x_9142 = x_9135 & x_9141;
assign x_9143 = x_2487 & x_2488;
assign x_9144 = x_2486 & x_9143;
assign x_9145 = x_2489 & x_2490;
assign x_9146 = x_2491 & x_2492;
assign x_9147 = x_9145 & x_9146;
assign x_9148 = x_9144 & x_9147;
assign x_9149 = x_2494 & x_2495;
assign x_9150 = x_2493 & x_9149;
assign x_9151 = x_2496 & x_2497;
assign x_9152 = x_2498 & x_2499;
assign x_9153 = x_9151 & x_9152;
assign x_9154 = x_9150 & x_9153;
assign x_9155 = x_9148 & x_9154;
assign x_9156 = x_9142 & x_9155;
assign x_9157 = x_9130 & x_9156;
assign x_9158 = x_9105 & x_9157;
assign x_9159 = x_9054 & x_9158;
assign x_9160 = x_8951 & x_9159;
assign x_9161 = x_8744 & x_9160;
assign x_9162 = x_2501 & x_2502;
assign x_9163 = x_2500 & x_9162;
assign x_9164 = x_2504 & x_2505;
assign x_9165 = x_2503 & x_9164;
assign x_9166 = x_9163 & x_9165;
assign x_9167 = x_2507 & x_2508;
assign x_9168 = x_2506 & x_9167;
assign x_9169 = x_2509 & x_2510;
assign x_9170 = x_2511 & x_2512;
assign x_9171 = x_9169 & x_9170;
assign x_9172 = x_9168 & x_9171;
assign x_9173 = x_9166 & x_9172;
assign x_9174 = x_2514 & x_2515;
assign x_9175 = x_2513 & x_9174;
assign x_9176 = x_2517 & x_2518;
assign x_9177 = x_2516 & x_9176;
assign x_9178 = x_9175 & x_9177;
assign x_9179 = x_2520 & x_2521;
assign x_9180 = x_2519 & x_9179;
assign x_9181 = x_2522 & x_2523;
assign x_9182 = x_2524 & x_2525;
assign x_9183 = x_9181 & x_9182;
assign x_9184 = x_9180 & x_9183;
assign x_9185 = x_9178 & x_9184;
assign x_9186 = x_9173 & x_9185;
assign x_9187 = x_2527 & x_2528;
assign x_9188 = x_2526 & x_9187;
assign x_9189 = x_2530 & x_2531;
assign x_9190 = x_2529 & x_9189;
assign x_9191 = x_9188 & x_9190;
assign x_9192 = x_2533 & x_2534;
assign x_9193 = x_2532 & x_9192;
assign x_9194 = x_2535 & x_2536;
assign x_9195 = x_2537 & x_2538;
assign x_9196 = x_9194 & x_9195;
assign x_9197 = x_9193 & x_9196;
assign x_9198 = x_9191 & x_9197;
assign x_9199 = x_2540 & x_2541;
assign x_9200 = x_2539 & x_9199;
assign x_9201 = x_2543 & x_2544;
assign x_9202 = x_2542 & x_9201;
assign x_9203 = x_9200 & x_9202;
assign x_9204 = x_2546 & x_2547;
assign x_9205 = x_2545 & x_9204;
assign x_9206 = x_2548 & x_2549;
assign x_9207 = x_2550 & x_2551;
assign x_9208 = x_9206 & x_9207;
assign x_9209 = x_9205 & x_9208;
assign x_9210 = x_9203 & x_9209;
assign x_9211 = x_9198 & x_9210;
assign x_9212 = x_9186 & x_9211;
assign x_9213 = x_2553 & x_2554;
assign x_9214 = x_2552 & x_9213;
assign x_9215 = x_2556 & x_2557;
assign x_9216 = x_2555 & x_9215;
assign x_9217 = x_9214 & x_9216;
assign x_9218 = x_2559 & x_2560;
assign x_9219 = x_2558 & x_9218;
assign x_9220 = x_2561 & x_2562;
assign x_9221 = x_2563 & x_2564;
assign x_9222 = x_9220 & x_9221;
assign x_9223 = x_9219 & x_9222;
assign x_9224 = x_9217 & x_9223;
assign x_9225 = x_2566 & x_2567;
assign x_9226 = x_2565 & x_9225;
assign x_9227 = x_2569 & x_2570;
assign x_9228 = x_2568 & x_9227;
assign x_9229 = x_9226 & x_9228;
assign x_9230 = x_2572 & x_2573;
assign x_9231 = x_2571 & x_9230;
assign x_9232 = x_2574 & x_2575;
assign x_9233 = x_2576 & x_2577;
assign x_9234 = x_9232 & x_9233;
assign x_9235 = x_9231 & x_9234;
assign x_9236 = x_9229 & x_9235;
assign x_9237 = x_9224 & x_9236;
assign x_9238 = x_2579 & x_2580;
assign x_9239 = x_2578 & x_9238;
assign x_9240 = x_2582 & x_2583;
assign x_9241 = x_2581 & x_9240;
assign x_9242 = x_9239 & x_9241;
assign x_9243 = x_2585 & x_2586;
assign x_9244 = x_2584 & x_9243;
assign x_9245 = x_2587 & x_2588;
assign x_9246 = x_2589 & x_2590;
assign x_9247 = x_9245 & x_9246;
assign x_9248 = x_9244 & x_9247;
assign x_9249 = x_9242 & x_9248;
assign x_9250 = x_2592 & x_2593;
assign x_9251 = x_2591 & x_9250;
assign x_9252 = x_2595 & x_2596;
assign x_9253 = x_2594 & x_9252;
assign x_9254 = x_9251 & x_9253;
assign x_9255 = x_2598 & x_2599;
assign x_9256 = x_2597 & x_9255;
assign x_9257 = x_2600 & x_2601;
assign x_9258 = x_2602 & x_2603;
assign x_9259 = x_9257 & x_9258;
assign x_9260 = x_9256 & x_9259;
assign x_9261 = x_9254 & x_9260;
assign x_9262 = x_9249 & x_9261;
assign x_9263 = x_9237 & x_9262;
assign x_9264 = x_9212 & x_9263;
assign x_9265 = x_2605 & x_2606;
assign x_9266 = x_2604 & x_9265;
assign x_9267 = x_2608 & x_2609;
assign x_9268 = x_2607 & x_9267;
assign x_9269 = x_9266 & x_9268;
assign x_9270 = x_2611 & x_2612;
assign x_9271 = x_2610 & x_9270;
assign x_9272 = x_2613 & x_2614;
assign x_9273 = x_2615 & x_2616;
assign x_9274 = x_9272 & x_9273;
assign x_9275 = x_9271 & x_9274;
assign x_9276 = x_9269 & x_9275;
assign x_9277 = x_2618 & x_2619;
assign x_9278 = x_2617 & x_9277;
assign x_9279 = x_2621 & x_2622;
assign x_9280 = x_2620 & x_9279;
assign x_9281 = x_9278 & x_9280;
assign x_9282 = x_2624 & x_2625;
assign x_9283 = x_2623 & x_9282;
assign x_9284 = x_2626 & x_2627;
assign x_9285 = x_2628 & x_2629;
assign x_9286 = x_9284 & x_9285;
assign x_9287 = x_9283 & x_9286;
assign x_9288 = x_9281 & x_9287;
assign x_9289 = x_9276 & x_9288;
assign x_9290 = x_2631 & x_2632;
assign x_9291 = x_2630 & x_9290;
assign x_9292 = x_2634 & x_2635;
assign x_9293 = x_2633 & x_9292;
assign x_9294 = x_9291 & x_9293;
assign x_9295 = x_2637 & x_2638;
assign x_9296 = x_2636 & x_9295;
assign x_9297 = x_2639 & x_2640;
assign x_9298 = x_2641 & x_2642;
assign x_9299 = x_9297 & x_9298;
assign x_9300 = x_9296 & x_9299;
assign x_9301 = x_9294 & x_9300;
assign x_9302 = x_2644 & x_2645;
assign x_9303 = x_2643 & x_9302;
assign x_9304 = x_2647 & x_2648;
assign x_9305 = x_2646 & x_9304;
assign x_9306 = x_9303 & x_9305;
assign x_9307 = x_2650 & x_2651;
assign x_9308 = x_2649 & x_9307;
assign x_9309 = x_2652 & x_2653;
assign x_9310 = x_2654 & x_2655;
assign x_9311 = x_9309 & x_9310;
assign x_9312 = x_9308 & x_9311;
assign x_9313 = x_9306 & x_9312;
assign x_9314 = x_9301 & x_9313;
assign x_9315 = x_9289 & x_9314;
assign x_9316 = x_2657 & x_2658;
assign x_9317 = x_2656 & x_9316;
assign x_9318 = x_2660 & x_2661;
assign x_9319 = x_2659 & x_9318;
assign x_9320 = x_9317 & x_9319;
assign x_9321 = x_2663 & x_2664;
assign x_9322 = x_2662 & x_9321;
assign x_9323 = x_2665 & x_2666;
assign x_9324 = x_2667 & x_2668;
assign x_9325 = x_9323 & x_9324;
assign x_9326 = x_9322 & x_9325;
assign x_9327 = x_9320 & x_9326;
assign x_9328 = x_2670 & x_2671;
assign x_9329 = x_2669 & x_9328;
assign x_9330 = x_2673 & x_2674;
assign x_9331 = x_2672 & x_9330;
assign x_9332 = x_9329 & x_9331;
assign x_9333 = x_2676 & x_2677;
assign x_9334 = x_2675 & x_9333;
assign x_9335 = x_2678 & x_2679;
assign x_9336 = x_2680 & x_2681;
assign x_9337 = x_9335 & x_9336;
assign x_9338 = x_9334 & x_9337;
assign x_9339 = x_9332 & x_9338;
assign x_9340 = x_9327 & x_9339;
assign x_9341 = x_2683 & x_2684;
assign x_9342 = x_2682 & x_9341;
assign x_9343 = x_2686 & x_2687;
assign x_9344 = x_2685 & x_9343;
assign x_9345 = x_9342 & x_9344;
assign x_9346 = x_2689 & x_2690;
assign x_9347 = x_2688 & x_9346;
assign x_9348 = x_2691 & x_2692;
assign x_9349 = x_2693 & x_2694;
assign x_9350 = x_9348 & x_9349;
assign x_9351 = x_9347 & x_9350;
assign x_9352 = x_9345 & x_9351;
assign x_9353 = x_2696 & x_2697;
assign x_9354 = x_2695 & x_9353;
assign x_9355 = x_2699 & x_2700;
assign x_9356 = x_2698 & x_9355;
assign x_9357 = x_9354 & x_9356;
assign x_9358 = x_2702 & x_2703;
assign x_9359 = x_2701 & x_9358;
assign x_9360 = x_2704 & x_2705;
assign x_9361 = x_2706 & x_2707;
assign x_9362 = x_9360 & x_9361;
assign x_9363 = x_9359 & x_9362;
assign x_9364 = x_9357 & x_9363;
assign x_9365 = x_9352 & x_9364;
assign x_9366 = x_9340 & x_9365;
assign x_9367 = x_9315 & x_9366;
assign x_9368 = x_9264 & x_9367;
assign x_9369 = x_2709 & x_2710;
assign x_9370 = x_2708 & x_9369;
assign x_9371 = x_2712 & x_2713;
assign x_9372 = x_2711 & x_9371;
assign x_9373 = x_9370 & x_9372;
assign x_9374 = x_2715 & x_2716;
assign x_9375 = x_2714 & x_9374;
assign x_9376 = x_2717 & x_2718;
assign x_9377 = x_2719 & x_2720;
assign x_9378 = x_9376 & x_9377;
assign x_9379 = x_9375 & x_9378;
assign x_9380 = x_9373 & x_9379;
assign x_9381 = x_2722 & x_2723;
assign x_9382 = x_2721 & x_9381;
assign x_9383 = x_2725 & x_2726;
assign x_9384 = x_2724 & x_9383;
assign x_9385 = x_9382 & x_9384;
assign x_9386 = x_2728 & x_2729;
assign x_9387 = x_2727 & x_9386;
assign x_9388 = x_2730 & x_2731;
assign x_9389 = x_2732 & x_2733;
assign x_9390 = x_9388 & x_9389;
assign x_9391 = x_9387 & x_9390;
assign x_9392 = x_9385 & x_9391;
assign x_9393 = x_9380 & x_9392;
assign x_9394 = x_2735 & x_2736;
assign x_9395 = x_2734 & x_9394;
assign x_9396 = x_2738 & x_2739;
assign x_9397 = x_2737 & x_9396;
assign x_9398 = x_9395 & x_9397;
assign x_9399 = x_2741 & x_2742;
assign x_9400 = x_2740 & x_9399;
assign x_9401 = x_2743 & x_2744;
assign x_9402 = x_2745 & x_2746;
assign x_9403 = x_9401 & x_9402;
assign x_9404 = x_9400 & x_9403;
assign x_9405 = x_9398 & x_9404;
assign x_9406 = x_2748 & x_2749;
assign x_9407 = x_2747 & x_9406;
assign x_9408 = x_2751 & x_2752;
assign x_9409 = x_2750 & x_9408;
assign x_9410 = x_9407 & x_9409;
assign x_9411 = x_2754 & x_2755;
assign x_9412 = x_2753 & x_9411;
assign x_9413 = x_2756 & x_2757;
assign x_9414 = x_2758 & x_2759;
assign x_9415 = x_9413 & x_9414;
assign x_9416 = x_9412 & x_9415;
assign x_9417 = x_9410 & x_9416;
assign x_9418 = x_9405 & x_9417;
assign x_9419 = x_9393 & x_9418;
assign x_9420 = x_2761 & x_2762;
assign x_9421 = x_2760 & x_9420;
assign x_9422 = x_2764 & x_2765;
assign x_9423 = x_2763 & x_9422;
assign x_9424 = x_9421 & x_9423;
assign x_9425 = x_2767 & x_2768;
assign x_9426 = x_2766 & x_9425;
assign x_9427 = x_2769 & x_2770;
assign x_9428 = x_2771 & x_2772;
assign x_9429 = x_9427 & x_9428;
assign x_9430 = x_9426 & x_9429;
assign x_9431 = x_9424 & x_9430;
assign x_9432 = x_2774 & x_2775;
assign x_9433 = x_2773 & x_9432;
assign x_9434 = x_2777 & x_2778;
assign x_9435 = x_2776 & x_9434;
assign x_9436 = x_9433 & x_9435;
assign x_9437 = x_2780 & x_2781;
assign x_9438 = x_2779 & x_9437;
assign x_9439 = x_2782 & x_2783;
assign x_9440 = x_2784 & x_2785;
assign x_9441 = x_9439 & x_9440;
assign x_9442 = x_9438 & x_9441;
assign x_9443 = x_9436 & x_9442;
assign x_9444 = x_9431 & x_9443;
assign x_9445 = x_2787 & x_2788;
assign x_9446 = x_2786 & x_9445;
assign x_9447 = x_2790 & x_2791;
assign x_9448 = x_2789 & x_9447;
assign x_9449 = x_9446 & x_9448;
assign x_9450 = x_2793 & x_2794;
assign x_9451 = x_2792 & x_9450;
assign x_9452 = x_2795 & x_2796;
assign x_9453 = x_2797 & x_2798;
assign x_9454 = x_9452 & x_9453;
assign x_9455 = x_9451 & x_9454;
assign x_9456 = x_9449 & x_9455;
assign x_9457 = x_2800 & x_2801;
assign x_9458 = x_2799 & x_9457;
assign x_9459 = x_2803 & x_2804;
assign x_9460 = x_2802 & x_9459;
assign x_9461 = x_9458 & x_9460;
assign x_9462 = x_2806 & x_2807;
assign x_9463 = x_2805 & x_9462;
assign x_9464 = x_2808 & x_2809;
assign x_9465 = x_2810 & x_2811;
assign x_9466 = x_9464 & x_9465;
assign x_9467 = x_9463 & x_9466;
assign x_9468 = x_9461 & x_9467;
assign x_9469 = x_9456 & x_9468;
assign x_9470 = x_9444 & x_9469;
assign x_9471 = x_9419 & x_9470;
assign x_9472 = x_2813 & x_2814;
assign x_9473 = x_2812 & x_9472;
assign x_9474 = x_2816 & x_2817;
assign x_9475 = x_2815 & x_9474;
assign x_9476 = x_9473 & x_9475;
assign x_9477 = x_2819 & x_2820;
assign x_9478 = x_2818 & x_9477;
assign x_9479 = x_2821 & x_2822;
assign x_9480 = x_2823 & x_2824;
assign x_9481 = x_9479 & x_9480;
assign x_9482 = x_9478 & x_9481;
assign x_9483 = x_9476 & x_9482;
assign x_9484 = x_2826 & x_2827;
assign x_9485 = x_2825 & x_9484;
assign x_9486 = x_2829 & x_2830;
assign x_9487 = x_2828 & x_9486;
assign x_9488 = x_9485 & x_9487;
assign x_9489 = x_2832 & x_2833;
assign x_9490 = x_2831 & x_9489;
assign x_9491 = x_2834 & x_2835;
assign x_9492 = x_2836 & x_2837;
assign x_9493 = x_9491 & x_9492;
assign x_9494 = x_9490 & x_9493;
assign x_9495 = x_9488 & x_9494;
assign x_9496 = x_9483 & x_9495;
assign x_9497 = x_2839 & x_2840;
assign x_9498 = x_2838 & x_9497;
assign x_9499 = x_2842 & x_2843;
assign x_9500 = x_2841 & x_9499;
assign x_9501 = x_9498 & x_9500;
assign x_9502 = x_2845 & x_2846;
assign x_9503 = x_2844 & x_9502;
assign x_9504 = x_2847 & x_2848;
assign x_9505 = x_2849 & x_2850;
assign x_9506 = x_9504 & x_9505;
assign x_9507 = x_9503 & x_9506;
assign x_9508 = x_9501 & x_9507;
assign x_9509 = x_2852 & x_2853;
assign x_9510 = x_2851 & x_9509;
assign x_9511 = x_2855 & x_2856;
assign x_9512 = x_2854 & x_9511;
assign x_9513 = x_9510 & x_9512;
assign x_9514 = x_2858 & x_2859;
assign x_9515 = x_2857 & x_9514;
assign x_9516 = x_2860 & x_2861;
assign x_9517 = x_2862 & x_2863;
assign x_9518 = x_9516 & x_9517;
assign x_9519 = x_9515 & x_9518;
assign x_9520 = x_9513 & x_9519;
assign x_9521 = x_9508 & x_9520;
assign x_9522 = x_9496 & x_9521;
assign x_9523 = x_2865 & x_2866;
assign x_9524 = x_2864 & x_9523;
assign x_9525 = x_2868 & x_2869;
assign x_9526 = x_2867 & x_9525;
assign x_9527 = x_9524 & x_9526;
assign x_9528 = x_2871 & x_2872;
assign x_9529 = x_2870 & x_9528;
assign x_9530 = x_2873 & x_2874;
assign x_9531 = x_2875 & x_2876;
assign x_9532 = x_9530 & x_9531;
assign x_9533 = x_9529 & x_9532;
assign x_9534 = x_9527 & x_9533;
assign x_9535 = x_2878 & x_2879;
assign x_9536 = x_2877 & x_9535;
assign x_9537 = x_2881 & x_2882;
assign x_9538 = x_2880 & x_9537;
assign x_9539 = x_9536 & x_9538;
assign x_9540 = x_2884 & x_2885;
assign x_9541 = x_2883 & x_9540;
assign x_9542 = x_2886 & x_2887;
assign x_9543 = x_2888 & x_2889;
assign x_9544 = x_9542 & x_9543;
assign x_9545 = x_9541 & x_9544;
assign x_9546 = x_9539 & x_9545;
assign x_9547 = x_9534 & x_9546;
assign x_9548 = x_2891 & x_2892;
assign x_9549 = x_2890 & x_9548;
assign x_9550 = x_2894 & x_2895;
assign x_9551 = x_2893 & x_9550;
assign x_9552 = x_9549 & x_9551;
assign x_9553 = x_2897 & x_2898;
assign x_9554 = x_2896 & x_9553;
assign x_9555 = x_2899 & x_2900;
assign x_9556 = x_2901 & x_2902;
assign x_9557 = x_9555 & x_9556;
assign x_9558 = x_9554 & x_9557;
assign x_9559 = x_9552 & x_9558;
assign x_9560 = x_2904 & x_2905;
assign x_9561 = x_2903 & x_9560;
assign x_9562 = x_2907 & x_2908;
assign x_9563 = x_2906 & x_9562;
assign x_9564 = x_9561 & x_9563;
assign x_9565 = x_2910 & x_2911;
assign x_9566 = x_2909 & x_9565;
assign x_9567 = x_2912 & x_2913;
assign x_9568 = x_2914 & x_2915;
assign x_9569 = x_9567 & x_9568;
assign x_9570 = x_9566 & x_9569;
assign x_9571 = x_9564 & x_9570;
assign x_9572 = x_9559 & x_9571;
assign x_9573 = x_9547 & x_9572;
assign x_9574 = x_9522 & x_9573;
assign x_9575 = x_9471 & x_9574;
assign x_9576 = x_9368 & x_9575;
assign x_9577 = x_2917 & x_2918;
assign x_9578 = x_2916 & x_9577;
assign x_9579 = x_2920 & x_2921;
assign x_9580 = x_2919 & x_9579;
assign x_9581 = x_9578 & x_9580;
assign x_9582 = x_2923 & x_2924;
assign x_9583 = x_2922 & x_9582;
assign x_9584 = x_2925 & x_2926;
assign x_9585 = x_2927 & x_2928;
assign x_9586 = x_9584 & x_9585;
assign x_9587 = x_9583 & x_9586;
assign x_9588 = x_9581 & x_9587;
assign x_9589 = x_2930 & x_2931;
assign x_9590 = x_2929 & x_9589;
assign x_9591 = x_2933 & x_2934;
assign x_9592 = x_2932 & x_9591;
assign x_9593 = x_9590 & x_9592;
assign x_9594 = x_2936 & x_2937;
assign x_9595 = x_2935 & x_9594;
assign x_9596 = x_2938 & x_2939;
assign x_9597 = x_2940 & x_2941;
assign x_9598 = x_9596 & x_9597;
assign x_9599 = x_9595 & x_9598;
assign x_9600 = x_9593 & x_9599;
assign x_9601 = x_9588 & x_9600;
assign x_9602 = x_2943 & x_2944;
assign x_9603 = x_2942 & x_9602;
assign x_9604 = x_2946 & x_2947;
assign x_9605 = x_2945 & x_9604;
assign x_9606 = x_9603 & x_9605;
assign x_9607 = x_2949 & x_2950;
assign x_9608 = x_2948 & x_9607;
assign x_9609 = x_2951 & x_2952;
assign x_9610 = x_2953 & x_2954;
assign x_9611 = x_9609 & x_9610;
assign x_9612 = x_9608 & x_9611;
assign x_9613 = x_9606 & x_9612;
assign x_9614 = x_2956 & x_2957;
assign x_9615 = x_2955 & x_9614;
assign x_9616 = x_2959 & x_2960;
assign x_9617 = x_2958 & x_9616;
assign x_9618 = x_9615 & x_9617;
assign x_9619 = x_2962 & x_2963;
assign x_9620 = x_2961 & x_9619;
assign x_9621 = x_2964 & x_2965;
assign x_9622 = x_2966 & x_2967;
assign x_9623 = x_9621 & x_9622;
assign x_9624 = x_9620 & x_9623;
assign x_9625 = x_9618 & x_9624;
assign x_9626 = x_9613 & x_9625;
assign x_9627 = x_9601 & x_9626;
assign x_9628 = x_2969 & x_2970;
assign x_9629 = x_2968 & x_9628;
assign x_9630 = x_2972 & x_2973;
assign x_9631 = x_2971 & x_9630;
assign x_9632 = x_9629 & x_9631;
assign x_9633 = x_2975 & x_2976;
assign x_9634 = x_2974 & x_9633;
assign x_9635 = x_2977 & x_2978;
assign x_9636 = x_2979 & x_2980;
assign x_9637 = x_9635 & x_9636;
assign x_9638 = x_9634 & x_9637;
assign x_9639 = x_9632 & x_9638;
assign x_9640 = x_2982 & x_2983;
assign x_9641 = x_2981 & x_9640;
assign x_9642 = x_2985 & x_2986;
assign x_9643 = x_2984 & x_9642;
assign x_9644 = x_9641 & x_9643;
assign x_9645 = x_2988 & x_2989;
assign x_9646 = x_2987 & x_9645;
assign x_9647 = x_2990 & x_2991;
assign x_9648 = x_2992 & x_2993;
assign x_9649 = x_9647 & x_9648;
assign x_9650 = x_9646 & x_9649;
assign x_9651 = x_9644 & x_9650;
assign x_9652 = x_9639 & x_9651;
assign x_9653 = x_2995 & x_2996;
assign x_9654 = x_2994 & x_9653;
assign x_9655 = x_2998 & x_2999;
assign x_9656 = x_2997 & x_9655;
assign x_9657 = x_9654 & x_9656;
assign x_9658 = x_3001 & x_3002;
assign x_9659 = x_3000 & x_9658;
assign x_9660 = x_3003 & x_3004;
assign x_9661 = x_3005 & x_3006;
assign x_9662 = x_9660 & x_9661;
assign x_9663 = x_9659 & x_9662;
assign x_9664 = x_9657 & x_9663;
assign x_9665 = x_3008 & x_3009;
assign x_9666 = x_3007 & x_9665;
assign x_9667 = x_3011 & x_3012;
assign x_9668 = x_3010 & x_9667;
assign x_9669 = x_9666 & x_9668;
assign x_9670 = x_3014 & x_3015;
assign x_9671 = x_3013 & x_9670;
assign x_9672 = x_3016 & x_3017;
assign x_9673 = x_3018 & x_3019;
assign x_9674 = x_9672 & x_9673;
assign x_9675 = x_9671 & x_9674;
assign x_9676 = x_9669 & x_9675;
assign x_9677 = x_9664 & x_9676;
assign x_9678 = x_9652 & x_9677;
assign x_9679 = x_9627 & x_9678;
assign x_9680 = x_3021 & x_3022;
assign x_9681 = x_3020 & x_9680;
assign x_9682 = x_3024 & x_3025;
assign x_9683 = x_3023 & x_9682;
assign x_9684 = x_9681 & x_9683;
assign x_9685 = x_3027 & x_3028;
assign x_9686 = x_3026 & x_9685;
assign x_9687 = x_3029 & x_3030;
assign x_9688 = x_3031 & x_3032;
assign x_9689 = x_9687 & x_9688;
assign x_9690 = x_9686 & x_9689;
assign x_9691 = x_9684 & x_9690;
assign x_9692 = x_3034 & x_3035;
assign x_9693 = x_3033 & x_9692;
assign x_9694 = x_3037 & x_3038;
assign x_9695 = x_3036 & x_9694;
assign x_9696 = x_9693 & x_9695;
assign x_9697 = x_3040 & x_3041;
assign x_9698 = x_3039 & x_9697;
assign x_9699 = x_3042 & x_3043;
assign x_9700 = x_3044 & x_3045;
assign x_9701 = x_9699 & x_9700;
assign x_9702 = x_9698 & x_9701;
assign x_9703 = x_9696 & x_9702;
assign x_9704 = x_9691 & x_9703;
assign x_9705 = x_3047 & x_3048;
assign x_9706 = x_3046 & x_9705;
assign x_9707 = x_3050 & x_3051;
assign x_9708 = x_3049 & x_9707;
assign x_9709 = x_9706 & x_9708;
assign x_9710 = x_3053 & x_3054;
assign x_9711 = x_3052 & x_9710;
assign x_9712 = x_3055 & x_3056;
assign x_9713 = x_3057 & x_3058;
assign x_9714 = x_9712 & x_9713;
assign x_9715 = x_9711 & x_9714;
assign x_9716 = x_9709 & x_9715;
assign x_9717 = x_3060 & x_3061;
assign x_9718 = x_3059 & x_9717;
assign x_9719 = x_3063 & x_3064;
assign x_9720 = x_3062 & x_9719;
assign x_9721 = x_9718 & x_9720;
assign x_9722 = x_3066 & x_3067;
assign x_9723 = x_3065 & x_9722;
assign x_9724 = x_3068 & x_3069;
assign x_9725 = x_3070 & x_3071;
assign x_9726 = x_9724 & x_9725;
assign x_9727 = x_9723 & x_9726;
assign x_9728 = x_9721 & x_9727;
assign x_9729 = x_9716 & x_9728;
assign x_9730 = x_9704 & x_9729;
assign x_9731 = x_3073 & x_3074;
assign x_9732 = x_3072 & x_9731;
assign x_9733 = x_3076 & x_3077;
assign x_9734 = x_3075 & x_9733;
assign x_9735 = x_9732 & x_9734;
assign x_9736 = x_3079 & x_3080;
assign x_9737 = x_3078 & x_9736;
assign x_9738 = x_3081 & x_3082;
assign x_9739 = x_3083 & x_3084;
assign x_9740 = x_9738 & x_9739;
assign x_9741 = x_9737 & x_9740;
assign x_9742 = x_9735 & x_9741;
assign x_9743 = x_3086 & x_3087;
assign x_9744 = x_3085 & x_9743;
assign x_9745 = x_3089 & x_3090;
assign x_9746 = x_3088 & x_9745;
assign x_9747 = x_9744 & x_9746;
assign x_9748 = x_3092 & x_3093;
assign x_9749 = x_3091 & x_9748;
assign x_9750 = x_3094 & x_3095;
assign x_9751 = x_3096 & x_3097;
assign x_9752 = x_9750 & x_9751;
assign x_9753 = x_9749 & x_9752;
assign x_9754 = x_9747 & x_9753;
assign x_9755 = x_9742 & x_9754;
assign x_9756 = x_3099 & x_3100;
assign x_9757 = x_3098 & x_9756;
assign x_9758 = x_3102 & x_3103;
assign x_9759 = x_3101 & x_9758;
assign x_9760 = x_9757 & x_9759;
assign x_9761 = x_3105 & x_3106;
assign x_9762 = x_3104 & x_9761;
assign x_9763 = x_3107 & x_3108;
assign x_9764 = x_3109 & x_3110;
assign x_9765 = x_9763 & x_9764;
assign x_9766 = x_9762 & x_9765;
assign x_9767 = x_9760 & x_9766;
assign x_9768 = x_3112 & x_3113;
assign x_9769 = x_3111 & x_9768;
assign x_9770 = x_3115 & x_3116;
assign x_9771 = x_3114 & x_9770;
assign x_9772 = x_9769 & x_9771;
assign x_9773 = x_3118 & x_3119;
assign x_9774 = x_3117 & x_9773;
assign x_9775 = x_3120 & x_3121;
assign x_9776 = x_3122 & x_3123;
assign x_9777 = x_9775 & x_9776;
assign x_9778 = x_9774 & x_9777;
assign x_9779 = x_9772 & x_9778;
assign x_9780 = x_9767 & x_9779;
assign x_9781 = x_9755 & x_9780;
assign x_9782 = x_9730 & x_9781;
assign x_9783 = x_9679 & x_9782;
assign x_9784 = x_3125 & x_3126;
assign x_9785 = x_3124 & x_9784;
assign x_9786 = x_3128 & x_3129;
assign x_9787 = x_3127 & x_9786;
assign x_9788 = x_9785 & x_9787;
assign x_9789 = x_3131 & x_3132;
assign x_9790 = x_3130 & x_9789;
assign x_9791 = x_3133 & x_3134;
assign x_9792 = x_3135 & x_3136;
assign x_9793 = x_9791 & x_9792;
assign x_9794 = x_9790 & x_9793;
assign x_9795 = x_9788 & x_9794;
assign x_9796 = x_3138 & x_3139;
assign x_9797 = x_3137 & x_9796;
assign x_9798 = x_3141 & x_3142;
assign x_9799 = x_3140 & x_9798;
assign x_9800 = x_9797 & x_9799;
assign x_9801 = x_3144 & x_3145;
assign x_9802 = x_3143 & x_9801;
assign x_9803 = x_3146 & x_3147;
assign x_9804 = x_3148 & x_3149;
assign x_9805 = x_9803 & x_9804;
assign x_9806 = x_9802 & x_9805;
assign x_9807 = x_9800 & x_9806;
assign x_9808 = x_9795 & x_9807;
assign x_9809 = x_3151 & x_3152;
assign x_9810 = x_3150 & x_9809;
assign x_9811 = x_3154 & x_3155;
assign x_9812 = x_3153 & x_9811;
assign x_9813 = x_9810 & x_9812;
assign x_9814 = x_3157 & x_3158;
assign x_9815 = x_3156 & x_9814;
assign x_9816 = x_3159 & x_3160;
assign x_9817 = x_3161 & x_3162;
assign x_9818 = x_9816 & x_9817;
assign x_9819 = x_9815 & x_9818;
assign x_9820 = x_9813 & x_9819;
assign x_9821 = x_3164 & x_3165;
assign x_9822 = x_3163 & x_9821;
assign x_9823 = x_3167 & x_3168;
assign x_9824 = x_3166 & x_9823;
assign x_9825 = x_9822 & x_9824;
assign x_9826 = x_3170 & x_3171;
assign x_9827 = x_3169 & x_9826;
assign x_9828 = x_3172 & x_3173;
assign x_9829 = x_3174 & x_3175;
assign x_9830 = x_9828 & x_9829;
assign x_9831 = x_9827 & x_9830;
assign x_9832 = x_9825 & x_9831;
assign x_9833 = x_9820 & x_9832;
assign x_9834 = x_9808 & x_9833;
assign x_9835 = x_3177 & x_3178;
assign x_9836 = x_3176 & x_9835;
assign x_9837 = x_3180 & x_3181;
assign x_9838 = x_3179 & x_9837;
assign x_9839 = x_9836 & x_9838;
assign x_9840 = x_3183 & x_3184;
assign x_9841 = x_3182 & x_9840;
assign x_9842 = x_3185 & x_3186;
assign x_9843 = x_3187 & x_3188;
assign x_9844 = x_9842 & x_9843;
assign x_9845 = x_9841 & x_9844;
assign x_9846 = x_9839 & x_9845;
assign x_9847 = x_3190 & x_3191;
assign x_9848 = x_3189 & x_9847;
assign x_9849 = x_3193 & x_3194;
assign x_9850 = x_3192 & x_9849;
assign x_9851 = x_9848 & x_9850;
assign x_9852 = x_3196 & x_3197;
assign x_9853 = x_3195 & x_9852;
assign x_9854 = x_3198 & x_3199;
assign x_9855 = x_3200 & x_3201;
assign x_9856 = x_9854 & x_9855;
assign x_9857 = x_9853 & x_9856;
assign x_9858 = x_9851 & x_9857;
assign x_9859 = x_9846 & x_9858;
assign x_9860 = x_3203 & x_3204;
assign x_9861 = x_3202 & x_9860;
assign x_9862 = x_3206 & x_3207;
assign x_9863 = x_3205 & x_9862;
assign x_9864 = x_9861 & x_9863;
assign x_9865 = x_3209 & x_3210;
assign x_9866 = x_3208 & x_9865;
assign x_9867 = x_3211 & x_3212;
assign x_9868 = x_3213 & x_3214;
assign x_9869 = x_9867 & x_9868;
assign x_9870 = x_9866 & x_9869;
assign x_9871 = x_9864 & x_9870;
assign x_9872 = x_3216 & x_3217;
assign x_9873 = x_3215 & x_9872;
assign x_9874 = x_3219 & x_3220;
assign x_9875 = x_3218 & x_9874;
assign x_9876 = x_9873 & x_9875;
assign x_9877 = x_3222 & x_3223;
assign x_9878 = x_3221 & x_9877;
assign x_9879 = x_3224 & x_3225;
assign x_9880 = x_3226 & x_3227;
assign x_9881 = x_9879 & x_9880;
assign x_9882 = x_9878 & x_9881;
assign x_9883 = x_9876 & x_9882;
assign x_9884 = x_9871 & x_9883;
assign x_9885 = x_9859 & x_9884;
assign x_9886 = x_9834 & x_9885;
assign x_9887 = x_3229 & x_3230;
assign x_9888 = x_3228 & x_9887;
assign x_9889 = x_3232 & x_3233;
assign x_9890 = x_3231 & x_9889;
assign x_9891 = x_9888 & x_9890;
assign x_9892 = x_3235 & x_3236;
assign x_9893 = x_3234 & x_9892;
assign x_9894 = x_3237 & x_3238;
assign x_9895 = x_3239 & x_3240;
assign x_9896 = x_9894 & x_9895;
assign x_9897 = x_9893 & x_9896;
assign x_9898 = x_9891 & x_9897;
assign x_9899 = x_3242 & x_3243;
assign x_9900 = x_3241 & x_9899;
assign x_9901 = x_3245 & x_3246;
assign x_9902 = x_3244 & x_9901;
assign x_9903 = x_9900 & x_9902;
assign x_9904 = x_3248 & x_3249;
assign x_9905 = x_3247 & x_9904;
assign x_9906 = x_3250 & x_3251;
assign x_9907 = x_3252 & x_3253;
assign x_9908 = x_9906 & x_9907;
assign x_9909 = x_9905 & x_9908;
assign x_9910 = x_9903 & x_9909;
assign x_9911 = x_9898 & x_9910;
assign x_9912 = x_3255 & x_3256;
assign x_9913 = x_3254 & x_9912;
assign x_9914 = x_3258 & x_3259;
assign x_9915 = x_3257 & x_9914;
assign x_9916 = x_9913 & x_9915;
assign x_9917 = x_3261 & x_3262;
assign x_9918 = x_3260 & x_9917;
assign x_9919 = x_3263 & x_3264;
assign x_9920 = x_3265 & x_3266;
assign x_9921 = x_9919 & x_9920;
assign x_9922 = x_9918 & x_9921;
assign x_9923 = x_9916 & x_9922;
assign x_9924 = x_3268 & x_3269;
assign x_9925 = x_3267 & x_9924;
assign x_9926 = x_3271 & x_3272;
assign x_9927 = x_3270 & x_9926;
assign x_9928 = x_9925 & x_9927;
assign x_9929 = x_3274 & x_3275;
assign x_9930 = x_3273 & x_9929;
assign x_9931 = x_3276 & x_3277;
assign x_9932 = x_3278 & x_3279;
assign x_9933 = x_9931 & x_9932;
assign x_9934 = x_9930 & x_9933;
assign x_9935 = x_9928 & x_9934;
assign x_9936 = x_9923 & x_9935;
assign x_9937 = x_9911 & x_9936;
assign x_9938 = x_3281 & x_3282;
assign x_9939 = x_3280 & x_9938;
assign x_9940 = x_3284 & x_3285;
assign x_9941 = x_3283 & x_9940;
assign x_9942 = x_9939 & x_9941;
assign x_9943 = x_3287 & x_3288;
assign x_9944 = x_3286 & x_9943;
assign x_9945 = x_3289 & x_3290;
assign x_9946 = x_3291 & x_3292;
assign x_9947 = x_9945 & x_9946;
assign x_9948 = x_9944 & x_9947;
assign x_9949 = x_9942 & x_9948;
assign x_9950 = x_3294 & x_3295;
assign x_9951 = x_3293 & x_9950;
assign x_9952 = x_3297 & x_3298;
assign x_9953 = x_3296 & x_9952;
assign x_9954 = x_9951 & x_9953;
assign x_9955 = x_3300 & x_3301;
assign x_9956 = x_3299 & x_9955;
assign x_9957 = x_3302 & x_3303;
assign x_9958 = x_3304 & x_3305;
assign x_9959 = x_9957 & x_9958;
assign x_9960 = x_9956 & x_9959;
assign x_9961 = x_9954 & x_9960;
assign x_9962 = x_9949 & x_9961;
assign x_9963 = x_3307 & x_3308;
assign x_9964 = x_3306 & x_9963;
assign x_9965 = x_3310 & x_3311;
assign x_9966 = x_3309 & x_9965;
assign x_9967 = x_9964 & x_9966;
assign x_9968 = x_3313 & x_3314;
assign x_9969 = x_3312 & x_9968;
assign x_9970 = x_3315 & x_3316;
assign x_9971 = x_3317 & x_3318;
assign x_9972 = x_9970 & x_9971;
assign x_9973 = x_9969 & x_9972;
assign x_9974 = x_9967 & x_9973;
assign x_9975 = x_3320 & x_3321;
assign x_9976 = x_3319 & x_9975;
assign x_9977 = x_3322 & x_3323;
assign x_9978 = x_3324 & x_3325;
assign x_9979 = x_9977 & x_9978;
assign x_9980 = x_9976 & x_9979;
assign x_9981 = x_3327 & x_3328;
assign x_9982 = x_3326 & x_9981;
assign x_9983 = x_3329 & x_3330;
assign x_9984 = x_3331 & x_3332;
assign x_9985 = x_9983 & x_9984;
assign x_9986 = x_9982 & x_9985;
assign x_9987 = x_9980 & x_9986;
assign x_9988 = x_9974 & x_9987;
assign x_9989 = x_9962 & x_9988;
assign x_9990 = x_9937 & x_9989;
assign x_9991 = x_9886 & x_9990;
assign x_9992 = x_9783 & x_9991;
assign x_9993 = x_9576 & x_9992;
assign x_9994 = x_9161 & x_9993;
assign x_9995 = x_8329 & x_9994;
assign x_9996 = x_3334 & x_3335;
assign x_9997 = x_3333 & x_9996;
assign x_9998 = x_3337 & x_3338;
assign x_9999 = x_3336 & x_9998;
assign x_10000 = x_9997 & x_9999;
assign x_10001 = x_3340 & x_3341;
assign x_10002 = x_3339 & x_10001;
assign x_10003 = x_3342 & x_3343;
assign x_10004 = x_3344 & x_3345;
assign x_10005 = x_10003 & x_10004;
assign x_10006 = x_10002 & x_10005;
assign x_10007 = x_10000 & x_10006;
assign x_10008 = x_3347 & x_3348;
assign x_10009 = x_3346 & x_10008;
assign x_10010 = x_3350 & x_3351;
assign x_10011 = x_3349 & x_10010;
assign x_10012 = x_10009 & x_10011;
assign x_10013 = x_3353 & x_3354;
assign x_10014 = x_3352 & x_10013;
assign x_10015 = x_3355 & x_3356;
assign x_10016 = x_3357 & x_3358;
assign x_10017 = x_10015 & x_10016;
assign x_10018 = x_10014 & x_10017;
assign x_10019 = x_10012 & x_10018;
assign x_10020 = x_10007 & x_10019;
assign x_10021 = x_3360 & x_3361;
assign x_10022 = x_3359 & x_10021;
assign x_10023 = x_3363 & x_3364;
assign x_10024 = x_3362 & x_10023;
assign x_10025 = x_10022 & x_10024;
assign x_10026 = x_3366 & x_3367;
assign x_10027 = x_3365 & x_10026;
assign x_10028 = x_3368 & x_3369;
assign x_10029 = x_3370 & x_3371;
assign x_10030 = x_10028 & x_10029;
assign x_10031 = x_10027 & x_10030;
assign x_10032 = x_10025 & x_10031;
assign x_10033 = x_3373 & x_3374;
assign x_10034 = x_3372 & x_10033;
assign x_10035 = x_3376 & x_3377;
assign x_10036 = x_3375 & x_10035;
assign x_10037 = x_10034 & x_10036;
assign x_10038 = x_3379 & x_3380;
assign x_10039 = x_3378 & x_10038;
assign x_10040 = x_3381 & x_3382;
assign x_10041 = x_3383 & x_3384;
assign x_10042 = x_10040 & x_10041;
assign x_10043 = x_10039 & x_10042;
assign x_10044 = x_10037 & x_10043;
assign x_10045 = x_10032 & x_10044;
assign x_10046 = x_10020 & x_10045;
assign x_10047 = x_3386 & x_3387;
assign x_10048 = x_3385 & x_10047;
assign x_10049 = x_3389 & x_3390;
assign x_10050 = x_3388 & x_10049;
assign x_10051 = x_10048 & x_10050;
assign x_10052 = x_3392 & x_3393;
assign x_10053 = x_3391 & x_10052;
assign x_10054 = x_3394 & x_3395;
assign x_10055 = x_3396 & x_3397;
assign x_10056 = x_10054 & x_10055;
assign x_10057 = x_10053 & x_10056;
assign x_10058 = x_10051 & x_10057;
assign x_10059 = x_3399 & x_3400;
assign x_10060 = x_3398 & x_10059;
assign x_10061 = x_3402 & x_3403;
assign x_10062 = x_3401 & x_10061;
assign x_10063 = x_10060 & x_10062;
assign x_10064 = x_3405 & x_3406;
assign x_10065 = x_3404 & x_10064;
assign x_10066 = x_3407 & x_3408;
assign x_10067 = x_3409 & x_3410;
assign x_10068 = x_10066 & x_10067;
assign x_10069 = x_10065 & x_10068;
assign x_10070 = x_10063 & x_10069;
assign x_10071 = x_10058 & x_10070;
assign x_10072 = x_3412 & x_3413;
assign x_10073 = x_3411 & x_10072;
assign x_10074 = x_3415 & x_3416;
assign x_10075 = x_3414 & x_10074;
assign x_10076 = x_10073 & x_10075;
assign x_10077 = x_3418 & x_3419;
assign x_10078 = x_3417 & x_10077;
assign x_10079 = x_3420 & x_3421;
assign x_10080 = x_3422 & x_3423;
assign x_10081 = x_10079 & x_10080;
assign x_10082 = x_10078 & x_10081;
assign x_10083 = x_10076 & x_10082;
assign x_10084 = x_3425 & x_3426;
assign x_10085 = x_3424 & x_10084;
assign x_10086 = x_3428 & x_3429;
assign x_10087 = x_3427 & x_10086;
assign x_10088 = x_10085 & x_10087;
assign x_10089 = x_3431 & x_3432;
assign x_10090 = x_3430 & x_10089;
assign x_10091 = x_3433 & x_3434;
assign x_10092 = x_3435 & x_3436;
assign x_10093 = x_10091 & x_10092;
assign x_10094 = x_10090 & x_10093;
assign x_10095 = x_10088 & x_10094;
assign x_10096 = x_10083 & x_10095;
assign x_10097 = x_10071 & x_10096;
assign x_10098 = x_10046 & x_10097;
assign x_10099 = x_3438 & x_3439;
assign x_10100 = x_3437 & x_10099;
assign x_10101 = x_3441 & x_3442;
assign x_10102 = x_3440 & x_10101;
assign x_10103 = x_10100 & x_10102;
assign x_10104 = x_3444 & x_3445;
assign x_10105 = x_3443 & x_10104;
assign x_10106 = x_3446 & x_3447;
assign x_10107 = x_3448 & x_3449;
assign x_10108 = x_10106 & x_10107;
assign x_10109 = x_10105 & x_10108;
assign x_10110 = x_10103 & x_10109;
assign x_10111 = x_3451 & x_3452;
assign x_10112 = x_3450 & x_10111;
assign x_10113 = x_3454 & x_3455;
assign x_10114 = x_3453 & x_10113;
assign x_10115 = x_10112 & x_10114;
assign x_10116 = x_3457 & x_3458;
assign x_10117 = x_3456 & x_10116;
assign x_10118 = x_3459 & x_3460;
assign x_10119 = x_3461 & x_3462;
assign x_10120 = x_10118 & x_10119;
assign x_10121 = x_10117 & x_10120;
assign x_10122 = x_10115 & x_10121;
assign x_10123 = x_10110 & x_10122;
assign x_10124 = x_3464 & x_3465;
assign x_10125 = x_3463 & x_10124;
assign x_10126 = x_3467 & x_3468;
assign x_10127 = x_3466 & x_10126;
assign x_10128 = x_10125 & x_10127;
assign x_10129 = x_3470 & x_3471;
assign x_10130 = x_3469 & x_10129;
assign x_10131 = x_3472 & x_3473;
assign x_10132 = x_3474 & x_3475;
assign x_10133 = x_10131 & x_10132;
assign x_10134 = x_10130 & x_10133;
assign x_10135 = x_10128 & x_10134;
assign x_10136 = x_3477 & x_3478;
assign x_10137 = x_3476 & x_10136;
assign x_10138 = x_3480 & x_3481;
assign x_10139 = x_3479 & x_10138;
assign x_10140 = x_10137 & x_10139;
assign x_10141 = x_3483 & x_3484;
assign x_10142 = x_3482 & x_10141;
assign x_10143 = x_3485 & x_3486;
assign x_10144 = x_3487 & x_3488;
assign x_10145 = x_10143 & x_10144;
assign x_10146 = x_10142 & x_10145;
assign x_10147 = x_10140 & x_10146;
assign x_10148 = x_10135 & x_10147;
assign x_10149 = x_10123 & x_10148;
assign x_10150 = x_3490 & x_3491;
assign x_10151 = x_3489 & x_10150;
assign x_10152 = x_3493 & x_3494;
assign x_10153 = x_3492 & x_10152;
assign x_10154 = x_10151 & x_10153;
assign x_10155 = x_3496 & x_3497;
assign x_10156 = x_3495 & x_10155;
assign x_10157 = x_3498 & x_3499;
assign x_10158 = x_3500 & x_3501;
assign x_10159 = x_10157 & x_10158;
assign x_10160 = x_10156 & x_10159;
assign x_10161 = x_10154 & x_10160;
assign x_10162 = x_3503 & x_3504;
assign x_10163 = x_3502 & x_10162;
assign x_10164 = x_3506 & x_3507;
assign x_10165 = x_3505 & x_10164;
assign x_10166 = x_10163 & x_10165;
assign x_10167 = x_3509 & x_3510;
assign x_10168 = x_3508 & x_10167;
assign x_10169 = x_3511 & x_3512;
assign x_10170 = x_3513 & x_3514;
assign x_10171 = x_10169 & x_10170;
assign x_10172 = x_10168 & x_10171;
assign x_10173 = x_10166 & x_10172;
assign x_10174 = x_10161 & x_10173;
assign x_10175 = x_3516 & x_3517;
assign x_10176 = x_3515 & x_10175;
assign x_10177 = x_3519 & x_3520;
assign x_10178 = x_3518 & x_10177;
assign x_10179 = x_10176 & x_10178;
assign x_10180 = x_3522 & x_3523;
assign x_10181 = x_3521 & x_10180;
assign x_10182 = x_3524 & x_3525;
assign x_10183 = x_3526 & x_3527;
assign x_10184 = x_10182 & x_10183;
assign x_10185 = x_10181 & x_10184;
assign x_10186 = x_10179 & x_10185;
assign x_10187 = x_3529 & x_3530;
assign x_10188 = x_3528 & x_10187;
assign x_10189 = x_3532 & x_3533;
assign x_10190 = x_3531 & x_10189;
assign x_10191 = x_10188 & x_10190;
assign x_10192 = x_3535 & x_3536;
assign x_10193 = x_3534 & x_10192;
assign x_10194 = x_3537 & x_3538;
assign x_10195 = x_3539 & x_3540;
assign x_10196 = x_10194 & x_10195;
assign x_10197 = x_10193 & x_10196;
assign x_10198 = x_10191 & x_10197;
assign x_10199 = x_10186 & x_10198;
assign x_10200 = x_10174 & x_10199;
assign x_10201 = x_10149 & x_10200;
assign x_10202 = x_10098 & x_10201;
assign x_10203 = x_3542 & x_3543;
assign x_10204 = x_3541 & x_10203;
assign x_10205 = x_3545 & x_3546;
assign x_10206 = x_3544 & x_10205;
assign x_10207 = x_10204 & x_10206;
assign x_10208 = x_3548 & x_3549;
assign x_10209 = x_3547 & x_10208;
assign x_10210 = x_3550 & x_3551;
assign x_10211 = x_3552 & x_3553;
assign x_10212 = x_10210 & x_10211;
assign x_10213 = x_10209 & x_10212;
assign x_10214 = x_10207 & x_10213;
assign x_10215 = x_3555 & x_3556;
assign x_10216 = x_3554 & x_10215;
assign x_10217 = x_3558 & x_3559;
assign x_10218 = x_3557 & x_10217;
assign x_10219 = x_10216 & x_10218;
assign x_10220 = x_3561 & x_3562;
assign x_10221 = x_3560 & x_10220;
assign x_10222 = x_3563 & x_3564;
assign x_10223 = x_3565 & x_3566;
assign x_10224 = x_10222 & x_10223;
assign x_10225 = x_10221 & x_10224;
assign x_10226 = x_10219 & x_10225;
assign x_10227 = x_10214 & x_10226;
assign x_10228 = x_3568 & x_3569;
assign x_10229 = x_3567 & x_10228;
assign x_10230 = x_3571 & x_3572;
assign x_10231 = x_3570 & x_10230;
assign x_10232 = x_10229 & x_10231;
assign x_10233 = x_3574 & x_3575;
assign x_10234 = x_3573 & x_10233;
assign x_10235 = x_3576 & x_3577;
assign x_10236 = x_3578 & x_3579;
assign x_10237 = x_10235 & x_10236;
assign x_10238 = x_10234 & x_10237;
assign x_10239 = x_10232 & x_10238;
assign x_10240 = x_3581 & x_3582;
assign x_10241 = x_3580 & x_10240;
assign x_10242 = x_3584 & x_3585;
assign x_10243 = x_3583 & x_10242;
assign x_10244 = x_10241 & x_10243;
assign x_10245 = x_3587 & x_3588;
assign x_10246 = x_3586 & x_10245;
assign x_10247 = x_3589 & x_3590;
assign x_10248 = x_3591 & x_3592;
assign x_10249 = x_10247 & x_10248;
assign x_10250 = x_10246 & x_10249;
assign x_10251 = x_10244 & x_10250;
assign x_10252 = x_10239 & x_10251;
assign x_10253 = x_10227 & x_10252;
assign x_10254 = x_3594 & x_3595;
assign x_10255 = x_3593 & x_10254;
assign x_10256 = x_3597 & x_3598;
assign x_10257 = x_3596 & x_10256;
assign x_10258 = x_10255 & x_10257;
assign x_10259 = x_3600 & x_3601;
assign x_10260 = x_3599 & x_10259;
assign x_10261 = x_3602 & x_3603;
assign x_10262 = x_3604 & x_3605;
assign x_10263 = x_10261 & x_10262;
assign x_10264 = x_10260 & x_10263;
assign x_10265 = x_10258 & x_10264;
assign x_10266 = x_3607 & x_3608;
assign x_10267 = x_3606 & x_10266;
assign x_10268 = x_3610 & x_3611;
assign x_10269 = x_3609 & x_10268;
assign x_10270 = x_10267 & x_10269;
assign x_10271 = x_3613 & x_3614;
assign x_10272 = x_3612 & x_10271;
assign x_10273 = x_3615 & x_3616;
assign x_10274 = x_3617 & x_3618;
assign x_10275 = x_10273 & x_10274;
assign x_10276 = x_10272 & x_10275;
assign x_10277 = x_10270 & x_10276;
assign x_10278 = x_10265 & x_10277;
assign x_10279 = x_3620 & x_3621;
assign x_10280 = x_3619 & x_10279;
assign x_10281 = x_3623 & x_3624;
assign x_10282 = x_3622 & x_10281;
assign x_10283 = x_10280 & x_10282;
assign x_10284 = x_3626 & x_3627;
assign x_10285 = x_3625 & x_10284;
assign x_10286 = x_3628 & x_3629;
assign x_10287 = x_3630 & x_3631;
assign x_10288 = x_10286 & x_10287;
assign x_10289 = x_10285 & x_10288;
assign x_10290 = x_10283 & x_10289;
assign x_10291 = x_3633 & x_3634;
assign x_10292 = x_3632 & x_10291;
assign x_10293 = x_3636 & x_3637;
assign x_10294 = x_3635 & x_10293;
assign x_10295 = x_10292 & x_10294;
assign x_10296 = x_3639 & x_3640;
assign x_10297 = x_3638 & x_10296;
assign x_10298 = x_3641 & x_3642;
assign x_10299 = x_3643 & x_3644;
assign x_10300 = x_10298 & x_10299;
assign x_10301 = x_10297 & x_10300;
assign x_10302 = x_10295 & x_10301;
assign x_10303 = x_10290 & x_10302;
assign x_10304 = x_10278 & x_10303;
assign x_10305 = x_10253 & x_10304;
assign x_10306 = x_3646 & x_3647;
assign x_10307 = x_3645 & x_10306;
assign x_10308 = x_3649 & x_3650;
assign x_10309 = x_3648 & x_10308;
assign x_10310 = x_10307 & x_10309;
assign x_10311 = x_3652 & x_3653;
assign x_10312 = x_3651 & x_10311;
assign x_10313 = x_3654 & x_3655;
assign x_10314 = x_3656 & x_3657;
assign x_10315 = x_10313 & x_10314;
assign x_10316 = x_10312 & x_10315;
assign x_10317 = x_10310 & x_10316;
assign x_10318 = x_3659 & x_3660;
assign x_10319 = x_3658 & x_10318;
assign x_10320 = x_3662 & x_3663;
assign x_10321 = x_3661 & x_10320;
assign x_10322 = x_10319 & x_10321;
assign x_10323 = x_3665 & x_3666;
assign x_10324 = x_3664 & x_10323;
assign x_10325 = x_3667 & x_3668;
assign x_10326 = x_3669 & x_3670;
assign x_10327 = x_10325 & x_10326;
assign x_10328 = x_10324 & x_10327;
assign x_10329 = x_10322 & x_10328;
assign x_10330 = x_10317 & x_10329;
assign x_10331 = x_3672 & x_3673;
assign x_10332 = x_3671 & x_10331;
assign x_10333 = x_3675 & x_3676;
assign x_10334 = x_3674 & x_10333;
assign x_10335 = x_10332 & x_10334;
assign x_10336 = x_3678 & x_3679;
assign x_10337 = x_3677 & x_10336;
assign x_10338 = x_3680 & x_3681;
assign x_10339 = x_3682 & x_3683;
assign x_10340 = x_10338 & x_10339;
assign x_10341 = x_10337 & x_10340;
assign x_10342 = x_10335 & x_10341;
assign x_10343 = x_3685 & x_3686;
assign x_10344 = x_3684 & x_10343;
assign x_10345 = x_3688 & x_3689;
assign x_10346 = x_3687 & x_10345;
assign x_10347 = x_10344 & x_10346;
assign x_10348 = x_3691 & x_3692;
assign x_10349 = x_3690 & x_10348;
assign x_10350 = x_3693 & x_3694;
assign x_10351 = x_3695 & x_3696;
assign x_10352 = x_10350 & x_10351;
assign x_10353 = x_10349 & x_10352;
assign x_10354 = x_10347 & x_10353;
assign x_10355 = x_10342 & x_10354;
assign x_10356 = x_10330 & x_10355;
assign x_10357 = x_3698 & x_3699;
assign x_10358 = x_3697 & x_10357;
assign x_10359 = x_3701 & x_3702;
assign x_10360 = x_3700 & x_10359;
assign x_10361 = x_10358 & x_10360;
assign x_10362 = x_3704 & x_3705;
assign x_10363 = x_3703 & x_10362;
assign x_10364 = x_3706 & x_3707;
assign x_10365 = x_3708 & x_3709;
assign x_10366 = x_10364 & x_10365;
assign x_10367 = x_10363 & x_10366;
assign x_10368 = x_10361 & x_10367;
assign x_10369 = x_3711 & x_3712;
assign x_10370 = x_3710 & x_10369;
assign x_10371 = x_3714 & x_3715;
assign x_10372 = x_3713 & x_10371;
assign x_10373 = x_10370 & x_10372;
assign x_10374 = x_3717 & x_3718;
assign x_10375 = x_3716 & x_10374;
assign x_10376 = x_3719 & x_3720;
assign x_10377 = x_3721 & x_3722;
assign x_10378 = x_10376 & x_10377;
assign x_10379 = x_10375 & x_10378;
assign x_10380 = x_10373 & x_10379;
assign x_10381 = x_10368 & x_10380;
assign x_10382 = x_3724 & x_3725;
assign x_10383 = x_3723 & x_10382;
assign x_10384 = x_3727 & x_3728;
assign x_10385 = x_3726 & x_10384;
assign x_10386 = x_10383 & x_10385;
assign x_10387 = x_3730 & x_3731;
assign x_10388 = x_3729 & x_10387;
assign x_10389 = x_3732 & x_3733;
assign x_10390 = x_3734 & x_3735;
assign x_10391 = x_10389 & x_10390;
assign x_10392 = x_10388 & x_10391;
assign x_10393 = x_10386 & x_10392;
assign x_10394 = x_3737 & x_3738;
assign x_10395 = x_3736 & x_10394;
assign x_10396 = x_3740 & x_3741;
assign x_10397 = x_3739 & x_10396;
assign x_10398 = x_10395 & x_10397;
assign x_10399 = x_3743 & x_3744;
assign x_10400 = x_3742 & x_10399;
assign x_10401 = x_3745 & x_3746;
assign x_10402 = x_3747 & x_3748;
assign x_10403 = x_10401 & x_10402;
assign x_10404 = x_10400 & x_10403;
assign x_10405 = x_10398 & x_10404;
assign x_10406 = x_10393 & x_10405;
assign x_10407 = x_10381 & x_10406;
assign x_10408 = x_10356 & x_10407;
assign x_10409 = x_10305 & x_10408;
assign x_10410 = x_10202 & x_10409;
assign x_10411 = x_3750 & x_3751;
assign x_10412 = x_3749 & x_10411;
assign x_10413 = x_3753 & x_3754;
assign x_10414 = x_3752 & x_10413;
assign x_10415 = x_10412 & x_10414;
assign x_10416 = x_3756 & x_3757;
assign x_10417 = x_3755 & x_10416;
assign x_10418 = x_3758 & x_3759;
assign x_10419 = x_3760 & x_3761;
assign x_10420 = x_10418 & x_10419;
assign x_10421 = x_10417 & x_10420;
assign x_10422 = x_10415 & x_10421;
assign x_10423 = x_3763 & x_3764;
assign x_10424 = x_3762 & x_10423;
assign x_10425 = x_3766 & x_3767;
assign x_10426 = x_3765 & x_10425;
assign x_10427 = x_10424 & x_10426;
assign x_10428 = x_3769 & x_3770;
assign x_10429 = x_3768 & x_10428;
assign x_10430 = x_3771 & x_3772;
assign x_10431 = x_3773 & x_3774;
assign x_10432 = x_10430 & x_10431;
assign x_10433 = x_10429 & x_10432;
assign x_10434 = x_10427 & x_10433;
assign x_10435 = x_10422 & x_10434;
assign x_10436 = x_3776 & x_3777;
assign x_10437 = x_3775 & x_10436;
assign x_10438 = x_3779 & x_3780;
assign x_10439 = x_3778 & x_10438;
assign x_10440 = x_10437 & x_10439;
assign x_10441 = x_3782 & x_3783;
assign x_10442 = x_3781 & x_10441;
assign x_10443 = x_3784 & x_3785;
assign x_10444 = x_3786 & x_3787;
assign x_10445 = x_10443 & x_10444;
assign x_10446 = x_10442 & x_10445;
assign x_10447 = x_10440 & x_10446;
assign x_10448 = x_3789 & x_3790;
assign x_10449 = x_3788 & x_10448;
assign x_10450 = x_3792 & x_3793;
assign x_10451 = x_3791 & x_10450;
assign x_10452 = x_10449 & x_10451;
assign x_10453 = x_3795 & x_3796;
assign x_10454 = x_3794 & x_10453;
assign x_10455 = x_3797 & x_3798;
assign x_10456 = x_3799 & x_3800;
assign x_10457 = x_10455 & x_10456;
assign x_10458 = x_10454 & x_10457;
assign x_10459 = x_10452 & x_10458;
assign x_10460 = x_10447 & x_10459;
assign x_10461 = x_10435 & x_10460;
assign x_10462 = x_3802 & x_3803;
assign x_10463 = x_3801 & x_10462;
assign x_10464 = x_3805 & x_3806;
assign x_10465 = x_3804 & x_10464;
assign x_10466 = x_10463 & x_10465;
assign x_10467 = x_3808 & x_3809;
assign x_10468 = x_3807 & x_10467;
assign x_10469 = x_3810 & x_3811;
assign x_10470 = x_3812 & x_3813;
assign x_10471 = x_10469 & x_10470;
assign x_10472 = x_10468 & x_10471;
assign x_10473 = x_10466 & x_10472;
assign x_10474 = x_3815 & x_3816;
assign x_10475 = x_3814 & x_10474;
assign x_10476 = x_3818 & x_3819;
assign x_10477 = x_3817 & x_10476;
assign x_10478 = x_10475 & x_10477;
assign x_10479 = x_3821 & x_3822;
assign x_10480 = x_3820 & x_10479;
assign x_10481 = x_3823 & x_3824;
assign x_10482 = x_3825 & x_3826;
assign x_10483 = x_10481 & x_10482;
assign x_10484 = x_10480 & x_10483;
assign x_10485 = x_10478 & x_10484;
assign x_10486 = x_10473 & x_10485;
assign x_10487 = x_3828 & x_3829;
assign x_10488 = x_3827 & x_10487;
assign x_10489 = x_3831 & x_3832;
assign x_10490 = x_3830 & x_10489;
assign x_10491 = x_10488 & x_10490;
assign x_10492 = x_3834 & x_3835;
assign x_10493 = x_3833 & x_10492;
assign x_10494 = x_3836 & x_3837;
assign x_10495 = x_3838 & x_3839;
assign x_10496 = x_10494 & x_10495;
assign x_10497 = x_10493 & x_10496;
assign x_10498 = x_10491 & x_10497;
assign x_10499 = x_3841 & x_3842;
assign x_10500 = x_3840 & x_10499;
assign x_10501 = x_3844 & x_3845;
assign x_10502 = x_3843 & x_10501;
assign x_10503 = x_10500 & x_10502;
assign x_10504 = x_3847 & x_3848;
assign x_10505 = x_3846 & x_10504;
assign x_10506 = x_3849 & x_3850;
assign x_10507 = x_3851 & x_3852;
assign x_10508 = x_10506 & x_10507;
assign x_10509 = x_10505 & x_10508;
assign x_10510 = x_10503 & x_10509;
assign x_10511 = x_10498 & x_10510;
assign x_10512 = x_10486 & x_10511;
assign x_10513 = x_10461 & x_10512;
assign x_10514 = x_3854 & x_3855;
assign x_10515 = x_3853 & x_10514;
assign x_10516 = x_3857 & x_3858;
assign x_10517 = x_3856 & x_10516;
assign x_10518 = x_10515 & x_10517;
assign x_10519 = x_3860 & x_3861;
assign x_10520 = x_3859 & x_10519;
assign x_10521 = x_3862 & x_3863;
assign x_10522 = x_3864 & x_3865;
assign x_10523 = x_10521 & x_10522;
assign x_10524 = x_10520 & x_10523;
assign x_10525 = x_10518 & x_10524;
assign x_10526 = x_3867 & x_3868;
assign x_10527 = x_3866 & x_10526;
assign x_10528 = x_3870 & x_3871;
assign x_10529 = x_3869 & x_10528;
assign x_10530 = x_10527 & x_10529;
assign x_10531 = x_3873 & x_3874;
assign x_10532 = x_3872 & x_10531;
assign x_10533 = x_3875 & x_3876;
assign x_10534 = x_3877 & x_3878;
assign x_10535 = x_10533 & x_10534;
assign x_10536 = x_10532 & x_10535;
assign x_10537 = x_10530 & x_10536;
assign x_10538 = x_10525 & x_10537;
assign x_10539 = x_3880 & x_3881;
assign x_10540 = x_3879 & x_10539;
assign x_10541 = x_3883 & x_3884;
assign x_10542 = x_3882 & x_10541;
assign x_10543 = x_10540 & x_10542;
assign x_10544 = x_3886 & x_3887;
assign x_10545 = x_3885 & x_10544;
assign x_10546 = x_3888 & x_3889;
assign x_10547 = x_3890 & x_3891;
assign x_10548 = x_10546 & x_10547;
assign x_10549 = x_10545 & x_10548;
assign x_10550 = x_10543 & x_10549;
assign x_10551 = x_3893 & x_3894;
assign x_10552 = x_3892 & x_10551;
assign x_10553 = x_3896 & x_3897;
assign x_10554 = x_3895 & x_10553;
assign x_10555 = x_10552 & x_10554;
assign x_10556 = x_3899 & x_3900;
assign x_10557 = x_3898 & x_10556;
assign x_10558 = x_3901 & x_3902;
assign x_10559 = x_3903 & x_3904;
assign x_10560 = x_10558 & x_10559;
assign x_10561 = x_10557 & x_10560;
assign x_10562 = x_10555 & x_10561;
assign x_10563 = x_10550 & x_10562;
assign x_10564 = x_10538 & x_10563;
assign x_10565 = x_3906 & x_3907;
assign x_10566 = x_3905 & x_10565;
assign x_10567 = x_3909 & x_3910;
assign x_10568 = x_3908 & x_10567;
assign x_10569 = x_10566 & x_10568;
assign x_10570 = x_3912 & x_3913;
assign x_10571 = x_3911 & x_10570;
assign x_10572 = x_3914 & x_3915;
assign x_10573 = x_3916 & x_3917;
assign x_10574 = x_10572 & x_10573;
assign x_10575 = x_10571 & x_10574;
assign x_10576 = x_10569 & x_10575;
assign x_10577 = x_3919 & x_3920;
assign x_10578 = x_3918 & x_10577;
assign x_10579 = x_3922 & x_3923;
assign x_10580 = x_3921 & x_10579;
assign x_10581 = x_10578 & x_10580;
assign x_10582 = x_3925 & x_3926;
assign x_10583 = x_3924 & x_10582;
assign x_10584 = x_3927 & x_3928;
assign x_10585 = x_3929 & x_3930;
assign x_10586 = x_10584 & x_10585;
assign x_10587 = x_10583 & x_10586;
assign x_10588 = x_10581 & x_10587;
assign x_10589 = x_10576 & x_10588;
assign x_10590 = x_3932 & x_3933;
assign x_10591 = x_3931 & x_10590;
assign x_10592 = x_3935 & x_3936;
assign x_10593 = x_3934 & x_10592;
assign x_10594 = x_10591 & x_10593;
assign x_10595 = x_3938 & x_3939;
assign x_10596 = x_3937 & x_10595;
assign x_10597 = x_3940 & x_3941;
assign x_10598 = x_3942 & x_3943;
assign x_10599 = x_10597 & x_10598;
assign x_10600 = x_10596 & x_10599;
assign x_10601 = x_10594 & x_10600;
assign x_10602 = x_3945 & x_3946;
assign x_10603 = x_3944 & x_10602;
assign x_10604 = x_3948 & x_3949;
assign x_10605 = x_3947 & x_10604;
assign x_10606 = x_10603 & x_10605;
assign x_10607 = x_3951 & x_3952;
assign x_10608 = x_3950 & x_10607;
assign x_10609 = x_3953 & x_3954;
assign x_10610 = x_3955 & x_3956;
assign x_10611 = x_10609 & x_10610;
assign x_10612 = x_10608 & x_10611;
assign x_10613 = x_10606 & x_10612;
assign x_10614 = x_10601 & x_10613;
assign x_10615 = x_10589 & x_10614;
assign x_10616 = x_10564 & x_10615;
assign x_10617 = x_10513 & x_10616;
assign x_10618 = x_3958 & x_3959;
assign x_10619 = x_3957 & x_10618;
assign x_10620 = x_3961 & x_3962;
assign x_10621 = x_3960 & x_10620;
assign x_10622 = x_10619 & x_10621;
assign x_10623 = x_3964 & x_3965;
assign x_10624 = x_3963 & x_10623;
assign x_10625 = x_3966 & x_3967;
assign x_10626 = x_3968 & x_3969;
assign x_10627 = x_10625 & x_10626;
assign x_10628 = x_10624 & x_10627;
assign x_10629 = x_10622 & x_10628;
assign x_10630 = x_3971 & x_3972;
assign x_10631 = x_3970 & x_10630;
assign x_10632 = x_3974 & x_3975;
assign x_10633 = x_3973 & x_10632;
assign x_10634 = x_10631 & x_10633;
assign x_10635 = x_3977 & x_3978;
assign x_10636 = x_3976 & x_10635;
assign x_10637 = x_3979 & x_3980;
assign x_10638 = x_3981 & x_3982;
assign x_10639 = x_10637 & x_10638;
assign x_10640 = x_10636 & x_10639;
assign x_10641 = x_10634 & x_10640;
assign x_10642 = x_10629 & x_10641;
assign x_10643 = x_3984 & x_3985;
assign x_10644 = x_3983 & x_10643;
assign x_10645 = x_3987 & x_3988;
assign x_10646 = x_3986 & x_10645;
assign x_10647 = x_10644 & x_10646;
assign x_10648 = x_3990 & x_3991;
assign x_10649 = x_3989 & x_10648;
assign x_10650 = x_3992 & x_3993;
assign x_10651 = x_3994 & x_3995;
assign x_10652 = x_10650 & x_10651;
assign x_10653 = x_10649 & x_10652;
assign x_10654 = x_10647 & x_10653;
assign x_10655 = x_3997 & x_3998;
assign x_10656 = x_3996 & x_10655;
assign x_10657 = x_4000 & x_4001;
assign x_10658 = x_3999 & x_10657;
assign x_10659 = x_10656 & x_10658;
assign x_10660 = x_4003 & x_4004;
assign x_10661 = x_4002 & x_10660;
assign x_10662 = x_4005 & x_4006;
assign x_10663 = x_4007 & x_4008;
assign x_10664 = x_10662 & x_10663;
assign x_10665 = x_10661 & x_10664;
assign x_10666 = x_10659 & x_10665;
assign x_10667 = x_10654 & x_10666;
assign x_10668 = x_10642 & x_10667;
assign x_10669 = x_4010 & x_4011;
assign x_10670 = x_4009 & x_10669;
assign x_10671 = x_4013 & x_4014;
assign x_10672 = x_4012 & x_10671;
assign x_10673 = x_10670 & x_10672;
assign x_10674 = x_4016 & x_4017;
assign x_10675 = x_4015 & x_10674;
assign x_10676 = x_4018 & x_4019;
assign x_10677 = x_4020 & x_4021;
assign x_10678 = x_10676 & x_10677;
assign x_10679 = x_10675 & x_10678;
assign x_10680 = x_10673 & x_10679;
assign x_10681 = x_4023 & x_4024;
assign x_10682 = x_4022 & x_10681;
assign x_10683 = x_4026 & x_4027;
assign x_10684 = x_4025 & x_10683;
assign x_10685 = x_10682 & x_10684;
assign x_10686 = x_4029 & x_4030;
assign x_10687 = x_4028 & x_10686;
assign x_10688 = x_4031 & x_4032;
assign x_10689 = x_4033 & x_4034;
assign x_10690 = x_10688 & x_10689;
assign x_10691 = x_10687 & x_10690;
assign x_10692 = x_10685 & x_10691;
assign x_10693 = x_10680 & x_10692;
assign x_10694 = x_4036 & x_4037;
assign x_10695 = x_4035 & x_10694;
assign x_10696 = x_4039 & x_4040;
assign x_10697 = x_4038 & x_10696;
assign x_10698 = x_10695 & x_10697;
assign x_10699 = x_4042 & x_4043;
assign x_10700 = x_4041 & x_10699;
assign x_10701 = x_4044 & x_4045;
assign x_10702 = x_4046 & x_4047;
assign x_10703 = x_10701 & x_10702;
assign x_10704 = x_10700 & x_10703;
assign x_10705 = x_10698 & x_10704;
assign x_10706 = x_4049 & x_4050;
assign x_10707 = x_4048 & x_10706;
assign x_10708 = x_4052 & x_4053;
assign x_10709 = x_4051 & x_10708;
assign x_10710 = x_10707 & x_10709;
assign x_10711 = x_4055 & x_4056;
assign x_10712 = x_4054 & x_10711;
assign x_10713 = x_4057 & x_4058;
assign x_10714 = x_4059 & x_4060;
assign x_10715 = x_10713 & x_10714;
assign x_10716 = x_10712 & x_10715;
assign x_10717 = x_10710 & x_10716;
assign x_10718 = x_10705 & x_10717;
assign x_10719 = x_10693 & x_10718;
assign x_10720 = x_10668 & x_10719;
assign x_10721 = x_4062 & x_4063;
assign x_10722 = x_4061 & x_10721;
assign x_10723 = x_4065 & x_4066;
assign x_10724 = x_4064 & x_10723;
assign x_10725 = x_10722 & x_10724;
assign x_10726 = x_4068 & x_4069;
assign x_10727 = x_4067 & x_10726;
assign x_10728 = x_4070 & x_4071;
assign x_10729 = x_4072 & x_4073;
assign x_10730 = x_10728 & x_10729;
assign x_10731 = x_10727 & x_10730;
assign x_10732 = x_10725 & x_10731;
assign x_10733 = x_4075 & x_4076;
assign x_10734 = x_4074 & x_10733;
assign x_10735 = x_4078 & x_4079;
assign x_10736 = x_4077 & x_10735;
assign x_10737 = x_10734 & x_10736;
assign x_10738 = x_4081 & x_4082;
assign x_10739 = x_4080 & x_10738;
assign x_10740 = x_4083 & x_4084;
assign x_10741 = x_4085 & x_4086;
assign x_10742 = x_10740 & x_10741;
assign x_10743 = x_10739 & x_10742;
assign x_10744 = x_10737 & x_10743;
assign x_10745 = x_10732 & x_10744;
assign x_10746 = x_4088 & x_4089;
assign x_10747 = x_4087 & x_10746;
assign x_10748 = x_4091 & x_4092;
assign x_10749 = x_4090 & x_10748;
assign x_10750 = x_10747 & x_10749;
assign x_10751 = x_4094 & x_4095;
assign x_10752 = x_4093 & x_10751;
assign x_10753 = x_4096 & x_4097;
assign x_10754 = x_4098 & x_4099;
assign x_10755 = x_10753 & x_10754;
assign x_10756 = x_10752 & x_10755;
assign x_10757 = x_10750 & x_10756;
assign x_10758 = x_4101 & x_4102;
assign x_10759 = x_4100 & x_10758;
assign x_10760 = x_4104 & x_4105;
assign x_10761 = x_4103 & x_10760;
assign x_10762 = x_10759 & x_10761;
assign x_10763 = x_4107 & x_4108;
assign x_10764 = x_4106 & x_10763;
assign x_10765 = x_4109 & x_4110;
assign x_10766 = x_4111 & x_4112;
assign x_10767 = x_10765 & x_10766;
assign x_10768 = x_10764 & x_10767;
assign x_10769 = x_10762 & x_10768;
assign x_10770 = x_10757 & x_10769;
assign x_10771 = x_10745 & x_10770;
assign x_10772 = x_4114 & x_4115;
assign x_10773 = x_4113 & x_10772;
assign x_10774 = x_4117 & x_4118;
assign x_10775 = x_4116 & x_10774;
assign x_10776 = x_10773 & x_10775;
assign x_10777 = x_4120 & x_4121;
assign x_10778 = x_4119 & x_10777;
assign x_10779 = x_4122 & x_4123;
assign x_10780 = x_4124 & x_4125;
assign x_10781 = x_10779 & x_10780;
assign x_10782 = x_10778 & x_10781;
assign x_10783 = x_10776 & x_10782;
assign x_10784 = x_4127 & x_4128;
assign x_10785 = x_4126 & x_10784;
assign x_10786 = x_4130 & x_4131;
assign x_10787 = x_4129 & x_10786;
assign x_10788 = x_10785 & x_10787;
assign x_10789 = x_4133 & x_4134;
assign x_10790 = x_4132 & x_10789;
assign x_10791 = x_4135 & x_4136;
assign x_10792 = x_4137 & x_4138;
assign x_10793 = x_10791 & x_10792;
assign x_10794 = x_10790 & x_10793;
assign x_10795 = x_10788 & x_10794;
assign x_10796 = x_10783 & x_10795;
assign x_10797 = x_4140 & x_4141;
assign x_10798 = x_4139 & x_10797;
assign x_10799 = x_4143 & x_4144;
assign x_10800 = x_4142 & x_10799;
assign x_10801 = x_10798 & x_10800;
assign x_10802 = x_4146 & x_4147;
assign x_10803 = x_4145 & x_10802;
assign x_10804 = x_4148 & x_4149;
assign x_10805 = x_4150 & x_4151;
assign x_10806 = x_10804 & x_10805;
assign x_10807 = x_10803 & x_10806;
assign x_10808 = x_10801 & x_10807;
assign x_10809 = x_4153 & x_4154;
assign x_10810 = x_4152 & x_10809;
assign x_10811 = x_4155 & x_4156;
assign x_10812 = x_4157 & x_4158;
assign x_10813 = x_10811 & x_10812;
assign x_10814 = x_10810 & x_10813;
assign x_10815 = x_4160 & x_4161;
assign x_10816 = x_4159 & x_10815;
assign x_10817 = x_4162 & x_4163;
assign x_10818 = x_4164 & x_4165;
assign x_10819 = x_10817 & x_10818;
assign x_10820 = x_10816 & x_10819;
assign x_10821 = x_10814 & x_10820;
assign x_10822 = x_10808 & x_10821;
assign x_10823 = x_10796 & x_10822;
assign x_10824 = x_10771 & x_10823;
assign x_10825 = x_10720 & x_10824;
assign x_10826 = x_10617 & x_10825;
assign x_10827 = x_10410 & x_10826;
assign x_10828 = x_4167 & x_4168;
assign x_10829 = x_4166 & x_10828;
assign x_10830 = x_4170 & x_4171;
assign x_10831 = x_4169 & x_10830;
assign x_10832 = x_10829 & x_10831;
assign x_10833 = x_4173 & x_4174;
assign x_10834 = x_4172 & x_10833;
assign x_10835 = x_4175 & x_4176;
assign x_10836 = x_4177 & x_4178;
assign x_10837 = x_10835 & x_10836;
assign x_10838 = x_10834 & x_10837;
assign x_10839 = x_10832 & x_10838;
assign x_10840 = x_4180 & x_4181;
assign x_10841 = x_4179 & x_10840;
assign x_10842 = x_4183 & x_4184;
assign x_10843 = x_4182 & x_10842;
assign x_10844 = x_10841 & x_10843;
assign x_10845 = x_4186 & x_4187;
assign x_10846 = x_4185 & x_10845;
assign x_10847 = x_4188 & x_4189;
assign x_10848 = x_4190 & x_4191;
assign x_10849 = x_10847 & x_10848;
assign x_10850 = x_10846 & x_10849;
assign x_10851 = x_10844 & x_10850;
assign x_10852 = x_10839 & x_10851;
assign x_10853 = x_4193 & x_4194;
assign x_10854 = x_4192 & x_10853;
assign x_10855 = x_4196 & x_4197;
assign x_10856 = x_4195 & x_10855;
assign x_10857 = x_10854 & x_10856;
assign x_10858 = x_4199 & x_4200;
assign x_10859 = x_4198 & x_10858;
assign x_10860 = x_4201 & x_4202;
assign x_10861 = x_4203 & x_4204;
assign x_10862 = x_10860 & x_10861;
assign x_10863 = x_10859 & x_10862;
assign x_10864 = x_10857 & x_10863;
assign x_10865 = x_4206 & x_4207;
assign x_10866 = x_4205 & x_10865;
assign x_10867 = x_4209 & x_4210;
assign x_10868 = x_4208 & x_10867;
assign x_10869 = x_10866 & x_10868;
assign x_10870 = x_4212 & x_4213;
assign x_10871 = x_4211 & x_10870;
assign x_10872 = x_4214 & x_4215;
assign x_10873 = x_4216 & x_4217;
assign x_10874 = x_10872 & x_10873;
assign x_10875 = x_10871 & x_10874;
assign x_10876 = x_10869 & x_10875;
assign x_10877 = x_10864 & x_10876;
assign x_10878 = x_10852 & x_10877;
assign x_10879 = x_4219 & x_4220;
assign x_10880 = x_4218 & x_10879;
assign x_10881 = x_4222 & x_4223;
assign x_10882 = x_4221 & x_10881;
assign x_10883 = x_10880 & x_10882;
assign x_10884 = x_4225 & x_4226;
assign x_10885 = x_4224 & x_10884;
assign x_10886 = x_4227 & x_4228;
assign x_10887 = x_4229 & x_4230;
assign x_10888 = x_10886 & x_10887;
assign x_10889 = x_10885 & x_10888;
assign x_10890 = x_10883 & x_10889;
assign x_10891 = x_4232 & x_4233;
assign x_10892 = x_4231 & x_10891;
assign x_10893 = x_4235 & x_4236;
assign x_10894 = x_4234 & x_10893;
assign x_10895 = x_10892 & x_10894;
assign x_10896 = x_4238 & x_4239;
assign x_10897 = x_4237 & x_10896;
assign x_10898 = x_4240 & x_4241;
assign x_10899 = x_4242 & x_4243;
assign x_10900 = x_10898 & x_10899;
assign x_10901 = x_10897 & x_10900;
assign x_10902 = x_10895 & x_10901;
assign x_10903 = x_10890 & x_10902;
assign x_10904 = x_4245 & x_4246;
assign x_10905 = x_4244 & x_10904;
assign x_10906 = x_4248 & x_4249;
assign x_10907 = x_4247 & x_10906;
assign x_10908 = x_10905 & x_10907;
assign x_10909 = x_4251 & x_4252;
assign x_10910 = x_4250 & x_10909;
assign x_10911 = x_4253 & x_4254;
assign x_10912 = x_4255 & x_4256;
assign x_10913 = x_10911 & x_10912;
assign x_10914 = x_10910 & x_10913;
assign x_10915 = x_10908 & x_10914;
assign x_10916 = x_4258 & x_4259;
assign x_10917 = x_4257 & x_10916;
assign x_10918 = x_4261 & x_4262;
assign x_10919 = x_4260 & x_10918;
assign x_10920 = x_10917 & x_10919;
assign x_10921 = x_4264 & x_4265;
assign x_10922 = x_4263 & x_10921;
assign x_10923 = x_4266 & x_4267;
assign x_10924 = x_4268 & x_4269;
assign x_10925 = x_10923 & x_10924;
assign x_10926 = x_10922 & x_10925;
assign x_10927 = x_10920 & x_10926;
assign x_10928 = x_10915 & x_10927;
assign x_10929 = x_10903 & x_10928;
assign x_10930 = x_10878 & x_10929;
assign x_10931 = x_4271 & x_4272;
assign x_10932 = x_4270 & x_10931;
assign x_10933 = x_4274 & x_4275;
assign x_10934 = x_4273 & x_10933;
assign x_10935 = x_10932 & x_10934;
assign x_10936 = x_4277 & x_4278;
assign x_10937 = x_4276 & x_10936;
assign x_10938 = x_4279 & x_4280;
assign x_10939 = x_4281 & x_4282;
assign x_10940 = x_10938 & x_10939;
assign x_10941 = x_10937 & x_10940;
assign x_10942 = x_10935 & x_10941;
assign x_10943 = x_4284 & x_4285;
assign x_10944 = x_4283 & x_10943;
assign x_10945 = x_4287 & x_4288;
assign x_10946 = x_4286 & x_10945;
assign x_10947 = x_10944 & x_10946;
assign x_10948 = x_4290 & x_4291;
assign x_10949 = x_4289 & x_10948;
assign x_10950 = x_4292 & x_4293;
assign x_10951 = x_4294 & x_4295;
assign x_10952 = x_10950 & x_10951;
assign x_10953 = x_10949 & x_10952;
assign x_10954 = x_10947 & x_10953;
assign x_10955 = x_10942 & x_10954;
assign x_10956 = x_4297 & x_4298;
assign x_10957 = x_4296 & x_10956;
assign x_10958 = x_4300 & x_4301;
assign x_10959 = x_4299 & x_10958;
assign x_10960 = x_10957 & x_10959;
assign x_10961 = x_4303 & x_4304;
assign x_10962 = x_4302 & x_10961;
assign x_10963 = x_4305 & x_4306;
assign x_10964 = x_4307 & x_4308;
assign x_10965 = x_10963 & x_10964;
assign x_10966 = x_10962 & x_10965;
assign x_10967 = x_10960 & x_10966;
assign x_10968 = x_4310 & x_4311;
assign x_10969 = x_4309 & x_10968;
assign x_10970 = x_4313 & x_4314;
assign x_10971 = x_4312 & x_10970;
assign x_10972 = x_10969 & x_10971;
assign x_10973 = x_4316 & x_4317;
assign x_10974 = x_4315 & x_10973;
assign x_10975 = x_4318 & x_4319;
assign x_10976 = x_4320 & x_4321;
assign x_10977 = x_10975 & x_10976;
assign x_10978 = x_10974 & x_10977;
assign x_10979 = x_10972 & x_10978;
assign x_10980 = x_10967 & x_10979;
assign x_10981 = x_10955 & x_10980;
assign x_10982 = x_4323 & x_4324;
assign x_10983 = x_4322 & x_10982;
assign x_10984 = x_4326 & x_4327;
assign x_10985 = x_4325 & x_10984;
assign x_10986 = x_10983 & x_10985;
assign x_10987 = x_4329 & x_4330;
assign x_10988 = x_4328 & x_10987;
assign x_10989 = x_4331 & x_4332;
assign x_10990 = x_4333 & x_4334;
assign x_10991 = x_10989 & x_10990;
assign x_10992 = x_10988 & x_10991;
assign x_10993 = x_10986 & x_10992;
assign x_10994 = x_4336 & x_4337;
assign x_10995 = x_4335 & x_10994;
assign x_10996 = x_4339 & x_4340;
assign x_10997 = x_4338 & x_10996;
assign x_10998 = x_10995 & x_10997;
assign x_10999 = x_4342 & x_4343;
assign x_11000 = x_4341 & x_10999;
assign x_11001 = x_4344 & x_4345;
assign x_11002 = x_4346 & x_4347;
assign x_11003 = x_11001 & x_11002;
assign x_11004 = x_11000 & x_11003;
assign x_11005 = x_10998 & x_11004;
assign x_11006 = x_10993 & x_11005;
assign x_11007 = x_4349 & x_4350;
assign x_11008 = x_4348 & x_11007;
assign x_11009 = x_4352 & x_4353;
assign x_11010 = x_4351 & x_11009;
assign x_11011 = x_11008 & x_11010;
assign x_11012 = x_4355 & x_4356;
assign x_11013 = x_4354 & x_11012;
assign x_11014 = x_4357 & x_4358;
assign x_11015 = x_4359 & x_4360;
assign x_11016 = x_11014 & x_11015;
assign x_11017 = x_11013 & x_11016;
assign x_11018 = x_11011 & x_11017;
assign x_11019 = x_4362 & x_4363;
assign x_11020 = x_4361 & x_11019;
assign x_11021 = x_4365 & x_4366;
assign x_11022 = x_4364 & x_11021;
assign x_11023 = x_11020 & x_11022;
assign x_11024 = x_4368 & x_4369;
assign x_11025 = x_4367 & x_11024;
assign x_11026 = x_4370 & x_4371;
assign x_11027 = x_4372 & x_4373;
assign x_11028 = x_11026 & x_11027;
assign x_11029 = x_11025 & x_11028;
assign x_11030 = x_11023 & x_11029;
assign x_11031 = x_11018 & x_11030;
assign x_11032 = x_11006 & x_11031;
assign x_11033 = x_10981 & x_11032;
assign x_11034 = x_10930 & x_11033;
assign x_11035 = x_4375 & x_4376;
assign x_11036 = x_4374 & x_11035;
assign x_11037 = x_4378 & x_4379;
assign x_11038 = x_4377 & x_11037;
assign x_11039 = x_11036 & x_11038;
assign x_11040 = x_4381 & x_4382;
assign x_11041 = x_4380 & x_11040;
assign x_11042 = x_4383 & x_4384;
assign x_11043 = x_4385 & x_4386;
assign x_11044 = x_11042 & x_11043;
assign x_11045 = x_11041 & x_11044;
assign x_11046 = x_11039 & x_11045;
assign x_11047 = x_4388 & x_4389;
assign x_11048 = x_4387 & x_11047;
assign x_11049 = x_4391 & x_4392;
assign x_11050 = x_4390 & x_11049;
assign x_11051 = x_11048 & x_11050;
assign x_11052 = x_4394 & x_4395;
assign x_11053 = x_4393 & x_11052;
assign x_11054 = x_4396 & x_4397;
assign x_11055 = x_4398 & x_4399;
assign x_11056 = x_11054 & x_11055;
assign x_11057 = x_11053 & x_11056;
assign x_11058 = x_11051 & x_11057;
assign x_11059 = x_11046 & x_11058;
assign x_11060 = x_4401 & x_4402;
assign x_11061 = x_4400 & x_11060;
assign x_11062 = x_4404 & x_4405;
assign x_11063 = x_4403 & x_11062;
assign x_11064 = x_11061 & x_11063;
assign x_11065 = x_4407 & x_4408;
assign x_11066 = x_4406 & x_11065;
assign x_11067 = x_4409 & x_4410;
assign x_11068 = x_4411 & x_4412;
assign x_11069 = x_11067 & x_11068;
assign x_11070 = x_11066 & x_11069;
assign x_11071 = x_11064 & x_11070;
assign x_11072 = x_4414 & x_4415;
assign x_11073 = x_4413 & x_11072;
assign x_11074 = x_4417 & x_4418;
assign x_11075 = x_4416 & x_11074;
assign x_11076 = x_11073 & x_11075;
assign x_11077 = x_4420 & x_4421;
assign x_11078 = x_4419 & x_11077;
assign x_11079 = x_4422 & x_4423;
assign x_11080 = x_4424 & x_4425;
assign x_11081 = x_11079 & x_11080;
assign x_11082 = x_11078 & x_11081;
assign x_11083 = x_11076 & x_11082;
assign x_11084 = x_11071 & x_11083;
assign x_11085 = x_11059 & x_11084;
assign x_11086 = x_4427 & x_4428;
assign x_11087 = x_4426 & x_11086;
assign x_11088 = x_4430 & x_4431;
assign x_11089 = x_4429 & x_11088;
assign x_11090 = x_11087 & x_11089;
assign x_11091 = x_4433 & x_4434;
assign x_11092 = x_4432 & x_11091;
assign x_11093 = x_4435 & x_4436;
assign x_11094 = x_4437 & x_4438;
assign x_11095 = x_11093 & x_11094;
assign x_11096 = x_11092 & x_11095;
assign x_11097 = x_11090 & x_11096;
assign x_11098 = x_4440 & x_4441;
assign x_11099 = x_4439 & x_11098;
assign x_11100 = x_4443 & x_4444;
assign x_11101 = x_4442 & x_11100;
assign x_11102 = x_11099 & x_11101;
assign x_11103 = x_4446 & x_4447;
assign x_11104 = x_4445 & x_11103;
assign x_11105 = x_4448 & x_4449;
assign x_11106 = x_4450 & x_4451;
assign x_11107 = x_11105 & x_11106;
assign x_11108 = x_11104 & x_11107;
assign x_11109 = x_11102 & x_11108;
assign x_11110 = x_11097 & x_11109;
assign x_11111 = x_4453 & x_4454;
assign x_11112 = x_4452 & x_11111;
assign x_11113 = x_4456 & x_4457;
assign x_11114 = x_4455 & x_11113;
assign x_11115 = x_11112 & x_11114;
assign x_11116 = x_4459 & x_4460;
assign x_11117 = x_4458 & x_11116;
assign x_11118 = x_4461 & x_4462;
assign x_11119 = x_4463 & x_4464;
assign x_11120 = x_11118 & x_11119;
assign x_11121 = x_11117 & x_11120;
assign x_11122 = x_11115 & x_11121;
assign x_11123 = x_4466 & x_4467;
assign x_11124 = x_4465 & x_11123;
assign x_11125 = x_4469 & x_4470;
assign x_11126 = x_4468 & x_11125;
assign x_11127 = x_11124 & x_11126;
assign x_11128 = x_4472 & x_4473;
assign x_11129 = x_4471 & x_11128;
assign x_11130 = x_4474 & x_4475;
assign x_11131 = x_4476 & x_4477;
assign x_11132 = x_11130 & x_11131;
assign x_11133 = x_11129 & x_11132;
assign x_11134 = x_11127 & x_11133;
assign x_11135 = x_11122 & x_11134;
assign x_11136 = x_11110 & x_11135;
assign x_11137 = x_11085 & x_11136;
assign x_11138 = x_4479 & x_4480;
assign x_11139 = x_4478 & x_11138;
assign x_11140 = x_4482 & x_4483;
assign x_11141 = x_4481 & x_11140;
assign x_11142 = x_11139 & x_11141;
assign x_11143 = x_4485 & x_4486;
assign x_11144 = x_4484 & x_11143;
assign x_11145 = x_4487 & x_4488;
assign x_11146 = x_4489 & x_4490;
assign x_11147 = x_11145 & x_11146;
assign x_11148 = x_11144 & x_11147;
assign x_11149 = x_11142 & x_11148;
assign x_11150 = x_4492 & x_4493;
assign x_11151 = x_4491 & x_11150;
assign x_11152 = x_4495 & x_4496;
assign x_11153 = x_4494 & x_11152;
assign x_11154 = x_11151 & x_11153;
assign x_11155 = x_4498 & x_4499;
assign x_11156 = x_4497 & x_11155;
assign x_11157 = x_4500 & x_4501;
assign x_11158 = x_4502 & x_4503;
assign x_11159 = x_11157 & x_11158;
assign x_11160 = x_11156 & x_11159;
assign x_11161 = x_11154 & x_11160;
assign x_11162 = x_11149 & x_11161;
assign x_11163 = x_4505 & x_4506;
assign x_11164 = x_4504 & x_11163;
assign x_11165 = x_4508 & x_4509;
assign x_11166 = x_4507 & x_11165;
assign x_11167 = x_11164 & x_11166;
assign x_11168 = x_4511 & x_4512;
assign x_11169 = x_4510 & x_11168;
assign x_11170 = x_4513 & x_4514;
assign x_11171 = x_4515 & x_4516;
assign x_11172 = x_11170 & x_11171;
assign x_11173 = x_11169 & x_11172;
assign x_11174 = x_11167 & x_11173;
assign x_11175 = x_4518 & x_4519;
assign x_11176 = x_4517 & x_11175;
assign x_11177 = x_4521 & x_4522;
assign x_11178 = x_4520 & x_11177;
assign x_11179 = x_11176 & x_11178;
assign x_11180 = x_4524 & x_4525;
assign x_11181 = x_4523 & x_11180;
assign x_11182 = x_4526 & x_4527;
assign x_11183 = x_4528 & x_4529;
assign x_11184 = x_11182 & x_11183;
assign x_11185 = x_11181 & x_11184;
assign x_11186 = x_11179 & x_11185;
assign x_11187 = x_11174 & x_11186;
assign x_11188 = x_11162 & x_11187;
assign x_11189 = x_4531 & x_4532;
assign x_11190 = x_4530 & x_11189;
assign x_11191 = x_4534 & x_4535;
assign x_11192 = x_4533 & x_11191;
assign x_11193 = x_11190 & x_11192;
assign x_11194 = x_4537 & x_4538;
assign x_11195 = x_4536 & x_11194;
assign x_11196 = x_4539 & x_4540;
assign x_11197 = x_4541 & x_4542;
assign x_11198 = x_11196 & x_11197;
assign x_11199 = x_11195 & x_11198;
assign x_11200 = x_11193 & x_11199;
assign x_11201 = x_4544 & x_4545;
assign x_11202 = x_4543 & x_11201;
assign x_11203 = x_4547 & x_4548;
assign x_11204 = x_4546 & x_11203;
assign x_11205 = x_11202 & x_11204;
assign x_11206 = x_4550 & x_4551;
assign x_11207 = x_4549 & x_11206;
assign x_11208 = x_4552 & x_4553;
assign x_11209 = x_4554 & x_4555;
assign x_11210 = x_11208 & x_11209;
assign x_11211 = x_11207 & x_11210;
assign x_11212 = x_11205 & x_11211;
assign x_11213 = x_11200 & x_11212;
assign x_11214 = x_4557 & x_4558;
assign x_11215 = x_4556 & x_11214;
assign x_11216 = x_4560 & x_4561;
assign x_11217 = x_4559 & x_11216;
assign x_11218 = x_11215 & x_11217;
assign x_11219 = x_4563 & x_4564;
assign x_11220 = x_4562 & x_11219;
assign x_11221 = x_4565 & x_4566;
assign x_11222 = x_4567 & x_4568;
assign x_11223 = x_11221 & x_11222;
assign x_11224 = x_11220 & x_11223;
assign x_11225 = x_11218 & x_11224;
assign x_11226 = x_4570 & x_4571;
assign x_11227 = x_4569 & x_11226;
assign x_11228 = x_4573 & x_4574;
assign x_11229 = x_4572 & x_11228;
assign x_11230 = x_11227 & x_11229;
assign x_11231 = x_4576 & x_4577;
assign x_11232 = x_4575 & x_11231;
assign x_11233 = x_4578 & x_4579;
assign x_11234 = x_4580 & x_4581;
assign x_11235 = x_11233 & x_11234;
assign x_11236 = x_11232 & x_11235;
assign x_11237 = x_11230 & x_11236;
assign x_11238 = x_11225 & x_11237;
assign x_11239 = x_11213 & x_11238;
assign x_11240 = x_11188 & x_11239;
assign x_11241 = x_11137 & x_11240;
assign x_11242 = x_11034 & x_11241;
assign x_11243 = x_4583 & x_4584;
assign x_11244 = x_4582 & x_11243;
assign x_11245 = x_4586 & x_4587;
assign x_11246 = x_4585 & x_11245;
assign x_11247 = x_11244 & x_11246;
assign x_11248 = x_4589 & x_4590;
assign x_11249 = x_4588 & x_11248;
assign x_11250 = x_4591 & x_4592;
assign x_11251 = x_4593 & x_4594;
assign x_11252 = x_11250 & x_11251;
assign x_11253 = x_11249 & x_11252;
assign x_11254 = x_11247 & x_11253;
assign x_11255 = x_4596 & x_4597;
assign x_11256 = x_4595 & x_11255;
assign x_11257 = x_4599 & x_4600;
assign x_11258 = x_4598 & x_11257;
assign x_11259 = x_11256 & x_11258;
assign x_11260 = x_4602 & x_4603;
assign x_11261 = x_4601 & x_11260;
assign x_11262 = x_4604 & x_4605;
assign x_11263 = x_4606 & x_4607;
assign x_11264 = x_11262 & x_11263;
assign x_11265 = x_11261 & x_11264;
assign x_11266 = x_11259 & x_11265;
assign x_11267 = x_11254 & x_11266;
assign x_11268 = x_4609 & x_4610;
assign x_11269 = x_4608 & x_11268;
assign x_11270 = x_4612 & x_4613;
assign x_11271 = x_4611 & x_11270;
assign x_11272 = x_11269 & x_11271;
assign x_11273 = x_4615 & x_4616;
assign x_11274 = x_4614 & x_11273;
assign x_11275 = x_4617 & x_4618;
assign x_11276 = x_4619 & x_4620;
assign x_11277 = x_11275 & x_11276;
assign x_11278 = x_11274 & x_11277;
assign x_11279 = x_11272 & x_11278;
assign x_11280 = x_4622 & x_4623;
assign x_11281 = x_4621 & x_11280;
assign x_11282 = x_4625 & x_4626;
assign x_11283 = x_4624 & x_11282;
assign x_11284 = x_11281 & x_11283;
assign x_11285 = x_4628 & x_4629;
assign x_11286 = x_4627 & x_11285;
assign x_11287 = x_4630 & x_4631;
assign x_11288 = x_4632 & x_4633;
assign x_11289 = x_11287 & x_11288;
assign x_11290 = x_11286 & x_11289;
assign x_11291 = x_11284 & x_11290;
assign x_11292 = x_11279 & x_11291;
assign x_11293 = x_11267 & x_11292;
assign x_11294 = x_4635 & x_4636;
assign x_11295 = x_4634 & x_11294;
assign x_11296 = x_4638 & x_4639;
assign x_11297 = x_4637 & x_11296;
assign x_11298 = x_11295 & x_11297;
assign x_11299 = x_4641 & x_4642;
assign x_11300 = x_4640 & x_11299;
assign x_11301 = x_4643 & x_4644;
assign x_11302 = x_4645 & x_4646;
assign x_11303 = x_11301 & x_11302;
assign x_11304 = x_11300 & x_11303;
assign x_11305 = x_11298 & x_11304;
assign x_11306 = x_4648 & x_4649;
assign x_11307 = x_4647 & x_11306;
assign x_11308 = x_4651 & x_4652;
assign x_11309 = x_4650 & x_11308;
assign x_11310 = x_11307 & x_11309;
assign x_11311 = x_4654 & x_4655;
assign x_11312 = x_4653 & x_11311;
assign x_11313 = x_4656 & x_4657;
assign x_11314 = x_4658 & x_4659;
assign x_11315 = x_11313 & x_11314;
assign x_11316 = x_11312 & x_11315;
assign x_11317 = x_11310 & x_11316;
assign x_11318 = x_11305 & x_11317;
assign x_11319 = x_4661 & x_4662;
assign x_11320 = x_4660 & x_11319;
assign x_11321 = x_4664 & x_4665;
assign x_11322 = x_4663 & x_11321;
assign x_11323 = x_11320 & x_11322;
assign x_11324 = x_4667 & x_4668;
assign x_11325 = x_4666 & x_11324;
assign x_11326 = x_4669 & x_4670;
assign x_11327 = x_4671 & x_4672;
assign x_11328 = x_11326 & x_11327;
assign x_11329 = x_11325 & x_11328;
assign x_11330 = x_11323 & x_11329;
assign x_11331 = x_4674 & x_4675;
assign x_11332 = x_4673 & x_11331;
assign x_11333 = x_4677 & x_4678;
assign x_11334 = x_4676 & x_11333;
assign x_11335 = x_11332 & x_11334;
assign x_11336 = x_4680 & x_4681;
assign x_11337 = x_4679 & x_11336;
assign x_11338 = x_4682 & x_4683;
assign x_11339 = x_4684 & x_4685;
assign x_11340 = x_11338 & x_11339;
assign x_11341 = x_11337 & x_11340;
assign x_11342 = x_11335 & x_11341;
assign x_11343 = x_11330 & x_11342;
assign x_11344 = x_11318 & x_11343;
assign x_11345 = x_11293 & x_11344;
assign x_11346 = x_4687 & x_4688;
assign x_11347 = x_4686 & x_11346;
assign x_11348 = x_4690 & x_4691;
assign x_11349 = x_4689 & x_11348;
assign x_11350 = x_11347 & x_11349;
assign x_11351 = x_4693 & x_4694;
assign x_11352 = x_4692 & x_11351;
assign x_11353 = x_4695 & x_4696;
assign x_11354 = x_4697 & x_4698;
assign x_11355 = x_11353 & x_11354;
assign x_11356 = x_11352 & x_11355;
assign x_11357 = x_11350 & x_11356;
assign x_11358 = x_4700 & x_4701;
assign x_11359 = x_4699 & x_11358;
assign x_11360 = x_4703 & x_4704;
assign x_11361 = x_4702 & x_11360;
assign x_11362 = x_11359 & x_11361;
assign x_11363 = x_4706 & x_4707;
assign x_11364 = x_4705 & x_11363;
assign x_11365 = x_4708 & x_4709;
assign x_11366 = x_4710 & x_4711;
assign x_11367 = x_11365 & x_11366;
assign x_11368 = x_11364 & x_11367;
assign x_11369 = x_11362 & x_11368;
assign x_11370 = x_11357 & x_11369;
assign x_11371 = x_4713 & x_4714;
assign x_11372 = x_4712 & x_11371;
assign x_11373 = x_4716 & x_4717;
assign x_11374 = x_4715 & x_11373;
assign x_11375 = x_11372 & x_11374;
assign x_11376 = x_4719 & x_4720;
assign x_11377 = x_4718 & x_11376;
assign x_11378 = x_4721 & x_4722;
assign x_11379 = x_4723 & x_4724;
assign x_11380 = x_11378 & x_11379;
assign x_11381 = x_11377 & x_11380;
assign x_11382 = x_11375 & x_11381;
assign x_11383 = x_4726 & x_4727;
assign x_11384 = x_4725 & x_11383;
assign x_11385 = x_4729 & x_4730;
assign x_11386 = x_4728 & x_11385;
assign x_11387 = x_11384 & x_11386;
assign x_11388 = x_4732 & x_4733;
assign x_11389 = x_4731 & x_11388;
assign x_11390 = x_4734 & x_4735;
assign x_11391 = x_4736 & x_4737;
assign x_11392 = x_11390 & x_11391;
assign x_11393 = x_11389 & x_11392;
assign x_11394 = x_11387 & x_11393;
assign x_11395 = x_11382 & x_11394;
assign x_11396 = x_11370 & x_11395;
assign x_11397 = x_4739 & x_4740;
assign x_11398 = x_4738 & x_11397;
assign x_11399 = x_4742 & x_4743;
assign x_11400 = x_4741 & x_11399;
assign x_11401 = x_11398 & x_11400;
assign x_11402 = x_4745 & x_4746;
assign x_11403 = x_4744 & x_11402;
assign x_11404 = x_4747 & x_4748;
assign x_11405 = x_4749 & x_4750;
assign x_11406 = x_11404 & x_11405;
assign x_11407 = x_11403 & x_11406;
assign x_11408 = x_11401 & x_11407;
assign x_11409 = x_4752 & x_4753;
assign x_11410 = x_4751 & x_11409;
assign x_11411 = x_4755 & x_4756;
assign x_11412 = x_4754 & x_11411;
assign x_11413 = x_11410 & x_11412;
assign x_11414 = x_4758 & x_4759;
assign x_11415 = x_4757 & x_11414;
assign x_11416 = x_4760 & x_4761;
assign x_11417 = x_4762 & x_4763;
assign x_11418 = x_11416 & x_11417;
assign x_11419 = x_11415 & x_11418;
assign x_11420 = x_11413 & x_11419;
assign x_11421 = x_11408 & x_11420;
assign x_11422 = x_4765 & x_4766;
assign x_11423 = x_4764 & x_11422;
assign x_11424 = x_4768 & x_4769;
assign x_11425 = x_4767 & x_11424;
assign x_11426 = x_11423 & x_11425;
assign x_11427 = x_4771 & x_4772;
assign x_11428 = x_4770 & x_11427;
assign x_11429 = x_4773 & x_4774;
assign x_11430 = x_4775 & x_4776;
assign x_11431 = x_11429 & x_11430;
assign x_11432 = x_11428 & x_11431;
assign x_11433 = x_11426 & x_11432;
assign x_11434 = x_4778 & x_4779;
assign x_11435 = x_4777 & x_11434;
assign x_11436 = x_4781 & x_4782;
assign x_11437 = x_4780 & x_11436;
assign x_11438 = x_11435 & x_11437;
assign x_11439 = x_4784 & x_4785;
assign x_11440 = x_4783 & x_11439;
assign x_11441 = x_4786 & x_4787;
assign x_11442 = x_4788 & x_4789;
assign x_11443 = x_11441 & x_11442;
assign x_11444 = x_11440 & x_11443;
assign x_11445 = x_11438 & x_11444;
assign x_11446 = x_11433 & x_11445;
assign x_11447 = x_11421 & x_11446;
assign x_11448 = x_11396 & x_11447;
assign x_11449 = x_11345 & x_11448;
assign x_11450 = x_4791 & x_4792;
assign x_11451 = x_4790 & x_11450;
assign x_11452 = x_4794 & x_4795;
assign x_11453 = x_4793 & x_11452;
assign x_11454 = x_11451 & x_11453;
assign x_11455 = x_4797 & x_4798;
assign x_11456 = x_4796 & x_11455;
assign x_11457 = x_4799 & x_4800;
assign x_11458 = x_4801 & x_4802;
assign x_11459 = x_11457 & x_11458;
assign x_11460 = x_11456 & x_11459;
assign x_11461 = x_11454 & x_11460;
assign x_11462 = x_4804 & x_4805;
assign x_11463 = x_4803 & x_11462;
assign x_11464 = x_4807 & x_4808;
assign x_11465 = x_4806 & x_11464;
assign x_11466 = x_11463 & x_11465;
assign x_11467 = x_4810 & x_4811;
assign x_11468 = x_4809 & x_11467;
assign x_11469 = x_4812 & x_4813;
assign x_11470 = x_4814 & x_4815;
assign x_11471 = x_11469 & x_11470;
assign x_11472 = x_11468 & x_11471;
assign x_11473 = x_11466 & x_11472;
assign x_11474 = x_11461 & x_11473;
assign x_11475 = x_4817 & x_4818;
assign x_11476 = x_4816 & x_11475;
assign x_11477 = x_4820 & x_4821;
assign x_11478 = x_4819 & x_11477;
assign x_11479 = x_11476 & x_11478;
assign x_11480 = x_4823 & x_4824;
assign x_11481 = x_4822 & x_11480;
assign x_11482 = x_4825 & x_4826;
assign x_11483 = x_4827 & x_4828;
assign x_11484 = x_11482 & x_11483;
assign x_11485 = x_11481 & x_11484;
assign x_11486 = x_11479 & x_11485;
assign x_11487 = x_4830 & x_4831;
assign x_11488 = x_4829 & x_11487;
assign x_11489 = x_4833 & x_4834;
assign x_11490 = x_4832 & x_11489;
assign x_11491 = x_11488 & x_11490;
assign x_11492 = x_4836 & x_4837;
assign x_11493 = x_4835 & x_11492;
assign x_11494 = x_4838 & x_4839;
assign x_11495 = x_4840 & x_4841;
assign x_11496 = x_11494 & x_11495;
assign x_11497 = x_11493 & x_11496;
assign x_11498 = x_11491 & x_11497;
assign x_11499 = x_11486 & x_11498;
assign x_11500 = x_11474 & x_11499;
assign x_11501 = x_4843 & x_4844;
assign x_11502 = x_4842 & x_11501;
assign x_11503 = x_4846 & x_4847;
assign x_11504 = x_4845 & x_11503;
assign x_11505 = x_11502 & x_11504;
assign x_11506 = x_4849 & x_4850;
assign x_11507 = x_4848 & x_11506;
assign x_11508 = x_4851 & x_4852;
assign x_11509 = x_4853 & x_4854;
assign x_11510 = x_11508 & x_11509;
assign x_11511 = x_11507 & x_11510;
assign x_11512 = x_11505 & x_11511;
assign x_11513 = x_4856 & x_4857;
assign x_11514 = x_4855 & x_11513;
assign x_11515 = x_4859 & x_4860;
assign x_11516 = x_4858 & x_11515;
assign x_11517 = x_11514 & x_11516;
assign x_11518 = x_4862 & x_4863;
assign x_11519 = x_4861 & x_11518;
assign x_11520 = x_4864 & x_4865;
assign x_11521 = x_4866 & x_4867;
assign x_11522 = x_11520 & x_11521;
assign x_11523 = x_11519 & x_11522;
assign x_11524 = x_11517 & x_11523;
assign x_11525 = x_11512 & x_11524;
assign x_11526 = x_4869 & x_4870;
assign x_11527 = x_4868 & x_11526;
assign x_11528 = x_4872 & x_4873;
assign x_11529 = x_4871 & x_11528;
assign x_11530 = x_11527 & x_11529;
assign x_11531 = x_4875 & x_4876;
assign x_11532 = x_4874 & x_11531;
assign x_11533 = x_4877 & x_4878;
assign x_11534 = x_4879 & x_4880;
assign x_11535 = x_11533 & x_11534;
assign x_11536 = x_11532 & x_11535;
assign x_11537 = x_11530 & x_11536;
assign x_11538 = x_4882 & x_4883;
assign x_11539 = x_4881 & x_11538;
assign x_11540 = x_4885 & x_4886;
assign x_11541 = x_4884 & x_11540;
assign x_11542 = x_11539 & x_11541;
assign x_11543 = x_4888 & x_4889;
assign x_11544 = x_4887 & x_11543;
assign x_11545 = x_4890 & x_4891;
assign x_11546 = x_4892 & x_4893;
assign x_11547 = x_11545 & x_11546;
assign x_11548 = x_11544 & x_11547;
assign x_11549 = x_11542 & x_11548;
assign x_11550 = x_11537 & x_11549;
assign x_11551 = x_11525 & x_11550;
assign x_11552 = x_11500 & x_11551;
assign x_11553 = x_4895 & x_4896;
assign x_11554 = x_4894 & x_11553;
assign x_11555 = x_4898 & x_4899;
assign x_11556 = x_4897 & x_11555;
assign x_11557 = x_11554 & x_11556;
assign x_11558 = x_4901 & x_4902;
assign x_11559 = x_4900 & x_11558;
assign x_11560 = x_4903 & x_4904;
assign x_11561 = x_4905 & x_4906;
assign x_11562 = x_11560 & x_11561;
assign x_11563 = x_11559 & x_11562;
assign x_11564 = x_11557 & x_11563;
assign x_11565 = x_4908 & x_4909;
assign x_11566 = x_4907 & x_11565;
assign x_11567 = x_4911 & x_4912;
assign x_11568 = x_4910 & x_11567;
assign x_11569 = x_11566 & x_11568;
assign x_11570 = x_4914 & x_4915;
assign x_11571 = x_4913 & x_11570;
assign x_11572 = x_4916 & x_4917;
assign x_11573 = x_4918 & x_4919;
assign x_11574 = x_11572 & x_11573;
assign x_11575 = x_11571 & x_11574;
assign x_11576 = x_11569 & x_11575;
assign x_11577 = x_11564 & x_11576;
assign x_11578 = x_4921 & x_4922;
assign x_11579 = x_4920 & x_11578;
assign x_11580 = x_4924 & x_4925;
assign x_11581 = x_4923 & x_11580;
assign x_11582 = x_11579 & x_11581;
assign x_11583 = x_4927 & x_4928;
assign x_11584 = x_4926 & x_11583;
assign x_11585 = x_4929 & x_4930;
assign x_11586 = x_4931 & x_4932;
assign x_11587 = x_11585 & x_11586;
assign x_11588 = x_11584 & x_11587;
assign x_11589 = x_11582 & x_11588;
assign x_11590 = x_4934 & x_4935;
assign x_11591 = x_4933 & x_11590;
assign x_11592 = x_4937 & x_4938;
assign x_11593 = x_4936 & x_11592;
assign x_11594 = x_11591 & x_11593;
assign x_11595 = x_4940 & x_4941;
assign x_11596 = x_4939 & x_11595;
assign x_11597 = x_4942 & x_4943;
assign x_11598 = x_4944 & x_4945;
assign x_11599 = x_11597 & x_11598;
assign x_11600 = x_11596 & x_11599;
assign x_11601 = x_11594 & x_11600;
assign x_11602 = x_11589 & x_11601;
assign x_11603 = x_11577 & x_11602;
assign x_11604 = x_4947 & x_4948;
assign x_11605 = x_4946 & x_11604;
assign x_11606 = x_4950 & x_4951;
assign x_11607 = x_4949 & x_11606;
assign x_11608 = x_11605 & x_11607;
assign x_11609 = x_4953 & x_4954;
assign x_11610 = x_4952 & x_11609;
assign x_11611 = x_4955 & x_4956;
assign x_11612 = x_4957 & x_4958;
assign x_11613 = x_11611 & x_11612;
assign x_11614 = x_11610 & x_11613;
assign x_11615 = x_11608 & x_11614;
assign x_11616 = x_4960 & x_4961;
assign x_11617 = x_4959 & x_11616;
assign x_11618 = x_4963 & x_4964;
assign x_11619 = x_4962 & x_11618;
assign x_11620 = x_11617 & x_11619;
assign x_11621 = x_4966 & x_4967;
assign x_11622 = x_4965 & x_11621;
assign x_11623 = x_4968 & x_4969;
assign x_11624 = x_4970 & x_4971;
assign x_11625 = x_11623 & x_11624;
assign x_11626 = x_11622 & x_11625;
assign x_11627 = x_11620 & x_11626;
assign x_11628 = x_11615 & x_11627;
assign x_11629 = x_4973 & x_4974;
assign x_11630 = x_4972 & x_11629;
assign x_11631 = x_4976 & x_4977;
assign x_11632 = x_4975 & x_11631;
assign x_11633 = x_11630 & x_11632;
assign x_11634 = x_4979 & x_4980;
assign x_11635 = x_4978 & x_11634;
assign x_11636 = x_4981 & x_4982;
assign x_11637 = x_4983 & x_4984;
assign x_11638 = x_11636 & x_11637;
assign x_11639 = x_11635 & x_11638;
assign x_11640 = x_11633 & x_11639;
assign x_11641 = x_4986 & x_4987;
assign x_11642 = x_4985 & x_11641;
assign x_11643 = x_4988 & x_4989;
assign x_11644 = x_4990 & x_4991;
assign x_11645 = x_11643 & x_11644;
assign x_11646 = x_11642 & x_11645;
assign x_11647 = x_4993 & x_4994;
assign x_11648 = x_4992 & x_11647;
assign x_11649 = x_4995 & x_4996;
assign x_11650 = x_4997 & x_4998;
assign x_11651 = x_11649 & x_11650;
assign x_11652 = x_11648 & x_11651;
assign x_11653 = x_11646 & x_11652;
assign x_11654 = x_11640 & x_11653;
assign x_11655 = x_11628 & x_11654;
assign x_11656 = x_11603 & x_11655;
assign x_11657 = x_11552 & x_11656;
assign x_11658 = x_11449 & x_11657;
assign x_11659 = x_11242 & x_11658;
assign x_11660 = x_10827 & x_11659;
assign x_11661 = x_5000 & x_5001;
assign x_11662 = x_4999 & x_11661;
assign x_11663 = x_5003 & x_5004;
assign x_11664 = x_5002 & x_11663;
assign x_11665 = x_11662 & x_11664;
assign x_11666 = x_5006 & x_5007;
assign x_11667 = x_5005 & x_11666;
assign x_11668 = x_5008 & x_5009;
assign x_11669 = x_5010 & x_5011;
assign x_11670 = x_11668 & x_11669;
assign x_11671 = x_11667 & x_11670;
assign x_11672 = x_11665 & x_11671;
assign x_11673 = x_5013 & x_5014;
assign x_11674 = x_5012 & x_11673;
assign x_11675 = x_5016 & x_5017;
assign x_11676 = x_5015 & x_11675;
assign x_11677 = x_11674 & x_11676;
assign x_11678 = x_5019 & x_5020;
assign x_11679 = x_5018 & x_11678;
assign x_11680 = x_5021 & x_5022;
assign x_11681 = x_5023 & x_5024;
assign x_11682 = x_11680 & x_11681;
assign x_11683 = x_11679 & x_11682;
assign x_11684 = x_11677 & x_11683;
assign x_11685 = x_11672 & x_11684;
assign x_11686 = x_5026 & x_5027;
assign x_11687 = x_5025 & x_11686;
assign x_11688 = x_5029 & x_5030;
assign x_11689 = x_5028 & x_11688;
assign x_11690 = x_11687 & x_11689;
assign x_11691 = x_5032 & x_5033;
assign x_11692 = x_5031 & x_11691;
assign x_11693 = x_5034 & x_5035;
assign x_11694 = x_5036 & x_5037;
assign x_11695 = x_11693 & x_11694;
assign x_11696 = x_11692 & x_11695;
assign x_11697 = x_11690 & x_11696;
assign x_11698 = x_5039 & x_5040;
assign x_11699 = x_5038 & x_11698;
assign x_11700 = x_5042 & x_5043;
assign x_11701 = x_5041 & x_11700;
assign x_11702 = x_11699 & x_11701;
assign x_11703 = x_5045 & x_5046;
assign x_11704 = x_5044 & x_11703;
assign x_11705 = x_5047 & x_5048;
assign x_11706 = x_5049 & x_5050;
assign x_11707 = x_11705 & x_11706;
assign x_11708 = x_11704 & x_11707;
assign x_11709 = x_11702 & x_11708;
assign x_11710 = x_11697 & x_11709;
assign x_11711 = x_11685 & x_11710;
assign x_11712 = x_5052 & x_5053;
assign x_11713 = x_5051 & x_11712;
assign x_11714 = x_5055 & x_5056;
assign x_11715 = x_5054 & x_11714;
assign x_11716 = x_11713 & x_11715;
assign x_11717 = x_5058 & x_5059;
assign x_11718 = x_5057 & x_11717;
assign x_11719 = x_5060 & x_5061;
assign x_11720 = x_5062 & x_5063;
assign x_11721 = x_11719 & x_11720;
assign x_11722 = x_11718 & x_11721;
assign x_11723 = x_11716 & x_11722;
assign x_11724 = x_5065 & x_5066;
assign x_11725 = x_5064 & x_11724;
assign x_11726 = x_5068 & x_5069;
assign x_11727 = x_5067 & x_11726;
assign x_11728 = x_11725 & x_11727;
assign x_11729 = x_5071 & x_5072;
assign x_11730 = x_5070 & x_11729;
assign x_11731 = x_5073 & x_5074;
assign x_11732 = x_5075 & x_5076;
assign x_11733 = x_11731 & x_11732;
assign x_11734 = x_11730 & x_11733;
assign x_11735 = x_11728 & x_11734;
assign x_11736 = x_11723 & x_11735;
assign x_11737 = x_5078 & x_5079;
assign x_11738 = x_5077 & x_11737;
assign x_11739 = x_5081 & x_5082;
assign x_11740 = x_5080 & x_11739;
assign x_11741 = x_11738 & x_11740;
assign x_11742 = x_5084 & x_5085;
assign x_11743 = x_5083 & x_11742;
assign x_11744 = x_5086 & x_5087;
assign x_11745 = x_5088 & x_5089;
assign x_11746 = x_11744 & x_11745;
assign x_11747 = x_11743 & x_11746;
assign x_11748 = x_11741 & x_11747;
assign x_11749 = x_5091 & x_5092;
assign x_11750 = x_5090 & x_11749;
assign x_11751 = x_5094 & x_5095;
assign x_11752 = x_5093 & x_11751;
assign x_11753 = x_11750 & x_11752;
assign x_11754 = x_5097 & x_5098;
assign x_11755 = x_5096 & x_11754;
assign x_11756 = x_5099 & x_5100;
assign x_11757 = x_5101 & x_5102;
assign x_11758 = x_11756 & x_11757;
assign x_11759 = x_11755 & x_11758;
assign x_11760 = x_11753 & x_11759;
assign x_11761 = x_11748 & x_11760;
assign x_11762 = x_11736 & x_11761;
assign x_11763 = x_11711 & x_11762;
assign x_11764 = x_5104 & x_5105;
assign x_11765 = x_5103 & x_11764;
assign x_11766 = x_5107 & x_5108;
assign x_11767 = x_5106 & x_11766;
assign x_11768 = x_11765 & x_11767;
assign x_11769 = x_5110 & x_5111;
assign x_11770 = x_5109 & x_11769;
assign x_11771 = x_5112 & x_5113;
assign x_11772 = x_5114 & x_5115;
assign x_11773 = x_11771 & x_11772;
assign x_11774 = x_11770 & x_11773;
assign x_11775 = x_11768 & x_11774;
assign x_11776 = x_5117 & x_5118;
assign x_11777 = x_5116 & x_11776;
assign x_11778 = x_5120 & x_5121;
assign x_11779 = x_5119 & x_11778;
assign x_11780 = x_11777 & x_11779;
assign x_11781 = x_5123 & x_5124;
assign x_11782 = x_5122 & x_11781;
assign x_11783 = x_5125 & x_5126;
assign x_11784 = x_5127 & x_5128;
assign x_11785 = x_11783 & x_11784;
assign x_11786 = x_11782 & x_11785;
assign x_11787 = x_11780 & x_11786;
assign x_11788 = x_11775 & x_11787;
assign x_11789 = x_5130 & x_5131;
assign x_11790 = x_5129 & x_11789;
assign x_11791 = x_5133 & x_5134;
assign x_11792 = x_5132 & x_11791;
assign x_11793 = x_11790 & x_11792;
assign x_11794 = x_5136 & x_5137;
assign x_11795 = x_5135 & x_11794;
assign x_11796 = x_5138 & x_5139;
assign x_11797 = x_5140 & x_5141;
assign x_11798 = x_11796 & x_11797;
assign x_11799 = x_11795 & x_11798;
assign x_11800 = x_11793 & x_11799;
assign x_11801 = x_5143 & x_5144;
assign x_11802 = x_5142 & x_11801;
assign x_11803 = x_5146 & x_5147;
assign x_11804 = x_5145 & x_11803;
assign x_11805 = x_11802 & x_11804;
assign x_11806 = x_5149 & x_5150;
assign x_11807 = x_5148 & x_11806;
assign x_11808 = x_5151 & x_5152;
assign x_11809 = x_5153 & x_5154;
assign x_11810 = x_11808 & x_11809;
assign x_11811 = x_11807 & x_11810;
assign x_11812 = x_11805 & x_11811;
assign x_11813 = x_11800 & x_11812;
assign x_11814 = x_11788 & x_11813;
assign x_11815 = x_5156 & x_5157;
assign x_11816 = x_5155 & x_11815;
assign x_11817 = x_5159 & x_5160;
assign x_11818 = x_5158 & x_11817;
assign x_11819 = x_11816 & x_11818;
assign x_11820 = x_5162 & x_5163;
assign x_11821 = x_5161 & x_11820;
assign x_11822 = x_5164 & x_5165;
assign x_11823 = x_5166 & x_5167;
assign x_11824 = x_11822 & x_11823;
assign x_11825 = x_11821 & x_11824;
assign x_11826 = x_11819 & x_11825;
assign x_11827 = x_5169 & x_5170;
assign x_11828 = x_5168 & x_11827;
assign x_11829 = x_5172 & x_5173;
assign x_11830 = x_5171 & x_11829;
assign x_11831 = x_11828 & x_11830;
assign x_11832 = x_5175 & x_5176;
assign x_11833 = x_5174 & x_11832;
assign x_11834 = x_5177 & x_5178;
assign x_11835 = x_5179 & x_5180;
assign x_11836 = x_11834 & x_11835;
assign x_11837 = x_11833 & x_11836;
assign x_11838 = x_11831 & x_11837;
assign x_11839 = x_11826 & x_11838;
assign x_11840 = x_5182 & x_5183;
assign x_11841 = x_5181 & x_11840;
assign x_11842 = x_5185 & x_5186;
assign x_11843 = x_5184 & x_11842;
assign x_11844 = x_11841 & x_11843;
assign x_11845 = x_5188 & x_5189;
assign x_11846 = x_5187 & x_11845;
assign x_11847 = x_5190 & x_5191;
assign x_11848 = x_5192 & x_5193;
assign x_11849 = x_11847 & x_11848;
assign x_11850 = x_11846 & x_11849;
assign x_11851 = x_11844 & x_11850;
assign x_11852 = x_5195 & x_5196;
assign x_11853 = x_5194 & x_11852;
assign x_11854 = x_5198 & x_5199;
assign x_11855 = x_5197 & x_11854;
assign x_11856 = x_11853 & x_11855;
assign x_11857 = x_5201 & x_5202;
assign x_11858 = x_5200 & x_11857;
assign x_11859 = x_5203 & x_5204;
assign x_11860 = x_5205 & x_5206;
assign x_11861 = x_11859 & x_11860;
assign x_11862 = x_11858 & x_11861;
assign x_11863 = x_11856 & x_11862;
assign x_11864 = x_11851 & x_11863;
assign x_11865 = x_11839 & x_11864;
assign x_11866 = x_11814 & x_11865;
assign x_11867 = x_11763 & x_11866;
assign x_11868 = x_5208 & x_5209;
assign x_11869 = x_5207 & x_11868;
assign x_11870 = x_5211 & x_5212;
assign x_11871 = x_5210 & x_11870;
assign x_11872 = x_11869 & x_11871;
assign x_11873 = x_5214 & x_5215;
assign x_11874 = x_5213 & x_11873;
assign x_11875 = x_5216 & x_5217;
assign x_11876 = x_5218 & x_5219;
assign x_11877 = x_11875 & x_11876;
assign x_11878 = x_11874 & x_11877;
assign x_11879 = x_11872 & x_11878;
assign x_11880 = x_5221 & x_5222;
assign x_11881 = x_5220 & x_11880;
assign x_11882 = x_5224 & x_5225;
assign x_11883 = x_5223 & x_11882;
assign x_11884 = x_11881 & x_11883;
assign x_11885 = x_5227 & x_5228;
assign x_11886 = x_5226 & x_11885;
assign x_11887 = x_5229 & x_5230;
assign x_11888 = x_5231 & x_5232;
assign x_11889 = x_11887 & x_11888;
assign x_11890 = x_11886 & x_11889;
assign x_11891 = x_11884 & x_11890;
assign x_11892 = x_11879 & x_11891;
assign x_11893 = x_5234 & x_5235;
assign x_11894 = x_5233 & x_11893;
assign x_11895 = x_5237 & x_5238;
assign x_11896 = x_5236 & x_11895;
assign x_11897 = x_11894 & x_11896;
assign x_11898 = x_5240 & x_5241;
assign x_11899 = x_5239 & x_11898;
assign x_11900 = x_5242 & x_5243;
assign x_11901 = x_5244 & x_5245;
assign x_11902 = x_11900 & x_11901;
assign x_11903 = x_11899 & x_11902;
assign x_11904 = x_11897 & x_11903;
assign x_11905 = x_5247 & x_5248;
assign x_11906 = x_5246 & x_11905;
assign x_11907 = x_5250 & x_5251;
assign x_11908 = x_5249 & x_11907;
assign x_11909 = x_11906 & x_11908;
assign x_11910 = x_5253 & x_5254;
assign x_11911 = x_5252 & x_11910;
assign x_11912 = x_5255 & x_5256;
assign x_11913 = x_5257 & x_5258;
assign x_11914 = x_11912 & x_11913;
assign x_11915 = x_11911 & x_11914;
assign x_11916 = x_11909 & x_11915;
assign x_11917 = x_11904 & x_11916;
assign x_11918 = x_11892 & x_11917;
assign x_11919 = x_5260 & x_5261;
assign x_11920 = x_5259 & x_11919;
assign x_11921 = x_5263 & x_5264;
assign x_11922 = x_5262 & x_11921;
assign x_11923 = x_11920 & x_11922;
assign x_11924 = x_5266 & x_5267;
assign x_11925 = x_5265 & x_11924;
assign x_11926 = x_5268 & x_5269;
assign x_11927 = x_5270 & x_5271;
assign x_11928 = x_11926 & x_11927;
assign x_11929 = x_11925 & x_11928;
assign x_11930 = x_11923 & x_11929;
assign x_11931 = x_5273 & x_5274;
assign x_11932 = x_5272 & x_11931;
assign x_11933 = x_5276 & x_5277;
assign x_11934 = x_5275 & x_11933;
assign x_11935 = x_11932 & x_11934;
assign x_11936 = x_5279 & x_5280;
assign x_11937 = x_5278 & x_11936;
assign x_11938 = x_5281 & x_5282;
assign x_11939 = x_5283 & x_5284;
assign x_11940 = x_11938 & x_11939;
assign x_11941 = x_11937 & x_11940;
assign x_11942 = x_11935 & x_11941;
assign x_11943 = x_11930 & x_11942;
assign x_11944 = x_5286 & x_5287;
assign x_11945 = x_5285 & x_11944;
assign x_11946 = x_5289 & x_5290;
assign x_11947 = x_5288 & x_11946;
assign x_11948 = x_11945 & x_11947;
assign x_11949 = x_5292 & x_5293;
assign x_11950 = x_5291 & x_11949;
assign x_11951 = x_5294 & x_5295;
assign x_11952 = x_5296 & x_5297;
assign x_11953 = x_11951 & x_11952;
assign x_11954 = x_11950 & x_11953;
assign x_11955 = x_11948 & x_11954;
assign x_11956 = x_5299 & x_5300;
assign x_11957 = x_5298 & x_11956;
assign x_11958 = x_5302 & x_5303;
assign x_11959 = x_5301 & x_11958;
assign x_11960 = x_11957 & x_11959;
assign x_11961 = x_5305 & x_5306;
assign x_11962 = x_5304 & x_11961;
assign x_11963 = x_5307 & x_5308;
assign x_11964 = x_5309 & x_5310;
assign x_11965 = x_11963 & x_11964;
assign x_11966 = x_11962 & x_11965;
assign x_11967 = x_11960 & x_11966;
assign x_11968 = x_11955 & x_11967;
assign x_11969 = x_11943 & x_11968;
assign x_11970 = x_11918 & x_11969;
assign x_11971 = x_5312 & x_5313;
assign x_11972 = x_5311 & x_11971;
assign x_11973 = x_5315 & x_5316;
assign x_11974 = x_5314 & x_11973;
assign x_11975 = x_11972 & x_11974;
assign x_11976 = x_5318 & x_5319;
assign x_11977 = x_5317 & x_11976;
assign x_11978 = x_5320 & x_5321;
assign x_11979 = x_5322 & x_5323;
assign x_11980 = x_11978 & x_11979;
assign x_11981 = x_11977 & x_11980;
assign x_11982 = x_11975 & x_11981;
assign x_11983 = x_5325 & x_5326;
assign x_11984 = x_5324 & x_11983;
assign x_11985 = x_5328 & x_5329;
assign x_11986 = x_5327 & x_11985;
assign x_11987 = x_11984 & x_11986;
assign x_11988 = x_5331 & x_5332;
assign x_11989 = x_5330 & x_11988;
assign x_11990 = x_5333 & x_5334;
assign x_11991 = x_5335 & x_5336;
assign x_11992 = x_11990 & x_11991;
assign x_11993 = x_11989 & x_11992;
assign x_11994 = x_11987 & x_11993;
assign x_11995 = x_11982 & x_11994;
assign x_11996 = x_5338 & x_5339;
assign x_11997 = x_5337 & x_11996;
assign x_11998 = x_5341 & x_5342;
assign x_11999 = x_5340 & x_11998;
assign x_12000 = x_11997 & x_11999;
assign x_12001 = x_5344 & x_5345;
assign x_12002 = x_5343 & x_12001;
assign x_12003 = x_5346 & x_5347;
assign x_12004 = x_5348 & x_5349;
assign x_12005 = x_12003 & x_12004;
assign x_12006 = x_12002 & x_12005;
assign x_12007 = x_12000 & x_12006;
assign x_12008 = x_5351 & x_5352;
assign x_12009 = x_5350 & x_12008;
assign x_12010 = x_5354 & x_5355;
assign x_12011 = x_5353 & x_12010;
assign x_12012 = x_12009 & x_12011;
assign x_12013 = x_5357 & x_5358;
assign x_12014 = x_5356 & x_12013;
assign x_12015 = x_5359 & x_5360;
assign x_12016 = x_5361 & x_5362;
assign x_12017 = x_12015 & x_12016;
assign x_12018 = x_12014 & x_12017;
assign x_12019 = x_12012 & x_12018;
assign x_12020 = x_12007 & x_12019;
assign x_12021 = x_11995 & x_12020;
assign x_12022 = x_5364 & x_5365;
assign x_12023 = x_5363 & x_12022;
assign x_12024 = x_5367 & x_5368;
assign x_12025 = x_5366 & x_12024;
assign x_12026 = x_12023 & x_12025;
assign x_12027 = x_5370 & x_5371;
assign x_12028 = x_5369 & x_12027;
assign x_12029 = x_5372 & x_5373;
assign x_12030 = x_5374 & x_5375;
assign x_12031 = x_12029 & x_12030;
assign x_12032 = x_12028 & x_12031;
assign x_12033 = x_12026 & x_12032;
assign x_12034 = x_5377 & x_5378;
assign x_12035 = x_5376 & x_12034;
assign x_12036 = x_5380 & x_5381;
assign x_12037 = x_5379 & x_12036;
assign x_12038 = x_12035 & x_12037;
assign x_12039 = x_5383 & x_5384;
assign x_12040 = x_5382 & x_12039;
assign x_12041 = x_5385 & x_5386;
assign x_12042 = x_5387 & x_5388;
assign x_12043 = x_12041 & x_12042;
assign x_12044 = x_12040 & x_12043;
assign x_12045 = x_12038 & x_12044;
assign x_12046 = x_12033 & x_12045;
assign x_12047 = x_5390 & x_5391;
assign x_12048 = x_5389 & x_12047;
assign x_12049 = x_5393 & x_5394;
assign x_12050 = x_5392 & x_12049;
assign x_12051 = x_12048 & x_12050;
assign x_12052 = x_5396 & x_5397;
assign x_12053 = x_5395 & x_12052;
assign x_12054 = x_5398 & x_5399;
assign x_12055 = x_5400 & x_5401;
assign x_12056 = x_12054 & x_12055;
assign x_12057 = x_12053 & x_12056;
assign x_12058 = x_12051 & x_12057;
assign x_12059 = x_5403 & x_5404;
assign x_12060 = x_5402 & x_12059;
assign x_12061 = x_5406 & x_5407;
assign x_12062 = x_5405 & x_12061;
assign x_12063 = x_12060 & x_12062;
assign x_12064 = x_5409 & x_5410;
assign x_12065 = x_5408 & x_12064;
assign x_12066 = x_5411 & x_5412;
assign x_12067 = x_5413 & x_5414;
assign x_12068 = x_12066 & x_12067;
assign x_12069 = x_12065 & x_12068;
assign x_12070 = x_12063 & x_12069;
assign x_12071 = x_12058 & x_12070;
assign x_12072 = x_12046 & x_12071;
assign x_12073 = x_12021 & x_12072;
assign x_12074 = x_11970 & x_12073;
assign x_12075 = x_11867 & x_12074;
assign x_12076 = x_5416 & x_5417;
assign x_12077 = x_5415 & x_12076;
assign x_12078 = x_5419 & x_5420;
assign x_12079 = x_5418 & x_12078;
assign x_12080 = x_12077 & x_12079;
assign x_12081 = x_5422 & x_5423;
assign x_12082 = x_5421 & x_12081;
assign x_12083 = x_5424 & x_5425;
assign x_12084 = x_5426 & x_5427;
assign x_12085 = x_12083 & x_12084;
assign x_12086 = x_12082 & x_12085;
assign x_12087 = x_12080 & x_12086;
assign x_12088 = x_5429 & x_5430;
assign x_12089 = x_5428 & x_12088;
assign x_12090 = x_5432 & x_5433;
assign x_12091 = x_5431 & x_12090;
assign x_12092 = x_12089 & x_12091;
assign x_12093 = x_5435 & x_5436;
assign x_12094 = x_5434 & x_12093;
assign x_12095 = x_5437 & x_5438;
assign x_12096 = x_5439 & x_5440;
assign x_12097 = x_12095 & x_12096;
assign x_12098 = x_12094 & x_12097;
assign x_12099 = x_12092 & x_12098;
assign x_12100 = x_12087 & x_12099;
assign x_12101 = x_5442 & x_5443;
assign x_12102 = x_5441 & x_12101;
assign x_12103 = x_5445 & x_5446;
assign x_12104 = x_5444 & x_12103;
assign x_12105 = x_12102 & x_12104;
assign x_12106 = x_5448 & x_5449;
assign x_12107 = x_5447 & x_12106;
assign x_12108 = x_5450 & x_5451;
assign x_12109 = x_5452 & x_5453;
assign x_12110 = x_12108 & x_12109;
assign x_12111 = x_12107 & x_12110;
assign x_12112 = x_12105 & x_12111;
assign x_12113 = x_5455 & x_5456;
assign x_12114 = x_5454 & x_12113;
assign x_12115 = x_5458 & x_5459;
assign x_12116 = x_5457 & x_12115;
assign x_12117 = x_12114 & x_12116;
assign x_12118 = x_5461 & x_5462;
assign x_12119 = x_5460 & x_12118;
assign x_12120 = x_5463 & x_5464;
assign x_12121 = x_5465 & x_5466;
assign x_12122 = x_12120 & x_12121;
assign x_12123 = x_12119 & x_12122;
assign x_12124 = x_12117 & x_12123;
assign x_12125 = x_12112 & x_12124;
assign x_12126 = x_12100 & x_12125;
assign x_12127 = x_5468 & x_5469;
assign x_12128 = x_5467 & x_12127;
assign x_12129 = x_5471 & x_5472;
assign x_12130 = x_5470 & x_12129;
assign x_12131 = x_12128 & x_12130;
assign x_12132 = x_5474 & x_5475;
assign x_12133 = x_5473 & x_12132;
assign x_12134 = x_5476 & x_5477;
assign x_12135 = x_5478 & x_5479;
assign x_12136 = x_12134 & x_12135;
assign x_12137 = x_12133 & x_12136;
assign x_12138 = x_12131 & x_12137;
assign x_12139 = x_5481 & x_5482;
assign x_12140 = x_5480 & x_12139;
assign x_12141 = x_5484 & x_5485;
assign x_12142 = x_5483 & x_12141;
assign x_12143 = x_12140 & x_12142;
assign x_12144 = x_5487 & x_5488;
assign x_12145 = x_5486 & x_12144;
assign x_12146 = x_5489 & x_5490;
assign x_12147 = x_5491 & x_5492;
assign x_12148 = x_12146 & x_12147;
assign x_12149 = x_12145 & x_12148;
assign x_12150 = x_12143 & x_12149;
assign x_12151 = x_12138 & x_12150;
assign x_12152 = x_5494 & x_5495;
assign x_12153 = x_5493 & x_12152;
assign x_12154 = x_5497 & x_5498;
assign x_12155 = x_5496 & x_12154;
assign x_12156 = x_12153 & x_12155;
assign x_12157 = x_5500 & x_5501;
assign x_12158 = x_5499 & x_12157;
assign x_12159 = x_5502 & x_5503;
assign x_12160 = x_5504 & x_5505;
assign x_12161 = x_12159 & x_12160;
assign x_12162 = x_12158 & x_12161;
assign x_12163 = x_12156 & x_12162;
assign x_12164 = x_5507 & x_5508;
assign x_12165 = x_5506 & x_12164;
assign x_12166 = x_5510 & x_5511;
assign x_12167 = x_5509 & x_12166;
assign x_12168 = x_12165 & x_12167;
assign x_12169 = x_5513 & x_5514;
assign x_12170 = x_5512 & x_12169;
assign x_12171 = x_5515 & x_5516;
assign x_12172 = x_5517 & x_5518;
assign x_12173 = x_12171 & x_12172;
assign x_12174 = x_12170 & x_12173;
assign x_12175 = x_12168 & x_12174;
assign x_12176 = x_12163 & x_12175;
assign x_12177 = x_12151 & x_12176;
assign x_12178 = x_12126 & x_12177;
assign x_12179 = x_5520 & x_5521;
assign x_12180 = x_5519 & x_12179;
assign x_12181 = x_5523 & x_5524;
assign x_12182 = x_5522 & x_12181;
assign x_12183 = x_12180 & x_12182;
assign x_12184 = x_5526 & x_5527;
assign x_12185 = x_5525 & x_12184;
assign x_12186 = x_5528 & x_5529;
assign x_12187 = x_5530 & x_5531;
assign x_12188 = x_12186 & x_12187;
assign x_12189 = x_12185 & x_12188;
assign x_12190 = x_12183 & x_12189;
assign x_12191 = x_5533 & x_5534;
assign x_12192 = x_5532 & x_12191;
assign x_12193 = x_5536 & x_5537;
assign x_12194 = x_5535 & x_12193;
assign x_12195 = x_12192 & x_12194;
assign x_12196 = x_5539 & x_5540;
assign x_12197 = x_5538 & x_12196;
assign x_12198 = x_5541 & x_5542;
assign x_12199 = x_5543 & x_5544;
assign x_12200 = x_12198 & x_12199;
assign x_12201 = x_12197 & x_12200;
assign x_12202 = x_12195 & x_12201;
assign x_12203 = x_12190 & x_12202;
assign x_12204 = x_5546 & x_5547;
assign x_12205 = x_5545 & x_12204;
assign x_12206 = x_5549 & x_5550;
assign x_12207 = x_5548 & x_12206;
assign x_12208 = x_12205 & x_12207;
assign x_12209 = x_5552 & x_5553;
assign x_12210 = x_5551 & x_12209;
assign x_12211 = x_5554 & x_5555;
assign x_12212 = x_5556 & x_5557;
assign x_12213 = x_12211 & x_12212;
assign x_12214 = x_12210 & x_12213;
assign x_12215 = x_12208 & x_12214;
assign x_12216 = x_5559 & x_5560;
assign x_12217 = x_5558 & x_12216;
assign x_12218 = x_5562 & x_5563;
assign x_12219 = x_5561 & x_12218;
assign x_12220 = x_12217 & x_12219;
assign x_12221 = x_5565 & x_5566;
assign x_12222 = x_5564 & x_12221;
assign x_12223 = x_5567 & x_5568;
assign x_12224 = x_5569 & x_5570;
assign x_12225 = x_12223 & x_12224;
assign x_12226 = x_12222 & x_12225;
assign x_12227 = x_12220 & x_12226;
assign x_12228 = x_12215 & x_12227;
assign x_12229 = x_12203 & x_12228;
assign x_12230 = x_5572 & x_5573;
assign x_12231 = x_5571 & x_12230;
assign x_12232 = x_5575 & x_5576;
assign x_12233 = x_5574 & x_12232;
assign x_12234 = x_12231 & x_12233;
assign x_12235 = x_5578 & x_5579;
assign x_12236 = x_5577 & x_12235;
assign x_12237 = x_5580 & x_5581;
assign x_12238 = x_5582 & x_5583;
assign x_12239 = x_12237 & x_12238;
assign x_12240 = x_12236 & x_12239;
assign x_12241 = x_12234 & x_12240;
assign x_12242 = x_5585 & x_5586;
assign x_12243 = x_5584 & x_12242;
assign x_12244 = x_5588 & x_5589;
assign x_12245 = x_5587 & x_12244;
assign x_12246 = x_12243 & x_12245;
assign x_12247 = x_5591 & x_5592;
assign x_12248 = x_5590 & x_12247;
assign x_12249 = x_5593 & x_5594;
assign x_12250 = x_5595 & x_5596;
assign x_12251 = x_12249 & x_12250;
assign x_12252 = x_12248 & x_12251;
assign x_12253 = x_12246 & x_12252;
assign x_12254 = x_12241 & x_12253;
assign x_12255 = x_5598 & x_5599;
assign x_12256 = x_5597 & x_12255;
assign x_12257 = x_5601 & x_5602;
assign x_12258 = x_5600 & x_12257;
assign x_12259 = x_12256 & x_12258;
assign x_12260 = x_5604 & x_5605;
assign x_12261 = x_5603 & x_12260;
assign x_12262 = x_5606 & x_5607;
assign x_12263 = x_5608 & x_5609;
assign x_12264 = x_12262 & x_12263;
assign x_12265 = x_12261 & x_12264;
assign x_12266 = x_12259 & x_12265;
assign x_12267 = x_5611 & x_5612;
assign x_12268 = x_5610 & x_12267;
assign x_12269 = x_5614 & x_5615;
assign x_12270 = x_5613 & x_12269;
assign x_12271 = x_12268 & x_12270;
assign x_12272 = x_5617 & x_5618;
assign x_12273 = x_5616 & x_12272;
assign x_12274 = x_5619 & x_5620;
assign x_12275 = x_5621 & x_5622;
assign x_12276 = x_12274 & x_12275;
assign x_12277 = x_12273 & x_12276;
assign x_12278 = x_12271 & x_12277;
assign x_12279 = x_12266 & x_12278;
assign x_12280 = x_12254 & x_12279;
assign x_12281 = x_12229 & x_12280;
assign x_12282 = x_12178 & x_12281;
assign x_12283 = x_5624 & x_5625;
assign x_12284 = x_5623 & x_12283;
assign x_12285 = x_5627 & x_5628;
assign x_12286 = x_5626 & x_12285;
assign x_12287 = x_12284 & x_12286;
assign x_12288 = x_5630 & x_5631;
assign x_12289 = x_5629 & x_12288;
assign x_12290 = x_5632 & x_5633;
assign x_12291 = x_5634 & x_5635;
assign x_12292 = x_12290 & x_12291;
assign x_12293 = x_12289 & x_12292;
assign x_12294 = x_12287 & x_12293;
assign x_12295 = x_5637 & x_5638;
assign x_12296 = x_5636 & x_12295;
assign x_12297 = x_5640 & x_5641;
assign x_12298 = x_5639 & x_12297;
assign x_12299 = x_12296 & x_12298;
assign x_12300 = x_5643 & x_5644;
assign x_12301 = x_5642 & x_12300;
assign x_12302 = x_5645 & x_5646;
assign x_12303 = x_5647 & x_5648;
assign x_12304 = x_12302 & x_12303;
assign x_12305 = x_12301 & x_12304;
assign x_12306 = x_12299 & x_12305;
assign x_12307 = x_12294 & x_12306;
assign x_12308 = x_5650 & x_5651;
assign x_12309 = x_5649 & x_12308;
assign x_12310 = x_5653 & x_5654;
assign x_12311 = x_5652 & x_12310;
assign x_12312 = x_12309 & x_12311;
assign x_12313 = x_5656 & x_5657;
assign x_12314 = x_5655 & x_12313;
assign x_12315 = x_5658 & x_5659;
assign x_12316 = x_5660 & x_5661;
assign x_12317 = x_12315 & x_12316;
assign x_12318 = x_12314 & x_12317;
assign x_12319 = x_12312 & x_12318;
assign x_12320 = x_5663 & x_5664;
assign x_12321 = x_5662 & x_12320;
assign x_12322 = x_5666 & x_5667;
assign x_12323 = x_5665 & x_12322;
assign x_12324 = x_12321 & x_12323;
assign x_12325 = x_5669 & x_5670;
assign x_12326 = x_5668 & x_12325;
assign x_12327 = x_5671 & x_5672;
assign x_12328 = x_5673 & x_5674;
assign x_12329 = x_12327 & x_12328;
assign x_12330 = x_12326 & x_12329;
assign x_12331 = x_12324 & x_12330;
assign x_12332 = x_12319 & x_12331;
assign x_12333 = x_12307 & x_12332;
assign x_12334 = x_5676 & x_5677;
assign x_12335 = x_5675 & x_12334;
assign x_12336 = x_5679 & x_5680;
assign x_12337 = x_5678 & x_12336;
assign x_12338 = x_12335 & x_12337;
assign x_12339 = x_5682 & x_5683;
assign x_12340 = x_5681 & x_12339;
assign x_12341 = x_5684 & x_5685;
assign x_12342 = x_5686 & x_5687;
assign x_12343 = x_12341 & x_12342;
assign x_12344 = x_12340 & x_12343;
assign x_12345 = x_12338 & x_12344;
assign x_12346 = x_5689 & x_5690;
assign x_12347 = x_5688 & x_12346;
assign x_12348 = x_5692 & x_5693;
assign x_12349 = x_5691 & x_12348;
assign x_12350 = x_12347 & x_12349;
assign x_12351 = x_5695 & x_5696;
assign x_12352 = x_5694 & x_12351;
assign x_12353 = x_5697 & x_5698;
assign x_12354 = x_5699 & x_5700;
assign x_12355 = x_12353 & x_12354;
assign x_12356 = x_12352 & x_12355;
assign x_12357 = x_12350 & x_12356;
assign x_12358 = x_12345 & x_12357;
assign x_12359 = x_5702 & x_5703;
assign x_12360 = x_5701 & x_12359;
assign x_12361 = x_5705 & x_5706;
assign x_12362 = x_5704 & x_12361;
assign x_12363 = x_12360 & x_12362;
assign x_12364 = x_5708 & x_5709;
assign x_12365 = x_5707 & x_12364;
assign x_12366 = x_5710 & x_5711;
assign x_12367 = x_5712 & x_5713;
assign x_12368 = x_12366 & x_12367;
assign x_12369 = x_12365 & x_12368;
assign x_12370 = x_12363 & x_12369;
assign x_12371 = x_5715 & x_5716;
assign x_12372 = x_5714 & x_12371;
assign x_12373 = x_5718 & x_5719;
assign x_12374 = x_5717 & x_12373;
assign x_12375 = x_12372 & x_12374;
assign x_12376 = x_5721 & x_5722;
assign x_12377 = x_5720 & x_12376;
assign x_12378 = x_5723 & x_5724;
assign x_12379 = x_5725 & x_5726;
assign x_12380 = x_12378 & x_12379;
assign x_12381 = x_12377 & x_12380;
assign x_12382 = x_12375 & x_12381;
assign x_12383 = x_12370 & x_12382;
assign x_12384 = x_12358 & x_12383;
assign x_12385 = x_12333 & x_12384;
assign x_12386 = x_5728 & x_5729;
assign x_12387 = x_5727 & x_12386;
assign x_12388 = x_5731 & x_5732;
assign x_12389 = x_5730 & x_12388;
assign x_12390 = x_12387 & x_12389;
assign x_12391 = x_5734 & x_5735;
assign x_12392 = x_5733 & x_12391;
assign x_12393 = x_5736 & x_5737;
assign x_12394 = x_5738 & x_5739;
assign x_12395 = x_12393 & x_12394;
assign x_12396 = x_12392 & x_12395;
assign x_12397 = x_12390 & x_12396;
assign x_12398 = x_5741 & x_5742;
assign x_12399 = x_5740 & x_12398;
assign x_12400 = x_5744 & x_5745;
assign x_12401 = x_5743 & x_12400;
assign x_12402 = x_12399 & x_12401;
assign x_12403 = x_5747 & x_5748;
assign x_12404 = x_5746 & x_12403;
assign x_12405 = x_5749 & x_5750;
assign x_12406 = x_5751 & x_5752;
assign x_12407 = x_12405 & x_12406;
assign x_12408 = x_12404 & x_12407;
assign x_12409 = x_12402 & x_12408;
assign x_12410 = x_12397 & x_12409;
assign x_12411 = x_5754 & x_5755;
assign x_12412 = x_5753 & x_12411;
assign x_12413 = x_5757 & x_5758;
assign x_12414 = x_5756 & x_12413;
assign x_12415 = x_12412 & x_12414;
assign x_12416 = x_5760 & x_5761;
assign x_12417 = x_5759 & x_12416;
assign x_12418 = x_5762 & x_5763;
assign x_12419 = x_5764 & x_5765;
assign x_12420 = x_12418 & x_12419;
assign x_12421 = x_12417 & x_12420;
assign x_12422 = x_12415 & x_12421;
assign x_12423 = x_5767 & x_5768;
assign x_12424 = x_5766 & x_12423;
assign x_12425 = x_5770 & x_5771;
assign x_12426 = x_5769 & x_12425;
assign x_12427 = x_12424 & x_12426;
assign x_12428 = x_5773 & x_5774;
assign x_12429 = x_5772 & x_12428;
assign x_12430 = x_5775 & x_5776;
assign x_12431 = x_5777 & x_5778;
assign x_12432 = x_12430 & x_12431;
assign x_12433 = x_12429 & x_12432;
assign x_12434 = x_12427 & x_12433;
assign x_12435 = x_12422 & x_12434;
assign x_12436 = x_12410 & x_12435;
assign x_12437 = x_5780 & x_5781;
assign x_12438 = x_5779 & x_12437;
assign x_12439 = x_5783 & x_5784;
assign x_12440 = x_5782 & x_12439;
assign x_12441 = x_12438 & x_12440;
assign x_12442 = x_5786 & x_5787;
assign x_12443 = x_5785 & x_12442;
assign x_12444 = x_5788 & x_5789;
assign x_12445 = x_5790 & x_5791;
assign x_12446 = x_12444 & x_12445;
assign x_12447 = x_12443 & x_12446;
assign x_12448 = x_12441 & x_12447;
assign x_12449 = x_5793 & x_5794;
assign x_12450 = x_5792 & x_12449;
assign x_12451 = x_5796 & x_5797;
assign x_12452 = x_5795 & x_12451;
assign x_12453 = x_12450 & x_12452;
assign x_12454 = x_5799 & x_5800;
assign x_12455 = x_5798 & x_12454;
assign x_12456 = x_5801 & x_5802;
assign x_12457 = x_5803 & x_5804;
assign x_12458 = x_12456 & x_12457;
assign x_12459 = x_12455 & x_12458;
assign x_12460 = x_12453 & x_12459;
assign x_12461 = x_12448 & x_12460;
assign x_12462 = x_5806 & x_5807;
assign x_12463 = x_5805 & x_12462;
assign x_12464 = x_5809 & x_5810;
assign x_12465 = x_5808 & x_12464;
assign x_12466 = x_12463 & x_12465;
assign x_12467 = x_5812 & x_5813;
assign x_12468 = x_5811 & x_12467;
assign x_12469 = x_5814 & x_5815;
assign x_12470 = x_5816 & x_5817;
assign x_12471 = x_12469 & x_12470;
assign x_12472 = x_12468 & x_12471;
assign x_12473 = x_12466 & x_12472;
assign x_12474 = x_5819 & x_5820;
assign x_12475 = x_5818 & x_12474;
assign x_12476 = x_5821 & x_5822;
assign x_12477 = x_5823 & x_5824;
assign x_12478 = x_12476 & x_12477;
assign x_12479 = x_12475 & x_12478;
assign x_12480 = x_5826 & x_5827;
assign x_12481 = x_5825 & x_12480;
assign x_12482 = x_5828 & x_5829;
assign x_12483 = x_5830 & x_5831;
assign x_12484 = x_12482 & x_12483;
assign x_12485 = x_12481 & x_12484;
assign x_12486 = x_12479 & x_12485;
assign x_12487 = x_12473 & x_12486;
assign x_12488 = x_12461 & x_12487;
assign x_12489 = x_12436 & x_12488;
assign x_12490 = x_12385 & x_12489;
assign x_12491 = x_12282 & x_12490;
assign x_12492 = x_12075 & x_12491;
assign x_12493 = x_5833 & x_5834;
assign x_12494 = x_5832 & x_12493;
assign x_12495 = x_5836 & x_5837;
assign x_12496 = x_5835 & x_12495;
assign x_12497 = x_12494 & x_12496;
assign x_12498 = x_5839 & x_5840;
assign x_12499 = x_5838 & x_12498;
assign x_12500 = x_5841 & x_5842;
assign x_12501 = x_5843 & x_5844;
assign x_12502 = x_12500 & x_12501;
assign x_12503 = x_12499 & x_12502;
assign x_12504 = x_12497 & x_12503;
assign x_12505 = x_5846 & x_5847;
assign x_12506 = x_5845 & x_12505;
assign x_12507 = x_5849 & x_5850;
assign x_12508 = x_5848 & x_12507;
assign x_12509 = x_12506 & x_12508;
assign x_12510 = x_5852 & x_5853;
assign x_12511 = x_5851 & x_12510;
assign x_12512 = x_5854 & x_5855;
assign x_12513 = x_5856 & x_5857;
assign x_12514 = x_12512 & x_12513;
assign x_12515 = x_12511 & x_12514;
assign x_12516 = x_12509 & x_12515;
assign x_12517 = x_12504 & x_12516;
assign x_12518 = x_5859 & x_5860;
assign x_12519 = x_5858 & x_12518;
assign x_12520 = x_5862 & x_5863;
assign x_12521 = x_5861 & x_12520;
assign x_12522 = x_12519 & x_12521;
assign x_12523 = x_5865 & x_5866;
assign x_12524 = x_5864 & x_12523;
assign x_12525 = x_5867 & x_5868;
assign x_12526 = x_5869 & x_5870;
assign x_12527 = x_12525 & x_12526;
assign x_12528 = x_12524 & x_12527;
assign x_12529 = x_12522 & x_12528;
assign x_12530 = x_5872 & x_5873;
assign x_12531 = x_5871 & x_12530;
assign x_12532 = x_5875 & x_5876;
assign x_12533 = x_5874 & x_12532;
assign x_12534 = x_12531 & x_12533;
assign x_12535 = x_5878 & x_5879;
assign x_12536 = x_5877 & x_12535;
assign x_12537 = x_5880 & x_5881;
assign x_12538 = x_5882 & x_5883;
assign x_12539 = x_12537 & x_12538;
assign x_12540 = x_12536 & x_12539;
assign x_12541 = x_12534 & x_12540;
assign x_12542 = x_12529 & x_12541;
assign x_12543 = x_12517 & x_12542;
assign x_12544 = x_5885 & x_5886;
assign x_12545 = x_5884 & x_12544;
assign x_12546 = x_5888 & x_5889;
assign x_12547 = x_5887 & x_12546;
assign x_12548 = x_12545 & x_12547;
assign x_12549 = x_5891 & x_5892;
assign x_12550 = x_5890 & x_12549;
assign x_12551 = x_5893 & x_5894;
assign x_12552 = x_5895 & x_5896;
assign x_12553 = x_12551 & x_12552;
assign x_12554 = x_12550 & x_12553;
assign x_12555 = x_12548 & x_12554;
assign x_12556 = x_5898 & x_5899;
assign x_12557 = x_5897 & x_12556;
assign x_12558 = x_5901 & x_5902;
assign x_12559 = x_5900 & x_12558;
assign x_12560 = x_12557 & x_12559;
assign x_12561 = x_5904 & x_5905;
assign x_12562 = x_5903 & x_12561;
assign x_12563 = x_5906 & x_5907;
assign x_12564 = x_5908 & x_5909;
assign x_12565 = x_12563 & x_12564;
assign x_12566 = x_12562 & x_12565;
assign x_12567 = x_12560 & x_12566;
assign x_12568 = x_12555 & x_12567;
assign x_12569 = x_5911 & x_5912;
assign x_12570 = x_5910 & x_12569;
assign x_12571 = x_5914 & x_5915;
assign x_12572 = x_5913 & x_12571;
assign x_12573 = x_12570 & x_12572;
assign x_12574 = x_5917 & x_5918;
assign x_12575 = x_5916 & x_12574;
assign x_12576 = x_5919 & x_5920;
assign x_12577 = x_5921 & x_5922;
assign x_12578 = x_12576 & x_12577;
assign x_12579 = x_12575 & x_12578;
assign x_12580 = x_12573 & x_12579;
assign x_12581 = x_5924 & x_5925;
assign x_12582 = x_5923 & x_12581;
assign x_12583 = x_5927 & x_5928;
assign x_12584 = x_5926 & x_12583;
assign x_12585 = x_12582 & x_12584;
assign x_12586 = x_5930 & x_5931;
assign x_12587 = x_5929 & x_12586;
assign x_12588 = x_5932 & x_5933;
assign x_12589 = x_5934 & x_5935;
assign x_12590 = x_12588 & x_12589;
assign x_12591 = x_12587 & x_12590;
assign x_12592 = x_12585 & x_12591;
assign x_12593 = x_12580 & x_12592;
assign x_12594 = x_12568 & x_12593;
assign x_12595 = x_12543 & x_12594;
assign x_12596 = x_5937 & x_5938;
assign x_12597 = x_5936 & x_12596;
assign x_12598 = x_5940 & x_5941;
assign x_12599 = x_5939 & x_12598;
assign x_12600 = x_12597 & x_12599;
assign x_12601 = x_5943 & x_5944;
assign x_12602 = x_5942 & x_12601;
assign x_12603 = x_5945 & x_5946;
assign x_12604 = x_5947 & x_5948;
assign x_12605 = x_12603 & x_12604;
assign x_12606 = x_12602 & x_12605;
assign x_12607 = x_12600 & x_12606;
assign x_12608 = x_5950 & x_5951;
assign x_12609 = x_5949 & x_12608;
assign x_12610 = x_5953 & x_5954;
assign x_12611 = x_5952 & x_12610;
assign x_12612 = x_12609 & x_12611;
assign x_12613 = x_5956 & x_5957;
assign x_12614 = x_5955 & x_12613;
assign x_12615 = x_5958 & x_5959;
assign x_12616 = x_5960 & x_5961;
assign x_12617 = x_12615 & x_12616;
assign x_12618 = x_12614 & x_12617;
assign x_12619 = x_12612 & x_12618;
assign x_12620 = x_12607 & x_12619;
assign x_12621 = x_5963 & x_5964;
assign x_12622 = x_5962 & x_12621;
assign x_12623 = x_5966 & x_5967;
assign x_12624 = x_5965 & x_12623;
assign x_12625 = x_12622 & x_12624;
assign x_12626 = x_5969 & x_5970;
assign x_12627 = x_5968 & x_12626;
assign x_12628 = x_5971 & x_5972;
assign x_12629 = x_5973 & x_5974;
assign x_12630 = x_12628 & x_12629;
assign x_12631 = x_12627 & x_12630;
assign x_12632 = x_12625 & x_12631;
assign x_12633 = x_5976 & x_5977;
assign x_12634 = x_5975 & x_12633;
assign x_12635 = x_5979 & x_5980;
assign x_12636 = x_5978 & x_12635;
assign x_12637 = x_12634 & x_12636;
assign x_12638 = x_5982 & x_5983;
assign x_12639 = x_5981 & x_12638;
assign x_12640 = x_5984 & x_5985;
assign x_12641 = x_5986 & x_5987;
assign x_12642 = x_12640 & x_12641;
assign x_12643 = x_12639 & x_12642;
assign x_12644 = x_12637 & x_12643;
assign x_12645 = x_12632 & x_12644;
assign x_12646 = x_12620 & x_12645;
assign x_12647 = x_5989 & x_5990;
assign x_12648 = x_5988 & x_12647;
assign x_12649 = x_5992 & x_5993;
assign x_12650 = x_5991 & x_12649;
assign x_12651 = x_12648 & x_12650;
assign x_12652 = x_5995 & x_5996;
assign x_12653 = x_5994 & x_12652;
assign x_12654 = x_5997 & x_5998;
assign x_12655 = x_5999 & x_6000;
assign x_12656 = x_12654 & x_12655;
assign x_12657 = x_12653 & x_12656;
assign x_12658 = x_12651 & x_12657;
assign x_12659 = x_6002 & x_6003;
assign x_12660 = x_6001 & x_12659;
assign x_12661 = x_6005 & x_6006;
assign x_12662 = x_6004 & x_12661;
assign x_12663 = x_12660 & x_12662;
assign x_12664 = x_6008 & x_6009;
assign x_12665 = x_6007 & x_12664;
assign x_12666 = x_6010 & x_6011;
assign x_12667 = x_6012 & x_6013;
assign x_12668 = x_12666 & x_12667;
assign x_12669 = x_12665 & x_12668;
assign x_12670 = x_12663 & x_12669;
assign x_12671 = x_12658 & x_12670;
assign x_12672 = x_6015 & x_6016;
assign x_12673 = x_6014 & x_12672;
assign x_12674 = x_6018 & x_6019;
assign x_12675 = x_6017 & x_12674;
assign x_12676 = x_12673 & x_12675;
assign x_12677 = x_6021 & x_6022;
assign x_12678 = x_6020 & x_12677;
assign x_12679 = x_6023 & x_6024;
assign x_12680 = x_6025 & x_6026;
assign x_12681 = x_12679 & x_12680;
assign x_12682 = x_12678 & x_12681;
assign x_12683 = x_12676 & x_12682;
assign x_12684 = x_6028 & x_6029;
assign x_12685 = x_6027 & x_12684;
assign x_12686 = x_6031 & x_6032;
assign x_12687 = x_6030 & x_12686;
assign x_12688 = x_12685 & x_12687;
assign x_12689 = x_6034 & x_6035;
assign x_12690 = x_6033 & x_12689;
assign x_12691 = x_6036 & x_6037;
assign x_12692 = x_6038 & x_6039;
assign x_12693 = x_12691 & x_12692;
assign x_12694 = x_12690 & x_12693;
assign x_12695 = x_12688 & x_12694;
assign x_12696 = x_12683 & x_12695;
assign x_12697 = x_12671 & x_12696;
assign x_12698 = x_12646 & x_12697;
assign x_12699 = x_12595 & x_12698;
assign x_12700 = x_6041 & x_6042;
assign x_12701 = x_6040 & x_12700;
assign x_12702 = x_6044 & x_6045;
assign x_12703 = x_6043 & x_12702;
assign x_12704 = x_12701 & x_12703;
assign x_12705 = x_6047 & x_6048;
assign x_12706 = x_6046 & x_12705;
assign x_12707 = x_6049 & x_6050;
assign x_12708 = x_6051 & x_6052;
assign x_12709 = x_12707 & x_12708;
assign x_12710 = x_12706 & x_12709;
assign x_12711 = x_12704 & x_12710;
assign x_12712 = x_6054 & x_6055;
assign x_12713 = x_6053 & x_12712;
assign x_12714 = x_6057 & x_6058;
assign x_12715 = x_6056 & x_12714;
assign x_12716 = x_12713 & x_12715;
assign x_12717 = x_6060 & x_6061;
assign x_12718 = x_6059 & x_12717;
assign x_12719 = x_6062 & x_6063;
assign x_12720 = x_6064 & x_6065;
assign x_12721 = x_12719 & x_12720;
assign x_12722 = x_12718 & x_12721;
assign x_12723 = x_12716 & x_12722;
assign x_12724 = x_12711 & x_12723;
assign x_12725 = x_6067 & x_6068;
assign x_12726 = x_6066 & x_12725;
assign x_12727 = x_6070 & x_6071;
assign x_12728 = x_6069 & x_12727;
assign x_12729 = x_12726 & x_12728;
assign x_12730 = x_6073 & x_6074;
assign x_12731 = x_6072 & x_12730;
assign x_12732 = x_6075 & x_6076;
assign x_12733 = x_6077 & x_6078;
assign x_12734 = x_12732 & x_12733;
assign x_12735 = x_12731 & x_12734;
assign x_12736 = x_12729 & x_12735;
assign x_12737 = x_6080 & x_6081;
assign x_12738 = x_6079 & x_12737;
assign x_12739 = x_6083 & x_6084;
assign x_12740 = x_6082 & x_12739;
assign x_12741 = x_12738 & x_12740;
assign x_12742 = x_6086 & x_6087;
assign x_12743 = x_6085 & x_12742;
assign x_12744 = x_6088 & x_6089;
assign x_12745 = x_6090 & x_6091;
assign x_12746 = x_12744 & x_12745;
assign x_12747 = x_12743 & x_12746;
assign x_12748 = x_12741 & x_12747;
assign x_12749 = x_12736 & x_12748;
assign x_12750 = x_12724 & x_12749;
assign x_12751 = x_6093 & x_6094;
assign x_12752 = x_6092 & x_12751;
assign x_12753 = x_6096 & x_6097;
assign x_12754 = x_6095 & x_12753;
assign x_12755 = x_12752 & x_12754;
assign x_12756 = x_6099 & x_6100;
assign x_12757 = x_6098 & x_12756;
assign x_12758 = x_6101 & x_6102;
assign x_12759 = x_6103 & x_6104;
assign x_12760 = x_12758 & x_12759;
assign x_12761 = x_12757 & x_12760;
assign x_12762 = x_12755 & x_12761;
assign x_12763 = x_6106 & x_6107;
assign x_12764 = x_6105 & x_12763;
assign x_12765 = x_6109 & x_6110;
assign x_12766 = x_6108 & x_12765;
assign x_12767 = x_12764 & x_12766;
assign x_12768 = x_6112 & x_6113;
assign x_12769 = x_6111 & x_12768;
assign x_12770 = x_6114 & x_6115;
assign x_12771 = x_6116 & x_6117;
assign x_12772 = x_12770 & x_12771;
assign x_12773 = x_12769 & x_12772;
assign x_12774 = x_12767 & x_12773;
assign x_12775 = x_12762 & x_12774;
assign x_12776 = x_6119 & x_6120;
assign x_12777 = x_6118 & x_12776;
assign x_12778 = x_6122 & x_6123;
assign x_12779 = x_6121 & x_12778;
assign x_12780 = x_12777 & x_12779;
assign x_12781 = x_6125 & x_6126;
assign x_12782 = x_6124 & x_12781;
assign x_12783 = x_6127 & x_6128;
assign x_12784 = x_6129 & x_6130;
assign x_12785 = x_12783 & x_12784;
assign x_12786 = x_12782 & x_12785;
assign x_12787 = x_12780 & x_12786;
assign x_12788 = x_6132 & x_6133;
assign x_12789 = x_6131 & x_12788;
assign x_12790 = x_6135 & x_6136;
assign x_12791 = x_6134 & x_12790;
assign x_12792 = x_12789 & x_12791;
assign x_12793 = x_6138 & x_6139;
assign x_12794 = x_6137 & x_12793;
assign x_12795 = x_6140 & x_6141;
assign x_12796 = x_6142 & x_6143;
assign x_12797 = x_12795 & x_12796;
assign x_12798 = x_12794 & x_12797;
assign x_12799 = x_12792 & x_12798;
assign x_12800 = x_12787 & x_12799;
assign x_12801 = x_12775 & x_12800;
assign x_12802 = x_12750 & x_12801;
assign x_12803 = x_6145 & x_6146;
assign x_12804 = x_6144 & x_12803;
assign x_12805 = x_6148 & x_6149;
assign x_12806 = x_6147 & x_12805;
assign x_12807 = x_12804 & x_12806;
assign x_12808 = x_6151 & x_6152;
assign x_12809 = x_6150 & x_12808;
assign x_12810 = x_6153 & x_6154;
assign x_12811 = x_6155 & x_6156;
assign x_12812 = x_12810 & x_12811;
assign x_12813 = x_12809 & x_12812;
assign x_12814 = x_12807 & x_12813;
assign x_12815 = x_6158 & x_6159;
assign x_12816 = x_6157 & x_12815;
assign x_12817 = x_6161 & x_6162;
assign x_12818 = x_6160 & x_12817;
assign x_12819 = x_12816 & x_12818;
assign x_12820 = x_6164 & x_6165;
assign x_12821 = x_6163 & x_12820;
assign x_12822 = x_6166 & x_6167;
assign x_12823 = x_6168 & x_6169;
assign x_12824 = x_12822 & x_12823;
assign x_12825 = x_12821 & x_12824;
assign x_12826 = x_12819 & x_12825;
assign x_12827 = x_12814 & x_12826;
assign x_12828 = x_6171 & x_6172;
assign x_12829 = x_6170 & x_12828;
assign x_12830 = x_6174 & x_6175;
assign x_12831 = x_6173 & x_12830;
assign x_12832 = x_12829 & x_12831;
assign x_12833 = x_6177 & x_6178;
assign x_12834 = x_6176 & x_12833;
assign x_12835 = x_6179 & x_6180;
assign x_12836 = x_6181 & x_6182;
assign x_12837 = x_12835 & x_12836;
assign x_12838 = x_12834 & x_12837;
assign x_12839 = x_12832 & x_12838;
assign x_12840 = x_6184 & x_6185;
assign x_12841 = x_6183 & x_12840;
assign x_12842 = x_6187 & x_6188;
assign x_12843 = x_6186 & x_12842;
assign x_12844 = x_12841 & x_12843;
assign x_12845 = x_6190 & x_6191;
assign x_12846 = x_6189 & x_12845;
assign x_12847 = x_6192 & x_6193;
assign x_12848 = x_6194 & x_6195;
assign x_12849 = x_12847 & x_12848;
assign x_12850 = x_12846 & x_12849;
assign x_12851 = x_12844 & x_12850;
assign x_12852 = x_12839 & x_12851;
assign x_12853 = x_12827 & x_12852;
assign x_12854 = x_6197 & x_6198;
assign x_12855 = x_6196 & x_12854;
assign x_12856 = x_6200 & x_6201;
assign x_12857 = x_6199 & x_12856;
assign x_12858 = x_12855 & x_12857;
assign x_12859 = x_6203 & x_6204;
assign x_12860 = x_6202 & x_12859;
assign x_12861 = x_6205 & x_6206;
assign x_12862 = x_6207 & x_6208;
assign x_12863 = x_12861 & x_12862;
assign x_12864 = x_12860 & x_12863;
assign x_12865 = x_12858 & x_12864;
assign x_12866 = x_6210 & x_6211;
assign x_12867 = x_6209 & x_12866;
assign x_12868 = x_6213 & x_6214;
assign x_12869 = x_6212 & x_12868;
assign x_12870 = x_12867 & x_12869;
assign x_12871 = x_6216 & x_6217;
assign x_12872 = x_6215 & x_12871;
assign x_12873 = x_6218 & x_6219;
assign x_12874 = x_6220 & x_6221;
assign x_12875 = x_12873 & x_12874;
assign x_12876 = x_12872 & x_12875;
assign x_12877 = x_12870 & x_12876;
assign x_12878 = x_12865 & x_12877;
assign x_12879 = x_6223 & x_6224;
assign x_12880 = x_6222 & x_12879;
assign x_12881 = x_6226 & x_6227;
assign x_12882 = x_6225 & x_12881;
assign x_12883 = x_12880 & x_12882;
assign x_12884 = x_6229 & x_6230;
assign x_12885 = x_6228 & x_12884;
assign x_12886 = x_6231 & x_6232;
assign x_12887 = x_6233 & x_6234;
assign x_12888 = x_12886 & x_12887;
assign x_12889 = x_12885 & x_12888;
assign x_12890 = x_12883 & x_12889;
assign x_12891 = x_6236 & x_6237;
assign x_12892 = x_6235 & x_12891;
assign x_12893 = x_6239 & x_6240;
assign x_12894 = x_6238 & x_12893;
assign x_12895 = x_12892 & x_12894;
assign x_12896 = x_6242 & x_6243;
assign x_12897 = x_6241 & x_12896;
assign x_12898 = x_6244 & x_6245;
assign x_12899 = x_6246 & x_6247;
assign x_12900 = x_12898 & x_12899;
assign x_12901 = x_12897 & x_12900;
assign x_12902 = x_12895 & x_12901;
assign x_12903 = x_12890 & x_12902;
assign x_12904 = x_12878 & x_12903;
assign x_12905 = x_12853 & x_12904;
assign x_12906 = x_12802 & x_12905;
assign x_12907 = x_12699 & x_12906;
assign x_12908 = x_6249 & x_6250;
assign x_12909 = x_6248 & x_12908;
assign x_12910 = x_6252 & x_6253;
assign x_12911 = x_6251 & x_12910;
assign x_12912 = x_12909 & x_12911;
assign x_12913 = x_6255 & x_6256;
assign x_12914 = x_6254 & x_12913;
assign x_12915 = x_6257 & x_6258;
assign x_12916 = x_6259 & x_6260;
assign x_12917 = x_12915 & x_12916;
assign x_12918 = x_12914 & x_12917;
assign x_12919 = x_12912 & x_12918;
assign x_12920 = x_6262 & x_6263;
assign x_12921 = x_6261 & x_12920;
assign x_12922 = x_6265 & x_6266;
assign x_12923 = x_6264 & x_12922;
assign x_12924 = x_12921 & x_12923;
assign x_12925 = x_6268 & x_6269;
assign x_12926 = x_6267 & x_12925;
assign x_12927 = x_6270 & x_6271;
assign x_12928 = x_6272 & x_6273;
assign x_12929 = x_12927 & x_12928;
assign x_12930 = x_12926 & x_12929;
assign x_12931 = x_12924 & x_12930;
assign x_12932 = x_12919 & x_12931;
assign x_12933 = x_6275 & x_6276;
assign x_12934 = x_6274 & x_12933;
assign x_12935 = x_6278 & x_6279;
assign x_12936 = x_6277 & x_12935;
assign x_12937 = x_12934 & x_12936;
assign x_12938 = x_6281 & x_6282;
assign x_12939 = x_6280 & x_12938;
assign x_12940 = x_6283 & x_6284;
assign x_12941 = x_6285 & x_6286;
assign x_12942 = x_12940 & x_12941;
assign x_12943 = x_12939 & x_12942;
assign x_12944 = x_12937 & x_12943;
assign x_12945 = x_6288 & x_6289;
assign x_12946 = x_6287 & x_12945;
assign x_12947 = x_6291 & x_6292;
assign x_12948 = x_6290 & x_12947;
assign x_12949 = x_12946 & x_12948;
assign x_12950 = x_6294 & x_6295;
assign x_12951 = x_6293 & x_12950;
assign x_12952 = x_6296 & x_6297;
assign x_12953 = x_6298 & x_6299;
assign x_12954 = x_12952 & x_12953;
assign x_12955 = x_12951 & x_12954;
assign x_12956 = x_12949 & x_12955;
assign x_12957 = x_12944 & x_12956;
assign x_12958 = x_12932 & x_12957;
assign x_12959 = x_6301 & x_6302;
assign x_12960 = x_6300 & x_12959;
assign x_12961 = x_6304 & x_6305;
assign x_12962 = x_6303 & x_12961;
assign x_12963 = x_12960 & x_12962;
assign x_12964 = x_6307 & x_6308;
assign x_12965 = x_6306 & x_12964;
assign x_12966 = x_6309 & x_6310;
assign x_12967 = x_6311 & x_6312;
assign x_12968 = x_12966 & x_12967;
assign x_12969 = x_12965 & x_12968;
assign x_12970 = x_12963 & x_12969;
assign x_12971 = x_6314 & x_6315;
assign x_12972 = x_6313 & x_12971;
assign x_12973 = x_6317 & x_6318;
assign x_12974 = x_6316 & x_12973;
assign x_12975 = x_12972 & x_12974;
assign x_12976 = x_6320 & x_6321;
assign x_12977 = x_6319 & x_12976;
assign x_12978 = x_6322 & x_6323;
assign x_12979 = x_6324 & x_6325;
assign x_12980 = x_12978 & x_12979;
assign x_12981 = x_12977 & x_12980;
assign x_12982 = x_12975 & x_12981;
assign x_12983 = x_12970 & x_12982;
assign x_12984 = x_6327 & x_6328;
assign x_12985 = x_6326 & x_12984;
assign x_12986 = x_6330 & x_6331;
assign x_12987 = x_6329 & x_12986;
assign x_12988 = x_12985 & x_12987;
assign x_12989 = x_6333 & x_6334;
assign x_12990 = x_6332 & x_12989;
assign x_12991 = x_6335 & x_6336;
assign x_12992 = x_6337 & x_6338;
assign x_12993 = x_12991 & x_12992;
assign x_12994 = x_12990 & x_12993;
assign x_12995 = x_12988 & x_12994;
assign x_12996 = x_6340 & x_6341;
assign x_12997 = x_6339 & x_12996;
assign x_12998 = x_6343 & x_6344;
assign x_12999 = x_6342 & x_12998;
assign x_13000 = x_12997 & x_12999;
assign x_13001 = x_6346 & x_6347;
assign x_13002 = x_6345 & x_13001;
assign x_13003 = x_6348 & x_6349;
assign x_13004 = x_6350 & x_6351;
assign x_13005 = x_13003 & x_13004;
assign x_13006 = x_13002 & x_13005;
assign x_13007 = x_13000 & x_13006;
assign x_13008 = x_12995 & x_13007;
assign x_13009 = x_12983 & x_13008;
assign x_13010 = x_12958 & x_13009;
assign x_13011 = x_6353 & x_6354;
assign x_13012 = x_6352 & x_13011;
assign x_13013 = x_6356 & x_6357;
assign x_13014 = x_6355 & x_13013;
assign x_13015 = x_13012 & x_13014;
assign x_13016 = x_6359 & x_6360;
assign x_13017 = x_6358 & x_13016;
assign x_13018 = x_6361 & x_6362;
assign x_13019 = x_6363 & x_6364;
assign x_13020 = x_13018 & x_13019;
assign x_13021 = x_13017 & x_13020;
assign x_13022 = x_13015 & x_13021;
assign x_13023 = x_6366 & x_6367;
assign x_13024 = x_6365 & x_13023;
assign x_13025 = x_6369 & x_6370;
assign x_13026 = x_6368 & x_13025;
assign x_13027 = x_13024 & x_13026;
assign x_13028 = x_6372 & x_6373;
assign x_13029 = x_6371 & x_13028;
assign x_13030 = x_6374 & x_6375;
assign x_13031 = x_6376 & x_6377;
assign x_13032 = x_13030 & x_13031;
assign x_13033 = x_13029 & x_13032;
assign x_13034 = x_13027 & x_13033;
assign x_13035 = x_13022 & x_13034;
assign x_13036 = x_6379 & x_6380;
assign x_13037 = x_6378 & x_13036;
assign x_13038 = x_6382 & x_6383;
assign x_13039 = x_6381 & x_13038;
assign x_13040 = x_13037 & x_13039;
assign x_13041 = x_6385 & x_6386;
assign x_13042 = x_6384 & x_13041;
assign x_13043 = x_6387 & x_6388;
assign x_13044 = x_6389 & x_6390;
assign x_13045 = x_13043 & x_13044;
assign x_13046 = x_13042 & x_13045;
assign x_13047 = x_13040 & x_13046;
assign x_13048 = x_6392 & x_6393;
assign x_13049 = x_6391 & x_13048;
assign x_13050 = x_6395 & x_6396;
assign x_13051 = x_6394 & x_13050;
assign x_13052 = x_13049 & x_13051;
assign x_13053 = x_6398 & x_6399;
assign x_13054 = x_6397 & x_13053;
assign x_13055 = x_6400 & x_6401;
assign x_13056 = x_6402 & x_6403;
assign x_13057 = x_13055 & x_13056;
assign x_13058 = x_13054 & x_13057;
assign x_13059 = x_13052 & x_13058;
assign x_13060 = x_13047 & x_13059;
assign x_13061 = x_13035 & x_13060;
assign x_13062 = x_6405 & x_6406;
assign x_13063 = x_6404 & x_13062;
assign x_13064 = x_6408 & x_6409;
assign x_13065 = x_6407 & x_13064;
assign x_13066 = x_13063 & x_13065;
assign x_13067 = x_6411 & x_6412;
assign x_13068 = x_6410 & x_13067;
assign x_13069 = x_6413 & x_6414;
assign x_13070 = x_6415 & x_6416;
assign x_13071 = x_13069 & x_13070;
assign x_13072 = x_13068 & x_13071;
assign x_13073 = x_13066 & x_13072;
assign x_13074 = x_6418 & x_6419;
assign x_13075 = x_6417 & x_13074;
assign x_13076 = x_6421 & x_6422;
assign x_13077 = x_6420 & x_13076;
assign x_13078 = x_13075 & x_13077;
assign x_13079 = x_6424 & x_6425;
assign x_13080 = x_6423 & x_13079;
assign x_13081 = x_6426 & x_6427;
assign x_13082 = x_6428 & x_6429;
assign x_13083 = x_13081 & x_13082;
assign x_13084 = x_13080 & x_13083;
assign x_13085 = x_13078 & x_13084;
assign x_13086 = x_13073 & x_13085;
assign x_13087 = x_6431 & x_6432;
assign x_13088 = x_6430 & x_13087;
assign x_13089 = x_6434 & x_6435;
assign x_13090 = x_6433 & x_13089;
assign x_13091 = x_13088 & x_13090;
assign x_13092 = x_6437 & x_6438;
assign x_13093 = x_6436 & x_13092;
assign x_13094 = x_6439 & x_6440;
assign x_13095 = x_6441 & x_6442;
assign x_13096 = x_13094 & x_13095;
assign x_13097 = x_13093 & x_13096;
assign x_13098 = x_13091 & x_13097;
assign x_13099 = x_6444 & x_6445;
assign x_13100 = x_6443 & x_13099;
assign x_13101 = x_6447 & x_6448;
assign x_13102 = x_6446 & x_13101;
assign x_13103 = x_13100 & x_13102;
assign x_13104 = x_6450 & x_6451;
assign x_13105 = x_6449 & x_13104;
assign x_13106 = x_6452 & x_6453;
assign x_13107 = x_6454 & x_6455;
assign x_13108 = x_13106 & x_13107;
assign x_13109 = x_13105 & x_13108;
assign x_13110 = x_13103 & x_13109;
assign x_13111 = x_13098 & x_13110;
assign x_13112 = x_13086 & x_13111;
assign x_13113 = x_13061 & x_13112;
assign x_13114 = x_13010 & x_13113;
assign x_13115 = x_6457 & x_6458;
assign x_13116 = x_6456 & x_13115;
assign x_13117 = x_6460 & x_6461;
assign x_13118 = x_6459 & x_13117;
assign x_13119 = x_13116 & x_13118;
assign x_13120 = x_6463 & x_6464;
assign x_13121 = x_6462 & x_13120;
assign x_13122 = x_6465 & x_6466;
assign x_13123 = x_6467 & x_6468;
assign x_13124 = x_13122 & x_13123;
assign x_13125 = x_13121 & x_13124;
assign x_13126 = x_13119 & x_13125;
assign x_13127 = x_6470 & x_6471;
assign x_13128 = x_6469 & x_13127;
assign x_13129 = x_6473 & x_6474;
assign x_13130 = x_6472 & x_13129;
assign x_13131 = x_13128 & x_13130;
assign x_13132 = x_6476 & x_6477;
assign x_13133 = x_6475 & x_13132;
assign x_13134 = x_6478 & x_6479;
assign x_13135 = x_6480 & x_6481;
assign x_13136 = x_13134 & x_13135;
assign x_13137 = x_13133 & x_13136;
assign x_13138 = x_13131 & x_13137;
assign x_13139 = x_13126 & x_13138;
assign x_13140 = x_6483 & x_6484;
assign x_13141 = x_6482 & x_13140;
assign x_13142 = x_6486 & x_6487;
assign x_13143 = x_6485 & x_13142;
assign x_13144 = x_13141 & x_13143;
assign x_13145 = x_6489 & x_6490;
assign x_13146 = x_6488 & x_13145;
assign x_13147 = x_6491 & x_6492;
assign x_13148 = x_6493 & x_6494;
assign x_13149 = x_13147 & x_13148;
assign x_13150 = x_13146 & x_13149;
assign x_13151 = x_13144 & x_13150;
assign x_13152 = x_6496 & x_6497;
assign x_13153 = x_6495 & x_13152;
assign x_13154 = x_6499 & x_6500;
assign x_13155 = x_6498 & x_13154;
assign x_13156 = x_13153 & x_13155;
assign x_13157 = x_6502 & x_6503;
assign x_13158 = x_6501 & x_13157;
assign x_13159 = x_6504 & x_6505;
assign x_13160 = x_6506 & x_6507;
assign x_13161 = x_13159 & x_13160;
assign x_13162 = x_13158 & x_13161;
assign x_13163 = x_13156 & x_13162;
assign x_13164 = x_13151 & x_13163;
assign x_13165 = x_13139 & x_13164;
assign x_13166 = x_6509 & x_6510;
assign x_13167 = x_6508 & x_13166;
assign x_13168 = x_6512 & x_6513;
assign x_13169 = x_6511 & x_13168;
assign x_13170 = x_13167 & x_13169;
assign x_13171 = x_6515 & x_6516;
assign x_13172 = x_6514 & x_13171;
assign x_13173 = x_6517 & x_6518;
assign x_13174 = x_6519 & x_6520;
assign x_13175 = x_13173 & x_13174;
assign x_13176 = x_13172 & x_13175;
assign x_13177 = x_13170 & x_13176;
assign x_13178 = x_6522 & x_6523;
assign x_13179 = x_6521 & x_13178;
assign x_13180 = x_6525 & x_6526;
assign x_13181 = x_6524 & x_13180;
assign x_13182 = x_13179 & x_13181;
assign x_13183 = x_6528 & x_6529;
assign x_13184 = x_6527 & x_13183;
assign x_13185 = x_6530 & x_6531;
assign x_13186 = x_6532 & x_6533;
assign x_13187 = x_13185 & x_13186;
assign x_13188 = x_13184 & x_13187;
assign x_13189 = x_13182 & x_13188;
assign x_13190 = x_13177 & x_13189;
assign x_13191 = x_6535 & x_6536;
assign x_13192 = x_6534 & x_13191;
assign x_13193 = x_6538 & x_6539;
assign x_13194 = x_6537 & x_13193;
assign x_13195 = x_13192 & x_13194;
assign x_13196 = x_6541 & x_6542;
assign x_13197 = x_6540 & x_13196;
assign x_13198 = x_6543 & x_6544;
assign x_13199 = x_6545 & x_6546;
assign x_13200 = x_13198 & x_13199;
assign x_13201 = x_13197 & x_13200;
assign x_13202 = x_13195 & x_13201;
assign x_13203 = x_6548 & x_6549;
assign x_13204 = x_6547 & x_13203;
assign x_13205 = x_6551 & x_6552;
assign x_13206 = x_6550 & x_13205;
assign x_13207 = x_13204 & x_13206;
assign x_13208 = x_6554 & x_6555;
assign x_13209 = x_6553 & x_13208;
assign x_13210 = x_6556 & x_6557;
assign x_13211 = x_6558 & x_6559;
assign x_13212 = x_13210 & x_13211;
assign x_13213 = x_13209 & x_13212;
assign x_13214 = x_13207 & x_13213;
assign x_13215 = x_13202 & x_13214;
assign x_13216 = x_13190 & x_13215;
assign x_13217 = x_13165 & x_13216;
assign x_13218 = x_6561 & x_6562;
assign x_13219 = x_6560 & x_13218;
assign x_13220 = x_6564 & x_6565;
assign x_13221 = x_6563 & x_13220;
assign x_13222 = x_13219 & x_13221;
assign x_13223 = x_6567 & x_6568;
assign x_13224 = x_6566 & x_13223;
assign x_13225 = x_6569 & x_6570;
assign x_13226 = x_6571 & x_6572;
assign x_13227 = x_13225 & x_13226;
assign x_13228 = x_13224 & x_13227;
assign x_13229 = x_13222 & x_13228;
assign x_13230 = x_6574 & x_6575;
assign x_13231 = x_6573 & x_13230;
assign x_13232 = x_6577 & x_6578;
assign x_13233 = x_6576 & x_13232;
assign x_13234 = x_13231 & x_13233;
assign x_13235 = x_6580 & x_6581;
assign x_13236 = x_6579 & x_13235;
assign x_13237 = x_6582 & x_6583;
assign x_13238 = x_6584 & x_6585;
assign x_13239 = x_13237 & x_13238;
assign x_13240 = x_13236 & x_13239;
assign x_13241 = x_13234 & x_13240;
assign x_13242 = x_13229 & x_13241;
assign x_13243 = x_6587 & x_6588;
assign x_13244 = x_6586 & x_13243;
assign x_13245 = x_6590 & x_6591;
assign x_13246 = x_6589 & x_13245;
assign x_13247 = x_13244 & x_13246;
assign x_13248 = x_6593 & x_6594;
assign x_13249 = x_6592 & x_13248;
assign x_13250 = x_6595 & x_6596;
assign x_13251 = x_6597 & x_6598;
assign x_13252 = x_13250 & x_13251;
assign x_13253 = x_13249 & x_13252;
assign x_13254 = x_13247 & x_13253;
assign x_13255 = x_6600 & x_6601;
assign x_13256 = x_6599 & x_13255;
assign x_13257 = x_6603 & x_6604;
assign x_13258 = x_6602 & x_13257;
assign x_13259 = x_13256 & x_13258;
assign x_13260 = x_6606 & x_6607;
assign x_13261 = x_6605 & x_13260;
assign x_13262 = x_6608 & x_6609;
assign x_13263 = x_6610 & x_6611;
assign x_13264 = x_13262 & x_13263;
assign x_13265 = x_13261 & x_13264;
assign x_13266 = x_13259 & x_13265;
assign x_13267 = x_13254 & x_13266;
assign x_13268 = x_13242 & x_13267;
assign x_13269 = x_6613 & x_6614;
assign x_13270 = x_6612 & x_13269;
assign x_13271 = x_6616 & x_6617;
assign x_13272 = x_6615 & x_13271;
assign x_13273 = x_13270 & x_13272;
assign x_13274 = x_6619 & x_6620;
assign x_13275 = x_6618 & x_13274;
assign x_13276 = x_6621 & x_6622;
assign x_13277 = x_6623 & x_6624;
assign x_13278 = x_13276 & x_13277;
assign x_13279 = x_13275 & x_13278;
assign x_13280 = x_13273 & x_13279;
assign x_13281 = x_6626 & x_6627;
assign x_13282 = x_6625 & x_13281;
assign x_13283 = x_6629 & x_6630;
assign x_13284 = x_6628 & x_13283;
assign x_13285 = x_13282 & x_13284;
assign x_13286 = x_6632 & x_6633;
assign x_13287 = x_6631 & x_13286;
assign x_13288 = x_6634 & x_6635;
assign x_13289 = x_6636 & x_6637;
assign x_13290 = x_13288 & x_13289;
assign x_13291 = x_13287 & x_13290;
assign x_13292 = x_13285 & x_13291;
assign x_13293 = x_13280 & x_13292;
assign x_13294 = x_6639 & x_6640;
assign x_13295 = x_6638 & x_13294;
assign x_13296 = x_6642 & x_6643;
assign x_13297 = x_6641 & x_13296;
assign x_13298 = x_13295 & x_13297;
assign x_13299 = x_6645 & x_6646;
assign x_13300 = x_6644 & x_13299;
assign x_13301 = x_6647 & x_6648;
assign x_13302 = x_6649 & x_6650;
assign x_13303 = x_13301 & x_13302;
assign x_13304 = x_13300 & x_13303;
assign x_13305 = x_13298 & x_13304;
assign x_13306 = x_6652 & x_6653;
assign x_13307 = x_6651 & x_13306;
assign x_13308 = x_6654 & x_6655;
assign x_13309 = x_6656 & x_6657;
assign x_13310 = x_13308 & x_13309;
assign x_13311 = x_13307 & x_13310;
assign x_13312 = x_6659 & x_6660;
assign x_13313 = x_6658 & x_13312;
assign x_13314 = x_6661 & x_6662;
assign x_13315 = x_6663 & x_6664;
assign x_13316 = x_13314 & x_13315;
assign x_13317 = x_13313 & x_13316;
assign x_13318 = x_13311 & x_13317;
assign x_13319 = x_13305 & x_13318;
assign x_13320 = x_13293 & x_13319;
assign x_13321 = x_13268 & x_13320;
assign x_13322 = x_13217 & x_13321;
assign x_13323 = x_13114 & x_13322;
assign x_13324 = x_12907 & x_13323;
assign x_13325 = x_12492 & x_13324;
assign x_13326 = x_11660 & x_13325;
assign x_13327 = x_9995 & x_13326;
assign o_1 = x_13327;
endmodule
