// Benchmark "SKOLEMFORMULA" written by ABC on Wed May 18 01:46:03 2022

module SKOLEMFORMULA ( 
    i0, i1,
    i2, i3  );
  input  i0, i1;
  output i2, i3;
  assign i3 = ~i0;
  assign i2 = i0;
endmodule


