// Benchmark "SKOLEMFORMULA" written by ABC on Sun May 22 03:09:21 2022

module SKOLEMFORMULA ( 
    i0,
    i1  );
  input  i0;
  output i1;
  assign i1 = 1'b1;
endmodule


