// Benchmark "SKOLEMFORMULA" written by ABC on Fri May 20 21:06:53 2022

module SKOLEMFORMULA ( 
    i0,
    i1, i2  );
  input  i0;
  output i1, i2;
  assign i2 = 1'b1;
  assign i1 = i0;
endmodule


