module formula(x_0,i_1,i_2,i_3,x_4,x_5,x_6,i_7,i_8,i_9,i_10,i_11,i_12,out);
	input x_0;
	input i_1;
	input i_2;
	input i_3;
	input x_4;
	input x_5;
	input x_6;
	input i_7;
	input i_8;
	input i_9;
	input i_10;
	input i_11;
	input i_12;
	wire c1;
	wire carry1;
	wire c2;
	wire carry2;
	wire a1;
	wire a2;
	wire a3;
	wire c3;
	wire a4;
	wire c4;
	wire a5;
	wire c5;
	wire a6;
	wire c6;
	wire a7;
	output out;
	assign c1 = (x_0 ^ x_5);
	assign carry1 = (x_0 & x_5);
	assign c3 = ~i_9;
	assign c5 = (x_4 & i_10);
	assign c6 = (x_5 | i_11);
	assign c4 = (x_0 | i_12);
	assign a1 = ~((c1 ^ i_7));
	assign c2 = (((carry1 ^ x_4)) ^ x_6);
	assign carry2 = (((x_4 & x_6)) | ((carry1 & ((x_4 ^ x_6)))));
	assign a4 = ~((c3 ^ i_1));
	assign a6 = ~((i_11 ^ c5));
	assign a7 = ~((i_12 ^ c6));
	assign a5 = ~((i_10 ^ c4));
	assign a2 = ~((c2 ^ i_8));
	assign a3 = ~((carry2 ^ i_3));
	assign out = (((((((((((a1 & a2)) & a3)) & a4)) & a5)) & a6)) & a7);
endmodule
