// Benchmark "SKOLEMFORMULA" written by ABC on Wed May 18 12:51:36 2022

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5,
    i6, i7, i8, i9, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i20,
    i21, i22, i23, i24, i25, i26, i27, i28, i29, i30, i31  );
  input  i0, i1, i2, i3, i4, i5;
  output i6, i7, i8, i9, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19,
    i20, i21, i22, i23, i24, i25, i26, i27, i28, i29, i30, i31;
  wire n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
    n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
    n62, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
    n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
    n91, n92, n93, n94, n96, n97, n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n116, n117,
    n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
    n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n146, n147, n148, n149, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
    n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n183, n184, n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
    n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
    n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260, n261, n262, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n373, n374, n375, n376, n377, n378,
    n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n407, n408, n409, n410, n411, n412, n413, n414, n415,
    n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
    n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
    n440, n441, n442, n443, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n485, n486, n487, n488, n489,
    n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508, n510, n511, n512, n513, n514,
    n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n600, n601,
    n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620, n621, n622, n624, n625, n626,
    n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
    n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788;
  assign n34 = ~i2 & ~i3;
  assign n35 = ~i2 & i3;
  assign n36 = ~i5 & n35;
  assign n37 = ~i4 & n36;
  assign n38 = ~i1 & n37;
  assign n39 = ~n34 & ~n38;
  assign n40 = i4 & n36;
  assign n41 = n39 & ~n40;
  assign n42 = i5 & n35;
  assign n43 = i4 & n42;
  assign n44 = ~i1 & n43;
  assign n45 = n41 & ~n44;
  assign n46 = ~i1 & i2;
  assign n47 = ~i3 & n46;
  assign n48 = ~i5 & n47;
  assign n49 = n45 & ~n48;
  assign n50 = i5 & n47;
  assign n51 = ~i4 & n50;
  assign n52 = i0 & n51;
  assign n53 = n49 & ~n52;
  assign n54 = i1 & i2;
  assign n55 = ~i5 & n54;
  assign n56 = ~i3 & n55;
  assign n57 = n53 & ~n56;
  assign n58 = i5 & n54;
  assign n59 = ~i4 & n58;
  assign n60 = ~i0 & n59;
  assign n61 = n57 & ~n60;
  assign n62 = i4 & n58;
  assign i29 = ~n61 | n62;
  assign n64 = ~i3 & ~i4;
  assign n65 = ~i3 & i4;
  assign n66 = ~i1 & n65;
  assign n67 = ~n64 & ~n66;
  assign n68 = i1 & n65;
  assign n69 = i29 & n68;
  assign n70 = i2 & n69;
  assign n71 = n67 & ~n70;
  assign n72 = i3 & ~i5;
  assign n73 = ~i2 & n72;
  assign n74 = i4 & n73;
  assign n75 = i0 & n74;
  assign n76 = n71 & ~n75;
  assign n77 = i2 & n72;
  assign n78 = ~i29 & n77;
  assign n79 = n76 & ~n78;
  assign n80 = i29 & n77;
  assign n81 = i0 & n80;
  assign n82 = n79 & ~n81;
  assign n83 = i3 & i5;
  assign n84 = ~i2 & n83;
  assign n85 = n82 & ~n84;
  assign n86 = i2 & n83;
  assign n87 = ~i1 & n86;
  assign n88 = ~i0 & n87;
  assign n89 = n85 & ~n88;
  assign n90 = i0 & n87;
  assign n91 = i29 & n90;
  assign n92 = n89 & ~n91;
  assign n93 = i1 & n86;
  assign n94 = i0 & n93;
  assign i28 = ~n92 | n94;
  assign n96 = ~i5 & i29;
  assign n97 = ~i0 & n96;
  assign n98 = ~i4 & n97;
  assign n99 = ~i2 & n98;
  assign n100 = i2 & n98;
  assign n101 = ~n99 & ~n100;
  assign n102 = i4 & n97;
  assign n103 = ~i2 & n102;
  assign n104 = ~i3 & n103;
  assign n105 = n101 & ~n104;
  assign n106 = i0 & n96;
  assign n107 = n105 & ~n106;
  assign n108 = ~i0 & i5;
  assign n109 = n107 & ~n108;
  assign n110 = i0 & i5;
  assign n111 = ~i2 & n110;
  assign n112 = ~i29 & n111;
  assign n113 = n109 & ~n112;
  assign n114 = i2 & n110;
  assign i27 = ~n113 | n114;
  assign n116 = n108 & i27;
  assign n117 = ~i0 & ~i5;
  assign n118 = ~i27 & n117;
  assign n119 = i27 & n117;
  assign n120 = ~i1 & n119;
  assign n121 = ~i4 & n120;
  assign n122 = ~n118 & ~n121;
  assign n123 = i4 & n120;
  assign n124 = n122 & ~n123;
  assign n125 = i1 & n119;
  assign n126 = ~i2 & n125;
  assign n127 = i4 & n126;
  assign n128 = n124 & ~n127;
  assign n129 = n108 & ~i27;
  assign n130 = ~i3 & n129;
  assign n131 = n128 & ~n130;
  assign n132 = ~n116 & n131;
  assign n133 = i0 & ~i1;
  assign n134 = i2 & n133;
  assign n135 = ~i29 & n134;
  assign n136 = n132 & ~n135;
  assign n137 = i29 & n134;
  assign n138 = ~i3 & n137;
  assign n139 = i4 & n138;
  assign n140 = n136 & ~n139;
  assign n141 = i0 & i1;
  assign n142 = ~i28 & n141;
  assign n143 = n140 & ~n142;
  assign n144 = i28 & n141;
  assign n145 = ~i3 & n144;
  assign n146 = i27 & n145;
  assign n147 = i2 & n146;
  assign n148 = n143 & ~n147;
  assign n149 = i3 & n144;
  assign i26 = ~n148 | n149;
  assign n151 = ~i1 & ~i4;
  assign n152 = ~i27 & n151;
  assign n153 = i2 & n152;
  assign n154 = i27 & n151;
  assign n155 = i5 & n154;
  assign n156 = ~i29 & n155;
  assign n157 = ~i3 & n156;
  assign n158 = ~n153 & ~n157;
  assign n159 = i3 & n156;
  assign n160 = i0 & n159;
  assign n161 = n158 & ~n160;
  assign n162 = i1 & ~i4;
  assign n163 = ~i0 & n162;
  assign n164 = i26 & n163;
  assign n165 = ~i3 & n164;
  assign n166 = i2 & n165;
  assign n167 = n161 & ~n166;
  assign n168 = i3 & n164;
  assign n169 = n167 & ~n168;
  assign n170 = i0 & n162;
  assign n171 = n169 & ~n170;
  assign n172 = i4 & ~i5;
  assign n173 = ~i29 & n172;
  assign n174 = n171 & ~n173;
  assign n175 = i29 & n172;
  assign n176 = ~i2 & n175;
  assign n177 = n174 & ~n176;
  assign n178 = i2 & n175;
  assign n179 = ~i26 & n178;
  assign n180 = n177 & ~n179;
  assign n181 = i4 & i5;
  assign i25 = ~n180 | n181;
  assign n183 = ~i4 & ~i27;
  assign n184 = ~i4 & i27;
  assign n185 = ~i3 & n184;
  assign n186 = ~i26 & n185;
  assign n187 = ~n183 & ~n186;
  assign n188 = i26 & n185;
  assign n189 = i2 & n188;
  assign n190 = ~i0 & n189;
  assign n191 = n187 & ~n190;
  assign n192 = i3 & n184;
  assign n193 = i2 & n192;
  assign n194 = ~i0 & n193;
  assign n195 = n191 & ~n194;
  assign n196 = i4 & ~i25;
  assign n197 = n195 & ~n196;
  assign n198 = i4 & i25;
  assign n199 = ~i27 & n198;
  assign n200 = i0 & n199;
  assign n201 = ~i2 & n200;
  assign n202 = n197 & ~n201;
  assign n203 = i27 & n198;
  assign n204 = ~i26 & n203;
  assign n205 = n202 & ~n204;
  assign n206 = i26 & n203;
  assign n207 = ~i1 & n206;
  assign n208 = ~i5 & n207;
  assign n209 = n205 & ~n208;
  assign n210 = i5 & n207;
  assign n211 = i2 & n210;
  assign n212 = ~i3 & n211;
  assign n213 = n209 & ~n212;
  assign n214 = i1 & n206;
  assign n215 = i3 & n214;
  assign i24 = ~n213 | n215;
  assign n217 = ~i29 & i26;
  assign n218 = i3 & n217;
  assign n219 = ~i29 & ~i26;
  assign n220 = ~i4 & n219;
  assign n221 = ~i2 & n220;
  assign n222 = ~i0 & n221;
  assign n223 = i2 & n220;
  assign n224 = ~n222 & ~n223;
  assign n225 = ~i3 & n217;
  assign n226 = ~i5 & n225;
  assign n227 = n224 & ~n226;
  assign n228 = i5 & n225;
  assign n229 = i24 & n228;
  assign n230 = ~i4 & n229;
  assign n231 = n227 & ~n230;
  assign n232 = ~n218 & n231;
  assign n233 = ~i2 & i29;
  assign n234 = n232 & ~n233;
  assign n235 = i2 & i29;
  assign n236 = ~i25 & n235;
  assign n237 = ~i4 & n236;
  assign n238 = i0 & n237;
  assign n239 = n234 & ~n238;
  assign n240 = i4 & n236;
  assign n241 = n239 & ~n240;
  assign n242 = i25 & n235;
  assign i22 = ~n241 | n242;
  assign n244 = ~i1 & i4;
  assign n245 = ~i29 & n244;
  assign n246 = ~i27 & n245;
  assign n247 = i4 & ~n246;
  assign n248 = i29 & n244;
  assign n249 = ~i0 & n248;
  assign n250 = ~i28 & n249;
  assign n251 = n247 & ~n250;
  assign n252 = i0 & n248;
  assign n253 = n251 & ~n252;
  assign n254 = i1 & i4;
  assign n255 = ~i2 & n254;
  assign n256 = i22 & n255;
  assign n257 = ~i5 & n256;
  assign n258 = ~i28 & n257;
  assign n259 = n253 & ~n258;
  assign n260 = i5 & n256;
  assign n261 = n259 & ~n260;
  assign n262 = i2 & n254;
  assign i21 = ~n261 | n262;
  assign n264 = ~i4 & ~i24;
  assign n265 = ~i1 & n264;
  assign n266 = i28 & n265;
  assign n267 = i4 & ~i24;
  assign n268 = ~n266 & ~n267;
  assign n269 = ~i4 & i24;
  assign n270 = ~i5 & n269;
  assign n271 = n268 & ~n270;
  assign n272 = i5 & n269;
  assign n273 = ~i2 & n272;
  assign n274 = n271 & ~n273;
  assign n275 = i2 & n272;
  assign n276 = ~i25 & n275;
  assign n277 = n274 & ~n276;
  assign n278 = i4 & i24;
  assign n279 = ~i3 & n278;
  assign n280 = i27 & n279;
  assign n281 = ~i2 & n280;
  assign n282 = ~i1 & n281;
  assign n283 = n277 & ~n282;
  assign n284 = i2 & n280;
  assign n285 = n283 & ~n284;
  assign n286 = i3 & n278;
  assign n287 = i1 & n286;
  assign n288 = ~i28 & n287;
  assign i23 = ~n285 | n288;
  assign n290 = ~i2 & i23;
  assign n291 = ~i2 & ~i23;
  assign n292 = i27 & n291;
  assign n293 = i29 & n292;
  assign n294 = ~n290 & ~n293;
  assign n295 = i2 & ~i29;
  assign n296 = ~i5 & n295;
  assign n297 = ~i23 & n296;
  assign n298 = i3 & n297;
  assign n299 = n294 & ~n298;
  assign n300 = i5 & n295;
  assign n301 = ~i4 & n300;
  assign n302 = n299 & ~n301;
  assign n303 = i4 & n300;
  assign n304 = i22 & n303;
  assign n305 = n302 & ~n304;
  assign n306 = ~i28 & n235;
  assign n307 = i1 & n306;
  assign n308 = n305 & ~n307;
  assign n309 = i28 & n235;
  assign n310 = ~i5 & n309;
  assign i20 = ~n308 | n310;
  assign n312 = i3 & ~i26;
  assign n313 = ~i3 & ~i26;
  assign n314 = ~i1 & n313;
  assign n315 = i20 & n314;
  assign n316 = i1 & n313;
  assign n317 = ~i25 & n316;
  assign n318 = i22 & n317;
  assign n319 = ~n315 & ~n318;
  assign n320 = i25 & n316;
  assign n321 = n319 & ~n320;
  assign n322 = ~n312 & n321;
  assign n323 = ~i0 & i26;
  assign n324 = ~i25 & n323;
  assign n325 = n322 & ~n324;
  assign n326 = i25 & n323;
  assign n327 = ~i2 & n326;
  assign n328 = ~i5 & n327;
  assign n329 = i4 & n328;
  assign n330 = n325 & ~n329;
  assign n331 = i2 & n326;
  assign n332 = i21 & n331;
  assign n333 = n330 & ~n332;
  assign n334 = i0 & i26;
  assign n335 = ~i3 & n334;
  assign n336 = i21 & n335;
  assign n337 = ~i24 & n336;
  assign n338 = ~i23 & n337;
  assign n339 = n333 & ~n338;
  assign n340 = i24 & n336;
  assign n341 = n339 & ~n340;
  assign n342 = i3 & n334;
  assign i19 = ~n341 | n342;
  assign n344 = i28 & ~i27;
  assign n345 = ~i21 & n344;
  assign n346 = i28 & ~n345;
  assign n347 = i21 & n344;
  assign n348 = ~i29 & n347;
  assign n349 = ~i3 & n348;
  assign n350 = ~i20 & n349;
  assign n351 = ~i23 & n350;
  assign n352 = n346 & ~n351;
  assign n353 = i29 & n347;
  assign n354 = i25 & n353;
  assign n355 = n352 & ~n354;
  assign n356 = i28 & i27;
  assign n357 = ~i19 & n356;
  assign n358 = ~i29 & n357;
  assign n359 = n355 & ~n358;
  assign n360 = i29 & n357;
  assign n361 = ~i5 & n360;
  assign n362 = i0 & n361;
  assign n363 = n359 & ~n362;
  assign n364 = i19 & n356;
  assign n365 = ~i23 & n364;
  assign n366 = ~i2 & n365;
  assign n367 = ~i25 & n366;
  assign n368 = n363 & ~n367;
  assign n369 = i2 & n365;
  assign n370 = n368 & ~n369;
  assign n371 = i23 & n364;
  assign i18 = ~n370 | n371;
  assign n373 = i26 & ~i22;
  assign n374 = ~i26 & ~i18;
  assign n375 = ~i2 & n374;
  assign n376 = ~i25 & n375;
  assign n377 = ~i26 & i18;
  assign n378 = ~i5 & n377;
  assign n379 = ~i23 & n378;
  assign n380 = ~n376 & ~n379;
  assign n381 = i23 & n378;
  assign n382 = i21 & n381;
  assign n383 = n380 & ~n382;
  assign n384 = i5 & n377;
  assign n385 = n383 & ~n384;
  assign n386 = ~n373 & n385;
  assign n387 = i26 & i22;
  assign n388 = ~i2 & n387;
  assign n389 = ~i5 & n388;
  assign n390 = n386 & ~n389;
  assign n391 = i5 & n388;
  assign n392 = n390 & ~n391;
  assign n393 = i2 & n387;
  assign n394 = ~i27 & n393;
  assign n395 = ~i18 & n394;
  assign n396 = i1 & n395;
  assign n397 = n392 & ~n396;
  assign n398 = i18 & n394;
  assign n399 = n397 & ~n398;
  assign n400 = i27 & n393;
  assign n401 = ~i19 & n400;
  assign n402 = ~i18 & n401;
  assign n403 = n399 & ~n402;
  assign n404 = i19 & n400;
  assign n405 = i23 & n404;
  assign i17 = ~n403 | n405;
  assign n407 = ~i4 & ~i29;
  assign n408 = ~i19 & n407;
  assign n409 = i19 & n407;
  assign n410 = i2 & n409;
  assign n411 = ~i26 & n410;
  assign n412 = ~n408 & ~n411;
  assign n413 = i26 & n410;
  assign n414 = i20 & n413;
  assign n415 = i17 & n414;
  assign n416 = n412 & ~n415;
  assign n417 = ~i4 & i29;
  assign n418 = ~i17 & n417;
  assign n419 = n416 & ~n418;
  assign n420 = i17 & n417;
  assign n421 = ~i2 & n420;
  assign n422 = i28 & n421;
  assign n423 = n419 & ~n422;
  assign n424 = i2 & n420;
  assign n425 = ~i18 & n424;
  assign n426 = n423 & ~n425;
  assign n427 = i4 & ~i28;
  assign n428 = n426 & ~n427;
  assign n429 = i4 & i28;
  assign n430 = ~i25 & n429;
  assign n431 = n428 & ~n430;
  assign n432 = i25 & n429;
  assign n433 = ~i17 & n432;
  assign n434 = n431 & ~n433;
  assign n435 = i17 & n432;
  assign n436 = ~i20 & n435;
  assign n437 = ~i21 & n436;
  assign n438 = i19 & n437;
  assign n439 = n434 & ~n438;
  assign n440 = i21 & n436;
  assign n441 = n439 & ~n440;
  assign n442 = i20 & n435;
  assign n443 = ~i19 & n442;
  assign i16 = ~n441 | n443;
  assign n445 = ~i2 & ~i18;
  assign n446 = ~i0 & n445;
  assign n447 = ~i24 & n446;
  assign n448 = i21 & n447;
  assign n449 = i0 & n445;
  assign n450 = ~n448 & ~n449;
  assign n451 = ~i2 & i18;
  assign n452 = ~i26 & n451;
  assign n453 = ~i24 & n452;
  assign n454 = n450 & ~n453;
  assign n455 = i24 & n452;
  assign n456 = ~i17 & n455;
  assign n457 = n454 & ~n456;
  assign n458 = i17 & n455;
  assign n459 = ~i19 & n458;
  assign n460 = n457 & ~n459;
  assign n461 = i26 & n451;
  assign n462 = n460 & ~n461;
  assign n463 = i2 & ~i26;
  assign n464 = ~i5 & n463;
  assign n465 = n462 & ~n464;
  assign n466 = i5 & n463;
  assign n467 = ~i0 & n466;
  assign n468 = n465 & ~n467;
  assign n469 = i2 & i26;
  assign n470 = ~i16 & n469;
  assign n471 = ~i1 & n470;
  assign n472 = n468 & ~n471;
  assign n473 = i16 & n469;
  assign n474 = ~i19 & n473;
  assign n475 = ~i25 & n474;
  assign n476 = n472 & ~n475;
  assign n477 = i25 & n474;
  assign n478 = ~i20 & n477;
  assign n479 = ~i3 & n478;
  assign n480 = n476 & ~n479;
  assign n481 = i19 & n473;
  assign n482 = ~i4 & n481;
  assign n483 = ~i0 & n482;
  assign i15 = ~n480 | n483;
  assign n485 = ~i5 & ~i15;
  assign n486 = i16 & n485;
  assign n487 = ~i16 & n485;
  assign n488 = ~i19 & n487;
  assign n489 = ~n486 & ~n488;
  assign n490 = i5 & ~i15;
  assign n491 = ~i22 & n490;
  assign n492 = ~i4 & n491;
  assign n493 = n489 & ~n492;
  assign n494 = i22 & n490;
  assign n495 = ~i24 & n494;
  assign n496 = ~i19 & n495;
  assign n497 = n493 & ~n496;
  assign n498 = ~i1 & i15;
  assign n499 = n497 & ~n498;
  assign n500 = i1 & i15;
  assign n501 = ~i29 & n500;
  assign n502 = ~i27 & n501;
  assign n503 = n499 & ~n502;
  assign n504 = i29 & n500;
  assign n505 = ~i25 & n504;
  assign n506 = ~i5 & n505;
  assign n507 = n503 & ~n506;
  assign n508 = i25 & n504;
  assign i14 = ~n507 | n508;
  assign n510 = ~i0 & ~i21;
  assign n511 = i5 & n510;
  assign n512 = ~i4 & n511;
  assign n513 = i4 & n511;
  assign n514 = i18 & n513;
  assign n515 = ~n512 & ~n514;
  assign n516 = ~i0 & i21;
  assign n517 = ~i5 & n516;
  assign n518 = n515 & ~n517;
  assign n519 = i5 & n516;
  assign n520 = ~i25 & n519;
  assign n521 = i29 & n520;
  assign n522 = n518 & ~n521;
  assign n523 = i25 & n519;
  assign n524 = n522 & ~n523;
  assign n525 = i0 & ~i22;
  assign n526 = ~i14 & n525;
  assign n527 = n524 & ~n526;
  assign n528 = i0 & i22;
  assign n529 = ~i4 & n528;
  assign n530 = i27 & n529;
  assign n531 = i28 & n530;
  assign n532 = n527 & ~n531;
  assign n533 = i4 & n528;
  assign i13 = ~n532 | n533;
  assign n535 = ~i28 & ~i13;
  assign n536 = i28 & ~i13;
  assign n537 = ~i21 & n536;
  assign n538 = i20 & n537;
  assign n539 = ~n535 & ~n538;
  assign n540 = i21 & n536;
  assign n541 = ~i23 & n540;
  assign n542 = ~i22 & n541;
  assign n543 = n539 & ~n542;
  assign n544 = ~i21 & i13;
  assign n545 = i26 & n544;
  assign n546 = i15 & n545;
  assign n547 = n543 & ~n546;
  assign n548 = i21 & i13;
  assign n549 = ~i17 & n548;
  assign n550 = n547 & ~n549;
  assign n551 = i17 & n548;
  assign n552 = ~i29 & n551;
  assign n553 = ~i22 & n552;
  assign n554 = i16 & n553;
  assign n555 = n550 & ~n554;
  assign n556 = i22 & n552;
  assign n557 = n555 & ~n556;
  assign n558 = i29 & n551;
  assign n559 = ~i27 & n558;
  assign n560 = n557 & ~n559;
  assign n561 = i27 & n558;
  assign n562 = i1 & n561;
  assign n563 = i22 & n562;
  assign n564 = i26 & n563;
  assign i10 = ~n560 | n564;
  assign n566 = ~i2 & ~i28;
  assign n567 = ~i25 & n566;
  assign n568 = i25 & n566;
  assign n569 = ~i5 & n568;
  assign n570 = ~i10 & n569;
  assign n571 = i21 & n570;
  assign n572 = ~n567 & ~n571;
  assign n573 = i5 & n568;
  assign n574 = n572 & ~n573;
  assign n575 = ~i2 & i28;
  assign n576 = ~i22 & n575;
  assign n577 = ~i1 & n576;
  assign n578 = n574 & ~n577;
  assign n579 = i22 & n575;
  assign n580 = n578 & ~n579;
  assign n581 = ~i0 & n295;
  assign n582 = ~i16 & n581;
  assign n583 = i14 & n582;
  assign n584 = ~i27 & n583;
  assign n585 = n580 & ~n584;
  assign n586 = i16 & n581;
  assign n587 = n585 & ~n586;
  assign n588 = i0 & n295;
  assign n589 = ~i14 & n588;
  assign n590 = n587 & ~n589;
  assign n591 = ~i4 & n235;
  assign n592 = n590 & ~n591;
  assign n593 = i4 & n235;
  assign n594 = ~i26 & n593;
  assign n595 = n592 & ~n594;
  assign n596 = i26 & n593;
  assign n597 = i28 & n596;
  assign n598 = i5 & n597;
  assign i11 = ~n595 | n598;
  assign n600 = ~i25 & n407;
  assign n601 = i27 & n600;
  assign n602 = i25 & n407;
  assign n603 = ~n601 & ~n602;
  assign n604 = ~i1 & n417;
  assign n605 = ~i27 & n604;
  assign n606 = i13 & n605;
  assign n607 = n603 & ~n606;
  assign n608 = i27 & n604;
  assign n609 = n607 & ~n608;
  assign n610 = i1 & n417;
  assign n611 = ~i18 & n610;
  assign n612 = n609 & ~n611;
  assign n613 = i18 & n610;
  assign n614 = ~i11 & n613;
  assign n615 = n612 & ~n614;
  assign n616 = i4 & ~i20;
  assign n617 = ~i5 & n616;
  assign n618 = ~i26 & n617;
  assign n619 = n615 & ~n618;
  assign n620 = i5 & n616;
  assign n621 = n619 & ~n620;
  assign n622 = i4 & i20;
  assign i7 = ~n621 | n622;
  assign n624 = ~i1 & ~i27;
  assign n625 = ~i20 & n624;
  assign n626 = i18 & n625;
  assign n627 = ~i1 & i27;
  assign n628 = ~i29 & n627;
  assign n629 = ~i21 & n628;
  assign n630 = i14 & n629;
  assign n631 = ~n626 & ~n630;
  assign n632 = i29 & n627;
  assign n633 = ~i2 & n632;
  assign n634 = i11 & n633;
  assign n635 = ~i10 & n634;
  assign n636 = i5 & n635;
  assign n637 = n631 & ~n636;
  assign n638 = i10 & n634;
  assign n639 = n637 & ~n638;
  assign n640 = i2 & n632;
  assign n641 = n639 & ~n640;
  assign n642 = i1 & ~i17;
  assign n643 = ~i26 & n642;
  assign n644 = ~i7 & n643;
  assign n645 = n641 & ~n644;
  assign n646 = i26 & n642;
  assign n647 = n645 & ~n646;
  assign n648 = i1 & i17;
  assign n649 = ~i27 & n648;
  assign n650 = ~i24 & n649;
  assign n651 = ~i18 & n650;
  assign n652 = n647 & ~n651;
  assign n653 = i24 & n649;
  assign n654 = n652 & ~n653;
  assign n655 = i27 & n648;
  assign i12 = ~n654 | n655;
  assign n657 = ~i0 & ~i14;
  assign n658 = i4 & n657;
  assign n659 = ~i4 & n657;
  assign n660 = ~i17 & n659;
  assign n661 = ~n658 & ~n660;
  assign n662 = ~i16 & i14;
  assign n663 = n661 & ~n662;
  assign n664 = i16 & i14;
  assign n665 = ~i22 & n664;
  assign n666 = i19 & n665;
  assign n667 = i20 & n666;
  assign n668 = n663 & ~n667;
  assign n669 = i22 & n664;
  assign n670 = ~i1 & n669;
  assign n671 = ~i23 & n670;
  assign n672 = n668 & ~n671;
  assign n673 = i23 & n670;
  assign n674 = n672 & ~n673;
  assign n675 = i1 & n669;
  assign n676 = ~i12 & n675;
  assign n677 = ~i3 & n676;
  assign n678 = n674 & ~n677;
  assign n679 = i12 & n675;
  assign n680 = i21 & n679;
  assign i9 = ~n678 | n680;
  assign n682 = ~i24 & ~i19;
  assign n683 = ~i5 & n682;
  assign n684 = i24 & ~i19;
  assign n685 = ~i23 & n684;
  assign n686 = ~i20 & n685;
  assign n687 = i26 & n686;
  assign n688 = ~n683 & ~n687;
  assign n689 = i23 & n684;
  assign n690 = n688 & ~n689;
  assign n691 = ~i3 & i19;
  assign n692 = ~i5 & n691;
  assign n693 = n690 & ~n692;
  assign n694 = i5 & n691;
  assign n695 = ~i10 & n694;
  assign n696 = n693 & ~n695;
  assign n697 = i10 & n694;
  assign n698 = ~i23 & n697;
  assign n699 = i12 & n698;
  assign n700 = n696 & ~n699;
  assign n701 = i3 & i19;
  assign n702 = ~i13 & n701;
  assign n703 = i5 & n702;
  assign n704 = n700 & ~n703;
  assign n705 = i13 & n701;
  assign i8 = ~n704 | n705;
  assign n707 = ~i0 & i1;
  assign n708 = ~n133 & ~n707;
  assign n709 = i2 & n708;
  assign n710 = ~i2 & ~n708;
  assign n711 = ~n709 & ~n710;
  assign n712 = i3 & n711;
  assign n713 = ~i3 & ~n711;
  assign n714 = ~n712 & ~n713;
  assign n715 = i4 & n714;
  assign n716 = ~i4 & ~n714;
  assign n717 = ~n715 & ~n716;
  assign n718 = i5 & n717;
  assign n719 = ~i5 & ~n717;
  assign n720 = ~n718 & ~n719;
  assign n721 = i7 & ~n720;
  assign n722 = ~i7 & n720;
  assign n723 = ~n721 & ~n722;
  assign n724 = i8 & n723;
  assign n725 = ~i8 & ~n723;
  assign n726 = ~n724 & ~n725;
  assign n727 = i9 & n726;
  assign n728 = ~i9 & ~n726;
  assign n729 = ~n727 & ~n728;
  assign n730 = i10 & n729;
  assign n731 = ~i10 & ~n729;
  assign n732 = ~n730 & ~n731;
  assign n733 = i11 & n732;
  assign n734 = ~i11 & ~n732;
  assign n735 = ~n733 & ~n734;
  assign n736 = i12 & n735;
  assign n737 = ~i12 & ~n735;
  assign n738 = ~n736 & ~n737;
  assign n739 = i13 & n738;
  assign n740 = ~i13 & ~n738;
  assign n741 = ~n739 & ~n740;
  assign n742 = i14 & n741;
  assign n743 = ~i14 & ~n741;
  assign n744 = ~n742 & ~n743;
  assign n745 = i15 & n744;
  assign n746 = ~i15 & ~n744;
  assign n747 = ~n745 & ~n746;
  assign n748 = i16 & n747;
  assign n749 = ~i16 & ~n747;
  assign n750 = ~n748 & ~n749;
  assign n751 = i17 & n750;
  assign n752 = ~i17 & ~n750;
  assign n753 = ~n751 & ~n752;
  assign n754 = i18 & n753;
  assign n755 = ~i18 & ~n753;
  assign n756 = ~n754 & ~n755;
  assign n757 = i19 & n756;
  assign n758 = ~i19 & ~n756;
  assign n759 = ~n757 & ~n758;
  assign n760 = i20 & n759;
  assign n761 = ~i20 & ~n759;
  assign n762 = ~n760 & ~n761;
  assign n763 = i21 & n762;
  assign n764 = ~i21 & ~n762;
  assign n765 = ~n763 & ~n764;
  assign n766 = i22 & n765;
  assign n767 = ~i22 & ~n765;
  assign n768 = ~n766 & ~n767;
  assign n769 = i23 & n768;
  assign n770 = ~i23 & ~n768;
  assign n771 = ~n769 & ~n770;
  assign n772 = i24 & n771;
  assign n773 = ~i24 & ~n771;
  assign n774 = ~n772 & ~n773;
  assign n775 = i25 & n774;
  assign n776 = ~i25 & ~n774;
  assign n777 = ~n775 & ~n776;
  assign n778 = i26 & n777;
  assign n779 = ~i26 & ~n777;
  assign n780 = ~n778 & ~n779;
  assign n781 = i27 & n780;
  assign n782 = ~i27 & ~n780;
  assign n783 = ~n781 & ~n782;
  assign n784 = i28 & n783;
  assign n785 = ~i28 & ~n783;
  assign n786 = ~n784 & ~n785;
  assign n787 = i29 & n786;
  assign n788 = ~i29 & ~n786;
  assign i6 = n787 | n788;
  assign i30 = 1'b1;
  assign i31 = 1'b1;
endmodule


