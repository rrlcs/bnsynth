module formula(v_1,v_2,v_3,v_4,v_5,v_6,v_7,v_8,v_9,v_10,v_11,v_12,v_13,v_14,v_15,v_16,v_17,v_18,v_19,v_20,v_21,v_22,v_23,v_24,v_25,v_26,v_27,v_28,v_29,v_30,v_31,v_32,v_33,v_34,v_35,v_36,v_37,v_38,v_39,v_40,v_41,v_42,v_43,v_44,v_45,v_46,v_47,v_48,v_49,v_50,v_51,v_52,v_53,v_54,v_55,v_56,v_57,v_58,v_59,v_60,v_61,v_62,v_63,v_64,v_65,v_66,v_67,v_68,v_69,v_70,v_71,v_72,v_73,v_74,v_75,v_76,v_77,v_78,v_79,v_80,v_81,v_82,v_83,v_84,v_85,v_86,v_87,v_88,v_89,v_90,v_91,v_92,v_93,v_94,v_95,v_96,v_97,v_98,v_99,v_100,v_101,v_102,v_103,v_104,v_105,v_106,v_107,v_108,v_109,v_110,v_111,v_112,v_113,v_114,v_115,v_116,v_117,v_118,v_119,v_120,v_121,v_122,v_123,v_124,v_125,v_126,v_127,v_128,v_129,v_130,v_131,v_132,v_133,v_134,v_135,v_136,v_137,v_138,v_139,v_140,v_141,v_142,v_143,v_144,v_145,v_146,v_147,v_148,v_149,v_150,v_151,v_152,v_153,v_154,v_155,v_156,v_157,v_158,v_159,v_160,v_161,v_162,v_163,v_164,v_165,v_166,v_167,v_168,v_169,v_170,v_171,v_172,v_173,v_174,v_175,v_176,v_177,v_178,v_179,v_180,v_181,v_182,v_183,v_184,v_185,v_186,v_187,v_188,v_189,v_190,v_191,v_192,v_193,v_194,v_195,v_196,v_197,v_198,v_199,v_200,v_201,v_202,v_203,v_204,v_205,v_206,v_207,v_208,v_209,v_210,v_211,v_212,v_213,v_214,v_215,v_216,v_217,v_218,v_219,v_220,v_221,v_222,v_223,v_224,v_225,v_226,v_227,v_228,v_229,v_230,v_231,v_232,v_233,v_234,v_235,v_236,v_237,v_238,v_239,v_240,v_241,v_242,v_243,v_244,v_245,v_246,v_247,v_248,v_249,v_250,v_251,v_252,v_253,v_254,v_255,v_256,v_257,v_258,v_259,v_260,v_388,v_982,v_1582,o_1);
	input v_1;
	v_2;
	v_3;
	v_4;
	v_5;
	v_6;
	v_7;
	v_8;
	v_9;
	v_10;
	v_11;
	v_12;
	v_13;
	v_14;
	v_15;
	v_16;
	v_17;
	v_18;
	v_19;
	v_20;
	v_21;
	v_22;
	v_23;
	v_24;
	v_25;
	v_26;
	v_27;
	v_28;
	v_29;
	v_30;
	v_31;
	v_32;
	v_33;
	v_34;
	v_35;
	v_36;
	v_37;
	v_38;
	v_39;
	v_40;
	v_41;
	v_42;
	v_43;
	v_44;
	v_45;
	v_46;
	v_47;
	v_48;
	v_49;
	v_50;
	v_51;
	v_52;
	v_53;
	v_54;
	v_55;
	v_56;
	v_57;
	v_58;
	v_59;
	v_60;
	v_61;
	v_62;
	v_63;
	v_64;
	v_65;
	v_66;
	v_67;
	v_68;
	v_69;
	v_70;
	v_71;
	v_72;
	v_73;
	v_74;
	v_75;
	v_76;
	v_77;
	v_78;
	v_79;
	v_80;
	v_81;
	v_82;
	v_83;
	v_84;
	v_85;
	v_86;
	v_87;
	v_88;
	v_89;
	v_90;
	v_91;
	v_92;
	v_93;
	v_94;
	v_95;
	v_96;
	v_97;
	v_98;
	v_99;
	v_100;
	v_101;
	v_102;
	v_103;
	v_104;
	v_105;
	v_106;
	v_107;
	v_108;
	v_109;
	v_110;
	v_111;
	v_112;
	v_113;
	v_114;
	v_115;
	v_116;
	v_117;
	v_118;
	v_119;
	v_120;
	v_121;
	v_122;
	v_123;
	v_124;
	v_125;
	v_126;
	v_127;
	v_128;
	v_129;
	v_130;
	v_131;
	v_132;
	v_133;
	v_134;
	v_135;
	v_136;
	v_137;
	v_138;
	v_139;
	v_140;
	v_141;
	v_142;
	v_143;
	v_144;
	v_145;
	v_146;
	v_147;
	v_148;
	v_149;
	v_150;
	v_151;
	v_152;
	v_153;
	v_154;
	v_155;
	v_156;
	v_157;
	v_158;
	v_159;
	v_160;
	v_161;
	v_162;
	v_163;
	v_164;
	v_165;
	v_166;
	v_167;
	v_168;
	v_169;
	v_170;
	v_171;
	v_172;
	v_173;
	v_174;
	v_175;
	v_176;
	v_177;
	v_178;
	v_179;
	v_180;
	v_181;
	v_182;
	v_183;
	v_184;
	v_185;
	v_186;
	v_187;
	v_188;
	v_189;
	v_190;
	v_191;
	v_192;
	v_193;
	v_194;
	v_195;
	v_196;
	v_197;
	v_198;
	v_199;
	v_200;
	v_201;
	v_202;
	v_203;
	v_204;
	v_205;
	v_206;
	v_207;
	v_208;
	v_209;
	v_210;
	v_211;
	v_212;
	v_213;
	v_214;
	v_215;
	v_216;
	v_217;
	v_218;
	v_219;
	v_220;
	v_221;
	v_222;
	v_223;
	v_224;
	v_225;
	v_226;
	v_227;
	v_228;
	v_229;
	v_230;
	v_231;
	v_232;
	v_233;
	v_234;
	v_235;
	v_236;
	v_237;
	v_238;
	v_239;
	v_240;
	v_241;
	v_242;
	v_243;
	v_244;
	v_245;
	v_246;
	v_247;
	v_248;
	v_249;
	v_250;
	v_251;
	v_252;
	v_253;
	v_254;
	v_255;
	v_256;
	v_257;
	v_258;
	v_259;
	v_260;
	v_388;
	v_982;
	v_1582;
	wire v_261;
	wire v_262;
	wire v_263;
	wire v_264;
	wire v_265;
	wire v_266;
	wire v_267;
	wire v_268;
	wire v_269;
	wire v_270;
	wire v_271;
	wire v_272;
	wire v_273;
	wire v_274;
	wire v_275;
	wire v_276;
	wire v_277;
	wire v_278;
	wire v_279;
	wire v_280;
	wire v_281;
	wire v_282;
	wire v_283;
	wire v_284;
	wire v_285;
	wire v_286;
	wire v_287;
	wire v_288;
	wire v_289;
	wire v_290;
	wire v_291;
	wire v_292;
	wire v_293;
	wire v_294;
	wire v_295;
	wire v_296;
	wire v_297;
	wire v_298;
	wire v_299;
	wire v_300;
	wire v_301;
	wire v_302;
	wire v_303;
	wire v_304;
	wire v_305;
	wire v_306;
	wire v_307;
	wire v_308;
	wire v_309;
	wire v_310;
	wire v_311;
	wire v_312;
	wire v_313;
	wire v_314;
	wire v_315;
	wire v_316;
	wire v_317;
	wire v_318;
	wire v_319;
	wire v_320;
	wire v_321;
	wire v_322;
	wire v_323;
	wire v_324;
	wire v_325;
	wire v_326;
	wire v_327;
	wire v_328;
	wire v_329;
	wire v_330;
	wire v_331;
	wire v_332;
	wire v_333;
	wire v_334;
	wire v_335;
	wire v_336;
	wire v_337;
	wire v_338;
	wire v_339;
	wire v_340;
	wire v_341;
	wire v_342;
	wire v_343;
	wire v_344;
	wire v_345;
	wire v_346;
	wire v_347;
	wire v_348;
	wire v_349;
	wire v_350;
	wire v_351;
	wire v_352;
	wire v_353;
	wire v_354;
	wire v_355;
	wire v_356;
	wire v_357;
	wire v_358;
	wire v_359;
	wire v_360;
	wire v_361;
	wire v_362;
	wire v_363;
	wire v_364;
	wire v_365;
	wire v_366;
	wire v_367;
	wire v_368;
	wire v_369;
	wire v_370;
	wire v_371;
	wire v_372;
	wire v_373;
	wire v_374;
	wire v_375;
	wire v_376;
	wire v_377;
	wire v_378;
	wire v_379;
	wire v_380;
	wire v_381;
	wire v_382;
	wire v_383;
	wire v_384;
	wire v_385;
	wire v_386;
	wire v_387;
	wire v_389;
	wire v_390;
	wire v_391;
	wire v_392;
	wire v_393;
	wire v_394;
	wire v_395;
	wire v_396;
	wire v_397;
	wire v_398;
	wire v_399;
	wire v_400;
	wire v_401;
	wire v_402;
	wire v_403;
	wire v_404;
	wire v_405;
	wire v_406;
	wire v_407;
	wire v_408;
	wire v_409;
	wire v_410;
	wire v_411;
	wire v_412;
	wire v_413;
	wire v_414;
	wire v_415;
	wire v_416;
	wire v_417;
	wire v_418;
	wire v_419;
	wire v_420;
	wire v_421;
	wire v_422;
	wire v_423;
	wire v_424;
	wire v_425;
	wire v_426;
	wire v_427;
	wire v_428;
	wire v_429;
	wire v_430;
	wire v_431;
	wire v_432;
	wire v_433;
	wire v_434;
	wire v_435;
	wire v_436;
	wire v_437;
	wire v_438;
	wire v_439;
	wire v_440;
	wire v_441;
	wire v_442;
	wire v_443;
	wire v_444;
	wire v_445;
	wire v_446;
	wire v_447;
	wire v_448;
	wire v_449;
	wire v_450;
	wire v_451;
	wire v_452;
	wire v_453;
	wire v_454;
	wire v_455;
	wire v_456;
	wire v_457;
	wire v_458;
	wire v_459;
	wire v_460;
	wire v_461;
	wire v_462;
	wire v_463;
	wire v_464;
	wire v_465;
	wire v_466;
	wire v_467;
	wire v_468;
	wire v_469;
	wire v_470;
	wire v_471;
	wire v_472;
	wire v_473;
	wire v_474;
	wire v_475;
	wire v_476;
	wire v_477;
	wire v_478;
	wire v_479;
	wire v_480;
	wire v_481;
	wire v_482;
	wire v_483;
	wire v_484;
	wire v_485;
	wire v_486;
	wire v_487;
	wire v_488;
	wire v_489;
	wire v_490;
	wire v_491;
	wire v_492;
	wire v_493;
	wire v_494;
	wire v_495;
	wire v_496;
	wire v_497;
	wire v_498;
	wire v_499;
	wire v_500;
	wire v_501;
	wire v_502;
	wire v_503;
	wire v_504;
	wire v_505;
	wire v_506;
	wire v_507;
	wire v_508;
	wire v_509;
	wire v_510;
	wire v_511;
	wire v_512;
	wire v_513;
	wire v_514;
	wire v_515;
	wire v_516;
	wire v_517;
	wire v_518;
	wire v_519;
	wire v_520;
	wire v_521;
	wire v_522;
	wire v_523;
	wire v_524;
	wire v_525;
	wire v_526;
	wire v_527;
	wire v_528;
	wire v_529;
	wire v_530;
	wire v_531;
	wire v_532;
	wire v_533;
	wire v_534;
	wire v_535;
	wire v_536;
	wire v_537;
	wire v_538;
	wire v_539;
	wire v_540;
	wire v_541;
	wire v_542;
	wire v_543;
	wire v_544;
	wire v_545;
	wire v_546;
	wire v_547;
	wire v_548;
	wire v_549;
	wire v_550;
	wire v_551;
	wire v_552;
	wire v_553;
	wire v_554;
	wire v_555;
	wire v_556;
	wire v_557;
	wire v_558;
	wire v_559;
	wire v_560;
	wire v_561;
	wire v_562;
	wire v_563;
	wire v_564;
	wire v_565;
	wire v_566;
	wire v_567;
	wire v_568;
	wire v_569;
	wire v_570;
	wire v_571;
	wire v_572;
	wire v_573;
	wire v_574;
	wire v_575;
	wire v_576;
	wire v_577;
	wire v_578;
	wire v_579;
	wire v_580;
	wire v_581;
	wire v_582;
	wire v_583;
	wire v_584;
	wire v_585;
	wire v_586;
	wire v_587;
	wire v_588;
	wire v_589;
	wire v_590;
	wire v_591;
	wire v_592;
	wire v_593;
	wire v_594;
	wire v_595;
	wire v_596;
	wire v_597;
	wire v_598;
	wire v_599;
	wire v_600;
	wire v_601;
	wire v_602;
	wire v_603;
	wire v_604;
	wire v_605;
	wire v_606;
	wire v_607;
	wire v_608;
	wire v_609;
	wire v_610;
	wire v_611;
	wire v_612;
	wire v_613;
	wire v_614;
	wire v_615;
	wire v_616;
	wire v_617;
	wire v_618;
	wire v_619;
	wire v_620;
	wire v_621;
	wire v_622;
	wire v_623;
	wire v_624;
	wire v_625;
	wire v_626;
	wire v_627;
	wire v_628;
	wire v_629;
	wire v_630;
	wire v_631;
	wire v_632;
	wire v_633;
	wire v_634;
	wire v_635;
	wire v_636;
	wire v_637;
	wire v_638;
	wire v_639;
	wire v_640;
	wire v_641;
	wire v_642;
	wire v_643;
	wire v_644;
	wire v_645;
	wire v_646;
	wire v_647;
	wire v_648;
	wire v_649;
	wire v_650;
	wire v_651;
	wire v_652;
	wire v_653;
	wire v_654;
	wire v_655;
	wire v_656;
	wire v_657;
	wire v_658;
	wire v_659;
	wire v_660;
	wire v_661;
	wire v_662;
	wire v_663;
	wire v_664;
	wire v_665;
	wire v_666;
	wire v_667;
	wire v_668;
	wire v_669;
	wire v_670;
	wire v_671;
	wire v_672;
	wire v_673;
	wire v_674;
	wire v_675;
	wire v_676;
	wire v_677;
	wire v_678;
	wire v_679;
	wire v_680;
	wire v_681;
	wire v_682;
	wire v_683;
	wire v_684;
	wire v_685;
	wire v_686;
	wire v_687;
	wire v_688;
	wire v_689;
	wire v_690;
	wire v_691;
	wire v_692;
	wire v_693;
	wire v_694;
	wire v_695;
	wire v_696;
	wire v_697;
	wire v_698;
	wire v_699;
	wire v_700;
	wire v_701;
	wire v_702;
	wire v_703;
	wire v_704;
	wire v_705;
	wire v_706;
	wire v_707;
	wire v_708;
	wire v_709;
	wire v_710;
	wire v_711;
	wire v_712;
	wire v_713;
	wire v_714;
	wire v_715;
	wire v_716;
	wire v_717;
	wire v_718;
	wire v_719;
	wire v_720;
	wire v_721;
	wire v_722;
	wire v_723;
	wire v_724;
	wire v_725;
	wire v_726;
	wire v_727;
	wire v_728;
	wire v_729;
	wire v_730;
	wire v_731;
	wire v_732;
	wire v_733;
	wire v_734;
	wire v_735;
	wire v_736;
	wire v_737;
	wire v_738;
	wire v_739;
	wire v_740;
	wire v_741;
	wire v_742;
	wire v_743;
	wire v_744;
	wire v_745;
	wire v_746;
	wire v_747;
	wire v_748;
	wire v_749;
	wire v_750;
	wire v_751;
	wire v_752;
	wire v_753;
	wire v_754;
	wire v_755;
	wire v_756;
	wire v_757;
	wire v_758;
	wire v_759;
	wire v_760;
	wire v_761;
	wire v_762;
	wire v_763;
	wire v_764;
	wire v_765;
	wire v_766;
	wire v_767;
	wire v_768;
	wire v_769;
	wire v_770;
	wire v_771;
	wire v_772;
	wire v_773;
	wire v_774;
	wire v_775;
	wire v_776;
	wire v_777;
	wire v_778;
	wire v_779;
	wire v_780;
	wire v_781;
	wire v_782;
	wire v_783;
	wire v_784;
	wire v_785;
	wire v_786;
	wire v_787;
	wire v_788;
	wire v_789;
	wire v_790;
	wire v_791;
	wire v_792;
	wire v_793;
	wire v_794;
	wire v_795;
	wire v_796;
	wire v_797;
	wire v_798;
	wire v_799;
	wire v_800;
	wire v_801;
	wire v_802;
	wire v_803;
	wire v_804;
	wire v_805;
	wire v_806;
	wire v_807;
	wire v_808;
	wire v_809;
	wire v_810;
	wire v_811;
	wire v_812;
	wire v_813;
	wire v_814;
	wire v_815;
	wire v_816;
	wire v_817;
	wire v_818;
	wire v_819;
	wire v_820;
	wire v_821;
	wire v_822;
	wire v_823;
	wire v_824;
	wire v_825;
	wire v_826;
	wire v_827;
	wire v_828;
	wire v_829;
	wire v_830;
	wire v_831;
	wire v_832;
	wire v_833;
	wire v_834;
	wire v_835;
	wire v_836;
	wire v_837;
	wire v_838;
	wire v_839;
	wire v_840;
	wire v_841;
	wire v_842;
	wire v_843;
	wire v_844;
	wire v_845;
	wire v_846;
	wire v_847;
	wire v_848;
	wire v_849;
	wire v_850;
	wire v_851;
	wire v_852;
	wire v_853;
	wire v_854;
	wire v_855;
	wire v_856;
	wire v_857;
	wire v_858;
	wire v_859;
	wire v_860;
	wire v_861;
	wire v_862;
	wire v_863;
	wire v_864;
	wire v_865;
	wire v_866;
	wire v_867;
	wire v_868;
	wire v_869;
	wire v_870;
	wire v_871;
	wire v_872;
	wire v_873;
	wire v_874;
	wire v_875;
	wire v_876;
	wire v_877;
	wire v_878;
	wire v_879;
	wire v_880;
	wire v_881;
	wire v_882;
	wire v_883;
	wire v_884;
	wire v_885;
	wire v_886;
	wire v_887;
	wire v_888;
	wire v_889;
	wire v_890;
	wire v_891;
	wire v_892;
	wire v_893;
	wire v_894;
	wire v_895;
	wire v_896;
	wire v_897;
	wire v_898;
	wire v_899;
	wire v_900;
	wire v_901;
	wire v_902;
	wire v_903;
	wire v_904;
	wire v_905;
	wire v_906;
	wire v_907;
	wire v_908;
	wire v_909;
	wire v_910;
	wire v_911;
	wire v_912;
	wire v_913;
	wire v_914;
	wire v_915;
	wire v_916;
	wire v_917;
	wire v_918;
	wire v_919;
	wire v_920;
	wire v_921;
	wire v_922;
	wire v_923;
	wire v_924;
	wire v_925;
	wire v_926;
	wire v_927;
	wire v_928;
	wire v_929;
	wire v_930;
	wire v_931;
	wire v_932;
	wire v_933;
	wire v_934;
	wire v_935;
	wire v_936;
	wire v_937;
	wire v_938;
	wire v_939;
	wire v_940;
	wire v_941;
	wire v_942;
	wire v_943;
	wire v_944;
	wire v_945;
	wire v_946;
	wire v_947;
	wire v_948;
	wire v_949;
	wire v_950;
	wire v_951;
	wire v_952;
	wire v_953;
	wire v_954;
	wire v_955;
	wire v_956;
	wire v_957;
	wire v_958;
	wire v_959;
	wire v_960;
	wire v_961;
	wire v_962;
	wire v_963;
	wire v_964;
	wire v_965;
	wire v_966;
	wire v_967;
	wire v_968;
	wire v_969;
	wire v_970;
	wire v_971;
	wire v_972;
	wire v_973;
	wire v_974;
	wire v_975;
	wire v_976;
	wire v_977;
	wire v_978;
	wire v_979;
	wire v_980;
	wire v_981;
	wire v_983;
	wire v_984;
	wire v_985;
	wire v_986;
	wire v_987;
	wire v_988;
	wire v_989;
	wire v_990;
	wire v_991;
	wire v_992;
	wire v_993;
	wire v_994;
	wire v_995;
	wire v_996;
	wire v_997;
	wire v_998;
	wire v_999;
	wire v_1000;
	wire v_1001;
	wire v_1002;
	wire v_1003;
	wire v_1004;
	wire v_1005;
	wire v_1006;
	wire v_1007;
	wire v_1008;
	wire v_1009;
	wire v_1010;
	wire v_1011;
	wire v_1012;
	wire v_1013;
	wire v_1014;
	wire v_1015;
	wire v_1016;
	wire v_1017;
	wire v_1018;
	wire v_1019;
	wire v_1020;
	wire v_1021;
	wire v_1022;
	wire v_1023;
	wire v_1024;
	wire v_1025;
	wire v_1026;
	wire v_1027;
	wire v_1028;
	wire v_1029;
	wire v_1030;
	wire v_1031;
	wire v_1032;
	wire v_1033;
	wire v_1034;
	wire v_1035;
	wire v_1036;
	wire v_1037;
	wire v_1038;
	wire v_1039;
	wire v_1040;
	wire v_1041;
	wire v_1042;
	wire v_1043;
	wire v_1044;
	wire v_1045;
	wire v_1046;
	wire v_1047;
	wire v_1048;
	wire v_1049;
	wire v_1050;
	wire v_1051;
	wire v_1052;
	wire v_1053;
	wire v_1054;
	wire v_1055;
	wire v_1056;
	wire v_1057;
	wire v_1058;
	wire v_1059;
	wire v_1060;
	wire v_1061;
	wire v_1062;
	wire v_1063;
	wire v_1064;
	wire v_1065;
	wire v_1066;
	wire v_1067;
	wire v_1068;
	wire v_1069;
	wire v_1070;
	wire v_1071;
	wire v_1072;
	wire v_1073;
	wire v_1074;
	wire v_1075;
	wire v_1076;
	wire v_1077;
	wire v_1078;
	wire v_1079;
	wire v_1080;
	wire v_1081;
	wire v_1082;
	wire v_1083;
	wire v_1084;
	wire v_1085;
	wire v_1086;
	wire v_1087;
	wire v_1088;
	wire v_1089;
	wire v_1090;
	wire v_1091;
	wire v_1092;
	wire v_1093;
	wire v_1094;
	wire v_1095;
	wire v_1096;
	wire v_1097;
	wire v_1098;
	wire v_1099;
	wire v_1100;
	wire v_1101;
	wire v_1102;
	wire v_1103;
	wire v_1104;
	wire v_1105;
	wire v_1106;
	wire v_1107;
	wire v_1108;
	wire v_1109;
	wire v_1110;
	wire v_1111;
	wire v_1112;
	wire v_1113;
	wire v_1114;
	wire v_1115;
	wire v_1116;
	wire v_1117;
	wire v_1118;
	wire v_1119;
	wire v_1120;
	wire v_1121;
	wire v_1122;
	wire v_1123;
	wire v_1124;
	wire v_1125;
	wire v_1126;
	wire v_1127;
	wire v_1128;
	wire v_1129;
	wire v_1130;
	wire v_1131;
	wire v_1132;
	wire v_1133;
	wire v_1134;
	wire v_1135;
	wire v_1136;
	wire v_1137;
	wire v_1138;
	wire v_1139;
	wire v_1140;
	wire v_1141;
	wire v_1142;
	wire v_1143;
	wire v_1144;
	wire v_1145;
	wire v_1146;
	wire v_1147;
	wire v_1148;
	wire v_1149;
	wire v_1150;
	wire v_1151;
	wire v_1152;
	wire v_1153;
	wire v_1154;
	wire v_1155;
	wire v_1156;
	wire v_1157;
	wire v_1158;
	wire v_1159;
	wire v_1160;
	wire v_1161;
	wire v_1162;
	wire v_1163;
	wire v_1164;
	wire v_1165;
	wire v_1166;
	wire v_1167;
	wire v_1168;
	wire v_1169;
	wire v_1170;
	wire v_1171;
	wire v_1172;
	wire v_1173;
	wire v_1174;
	wire v_1175;
	wire v_1176;
	wire v_1177;
	wire v_1178;
	wire v_1179;
	wire v_1180;
	wire v_1181;
	wire v_1182;
	wire v_1183;
	wire v_1184;
	wire v_1185;
	wire v_1186;
	wire v_1187;
	wire v_1188;
	wire v_1189;
	wire v_1190;
	wire v_1191;
	wire v_1192;
	wire v_1193;
	wire v_1194;
	wire v_1195;
	wire v_1196;
	wire v_1197;
	wire v_1198;
	wire v_1199;
	wire v_1200;
	wire v_1201;
	wire v_1202;
	wire v_1203;
	wire v_1204;
	wire v_1205;
	wire v_1206;
	wire v_1207;
	wire v_1208;
	wire v_1209;
	wire v_1210;
	wire v_1211;
	wire v_1212;
	wire v_1213;
	wire v_1214;
	wire v_1215;
	wire v_1216;
	wire v_1217;
	wire v_1218;
	wire v_1219;
	wire v_1220;
	wire v_1221;
	wire v_1222;
	wire v_1223;
	wire v_1224;
	wire v_1225;
	wire v_1226;
	wire v_1227;
	wire v_1228;
	wire v_1229;
	wire v_1230;
	wire v_1231;
	wire v_1232;
	wire v_1233;
	wire v_1234;
	wire v_1235;
	wire v_1236;
	wire v_1237;
	wire v_1238;
	wire v_1239;
	wire v_1240;
	wire v_1241;
	wire v_1242;
	wire v_1243;
	wire v_1244;
	wire v_1245;
	wire v_1246;
	wire v_1247;
	wire v_1248;
	wire v_1249;
	wire v_1250;
	wire v_1251;
	wire v_1252;
	wire v_1253;
	wire v_1254;
	wire v_1255;
	wire v_1256;
	wire v_1257;
	wire v_1258;
	wire v_1259;
	wire v_1260;
	wire v_1261;
	wire v_1262;
	wire v_1263;
	wire v_1264;
	wire v_1265;
	wire v_1266;
	wire v_1267;
	wire v_1268;
	wire v_1269;
	wire v_1270;
	wire v_1271;
	wire v_1272;
	wire v_1273;
	wire v_1274;
	wire v_1275;
	wire v_1276;
	wire v_1277;
	wire v_1278;
	wire v_1279;
	wire v_1280;
	wire v_1281;
	wire v_1282;
	wire v_1283;
	wire v_1284;
	wire v_1285;
	wire v_1286;
	wire v_1287;
	wire v_1288;
	wire v_1289;
	wire v_1290;
	wire v_1291;
	wire v_1292;
	wire v_1293;
	wire v_1294;
	wire v_1295;
	wire v_1296;
	wire v_1297;
	wire v_1298;
	wire v_1299;
	wire v_1300;
	wire v_1301;
	wire v_1302;
	wire v_1303;
	wire v_1304;
	wire v_1305;
	wire v_1306;
	wire v_1307;
	wire v_1308;
	wire v_1309;
	wire v_1310;
	wire v_1311;
	wire v_1312;
	wire v_1313;
	wire v_1314;
	wire v_1315;
	wire v_1316;
	wire v_1317;
	wire v_1318;
	wire v_1319;
	wire v_1320;
	wire v_1321;
	wire v_1322;
	wire v_1323;
	wire v_1324;
	wire v_1325;
	wire v_1326;
	wire v_1327;
	wire v_1328;
	wire v_1329;
	wire v_1330;
	wire v_1331;
	wire v_1332;
	wire v_1333;
	wire v_1334;
	wire v_1335;
	wire v_1336;
	wire v_1337;
	wire v_1338;
	wire v_1339;
	wire v_1340;
	wire v_1341;
	wire v_1342;
	wire v_1343;
	wire v_1344;
	wire v_1345;
	wire v_1346;
	wire v_1347;
	wire v_1348;
	wire v_1349;
	wire v_1350;
	wire v_1351;
	wire v_1352;
	wire v_1353;
	wire v_1354;
	wire v_1355;
	wire v_1356;
	wire v_1357;
	wire v_1358;
	wire v_1359;
	wire v_1360;
	wire v_1361;
	wire v_1362;
	wire v_1363;
	wire v_1364;
	wire v_1365;
	wire v_1366;
	wire v_1367;
	wire v_1368;
	wire v_1369;
	wire v_1370;
	wire v_1371;
	wire v_1372;
	wire v_1373;
	wire v_1374;
	wire v_1375;
	wire v_1376;
	wire v_1377;
	wire v_1378;
	wire v_1379;
	wire v_1380;
	wire v_1381;
	wire v_1382;
	wire v_1383;
	wire v_1384;
	wire v_1385;
	wire v_1386;
	wire v_1387;
	wire v_1388;
	wire v_1389;
	wire v_1390;
	wire v_1391;
	wire v_1392;
	wire v_1393;
	wire v_1394;
	wire v_1395;
	wire v_1396;
	wire v_1397;
	wire v_1398;
	wire v_1399;
	wire v_1400;
	wire v_1401;
	wire v_1402;
	wire v_1403;
	wire v_1404;
	wire v_1405;
	wire v_1406;
	wire v_1407;
	wire v_1408;
	wire v_1409;
	wire v_1410;
	wire v_1411;
	wire v_1412;
	wire v_1413;
	wire v_1414;
	wire v_1415;
	wire v_1416;
	wire v_1417;
	wire v_1418;
	wire v_1419;
	wire v_1420;
	wire v_1421;
	wire v_1422;
	wire v_1423;
	wire v_1424;
	wire v_1425;
	wire v_1426;
	wire v_1427;
	wire v_1428;
	wire v_1429;
	wire v_1430;
	wire v_1431;
	wire v_1432;
	wire v_1433;
	wire v_1434;
	wire v_1435;
	wire v_1436;
	wire v_1437;
	wire v_1438;
	wire v_1439;
	wire v_1440;
	wire v_1441;
	wire v_1442;
	wire v_1443;
	wire v_1444;
	wire v_1445;
	wire v_1446;
	wire v_1447;
	wire v_1448;
	wire v_1449;
	wire v_1450;
	wire v_1451;
	wire v_1452;
	wire v_1453;
	wire v_1454;
	wire v_1455;
	wire v_1456;
	wire v_1457;
	wire v_1458;
	wire v_1459;
	wire v_1460;
	wire v_1461;
	wire v_1462;
	wire v_1463;
	wire v_1464;
	wire v_1465;
	wire v_1466;
	wire v_1467;
	wire v_1468;
	wire v_1469;
	wire v_1470;
	wire v_1471;
	wire v_1472;
	wire v_1473;
	wire v_1474;
	wire v_1475;
	wire v_1476;
	wire v_1477;
	wire v_1478;
	wire v_1479;
	wire v_1480;
	wire v_1481;
	wire v_1482;
	wire v_1483;
	wire v_1484;
	wire v_1485;
	wire v_1486;
	wire v_1487;
	wire v_1488;
	wire v_1489;
	wire v_1490;
	wire v_1491;
	wire v_1492;
	wire v_1493;
	wire v_1494;
	wire v_1495;
	wire v_1496;
	wire v_1497;
	wire v_1498;
	wire v_1499;
	wire v_1500;
	wire v_1501;
	wire v_1502;
	wire v_1503;
	wire v_1504;
	wire v_1505;
	wire v_1506;
	wire v_1507;
	wire v_1508;
	wire v_1509;
	wire v_1510;
	wire v_1511;
	wire v_1512;
	wire v_1513;
	wire v_1514;
	wire v_1515;
	wire v_1516;
	wire v_1517;
	wire v_1518;
	wire v_1519;
	wire v_1520;
	wire v_1521;
	wire v_1522;
	wire v_1523;
	wire v_1524;
	wire v_1525;
	wire v_1526;
	wire v_1527;
	wire v_1528;
	wire v_1529;
	wire v_1530;
	wire v_1531;
	wire v_1532;
	wire v_1533;
	wire v_1534;
	wire v_1535;
	wire v_1536;
	wire v_1537;
	wire v_1538;
	wire v_1539;
	wire v_1540;
	wire v_1541;
	wire v_1542;
	wire v_1543;
	wire v_1544;
	wire v_1545;
	wire v_1546;
	wire v_1547;
	wire v_1548;
	wire v_1549;
	wire v_1550;
	wire v_1551;
	wire v_1552;
	wire v_1553;
	wire v_1554;
	wire v_1555;
	wire v_1556;
	wire v_1557;
	wire v_1558;
	wire v_1559;
	wire v_1560;
	wire v_1561;
	wire v_1562;
	wire v_1563;
	wire v_1564;
	wire v_1565;
	wire v_1566;
	wire v_1567;
	wire v_1568;
	wire v_1569;
	wire v_1570;
	wire v_1571;
	wire v_1572;
	wire v_1573;
	wire v_1574;
	wire v_1575;
	wire v_1576;
	wire v_1577;
	wire v_1578;
	wire v_1579;
	wire v_1580;
	wire v_1581;
	wire v_1583;
	wire v_1584;
	wire v_1585;
	wire v_1586;
	wire v_1587;
	wire v_1588;
	wire v_1589;
	wire v_1590;
	wire v_1591;
	wire v_1592;
	wire v_1593;
	wire v_1594;
	wire v_1595;
	wire v_1596;
	wire v_1597;
	wire v_1598;
	wire v_1599;
	wire v_1600;
	wire v_1601;
	wire v_1602;
	wire v_1603;
	wire v_1604;
	wire v_1605;
	wire v_1606;
	wire v_1607;
	wire v_1608;
	wire v_1609;
	wire v_1610;
	wire v_1611;
	wire v_1612;
	wire v_1613;
	wire v_1614;
	wire v_1615;
	wire v_1616;
	wire v_1617;
	wire v_1618;
	wire v_1619;
	wire v_1620;
	wire v_1621;
	wire v_1622;
	wire v_1623;
	wire v_1624;
	wire v_1625;
	wire v_1626;
	wire v_1627;
	wire v_1628;
	wire v_1629;
	wire v_1630;
	wire v_1631;
	wire v_1632;
	wire v_1633;
	wire v_1634;
	wire v_1635;
	wire v_1636;
	wire v_1637;
	wire v_1638;
	wire v_1639;
	wire v_1640;
	wire v_1641;
	wire v_1642;
	wire v_1643;
	wire v_1644;
	wire v_1645;
	wire v_1646;
	wire v_1647;
	wire v_1648;
	wire v_1649;
	wire v_1650;
	wire v_1651;
	wire v_1652;
	wire v_1653;
	wire v_1654;
	wire v_1655;
	wire v_1656;
	wire v_1657;
	wire v_1658;
	wire v_1659;
	wire v_1660;
	wire v_1661;
	wire v_1662;
	wire v_1663;
	wire v_1664;
	wire v_1665;
	wire v_1666;
	wire v_1667;
	wire v_1668;
	wire v_1669;
	wire v_1670;
	wire v_1671;
	wire v_1672;
	wire v_1673;
	wire v_1674;
	wire v_1675;
	wire v_1676;
	wire v_1677;
	wire v_1678;
	wire v_1679;
	wire v_1680;
	wire v_1681;
	wire v_1682;
	wire v_1683;
	wire v_1684;
	wire v_1685;
	wire v_1686;
	wire v_1687;
	wire v_1688;
	wire v_1689;
	wire v_1690;
	wire v_1691;
	wire v_1692;
	wire v_1693;
	wire v_1694;
	wire v_1695;
	wire v_1696;
	wire v_1697;
	wire v_1698;
	wire v_1699;
	wire v_1700;
	wire v_1701;
	wire v_1702;
	wire v_1703;
	wire v_1704;
	wire v_1705;
	wire v_1706;
	wire v_1707;
	wire v_1708;
	wire v_1709;
	wire v_1710;
	wire v_1711;
	wire v_1712;
	wire v_1713;
	wire v_1714;
	wire v_1715;
	wire v_1716;
	wire v_1717;
	wire v_1718;
	wire v_1719;
	wire v_1720;
	wire v_1721;
	wire v_1722;
	wire v_1723;
	wire v_1724;
	wire v_1725;
	wire v_1726;
	wire v_1727;
	wire v_1728;
	wire v_1729;
	wire v_1730;
	wire v_1731;
	wire v_1732;
	wire v_1733;
	wire v_1734;
	wire v_1735;
	wire v_1736;
	wire v_1737;
	wire v_1738;
	wire v_1739;
	wire v_1740;
	wire v_1741;
	wire v_1742;
	wire v_1743;
	wire v_1744;
	wire v_1745;
	wire v_1746;
	wire v_1747;
	wire v_1748;
	wire v_1749;
	wire v_1750;
	wire v_1751;
	wire v_1752;
	wire v_1753;
	wire v_1754;
	wire v_1755;
	wire v_1756;
	wire v_1757;
	wire v_1758;
	wire v_1759;
	wire v_1760;
	wire v_1761;
	wire v_1762;
	wire v_1763;
	wire v_1764;
	wire v_1765;
	wire v_1766;
	wire v_1767;
	wire v_1768;
	wire v_1769;
	wire v_1770;
	wire v_1771;
	wire v_1772;
	wire v_1773;
	wire v_1774;
	wire v_1775;
	wire v_1776;
	wire v_1777;
	wire v_1778;
	wire v_1779;
	wire v_1780;
	wire v_1781;
	wire v_1782;
	wire v_1783;
	wire v_1784;
	wire v_1785;
	wire v_1786;
	wire v_1787;
	wire v_1788;
	wire v_1789;
	wire v_1790;
	wire v_1791;
	wire v_1792;
	wire v_1793;
	wire v_1794;
	wire v_1795;
	wire v_1796;
	wire v_1797;
	wire v_1798;
	wire v_1799;
	wire v_1800;
	wire v_1801;
	wire v_1802;
	wire v_1803;
	wire v_1804;
	wire v_1805;
	wire v_1806;
	wire v_1807;
	wire v_1808;
	wire v_1809;
	wire v_1810;
	wire v_1811;
	wire v_1812;
	wire v_1813;
	wire v_1814;
	wire v_1815;
	wire v_1816;
	wire v_1817;
	wire v_1818;
	wire v_1819;
	wire v_1820;
	wire v_1821;
	wire v_1822;
	wire v_1823;
	wire v_1824;
	wire v_1825;
	wire v_1826;
	wire v_1827;
	wire v_1828;
	wire v_1829;
	wire v_1830;
	wire v_1831;
	wire v_1832;
	wire v_1833;
	wire v_1834;
	wire v_1835;
	wire v_1836;
	wire v_1837;
	wire v_1838;
	wire v_1839;
	wire v_1840;
	wire v_1841;
	wire v_1842;
	wire v_1843;
	wire v_1844;
	wire v_1845;
	wire v_1846;
	wire v_1847;
	wire v_1848;
	wire v_1849;
	wire v_1850;
	wire v_1851;
	wire v_1852;
	wire v_1853;
	wire v_1854;
	wire v_1855;
	wire v_1856;
	wire v_1857;
	wire v_1858;
	wire v_1859;
	wire v_1860;
	wire v_1861;
	wire v_1862;
	wire v_1863;
	wire v_1864;
	wire v_1865;
	wire v_1866;
	wire v_1867;
	wire v_1868;
	wire v_1869;
	wire v_1870;
	wire v_1871;
	wire v_1872;
	wire v_1873;
	wire v_1874;
	wire v_1875;
	wire v_1876;
	wire v_1877;
	wire v_1878;
	wire v_1879;
	wire v_1880;
	wire v_1881;
	wire v_1882;
	wire v_1883;
	wire v_1884;
	wire v_1885;
	wire v_1886;
	wire v_1887;
	wire v_1888;
	wire v_1889;
	wire v_1890;
	wire v_1891;
	wire v_1892;
	wire v_1893;
	wire v_1894;
	wire v_1895;
	wire v_1896;
	wire v_1897;
	wire v_1898;
	wire v_1899;
	wire v_1900;
	wire v_1901;
	wire v_1902;
	wire v_1903;
	wire v_1904;
	wire v_1905;
	wire v_1906;
	wire v_1907;
	wire v_1908;
	wire v_1909;
	wire v_1910;
	wire v_1911;
	wire v_1912;
	wire v_1913;
	wire v_1914;
	wire v_1915;
	wire v_1916;
	wire v_1917;
	wire v_1918;
	wire v_1919;
	wire v_1920;
	wire v_1921;
	wire v_1922;
	wire v_1923;
	wire v_1924;
	wire v_1925;
	wire v_1926;
	wire v_1927;
	wire v_1928;
	wire v_1929;
	wire v_1930;
	wire v_1931;
	wire v_1932;
	wire v_1933;
	wire v_1934;
	wire v_1935;
	wire v_1936;
	wire v_1937;
	wire v_1938;
	wire v_1939;
	wire v_1940;
	wire v_1941;
	wire v_1942;
	wire v_1943;
	wire v_1944;
	wire v_1945;
	wire v_1946;
	wire v_1947;
	wire v_1948;
	wire v_1949;
	wire v_1950;
	wire v_1951;
	wire v_1952;
	wire v_1953;
	wire v_1954;
	wire v_1955;
	wire v_1956;
	wire v_1957;
	wire v_1958;
	wire v_1959;
	wire v_1960;
	wire v_1961;
	wire v_1962;
	wire v_1963;
	wire v_1964;
	wire v_1965;
	wire v_1966;
	wire v_1967;
	wire v_1968;
	wire v_1969;
	wire v_1970;
	wire v_1971;
	wire v_1972;
	wire v_1973;
	wire v_1974;
	wire v_1975;
	wire v_1976;
	wire v_1977;
	wire v_1978;
	wire v_1979;
	wire v_1980;
	wire v_1981;
	wire v_1982;
	wire v_1983;
	wire v_1984;
	wire v_1985;
	wire v_1986;
	wire v_1987;
	wire v_1988;
	wire v_1989;
	wire v_1990;
	wire v_1991;
	wire v_1992;
	wire v_1993;
	wire v_1994;
	wire v_1995;
	wire v_1996;
	wire v_1997;
	wire v_1998;
	wire v_1999;
	wire v_2000;
	wire v_2001;
	wire v_2002;
	wire v_2003;
	wire v_2004;
	wire v_2005;
	wire v_2006;
	wire v_2007;
	wire v_2008;
	wire v_2009;
	wire v_2010;
	wire v_2011;
	wire v_2012;
	wire v_2013;
	wire v_2014;
	wire v_2015;
	wire v_2016;
	wire v_2017;
	wire v_2018;
	wire v_2019;
	wire v_2020;
	wire v_2021;
	wire v_2022;
	wire v_2023;
	wire v_2024;
	wire v_2025;
	wire v_2026;
	wire v_2027;
	wire v_2028;
	wire v_2029;
	wire v_2030;
	wire v_2031;
	wire v_2032;
	wire v_2033;
	wire v_2034;
	wire v_2035;
	wire v_2036;
	wire v_2037;
	wire v_2038;
	wire v_2039;
	wire v_2040;
	wire v_2041;
	wire v_2042;
	wire v_2043;
	wire v_2044;
	wire v_2045;
	wire v_2046;
	wire v_2047;
	wire v_2048;
	wire v_2049;
	wire v_2050;
	wire v_2051;
	wire v_2052;
	wire v_2053;
	wire v_2054;
	wire v_2055;
	wire v_2056;
	wire v_2057;
	wire v_2058;
	wire v_2059;
	wire v_2060;
	wire v_2061;
	wire v_2062;
	wire v_2063;
	wire v_2064;
	wire v_2065;
	wire v_2066;
	wire v_2067;
	wire v_2068;
	wire v_2069;
	wire v_2070;
	wire v_2071;
	wire v_2072;
	wire v_2073;
	wire v_2074;
	wire v_2075;
	wire v_2076;
	wire v_2077;
	wire v_2078;
	wire v_2079;
	wire v_2080;
	wire v_2081;
	wire v_2082;
	wire v_2083;
	wire v_2084;
	wire v_2085;
	wire v_2086;
	wire v_2087;
	wire v_2088;
	wire v_2089;
	wire v_2090;
	wire v_2091;
	wire v_2092;
	wire v_2093;
	wire v_2094;
	wire v_2095;
	wire v_2096;
	wire v_2097;
	wire v_2098;
	wire v_2099;
	wire v_2100;
	wire v_2101;
	wire v_2102;
	wire v_2103;
	wire v_2104;
	wire v_2105;
	wire v_2106;
	wire v_2107;
	wire v_2108;
	wire v_2109;
	wire v_2110;
	wire v_2111;
	wire v_2112;
	wire v_2113;
	wire v_2114;
	wire v_2115;
	wire v_2116;
	wire v_2117;
	wire v_2118;
	wire v_2119;
	wire v_2120;
	wire v_2121;
	wire v_2122;
	wire v_2123;
	wire v_2124;
	wire v_2125;
	wire v_2126;
	wire v_2127;
	wire v_2128;
	wire v_2129;
	wire v_2130;
	wire v_2131;
	wire v_2132;
	wire v_2133;
	wire v_2134;
	wire v_2135;
	wire v_2136;
	wire v_2137;
	wire v_2138;
	wire v_2139;
	wire v_2140;
	wire v_2141;
	wire v_2142;
	wire v_2143;
	wire v_2144;
	wire v_2145;
	wire v_2146;
	wire v_2147;
	wire v_2148;
	wire v_2149;
	wire v_2150;
	wire v_2151;
	wire v_2152;
	wire v_2153;
	wire v_2154;
	wire v_2155;
	wire v_2156;
	wire v_2157;
	wire v_2158;
	wire v_2159;
	wire v_2160;
	wire v_2161;
	wire v_2162;
	wire v_2163;
	wire v_2164;
	wire v_2165;
	wire v_2166;
	wire v_2167;
	wire v_2168;
	wire v_2169;
	wire v_2170;
	wire v_2171;
	wire v_2172;
	wire v_2173;
	wire v_2174;
	wire v_2175;
	wire v_2176;
	wire v_2177;
	wire v_2178;
	wire v_2179;
	wire v_2180;
	wire v_2181;
	wire v_2182;
	wire v_2183;
	wire v_2184;
	wire v_2185;
	wire v_2186;
	wire v_2187;
	wire v_2188;
	wire v_2189;
	wire v_2190;
	wire v_2191;
	wire v_2192;
	wire v_2193;
	wire v_2194;
	wire v_2195;
	wire v_2196;
	wire v_2197;
	wire v_2198;
	wire v_2199;
	wire v_2200;
	wire v_2201;
	wire v_2202;
	wire v_2203;
	wire v_2204;
	wire v_2205;
	wire v_2206;
	wire v_2207;
	wire v_2208;
	wire v_2209;
	wire v_2210;
	wire v_2211;
	wire v_2212;
	wire v_2213;
	wire v_2214;
	wire v_2215;
	wire v_2216;
	wire v_2217;
	wire v_2218;
	wire v_2219;
	wire v_2220;
	wire v_2221;
	wire x_1;
	wire x_2;
	wire x_3;
	wire x_4;
	wire x_5;
	wire x_6;
	wire x_7;
	output o_1;
	assign v_2159 = (((((((~v_3 & ~v_4)) & ~v_5)) & ~v_6)) & ~v_7);
	assign v_2160 = (((~v_8 & ~v_9)) & ~v_10);
	assign v_267 = (~v_11 & v_2);
	assign v_266 = (~v_11 & v_1);
	assign v_270 = v_1);
	assign v_327 = (~v_13 & v_10);
	assign v_324 = (~v_13 & v_9);
	assign v_321 = (~v_13 & v_8);
	assign v_318 = (~v_13 & v_7);
	assign v_315 = (~v_13 & v_6);
	assign v_312 = (~v_13 & v_5);
	assign v_309 = (~v_13 & v_4);
	assign v_306 = (~v_13 & v_3);
	assign v_2163 = (((((((~v_1 & ~v_2)) & ~v_11)) & ~v_12)) & ~v_13);
	assign v_347 = ~v_1);
	assign v_407 = v_1);
	assign v_446 = (~v_1 & v_14);
	assign v_449 = (~v_1 & v_15);
	assign v_452 = (~v_1 & v_16);
	assign v_455 = (~v_1 & v_17);
	assign v_458 = (~v_1 & v_18);
	assign v_2161 = (((((((~v_14 & ~v_15)) & ~v_16)) & ~v_17)) & ~v_18);
	assign v_461 = (~v_1 & v_19);
	assign v_464 = (~v_1 & v_20);
	assign v_467 = (~v_1 & v_21);
	assign v_470 = (~v_1 & v_22);
	assign v_473 = (~v_1 & v_23);
	assign v_2162 = (((((((~v_19 & ~v_20)) & ~v_21)) & ~v_22)) & ~v_23);
	assign v_486 = v_2);
	assign v_263 = (((((~v_24 & ~v_25)) & ~v_26)) & ~v_27);
	assign v_264 = (((((~v_31 & ~v_32)) & ~v_33)) & ~v_34);
	assign v_689 = (~v_13 & v_36);
	assign v_2164 = (((((((~v_28 & ~v_29)) & ~v_30)) & ~v_35)) & ~v_36);
	assign v_620 = (v_38 & v_34);
	assign v_617 = (v_38 & v_33);
	assign v_614 = (v_38 & v_32);
	assign v_611 = (v_38 & v_31);
	assign v_511 = (v_38 & v_27);
	assign v_508 = (v_38 & v_26);
	assign v_505 = (v_38 & v_25);
	assign v_502 = (v_38 & v_24);
	assign v_631 = (v_38 & v_34);
	assign v_628 = (v_38 & v_33);
	assign v_625 = (v_38 & v_32);
	assign v_622 = (v_38 & v_31);
	assign v_522 = (v_38 & v_27);
	assign v_519 = (v_38 & v_26);
	assign v_516 = (v_38 & v_25);
	assign v_513 = (v_38 & v_24);
	assign v_579 = (v_38 & v_29);
	assign v_566 = (v_38 & v_28);
	assign v_677 = (~v_38 & v_35);
	assign v_567 = (v_38 & v_28);
	assign v_643 = (~v_38 & v_34);
	assign v_640 = (~v_38 & v_33);
	assign v_637 = (~v_38 & v_32);
	assign v_634 = (~v_38 & v_31);
	assign v_534 = (~v_38 & v_27);
	assign v_531 = (~v_38 & v_26);
	assign v_528 = (~v_38 & v_25);
	assign v_525 = (~v_38 & v_24);
	assign v_679 = (~v_38 & v_35);
	assign v_585 = (~v_38 & v_29);
	assign v_655 = (v_38 & v_34);
	assign v_652 = (v_38 & v_33);
	assign v_649 = (v_38 & v_32);
	assign v_646 = (v_38 & v_31);
	assign v_546 = (v_38 & v_27);
	assign v_543 = (v_38 & v_26);
	assign v_540 = (v_38 & v_25);
	assign v_537 = (v_38 & v_24);
	assign v_682 = (v_38 & v_35);
	assign v_588 = (v_38 & v_29);
	assign v_572 = (v_38 & v_28);
	assign v_667 = (~v_38 & v_34);
	assign v_664 = (~v_38 & v_33);
	assign v_661 = (~v_38 & v_32);
	assign v_658 = (~v_38 & v_31);
	assign v_558 = (~v_38 & v_27);
	assign v_555 = (~v_38 & v_26);
	assign v_552 = (~v_38 & v_25);
	assign v_549 = (~v_38 & v_24);
	assign v_591 = (~v_38 & v_29);
	assign v_575 = (~v_38 & v_28);
	assign v_601 = (v_39 & v_30);
	assign v_603 = (v_39 & v_30);
	assign v_606 = (~v_39 & v_30);
	assign v_750 = (~v_11 & v_40);
	assign v_393 = (v_40 & v_12);
	assign v_400 = (~v_40 & v_13);
	assign v_396 = (~v_40 & v_12);
	assign v_695 = (~v_41 & v_3);
	assign v_697 = (v_41 & v_4);
	assign v_762 = v_4);
	assign v_700 = (~v_41 & v_5);
	assign v_703 = (v_41 & v_6);
	assign v_706 = (~v_41 & v_7);
	assign v_709 = (v_41 & v_8);
	assign v_712 = (~v_41 & v_9);
	assign v_715 = (v_41 & v_10);
	assign v_779 = (~v_1 & v_41);
	assign v_595 = (v_42 & v_30);
	assign v_786 = (v_39 & v_42);
	assign v_788 = (v_39 & v_42);
	assign v_791 = (~v_39 & v_42);
	assign v_2165 = (((((((~v_37 & ~v_38)) & ~v_39)) & ~v_40)) & ~v_42);
	assign v_724 = (~v_43 & v_38);
	assign v_795 = (~v_42 & v_43);
	assign v_800 = (v_39 & v_43);
	assign v_802 = (v_39 & v_43);
	assign v_811 = (~v_43 & v_44);
	assign v_813 = (~v_38 & v_44);
	assign v_815 = (~v_38 & v_44);
	assign v_820 = (~v_38 & v_44);
	assign v_823 = (v_38 & v_44);
	assign v_826 = (~v_38 & v_44);
	assign v_829 = (v_38 & v_44);
	assign v_805 = (~v_44 & v_43);
	assign v_832 = (~v_38 & v_44);
	assign v_746 = (~v_39 & v_44);
	assign v_836 = (~v_11 & v_45);
	assign v_796 = (~v_45 & v_43);
	assign v_783 = (~v_42 & v_45);
	assign v_782 = (~v_45 & v_42);
	assign v_597 = (~v_45 & v_30);
	assign v_839 = (~v_40 & v_45);
	assign v_841 = (~v_40 & v_45);
	assign v_742 = (~v_39 & v_45);
	assign v_844 = (v_40 & v_45);
	assign v_849 = (v_45 & v_46);
	assign v_851 = (v_39 & v_46);
	assign v_401 = (~v_46 & v_13);
	assign v_855 = (~v_39 & v_46);
	assign v_757 = (~v_40 & v_46);
	assign v_861 = (~v_66 & v_49);
	assign v_860 = (~v_66 & v_47);
	assign v_392 = v_6);
	assign v_864 = v_6);
	assign v_921 = (~v_68 & v_57);
	assign v_918 = (~v_68 & v_56);
	assign v_915 = (~v_68 & v_55);
	assign v_912 = (~v_68 & v_54);
	assign v_909 = (~v_68 & v_53);
	assign v_906 = (~v_68 & v_52);
	assign v_903 = (~v_68 & v_51);
	assign v_900 = (~v_68 & v_50);
	assign v_941 = ~v_6);
	assign v_1001 = v_6);
	assign v_1040 = (~v_47 & v_69);
	assign v_1043 = (~v_47 & v_70);
	assign v_1046 = (~v_47 & v_71);
	assign v_1049 = (~v_47 & v_72);
	assign v_1052 = (~v_47 & v_73);
	assign v_1055 = (~v_47 & v_74);
	assign v_1058 = (~v_47 & v_75);
	assign v_1061 = (~v_47 & v_76);
	assign v_1064 = (~v_47 & v_77);
	assign v_1067 = (~v_47 & v_78);
	assign v_1080 = v_7);
	assign v_580 = (v_85 & v_29);
	assign v_675 = (v_85 & v_35);
	assign v_732 = (v_38 & v_85);
	assign v_1283 = (~v_68 & v_92);
	assign v_1214 = (v_94 & v_90);
	assign v_1211 = (v_94 & v_89);
	assign v_1208 = (v_94 & v_88);
	assign v_1205 = (v_94 & v_87);
	assign v_1105 = (v_94 & v_82);
	assign v_1102 = (v_94 & v_81);
	assign v_1099 = (v_94 & v_80);
	assign v_1096 = (v_94 & v_79);
	assign v_1225 = (v_94 & v_90);
	assign v_1222 = (v_94 & v_89);
	assign v_1219 = (v_94 & v_88);
	assign v_1216 = (v_94 & v_87);
	assign v_1116 = (v_94 & v_82);
	assign v_1113 = (v_94 & v_81);
	assign v_1110 = (v_94 & v_80);
	assign v_1107 = (v_94 & v_79);
	assign v_1173 = (v_94 & v_84);
	assign v_1160 = (v_94 & v_83);
	assign v_1271 = (~v_94 & v_91);
	assign v_1161 = (v_94 & v_83);
	assign v_1237 = (~v_94 & v_90);
	assign v_1234 = (~v_94 & v_89);
	assign v_1231 = (~v_94 & v_88);
	assign v_1228 = (~v_94 & v_87);
	assign v_1128 = (~v_94 & v_82);
	assign v_1125 = (~v_94 & v_81);
	assign v_1122 = (~v_94 & v_80);
	assign v_1119 = (~v_94 & v_79);
	assign v_1273 = (~v_94 & v_91);
	assign v_1179 = (~v_94 & v_84);
	assign v_1249 = (v_94 & v_90);
	assign v_1246 = (v_94 & v_89);
	assign v_1243 = (v_94 & v_88);
	assign v_1240 = (v_94 & v_87);
	assign v_1140 = (v_94 & v_82);
	assign v_1137 = (v_94 & v_81);
	assign v_1134 = (v_94 & v_80);
	assign v_1131 = (v_94 & v_79);
	assign v_1276 = (v_94 & v_91);
	assign v_1182 = (v_94 & v_84);
	assign v_1166 = (v_94 & v_83);
	assign v_1261 = (~v_94 & v_90);
	assign v_1258 = (~v_94 & v_89);
	assign v_1255 = (~v_94 & v_88);
	assign v_1252 = (~v_94 & v_87);
	assign v_1152 = (~v_94 & v_82);
	assign v_1149 = (~v_94 & v_81);
	assign v_1146 = (~v_94 & v_80);
	assign v_1143 = (~v_94 & v_79);
	assign v_1185 = (~v_94 & v_84);
	assign v_1169 = (~v_94 & v_83);
	assign v_1195 = (v_95 & v_86);
	assign v_1197 = (v_95 & v_86);
	assign v_1200 = (~v_95 & v_86);
	assign v_1344 = (~v_66 & v_96);
	assign v_987 = (v_96 & v_67);
	assign v_994 = (~v_96 & v_68);
	assign v_990 = (~v_96 & v_67);
	assign v_1289 = (~v_97 & v_50);
	assign v_1291 = (v_97 & v_51);
	assign v_1356 = v_9);
	assign v_1294 = (~v_97 & v_52);
	assign v_1297 = (v_97 & v_53);
	assign v_1300 = (~v_97 & v_54);
	assign v_1303 = (v_97 & v_55);
	assign v_1306 = (~v_97 & v_56);
	assign v_1309 = (v_97 & v_57);
	assign v_1373 = (~v_47 & v_97);
	assign v_1189 = (v_98 & v_86);
	assign v_1380 = (v_95 & v_98);
	assign v_1382 = (v_95 & v_98);
	assign v_1385 = (~v_95 & v_98);
	assign v_1318 = (~v_99 & v_94);
	assign v_1389 = (~v_98 & v_99);
	assign v_1394 = (v_95 & v_99);
	assign v_1396 = (v_95 & v_99);
	assign v_1405 = (~v_99 & v_100);
	assign v_1407 = (~v_94 & v_100);
	assign v_1409 = (~v_94 & v_100);
	assign v_1414 = (~v_94 & v_100);
	assign v_1417 = (v_94 & v_100);
	assign v_1420 = (~v_94 & v_100);
	assign v_1423 = (v_94 & v_100);
	assign v_1399 = (~v_100 & v_99);
	assign v_1426 = (~v_94 & v_100);
	assign v_1340 = (~v_95 & v_100);
	assign v_1430 = (~v_66 & v_101);
	assign v_1390 = (~v_101 & v_99);
	assign v_1377 = (~v_98 & v_101);
	assign v_1376 = (~v_101 & v_98);
	assign v_1191 = (~v_101 & v_86);
	assign v_1433 = (~v_96 & v_101);
	assign v_1435 = (~v_96 & v_101);
	assign v_1336 = (~v_95 & v_101);
	assign v_1438 = (v_96 & v_101);
	assign v_1443 = (v_101 & v_102);
	assign v_1445 = (v_95 & v_102);
	assign v_995 = (~v_102 & v_68);
	assign v_1449 = (~v_95 & v_102);
	assign v_1351 = (~v_96 & v_102);
	assign v_986 = v_12);
	assign v_1174 = (v_141 & v_84);
	assign v_1269 = (v_141 & v_91);
	assign v_1326 = (v_94 & v_141);
	assign v_2055 = (v_159 ^ v_103);
	assign v_2056 = (v_160 ^ v_105);
	assign v_2057 = (v_161 ^ v_106);
	assign v_2058 = (v_162 ^ v_107);
	assign v_2059 = (v_163 ^ v_108);
	assign v_2060 = (v_164 ^ v_109);
	assign v_2061 = (v_165 ^ v_110);
	assign v_2186 = (((((((~v_161 & ~v_162)) & ~v_163)) & ~v_164)) & ~v_165);
	assign v_2062 = (v_166 ^ v_111);
	assign v_2063 = (v_167 ^ v_112);
	assign v_2064 = (v_168 ^ v_113);
	assign v_2187 = (((~v_166 & ~v_167)) & ~v_168);
	assign v_1461 = (~v_169 & v_160);
	assign v_1460 = (~v_169 & v_159);
	assign v_2066 = (v_169 ^ v_122);
	assign v_2067 = (v_170 ^ v_123);
	assign v_1464 = v_17);
	assign v_1521 = (~v_171 & v_168);
	assign v_1518 = (~v_171 & v_167);
	assign v_1515 = (~v_171 & v_166);
	assign v_1512 = (~v_171 & v_165);
	assign v_1509 = (~v_171 & v_164);
	assign v_1506 = (~v_171 & v_163);
	assign v_1503 = (~v_171 & v_162);
	assign v_1500 = (~v_171 & v_161);
	assign v_2068 = (v_171 ^ v_124);
	assign v_2190 = (((((((~v_159 & ~v_160)) & ~v_169)) & ~v_170)) & ~v_171);
	assign v_1541 = ~v_17);
	assign v_1601 = v_17);
	assign v_1640 = (~v_159 & v_172);
	assign v_2069 = (v_172 ^ v_125);
	assign v_1643 = (~v_159 & v_173);
	assign v_2070 = (v_173 ^ v_126);
	assign v_1646 = (~v_159 & v_174);
	assign v_2071 = (v_174 ^ v_127);
	assign v_1649 = (~v_159 & v_175);
	assign v_2072 = (v_175 ^ v_128);
	assign v_1652 = (~v_159 & v_176);
	assign v_2073 = (v_176 ^ v_129);
	assign v_2188 = (((((((~v_172 & ~v_173)) & ~v_174)) & ~v_175)) & ~v_176);
	assign v_1655 = (~v_159 & v_177);
	assign v_2074 = (v_177 ^ v_130);
	assign v_1658 = (~v_159 & v_178);
	assign v_2075 = (v_178 ^ v_131);
	assign v_1661 = (~v_159 & v_179);
	assign v_2076 = (v_179 ^ v_132);
	assign v_1664 = (~v_159 & v_180);
	assign v_2077 = (v_180 ^ v_133);
	assign v_1667 = (~v_159 & v_181);
	assign v_2078 = (v_181 ^ v_134);
	assign v_2189 = (((((((~v_177 & ~v_178)) & ~v_179)) & ~v_180)) & ~v_181);
	assign v_1680 = v_18);
	assign v_2080 = (v_182 ^ v_135);
	assign v_2081 = (v_183 ^ v_136);
	assign v_2082 = (v_184 ^ v_137);
	assign v_2083 = (v_185 ^ v_138);
	assign v_1457 = (((((~v_182 & ~v_183)) & ~v_184)) & ~v_185);
	assign v_2085 = (v_186 ^ v_139);
	assign v_2086 = (v_187 ^ v_140);
	assign v_2087 = (v_188 ^ v_142);
	assign v_2088 = (v_189 ^ v_143);
	assign v_2089 = (v_190 ^ v_144);
	assign v_2090 = (v_191 ^ v_145);
	assign v_2091 = (v_192 ^ v_146);
	assign v_1458 = (((((~v_189 & ~v_190)) & ~v_191)) & ~v_192);
	assign v_2093 = (v_193 ^ v_147);
	assign v_1883 = (~v_171 & v_194);
	assign v_2094 = (v_194 ^ v_148);
	assign v_2191 = (((((((~v_186 & ~v_187)) & ~v_188)) & ~v_193)) & ~v_194);
	assign v_2095 = (v_195 ^ v_149);
	assign v_1814 = (v_196 & v_192);
	assign v_1811 = (v_196 & v_191);
	assign v_1808 = (v_196 & v_190);
	assign v_1805 = (v_196 & v_189);
	assign v_1705 = (v_196 & v_185);
	assign v_1702 = (v_196 & v_184);
	assign v_1699 = (v_196 & v_183);
	assign v_1696 = (v_196 & v_182);
	assign v_1825 = (v_196 & v_192);
	assign v_1822 = (v_196 & v_191);
	assign v_1819 = (v_196 & v_190);
	assign v_1816 = (v_196 & v_189);
	assign v_1716 = (v_196 & v_185);
	assign v_1713 = (v_196 & v_184);
	assign v_1710 = (v_196 & v_183);
	assign v_1707 = (v_196 & v_182);
	assign v_1773 = (v_196 & v_187);
	assign v_1760 = (v_196 & v_186);
	assign v_1871 = (~v_196 & v_193);
	assign v_1761 = (v_196 & v_186);
	assign v_1837 = (~v_196 & v_192);
	assign v_1834 = (~v_196 & v_191);
	assign v_1831 = (~v_196 & v_190);
	assign v_1828 = (~v_196 & v_189);
	assign v_1728 = (~v_196 & v_185);
	assign v_1725 = (~v_196 & v_184);
	assign v_1722 = (~v_196 & v_183);
	assign v_1719 = (~v_196 & v_182);
	assign v_1873 = (~v_196 & v_193);
	assign v_1779 = (~v_196 & v_187);
	assign v_1849 = (v_196 & v_192);
	assign v_1846 = (v_196 & v_191);
	assign v_1843 = (v_196 & v_190);
	assign v_1840 = (v_196 & v_189);
	assign v_1740 = (v_196 & v_185);
	assign v_1737 = (v_196 & v_184);
	assign v_1734 = (v_196 & v_183);
	assign v_1731 = (v_196 & v_182);
	assign v_1876 = (v_196 & v_193);
	assign v_1782 = (v_196 & v_187);
	assign v_1766 = (v_196 & v_186);
	assign v_1861 = (~v_196 & v_192);
	assign v_1858 = (~v_196 & v_191);
	assign v_1855 = (~v_196 & v_190);
	assign v_1852 = (~v_196 & v_189);
	assign v_1752 = (~v_196 & v_185);
	assign v_1749 = (~v_196 & v_184);
	assign v_1746 = (~v_196 & v_183);
	assign v_1743 = (~v_196 & v_182);
	assign v_1785 = (~v_196 & v_187);
	assign v_1769 = (~v_196 & v_186);
	assign v_2096 = (v_196 ^ v_150);
	assign v_1795 = (v_197 & v_188);
	assign v_1797 = (v_197 & v_188);
	assign v_1800 = (~v_197 & v_188);
	assign v_2097 = (v_197 ^ v_151);
	assign v_1944 = (~v_169 & v_198);
	assign v_1587 = (v_198 & v_170);
	assign v_1594 = (~v_198 & v_171);
	assign v_1590 = (~v_198 & v_170);
	assign v_2098 = (v_198 ^ v_152);
	assign v_1889 = (~v_199 & v_161);
	assign v_1891 = (v_199 & v_162);
	assign v_1956 = v_19);
	assign v_1894 = (~v_199 & v_163);
	assign v_1897 = (v_199 & v_164);
	assign v_1900 = (~v_199 & v_165);
	assign v_1903 = (v_199 & v_166);
	assign v_1906 = (~v_199 & v_167);
	assign v_1909 = (v_199 & v_168);
	assign v_1973 = (~v_159 & v_199);
	assign v_2099 = (v_199 ^ v_153);
	assign v_1789 = (v_200 & v_188);
	assign v_1980 = (v_197 & v_200);
	assign v_1982 = (v_197 & v_200);
	assign v_1985 = (~v_197 & v_200);
	assign v_2100 = (v_200 ^ v_154);
	assign v_2192 = (((((((~v_195 & ~v_196)) & ~v_197)) & ~v_198)) & ~v_200);
	assign v_1918 = (~v_201 & v_196);
	assign v_1989 = (~v_200 & v_201);
	assign v_1994 = (v_197 & v_201);
	assign v_1996 = (v_197 & v_201);
	assign v_2101 = (v_201 ^ v_155);
	assign v_2005 = (~v_201 & v_202);
	assign v_2007 = (~v_196 & v_202);
	assign v_2009 = (~v_196 & v_202);
	assign v_2014 = (~v_196 & v_202);
	assign v_2017 = (v_196 & v_202);
	assign v_2020 = (~v_196 & v_202);
	assign v_2023 = (v_196 & v_202);
	assign v_1999 = (~v_202 & v_201);
	assign v_2026 = (~v_196 & v_202);
	assign v_1940 = (~v_197 & v_202);
	assign v_2102 = (v_202 ^ v_156);
	assign v_2030 = (~v_169 & v_203);
	assign v_1990 = (~v_203 & v_201);
	assign v_1977 = (~v_200 & v_203);
	assign v_1976 = (~v_203 & v_200);
	assign v_1791 = (~v_203 & v_188);
	assign v_2033 = (~v_198 & v_203);
	assign v_2035 = (~v_198 & v_203);
	assign v_1936 = (~v_197 & v_203);
	assign v_2038 = (v_198 & v_203);
	assign v_2103 = (v_203 ^ v_157);
	assign v_2043 = (v_203 & v_204);
	assign v_2045 = (v_197 & v_204);
	assign v_1595 = (~v_204 & v_171);
	assign v_2049 = (~v_197 & v_204);
	assign v_1951 = (~v_198 & v_204);
	assign v_2104 = (v_204 ^ v_158);
	assign v_2106 = (v_205 ^ v_103);
	assign v_2107 = (v_207 ^ v_105);
	assign v_2108 = (v_208 ^ v_106);
	assign v_2109 = (v_209 ^ v_107);
	assign v_2110 = (v_210 ^ v_108);
	assign v_2111 = (v_211 ^ v_109);
	assign v_2112 = (v_212 ^ v_110);
	assign v_2113 = (v_213 ^ v_111);
	assign v_2114 = (v_214 ^ v_112);
	assign v_2115 = (v_215 ^ v_113);
	assign v_2117 = (v_224 ^ v_122);
	assign v_1586 = v_22);
	assign v_2118 = (v_225 ^ v_123);
	assign v_2119 = (v_226 ^ v_124);
	assign v_2120 = (v_227 ^ v_125);
	assign v_2121 = (v_228 ^ v_126);
	assign v_2122 = (v_229 ^ v_127);
	assign v_2123 = (v_230 ^ v_128);
	assign v_2124 = (v_231 ^ v_129);
	assign v_2125 = (v_232 ^ v_130);
	assign v_2126 = (v_233 ^ v_131);
	assign v_2127 = (v_234 ^ v_132);
	assign v_2128 = (v_235 ^ v_133);
	assign v_2129 = (v_236 ^ v_134);
	assign v_2131 = (v_237 ^ v_135);
	assign v_2132 = (v_238 ^ v_136);
	assign v_2133 = (v_239 ^ v_137);
	assign v_2134 = (v_240 ^ v_138);
	assign v_2136 = (v_241 ^ v_139);
	assign v_2137 = (v_242 ^ v_140);
	assign v_1774 = (v_243 & v_187);
	assign v_1869 = (v_243 & v_193);
	assign v_1926 = (v_196 & v_243);
	assign v_2138 = (v_244 ^ v_142);
	assign v_2139 = (v_245 ^ v_143);
	assign v_2140 = (v_246 ^ v_144);
	assign v_2141 = (v_247 ^ v_145);
	assign v_2142 = (v_248 ^ v_146);
	assign v_2144 = (v_249 ^ v_147);
	assign v_2145 = (v_250 ^ v_148);
	assign v_2146 = (v_251 ^ v_149);
	assign v_2147 = (v_252 ^ v_150);
	assign v_2148 = (v_253 ^ v_151);
	assign v_2149 = (v_254 ^ v_152);
	assign v_2150 = (v_255 ^ v_153);
	assign v_2151 = (v_256 ^ v_154);
	assign v_2152 = (v_257 ^ v_155);
	assign v_2153 = (v_258 ^ v_156);
	assign v_2154 = (v_259 ^ v_157);
	assign v_2155 = (v_260 ^ v_158);
	assign v_261 = (v_2159 & v_2160);
	assign v_268 = (v_11 | v_267);
	assign v_277 = (~v_12 & v_266);
	assign v_348 = (~v_15 & v_347);
	assign v_409 = (v_15 & v_407);
	assign v_408 = (v_407 ^ v_15);
	assign v_262 = (v_2161 & v_2162);
	assign v_488 = (v_25 & v_486);
	assign v_487 = (v_486 ^ v_25);
	assign v_583 = (~v_38 & v_579);
	assign v_568 = (~v_38 & v_566);
	assign v_751 = (v_40 & v_750);
	assign v_394 = (~v_40 & v_393);
	assign v_404 = (v_40 & v_400);
	assign v_696 = (v_695 | v_41);
	assign v_763 = (~v_41 & v_762);
	assign v_596 = (v_595 | ~v_42);
	assign v_726 = v_72);
	assign v_797 = (v_45 & v_795);
	assign v_812 = (v_38 & v_811);
	assign v_806 = (v_44 | v_805);
	assign v_837 = (v_11 | v_836);
	assign v_784 = (v_782 | v_783);
	assign v_744 = v_74);
	assign v_850 = (~v_39 & v_849);
	assign v_402 = (v_46 | v_401);
	assign v_862 = (v_66 | v_861);
	assign v_871 = (~v_67 & v_860);
	assign v_942 = (~v_70 & v_941);
	assign v_1003 = (v_70 & v_1001);
	assign v_1002 = (v_1001 ^ v_70);
	assign v_1082 = (v_80 & v_1080);
	assign v_1081 = (v_1080 ^ v_80);
	assign v_581 = (v_580 | ~v_85);
	assign v_676 = (v_38 & v_675);
	assign v_1177 = (~v_94 & v_1173);
	assign v_1162 = (~v_94 & v_1160);
	assign v_1345 = (v_96 & v_1344);
	assign v_988 = (~v_96 & v_987);
	assign v_998 = (v_96 & v_994);
	assign v_1290 = (v_1289 | v_97);
	assign v_1357 = (~v_97 & v_1356);
	assign v_1190 = (v_1189 | ~v_98);
	assign v_1320 = v_131);
	assign v_1391 = (v_101 & v_1389);
	assign v_1406 = (v_94 & v_1405);
	assign v_1400 = (v_100 | v_1399);
	assign v_1431 = (v_66 | v_1430);
	assign v_1378 = (v_1376 | v_1377);
	assign v_1338 = v_133);
	assign v_1444 = (~v_95 & v_1443);
	assign v_996 = (v_102 | v_995);
	assign v_1175 = (v_1174 | ~v_141);
	assign v_1270 = (v_94 & v_1269);
	assign v_2204 = (((((((~v_2057 & ~v_2058)) & ~v_2059)) & ~v_2060)) & ~v_2061);
	assign v_2205 = (((~v_2062 & ~v_2063)) & ~v_2064);
	assign v_1455 = (v_2186 & v_2187);
	assign v_1462 = (v_169 | v_1461);
	assign v_1471 = (~v_170 & v_1460);
	assign v_2208 = (((((((~v_2055 & ~v_2056)) & ~v_2066)) & ~v_2067)) & ~v_2068);
	assign v_1542 = (~v_173 & v_1541);
	assign v_1603 = (v_173 & v_1601);
	assign v_1602 = (v_1601 ^ v_173);
	assign v_2206 = (((((((~v_2069 & ~v_2070)) & ~v_2071)) & ~v_2072)) & ~v_2073);
	assign v_2207 = (((((((~v_2074 & ~v_2075)) & ~v_2076)) & ~v_2077)) & ~v_2078);
	assign v_1456 = (v_2188 & v_2189);
	assign v_1682 = (v_183 & v_1680);
	assign v_1681 = (v_1680 ^ v_183);
	assign v_2084 = (((((~v_2080 & ~v_2081)) & ~v_2082)) & ~v_2083);
	assign v_2092 = (((((~v_2088 & ~v_2089)) & ~v_2090)) & ~v_2091);
	assign v_2209 = (((((((~v_2085 & ~v_2086)) & ~v_2087)) & ~v_2093)) & ~v_2094);
	assign v_1777 = (~v_196 & v_1773);
	assign v_1762 = (~v_196 & v_1760);
	assign v_1945 = (v_198 & v_1944);
	assign v_1588 = (~v_198 & v_1587);
	assign v_1598 = (v_198 & v_1594);
	assign v_1890 = (v_1889 | v_199);
	assign v_1957 = (~v_199 & v_1956);
	assign v_2210 = (((((((~v_2095 & ~v_2096)) & ~v_2097)) & ~v_2098)) & ~v_2099);
	assign v_1790 = (v_1789 | ~v_200);
	assign v_1920 = v_191);
	assign v_1991 = (v_203 & v_1989);
	assign v_2006 = (v_196 & v_2005);
	assign v_2000 = (v_202 | v_1999);
	assign v_2031 = (v_169 | v_2030);
	assign v_1978 = (v_1976 | v_1977);
	assign v_1938 = v_193);
	assign v_2044 = (~v_197 & v_2043);
	assign v_1596 = (v_204 | v_1595);
	assign v_2211 = (((((((~v_2100 & ~v_2101)) & ~v_2102)) & ~v_2103)) & ~v_2104);
	assign v_2213 = (((((((~v_2108 & ~v_2109)) & ~v_2110)) & ~v_2111)) & ~v_2112);
	assign v_2214 = (((~v_2113 & ~v_2114)) & ~v_2115);
	assign v_2217 = (((((((~v_2106 & ~v_2107)) & ~v_2117)) & ~v_2118)) & ~v_2119);
	assign v_2215 = (((((((~v_2120 & ~v_2121)) & ~v_2122)) & ~v_2123)) & ~v_2124);
	assign v_2216 = (((((((~v_2125 & ~v_2126)) & ~v_2127)) & ~v_2128)) & ~v_2129);
	assign v_2135 = (((((~v_2131 & ~v_2132)) & ~v_2133)) & ~v_2134);
	assign v_1775 = (v_1774 | ~v_243);
	assign v_1870 = (v_196 & v_1869);
	assign v_2143 = (((((~v_2139 & ~v_2140)) & ~v_2141)) & ~v_2142);
	assign v_2218 = (((((((~v_2136 & ~v_2137)) & ~v_2138)) & ~v_2144)) & ~v_2145);
	assign v_2219 = (((((((~v_2146 & ~v_2147)) & ~v_2148)) & ~v_2149)) & ~v_2150);
	assign v_2220 = (((((((~v_2151 & ~v_2152)) & ~v_2153)) & ~v_2154)) & ~v_2155);
	assign v_2166 = (((((((~v_43 & ~v_44)) & ~v_45)) & ~v_46)) & v_261);
	assign v_271 = (~v_13 & v_268);
	assign v_303 = (v_268 & v_10);
	assign v_302 = (~v_268 & v_65);
	assign v_300 = (v_268 & v_9);
	assign v_299 = (~v_268 & v_64);
	assign v_297 = (v_268 & v_8);
	assign v_296 = (~v_268 & v_63);
	assign v_294 = (v_268 & v_7);
	assign v_293 = (~v_268 & v_62);
	assign v_291 = (v_268 & v_6);
	assign v_290 = (~v_268 & v_61);
	assign v_288 = (v_268 & v_5);
	assign v_287 = (~v_268 & v_60);
	assign v_285 = (v_268 & v_4);
	assign v_284 = (~v_268 & v_59);
	assign v_282 = (v_268 & v_3);
	assign v_281 = (~v_268 & v_58);
	assign v_688 = (v_13 & v_268);
	assign v_349 = v_34);
	assign v_410 = v_40);
	assign v_2167 = (((((v_262 & v_263)) & v_264)) & v_41);
	assign v_489 = v_48);
	assign v_569 = (v_567 | v_568);
	assign v_753 = v_75);
	assign v_395 = (v_40 | v_394);
	assign v_698 = (~v_41 & v_696);
	assign v_764 = (v_41 & v_763);
	assign v_598 = (v_45 & v_596);
	assign v_727 = (v_38 & v_726);
	assign v_798 = (v_796 | v_797);
	assign v_814 = (v_812 | v_813);
	assign v_807 = (~v_39 & v_806);
	assign v_838 = (v_40 & v_837);
	assign v_785 = (~v_39 & v_784);
	assign v_745 = (~v_39 & v_744);
	assign v_852 = (v_850 | v_851);
	assign v_403 = (~v_40 & v_402);
	assign v_865 = (~v_68 & v_862);
	assign v_897 = (v_862 & v_57);
	assign v_896 = (~v_862 & v_121);
	assign v_894 = (v_862 & v_56);
	assign v_893 = (~v_862 & v_120);
	assign v_891 = (v_862 & v_55);
	assign v_890 = (~v_862 & v_119);
	assign v_888 = (v_862 & v_54);
	assign v_887 = (~v_862 & v_118);
	assign v_885 = (v_862 & v_53);
	assign v_884 = (~v_862 & v_117);
	assign v_882 = (v_862 & v_52);
	assign v_881 = (~v_862 & v_116);
	assign v_879 = (v_862 & v_51);
	assign v_878 = (~v_862 & v_115);
	assign v_876 = (v_862 & v_50);
	assign v_875 = (~v_862 & v_114);
	assign v_1282 = (v_68 & v_862);
	assign v_943 = v_94);
	assign v_1004 = v_100);
	assign v_1083 = v_108);
	assign v_582 = (v_38 & v_581);
	assign v_678 = (v_676 | v_677);
	assign v_1163 = (v_1161 | v_1162);
	assign v_1347 = v_134);
	assign v_989 = (v_96 | v_988);
	assign v_1292 = (~v_97 & v_1290);
	assign v_1358 = (v_97 & v_1357);
	assign v_1192 = (v_101 & v_1190);
	assign v_1321 = (v_94 & v_1320);
	assign v_1392 = (v_1390 | v_1391);
	assign v_1408 = (v_1406 | v_1407);
	assign v_1401 = (~v_95 & v_1400);
	assign v_1432 = (v_96 & v_1431);
	assign v_1379 = (~v_95 & v_1378);
	assign v_1339 = (~v_95 & v_1338);
	assign v_1446 = (v_1444 | v_1445);
	assign v_997 = (~v_96 & v_996);
	assign v_1176 = (v_94 & v_1175);
	assign v_1272 = (v_1270 | v_1271);
	assign v_2065 = (v_2204 & v_2205);
	assign v_2193 = (((((((~v_201 & ~v_202)) & ~v_203)) & ~v_204)) & v_1455);
	assign v_1465 = (~v_171 & v_1462);
	assign v_1497 = (v_1462 & v_168);
	assign v_1496 = (~v_1462 & v_223);
	assign v_1494 = (v_1462 & v_167);
	assign v_1493 = (~v_1462 & v_222);
	assign v_1491 = (v_1462 & v_166);
	assign v_1490 = (~v_1462 & v_221);
	assign v_1488 = (v_1462 & v_165);
	assign v_1487 = (~v_1462 & v_220);
	assign v_1485 = (v_1462 & v_164);
	assign v_1484 = (~v_1462 & v_219);
	assign v_1482 = (v_1462 & v_163);
	assign v_1481 = (~v_1462 & v_218);
	assign v_1479 = (v_1462 & v_162);
	assign v_1478 = (~v_1462 & v_217);
	assign v_1476 = (v_1462 & v_161);
	assign v_1475 = (~v_1462 & v_216);
	assign v_1882 = (v_171 & v_1462);
	assign v_1543 = v_154);
	assign v_1604 = v_160);
	assign v_2079 = (v_2206 & v_2207);
	assign v_2194 = (((((v_1456 & v_1457)) & v_1458)) & v_199);
	assign v_1683 = v_168);
	assign v_1763 = (v_1761 | v_1762);
	assign v_1947 = v_194);
	assign v_1589 = (v_198 | v_1588);
	assign v_1892 = (~v_199 & v_1890);
	assign v_1958 = (v_199 & v_1957);
	assign v_1792 = (v_203 & v_1790);
	assign v_1921 = (v_196 & v_1920);
	assign v_1992 = (v_1990 | v_1991);
	assign v_2008 = (v_2006 | v_2007);
	assign v_2001 = (~v_197 & v_2000);
	assign v_2032 = (v_198 & v_2031);
	assign v_1979 = (~v_197 & v_1978);
	assign v_1939 = (~v_197 & v_1938);
	assign v_2046 = (v_2044 | v_2045);
	assign v_1597 = (~v_198 & v_1596);
	assign v_2116 = (v_2213 & v_2214);
	assign v_2130 = (v_2215 & v_2216);
	assign v_1776 = (v_196 & v_1775);
	assign v_1872 = (v_1870 | v_1871);
	assign v_272 = (v_270 | v_271);
	assign v_304 = (v_302 | v_303);
	assign v_301 = (v_299 | v_300);
	assign v_298 = (v_296 | v_297);
	assign v_295 = (v_293 | v_294);
	assign v_292 = (v_290 | v_291);
	assign v_289 = (v_287 | v_288);
	assign v_286 = (v_284 | v_285);
	assign v_283 = (v_281 | v_282);
	assign v_690 = (v_688 | v_689);
	assign v_350 = (~v_16 & v_349);
	assign v_412 = (v_16 & v_410);
	assign v_411 = (v_410 ^ v_16);
	assign v_265 = (((((((v_2163 & v_2164)) & v_2165)) & v_2166)) & v_2167);
	assign v_491 = (v_26 & v_489);
	assign v_490 = (v_489 ^ v_26);
	assign v_570 = (v_38 & v_569);
	assign v_754 = (v_40 & v_753);
	assign v_397 = (v_40 & v_395);
	assign v_699 = (v_697 | v_698);
	assign v_765 = (v_764 | ~v_41);
	assign v_599 = (v_597 | v_598);
	assign v_728 = (v_727 | ~v_38);
	assign v_799 = (~v_39 & v_798);
	assign v_816 = (v_38 & v_814);
	assign v_840 = (v_838 | v_839);
	assign v_787 = (v_785 | v_786);
	assign v_747 = (v_39 & v_745);
	assign v_853 = (~v_39 & v_852);
	assign v_405 = (v_403 | v_404);
	assign v_866 = (v_864 | v_865);
	assign v_898 = (v_896 | v_897);
	assign v_895 = (v_893 | v_894);
	assign v_892 = (v_890 | v_891);
	assign v_889 = (v_887 | v_888);
	assign v_886 = (v_884 | v_885);
	assign v_883 = (v_881 | v_882);
	assign v_880 = (v_878 | v_879);
	assign v_877 = (v_875 | v_876);
	assign v_1284 = (v_1282 | v_1283);
	assign v_944 = (~v_71 & v_943);
	assign v_1006 = (v_71 & v_1004);
	assign v_1005 = (v_1004 ^ v_71);
	assign v_1085 = (v_81 & v_1083);
	assign v_1084 = (v_1083 ^ v_81);
	assign v_584 = (v_582 | v_583);
	assign v_680 = (v_38 & v_678);
	assign v_1164 = (v_94 & v_1163);
	assign v_1348 = (v_96 & v_1347);
	assign v_991 = (v_96 & v_989);
	assign v_1293 = (v_1291 | v_1292);
	assign v_1359 = (v_1358 | ~v_97);
	assign v_1193 = (v_1191 | v_1192);
	assign v_1322 = (v_1321 | ~v_94);
	assign v_1393 = (~v_95 & v_1392);
	assign v_1410 = (v_94 & v_1408);
	assign v_1434 = (v_1432 | v_1433);
	assign v_1381 = (v_1379 | v_1380);
	assign v_1341 = (v_95 & v_1339);
	assign v_1447 = (~v_95 & v_1446);
	assign v_999 = (v_997 | v_998);
	assign v_1178 = (v_1176 | v_1177);
	assign v_1274 = (v_94 & v_1272);
	assign v_1466 = (v_1464 | v_1465);
	assign v_1498 = (v_1496 | v_1497);
	assign v_1495 = (v_1493 | v_1494);
	assign v_1492 = (v_1490 | v_1491);
	assign v_1489 = (v_1487 | v_1488);
	assign v_1486 = (v_1484 | v_1485);
	assign v_1483 = (v_1481 | v_1482);
	assign v_1480 = (v_1478 | v_1479);
	assign v_1477 = (v_1475 | v_1476);
	assign v_1884 = (v_1882 | v_1883);
	assign v_1544 = (~v_174 & v_1543);
	assign v_1606 = (v_174 & v_1604);
	assign v_1605 = (v_1604 ^ v_174);
	assign v_2212 = (((((v_2065 & v_2079)) & v_2084)) & v_2092);
	assign v_1459 = (((((((v_2190 & v_2191)) & v_2192)) & v_2193)) & v_2194);
	assign v_1685 = (v_184 & v_1683);
	assign v_1684 = (v_1683 ^ v_184);
	assign v_1764 = (v_196 & v_1763);
	assign v_1948 = (v_198 & v_1947);
	assign v_1591 = (v_198 & v_1589);
	assign v_1893 = (v_1891 | v_1892);
	assign v_1959 = (v_1958 | ~v_199);
	assign v_1793 = (v_1791 | v_1792);
	assign v_1922 = (v_1921 | ~v_196);
	assign v_1993 = (~v_197 & v_1992);
	assign v_2010 = (v_196 & v_2008);
	assign v_2034 = (v_2032 | v_2033);
	assign v_1981 = (v_1979 | v_1980);
	assign v_1941 = (v_197 & v_1939);
	assign v_2047 = (~v_197 & v_2046);
	assign v_1599 = (v_1597 | v_1598);
	assign v_2221 = (((((v_2116 & v_2130)) & v_2135)) & v_2143);
	assign v_1778 = (v_1776 | v_1777);
	assign v_1874 = (v_196 & v_1872);
	assign v_273 = (~v_272 | ~v_48);
	assign v_280 = (v_272 ^ v_49);
	assign v_326 = (v_13 & v_304);
	assign v_323 = (v_13 & v_301);
	assign v_320 = (v_13 & v_298);
	assign v_317 = (v_13 & v_295);
	assign v_314 = (v_13 & v_292);
	assign v_311 = (v_13 & v_289);
	assign v_308 = (v_13 & v_286);
	assign v_305 = (v_13 & v_283);
	assign v_692 = (~v_12 & v_690);
	assign v_351 = v_35);
	assign v_413 = v_41);
	assign v_492 = v_49);
	assign v_571 = (v_570 | ~v_38);
	assign v_755 = (v_754 | ~v_40);
	assign v_398 = (v_396 | v_397);
	assign v_701 = (v_41 & v_699);
	assign v_766 = (~v_41 & v_765);
	assign v_600 = (~v_39 & v_599);
	assign v_729 = (~v_38 & v_728);
	assign v_801 = (v_799 | v_800);
	assign v_817 = (v_815 | v_816);
	assign v_842 = (v_40 & v_840);
	assign v_789 = (~v_39 & v_787);
	assign v_748 = (v_746 | v_747);
	assign v_854 = (v_39 | v_853);
	assign v_406 = (v_405 ^ v_68);
	assign v_867 = (~v_866 | ~v_104);
	assign v_874 = (v_866 ^ v_105);
	assign v_920 = (v_68 & v_898);
	assign v_917 = (v_68 & v_895);
	assign v_914 = (v_68 & v_892);
	assign v_911 = (v_68 & v_889);
	assign v_908 = (v_68 & v_886);
	assign v_905 = (v_68 & v_883);
	assign v_902 = (v_68 & v_880);
	assign v_899 = (v_68 & v_877);
	assign v_1286 = (~v_67 & v_1284);
	assign v_945 = v_94);
	assign v_1007 = v_100);
	assign v_1086 = v_108);
	assign v_586 = (v_38 & v_584);
	assign v_681 = (v_679 | v_680);
	assign v_1165 = (v_1164 | ~v_94);
	assign v_1349 = (v_1348 | ~v_96);
	assign v_992 = (v_990 | v_991);
	assign v_1295 = (v_97 & v_1293);
	assign v_1360 = (~v_97 & v_1359);
	assign v_1194 = (~v_95 & v_1193);
	assign v_1323 = (~v_94 & v_1322);
	assign v_1395 = (v_1393 | v_1394);
	assign v_1411 = (v_1409 | v_1410);
	assign v_1436 = (v_96 & v_1434);
	assign v_1383 = (~v_95 & v_1381);
	assign v_1342 = (v_1340 | v_1341);
	assign v_1448 = (v_95 | v_1447);
	assign v_1000 = (v_999 ^ v_124);
	assign v_1180 = (v_94 & v_1178);
	assign v_1275 = (v_1273 | v_1274);
	assign v_1467 = (~v_1466 | ~v_206);
	assign v_1474 = (v_1466 ^ v_207);
	assign v_1520 = (v_171 & v_1498);
	assign v_1517 = (v_171 & v_1495);
	assign v_1514 = (v_171 & v_1492);
	assign v_1511 = (v_171 & v_1489);
	assign v_1508 = (v_171 & v_1486);
	assign v_1505 = (v_171 & v_1483);
	assign v_1502 = (v_171 & v_1480);
	assign v_1499 = (v_171 & v_1477);
	assign v_1886 = (~v_170 & v_1884);
	assign v_1545 = v_154);
	assign v_1607 = v_160);
	assign v_2105 = (((((((v_2208 & v_2209)) & v_2210)) & v_2211)) & v_2212);
	assign v_1686 = v_168);
	assign v_1765 = (v_1764 | ~v_196);
	assign v_1949 = (v_1948 | ~v_198);
	assign v_1592 = (v_1590 | v_1591);
	assign v_1895 = (v_199 & v_1893);
	assign v_1960 = (~v_199 & v_1959);
	assign v_1794 = (~v_197 & v_1793);
	assign v_1923 = (~v_196 & v_1922);
	assign v_1995 = (v_1993 | v_1994);
	assign v_2011 = (v_2009 | v_2010);
	assign v_2036 = (v_198 & v_2034);
	assign v_1983 = (~v_197 & v_1981);
	assign v_1942 = (v_1940 | v_1941);
	assign v_2048 = (v_197 | v_2047);
	assign v_1600 = (v_1599 ^ v_226);
	assign v_2156 = (((((((v_2217 & v_2218)) & v_2219)) & v_2220)) & v_2221);
	assign v_1780 = (v_196 & v_1778);
	assign v_1875 = (v_1873 | v_1874);
	assign v_274 = (v_273 & v_266);
	assign v_691 = (v_12 & v_273);
	assign v_328 = (v_326 | v_327);
	assign v_325 = (v_323 | v_324);
	assign v_322 = (v_320 | v_321);
	assign v_319 = (v_317 | v_318);
	assign v_316 = (v_314 | v_315);
	assign v_313 = (v_311 | v_312);
	assign v_310 = (v_308 | v_309);
	assign v_307 = (v_305 | v_306);
	assign v_352 = (~v_17 & v_351);
	assign v_415 = (v_17 & v_413);
	assign v_414 = (v_413 ^ v_17);
	assign v_493 = (v_492 ^ v_27);
	assign v_494 = (v_27 & v_492);
	assign v_573 = (~v_38 & v_571);
	assign v_756 = (~v_40 & v_755);
	assign v_399 = (v_398 ^ v_67);
	assign v_702 = (v_700 | v_701);
	assign v_767 = (v_41 & v_766);
	assign v_602 = (v_600 | v_601);
	assign v_730 = (v_38 & v_729);
	assign v_803 = (~v_39 & v_801);
	assign v_818 = (~v_38 & v_817);
	assign v_843 = (v_841 | v_842);
	assign v_790 = (v_788 | v_789);
	assign v_749 = (v_748 ^ v_95);
	assign v_856 = (v_39 & v_854);
	assign v_868 = (v_867 & v_860);
	assign v_1285 = (v_67 & v_867);
	assign v_922 = (v_920 | v_921);
	assign v_919 = (v_917 | v_918);
	assign v_916 = (v_914 | v_915);
	assign v_913 = (v_911 | v_912);
	assign v_910 = (v_908 | v_909);
	assign v_907 = (v_905 | v_906);
	assign v_904 = (v_902 | v_903);
	assign v_901 = (v_899 | v_900);
	assign v_946 = (~v_72 & v_945);
	assign v_1009 = (v_72 & v_1007);
	assign v_1008 = (v_1007 ^ v_72);
	assign v_1087 = (v_1086 ^ v_82);
	assign v_1088 = (v_82 & v_1086);
	assign v_587 = (v_585 | v_586);
	assign v_683 = (~v_38 & v_681);
	assign v_1167 = (~v_94 & v_1165);
	assign v_1350 = (~v_96 & v_1349);
	assign v_993 = (v_992 ^ v_123);
	assign v_1296 = (v_1294 | v_1295);
	assign v_1361 = (v_97 & v_1360);
	assign v_1196 = (v_1194 | v_1195);
	assign v_1324 = (v_94 & v_1323);
	assign v_1397 = (~v_95 & v_1395);
	assign v_1412 = (~v_94 & v_1411);
	assign v_1437 = (v_1435 | v_1436);
	assign v_1384 = (v_1382 | v_1383);
	assign v_1343 = (v_1342 ^ v_151);
	assign v_1450 = (v_95 & v_1448);
	assign v_1181 = (v_1179 | v_1180);
	assign v_1277 = (~v_94 & v_1275);
	assign v_1468 = (v_1467 & v_1460);
	assign v_1885 = (v_170 & v_1467);
	assign v_1522 = (v_1520 | v_1521);
	assign v_1519 = (v_1517 | v_1518);
	assign v_1516 = (v_1514 | v_1515);
	assign v_1513 = (v_1511 | v_1512);
	assign v_1510 = (v_1508 | v_1509);
	assign v_1507 = (v_1505 | v_1506);
	assign v_1504 = (v_1502 | v_1503);
	assign v_1501 = (v_1499 | v_1500);
	assign v_1546 = (~v_175 & v_1545);
	assign v_1609 = (v_175 & v_1607);
	assign v_1608 = (v_1607 ^ v_175);
	assign v_1687 = (v_1686 ^ v_185);
	assign v_1688 = (v_185 & v_1686);
	assign v_1767 = (~v_196 & v_1765);
	assign v_1950 = (~v_198 & v_1949);
	assign v_1593 = (v_1592 ^ v_225);
	assign v_1896 = (v_1894 | v_1895);
	assign v_1961 = (v_199 & v_1960);
	assign v_1796 = (v_1794 | v_1795);
	assign v_1924 = (v_196 & v_1923);
	assign v_1997 = (~v_197 & v_1995);
	assign v_2012 = (~v_196 & v_2011);
	assign v_2037 = (v_2035 | v_2036);
	assign v_1984 = (v_1982 | v_1983);
	assign v_1943 = (v_1942 ^ v_253);
	assign v_2050 = (v_197 & v_2048);
	assign v_2157 = (v_2105 | v_2156);
	assign v_1781 = (v_1779 | v_1780);
	assign v_1877 = (~v_196 & v_1875);
	assign v_275 = (v_274 | ~v_273);
	assign v_693 = (v_691 | v_692);
	assign v_336 = (v_328 ^ v_57);
	assign v_335 = (v_325 ^ v_56);
	assign v_334 = (v_322 ^ v_55);
	assign v_333 = (v_319 ^ v_54);
	assign v_332 = (v_316 ^ v_53);
	assign v_331 = (v_313 ^ v_52);
	assign v_330 = (v_310 ^ v_51);
	assign v_329 = (v_307 ^ v_50);
	assign v_353 = (((v_351 | v_352)) | ~v_17);
	assign v_416 = v_41);
	assign v_496 = (((((~v_487 & ~v_490)) & v_24)) & v_493);
	assign v_495 = v_49);
	assign v_574 = (v_572 | v_573);
	assign v_758 = (v_40 & v_756);
	assign v_704 = (~v_41 & v_702);
	assign v_768 = (v_767 | ~v_41);
	assign v_604 = (~v_39 & v_602);
	assign v_731 = (v_730 | ~v_38);
	assign v_804 = (v_802 | v_803);
	assign v_819 = (v_38 | v_818);
	assign v_845 = (~v_40 & v_843);
	assign v_792 = (v_39 & v_790);
	assign v_857 = (v_855 | v_856);
	assign v_869 = (v_868 | ~v_867);
	assign v_1287 = (v_1285 | v_1286);
	assign v_930 = (v_922 ^ v_113);
	assign v_929 = (v_919 ^ v_112);
	assign v_928 = (v_916 ^ v_111);
	assign v_927 = (v_913 ^ v_110);
	assign v_926 = (v_910 ^ v_109);
	assign v_925 = (v_907 ^ v_108);
	assign v_924 = (v_904 ^ v_107);
	assign v_923 = (v_901 ^ v_106);
	assign v_947 = (((v_945 | v_946)) | ~v_72);
	assign v_1010 = v_100);
	assign v_1090 = (((((~v_1081 & ~v_1084)) & v_79)) & v_1087);
	assign v_1089 = v_108);
	assign v_589 = (~v_38 & v_587);
	assign v_684 = (v_682 | v_683);
	assign v_1168 = (v_1166 | v_1167);
	assign v_1352 = (v_96 & v_1350);
	assign v_1298 = (~v_97 & v_1296);
	assign v_1362 = (v_1361 | ~v_97);
	assign v_1198 = (~v_95 & v_1196);
	assign v_1325 = (v_1324 | ~v_94);
	assign v_1398 = (v_1396 | v_1397);
	assign v_1413 = (v_94 | v_1412);
	assign v_1439 = (~v_96 & v_1437);
	assign v_1386 = (v_95 & v_1384);
	assign v_1451 = (v_1449 | v_1450);
	assign v_1183 = (~v_94 & v_1181);
	assign v_1278 = (v_1276 | v_1277);
	assign v_1469 = (v_1468 | ~v_1467);
	assign v_1887 = (v_1885 | v_1886);
	assign v_1530 = (v_1522 ^ v_215);
	assign v_1529 = (v_1519 ^ v_214);
	assign v_1528 = (v_1516 ^ v_213);
	assign v_1527 = (v_1513 ^ v_212);
	assign v_1526 = (v_1510 ^ v_211);
	assign v_1525 = (v_1507 ^ v_210);
	assign v_1524 = (v_1504 ^ v_209);
	assign v_1523 = (v_1501 ^ v_208);
	assign v_1547 = (((v_1545 | v_1546)) | ~v_175);
	assign v_1610 = v_160);
	assign v_1690 = (((((~v_1681 & ~v_1684)) & v_182)) & v_1687);
	assign v_1689 = v_168);
	assign v_1768 = (v_1766 | v_1767);
	assign v_1952 = (v_198 & v_1950);
	assign v_1898 = (~v_199 & v_1896);
	assign v_1962 = (v_1961 | ~v_199);
	assign v_1798 = (~v_197 & v_1796);
	assign v_1925 = (v_1924 | ~v_196);
	assign v_1998 = (v_1996 | v_1997);
	assign v_2013 = (v_196 | v_2012);
	assign v_2039 = (~v_198 & v_2037);
	assign v_1986 = (v_197 & v_1984);
	assign v_2051 = (v_2049 | v_2050);
	assign v_1783 = (~v_196 & v_1781);
	assign v_1878 = (v_1876 | v_1877);
	assign v_276 = (v_12 & v_275);
	assign v_694 = (v_693 ^ v_92);
	assign v_2169 = (((~v_334 & ~v_335)) & ~v_336);
	assign v_2168 = (((((((~v_329 & ~v_330)) & ~v_331)) & ~v_332)) & ~v_333);
	assign v_354 = (~v_18 & v_353);
	assign v_418 = (v_18 & v_416);
	assign v_417 = (v_416 ^ v_18);
	assign v_500 = (~v_496 & v_493);
	assign v_499 = (~v_496 & v_490);
	assign v_498 = (~v_496 & v_487);
	assign v_497 = (~v_496 & ~v_24);
	assign v_576 = (v_38 & v_574);
	assign v_759 = (v_757 | v_758);
	assign v_705 = (v_703 | v_704);
	assign v_769 = (~v_41 & v_768);
	assign v_605 = (v_603 | v_604);
	assign v_733 = (~v_38 & v_731);
	assign v_808 = (v_39 & v_804);
	assign v_821 = (v_38 & v_819);
	assign v_846 = (v_844 | v_845);
	assign v_793 = (v_791 | v_792);
	assign v_858 = (v_857 ^ v_102);
	assign v_870 = (v_67 & v_869);
	assign v_1288 = (v_1287 ^ v_148);
	assign v_2178 = (((~v_928 & ~v_929)) & ~v_930);
	assign v_2177 = (((((((~v_923 & ~v_924)) & ~v_925)) & ~v_926)) & ~v_927);
	assign v_948 = (~v_73 & v_947);
	assign v_1012 = (v_73 & v_1010);
	assign v_1011 = (v_1010 ^ v_73);
	assign v_1094 = (~v_1090 & v_1087);
	assign v_1093 = (~v_1090 & v_1084);
	assign v_1092 = (~v_1090 & v_1081);
	assign v_1091 = (~v_1090 & ~v_79);
	assign v_590 = (v_588 | v_589);
	assign v_685 = (v_38 & v_684);
	assign v_1170 = (v_94 & v_1168);
	assign v_1353 = (v_1351 | v_1352);
	assign v_1299 = (v_1297 | v_1298);
	assign v_1363 = (~v_97 & v_1362);
	assign v_1199 = (v_1197 | v_1198);
	assign v_1327 = (~v_94 & v_1325);
	assign v_1402 = (v_95 & v_1398);
	assign v_1415 = (v_94 & v_1413);
	assign v_1440 = (v_1438 | v_1439);
	assign v_1387 = (v_1385 | v_1386);
	assign v_1452 = (v_1451 ^ v_158);
	assign v_1184 = (v_1182 | v_1183);
	assign v_1279 = (v_94 & v_1278);
	assign v_1470 = (v_170 & v_1469);
	assign v_1888 = (v_1887 ^ v_250);
	assign v_2196 = (((~v_1528 & ~v_1529)) & ~v_1530);
	assign v_2195 = (((((((~v_1523 & ~v_1524)) & ~v_1525)) & ~v_1526)) & ~v_1527);
	assign v_1548 = (~v_176 & v_1547);
	assign v_1612 = (v_176 & v_1610);
	assign v_1611 = (v_1610 ^ v_176);
	assign v_1694 = (~v_1690 & v_1687);
	assign v_1693 = (~v_1690 & v_1684);
	assign v_1692 = (~v_1690 & v_1681);
	assign v_1691 = (~v_1690 & ~v_182);
	assign v_1770 = (v_196 & v_1768);
	assign v_1953 = (v_1951 | v_1952);
	assign v_1899 = (v_1897 | v_1898);
	assign v_1963 = (~v_199 & v_1962);
	assign v_1799 = (v_1797 | v_1798);
	assign v_1927 = (~v_196 & v_1925);
	assign v_2002 = (v_197 & v_1998);
	assign v_2015 = (v_196 & v_2013);
	assign v_2040 = (v_2038 | v_2039);
	assign v_1987 = (v_1985 | v_1986);
	assign v_2052 = (v_2051 ^ v_260);
	assign v_1784 = (v_1782 | v_1783);
	assign v_1879 = (v_196 & v_1878);
	assign v_278 = (v_276 | v_277);
	assign v_337 = (v_2168 & v_2169);
	assign v_355 = v_35);
	assign v_419 = v_41);
	assign v_619 = (~v_38 & v_500);
	assign v_510 = (~v_38 & v_500);
	assign v_616 = (~v_38 & v_499);
	assign v_507 = (~v_38 & v_499);
	assign v_613 = (~v_38 & v_498);
	assign v_504 = (~v_38 & v_498);
	assign v_610 = (~v_38 & v_497);
	assign v_501 = (~v_38 & v_497);
	assign v_577 = (v_575 | v_576);
	assign v_760 = (v_759 ^ v_96);
	assign v_707 = (v_41 & v_705);
	assign v_770 = (v_41 & v_769);
	assign v_607 = (v_39 & v_605);
	assign v_734 = (v_732 | v_733);
	assign v_809 = (v_807 | v_808);
	assign v_822 = (v_820 | v_821);
	assign v_847 = (v_40 & v_846);
	assign v_794 = (v_793 ^ v_98);
	assign v_872 = (v_870 | v_871);
	assign v_931 = (v_2177 & v_2178);
	assign v_949 = v_94);
	assign v_1013 = v_101);
	assign v_1213 = (~v_94 & v_1094);
	assign v_1104 = (~v_94 & v_1094);
	assign v_1210 = (~v_94 & v_1093);
	assign v_1101 = (~v_94 & v_1093);
	assign v_1207 = (~v_94 & v_1092);
	assign v_1098 = (~v_94 & v_1092);
	assign v_1204 = (~v_94 & v_1091);
	assign v_1095 = (~v_94 & v_1091);
	assign v_592 = (v_38 & v_590);
	assign v_686 = (v_685 | ~v_38);
	assign v_1171 = (v_1169 | v_1170);
	assign v_1354 = (v_1353 ^ v_152);
	assign v_1301 = (v_97 & v_1299);
	assign v_1364 = (v_97 & v_1363);
	assign v_1201 = (v_95 & v_1199);
	assign v_1328 = (v_1326 | v_1327);
	assign v_1403 = (v_1401 | v_1402);
	assign v_1416 = (v_1414 | v_1415);
	assign v_1441 = (v_96 & v_1440);
	assign v_1388 = (v_1387 ^ v_154);
	assign v_1186 = (v_94 & v_1184);
	assign v_1280 = (v_1279 | ~v_94);
	assign v_1472 = (v_1470 | v_1471);
	assign v_1531 = (v_2195 & v_2196);
	assign v_1549 = v_154);
	assign v_1613 = v_161);
	assign v_1813 = (~v_196 & v_1694);
	assign v_1704 = (~v_196 & v_1694);
	assign v_1810 = (~v_196 & v_1693);
	assign v_1701 = (~v_196 & v_1693);
	assign v_1807 = (~v_196 & v_1692);
	assign v_1698 = (~v_196 & v_1692);
	assign v_1804 = (~v_196 & v_1691);
	assign v_1695 = (~v_196 & v_1691);
	assign v_1771 = (v_1769 | v_1770);
	assign v_1954 = (v_1953 ^ v_254);
	assign v_1901 = (v_199 & v_1899);
	assign v_1964 = (v_199 & v_1963);
	assign v_1801 = (v_197 & v_1799);
	assign v_1928 = (v_1926 | v_1927);
	assign v_2003 = (v_2001 | v_2002);
	assign v_2016 = (v_2014 | v_2015);
	assign v_2041 = (v_198 & v_2040);
	assign v_1988 = (v_1987 ^ v_256);
	assign v_1786 = (v_196 & v_1784);
	assign v_1880 = (v_1879 | ~v_196);
	assign v_279 = (v_278 ^ v_47);
	assign v_356 = (~v_19 & v_355);
	assign v_421 = (v_19 & v_419);
	assign v_420 = (v_419 ^ v_19);
	assign v_621 = (v_619 | v_620);
	assign v_512 = (v_510 | v_511);
	assign v_618 = (v_616 | v_617);
	assign v_509 = (v_507 | v_508);
	assign v_615 = (v_613 | v_614);
	assign v_506 = (v_504 | v_505);
	assign v_612 = (v_610 | v_611);
	assign v_503 = (v_501 | v_502);
	assign v_578 = (v_577 ^ v_83);
	assign v_708 = (v_706 | v_707);
	assign v_771 = (v_770 | ~v_41);
	assign v_608 = (v_606 | v_607);
	assign v_735 = (v_38 & v_734);
	assign v_810 = (v_809 ^ v_99);
	assign v_824 = (~v_38 & v_822);
	assign v_848 = (v_847 ^ v_101);
	assign v_873 = (v_872 ^ v_103);
	assign v_950 = (~v_74 & v_949);
	assign v_1015 = (v_74 & v_1013);
	assign v_1014 = (v_1013 ^ v_74);
	assign v_1215 = (v_1213 | v_1214);
	assign v_1106 = (v_1104 | v_1105);
	assign v_1212 = (v_1210 | v_1211);
	assign v_1103 = (v_1101 | v_1102);
	assign v_1209 = (v_1207 | v_1208);
	assign v_1100 = (v_1098 | v_1099);
	assign v_1206 = (v_1204 | v_1205);
	assign v_1097 = (v_1095 | v_1096);
	assign v_593 = (v_591 | v_592);
	assign v_687 = (v_686 ^ v_91);
	assign v_1172 = (v_1171 ^ v_139);
	assign v_1302 = (v_1300 | v_1301);
	assign v_1365 = (v_1364 | ~v_97);
	assign v_1202 = (v_1200 | v_1201);
	assign v_1329 = (v_94 & v_1328);
	assign v_1404 = (v_1403 ^ v_155);
	assign v_1418 = (~v_94 & v_1416);
	assign v_1442 = (v_1441 ^ v_157);
	assign v_1187 = (v_1185 | v_1186);
	assign v_1281 = (v_1280 ^ v_147);
	assign v_1473 = (v_1472 ^ v_205);
	assign v_1550 = (~v_177 & v_1549);
	assign v_1615 = (v_177 & v_1613);
	assign v_1614 = (v_1613 ^ v_177);
	assign v_1815 = (v_1813 | v_1814);
	assign v_1706 = (v_1704 | v_1705);
	assign v_1812 = (v_1810 | v_1811);
	assign v_1703 = (v_1701 | v_1702);
	assign v_1809 = (v_1807 | v_1808);
	assign v_1700 = (v_1698 | v_1699);
	assign v_1806 = (v_1804 | v_1805);
	assign v_1697 = (v_1695 | v_1696);
	assign v_1772 = (v_1771 ^ v_241);
	assign v_1902 = (v_1900 | v_1901);
	assign v_1965 = (v_1964 | ~v_199);
	assign v_1802 = (v_1800 | v_1801);
	assign v_1929 = (v_196 & v_1928);
	assign v_2004 = (v_2003 ^ v_257);
	assign v_2018 = (~v_196 & v_2016);
	assign v_2042 = (v_2041 ^ v_259);
	assign v_1787 = (v_1785 | v_1786);
	assign v_1881 = (v_1880 ^ v_249);
	assign v_2172 = (((((((~v_279 & ~v_280)) & ~v_392)) & ~v_399)) & ~v_406);
	assign v_357 = (((v_355 | v_356)) | ~v_19);
	assign v_422 = v_42);
	assign v_632 = (~v_38 & v_621);
	assign v_523 = (~v_38 & v_512);
	assign v_629 = (~v_38 & v_618);
	assign v_520 = (~v_38 & v_509);
	assign v_626 = (~v_38 & v_615);
	assign v_517 = (~v_38 & v_506);
	assign v_623 = (~v_38 & v_612);
	assign v_514 = (~v_38 & v_503);
	assign v_710 = (~v_41 & v_708);
	assign v_772 = (~v_41 & v_771);
	assign v_609 = (v_608 ^ v_86);
	assign v_736 = (v_735 | ~v_38);
	assign v_825 = (v_823 | v_824);
	assign v_2181 = (((((((~v_873 & ~v_874)) & ~v_986)) & ~v_993)) & ~v_1000);
	assign v_951 = (((v_949 | v_950)) | ~v_74);
	assign v_1016 = v_101);
	assign v_1226 = (~v_94 & v_1215);
	assign v_1117 = (~v_94 & v_1106);
	assign v_1223 = (~v_94 & v_1212);
	assign v_1114 = (~v_94 & v_1103);
	assign v_1220 = (~v_94 & v_1209);
	assign v_1111 = (~v_94 & v_1100);
	assign v_1217 = (~v_94 & v_1206);
	assign v_1108 = (~v_94 & v_1097);
	assign v_594 = (v_593 ^ v_84);
	assign v_1304 = (~v_97 & v_1302);
	assign v_1366 = (~v_97 & v_1365);
	assign v_1203 = (v_1202 ^ v_142);
	assign v_1330 = (v_1329 | ~v_94);
	assign v_1419 = (v_1417 | v_1418);
	assign v_1188 = (v_1187 ^ v_140);
	assign v_2199 = (((((((~v_1473 & ~v_1474)) & ~v_1586)) & ~v_1593)) & ~v_1600);
	assign v_1551 = (((v_1549 | v_1550)) | ~v_177);
	assign v_1616 = v_161);
	assign v_1826 = (~v_196 & v_1815);
	assign v_1717 = (~v_196 & v_1706);
	assign v_1823 = (~v_196 & v_1812);
	assign v_1714 = (~v_196 & v_1703);
	assign v_1820 = (~v_196 & v_1809);
	assign v_1711 = (~v_196 & v_1700);
	assign v_1817 = (~v_196 & v_1806);
	assign v_1708 = (~v_196 & v_1697);
	assign v_1904 = (~v_199 & v_1902);
	assign v_1966 = (~v_199 & v_1965);
	assign v_1803 = (v_1802 ^ v_244);
	assign v_1930 = (v_1929 | ~v_196);
	assign v_2019 = (v_2017 | v_2018);
	assign v_1788 = (v_1787 ^ v_242);
	assign v_358 = (~v_20 & v_357);
	assign v_424 = (v_20 & v_422);
	assign v_423 = (v_422 ^ v_20);
	assign v_633 = (v_631 | v_632);
	assign v_524 = (v_522 | v_523);
	assign v_630 = (v_628 | v_629);
	assign v_521 = (v_519 | v_520);
	assign v_627 = (v_625 | v_626);
	assign v_518 = (v_516 | v_517);
	assign v_624 = (v_622 | v_623);
	assign v_515 = (v_513 | v_514);
	assign v_711 = (v_709 | v_710);
	assign v_773 = (~v_41 & v_772);
	assign v_737 = (~v_38 & v_736);
	assign v_827 = (v_38 & v_825);
	assign v_952 = (~v_75 & v_951);
	assign v_1018 = (v_75 & v_1016);
	assign v_1017 = (v_1016 ^ v_75);
	assign v_1227 = (v_1225 | v_1226);
	assign v_1118 = (v_1116 | v_1117);
	assign v_1224 = (v_1222 | v_1223);
	assign v_1115 = (v_1113 | v_1114);
	assign v_1221 = (v_1219 | v_1220);
	assign v_1112 = (v_1110 | v_1111);
	assign v_1218 = (v_1216 | v_1217);
	assign v_1109 = (v_1107 | v_1108);
	assign v_2173 = (((((((~v_578 & ~v_594)) & ~v_609)) & ~v_687)) & ~v_694);
	assign v_1305 = (v_1303 | v_1304);
	assign v_1367 = (~v_97 & v_1366);
	assign v_1331 = (~v_94 & v_1330);
	assign v_1421 = (v_94 & v_1419);
	assign v_2182 = (((((((~v_1172 & ~v_1188)) & ~v_1203)) & ~v_1281)) & ~v_1288);
	assign v_1552 = (~v_178 & v_1551);
	assign v_1618 = (v_178 & v_1616);
	assign v_1617 = (v_1616 ^ v_178);
	assign v_1827 = (v_1825 | v_1826);
	assign v_1718 = (v_1716 | v_1717);
	assign v_1824 = (v_1822 | v_1823);
	assign v_1715 = (v_1713 | v_1714);
	assign v_1821 = (v_1819 | v_1820);
	assign v_1712 = (v_1710 | v_1711);
	assign v_1818 = (v_1816 | v_1817);
	assign v_1709 = (v_1707 | v_1708);
	assign v_1905 = (v_1903 | v_1904);
	assign v_1967 = (~v_199 & v_1966);
	assign v_1931 = (~v_196 & v_1930);
	assign v_2021 = (v_196 & v_2019);
	assign v_2200 = (((((((~v_1772 & ~v_1788)) & ~v_1803)) & ~v_1881)) & ~v_1888);
	assign v_359 = (((v_357 | v_358)) | ~v_20);
	assign v_425 = v_42);
	assign v_644 = (v_38 & v_633);
	assign v_535 = (v_38 & v_524);
	assign v_641 = (v_38 & v_630);
	assign v_532 = (v_38 & v_521);
	assign v_638 = (v_38 & v_627);
	assign v_529 = (v_38 & v_518);
	assign v_635 = (v_38 & v_624);
	assign v_526 = (v_38 & v_515);
	assign v_713 = (v_41 & v_711);
	assign v_774 = (v_41 | v_773);
	assign v_738 = (v_38 & v_737);
	assign v_828 = (v_826 | v_827);
	assign v_953 = (((v_951 | v_952)) | ~v_75);
	assign v_1019 = v_101);
	assign v_1238 = (v_94 & v_1227);
	assign v_1129 = (v_94 & v_1118);
	assign v_1235 = (v_94 & v_1224);
	assign v_1126 = (v_94 & v_1115);
	assign v_1232 = (v_94 & v_1221);
	assign v_1123 = (v_94 & v_1112);
	assign v_1229 = (v_94 & v_1218);
	assign v_1120 = (v_94 & v_1109);
	assign v_1307 = (v_97 & v_1305);
	assign v_1368 = (v_97 | v_1367);
	assign v_1332 = (v_94 & v_1331);
	assign v_1422 = (v_1420 | v_1421);
	assign v_1553 = (((v_1551 | v_1552)) | ~v_178);
	assign v_1619 = v_161);
	assign v_1838 = (v_196 & v_1827);
	assign v_1729 = (v_196 & v_1718);
	assign v_1835 = (v_196 & v_1824);
	assign v_1726 = (v_196 & v_1715);
	assign v_1832 = (v_196 & v_1821);
	assign v_1723 = (v_196 & v_1712);
	assign v_1829 = (v_196 & v_1818);
	assign v_1720 = (v_196 & v_1709);
	assign v_1907 = (v_199 & v_1905);
	assign v_1968 = (v_199 | v_1967);
	assign v_1932 = (v_196 & v_1931);
	assign v_2022 = (v_2020 | v_2021);
	assign v_360 = (~v_21 & v_359);
	assign v_427 = (v_21 & v_425);
	assign v_426 = (v_425 ^ v_21);
	assign v_645 = (v_643 | v_644);
	assign v_536 = (v_534 | v_535);
	assign v_642 = (v_640 | v_641);
	assign v_533 = (v_531 | v_532);
	assign v_639 = (v_637 | v_638);
	assign v_530 = (v_528 | v_529);
	assign v_636 = (v_634 | v_635);
	assign v_527 = (v_525 | v_526);
	assign v_714 = (v_712 | v_713);
	assign v_739 = (v_738 | ~v_38);
	assign v_830 = (~v_38 & v_828);
	assign v_954 = (~v_76 & v_953);
	assign v_1021 = (v_76 & v_1019);
	assign v_1020 = (v_1019 ^ v_76);
	assign v_1239 = (v_1237 | v_1238);
	assign v_1130 = (v_1128 | v_1129);
	assign v_1236 = (v_1234 | v_1235);
	assign v_1127 = (v_1125 | v_1126);
	assign v_1233 = (v_1231 | v_1232);
	assign v_1124 = (v_1122 | v_1123);
	assign v_1230 = (v_1228 | v_1229);
	assign v_1121 = (v_1119 | v_1120);
	assign v_1308 = (v_1306 | v_1307);
	assign v_1333 = (v_1332 | ~v_94);
	assign v_1424 = (~v_94 & v_1422);
	assign v_1554 = (~v_179 & v_1553);
	assign v_1621 = (v_179 & v_1619);
	assign v_1620 = (v_1619 ^ v_179);
	assign v_1839 = (v_1837 | v_1838);
	assign v_1730 = (v_1728 | v_1729);
	assign v_1836 = (v_1834 | v_1835);
	assign v_1727 = (v_1725 | v_1726);
	assign v_1833 = (v_1831 | v_1832);
	assign v_1724 = (v_1722 | v_1723);
	assign v_1830 = (v_1828 | v_1829);
	assign v_1721 = (v_1719 | v_1720);
	assign v_1908 = (v_1906 | v_1907);
	assign v_1933 = (v_1932 | ~v_196);
	assign v_2024 = (~v_196 & v_2022);
	assign v_361 = v_36);
	assign v_428 = v_42);
	assign v_656 = (~v_38 & v_645);
	assign v_547 = (~v_38 & v_536);
	assign v_653 = (~v_38 & v_642);
	assign v_544 = (~v_38 & v_533);
	assign v_650 = (~v_38 & v_639);
	assign v_541 = (~v_38 & v_530);
	assign v_647 = (~v_38 & v_636);
	assign v_538 = (~v_38 & v_527);
	assign v_716 = (~v_41 & v_714);
	assign v_740 = (v_739 ^ v_94);
	assign v_831 = (v_829 | v_830);
	assign v_955 = v_95);
	assign v_1022 = v_102);
	assign v_1250 = (~v_94 & v_1239);
	assign v_1141 = (~v_94 & v_1130);
	assign v_1247 = (~v_94 & v_1236);
	assign v_1138 = (~v_94 & v_1127);
	assign v_1244 = (~v_94 & v_1233);
	assign v_1135 = (~v_94 & v_1124);
	assign v_1241 = (~v_94 & v_1230);
	assign v_1132 = (~v_94 & v_1121);
	assign v_1310 = (~v_97 & v_1308);
	assign v_1334 = (v_1333 ^ v_150);
	assign v_1425 = (v_1423 | v_1424);
	assign v_1555 = v_155);
	assign v_1622 = v_162);
	assign v_1850 = (~v_196 & v_1839);
	assign v_1741 = (~v_196 & v_1730);
	assign v_1847 = (~v_196 & v_1836);
	assign v_1738 = (~v_196 & v_1727);
	assign v_1844 = (~v_196 & v_1833);
	assign v_1735 = (~v_196 & v_1724);
	assign v_1841 = (~v_196 & v_1830);
	assign v_1732 = (~v_196 & v_1721);
	assign v_1910 = (~v_199 & v_1908);
	assign v_1934 = (v_1933 ^ v_252);
	assign v_2025 = (v_2023 | v_2024);
	assign v_362 = (~v_22 & v_361);
	assign v_430 = (v_22 & v_428);
	assign v_429 = (v_428 ^ v_22);
	assign v_657 = (v_655 | v_656);
	assign v_548 = (v_546 | v_547);
	assign v_654 = (v_652 | v_653);
	assign v_545 = (v_543 | v_544);
	assign v_651 = (v_649 | v_650);
	assign v_542 = (v_540 | v_541);
	assign v_648 = (v_646 | v_647);
	assign v_539 = (v_537 | v_538);
	assign v_717 = (v_715 | v_716);
	assign v_833 = (v_38 & v_831);
	assign v_956 = (~v_77 & v_955);
	assign v_1024 = (v_77 & v_1022);
	assign v_1023 = (v_1022 ^ v_77);
	assign v_1251 = (v_1249 | v_1250);
	assign v_1142 = (v_1140 | v_1141);
	assign v_1248 = (v_1246 | v_1247);
	assign v_1139 = (v_1137 | v_1138);
	assign v_1245 = (v_1243 | v_1244);
	assign v_1136 = (v_1134 | v_1135);
	assign v_1242 = (v_1240 | v_1241);
	assign v_1133 = (v_1131 | v_1132);
	assign v_1311 = (v_1309 | v_1310);
	assign v_1427 = (v_94 & v_1425);
	assign v_1556 = (~v_180 & v_1555);
	assign v_1624 = (v_180 & v_1622);
	assign v_1623 = (v_1622 ^ v_180);
	assign v_1851 = (v_1849 | v_1850);
	assign v_1742 = (v_1740 | v_1741);
	assign v_1848 = (v_1846 | v_1847);
	assign v_1739 = (v_1737 | v_1738);
	assign v_1845 = (v_1843 | v_1844);
	assign v_1736 = (v_1734 | v_1735);
	assign v_1842 = (v_1840 | v_1841);
	assign v_1733 = (v_1731 | v_1732);
	assign v_1911 = (v_1909 | v_1910);
	assign v_2027 = (v_196 & v_2025);
	assign v_363 = v_36);
	assign v_431 = v_43);
	assign v_668 = (v_38 & v_657);
	assign v_559 = (v_38 & v_548);
	assign v_665 = (v_38 & v_654);
	assign v_556 = (v_38 & v_545);
	assign v_662 = (v_38 & v_651);
	assign v_553 = (v_38 & v_542);
	assign v_659 = (v_38 & v_648);
	assign v_550 = (v_38 & v_539);
	assign v_718 = (~v_41 & v_717);
	assign v_834 = (v_832 | v_833);
	assign v_957 = v_95);
	assign v_1025 = v_102);
	assign v_1262 = (v_94 & v_1251);
	assign v_1153 = (v_94 & v_1142);
	assign v_1259 = (v_94 & v_1248);
	assign v_1150 = (v_94 & v_1139);
	assign v_1256 = (v_94 & v_1245);
	assign v_1147 = (v_94 & v_1136);
	assign v_1253 = (v_94 & v_1242);
	assign v_1144 = (v_94 & v_1133);
	assign v_1312 = (~v_97 & v_1311);
	assign v_1428 = (v_1426 | v_1427);
	assign v_1557 = v_155);
	assign v_1625 = v_162);
	assign v_1862 = (v_196 & v_1851);
	assign v_1753 = (v_196 & v_1742);
	assign v_1859 = (v_196 & v_1848);
	assign v_1750 = (v_196 & v_1739);
	assign v_1856 = (v_196 & v_1845);
	assign v_1747 = (v_196 & v_1736);
	assign v_1853 = (v_196 & v_1842);
	assign v_1744 = (v_196 & v_1733);
	assign v_1912 = (~v_199 & v_1911);
	assign v_2028 = (v_2026 | v_2027);
	assign v_364 = (~v_23 & v_363);
	assign v_432 = (v_431 ^ v_23);
	assign v_433 = (v_23 & v_431);
	assign v_669 = (v_667 | v_668);
	assign v_560 = (v_558 | v_559);
	assign v_666 = (v_664 | v_665);
	assign v_557 = (v_555 | v_556);
	assign v_663 = (v_661 | v_662);
	assign v_554 = (v_552 | v_553);
	assign v_660 = (v_658 | v_659);
	assign v_551 = (v_549 | v_550);
	assign v_835 = (v_834 ^ v_100);
	assign v_958 = (~v_78 & v_957);
	assign v_1026 = (v_1025 ^ v_78);
	assign v_1027 = (v_78 & v_1025);
	assign v_1263 = (v_1261 | v_1262);
	assign v_1154 = (v_1152 | v_1153);
	assign v_1260 = (v_1258 | v_1259);
	assign v_1151 = (v_1149 | v_1150);
	assign v_1257 = (v_1255 | v_1256);
	assign v_1148 = (v_1146 | v_1147);
	assign v_1254 = (v_1252 | v_1253);
	assign v_1145 = (v_1143 | v_1144);
	assign v_1429 = (v_1428 ^ v_156);
	assign v_1558 = (~v_181 & v_1557);
	assign v_1626 = (v_1625 ^ v_181);
	assign v_1627 = (v_181 & v_1625);
	assign v_1863 = (v_1861 | v_1862);
	assign v_1754 = (v_1752 | v_1753);
	assign v_1860 = (v_1858 | v_1859);
	assign v_1751 = (v_1749 | v_1750);
	assign v_1857 = (v_1855 | v_1856);
	assign v_1748 = (v_1746 | v_1747);
	assign v_1854 = (v_1852 | v_1853);
	assign v_1745 = (v_1743 | v_1744);
	assign v_2029 = (v_2028 ^ v_258);
	assign v_365 = v_36);
	assign v_434 = v_43);
	assign v_673 = (v_669 ^ v_90);
	assign v_564 = (v_560 ^ v_82);
	assign v_672 = (v_666 ^ v_89);
	assign v_563 = (v_557 ^ v_81);
	assign v_671 = (v_663 ^ v_88);
	assign v_562 = (v_554 ^ v_80);
	assign v_670 = (v_660 ^ v_87);
	assign v_561 = (v_551 ^ v_79);
	assign v_2175 = (((((((~v_794 & ~v_810)) & ~v_835)) & ~v_848)) & ~v_858);
	assign v_959 = v_95);
	assign v_1028 = v_102);
	assign v_1267 = (v_1263 ^ v_146);
	assign v_1158 = (v_1154 ^ v_138);
	assign v_1266 = (v_1260 ^ v_145);
	assign v_1157 = (v_1151 ^ v_137);
	assign v_1265 = (v_1257 ^ v_144);
	assign v_1156 = (v_1148 ^ v_136);
	assign v_1264 = (v_1254 ^ v_143);
	assign v_1155 = (v_1145 ^ v_135);
	assign v_2184 = (((((((~v_1388 & ~v_1404)) & ~v_1429)) & ~v_1442)) & ~v_1452);
	assign v_1559 = v_155);
	assign v_1628 = v_162);
	assign v_1867 = (v_1863 ^ v_248);
	assign v_1758 = (v_1754 ^ v_240);
	assign v_1866 = (v_1860 ^ v_247);
	assign v_1757 = (v_1751 ^ v_239);
	assign v_1865 = (v_1857 ^ v_246);
	assign v_1756 = (v_1748 ^ v_238);
	assign v_1864 = (v_1854 ^ v_245);
	assign v_1755 = (v_1745 ^ v_237);
	assign v_2202 = (((((((~v_1988 & ~v_2004)) & ~v_2029)) & ~v_2042)) & ~v_2052);
	assign v_366 = v_36);
	assign v_674 = (((((~v_670 & ~v_671)) & ~v_672)) & ~v_673);
	assign v_565 = (((((~v_561 & ~v_562)) & ~v_563)) & ~v_564);
	assign v_960 = v_95);
	assign v_1268 = (((((~v_1264 & ~v_1265)) & ~v_1266)) & ~v_1267);
	assign v_1159 = (((((~v_1155 & ~v_1156)) & ~v_1157)) & ~v_1158);
	assign v_1560 = v_155);
	assign v_1868 = (((((~v_1864 & ~v_1865)) & ~v_1866)) & ~v_1867);
	assign v_1759 = (((((~v_1755 & ~v_1756)) & ~v_1757)) & ~v_1758);
	assign v_367 = v_36);
	assign v_961 = v_96);
	assign v_1561 = v_156);
	assign v_368 = v_36);
	assign v_962 = v_96);
	assign v_1562 = v_156);
	assign v_369 = v_36);
	assign v_963 = v_96);
	assign v_1563 = v_156);
	assign v_370 = v_36);
	assign v_964 = v_96);
	assign v_1564 = v_156);
	assign v_371 = v_37);
	assign v_965 = v_96);
	assign v_1565 = v_156);
	assign v_372 = v_37);
	assign v_966 = v_96);
	assign v_1566 = v_156);
	assign v_373 = v_37);
	assign v_967 = v_96);
	assign v_1567 = v_156);
	assign v_374 = v_37);
	assign v_968 = v_96);
	assign v_1568 = v_156);
	assign v_375 = v_37);
	assign v_969 = v_96);
	assign v_1569 = v_156);
	assign v_376 = v_37);
	assign v_970 = v_96);
	assign v_1570 = v_156);
	assign v_377 = v_37);
	assign v_971 = v_97);
	assign v_1571 = v_157);
	assign v_378 = v_37);
	assign v_972 = v_97);
	assign v_1572 = v_157);
	assign v_379 = v_37);
	assign v_973 = v_97);
	assign v_1573 = v_157);
	assign v_380 = v_37);
	assign v_974 = v_97);
	assign v_1574 = v_157);
	assign v_381 = v_38);
	assign v_975 = v_97);
	assign v_1575 = v_157);
	assign v_382 = v_38);
	assign v_976 = v_97);
	assign v_1576 = v_157);
	assign v_383 = v_38);
	assign v_977 = v_97);
	assign v_1577 = v_157);
	assign v_384 = v_38);
	assign v_978 = v_97);
	assign v_1578 = v_157);
	assign v_385 = v_38);
	assign v_979 = v_97);
	assign v_1579 = v_157);
	assign v_386 = v_38);
	assign v_980 = v_97);
	assign v_1580 = v_157);
	assign v_387 = v_38);
	assign v_981 = v_98);
	assign v_1581 = v_158);
	assign v_444 = (v_387 & v_432);
	assign v_443 = (v_387 & v_429);
	assign v_442 = (v_387 & v_426);
	assign v_441 = (v_387 & v_423);
	assign v_440 = (v_387 & v_420);
	assign v_439 = (v_387 & v_417);
	assign v_438 = (v_387 & v_414);
	assign v_437 = (v_387 & v_411);
	assign v_436 = (v_387 & v_408);
	assign v_435 = (~v_14 & v_387);
	assign v_776 = (v_387 & v_41);
	assign v_775 = (~v_387 & v_774);
	assign v_719 = (~v_387 & v_718);
	assign x_1 = (v_387 | ~v_388);
	assign v_1038 = (v_981 & v_1026);
	assign v_1037 = (v_981 & v_1023);
	assign v_1036 = (v_981 & v_1020);
	assign v_1035 = (v_981 & v_1017);
	assign v_1034 = (v_981 & v_1014);
	assign v_1033 = (v_981 & v_1011);
	assign v_1032 = (v_981 & v_1008);
	assign v_1031 = (v_981 & v_1005);
	assign v_1030 = (v_981 & v_1002);
	assign v_1029 = (~v_69 & v_981);
	assign v_1370 = (v_981 & v_97);
	assign v_1369 = (~v_981 & v_1368);
	assign v_1313 = (~v_981 & v_1312);
	assign x_2 = (v_981 | ~v_982);
	assign v_1638 = (v_1581 & v_1626);
	assign v_1637 = (v_1581 & v_1623);
	assign v_1636 = (v_1581 & v_1620);
	assign v_1635 = (v_1581 & v_1617);
	assign v_1634 = (v_1581 & v_1614);
	assign v_1633 = (v_1581 & v_1611);
	assign v_1632 = (v_1581 & v_1608);
	assign v_1631 = (v_1581 & v_1605);
	assign v_1630 = (v_1581 & v_1602);
	assign v_1629 = (~v_172 & v_1581);
	assign v_1970 = (v_1581 & v_199);
	assign v_1969 = (~v_1581 & v_1968);
	assign v_1913 = (~v_1581 & v_1912);
	assign x_3 = (v_1581 | ~v_1582);
	assign v_472 = (v_1 & v_444);
	assign v_469 = (v_1 & v_443);
	assign v_466 = (v_1 & v_442);
	assign v_463 = (v_1 & v_441);
	assign v_460 = (v_1 & v_440);
	assign v_457 = (v_1 & v_439);
	assign v_454 = (v_1 & v_438);
	assign v_451 = (v_1 & v_437);
	assign v_448 = (v_1 & v_436);
	assign v_445 = (v_1 & v_435);
	assign v_777 = (v_775 | v_776);
	assign v_720 = (v_719 | v_387);
	assign v_1066 = (v_47 & v_1038);
	assign v_1063 = (v_47 & v_1037);
	assign v_1060 = (v_47 & v_1036);
	assign v_1057 = (v_47 & v_1035);
	assign v_1054 = (v_47 & v_1034);
	assign v_1051 = (v_47 & v_1033);
	assign v_1048 = (v_47 & v_1032);
	assign v_1045 = (v_47 & v_1031);
	assign v_1042 = (v_47 & v_1030);
	assign v_1039 = (v_47 & v_1029);
	assign v_1371 = (v_1369 | v_1370);
	assign v_1314 = (v_1313 | v_981);
	assign x_5 = (x_1 & x_2);
	assign v_1666 = (v_159 & v_1638);
	assign v_1663 = (v_159 & v_1637);
	assign v_1660 = (v_159 & v_1636);
	assign v_1657 = (v_159 & v_1635);
	assign v_1654 = (v_159 & v_1634);
	assign v_1651 = (v_159 & v_1633);
	assign v_1648 = (v_159 & v_1632);
	assign v_1645 = (v_159 & v_1631);
	assign v_1642 = (v_159 & v_1630);
	assign v_1639 = (v_159 & v_1629);
	assign v_1971 = (v_1969 | v_1970);
	assign v_1914 = (v_1913 | v_1581);
	assign v_474 = (v_472 | v_473);
	assign v_471 = (v_469 | v_470);
	assign v_468 = (v_466 | v_467);
	assign v_465 = (v_463 | v_464);
	assign v_462 = (v_460 | v_461);
	assign v_459 = (v_457 | v_458);
	assign v_456 = (v_454 | v_455);
	assign v_453 = (v_451 | v_452);
	assign v_450 = (v_448 | v_449);
	assign v_447 = (v_445 | v_446);
	assign v_778 = (v_1 & v_777);
	assign v_721 = (v_1 & v_720);
	assign v_1068 = (v_1066 | v_1067);
	assign v_1065 = (v_1063 | v_1064);
	assign v_1062 = (v_1060 | v_1061);
	assign v_1059 = (v_1057 | v_1058);
	assign v_1056 = (v_1054 | v_1055);
	assign v_1053 = (v_1051 | v_1052);
	assign v_1050 = (v_1048 | v_1049);
	assign v_1047 = (v_1045 | v_1046);
	assign v_1044 = (v_1042 | v_1043);
	assign v_1041 = (v_1039 | v_1040);
	assign v_1372 = (v_47 & v_1371);
	assign v_1315 = (v_47 & v_1314);
	assign v_1668 = (v_1666 | v_1667);
	assign v_1665 = (v_1663 | v_1664);
	assign v_1662 = (v_1660 | v_1661);
	assign v_1659 = (v_1657 | v_1658);
	assign v_1656 = (v_1654 | v_1655);
	assign v_1653 = (v_1651 | v_1652);
	assign v_1650 = (v_1648 | v_1649);
	assign v_1647 = (v_1645 | v_1646);
	assign v_1644 = (v_1642 | v_1643);
	assign v_1641 = (v_1639 | v_1640);
	assign v_1972 = (v_159 & v_1971);
	assign v_1915 = (v_159 & v_1914);
	assign v_484 = (v_474 ^ v_78);
	assign v_483 = (v_471 ^ v_77);
	assign v_482 = (v_468 ^ v_76);
	assign v_481 = (v_465 ^ v_75);
	assign v_480 = (v_462 ^ v_74);
	assign v_479 = (v_459 ^ v_73);
	assign v_478 = (v_456 ^ v_72);
	assign v_477 = (v_453 ^ v_71);
	assign v_476 = (v_450 ^ v_70);
	assign v_475 = (v_447 ^ v_69);
	assign v_780 = (v_778 | v_779);
	assign v_722 = (v_721 | ~v_1);
	assign v_1078 = (v_1068 ^ v_134);
	assign v_1077 = (v_1065 ^ v_133);
	assign v_1076 = (v_1062 ^ v_132);
	assign v_1075 = (v_1059 ^ v_131);
	assign v_1074 = (v_1056 ^ v_130);
	assign v_1073 = (v_1053 ^ v_129);
	assign v_1072 = (v_1050 ^ v_128);
	assign v_1071 = (v_1047 ^ v_127);
	assign v_1070 = (v_1044 ^ v_126);
	assign v_1069 = (v_1041 ^ v_125);
	assign v_1374 = (v_1372 | v_1373);
	assign v_1316 = (v_1315 | ~v_47);
	assign v_1678 = (v_1668 ^ v_236);
	assign v_1677 = (v_1665 ^ v_235);
	assign v_1676 = (v_1662 ^ v_234);
	assign v_1675 = (v_1659 ^ v_233);
	assign v_1674 = (v_1656 ^ v_232);
	assign v_1673 = (v_1653 ^ v_231);
	assign v_1672 = (v_1650 ^ v_230);
	assign v_1671 = (v_1647 ^ v_229);
	assign v_1670 = (v_1644 ^ v_228);
	assign v_1669 = (v_1641 ^ v_227);
	assign v_1974 = (v_1972 | v_1973);
	assign v_1916 = (v_1915 | ~v_159);
	assign v_2171 = (((((((~v_480 & ~v_481)) & ~v_482)) & ~v_483)) & ~v_484);
	assign v_2170 = (((((((~v_475 & ~v_476)) & ~v_477)) & ~v_478)) & ~v_479);
	assign v_781 = (v_780 ^ v_97);
	assign v_723 = (v_722 ^ v_93);
	assign v_2180 = (((((((~v_1074 & ~v_1075)) & ~v_1076)) & ~v_1077)) & ~v_1078);
	assign v_2179 = (((((((~v_1069 & ~v_1070)) & ~v_1071)) & ~v_1072)) & ~v_1073);
	assign v_1375 = (v_1374 ^ v_153);
	assign v_1317 = (v_1316 ^ v_149);
	assign v_2198 = (((((((~v_1674 & ~v_1675)) & ~v_1676)) & ~v_1677)) & ~v_1678);
	assign v_2197 = (((((((~v_1669 & ~v_1670)) & ~v_1671)) & ~v_1672)) & ~v_1673);
	assign v_1975 = (v_1974 ^ v_255);
	assign v_1917 = (v_1916 ^ v_251);
	assign v_485 = (v_2170 & v_2171);
	assign v_2174 = (((((((~v_723 & ~v_740)) & ~v_749)) & ~v_760)) & ~v_781);
	assign v_1079 = (v_2179 & v_2180);
	assign v_2183 = (((((((~v_1317 & ~v_1334)) & ~v_1343)) & ~v_1354)) & ~v_1375);
	assign v_1679 = (v_2197 & v_2198);
	assign v_2201 = (((((((~v_1917 & ~v_1934)) & ~v_1943)) & ~v_1954)) & ~v_1975);
	assign v_2176 = (((((v_337 & v_485)) & v_565)) & v_674);
	assign v_2185 = (((((v_931 & v_1079)) & v_1159)) & v_1268);
	assign v_2203 = (((((v_1531 & v_1679)) & v_1759)) & v_1868);
	assign v_859 = (((((((v_2172 & v_2173)) & v_2174)) & v_2175)) & v_2176);
	assign v_1453 = (((((((v_2181 & v_2182)) & v_2183)) & v_2184)) & v_2185);
	assign v_2053 = (((((((v_2199 & v_2200)) & v_2201)) & v_2202)) & v_2203);
	assign v_1454 = (((v_265 & v_859)) & v_1453);
	assign v_2054 = (v_1459 & v_2053);
	assign v_2158 = (v_2054 & v_2157);
	assign x_4 = (v_2158 | ~v_1454);
	assign x_6 = (x_3 & x_4);
	assign x_7 = (x_5 & x_6);
	assign o_1 = x_);
endmodule
