module formula(v_1,v_2,v_3,v_4,v_5,v_6,v_7,v_8,v_9,v_10,v_11,v_12,v_13,v_14,v_15,v_16,v_17,v_18,v_19,v_20,v_21,v_22,v_23,v_24,v_25,v_26,v_27,v_28,v_29,v_30,v_31,v_32,v_33,v_34,v_35,v_36,v_37,v_38,v_39,v_40,v_41,v_42,v_43,v_44,v_45,v_46,v_47,v_48,v_49,v_50,v_51,v_52,v_53,v_54,v_55,v_56,o_1);
	input v_1;
	input v_2;
	input v_3;
	input v_4;
	input v_5;
	input v_6;
	input v_7;
	input v_8;
	input v_9;
	input v_10;
	input v_11;
	input v_12;
	input v_13;
	input v_14;
	input v_15;
	input v_16;
	input v_17;
	input v_18;
	input v_19;
	input v_20;
	input v_21;
	input v_22;
	input v_23;
	input v_24;
	input v_25;
	input v_26;
	input v_27;
	input v_28;
	input v_29;
	input v_30;
	input v_31;
	input v_32;
	input v_33;
	input v_34;
	input v_35;
	input v_36;
	input v_37;
	input v_38;
	input v_39;
	input v_40;
	input v_41;
	input v_42;
	input v_43;
	input v_44;
	input v_45;
	input v_46;
	input v_47;
	input v_48;
	input v_49;
	input v_50;
	input v_51;
	input v_52;
	input v_53;
	input v_54;
	input v_55;
	input v_56;
	wire v_57;
	wire v_58;
	wire v_59;
	wire v_60;
	wire v_61;
	wire v_62;
	wire v_63;
	wire v_64;
	wire v_65;
	wire v_66;
	wire v_67;
	wire v_68;
	wire v_69;
	wire v_70;
	wire v_71;
	wire v_72;
	wire v_73;
	wire v_74;
	wire v_75;
	wire v_76;
	wire v_77;
	wire v_78;
	wire v_79;
	wire v_80;
	wire v_81;
	wire v_82;
	wire v_83;
	wire v_84;
	wire v_85;
	wire v_86;
	wire v_87;
	wire v_88;
	wire v_89;
	wire v_90;
	wire v_91;
	wire v_92;
	wire v_93;
	wire v_94;
	wire v_95;
	wire v_96;
	wire v_97;
	wire v_98;
	wire v_99;
	wire v_100;
	wire v_101;
	wire v_102;
	wire v_103;
	wire v_104;
	wire v_105;
	wire v_106;
	wire v_107;
	wire v_108;
	wire v_109;
	wire v_110;
	wire v_111;
	wire v_112;
	wire v_113;
	wire v_114;
	wire v_115;
	wire v_116;
	wire v_117;
	wire v_118;
	wire v_119;
	wire v_120;
	wire v_121;
	wire v_122;
	wire v_123;
	wire v_124;
	wire v_125;
	wire v_126;
	wire v_127;
	wire v_128;
	wire v_129;
	wire v_130;
	wire v_131;
	wire v_132;
	wire v_133;
	wire v_134;
	wire v_135;
	wire v_136;
	wire v_137;
	wire v_138;
	wire v_139;
	wire v_140;
	wire v_141;
	wire v_142;
	wire v_143;
	wire v_144;
	wire v_145;
	wire v_146;
	wire v_147;
	wire v_148;
	wire v_149;
	wire v_150;
	wire v_151;
	wire v_152;
	wire v_153;
	wire v_154;
	wire v_155;
	wire v_156;
	wire v_157;
	wire v_158;
	wire v_159;
	wire v_160;
	wire v_161;
	wire v_162;
	wire v_163;
	wire v_164;
	wire v_165;
	wire v_166;
	wire v_167;
	wire v_168;
	wire v_169;
	wire v_170;
	wire v_171;
	wire v_172;
	wire v_173;
	wire v_174;
	wire v_175;
	wire v_176;
	wire v_177;
	wire v_178;
	wire v_179;
	wire v_180;
	wire v_181;
	wire v_182;
	wire v_183;
	wire v_184;
	wire v_185;
	wire v_186;
	wire v_187;
	wire v_188;
	wire v_189;
	wire v_190;
	wire v_191;
	wire v_192;
	wire v_193;
	wire v_194;
	wire v_195;
	wire v_196;
	wire v_197;
	wire v_198;
	wire v_199;
	wire v_200;
	wire v_201;
	wire v_202;
	wire v_203;
	wire v_204;
	wire v_205;
	wire v_206;
	wire v_207;
	wire v_208;
	wire v_209;
	wire v_210;
	wire v_211;
	wire v_212;
	wire v_213;
	wire v_214;
	wire v_215;
	wire v_216;
	wire v_217;
	wire v_218;
	wire v_219;
	wire v_220;
	wire v_221;
	wire v_222;
	wire v_223;
	wire v_224;
	wire v_225;
	wire v_226;
	wire v_227;
	wire v_228;
	wire v_229;
	wire v_230;
	wire v_231;
	wire v_232;
	wire v_233;
	wire v_234;
	wire v_235;
	wire v_236;
	wire v_237;
	wire v_238;
	wire v_239;
	wire v_240;
	wire v_241;
	wire v_242;
	wire v_243;
	wire v_244;
	wire v_245;
	wire v_246;
	wire v_247;
	wire v_248;
	wire v_249;
	wire v_250;
	wire v_251;
	wire v_252;
	wire v_253;
	wire v_254;
	wire v_255;
	wire v_256;
	wire v_257;
	wire v_258;
	wire v_259;
	wire v_260;
	wire v_261;
	wire v_262;
	wire v_263;
	wire v_264;
	wire v_265;
	wire v_266;
	wire v_267;
	wire v_268;
	wire v_269;
	wire v_270;
	wire v_271;
	wire v_272;
	wire v_273;
	wire v_274;
	wire v_275;
	wire v_276;
	wire v_277;
	wire v_278;
	wire v_279;
	wire v_280;
	wire v_281;
	wire v_282;
	wire v_283;
	wire v_284;
	wire v_285;
	wire v_286;
	wire v_287;
	wire v_288;
	wire v_289;
	wire v_290;
	wire v_291;
	wire v_292;
	wire v_293;
	wire v_294;
	wire v_295;
	wire v_296;
	wire v_297;
	wire v_298;
	wire v_299;
	wire v_300;
	wire v_301;
	wire v_302;
	wire v_303;
	wire v_304;
	wire v_305;
	wire v_306;
	wire v_307;
	wire v_308;
	wire v_309;
	wire v_310;
	wire v_311;
	wire v_312;
	wire v_313;
	wire v_314;
	wire v_315;
	wire v_316;
	wire v_317;
	wire v_318;
	wire v_319;
	wire x_1;
	output o_1;
	assign v_261 = v_44 ;
	assign v_241 = v_41 ;
	assign v_217 = v_36 ;
	assign v_197 = v_33 ;
	assign v_169 = v_20 ;
	assign v_149 = v_17 ;
	assign v_125 = v_12 ;
	assign v_105 = v_9 ;
	assign v_81 = v_4 ;
	assign v_61 = v_1 ;
	assign v_263 = (v_45 & v_261) ;
	assign v_243 = (v_42 & v_241) ;
	assign v_219 = (v_37 & v_217) ;
	assign v_199 = (v_34 & v_197) ;
	assign v_171 = (v_21 & v_169) ;
	assign v_151 = (v_18 & v_149) ;
	assign v_127 = (v_13 & v_125) ;
	assign v_107 = (v_10 & v_105) ;
	assign v_83 = (v_5 & v_81) ;
	assign v_63 = (v_2 & v_61) ;
	assign v_264 = v_263 ;
	assign v_244 = v_243 ;
	assign v_220 = v_219 ;
	assign v_200 = v_199 ;
	assign v_172 = v_171 ;
	assign v_152 = v_151 ;
	assign v_128 = v_127 ;
	assign v_108 = v_107 ;
	assign v_84 = v_83 ;
	assign v_64 = v_63 ;
	assign v_265 = (v_264 ^ v_46) ;
	assign v_240 = (v_48 ^ v_47) ;
	assign v_262 = (v_261 ^ v_45) ;
	assign v_245 = (v_244 ^ v_43) ;
	assign v_242 = (v_241 ^ v_42) ;
	assign v_221 = (v_220 ^ v_38) ;
	assign v_196 = (v_40 ^ v_39) ;
	assign v_218 = (v_217 ^ v_37) ;
	assign v_201 = (v_200 ^ v_35) ;
	assign v_198 = (v_197 ^ v_34) ;
	assign v_173 = (v_172 ^ v_22) ;
	assign v_148 = (v_24 ^ v_23) ;
	assign v_170 = (v_169 ^ v_21) ;
	assign v_153 = (v_152 ^ v_19) ;
	assign v_150 = (v_149 ^ v_18) ;
	assign v_129 = (v_128 ^ v_14) ;
	assign v_104 = (v_16 ^ v_15) ;
	assign v_126 = (v_125 ^ v_13) ;
	assign v_109 = (v_108 ^ v_11) ;
	assign v_106 = (v_105 ^ v_10) ;
	assign v_85 = (v_84 ^ v_6) ;
	assign v_60 = (v_8 ^ v_7) ;
	assign v_82 = (v_81 ^ v_5) ;
	assign v_65 = (v_64 ^ v_3) ;
	assign v_62 = (v_61 ^ v_2) ;
	assign v_275 = (v_240 & v_265) ;
	assign v_274 = (~v_240 & v_46) ;
	assign v_272 = (v_240 & v_262) ;
	assign v_271 = (~v_240 & v_45) ;
	assign v_269 = (~v_44 & v_240) ;
	assign v_268 = (~v_240 & v_44) ;
	assign v_255 = (v_240 & v_43) ;
	assign v_254 = (~v_240 & v_245) ;
	assign v_252 = (v_240 & v_42) ;
	assign v_251 = (~v_240 & v_242) ;
	assign v_249 = (v_240 & v_41) ;
	assign v_248 = (~v_240 & ~v_41) ;
	assign v_231 = (v_196 & v_221) ;
	assign v_230 = (~v_196 & v_38) ;
	assign v_228 = (v_196 & v_218) ;
	assign v_227 = (~v_196 & v_37) ;
	assign v_225 = (~v_36 & v_196) ;
	assign v_224 = (~v_196 & v_36) ;
	assign v_211 = (v_196 & v_35) ;
	assign v_210 = (~v_196 & v_201) ;
	assign v_208 = (v_196 & v_34) ;
	assign v_207 = (~v_196 & v_198) ;
	assign v_205 = (v_196 & v_33) ;
	assign v_204 = (~v_196 & ~v_33) ;
	assign v_183 = (v_148 & v_173) ;
	assign v_182 = (~v_148 & v_22) ;
	assign v_180 = (v_148 & v_170) ;
	assign v_179 = (~v_148 & v_21) ;
	assign v_177 = (~v_20 & v_148) ;
	assign v_176 = (~v_148 & v_20) ;
	assign v_163 = (v_148 & v_19) ;
	assign v_162 = (~v_148 & v_153) ;
	assign v_160 = (v_148 & v_18) ;
	assign v_159 = (~v_148 & v_150) ;
	assign v_157 = (v_148 & v_17) ;
	assign v_156 = (~v_148 & ~v_17) ;
	assign v_139 = (v_104 & v_129) ;
	assign v_138 = (~v_104 & v_14) ;
	assign v_136 = (v_104 & v_126) ;
	assign v_135 = (~v_104 & v_13) ;
	assign v_133 = (~v_12 & v_104) ;
	assign v_132 = (~v_104 & v_12) ;
	assign v_119 = (v_104 & v_11) ;
	assign v_118 = (~v_104 & v_109) ;
	assign v_116 = (v_104 & v_10) ;
	assign v_115 = (~v_104 & v_106) ;
	assign v_113 = (v_104 & v_9) ;
	assign v_112 = (~v_104 & ~v_9) ;
	assign v_95 = (v_60 & v_85) ;
	assign v_94 = (~v_60 & v_6) ;
	assign v_92 = (v_60 & v_82) ;
	assign v_91 = (~v_60 & v_5) ;
	assign v_89 = (~v_4 & v_60) ;
	assign v_88 = (~v_60 & v_4) ;
	assign v_75 = (v_60 & v_3) ;
	assign v_74 = (~v_60 & v_65) ;
	assign v_72 = (v_60 & v_2) ;
	assign v_71 = (~v_60 & v_62) ;
	assign v_69 = (v_60 & v_1) ;
	assign v_68 = (~v_60 & ~v_1) ;
	assign v_276 = (v_274 | v_275) ;
	assign v_273 = (v_271 | v_272) ;
	assign v_270 = (v_268 | v_269) ;
	assign v_256 = (v_254 | v_255) ;
	assign v_253 = (v_251 | v_252) ;
	assign v_250 = (v_248 | v_249) ;
	assign v_232 = (v_230 | v_231) ;
	assign v_229 = (v_227 | v_228) ;
	assign v_226 = (v_224 | v_225) ;
	assign v_212 = (v_210 | v_211) ;
	assign v_209 = (v_207 | v_208) ;
	assign v_206 = (v_204 | v_205) ;
	assign v_184 = (v_182 | v_183) ;
	assign v_181 = (v_179 | v_180) ;
	assign v_178 = (v_176 | v_177) ;
	assign v_164 = (v_162 | v_163) ;
	assign v_161 = (v_159 | v_160) ;
	assign v_158 = (v_156 | v_157) ;
	assign v_140 = (v_138 | v_139) ;
	assign v_137 = (v_135 | v_136) ;
	assign v_134 = (v_132 | v_133) ;
	assign v_120 = (v_118 | v_119) ;
	assign v_117 = (v_115 | v_116) ;
	assign v_114 = (v_112 | v_113) ;
	assign v_96 = (v_94 | v_95) ;
	assign v_93 = (v_91 | v_92) ;
	assign v_90 = (v_88 | v_89) ;
	assign v_76 = (v_74 | v_75) ;
	assign v_73 = (v_71 | v_72) ;
	assign v_70 = (v_68 | v_69) ;
	assign v_313 = (v_54 ^ v_30) ;
	assign v_312 = (v_53 ^ v_29) ;
	assign v_311 = (v_52 ^ v_28) ;
	assign v_309 = (v_51 ^ v_27) ;
	assign v_308 = (v_50 ^ v_26) ;
	assign v_307 = (v_49 ^ v_25) ;
	assign v_302 = (v_46 ^ v_30) ;
	assign v_301 = (v_45 ^ v_29) ;
	assign v_300 = (v_44 ^ v_28) ;
	assign v_298 = (v_43 ^ v_27) ;
	assign v_297 = (v_42 ^ v_26) ;
	assign v_296 = (v_41 ^ v_25) ;
	assign v_291 = (v_38 ^ v_30) ;
	assign v_290 = (v_37 ^ v_29) ;
	assign v_289 = (v_36 ^ v_28) ;
	assign v_287 = (v_35 ^ v_27) ;
	assign v_286 = (v_34 ^ v_26) ;
	assign v_285 = (v_33 ^ v_25) ;
	assign v_279 = (v_276 ^ v_54) ;
	assign v_278 = (v_273 ^ v_53) ;
	assign v_277 = (v_270 ^ v_52) ;
	assign v_259 = (v_256 ^ v_51) ;
	assign v_258 = (v_253 ^ v_50) ;
	assign v_257 = (v_250 ^ v_49) ;
	assign v_235 = (v_232 ^ v_46) ;
	assign v_234 = (v_229 ^ v_45) ;
	assign v_233 = (v_226 ^ v_44) ;
	assign v_215 = (v_212 ^ v_43) ;
	assign v_214 = (v_209 ^ v_42) ;
	assign v_213 = (v_206 ^ v_41) ;
	assign v_187 = (v_184 ^ v_30) ;
	assign v_186 = (v_181 ^ v_29) ;
	assign v_185 = (v_178 ^ v_28) ;
	assign v_167 = (v_164 ^ v_27) ;
	assign v_166 = (v_161 ^ v_26) ;
	assign v_165 = (v_158 ^ v_25) ;
	assign v_143 = (v_140 ^ v_22) ;
	assign v_142 = (v_137 ^ v_21) ;
	assign v_141 = (v_134 ^ v_20) ;
	assign v_123 = (v_120 ^ v_19) ;
	assign v_122 = (v_117 ^ v_18) ;
	assign v_121 = (v_114 ^ v_17) ;
	assign v_99 = (v_96 ^ v_14) ;
	assign v_98 = (v_93 ^ v_13) ;
	assign v_97 = (v_90 ^ v_12) ;
	assign v_79 = (v_76 ^ v_11) ;
	assign v_78 = (v_73 ^ v_10) ;
	assign v_77 = (v_70 ^ v_9) ;
	assign v_314 = ((~v_311 & ~v_312) & ~v_313) ;
	assign v_310 = ((~v_307 & ~v_308) & ~v_309) ;
	assign v_316 = (v_56 ^ v_32) ;
	assign v_315 = (v_55 ^ v_31) ;
	assign v_303 = ((~v_300 & ~v_301) & ~v_302) ;
	assign v_299 = ((~v_296 & ~v_297) & ~v_298) ;
	assign v_305 = (v_48 ^ v_32) ;
	assign v_304 = (v_47 ^ v_31) ;
	assign v_292 = ((~v_289 & ~v_290) & ~v_291) ;
	assign v_288 = ((~v_285 & ~v_286) & ~v_287) ;
	assign v_294 = (v_40 ^ v_32) ;
	assign v_293 = (v_39 ^ v_31) ;
	assign v_280 = ((~v_277 & ~v_278) & ~v_279) ;
	assign v_260 = ((~v_257 & ~v_258) & ~v_259) ;
	assign v_282 = (v_47 ^ v_56) ;
	assign v_281 = (~v_55 ^ v_48) ;
	assign v_236 = ((~v_233 & ~v_234) & ~v_235) ;
	assign v_216 = ((~v_213 & ~v_214) & ~v_215) ;
	assign v_238 = (v_39 ^ v_48) ;
	assign v_237 = (~v_47 ^ v_40) ;
	assign v_194 = ((~v_36 & ~v_37) & ~v_38) ;
	assign v_193 = ((~v_33 & ~v_34) & ~v_35) ;
	assign v_188 = ((~v_185 & ~v_186) & ~v_187) ;
	assign v_168 = ((~v_165 & ~v_166) & ~v_167) ;
	assign v_190 = (v_23 ^ v_32) ;
	assign v_189 = (~v_31 ^ v_24) ;
	assign v_144 = ((~v_141 & ~v_142) & ~v_143) ;
	assign v_124 = ((~v_121 & ~v_122) & ~v_123) ;
	assign v_146 = (v_15 ^ v_24) ;
	assign v_145 = (~v_23 ^ v_16) ;
	assign v_100 = ((~v_97 & ~v_98) & ~v_99) ;
	assign v_80 = ((~v_77 & ~v_78) & ~v_79) ;
	assign v_102 = (v_7 ^ v_16) ;
	assign v_101 = (~v_15 ^ v_8) ;
	assign v_58 = ((~v_4 & ~v_5) & ~v_6) ;
	assign v_57 = ((~v_1 & ~v_2) & ~v_3) ;
	assign v_317 = (((~v_315 & ~v_316) & v_310) & v_314) ;
	assign v_306 = (((~v_304 & ~v_305) & v_299) & v_303) ;
	assign v_295 = (((~v_293 & ~v_294) & v_288) & v_292) ;
	assign v_283 = (((~v_281 & ~v_282) & v_260) & v_280) ;
	assign v_239 = (((~v_237 & ~v_238) & v_216) & v_236) ;
	assign v_195 = (((~v_39 & ~v_40) & v_193) & v_194) ;
	assign v_191 = (((~v_189 & ~v_190) & v_168) & v_188) ;
	assign v_147 = (((~v_145 & ~v_146) & v_124) & v_144) ;
	assign v_103 = (((~v_101 & ~v_102) & v_80) & v_100) ;
	assign v_59 = (((~v_7 & ~v_8) & v_57) & v_58) ;
	assign v_318 = ((v_295 | v_306) | v_317) ;
	assign v_284 = ((v_195 & v_239) & v_283) ;
	assign v_192 = (((v_59 & v_103) & v_147) & v_191) ;
	assign v_319 = (v_284 & v_318) ;
	assign v_266 = (v_46 & v_264) ;
	assign v_246 = (v_43 & v_244) ;
	assign v_222 = (v_38 & v_220) ;
	assign v_202 = (v_35 & v_200) ;
	assign v_174 = (v_22 & v_172) ;
	assign v_154 = (v_19 & v_152) ;
	assign v_130 = (v_14 & v_128) ;
	assign v_110 = (v_11 & v_108) ;
	assign v_86 = (v_6 & v_84) ;
	assign v_66 = (v_3 & v_64) ;
	assign x_1 = (v_319 | ~v_192) ;
	assign v_267 = v_266 ;
	assign v_247 = v_246 ;
	assign v_223 = v_222 ;
	assign v_203 = v_202 ;
	assign v_175 = v_174 ;
	assign v_155 = v_154 ;
	assign v_131 = v_130 ;
	assign v_111 = v_110 ;
	assign v_87 = v_86 ;
	assign v_67 = v_66 ;
	assign o_1 = x_1 ;
endmodule
