// skolem function for order file variables
// Generated using findDep.cpp 
module stmt23_66_76 (v_2, v_3, v_4, v_5, v_7, v_8, v_213, v_214, v_219, v_221, v_225, v_227, v_229, v_230, v_232, v_234, v_236, v_237, v_239, v_241, v_243, v_245, v_247, v_249, v_251, v_254, v_255, v_262, v_264, v_268, v_272, v_274, v_279, v_280, v_281, v_283, v_286, v_288, v_292, v_293, v_295, v_297, v_298, v_303, v_308, v_309, v_311, v_312, v_316, v_318, v_322, v_324, v_326, v_333, v_334, v_336, v_338, v_340, v_345, v_346, v_348, v_350, v_352, v_354, v_357, v_359, v_360, v_362, v_364, v_366, v_370, v_372, v_373, v_375, v_377, v_379, v_381, v_385, v_389, v_391, v_392, v_394, v_396, v_398, v_400, v_406, v_410, v_411, v_413, v_415, v_417, v_419, v_422, v_424, v_425, v_427, v_429, v_431, v_435, v_437, v_438, v_440, v_442, v_444, v_446, v_450, v_454, v_456, v_457, v_459, v_461, v_463, v_465, v_471, v_475, v_477, v_481, v_486, v_489, v_491, v_493, v_494, v_496, v_498, v_500, v_501, v_503, v_505, v_507, v_509, v_511, v_513, v_515, v_518, v_519, v_526, v_528, v_532, v_537, v_542, v_543, v_547, v_549, v_551, v_555, v_559, v_561, v_563, v_565, v_569, v_571, v_573, v_574, v_578, v_583, v_584, v_586, v_589, v_591, v_594, v_600, v_601, v_605, v_607, v_609, v_613, v_617, v_619, v_621, v_623, v_627, v_629, v_631, v_632, v_636, v_641, v_643, v_645, v_647, v_649, v_663, v_666, v_669, v_670, v_672, v_674, v_675, v_680, v_682, v_684, v_685, v_687, v_690, v_692, v_695, v_700, v_705, v_706, v_707, v_711, v_713, v_715, v_719, v_723, v_724, v_726, v_727, v_729, v_731, v_733, v_735, v_738, v_739, v_742, v_746, v_747, v_751, v_753, v_755, v_759, v_760, v_764, v_766, v_768, v_772, v_775, v_776, v_780, v_782, v_784, v_788, v_792, v_798, v_799, v_800, v_801, v_805, v_809, v_811, v_815, v_817, v_822, v_823, v_824, v_828, v_832, v_834, v_838, v_840, v_845, v_846, v_847, v_851, v_855, v_857, v_861, v_863, v_868, v_869, v_870, v_872, v_879, v_880, v_881, v_882, v_886, v_890, v_892, v_896, v_898, v_903, v_904, v_905, v_909, v_913, v_915, v_919, v_921, v_926, v_927, v_928, v_932, v_936, v_938, v_942, v_944, v_949, v_950, v_951, v_953, v_960, v_961, v_962, v_963, v_967, v_971, v_973, v_977, v_979, v_984, v_985, v_986, v_990, v_994, v_996, v_1000, v_1002, v_1007, v_1008, v_1009, v_1013, v_1017, v_1019, v_1023, v_1025, v_1030, v_1031, v_1032, v_1034, v_1041, v_1042, v_1043, v_1047, v_1168, v_1169, v_1398, v_1402, v_1498, v_1814, v_1834, v_1885, v_1903, v_2137, v_2157, v_2208, v_2226, v_2338, v_2463, v_2483, v_2534, v_2552, v_2664, v_2789, v_2809, v_2860, v_2878, v_3114, v_3134, v_3185, v_3203, v_3315, v_3440, v_3460, v_3511, v_3529, v_3641, v_3646, v_3741, v_3932, v_4057, v_4077, v_4128, v_4146, v_4258, v_4259, v_4260, v_4261, v_4263, v_4264, v_4469, v_4470, v_4475, v_4477, v_4481, v_4483, v_4485, v_4486, v_4488, v_4490, v_4492, v_4493, v_4495, v_4497, v_4499, v_4501, v_4503, v_4505, v_4507, v_4510, v_4511, v_4518, v_4520, v_4524, v_4528, v_4530, v_4535, v_4536, v_4537, v_4539, v_4542, v_4544, v_4548, v_4549, v_4551, v_4553, v_4554, v_4559, v_4564, v_4565, v_4567, v_4568, v_4572, v_4574, v_4578, v_4580, v_4582, v_4589, v_4590, v_4592, v_4594, v_4596, v_4601, v_4602, v_4604, v_4606, v_4608, v_4610, v_4613, v_4615, v_4616, v_4618, v_4620, v_4622, v_4626, v_4628, v_4629, v_4631, v_4633, v_4635, v_4637, v_4641, v_4645, v_4647, v_4648, v_4650, v_4652, v_4654, v_4656, v_4662, v_4666, v_4667, v_4669, v_4671, v_4673, v_4675, v_4678, v_4680, v_4681, v_4683, v_4685, v_4687, v_4691, v_4693, v_4694, v_4696, v_4698, v_4700, v_4702, v_4706, v_4710, v_4712, v_4713, v_4715, v_4717, v_4719, v_4721, v_4727, v_4731, v_4733, v_4737, v_4742, v_4745, v_4747, v_4749, v_4750, v_4752, v_4754, v_4756, v_4757, v_4759, v_4761, v_4763, v_4765, v_4767, v_4769, v_4771, v_4774, v_4775, v_4782, v_4784, v_4788, v_4793, v_4798, v_4799, v_4803, v_4805, v_4807, v_4811, v_4815, v_4817, v_4819, v_4821, v_4825, v_4827, v_4829, v_4830, v_4834, v_4839, v_4840, v_4842, v_4845, v_4847, v_4850, v_4856, v_4857, v_4861, v_4863, v_4865, v_4869, v_4873, v_4875, v_4877, v_4879, v_4883, v_4885, v_4887, v_4888, v_4892, v_4897, v_4899, v_4901, v_4903, v_4905, v_4919, v_4922, v_4925, v_4926, v_4928, v_4930, v_4931, v_4936, v_4938, v_4940, v_4941, v_4943, v_4946, v_4948, v_4951, v_4956, v_4961, v_4962, v_4963, v_4967, v_4969, v_4971, v_4975, v_4979, v_4980, v_4982, v_4983, v_4985, v_4987, v_4989, v_4991, v_4994, v_4995, v_4998, v_5002, v_5003, v_5007, v_5009, v_5011, v_5015, v_5016, v_5020, v_5022, v_5024, v_5028, v_5031, v_5032, v_5036, v_5038, v_5040, v_5044, v_5048, v_5054, v_5055, v_5056, v_5060, v_5181, v_5182, v_5294, v_5298, v_5394, v_5605, v_5625, v_5676, v_5694, v_5823, v_5843, v_5894, v_5912, v_5919, v_6044, v_6064, v_6115, v_6133, v_6140, v_6265, v_6285, v_6336, v_6354, v_6485, v_6505, v_6556, v_6574, v_6581, v_6706, v_6726, v_6777, v_6795, v_6802, v_6807, v_6902, v_6988, v_7113, v_7133, v_7184, v_7202, o_1);
input v_2;
input v_3;
input v_4;
input v_5;
input v_7;
input v_8;
input v_213;
input v_214;
input v_219;
input v_221;
input v_225;
input v_227;
input v_229;
input v_230;
input v_232;
input v_234;
input v_236;
input v_237;
input v_239;
input v_241;
input v_243;
input v_245;
input v_247;
input v_249;
input v_251;
input v_254;
input v_255;
input v_262;
input v_264;
input v_268;
input v_272;
input v_274;
input v_279;
input v_280;
input v_281;
input v_283;
input v_286;
input v_288;
input v_292;
input v_293;
input v_295;
input v_297;
input v_298;
input v_303;
input v_308;
input v_309;
input v_311;
input v_312;
input v_316;
input v_318;
input v_322;
input v_324;
input v_326;
input v_333;
input v_334;
input v_336;
input v_338;
input v_340;
input v_345;
input v_346;
input v_348;
input v_350;
input v_352;
input v_354;
input v_357;
input v_359;
input v_360;
input v_362;
input v_364;
input v_366;
input v_370;
input v_372;
input v_373;
input v_375;
input v_377;
input v_379;
input v_381;
input v_385;
input v_389;
input v_391;
input v_392;
input v_394;
input v_396;
input v_398;
input v_400;
input v_406;
input v_410;
input v_411;
input v_413;
input v_415;
input v_417;
input v_419;
input v_422;
input v_424;
input v_425;
input v_427;
input v_429;
input v_431;
input v_435;
input v_437;
input v_438;
input v_440;
input v_442;
input v_444;
input v_446;
input v_450;
input v_454;
input v_456;
input v_457;
input v_459;
input v_461;
input v_463;
input v_465;
input v_471;
input v_475;
input v_477;
input v_481;
input v_486;
input v_489;
input v_491;
input v_493;
input v_494;
input v_496;
input v_498;
input v_500;
input v_501;
input v_503;
input v_505;
input v_507;
input v_509;
input v_511;
input v_513;
input v_515;
input v_518;
input v_519;
input v_526;
input v_528;
input v_532;
input v_537;
input v_542;
input v_543;
input v_547;
input v_549;
input v_551;
input v_555;
input v_559;
input v_561;
input v_563;
input v_565;
input v_569;
input v_571;
input v_573;
input v_574;
input v_578;
input v_583;
input v_584;
input v_586;
input v_589;
input v_591;
input v_594;
input v_600;
input v_601;
input v_605;
input v_607;
input v_609;
input v_613;
input v_617;
input v_619;
input v_621;
input v_623;
input v_627;
input v_629;
input v_631;
input v_632;
input v_636;
input v_641;
input v_643;
input v_645;
input v_647;
input v_649;
input v_663;
input v_666;
input v_669;
input v_670;
input v_672;
input v_674;
input v_675;
input v_680;
input v_682;
input v_684;
input v_685;
input v_687;
input v_690;
input v_692;
input v_695;
input v_700;
input v_705;
input v_706;
input v_707;
input v_711;
input v_713;
input v_715;
input v_719;
input v_723;
input v_724;
input v_726;
input v_727;
input v_729;
input v_731;
input v_733;
input v_735;
input v_738;
input v_739;
input v_742;
input v_746;
input v_747;
input v_751;
input v_753;
input v_755;
input v_759;
input v_760;
input v_764;
input v_766;
input v_768;
input v_772;
input v_775;
input v_776;
input v_780;
input v_782;
input v_784;
input v_788;
input v_792;
input v_798;
input v_799;
input v_800;
input v_801;
input v_805;
input v_809;
input v_811;
input v_815;
input v_817;
input v_822;
input v_823;
input v_824;
input v_828;
input v_832;
input v_834;
input v_838;
input v_840;
input v_845;
input v_846;
input v_847;
input v_851;
input v_855;
input v_857;
input v_861;
input v_863;
input v_868;
input v_869;
input v_870;
input v_872;
input v_879;
input v_880;
input v_881;
input v_882;
input v_886;
input v_890;
input v_892;
input v_896;
input v_898;
input v_903;
input v_904;
input v_905;
input v_909;
input v_913;
input v_915;
input v_919;
input v_921;
input v_926;
input v_927;
input v_928;
input v_932;
input v_936;
input v_938;
input v_942;
input v_944;
input v_949;
input v_950;
input v_951;
input v_953;
input v_960;
input v_961;
input v_962;
input v_963;
input v_967;
input v_971;
input v_973;
input v_977;
input v_979;
input v_984;
input v_985;
input v_986;
input v_990;
input v_994;
input v_996;
input v_1000;
input v_1002;
input v_1007;
input v_1008;
input v_1009;
input v_1013;
input v_1017;
input v_1019;
input v_1023;
input v_1025;
input v_1030;
input v_1031;
input v_1032;
input v_1034;
input v_1041;
input v_1042;
input v_1043;
input v_1047;
input v_1168;
input v_1169;
input v_1398;
input v_1402;
input v_1498;
input v_1814;
input v_1834;
input v_1885;
input v_1903;
input v_2137;
input v_2157;
input v_2208;
input v_2226;
input v_2338;
input v_2463;
input v_2483;
input v_2534;
input v_2552;
input v_2664;
input v_2789;
input v_2809;
input v_2860;
input v_2878;
input v_3114;
input v_3134;
input v_3185;
input v_3203;
input v_3315;
input v_3440;
input v_3460;
input v_3511;
input v_3529;
input v_3641;
input v_3646;
input v_3741;
input v_3932;
input v_4057;
input v_4077;
input v_4128;
input v_4146;
input v_4258;
input v_4259;
input v_4260;
input v_4261;
input v_4263;
input v_4264;
input v_4469;
input v_4470;
input v_4475;
input v_4477;
input v_4481;
input v_4483;
input v_4485;
input v_4486;
input v_4488;
input v_4490;
input v_4492;
input v_4493;
input v_4495;
input v_4497;
input v_4499;
input v_4501;
input v_4503;
input v_4505;
input v_4507;
input v_4510;
input v_4511;
input v_4518;
input v_4520;
input v_4524;
input v_4528;
input v_4530;
input v_4535;
input v_4536;
input v_4537;
input v_4539;
input v_4542;
input v_4544;
input v_4548;
input v_4549;
input v_4551;
input v_4553;
input v_4554;
input v_4559;
input v_4564;
input v_4565;
input v_4567;
input v_4568;
input v_4572;
input v_4574;
input v_4578;
input v_4580;
input v_4582;
input v_4589;
input v_4590;
input v_4592;
input v_4594;
input v_4596;
input v_4601;
input v_4602;
input v_4604;
input v_4606;
input v_4608;
input v_4610;
input v_4613;
input v_4615;
input v_4616;
input v_4618;
input v_4620;
input v_4622;
input v_4626;
input v_4628;
input v_4629;
input v_4631;
input v_4633;
input v_4635;
input v_4637;
input v_4641;
input v_4645;
input v_4647;
input v_4648;
input v_4650;
input v_4652;
input v_4654;
input v_4656;
input v_4662;
input v_4666;
input v_4667;
input v_4669;
input v_4671;
input v_4673;
input v_4675;
input v_4678;
input v_4680;
input v_4681;
input v_4683;
input v_4685;
input v_4687;
input v_4691;
input v_4693;
input v_4694;
input v_4696;
input v_4698;
input v_4700;
input v_4702;
input v_4706;
input v_4710;
input v_4712;
input v_4713;
input v_4715;
input v_4717;
input v_4719;
input v_4721;
input v_4727;
input v_4731;
input v_4733;
input v_4737;
input v_4742;
input v_4745;
input v_4747;
input v_4749;
input v_4750;
input v_4752;
input v_4754;
input v_4756;
input v_4757;
input v_4759;
input v_4761;
input v_4763;
input v_4765;
input v_4767;
input v_4769;
input v_4771;
input v_4774;
input v_4775;
input v_4782;
input v_4784;
input v_4788;
input v_4793;
input v_4798;
input v_4799;
input v_4803;
input v_4805;
input v_4807;
input v_4811;
input v_4815;
input v_4817;
input v_4819;
input v_4821;
input v_4825;
input v_4827;
input v_4829;
input v_4830;
input v_4834;
input v_4839;
input v_4840;
input v_4842;
input v_4845;
input v_4847;
input v_4850;
input v_4856;
input v_4857;
input v_4861;
input v_4863;
input v_4865;
input v_4869;
input v_4873;
input v_4875;
input v_4877;
input v_4879;
input v_4883;
input v_4885;
input v_4887;
input v_4888;
input v_4892;
input v_4897;
input v_4899;
input v_4901;
input v_4903;
input v_4905;
input v_4919;
input v_4922;
input v_4925;
input v_4926;
input v_4928;
input v_4930;
input v_4931;
input v_4936;
input v_4938;
input v_4940;
input v_4941;
input v_4943;
input v_4946;
input v_4948;
input v_4951;
input v_4956;
input v_4961;
input v_4962;
input v_4963;
input v_4967;
input v_4969;
input v_4971;
input v_4975;
input v_4979;
input v_4980;
input v_4982;
input v_4983;
input v_4985;
input v_4987;
input v_4989;
input v_4991;
input v_4994;
input v_4995;
input v_4998;
input v_5002;
input v_5003;
input v_5007;
input v_5009;
input v_5011;
input v_5015;
input v_5016;
input v_5020;
input v_5022;
input v_5024;
input v_5028;
input v_5031;
input v_5032;
input v_5036;
input v_5038;
input v_5040;
input v_5044;
input v_5048;
input v_5054;
input v_5055;
input v_5056;
input v_5060;
input v_5181;
input v_5182;
input v_5294;
input v_5298;
input v_5394;
input v_5605;
input v_5625;
input v_5676;
input v_5694;
input v_5823;
input v_5843;
input v_5894;
input v_5912;
input v_5919;
input v_6044;
input v_6064;
input v_6115;
input v_6133;
input v_6140;
input v_6265;
input v_6285;
input v_6336;
input v_6354;
input v_6485;
input v_6505;
input v_6556;
input v_6574;
input v_6581;
input v_6706;
input v_6726;
input v_6777;
input v_6795;
input v_6802;
input v_6807;
input v_6902;
input v_6988;
input v_7113;
input v_7133;
input v_7184;
input v_7202;
output o_1;
wire v_1;
wire v_6;
wire v_9;
wire v_10;
wire v_11;
wire v_12;
wire v_13;
wire v_14;
wire v_15;
wire v_16;
wire v_17;
wire v_18;
wire v_19;
wire v_20;
wire v_21;
wire v_22;
wire v_23;
wire v_24;
wire v_25;
wire v_26;
wire v_27;
wire v_28;
wire v_29;
wire v_30;
wire v_31;
wire v_32;
wire v_33;
wire v_34;
wire v_35;
wire v_36;
wire v_37;
wire v_38;
wire v_39;
wire v_40;
wire v_41;
wire v_42;
wire v_43;
wire v_44;
wire v_45;
wire v_46;
wire v_47;
wire v_48;
wire v_49;
wire v_50;
wire v_51;
wire v_52;
wire v_53;
wire v_54;
wire v_55;
wire v_56;
wire v_57;
wire v_58;
wire v_59;
wire v_60;
wire v_61;
wire v_62;
wire v_63;
wire v_64;
wire v_65;
wire v_66;
wire v_67;
wire v_68;
wire v_69;
wire v_70;
wire v_71;
wire v_72;
wire v_73;
wire v_74;
wire v_75;
wire v_76;
wire v_77;
wire v_78;
wire v_79;
wire v_80;
wire v_81;
wire v_82;
wire v_83;
wire v_84;
wire v_85;
wire v_86;
wire v_87;
wire v_88;
wire v_89;
wire v_90;
wire v_91;
wire v_92;
wire v_93;
wire v_94;
wire v_95;
wire v_96;
wire v_97;
wire v_98;
wire v_99;
wire v_100;
wire v_101;
wire v_102;
wire v_103;
wire v_104;
wire v_105;
wire v_106;
wire v_107;
wire v_108;
wire v_109;
wire v_110;
wire v_111;
wire v_112;
wire v_113;
wire v_114;
wire v_115;
wire v_116;
wire v_117;
wire v_118;
wire v_119;
wire v_120;
wire v_121;
wire v_122;
wire v_123;
wire v_124;
wire v_125;
wire v_126;
wire v_127;
wire v_128;
wire v_129;
wire v_130;
wire v_131;
wire v_132;
wire v_133;
wire v_134;
wire v_135;
wire v_136;
wire v_137;
wire v_138;
wire v_139;
wire v_140;
wire v_141;
wire v_142;
wire v_143;
wire v_144;
wire v_145;
wire v_146;
wire v_147;
wire v_148;
wire v_149;
wire v_150;
wire v_151;
wire v_152;
wire v_153;
wire v_154;
wire v_155;
wire v_156;
wire v_157;
wire v_158;
wire v_159;
wire v_160;
wire v_161;
wire v_162;
wire v_163;
wire v_164;
wire v_165;
wire v_166;
wire v_167;
wire v_168;
wire v_169;
wire v_170;
wire v_171;
wire v_172;
wire v_173;
wire v_174;
wire v_175;
wire v_176;
wire v_177;
wire v_178;
wire v_179;
wire v_180;
wire v_181;
wire v_182;
wire v_183;
wire v_184;
wire v_185;
wire v_186;
wire v_187;
wire v_188;
wire v_189;
wire v_190;
wire v_191;
wire v_192;
wire v_193;
wire v_194;
wire v_195;
wire v_196;
wire v_197;
wire v_198;
wire v_199;
wire v_200;
wire v_201;
wire v_202;
wire v_203;
wire v_204;
wire v_205;
wire v_206;
wire v_207;
wire v_208;
wire v_209;
wire v_210;
wire v_211;
wire v_212;
wire v_215;
wire v_216;
wire v_217;
wire v_218;
wire v_220;
wire v_222;
wire v_223;
wire v_224;
wire v_226;
wire v_228;
wire v_231;
wire v_233;
wire v_235;
wire v_238;
wire v_240;
wire v_242;
wire v_244;
wire v_246;
wire v_248;
wire v_250;
wire v_252;
wire v_253;
wire v_256;
wire v_257;
wire v_258;
wire v_259;
wire v_260;
wire v_261;
wire v_263;
wire v_265;
wire v_266;
wire v_267;
wire v_269;
wire v_270;
wire v_271;
wire v_273;
wire v_275;
wire v_276;
wire v_277;
wire v_278;
wire v_282;
wire v_284;
wire v_285;
wire v_287;
wire v_289;
wire v_290;
wire v_291;
wire v_294;
wire v_296;
wire v_299;
wire v_300;
wire v_301;
wire v_302;
wire v_304;
wire v_305;
wire v_306;
wire v_307;
wire v_310;
wire v_313;
wire v_314;
wire v_315;
wire v_317;
wire v_319;
wire v_320;
wire v_321;
wire v_323;
wire v_325;
wire v_327;
wire v_328;
wire v_329;
wire v_330;
wire v_331;
wire v_332;
wire v_335;
wire v_337;
wire v_339;
wire v_341;
wire v_342;
wire v_343;
wire v_344;
wire v_347;
wire v_349;
wire v_351;
wire v_353;
wire v_355;
wire v_356;
wire v_358;
wire v_361;
wire v_363;
wire v_365;
wire v_367;
wire v_368;
wire v_369;
wire v_371;
wire v_374;
wire v_376;
wire v_378;
wire v_380;
wire v_382;
wire v_383;
wire v_384;
wire v_386;
wire v_387;
wire v_388;
wire v_390;
wire v_393;
wire v_395;
wire v_397;
wire v_399;
wire v_401;
wire v_402;
wire v_403;
wire v_404;
wire v_405;
wire v_407;
wire v_408;
wire v_409;
wire v_412;
wire v_414;
wire v_416;
wire v_418;
wire v_420;
wire v_421;
wire v_423;
wire v_426;
wire v_428;
wire v_430;
wire v_432;
wire v_433;
wire v_434;
wire v_436;
wire v_439;
wire v_441;
wire v_443;
wire v_445;
wire v_447;
wire v_448;
wire v_449;
wire v_451;
wire v_452;
wire v_453;
wire v_455;
wire v_458;
wire v_460;
wire v_462;
wire v_464;
wire v_466;
wire v_467;
wire v_468;
wire v_469;
wire v_470;
wire v_472;
wire v_473;
wire v_474;
wire v_476;
wire v_478;
wire v_479;
wire v_480;
wire v_482;
wire v_483;
wire v_484;
wire v_485;
wire v_487;
wire v_488;
wire v_490;
wire v_492;
wire v_495;
wire v_497;
wire v_499;
wire v_502;
wire v_504;
wire v_506;
wire v_508;
wire v_510;
wire v_512;
wire v_514;
wire v_516;
wire v_517;
wire v_520;
wire v_521;
wire v_522;
wire v_523;
wire v_524;
wire v_525;
wire v_527;
wire v_529;
wire v_530;
wire v_531;
wire v_533;
wire v_534;
wire v_535;
wire v_536;
wire v_538;
wire v_539;
wire v_540;
wire v_541;
wire v_544;
wire v_545;
wire v_546;
wire v_548;
wire v_550;
wire v_552;
wire v_553;
wire v_554;
wire v_556;
wire v_557;
wire v_558;
wire v_560;
wire v_562;
wire v_564;
wire v_566;
wire v_567;
wire v_568;
wire v_570;
wire v_572;
wire v_575;
wire v_576;
wire v_577;
wire v_579;
wire v_580;
wire v_581;
wire v_582;
wire v_585;
wire v_587;
wire v_588;
wire v_590;
wire v_592;
wire v_593;
wire v_595;
wire v_596;
wire v_597;
wire v_598;
wire v_599;
wire v_602;
wire v_603;
wire v_604;
wire v_606;
wire v_608;
wire v_610;
wire v_611;
wire v_612;
wire v_614;
wire v_615;
wire v_616;
wire v_618;
wire v_620;
wire v_622;
wire v_624;
wire v_625;
wire v_626;
wire v_628;
wire v_630;
wire v_633;
wire v_634;
wire v_635;
wire v_637;
wire v_638;
wire v_639;
wire v_640;
wire v_642;
wire v_644;
wire v_646;
wire v_648;
wire v_650;
wire v_651;
wire v_652;
wire v_653;
wire v_654;
wire v_655;
wire v_656;
wire v_657;
wire v_658;
wire v_659;
wire v_660;
wire v_661;
wire v_662;
wire v_664;
wire v_665;
wire v_667;
wire v_668;
wire v_671;
wire v_673;
wire v_676;
wire v_677;
wire v_678;
wire v_679;
wire v_681;
wire v_683;
wire v_686;
wire v_688;
wire v_689;
wire v_691;
wire v_693;
wire v_694;
wire v_696;
wire v_697;
wire v_698;
wire v_699;
wire v_701;
wire v_702;
wire v_703;
wire v_704;
wire v_708;
wire v_709;
wire v_710;
wire v_712;
wire v_714;
wire v_716;
wire v_717;
wire v_718;
wire v_720;
wire v_721;
wire v_722;
wire v_725;
wire v_728;
wire v_730;
wire v_732;
wire v_734;
wire v_736;
wire v_737;
wire v_740;
wire v_741;
wire v_743;
wire v_744;
wire v_745;
wire v_748;
wire v_749;
wire v_750;
wire v_752;
wire v_754;
wire v_756;
wire v_757;
wire v_758;
wire v_761;
wire v_762;
wire v_763;
wire v_765;
wire v_767;
wire v_769;
wire v_770;
wire v_771;
wire v_773;
wire v_774;
wire v_777;
wire v_778;
wire v_779;
wire v_781;
wire v_783;
wire v_785;
wire v_786;
wire v_787;
wire v_789;
wire v_790;
wire v_791;
wire v_793;
wire v_794;
wire v_795;
wire v_796;
wire v_797;
wire v_802;
wire v_803;
wire v_804;
wire v_806;
wire v_807;
wire v_808;
wire v_810;
wire v_812;
wire v_813;
wire v_814;
wire v_816;
wire v_818;
wire v_819;
wire v_820;
wire v_821;
wire v_825;
wire v_826;
wire v_827;
wire v_829;
wire v_830;
wire v_831;
wire v_833;
wire v_835;
wire v_836;
wire v_837;
wire v_839;
wire v_841;
wire v_842;
wire v_843;
wire v_844;
wire v_848;
wire v_849;
wire v_850;
wire v_852;
wire v_853;
wire v_854;
wire v_856;
wire v_858;
wire v_859;
wire v_860;
wire v_862;
wire v_864;
wire v_865;
wire v_866;
wire v_867;
wire v_871;
wire v_873;
wire v_874;
wire v_875;
wire v_876;
wire v_877;
wire v_878;
wire v_883;
wire v_884;
wire v_885;
wire v_887;
wire v_888;
wire v_889;
wire v_891;
wire v_893;
wire v_894;
wire v_895;
wire v_897;
wire v_899;
wire v_900;
wire v_901;
wire v_902;
wire v_906;
wire v_907;
wire v_908;
wire v_910;
wire v_911;
wire v_912;
wire v_914;
wire v_916;
wire v_917;
wire v_918;
wire v_920;
wire v_922;
wire v_923;
wire v_924;
wire v_925;
wire v_929;
wire v_930;
wire v_931;
wire v_933;
wire v_934;
wire v_935;
wire v_937;
wire v_939;
wire v_940;
wire v_941;
wire v_943;
wire v_945;
wire v_946;
wire v_947;
wire v_948;
wire v_952;
wire v_954;
wire v_955;
wire v_956;
wire v_957;
wire v_958;
wire v_959;
wire v_964;
wire v_965;
wire v_966;
wire v_968;
wire v_969;
wire v_970;
wire v_972;
wire v_974;
wire v_975;
wire v_976;
wire v_978;
wire v_980;
wire v_981;
wire v_982;
wire v_983;
wire v_987;
wire v_988;
wire v_989;
wire v_991;
wire v_992;
wire v_993;
wire v_995;
wire v_997;
wire v_998;
wire v_999;
wire v_1001;
wire v_1003;
wire v_1004;
wire v_1005;
wire v_1006;
wire v_1010;
wire v_1011;
wire v_1012;
wire v_1014;
wire v_1015;
wire v_1016;
wire v_1018;
wire v_1020;
wire v_1021;
wire v_1022;
wire v_1024;
wire v_1026;
wire v_1027;
wire v_1028;
wire v_1029;
wire v_1033;
wire v_1035;
wire v_1036;
wire v_1037;
wire v_1038;
wire v_1039;
wire v_1040;
wire v_1044;
wire v_1045;
wire v_1046;
wire v_1048;
wire v_1049;
wire v_1050;
wire v_1051;
wire v_1052;
wire v_1053;
wire v_1054;
wire v_1055;
wire v_1056;
wire v_1057;
wire v_1058;
wire v_1059;
wire v_1060;
wire v_1061;
wire v_1062;
wire v_1063;
wire v_1064;
wire v_1065;
wire v_1066;
wire v_1067;
wire v_1068;
wire v_1069;
wire v_1070;
wire v_1071;
wire v_1072;
wire v_1073;
wire v_1074;
wire v_1075;
wire v_1076;
wire v_1077;
wire v_1078;
wire v_1079;
wire v_1080;
wire v_1081;
wire v_1082;
wire v_1083;
wire v_1084;
wire v_1085;
wire v_1086;
wire v_1087;
wire v_1088;
wire v_1089;
wire v_1090;
wire v_1091;
wire v_1092;
wire v_1093;
wire v_1094;
wire v_1095;
wire v_1096;
wire v_1097;
wire v_1098;
wire v_1099;
wire v_1100;
wire v_1101;
wire v_1102;
wire v_1103;
wire v_1104;
wire v_1105;
wire v_1106;
wire v_1107;
wire v_1108;
wire v_1109;
wire v_1110;
wire v_1111;
wire v_1112;
wire v_1113;
wire v_1114;
wire v_1115;
wire v_1116;
wire v_1117;
wire v_1118;
wire v_1119;
wire v_1120;
wire v_1121;
wire v_1122;
wire v_1123;
wire v_1124;
wire v_1125;
wire v_1126;
wire v_1127;
wire v_1128;
wire v_1129;
wire v_1130;
wire v_1131;
wire v_1132;
wire v_1133;
wire v_1134;
wire v_1135;
wire v_1136;
wire v_1137;
wire v_1138;
wire v_1139;
wire v_1140;
wire v_1141;
wire v_1142;
wire v_1143;
wire v_1144;
wire v_1145;
wire v_1146;
wire v_1147;
wire v_1148;
wire v_1149;
wire v_1150;
wire v_1151;
wire v_1152;
wire v_1153;
wire v_1154;
wire v_1155;
wire v_1156;
wire v_1157;
wire v_1158;
wire v_1159;
wire v_1160;
wire v_1161;
wire v_1162;
wire v_1163;
wire v_1164;
wire v_1165;
wire v_1166;
wire v_1167;
wire v_1170;
wire v_1171;
wire v_1172;
wire v_1173;
wire v_1174;
wire v_1175;
wire v_1176;
wire v_1177;
wire v_1178;
wire v_1179;
wire v_1180;
wire v_1181;
wire v_1182;
wire v_1183;
wire v_1184;
wire v_1185;
wire v_1186;
wire v_1187;
wire v_1188;
wire v_1189;
wire v_1190;
wire v_1191;
wire v_1192;
wire v_1193;
wire v_1194;
wire v_1195;
wire v_1196;
wire v_1197;
wire v_1198;
wire v_1199;
wire v_1200;
wire v_1201;
wire v_1202;
wire v_1203;
wire v_1204;
wire v_1205;
wire v_1206;
wire v_1207;
wire v_1208;
wire v_1209;
wire v_1210;
wire v_1211;
wire v_1212;
wire v_1213;
wire v_1214;
wire v_1215;
wire v_1216;
wire v_1217;
wire v_1218;
wire v_1219;
wire v_1220;
wire v_1221;
wire v_1222;
wire v_1223;
wire v_1224;
wire v_1225;
wire v_1226;
wire v_1227;
wire v_1228;
wire v_1229;
wire v_1230;
wire v_1231;
wire v_1232;
wire v_1233;
wire v_1234;
wire v_1235;
wire v_1236;
wire v_1237;
wire v_1238;
wire v_1239;
wire v_1240;
wire v_1241;
wire v_1242;
wire v_1243;
wire v_1244;
wire v_1245;
wire v_1246;
wire v_1247;
wire v_1248;
wire v_1249;
wire v_1250;
wire v_1251;
wire v_1252;
wire v_1253;
wire v_1254;
wire v_1255;
wire v_1256;
wire v_1257;
wire v_1258;
wire v_1259;
wire v_1260;
wire v_1261;
wire v_1262;
wire v_1263;
wire v_1264;
wire v_1265;
wire v_1266;
wire v_1267;
wire v_1268;
wire v_1269;
wire v_1270;
wire v_1271;
wire v_1272;
wire v_1273;
wire v_1274;
wire v_1275;
wire v_1276;
wire v_1277;
wire v_1278;
wire v_1279;
wire v_1280;
wire v_1281;
wire v_1282;
wire v_1283;
wire v_1284;
wire v_1285;
wire v_1286;
wire v_1287;
wire v_1288;
wire v_1289;
wire v_1290;
wire v_1291;
wire v_1292;
wire v_1293;
wire v_1294;
wire v_1295;
wire v_1296;
wire v_1297;
wire v_1298;
wire v_1299;
wire v_1300;
wire v_1301;
wire v_1302;
wire v_1303;
wire v_1304;
wire v_1305;
wire v_1306;
wire v_1307;
wire v_1308;
wire v_1309;
wire v_1310;
wire v_1311;
wire v_1312;
wire v_1313;
wire v_1314;
wire v_1315;
wire v_1316;
wire v_1317;
wire v_1318;
wire v_1319;
wire v_1320;
wire v_1321;
wire v_1322;
wire v_1323;
wire v_1324;
wire v_1325;
wire v_1326;
wire v_1327;
wire v_1328;
wire v_1329;
wire v_1330;
wire v_1331;
wire v_1332;
wire v_1333;
wire v_1334;
wire v_1335;
wire v_1336;
wire v_1337;
wire v_1338;
wire v_1339;
wire v_1340;
wire v_1341;
wire v_1342;
wire v_1343;
wire v_1344;
wire v_1345;
wire v_1346;
wire v_1347;
wire v_1348;
wire v_1349;
wire v_1350;
wire v_1351;
wire v_1352;
wire v_1353;
wire v_1354;
wire v_1355;
wire v_1356;
wire v_1357;
wire v_1358;
wire v_1359;
wire v_1360;
wire v_1361;
wire v_1362;
wire v_1363;
wire v_1364;
wire v_1365;
wire v_1366;
wire v_1367;
wire v_1368;
wire v_1369;
wire v_1370;
wire v_1371;
wire v_1372;
wire v_1373;
wire v_1374;
wire v_1375;
wire v_1376;
wire v_1377;
wire v_1378;
wire v_1379;
wire v_1380;
wire v_1381;
wire v_1382;
wire v_1383;
wire v_1384;
wire v_1385;
wire v_1386;
wire v_1387;
wire v_1388;
wire v_1389;
wire v_1390;
wire v_1391;
wire v_1392;
wire v_1393;
wire v_1394;
wire v_1395;
wire v_1396;
wire v_1397;
wire v_1399;
wire v_1400;
wire v_1401;
wire v_1403;
wire v_1404;
wire v_1405;
wire v_1406;
wire v_1407;
wire v_1408;
wire v_1409;
wire v_1410;
wire v_1411;
wire v_1412;
wire v_1413;
wire v_1414;
wire v_1415;
wire v_1416;
wire v_1417;
wire v_1418;
wire v_1419;
wire v_1420;
wire v_1421;
wire v_1422;
wire v_1423;
wire v_1424;
wire v_1425;
wire v_1426;
wire v_1427;
wire v_1428;
wire v_1429;
wire v_1430;
wire v_1431;
wire v_1432;
wire v_1433;
wire v_1434;
wire v_1435;
wire v_1436;
wire v_1437;
wire v_1438;
wire v_1439;
wire v_1440;
wire v_1441;
wire v_1442;
wire v_1443;
wire v_1444;
wire v_1445;
wire v_1446;
wire v_1447;
wire v_1448;
wire v_1449;
wire v_1450;
wire v_1451;
wire v_1452;
wire v_1453;
wire v_1454;
wire v_1455;
wire v_1456;
wire v_1457;
wire v_1458;
wire v_1459;
wire v_1460;
wire v_1461;
wire v_1462;
wire v_1463;
wire v_1464;
wire v_1465;
wire v_1466;
wire v_1467;
wire v_1468;
wire v_1469;
wire v_1470;
wire v_1471;
wire v_1472;
wire v_1473;
wire v_1474;
wire v_1475;
wire v_1476;
wire v_1477;
wire v_1478;
wire v_1479;
wire v_1480;
wire v_1481;
wire v_1482;
wire v_1483;
wire v_1484;
wire v_1485;
wire v_1486;
wire v_1487;
wire v_1488;
wire v_1489;
wire v_1490;
wire v_1491;
wire v_1492;
wire v_1493;
wire v_1494;
wire v_1495;
wire v_1496;
wire v_1497;
wire v_1499;
wire v_1500;
wire v_1501;
wire v_1502;
wire v_1503;
wire v_1504;
wire v_1505;
wire v_1506;
wire v_1507;
wire v_1508;
wire v_1509;
wire v_1510;
wire v_1511;
wire v_1512;
wire v_1513;
wire v_1514;
wire v_1515;
wire v_1516;
wire v_1517;
wire v_1518;
wire v_1519;
wire v_1520;
wire v_1521;
wire v_1522;
wire v_1523;
wire v_1524;
wire v_1525;
wire v_1526;
wire v_1527;
wire v_1528;
wire v_1529;
wire v_1530;
wire v_1531;
wire v_1532;
wire v_1533;
wire v_1534;
wire v_1535;
wire v_1536;
wire v_1537;
wire v_1538;
wire v_1539;
wire v_1540;
wire v_1541;
wire v_1542;
wire v_1543;
wire v_1544;
wire v_1545;
wire v_1546;
wire v_1547;
wire v_1548;
wire v_1549;
wire v_1550;
wire v_1551;
wire v_1552;
wire v_1553;
wire v_1554;
wire v_1555;
wire v_1556;
wire v_1557;
wire v_1558;
wire v_1559;
wire v_1560;
wire v_1561;
wire v_1562;
wire v_1563;
wire v_1564;
wire v_1565;
wire v_1566;
wire v_1567;
wire v_1568;
wire v_1569;
wire v_1570;
wire v_1571;
wire v_1572;
wire v_1573;
wire v_1574;
wire v_1575;
wire v_1576;
wire v_1577;
wire v_1578;
wire v_1579;
wire v_1580;
wire v_1581;
wire v_1582;
wire v_1583;
wire v_1584;
wire v_1585;
wire v_1586;
wire v_1587;
wire v_1588;
wire v_1589;
wire v_1590;
wire v_1591;
wire v_1592;
wire v_1593;
wire v_1594;
wire v_1595;
wire v_1596;
wire v_1597;
wire v_1598;
wire v_1599;
wire v_1600;
wire v_1601;
wire v_1602;
wire v_1603;
wire v_1604;
wire v_1605;
wire v_1606;
wire v_1607;
wire v_1608;
wire v_1609;
wire v_1610;
wire v_1611;
wire v_1612;
wire v_1613;
wire v_1614;
wire v_1615;
wire v_1616;
wire v_1617;
wire v_1618;
wire v_1619;
wire v_1620;
wire v_1621;
wire v_1622;
wire v_1623;
wire v_1624;
wire v_1625;
wire v_1626;
wire v_1627;
wire v_1628;
wire v_1629;
wire v_1630;
wire v_1631;
wire v_1632;
wire v_1633;
wire v_1634;
wire v_1635;
wire v_1636;
wire v_1637;
wire v_1638;
wire v_1639;
wire v_1640;
wire v_1641;
wire v_1642;
wire v_1643;
wire v_1644;
wire v_1645;
wire v_1646;
wire v_1647;
wire v_1648;
wire v_1649;
wire v_1650;
wire v_1651;
wire v_1652;
wire v_1653;
wire v_1654;
wire v_1655;
wire v_1656;
wire v_1657;
wire v_1658;
wire v_1659;
wire v_1660;
wire v_1661;
wire v_1662;
wire v_1663;
wire v_1664;
wire v_1665;
wire v_1666;
wire v_1667;
wire v_1668;
wire v_1669;
wire v_1670;
wire v_1671;
wire v_1672;
wire v_1673;
wire v_1674;
wire v_1675;
wire v_1676;
wire v_1677;
wire v_1678;
wire v_1679;
wire v_1680;
wire v_1681;
wire v_1682;
wire v_1683;
wire v_1684;
wire v_1685;
wire v_1686;
wire v_1687;
wire v_1688;
wire v_1689;
wire v_1690;
wire v_1691;
wire v_1692;
wire v_1693;
wire v_1694;
wire v_1695;
wire v_1696;
wire v_1697;
wire v_1698;
wire v_1699;
wire v_1700;
wire v_1701;
wire v_1702;
wire v_1703;
wire v_1704;
wire v_1705;
wire v_1706;
wire v_1707;
wire v_1708;
wire v_1709;
wire v_1710;
wire v_1711;
wire v_1712;
wire v_1713;
wire v_1714;
wire v_1715;
wire v_1716;
wire v_1717;
wire v_1718;
wire v_1719;
wire v_1720;
wire v_1721;
wire v_1722;
wire v_1723;
wire v_1724;
wire v_1725;
wire v_1726;
wire v_1727;
wire v_1728;
wire v_1729;
wire v_1730;
wire v_1731;
wire v_1732;
wire v_1733;
wire v_1734;
wire v_1735;
wire v_1736;
wire v_1737;
wire v_1738;
wire v_1739;
wire v_1740;
wire v_1741;
wire v_1742;
wire v_1743;
wire v_1744;
wire v_1745;
wire v_1746;
wire v_1747;
wire v_1748;
wire v_1749;
wire v_1750;
wire v_1751;
wire v_1752;
wire v_1753;
wire v_1754;
wire v_1755;
wire v_1756;
wire v_1757;
wire v_1758;
wire v_1759;
wire v_1760;
wire v_1761;
wire v_1762;
wire v_1763;
wire v_1764;
wire v_1765;
wire v_1766;
wire v_1767;
wire v_1768;
wire v_1769;
wire v_1770;
wire v_1771;
wire v_1772;
wire v_1773;
wire v_1774;
wire v_1775;
wire v_1776;
wire v_1777;
wire v_1778;
wire v_1779;
wire v_1780;
wire v_1781;
wire v_1782;
wire v_1783;
wire v_1784;
wire v_1785;
wire v_1786;
wire v_1787;
wire v_1788;
wire v_1789;
wire v_1790;
wire v_1791;
wire v_1792;
wire v_1793;
wire v_1794;
wire v_1795;
wire v_1796;
wire v_1797;
wire v_1798;
wire v_1799;
wire v_1800;
wire v_1801;
wire v_1802;
wire v_1803;
wire v_1804;
wire v_1805;
wire v_1806;
wire v_1807;
wire v_1808;
wire v_1809;
wire v_1810;
wire v_1811;
wire v_1812;
wire v_1813;
wire v_1815;
wire v_1816;
wire v_1817;
wire v_1818;
wire v_1819;
wire v_1820;
wire v_1821;
wire v_1822;
wire v_1823;
wire v_1824;
wire v_1825;
wire v_1826;
wire v_1827;
wire v_1828;
wire v_1829;
wire v_1830;
wire v_1831;
wire v_1832;
wire v_1833;
wire v_1835;
wire v_1836;
wire v_1837;
wire v_1838;
wire v_1839;
wire v_1840;
wire v_1841;
wire v_1842;
wire v_1843;
wire v_1844;
wire v_1845;
wire v_1846;
wire v_1847;
wire v_1848;
wire v_1849;
wire v_1850;
wire v_1851;
wire v_1852;
wire v_1853;
wire v_1854;
wire v_1855;
wire v_1856;
wire v_1857;
wire v_1858;
wire v_1859;
wire v_1860;
wire v_1861;
wire v_1862;
wire v_1863;
wire v_1864;
wire v_1865;
wire v_1866;
wire v_1867;
wire v_1868;
wire v_1869;
wire v_1870;
wire v_1871;
wire v_1872;
wire v_1873;
wire v_1874;
wire v_1875;
wire v_1876;
wire v_1877;
wire v_1878;
wire v_1879;
wire v_1880;
wire v_1881;
wire v_1882;
wire v_1883;
wire v_1884;
wire v_1886;
wire v_1887;
wire v_1888;
wire v_1889;
wire v_1890;
wire v_1891;
wire v_1892;
wire v_1893;
wire v_1894;
wire v_1895;
wire v_1896;
wire v_1897;
wire v_1898;
wire v_1899;
wire v_1900;
wire v_1901;
wire v_1902;
wire v_1904;
wire v_1905;
wire v_1906;
wire v_1907;
wire v_1908;
wire v_1909;
wire v_1910;
wire v_1911;
wire v_1912;
wire v_1913;
wire v_1914;
wire v_1915;
wire v_1916;
wire v_1917;
wire v_1918;
wire v_1919;
wire v_1920;
wire v_1921;
wire v_1922;
wire v_1923;
wire v_1924;
wire v_1925;
wire v_1926;
wire v_1927;
wire v_1928;
wire v_1929;
wire v_1930;
wire v_1931;
wire v_1932;
wire v_1933;
wire v_1934;
wire v_1935;
wire v_1936;
wire v_1937;
wire v_1938;
wire v_1939;
wire v_1940;
wire v_1941;
wire v_1942;
wire v_1943;
wire v_1944;
wire v_1945;
wire v_1946;
wire v_1947;
wire v_1948;
wire v_1949;
wire v_1950;
wire v_1951;
wire v_1952;
wire v_1953;
wire v_1954;
wire v_1955;
wire v_1956;
wire v_1957;
wire v_1958;
wire v_1959;
wire v_1960;
wire v_1961;
wire v_1962;
wire v_1963;
wire v_1964;
wire v_1965;
wire v_1966;
wire v_1967;
wire v_1968;
wire v_1969;
wire v_1970;
wire v_1971;
wire v_1972;
wire v_1973;
wire v_1974;
wire v_1975;
wire v_1976;
wire v_1977;
wire v_1978;
wire v_1979;
wire v_1980;
wire v_1981;
wire v_1982;
wire v_1983;
wire v_1984;
wire v_1985;
wire v_1986;
wire v_1987;
wire v_1988;
wire v_1989;
wire v_1990;
wire v_1991;
wire v_1992;
wire v_1993;
wire v_1994;
wire v_1995;
wire v_1996;
wire v_1997;
wire v_1998;
wire v_1999;
wire v_2000;
wire v_2001;
wire v_2002;
wire v_2003;
wire v_2004;
wire v_2005;
wire v_2006;
wire v_2007;
wire v_2008;
wire v_2009;
wire v_2010;
wire v_2011;
wire v_2012;
wire v_2013;
wire v_2014;
wire v_2015;
wire v_2016;
wire v_2017;
wire v_2018;
wire v_2019;
wire v_2020;
wire v_2021;
wire v_2022;
wire v_2023;
wire v_2024;
wire v_2025;
wire v_2026;
wire v_2027;
wire v_2028;
wire v_2029;
wire v_2030;
wire v_2031;
wire v_2032;
wire v_2033;
wire v_2034;
wire v_2035;
wire v_2036;
wire v_2037;
wire v_2038;
wire v_2039;
wire v_2040;
wire v_2041;
wire v_2042;
wire v_2043;
wire v_2044;
wire v_2045;
wire v_2046;
wire v_2047;
wire v_2048;
wire v_2049;
wire v_2050;
wire v_2051;
wire v_2052;
wire v_2053;
wire v_2054;
wire v_2055;
wire v_2056;
wire v_2057;
wire v_2058;
wire v_2059;
wire v_2060;
wire v_2061;
wire v_2062;
wire v_2063;
wire v_2064;
wire v_2065;
wire v_2066;
wire v_2067;
wire v_2068;
wire v_2069;
wire v_2070;
wire v_2071;
wire v_2072;
wire v_2073;
wire v_2074;
wire v_2075;
wire v_2076;
wire v_2077;
wire v_2078;
wire v_2079;
wire v_2080;
wire v_2081;
wire v_2082;
wire v_2083;
wire v_2084;
wire v_2085;
wire v_2086;
wire v_2087;
wire v_2088;
wire v_2089;
wire v_2090;
wire v_2091;
wire v_2092;
wire v_2093;
wire v_2094;
wire v_2095;
wire v_2096;
wire v_2097;
wire v_2098;
wire v_2099;
wire v_2100;
wire v_2101;
wire v_2102;
wire v_2103;
wire v_2104;
wire v_2105;
wire v_2106;
wire v_2107;
wire v_2108;
wire v_2109;
wire v_2110;
wire v_2111;
wire v_2112;
wire v_2113;
wire v_2114;
wire v_2115;
wire v_2116;
wire v_2117;
wire v_2118;
wire v_2119;
wire v_2120;
wire v_2121;
wire v_2122;
wire v_2123;
wire v_2124;
wire v_2125;
wire v_2126;
wire v_2127;
wire v_2128;
wire v_2129;
wire v_2130;
wire v_2131;
wire v_2132;
wire v_2133;
wire v_2134;
wire v_2135;
wire v_2136;
wire v_2138;
wire v_2139;
wire v_2140;
wire v_2141;
wire v_2142;
wire v_2143;
wire v_2144;
wire v_2145;
wire v_2146;
wire v_2147;
wire v_2148;
wire v_2149;
wire v_2150;
wire v_2151;
wire v_2152;
wire v_2153;
wire v_2154;
wire v_2155;
wire v_2156;
wire v_2158;
wire v_2159;
wire v_2160;
wire v_2161;
wire v_2162;
wire v_2163;
wire v_2164;
wire v_2165;
wire v_2166;
wire v_2167;
wire v_2168;
wire v_2169;
wire v_2170;
wire v_2171;
wire v_2172;
wire v_2173;
wire v_2174;
wire v_2175;
wire v_2176;
wire v_2177;
wire v_2178;
wire v_2179;
wire v_2180;
wire v_2181;
wire v_2182;
wire v_2183;
wire v_2184;
wire v_2185;
wire v_2186;
wire v_2187;
wire v_2188;
wire v_2189;
wire v_2190;
wire v_2191;
wire v_2192;
wire v_2193;
wire v_2194;
wire v_2195;
wire v_2196;
wire v_2197;
wire v_2198;
wire v_2199;
wire v_2200;
wire v_2201;
wire v_2202;
wire v_2203;
wire v_2204;
wire v_2205;
wire v_2206;
wire v_2207;
wire v_2209;
wire v_2210;
wire v_2211;
wire v_2212;
wire v_2213;
wire v_2214;
wire v_2215;
wire v_2216;
wire v_2217;
wire v_2218;
wire v_2219;
wire v_2220;
wire v_2221;
wire v_2222;
wire v_2223;
wire v_2224;
wire v_2225;
wire v_2227;
wire v_2228;
wire v_2229;
wire v_2230;
wire v_2231;
wire v_2232;
wire v_2233;
wire v_2234;
wire v_2235;
wire v_2236;
wire v_2237;
wire v_2238;
wire v_2239;
wire v_2240;
wire v_2241;
wire v_2242;
wire v_2243;
wire v_2244;
wire v_2245;
wire v_2246;
wire v_2247;
wire v_2248;
wire v_2249;
wire v_2250;
wire v_2251;
wire v_2252;
wire v_2253;
wire v_2254;
wire v_2255;
wire v_2256;
wire v_2257;
wire v_2258;
wire v_2259;
wire v_2260;
wire v_2261;
wire v_2262;
wire v_2263;
wire v_2264;
wire v_2265;
wire v_2266;
wire v_2267;
wire v_2268;
wire v_2269;
wire v_2270;
wire v_2271;
wire v_2272;
wire v_2273;
wire v_2274;
wire v_2275;
wire v_2276;
wire v_2277;
wire v_2278;
wire v_2279;
wire v_2280;
wire v_2281;
wire v_2282;
wire v_2283;
wire v_2284;
wire v_2285;
wire v_2286;
wire v_2287;
wire v_2288;
wire v_2289;
wire v_2290;
wire v_2291;
wire v_2292;
wire v_2293;
wire v_2294;
wire v_2295;
wire v_2296;
wire v_2297;
wire v_2298;
wire v_2299;
wire v_2300;
wire v_2301;
wire v_2302;
wire v_2303;
wire v_2304;
wire v_2305;
wire v_2306;
wire v_2307;
wire v_2308;
wire v_2309;
wire v_2310;
wire v_2311;
wire v_2312;
wire v_2313;
wire v_2314;
wire v_2315;
wire v_2316;
wire v_2317;
wire v_2318;
wire v_2319;
wire v_2320;
wire v_2321;
wire v_2322;
wire v_2323;
wire v_2324;
wire v_2325;
wire v_2326;
wire v_2327;
wire v_2328;
wire v_2329;
wire v_2330;
wire v_2331;
wire v_2332;
wire v_2333;
wire v_2334;
wire v_2335;
wire v_2336;
wire v_2337;
wire v_2339;
wire v_2340;
wire v_2341;
wire v_2342;
wire v_2343;
wire v_2344;
wire v_2345;
wire v_2346;
wire v_2347;
wire v_2348;
wire v_2349;
wire v_2350;
wire v_2351;
wire v_2352;
wire v_2353;
wire v_2354;
wire v_2355;
wire v_2356;
wire v_2357;
wire v_2358;
wire v_2359;
wire v_2360;
wire v_2361;
wire v_2362;
wire v_2363;
wire v_2364;
wire v_2365;
wire v_2366;
wire v_2367;
wire v_2368;
wire v_2369;
wire v_2370;
wire v_2371;
wire v_2372;
wire v_2373;
wire v_2374;
wire v_2375;
wire v_2376;
wire v_2377;
wire v_2378;
wire v_2379;
wire v_2380;
wire v_2381;
wire v_2382;
wire v_2383;
wire v_2384;
wire v_2385;
wire v_2386;
wire v_2387;
wire v_2388;
wire v_2389;
wire v_2390;
wire v_2391;
wire v_2392;
wire v_2393;
wire v_2394;
wire v_2395;
wire v_2396;
wire v_2397;
wire v_2398;
wire v_2399;
wire v_2400;
wire v_2401;
wire v_2402;
wire v_2403;
wire v_2404;
wire v_2405;
wire v_2406;
wire v_2407;
wire v_2408;
wire v_2409;
wire v_2410;
wire v_2411;
wire v_2412;
wire v_2413;
wire v_2414;
wire v_2415;
wire v_2416;
wire v_2417;
wire v_2418;
wire v_2419;
wire v_2420;
wire v_2421;
wire v_2422;
wire v_2423;
wire v_2424;
wire v_2425;
wire v_2426;
wire v_2427;
wire v_2428;
wire v_2429;
wire v_2430;
wire v_2431;
wire v_2432;
wire v_2433;
wire v_2434;
wire v_2435;
wire v_2436;
wire v_2437;
wire v_2438;
wire v_2439;
wire v_2440;
wire v_2441;
wire v_2442;
wire v_2443;
wire v_2444;
wire v_2445;
wire v_2446;
wire v_2447;
wire v_2448;
wire v_2449;
wire v_2450;
wire v_2451;
wire v_2452;
wire v_2453;
wire v_2454;
wire v_2455;
wire v_2456;
wire v_2457;
wire v_2458;
wire v_2459;
wire v_2460;
wire v_2461;
wire v_2462;
wire v_2464;
wire v_2465;
wire v_2466;
wire v_2467;
wire v_2468;
wire v_2469;
wire v_2470;
wire v_2471;
wire v_2472;
wire v_2473;
wire v_2474;
wire v_2475;
wire v_2476;
wire v_2477;
wire v_2478;
wire v_2479;
wire v_2480;
wire v_2481;
wire v_2482;
wire v_2484;
wire v_2485;
wire v_2486;
wire v_2487;
wire v_2488;
wire v_2489;
wire v_2490;
wire v_2491;
wire v_2492;
wire v_2493;
wire v_2494;
wire v_2495;
wire v_2496;
wire v_2497;
wire v_2498;
wire v_2499;
wire v_2500;
wire v_2501;
wire v_2502;
wire v_2503;
wire v_2504;
wire v_2505;
wire v_2506;
wire v_2507;
wire v_2508;
wire v_2509;
wire v_2510;
wire v_2511;
wire v_2512;
wire v_2513;
wire v_2514;
wire v_2515;
wire v_2516;
wire v_2517;
wire v_2518;
wire v_2519;
wire v_2520;
wire v_2521;
wire v_2522;
wire v_2523;
wire v_2524;
wire v_2525;
wire v_2526;
wire v_2527;
wire v_2528;
wire v_2529;
wire v_2530;
wire v_2531;
wire v_2532;
wire v_2533;
wire v_2535;
wire v_2536;
wire v_2537;
wire v_2538;
wire v_2539;
wire v_2540;
wire v_2541;
wire v_2542;
wire v_2543;
wire v_2544;
wire v_2545;
wire v_2546;
wire v_2547;
wire v_2548;
wire v_2549;
wire v_2550;
wire v_2551;
wire v_2553;
wire v_2554;
wire v_2555;
wire v_2556;
wire v_2557;
wire v_2558;
wire v_2559;
wire v_2560;
wire v_2561;
wire v_2562;
wire v_2563;
wire v_2564;
wire v_2565;
wire v_2566;
wire v_2567;
wire v_2568;
wire v_2569;
wire v_2570;
wire v_2571;
wire v_2572;
wire v_2573;
wire v_2574;
wire v_2575;
wire v_2576;
wire v_2577;
wire v_2578;
wire v_2579;
wire v_2580;
wire v_2581;
wire v_2582;
wire v_2583;
wire v_2584;
wire v_2585;
wire v_2586;
wire v_2587;
wire v_2588;
wire v_2589;
wire v_2590;
wire v_2591;
wire v_2592;
wire v_2593;
wire v_2594;
wire v_2595;
wire v_2596;
wire v_2597;
wire v_2598;
wire v_2599;
wire v_2600;
wire v_2601;
wire v_2602;
wire v_2603;
wire v_2604;
wire v_2605;
wire v_2606;
wire v_2607;
wire v_2608;
wire v_2609;
wire v_2610;
wire v_2611;
wire v_2612;
wire v_2613;
wire v_2614;
wire v_2615;
wire v_2616;
wire v_2617;
wire v_2618;
wire v_2619;
wire v_2620;
wire v_2621;
wire v_2622;
wire v_2623;
wire v_2624;
wire v_2625;
wire v_2626;
wire v_2627;
wire v_2628;
wire v_2629;
wire v_2630;
wire v_2631;
wire v_2632;
wire v_2633;
wire v_2634;
wire v_2635;
wire v_2636;
wire v_2637;
wire v_2638;
wire v_2639;
wire v_2640;
wire v_2641;
wire v_2642;
wire v_2643;
wire v_2644;
wire v_2645;
wire v_2646;
wire v_2647;
wire v_2648;
wire v_2649;
wire v_2650;
wire v_2651;
wire v_2652;
wire v_2653;
wire v_2654;
wire v_2655;
wire v_2656;
wire v_2657;
wire v_2658;
wire v_2659;
wire v_2660;
wire v_2661;
wire v_2662;
wire v_2663;
wire v_2665;
wire v_2666;
wire v_2667;
wire v_2668;
wire v_2669;
wire v_2670;
wire v_2671;
wire v_2672;
wire v_2673;
wire v_2674;
wire v_2675;
wire v_2676;
wire v_2677;
wire v_2678;
wire v_2679;
wire v_2680;
wire v_2681;
wire v_2682;
wire v_2683;
wire v_2684;
wire v_2685;
wire v_2686;
wire v_2687;
wire v_2688;
wire v_2689;
wire v_2690;
wire v_2691;
wire v_2692;
wire v_2693;
wire v_2694;
wire v_2695;
wire v_2696;
wire v_2697;
wire v_2698;
wire v_2699;
wire v_2700;
wire v_2701;
wire v_2702;
wire v_2703;
wire v_2704;
wire v_2705;
wire v_2706;
wire v_2707;
wire v_2708;
wire v_2709;
wire v_2710;
wire v_2711;
wire v_2712;
wire v_2713;
wire v_2714;
wire v_2715;
wire v_2716;
wire v_2717;
wire v_2718;
wire v_2719;
wire v_2720;
wire v_2721;
wire v_2722;
wire v_2723;
wire v_2724;
wire v_2725;
wire v_2726;
wire v_2727;
wire v_2728;
wire v_2729;
wire v_2730;
wire v_2731;
wire v_2732;
wire v_2733;
wire v_2734;
wire v_2735;
wire v_2736;
wire v_2737;
wire v_2738;
wire v_2739;
wire v_2740;
wire v_2741;
wire v_2742;
wire v_2743;
wire v_2744;
wire v_2745;
wire v_2746;
wire v_2747;
wire v_2748;
wire v_2749;
wire v_2750;
wire v_2751;
wire v_2752;
wire v_2753;
wire v_2754;
wire v_2755;
wire v_2756;
wire v_2757;
wire v_2758;
wire v_2759;
wire v_2760;
wire v_2761;
wire v_2762;
wire v_2763;
wire v_2764;
wire v_2765;
wire v_2766;
wire v_2767;
wire v_2768;
wire v_2769;
wire v_2770;
wire v_2771;
wire v_2772;
wire v_2773;
wire v_2774;
wire v_2775;
wire v_2776;
wire v_2777;
wire v_2778;
wire v_2779;
wire v_2780;
wire v_2781;
wire v_2782;
wire v_2783;
wire v_2784;
wire v_2785;
wire v_2786;
wire v_2787;
wire v_2788;
wire v_2790;
wire v_2791;
wire v_2792;
wire v_2793;
wire v_2794;
wire v_2795;
wire v_2796;
wire v_2797;
wire v_2798;
wire v_2799;
wire v_2800;
wire v_2801;
wire v_2802;
wire v_2803;
wire v_2804;
wire v_2805;
wire v_2806;
wire v_2807;
wire v_2808;
wire v_2810;
wire v_2811;
wire v_2812;
wire v_2813;
wire v_2814;
wire v_2815;
wire v_2816;
wire v_2817;
wire v_2818;
wire v_2819;
wire v_2820;
wire v_2821;
wire v_2822;
wire v_2823;
wire v_2824;
wire v_2825;
wire v_2826;
wire v_2827;
wire v_2828;
wire v_2829;
wire v_2830;
wire v_2831;
wire v_2832;
wire v_2833;
wire v_2834;
wire v_2835;
wire v_2836;
wire v_2837;
wire v_2838;
wire v_2839;
wire v_2840;
wire v_2841;
wire v_2842;
wire v_2843;
wire v_2844;
wire v_2845;
wire v_2846;
wire v_2847;
wire v_2848;
wire v_2849;
wire v_2850;
wire v_2851;
wire v_2852;
wire v_2853;
wire v_2854;
wire v_2855;
wire v_2856;
wire v_2857;
wire v_2858;
wire v_2859;
wire v_2861;
wire v_2862;
wire v_2863;
wire v_2864;
wire v_2865;
wire v_2866;
wire v_2867;
wire v_2868;
wire v_2869;
wire v_2870;
wire v_2871;
wire v_2872;
wire v_2873;
wire v_2874;
wire v_2875;
wire v_2876;
wire v_2877;
wire v_2879;
wire v_2880;
wire v_2881;
wire v_2882;
wire v_2883;
wire v_2884;
wire v_2885;
wire v_2886;
wire v_2887;
wire v_2888;
wire v_2889;
wire v_2890;
wire v_2891;
wire v_2892;
wire v_2893;
wire v_2894;
wire v_2895;
wire v_2896;
wire v_2897;
wire v_2898;
wire v_2899;
wire v_2900;
wire v_2901;
wire v_2902;
wire v_2903;
wire v_2904;
wire v_2905;
wire v_2906;
wire v_2907;
wire v_2908;
wire v_2909;
wire v_2910;
wire v_2911;
wire v_2912;
wire v_2913;
wire v_2914;
wire v_2915;
wire v_2916;
wire v_2917;
wire v_2918;
wire v_2919;
wire v_2920;
wire v_2921;
wire v_2922;
wire v_2923;
wire v_2924;
wire v_2925;
wire v_2926;
wire v_2927;
wire v_2928;
wire v_2929;
wire v_2930;
wire v_2931;
wire v_2932;
wire v_2933;
wire v_2934;
wire v_2935;
wire v_2936;
wire v_2937;
wire v_2938;
wire v_2939;
wire v_2940;
wire v_2941;
wire v_2942;
wire v_2943;
wire v_2944;
wire v_2945;
wire v_2946;
wire v_2947;
wire v_2948;
wire v_2949;
wire v_2950;
wire v_2951;
wire v_2952;
wire v_2953;
wire v_2954;
wire v_2955;
wire v_2956;
wire v_2957;
wire v_2958;
wire v_2959;
wire v_2960;
wire v_2961;
wire v_2962;
wire v_2963;
wire v_2964;
wire v_2965;
wire v_2966;
wire v_2967;
wire v_2968;
wire v_2969;
wire v_2970;
wire v_2971;
wire v_2972;
wire v_2973;
wire v_2974;
wire v_2975;
wire v_2976;
wire v_2977;
wire v_2978;
wire v_2979;
wire v_2980;
wire v_2981;
wire v_2982;
wire v_2983;
wire v_2984;
wire v_2985;
wire v_2986;
wire v_2987;
wire v_2988;
wire v_2989;
wire v_2990;
wire v_2991;
wire v_2992;
wire v_2993;
wire v_2994;
wire v_2995;
wire v_2996;
wire v_2997;
wire v_2998;
wire v_2999;
wire v_3000;
wire v_3001;
wire v_3002;
wire v_3003;
wire v_3004;
wire v_3005;
wire v_3006;
wire v_3007;
wire v_3008;
wire v_3009;
wire v_3010;
wire v_3011;
wire v_3012;
wire v_3013;
wire v_3014;
wire v_3015;
wire v_3016;
wire v_3017;
wire v_3018;
wire v_3019;
wire v_3020;
wire v_3021;
wire v_3022;
wire v_3023;
wire v_3024;
wire v_3025;
wire v_3026;
wire v_3027;
wire v_3028;
wire v_3029;
wire v_3030;
wire v_3031;
wire v_3032;
wire v_3033;
wire v_3034;
wire v_3035;
wire v_3036;
wire v_3037;
wire v_3038;
wire v_3039;
wire v_3040;
wire v_3041;
wire v_3042;
wire v_3043;
wire v_3044;
wire v_3045;
wire v_3046;
wire v_3047;
wire v_3048;
wire v_3049;
wire v_3050;
wire v_3051;
wire v_3052;
wire v_3053;
wire v_3054;
wire v_3055;
wire v_3056;
wire v_3057;
wire v_3058;
wire v_3059;
wire v_3060;
wire v_3061;
wire v_3062;
wire v_3063;
wire v_3064;
wire v_3065;
wire v_3066;
wire v_3067;
wire v_3068;
wire v_3069;
wire v_3070;
wire v_3071;
wire v_3072;
wire v_3073;
wire v_3074;
wire v_3075;
wire v_3076;
wire v_3077;
wire v_3078;
wire v_3079;
wire v_3080;
wire v_3081;
wire v_3082;
wire v_3083;
wire v_3084;
wire v_3085;
wire v_3086;
wire v_3087;
wire v_3088;
wire v_3089;
wire v_3090;
wire v_3091;
wire v_3092;
wire v_3093;
wire v_3094;
wire v_3095;
wire v_3096;
wire v_3097;
wire v_3098;
wire v_3099;
wire v_3100;
wire v_3101;
wire v_3102;
wire v_3103;
wire v_3104;
wire v_3105;
wire v_3106;
wire v_3107;
wire v_3108;
wire v_3109;
wire v_3110;
wire v_3111;
wire v_3112;
wire v_3113;
wire v_3115;
wire v_3116;
wire v_3117;
wire v_3118;
wire v_3119;
wire v_3120;
wire v_3121;
wire v_3122;
wire v_3123;
wire v_3124;
wire v_3125;
wire v_3126;
wire v_3127;
wire v_3128;
wire v_3129;
wire v_3130;
wire v_3131;
wire v_3132;
wire v_3133;
wire v_3135;
wire v_3136;
wire v_3137;
wire v_3138;
wire v_3139;
wire v_3140;
wire v_3141;
wire v_3142;
wire v_3143;
wire v_3144;
wire v_3145;
wire v_3146;
wire v_3147;
wire v_3148;
wire v_3149;
wire v_3150;
wire v_3151;
wire v_3152;
wire v_3153;
wire v_3154;
wire v_3155;
wire v_3156;
wire v_3157;
wire v_3158;
wire v_3159;
wire v_3160;
wire v_3161;
wire v_3162;
wire v_3163;
wire v_3164;
wire v_3165;
wire v_3166;
wire v_3167;
wire v_3168;
wire v_3169;
wire v_3170;
wire v_3171;
wire v_3172;
wire v_3173;
wire v_3174;
wire v_3175;
wire v_3176;
wire v_3177;
wire v_3178;
wire v_3179;
wire v_3180;
wire v_3181;
wire v_3182;
wire v_3183;
wire v_3184;
wire v_3186;
wire v_3187;
wire v_3188;
wire v_3189;
wire v_3190;
wire v_3191;
wire v_3192;
wire v_3193;
wire v_3194;
wire v_3195;
wire v_3196;
wire v_3197;
wire v_3198;
wire v_3199;
wire v_3200;
wire v_3201;
wire v_3202;
wire v_3204;
wire v_3205;
wire v_3206;
wire v_3207;
wire v_3208;
wire v_3209;
wire v_3210;
wire v_3211;
wire v_3212;
wire v_3213;
wire v_3214;
wire v_3215;
wire v_3216;
wire v_3217;
wire v_3218;
wire v_3219;
wire v_3220;
wire v_3221;
wire v_3222;
wire v_3223;
wire v_3224;
wire v_3225;
wire v_3226;
wire v_3227;
wire v_3228;
wire v_3229;
wire v_3230;
wire v_3231;
wire v_3232;
wire v_3233;
wire v_3234;
wire v_3235;
wire v_3236;
wire v_3237;
wire v_3238;
wire v_3239;
wire v_3240;
wire v_3241;
wire v_3242;
wire v_3243;
wire v_3244;
wire v_3245;
wire v_3246;
wire v_3247;
wire v_3248;
wire v_3249;
wire v_3250;
wire v_3251;
wire v_3252;
wire v_3253;
wire v_3254;
wire v_3255;
wire v_3256;
wire v_3257;
wire v_3258;
wire v_3259;
wire v_3260;
wire v_3261;
wire v_3262;
wire v_3263;
wire v_3264;
wire v_3265;
wire v_3266;
wire v_3267;
wire v_3268;
wire v_3269;
wire v_3270;
wire v_3271;
wire v_3272;
wire v_3273;
wire v_3274;
wire v_3275;
wire v_3276;
wire v_3277;
wire v_3278;
wire v_3279;
wire v_3280;
wire v_3281;
wire v_3282;
wire v_3283;
wire v_3284;
wire v_3285;
wire v_3286;
wire v_3287;
wire v_3288;
wire v_3289;
wire v_3290;
wire v_3291;
wire v_3292;
wire v_3293;
wire v_3294;
wire v_3295;
wire v_3296;
wire v_3297;
wire v_3298;
wire v_3299;
wire v_3300;
wire v_3301;
wire v_3302;
wire v_3303;
wire v_3304;
wire v_3305;
wire v_3306;
wire v_3307;
wire v_3308;
wire v_3309;
wire v_3310;
wire v_3311;
wire v_3312;
wire v_3313;
wire v_3314;
wire v_3316;
wire v_3317;
wire v_3318;
wire v_3319;
wire v_3320;
wire v_3321;
wire v_3322;
wire v_3323;
wire v_3324;
wire v_3325;
wire v_3326;
wire v_3327;
wire v_3328;
wire v_3329;
wire v_3330;
wire v_3331;
wire v_3332;
wire v_3333;
wire v_3334;
wire v_3335;
wire v_3336;
wire v_3337;
wire v_3338;
wire v_3339;
wire v_3340;
wire v_3341;
wire v_3342;
wire v_3343;
wire v_3344;
wire v_3345;
wire v_3346;
wire v_3347;
wire v_3348;
wire v_3349;
wire v_3350;
wire v_3351;
wire v_3352;
wire v_3353;
wire v_3354;
wire v_3355;
wire v_3356;
wire v_3357;
wire v_3358;
wire v_3359;
wire v_3360;
wire v_3361;
wire v_3362;
wire v_3363;
wire v_3364;
wire v_3365;
wire v_3366;
wire v_3367;
wire v_3368;
wire v_3369;
wire v_3370;
wire v_3371;
wire v_3372;
wire v_3373;
wire v_3374;
wire v_3375;
wire v_3376;
wire v_3377;
wire v_3378;
wire v_3379;
wire v_3380;
wire v_3381;
wire v_3382;
wire v_3383;
wire v_3384;
wire v_3385;
wire v_3386;
wire v_3387;
wire v_3388;
wire v_3389;
wire v_3390;
wire v_3391;
wire v_3392;
wire v_3393;
wire v_3394;
wire v_3395;
wire v_3396;
wire v_3397;
wire v_3398;
wire v_3399;
wire v_3400;
wire v_3401;
wire v_3402;
wire v_3403;
wire v_3404;
wire v_3405;
wire v_3406;
wire v_3407;
wire v_3408;
wire v_3409;
wire v_3410;
wire v_3411;
wire v_3412;
wire v_3413;
wire v_3414;
wire v_3415;
wire v_3416;
wire v_3417;
wire v_3418;
wire v_3419;
wire v_3420;
wire v_3421;
wire v_3422;
wire v_3423;
wire v_3424;
wire v_3425;
wire v_3426;
wire v_3427;
wire v_3428;
wire v_3429;
wire v_3430;
wire v_3431;
wire v_3432;
wire v_3433;
wire v_3434;
wire v_3435;
wire v_3436;
wire v_3437;
wire v_3438;
wire v_3439;
wire v_3441;
wire v_3442;
wire v_3443;
wire v_3444;
wire v_3445;
wire v_3446;
wire v_3447;
wire v_3448;
wire v_3449;
wire v_3450;
wire v_3451;
wire v_3452;
wire v_3453;
wire v_3454;
wire v_3455;
wire v_3456;
wire v_3457;
wire v_3458;
wire v_3459;
wire v_3461;
wire v_3462;
wire v_3463;
wire v_3464;
wire v_3465;
wire v_3466;
wire v_3467;
wire v_3468;
wire v_3469;
wire v_3470;
wire v_3471;
wire v_3472;
wire v_3473;
wire v_3474;
wire v_3475;
wire v_3476;
wire v_3477;
wire v_3478;
wire v_3479;
wire v_3480;
wire v_3481;
wire v_3482;
wire v_3483;
wire v_3484;
wire v_3485;
wire v_3486;
wire v_3487;
wire v_3488;
wire v_3489;
wire v_3490;
wire v_3491;
wire v_3492;
wire v_3493;
wire v_3494;
wire v_3495;
wire v_3496;
wire v_3497;
wire v_3498;
wire v_3499;
wire v_3500;
wire v_3501;
wire v_3502;
wire v_3503;
wire v_3504;
wire v_3505;
wire v_3506;
wire v_3507;
wire v_3508;
wire v_3509;
wire v_3510;
wire v_3512;
wire v_3513;
wire v_3514;
wire v_3515;
wire v_3516;
wire v_3517;
wire v_3518;
wire v_3519;
wire v_3520;
wire v_3521;
wire v_3522;
wire v_3523;
wire v_3524;
wire v_3525;
wire v_3526;
wire v_3527;
wire v_3528;
wire v_3530;
wire v_3531;
wire v_3532;
wire v_3533;
wire v_3534;
wire v_3535;
wire v_3536;
wire v_3537;
wire v_3538;
wire v_3539;
wire v_3540;
wire v_3541;
wire v_3542;
wire v_3543;
wire v_3544;
wire v_3545;
wire v_3546;
wire v_3547;
wire v_3548;
wire v_3549;
wire v_3550;
wire v_3551;
wire v_3552;
wire v_3553;
wire v_3554;
wire v_3555;
wire v_3556;
wire v_3557;
wire v_3558;
wire v_3559;
wire v_3560;
wire v_3561;
wire v_3562;
wire v_3563;
wire v_3564;
wire v_3565;
wire v_3566;
wire v_3567;
wire v_3568;
wire v_3569;
wire v_3570;
wire v_3571;
wire v_3572;
wire v_3573;
wire v_3574;
wire v_3575;
wire v_3576;
wire v_3577;
wire v_3578;
wire v_3579;
wire v_3580;
wire v_3581;
wire v_3582;
wire v_3583;
wire v_3584;
wire v_3585;
wire v_3586;
wire v_3587;
wire v_3588;
wire v_3589;
wire v_3590;
wire v_3591;
wire v_3592;
wire v_3593;
wire v_3594;
wire v_3595;
wire v_3596;
wire v_3597;
wire v_3598;
wire v_3599;
wire v_3600;
wire v_3601;
wire v_3602;
wire v_3603;
wire v_3604;
wire v_3605;
wire v_3606;
wire v_3607;
wire v_3608;
wire v_3609;
wire v_3610;
wire v_3611;
wire v_3612;
wire v_3613;
wire v_3614;
wire v_3615;
wire v_3616;
wire v_3617;
wire v_3618;
wire v_3619;
wire v_3620;
wire v_3621;
wire v_3622;
wire v_3623;
wire v_3624;
wire v_3625;
wire v_3626;
wire v_3627;
wire v_3628;
wire v_3629;
wire v_3630;
wire v_3631;
wire v_3632;
wire v_3633;
wire v_3634;
wire v_3635;
wire v_3636;
wire v_3637;
wire v_3638;
wire v_3639;
wire v_3640;
wire v_3642;
wire v_3643;
wire v_3644;
wire v_3645;
wire v_3647;
wire v_3648;
wire v_3649;
wire v_3650;
wire v_3651;
wire v_3652;
wire v_3653;
wire v_3654;
wire v_3655;
wire v_3656;
wire v_3657;
wire v_3658;
wire v_3659;
wire v_3660;
wire v_3661;
wire v_3662;
wire v_3663;
wire v_3664;
wire v_3665;
wire v_3666;
wire v_3667;
wire v_3668;
wire v_3669;
wire v_3670;
wire v_3671;
wire v_3672;
wire v_3673;
wire v_3674;
wire v_3675;
wire v_3676;
wire v_3677;
wire v_3678;
wire v_3679;
wire v_3680;
wire v_3681;
wire v_3682;
wire v_3683;
wire v_3684;
wire v_3685;
wire v_3686;
wire v_3687;
wire v_3688;
wire v_3689;
wire v_3690;
wire v_3691;
wire v_3692;
wire v_3693;
wire v_3694;
wire v_3695;
wire v_3696;
wire v_3697;
wire v_3698;
wire v_3699;
wire v_3700;
wire v_3701;
wire v_3702;
wire v_3703;
wire v_3704;
wire v_3705;
wire v_3706;
wire v_3707;
wire v_3708;
wire v_3709;
wire v_3710;
wire v_3711;
wire v_3712;
wire v_3713;
wire v_3714;
wire v_3715;
wire v_3716;
wire v_3717;
wire v_3718;
wire v_3719;
wire v_3720;
wire v_3721;
wire v_3722;
wire v_3723;
wire v_3724;
wire v_3725;
wire v_3726;
wire v_3727;
wire v_3728;
wire v_3729;
wire v_3730;
wire v_3731;
wire v_3732;
wire v_3733;
wire v_3734;
wire v_3735;
wire v_3736;
wire v_3737;
wire v_3738;
wire v_3739;
wire v_3740;
wire v_3742;
wire v_3743;
wire v_3744;
wire v_3745;
wire v_3746;
wire v_3747;
wire v_3748;
wire v_3749;
wire v_3750;
wire v_3751;
wire v_3752;
wire v_3753;
wire v_3754;
wire v_3755;
wire v_3756;
wire v_3757;
wire v_3758;
wire v_3759;
wire v_3760;
wire v_3761;
wire v_3762;
wire v_3763;
wire v_3764;
wire v_3765;
wire v_3766;
wire v_3767;
wire v_3768;
wire v_3769;
wire v_3770;
wire v_3771;
wire v_3772;
wire v_3773;
wire v_3774;
wire v_3775;
wire v_3776;
wire v_3777;
wire v_3778;
wire v_3779;
wire v_3780;
wire v_3781;
wire v_3782;
wire v_3783;
wire v_3784;
wire v_3785;
wire v_3786;
wire v_3787;
wire v_3788;
wire v_3789;
wire v_3790;
wire v_3791;
wire v_3792;
wire v_3793;
wire v_3794;
wire v_3795;
wire v_3796;
wire v_3797;
wire v_3798;
wire v_3799;
wire v_3800;
wire v_3801;
wire v_3802;
wire v_3803;
wire v_3804;
wire v_3805;
wire v_3806;
wire v_3807;
wire v_3808;
wire v_3809;
wire v_3810;
wire v_3811;
wire v_3812;
wire v_3813;
wire v_3814;
wire v_3815;
wire v_3816;
wire v_3817;
wire v_3818;
wire v_3819;
wire v_3820;
wire v_3821;
wire v_3822;
wire v_3823;
wire v_3824;
wire v_3825;
wire v_3826;
wire v_3827;
wire v_3828;
wire v_3829;
wire v_3830;
wire v_3831;
wire v_3832;
wire v_3833;
wire v_3834;
wire v_3835;
wire v_3836;
wire v_3837;
wire v_3838;
wire v_3839;
wire v_3840;
wire v_3841;
wire v_3842;
wire v_3843;
wire v_3844;
wire v_3845;
wire v_3846;
wire v_3847;
wire v_3848;
wire v_3849;
wire v_3850;
wire v_3851;
wire v_3852;
wire v_3853;
wire v_3854;
wire v_3855;
wire v_3856;
wire v_3857;
wire v_3858;
wire v_3859;
wire v_3860;
wire v_3861;
wire v_3862;
wire v_3863;
wire v_3864;
wire v_3865;
wire v_3866;
wire v_3867;
wire v_3868;
wire v_3869;
wire v_3870;
wire v_3871;
wire v_3872;
wire v_3873;
wire v_3874;
wire v_3875;
wire v_3876;
wire v_3877;
wire v_3878;
wire v_3879;
wire v_3880;
wire v_3881;
wire v_3882;
wire v_3883;
wire v_3884;
wire v_3885;
wire v_3886;
wire v_3887;
wire v_3888;
wire v_3889;
wire v_3890;
wire v_3891;
wire v_3892;
wire v_3893;
wire v_3894;
wire v_3895;
wire v_3896;
wire v_3897;
wire v_3898;
wire v_3899;
wire v_3900;
wire v_3901;
wire v_3902;
wire v_3903;
wire v_3904;
wire v_3905;
wire v_3906;
wire v_3907;
wire v_3908;
wire v_3909;
wire v_3910;
wire v_3911;
wire v_3912;
wire v_3913;
wire v_3914;
wire v_3915;
wire v_3916;
wire v_3917;
wire v_3918;
wire v_3919;
wire v_3920;
wire v_3921;
wire v_3922;
wire v_3923;
wire v_3924;
wire v_3925;
wire v_3926;
wire v_3927;
wire v_3928;
wire v_3929;
wire v_3930;
wire v_3931;
wire v_3933;
wire v_3934;
wire v_3935;
wire v_3936;
wire v_3937;
wire v_3938;
wire v_3939;
wire v_3940;
wire v_3941;
wire v_3942;
wire v_3943;
wire v_3944;
wire v_3945;
wire v_3946;
wire v_3947;
wire v_3948;
wire v_3949;
wire v_3950;
wire v_3951;
wire v_3952;
wire v_3953;
wire v_3954;
wire v_3955;
wire v_3956;
wire v_3957;
wire v_3958;
wire v_3959;
wire v_3960;
wire v_3961;
wire v_3962;
wire v_3963;
wire v_3964;
wire v_3965;
wire v_3966;
wire v_3967;
wire v_3968;
wire v_3969;
wire v_3970;
wire v_3971;
wire v_3972;
wire v_3973;
wire v_3974;
wire v_3975;
wire v_3976;
wire v_3977;
wire v_3978;
wire v_3979;
wire v_3980;
wire v_3981;
wire v_3982;
wire v_3983;
wire v_3984;
wire v_3985;
wire v_3986;
wire v_3987;
wire v_3988;
wire v_3989;
wire v_3990;
wire v_3991;
wire v_3992;
wire v_3993;
wire v_3994;
wire v_3995;
wire v_3996;
wire v_3997;
wire v_3998;
wire v_3999;
wire v_4000;
wire v_4001;
wire v_4002;
wire v_4003;
wire v_4004;
wire v_4005;
wire v_4006;
wire v_4007;
wire v_4008;
wire v_4009;
wire v_4010;
wire v_4011;
wire v_4012;
wire v_4013;
wire v_4014;
wire v_4015;
wire v_4016;
wire v_4017;
wire v_4018;
wire v_4019;
wire v_4020;
wire v_4021;
wire v_4022;
wire v_4023;
wire v_4024;
wire v_4025;
wire v_4026;
wire v_4027;
wire v_4028;
wire v_4029;
wire v_4030;
wire v_4031;
wire v_4032;
wire v_4033;
wire v_4034;
wire v_4035;
wire v_4036;
wire v_4037;
wire v_4038;
wire v_4039;
wire v_4040;
wire v_4041;
wire v_4042;
wire v_4043;
wire v_4044;
wire v_4045;
wire v_4046;
wire v_4047;
wire v_4048;
wire v_4049;
wire v_4050;
wire v_4051;
wire v_4052;
wire v_4053;
wire v_4054;
wire v_4055;
wire v_4056;
wire v_4058;
wire v_4059;
wire v_4060;
wire v_4061;
wire v_4062;
wire v_4063;
wire v_4064;
wire v_4065;
wire v_4066;
wire v_4067;
wire v_4068;
wire v_4069;
wire v_4070;
wire v_4071;
wire v_4072;
wire v_4073;
wire v_4074;
wire v_4075;
wire v_4076;
wire v_4078;
wire v_4079;
wire v_4080;
wire v_4081;
wire v_4082;
wire v_4083;
wire v_4084;
wire v_4085;
wire v_4086;
wire v_4087;
wire v_4088;
wire v_4089;
wire v_4090;
wire v_4091;
wire v_4092;
wire v_4093;
wire v_4094;
wire v_4095;
wire v_4096;
wire v_4097;
wire v_4098;
wire v_4099;
wire v_4100;
wire v_4101;
wire v_4102;
wire v_4103;
wire v_4104;
wire v_4105;
wire v_4106;
wire v_4107;
wire v_4108;
wire v_4109;
wire v_4110;
wire v_4111;
wire v_4112;
wire v_4113;
wire v_4114;
wire v_4115;
wire v_4116;
wire v_4117;
wire v_4118;
wire v_4119;
wire v_4120;
wire v_4121;
wire v_4122;
wire v_4123;
wire v_4124;
wire v_4125;
wire v_4126;
wire v_4127;
wire v_4129;
wire v_4130;
wire v_4131;
wire v_4132;
wire v_4133;
wire v_4134;
wire v_4135;
wire v_4136;
wire v_4137;
wire v_4138;
wire v_4139;
wire v_4140;
wire v_4141;
wire v_4142;
wire v_4143;
wire v_4144;
wire v_4145;
wire v_4147;
wire v_4148;
wire v_4149;
wire v_4150;
wire v_4151;
wire v_4152;
wire v_4153;
wire v_4154;
wire v_4155;
wire v_4156;
wire v_4157;
wire v_4158;
wire v_4159;
wire v_4160;
wire v_4161;
wire v_4162;
wire v_4163;
wire v_4164;
wire v_4165;
wire v_4166;
wire v_4167;
wire v_4168;
wire v_4169;
wire v_4170;
wire v_4171;
wire v_4172;
wire v_4173;
wire v_4174;
wire v_4175;
wire v_4176;
wire v_4177;
wire v_4178;
wire v_4179;
wire v_4180;
wire v_4181;
wire v_4182;
wire v_4183;
wire v_4184;
wire v_4185;
wire v_4186;
wire v_4187;
wire v_4188;
wire v_4189;
wire v_4190;
wire v_4191;
wire v_4192;
wire v_4193;
wire v_4194;
wire v_4195;
wire v_4196;
wire v_4197;
wire v_4198;
wire v_4199;
wire v_4200;
wire v_4201;
wire v_4202;
wire v_4203;
wire v_4204;
wire v_4205;
wire v_4206;
wire v_4207;
wire v_4208;
wire v_4209;
wire v_4210;
wire v_4211;
wire v_4212;
wire v_4213;
wire v_4214;
wire v_4215;
wire v_4216;
wire v_4217;
wire v_4218;
wire v_4219;
wire v_4220;
wire v_4221;
wire v_4222;
wire v_4223;
wire v_4224;
wire v_4225;
wire v_4226;
wire v_4227;
wire v_4228;
wire v_4229;
wire v_4230;
wire v_4231;
wire v_4232;
wire v_4233;
wire v_4234;
wire v_4235;
wire v_4236;
wire v_4237;
wire v_4238;
wire v_4239;
wire v_4240;
wire v_4241;
wire v_4242;
wire v_4243;
wire v_4244;
wire v_4245;
wire v_4246;
wire v_4247;
wire v_4248;
wire v_4249;
wire v_4250;
wire v_4251;
wire v_4252;
wire v_4253;
wire v_4254;
wire v_4255;
wire v_4256;
wire v_4257;
wire v_4262;
wire v_4265;
wire v_4266;
wire v_4267;
wire v_4268;
wire v_4269;
wire v_4270;
wire v_4271;
wire v_4272;
wire v_4273;
wire v_4274;
wire v_4275;
wire v_4276;
wire v_4277;
wire v_4278;
wire v_4279;
wire v_4280;
wire v_4281;
wire v_4282;
wire v_4283;
wire v_4284;
wire v_4285;
wire v_4286;
wire v_4287;
wire v_4288;
wire v_4289;
wire v_4290;
wire v_4291;
wire v_4292;
wire v_4293;
wire v_4294;
wire v_4295;
wire v_4296;
wire v_4297;
wire v_4298;
wire v_4299;
wire v_4300;
wire v_4301;
wire v_4302;
wire v_4303;
wire v_4304;
wire v_4305;
wire v_4306;
wire v_4307;
wire v_4308;
wire v_4309;
wire v_4310;
wire v_4311;
wire v_4312;
wire v_4313;
wire v_4314;
wire v_4315;
wire v_4316;
wire v_4317;
wire v_4318;
wire v_4319;
wire v_4320;
wire v_4321;
wire v_4322;
wire v_4323;
wire v_4324;
wire v_4325;
wire v_4326;
wire v_4327;
wire v_4328;
wire v_4329;
wire v_4330;
wire v_4331;
wire v_4332;
wire v_4333;
wire v_4334;
wire v_4335;
wire v_4336;
wire v_4337;
wire v_4338;
wire v_4339;
wire v_4340;
wire v_4341;
wire v_4342;
wire v_4343;
wire v_4344;
wire v_4345;
wire v_4346;
wire v_4347;
wire v_4348;
wire v_4349;
wire v_4350;
wire v_4351;
wire v_4352;
wire v_4353;
wire v_4354;
wire v_4355;
wire v_4356;
wire v_4357;
wire v_4358;
wire v_4359;
wire v_4360;
wire v_4361;
wire v_4362;
wire v_4363;
wire v_4364;
wire v_4365;
wire v_4366;
wire v_4367;
wire v_4368;
wire v_4369;
wire v_4370;
wire v_4371;
wire v_4372;
wire v_4373;
wire v_4374;
wire v_4375;
wire v_4376;
wire v_4377;
wire v_4378;
wire v_4379;
wire v_4380;
wire v_4381;
wire v_4382;
wire v_4383;
wire v_4384;
wire v_4385;
wire v_4386;
wire v_4387;
wire v_4388;
wire v_4389;
wire v_4390;
wire v_4391;
wire v_4392;
wire v_4393;
wire v_4394;
wire v_4395;
wire v_4396;
wire v_4397;
wire v_4398;
wire v_4399;
wire v_4400;
wire v_4401;
wire v_4402;
wire v_4403;
wire v_4404;
wire v_4405;
wire v_4406;
wire v_4407;
wire v_4408;
wire v_4409;
wire v_4410;
wire v_4411;
wire v_4412;
wire v_4413;
wire v_4414;
wire v_4415;
wire v_4416;
wire v_4417;
wire v_4418;
wire v_4419;
wire v_4420;
wire v_4421;
wire v_4422;
wire v_4423;
wire v_4424;
wire v_4425;
wire v_4426;
wire v_4427;
wire v_4428;
wire v_4429;
wire v_4430;
wire v_4431;
wire v_4432;
wire v_4433;
wire v_4434;
wire v_4435;
wire v_4436;
wire v_4437;
wire v_4438;
wire v_4439;
wire v_4440;
wire v_4441;
wire v_4442;
wire v_4443;
wire v_4444;
wire v_4445;
wire v_4446;
wire v_4447;
wire v_4448;
wire v_4449;
wire v_4450;
wire v_4451;
wire v_4452;
wire v_4453;
wire v_4454;
wire v_4455;
wire v_4456;
wire v_4457;
wire v_4458;
wire v_4459;
wire v_4460;
wire v_4461;
wire v_4462;
wire v_4463;
wire v_4464;
wire v_4465;
wire v_4466;
wire v_4467;
wire v_4468;
wire v_4471;
wire v_4472;
wire v_4473;
wire v_4474;
wire v_4476;
wire v_4478;
wire v_4479;
wire v_4480;
wire v_4482;
wire v_4484;
wire v_4487;
wire v_4489;
wire v_4491;
wire v_4494;
wire v_4496;
wire v_4498;
wire v_4500;
wire v_4502;
wire v_4504;
wire v_4506;
wire v_4508;
wire v_4509;
wire v_4512;
wire v_4513;
wire v_4514;
wire v_4515;
wire v_4516;
wire v_4517;
wire v_4519;
wire v_4521;
wire v_4522;
wire v_4523;
wire v_4525;
wire v_4526;
wire v_4527;
wire v_4529;
wire v_4531;
wire v_4532;
wire v_4533;
wire v_4534;
wire v_4538;
wire v_4540;
wire v_4541;
wire v_4543;
wire v_4545;
wire v_4546;
wire v_4547;
wire v_4550;
wire v_4552;
wire v_4555;
wire v_4556;
wire v_4557;
wire v_4558;
wire v_4560;
wire v_4561;
wire v_4562;
wire v_4563;
wire v_4566;
wire v_4569;
wire v_4570;
wire v_4571;
wire v_4573;
wire v_4575;
wire v_4576;
wire v_4577;
wire v_4579;
wire v_4581;
wire v_4583;
wire v_4584;
wire v_4585;
wire v_4586;
wire v_4587;
wire v_4588;
wire v_4591;
wire v_4593;
wire v_4595;
wire v_4597;
wire v_4598;
wire v_4599;
wire v_4600;
wire v_4603;
wire v_4605;
wire v_4607;
wire v_4609;
wire v_4611;
wire v_4612;
wire v_4614;
wire v_4617;
wire v_4619;
wire v_4621;
wire v_4623;
wire v_4624;
wire v_4625;
wire v_4627;
wire v_4630;
wire v_4632;
wire v_4634;
wire v_4636;
wire v_4638;
wire v_4639;
wire v_4640;
wire v_4642;
wire v_4643;
wire v_4644;
wire v_4646;
wire v_4649;
wire v_4651;
wire v_4653;
wire v_4655;
wire v_4657;
wire v_4658;
wire v_4659;
wire v_4660;
wire v_4661;
wire v_4663;
wire v_4664;
wire v_4665;
wire v_4668;
wire v_4670;
wire v_4672;
wire v_4674;
wire v_4676;
wire v_4677;
wire v_4679;
wire v_4682;
wire v_4684;
wire v_4686;
wire v_4688;
wire v_4689;
wire v_4690;
wire v_4692;
wire v_4695;
wire v_4697;
wire v_4699;
wire v_4701;
wire v_4703;
wire v_4704;
wire v_4705;
wire v_4707;
wire v_4708;
wire v_4709;
wire v_4711;
wire v_4714;
wire v_4716;
wire v_4718;
wire v_4720;
wire v_4722;
wire v_4723;
wire v_4724;
wire v_4725;
wire v_4726;
wire v_4728;
wire v_4729;
wire v_4730;
wire v_4732;
wire v_4734;
wire v_4735;
wire v_4736;
wire v_4738;
wire v_4739;
wire v_4740;
wire v_4741;
wire v_4743;
wire v_4744;
wire v_4746;
wire v_4748;
wire v_4751;
wire v_4753;
wire v_4755;
wire v_4758;
wire v_4760;
wire v_4762;
wire v_4764;
wire v_4766;
wire v_4768;
wire v_4770;
wire v_4772;
wire v_4773;
wire v_4776;
wire v_4777;
wire v_4778;
wire v_4779;
wire v_4780;
wire v_4781;
wire v_4783;
wire v_4785;
wire v_4786;
wire v_4787;
wire v_4789;
wire v_4790;
wire v_4791;
wire v_4792;
wire v_4794;
wire v_4795;
wire v_4796;
wire v_4797;
wire v_4800;
wire v_4801;
wire v_4802;
wire v_4804;
wire v_4806;
wire v_4808;
wire v_4809;
wire v_4810;
wire v_4812;
wire v_4813;
wire v_4814;
wire v_4816;
wire v_4818;
wire v_4820;
wire v_4822;
wire v_4823;
wire v_4824;
wire v_4826;
wire v_4828;
wire v_4831;
wire v_4832;
wire v_4833;
wire v_4835;
wire v_4836;
wire v_4837;
wire v_4838;
wire v_4841;
wire v_4843;
wire v_4844;
wire v_4846;
wire v_4848;
wire v_4849;
wire v_4851;
wire v_4852;
wire v_4853;
wire v_4854;
wire v_4855;
wire v_4858;
wire v_4859;
wire v_4860;
wire v_4862;
wire v_4864;
wire v_4866;
wire v_4867;
wire v_4868;
wire v_4870;
wire v_4871;
wire v_4872;
wire v_4874;
wire v_4876;
wire v_4878;
wire v_4880;
wire v_4881;
wire v_4882;
wire v_4884;
wire v_4886;
wire v_4889;
wire v_4890;
wire v_4891;
wire v_4893;
wire v_4894;
wire v_4895;
wire v_4896;
wire v_4898;
wire v_4900;
wire v_4902;
wire v_4904;
wire v_4906;
wire v_4907;
wire v_4908;
wire v_4909;
wire v_4910;
wire v_4911;
wire v_4912;
wire v_4913;
wire v_4914;
wire v_4915;
wire v_4916;
wire v_4917;
wire v_4918;
wire v_4920;
wire v_4921;
wire v_4923;
wire v_4924;
wire v_4927;
wire v_4929;
wire v_4932;
wire v_4933;
wire v_4934;
wire v_4935;
wire v_4937;
wire v_4939;
wire v_4942;
wire v_4944;
wire v_4945;
wire v_4947;
wire v_4949;
wire v_4950;
wire v_4952;
wire v_4953;
wire v_4954;
wire v_4955;
wire v_4957;
wire v_4958;
wire v_4959;
wire v_4960;
wire v_4964;
wire v_4965;
wire v_4966;
wire v_4968;
wire v_4970;
wire v_4972;
wire v_4973;
wire v_4974;
wire v_4976;
wire v_4977;
wire v_4978;
wire v_4981;
wire v_4984;
wire v_4986;
wire v_4988;
wire v_4990;
wire v_4992;
wire v_4993;
wire v_4996;
wire v_4997;
wire v_4999;
wire v_5000;
wire v_5001;
wire v_5004;
wire v_5005;
wire v_5006;
wire v_5008;
wire v_5010;
wire v_5012;
wire v_5013;
wire v_5014;
wire v_5017;
wire v_5018;
wire v_5019;
wire v_5021;
wire v_5023;
wire v_5025;
wire v_5026;
wire v_5027;
wire v_5029;
wire v_5030;
wire v_5033;
wire v_5034;
wire v_5035;
wire v_5037;
wire v_5039;
wire v_5041;
wire v_5042;
wire v_5043;
wire v_5045;
wire v_5046;
wire v_5047;
wire v_5049;
wire v_5050;
wire v_5051;
wire v_5052;
wire v_5053;
wire v_5057;
wire v_5058;
wire v_5059;
wire v_5061;
wire v_5062;
wire v_5063;
wire v_5064;
wire v_5065;
wire v_5066;
wire v_5067;
wire v_5068;
wire v_5069;
wire v_5070;
wire v_5071;
wire v_5072;
wire v_5073;
wire v_5074;
wire v_5075;
wire v_5076;
wire v_5077;
wire v_5078;
wire v_5079;
wire v_5080;
wire v_5081;
wire v_5082;
wire v_5083;
wire v_5084;
wire v_5085;
wire v_5086;
wire v_5087;
wire v_5088;
wire v_5089;
wire v_5090;
wire v_5091;
wire v_5092;
wire v_5093;
wire v_5094;
wire v_5095;
wire v_5096;
wire v_5097;
wire v_5098;
wire v_5099;
wire v_5100;
wire v_5101;
wire v_5102;
wire v_5103;
wire v_5104;
wire v_5105;
wire v_5106;
wire v_5107;
wire v_5108;
wire v_5109;
wire v_5110;
wire v_5111;
wire v_5112;
wire v_5113;
wire v_5114;
wire v_5115;
wire v_5116;
wire v_5117;
wire v_5118;
wire v_5119;
wire v_5120;
wire v_5121;
wire v_5122;
wire v_5123;
wire v_5124;
wire v_5125;
wire v_5126;
wire v_5127;
wire v_5128;
wire v_5129;
wire v_5130;
wire v_5131;
wire v_5132;
wire v_5133;
wire v_5134;
wire v_5135;
wire v_5136;
wire v_5137;
wire v_5138;
wire v_5139;
wire v_5140;
wire v_5141;
wire v_5142;
wire v_5143;
wire v_5144;
wire v_5145;
wire v_5146;
wire v_5147;
wire v_5148;
wire v_5149;
wire v_5150;
wire v_5151;
wire v_5152;
wire v_5153;
wire v_5154;
wire v_5155;
wire v_5156;
wire v_5157;
wire v_5158;
wire v_5159;
wire v_5160;
wire v_5161;
wire v_5162;
wire v_5163;
wire v_5164;
wire v_5165;
wire v_5166;
wire v_5167;
wire v_5168;
wire v_5169;
wire v_5170;
wire v_5171;
wire v_5172;
wire v_5173;
wire v_5174;
wire v_5175;
wire v_5176;
wire v_5177;
wire v_5178;
wire v_5179;
wire v_5180;
wire v_5183;
wire v_5184;
wire v_5185;
wire v_5186;
wire v_5187;
wire v_5188;
wire v_5189;
wire v_5190;
wire v_5191;
wire v_5192;
wire v_5193;
wire v_5194;
wire v_5195;
wire v_5196;
wire v_5197;
wire v_5198;
wire v_5199;
wire v_5200;
wire v_5201;
wire v_5202;
wire v_5203;
wire v_5204;
wire v_5205;
wire v_5206;
wire v_5207;
wire v_5208;
wire v_5209;
wire v_5210;
wire v_5211;
wire v_5212;
wire v_5213;
wire v_5214;
wire v_5215;
wire v_5216;
wire v_5217;
wire v_5218;
wire v_5219;
wire v_5220;
wire v_5221;
wire v_5222;
wire v_5223;
wire v_5224;
wire v_5225;
wire v_5226;
wire v_5227;
wire v_5228;
wire v_5229;
wire v_5230;
wire v_5231;
wire v_5232;
wire v_5233;
wire v_5234;
wire v_5235;
wire v_5236;
wire v_5237;
wire v_5238;
wire v_5239;
wire v_5240;
wire v_5241;
wire v_5242;
wire v_5243;
wire v_5244;
wire v_5245;
wire v_5246;
wire v_5247;
wire v_5248;
wire v_5249;
wire v_5250;
wire v_5251;
wire v_5252;
wire v_5253;
wire v_5254;
wire v_5255;
wire v_5256;
wire v_5257;
wire v_5258;
wire v_5259;
wire v_5260;
wire v_5261;
wire v_5262;
wire v_5263;
wire v_5264;
wire v_5265;
wire v_5266;
wire v_5267;
wire v_5268;
wire v_5269;
wire v_5270;
wire v_5271;
wire v_5272;
wire v_5273;
wire v_5274;
wire v_5275;
wire v_5276;
wire v_5277;
wire v_5278;
wire v_5279;
wire v_5280;
wire v_5281;
wire v_5282;
wire v_5283;
wire v_5284;
wire v_5285;
wire v_5286;
wire v_5287;
wire v_5288;
wire v_5289;
wire v_5290;
wire v_5291;
wire v_5292;
wire v_5293;
wire v_5295;
wire v_5296;
wire v_5297;
wire v_5299;
wire v_5300;
wire v_5301;
wire v_5302;
wire v_5303;
wire v_5304;
wire v_5305;
wire v_5306;
wire v_5307;
wire v_5308;
wire v_5309;
wire v_5310;
wire v_5311;
wire v_5312;
wire v_5313;
wire v_5314;
wire v_5315;
wire v_5316;
wire v_5317;
wire v_5318;
wire v_5319;
wire v_5320;
wire v_5321;
wire v_5322;
wire v_5323;
wire v_5324;
wire v_5325;
wire v_5326;
wire v_5327;
wire v_5328;
wire v_5329;
wire v_5330;
wire v_5331;
wire v_5332;
wire v_5333;
wire v_5334;
wire v_5335;
wire v_5336;
wire v_5337;
wire v_5338;
wire v_5339;
wire v_5340;
wire v_5341;
wire v_5342;
wire v_5343;
wire v_5344;
wire v_5345;
wire v_5346;
wire v_5347;
wire v_5348;
wire v_5349;
wire v_5350;
wire v_5351;
wire v_5352;
wire v_5353;
wire v_5354;
wire v_5355;
wire v_5356;
wire v_5357;
wire v_5358;
wire v_5359;
wire v_5360;
wire v_5361;
wire v_5362;
wire v_5363;
wire v_5364;
wire v_5365;
wire v_5366;
wire v_5367;
wire v_5368;
wire v_5369;
wire v_5370;
wire v_5371;
wire v_5372;
wire v_5373;
wire v_5374;
wire v_5375;
wire v_5376;
wire v_5377;
wire v_5378;
wire v_5379;
wire v_5380;
wire v_5381;
wire v_5382;
wire v_5383;
wire v_5384;
wire v_5385;
wire v_5386;
wire v_5387;
wire v_5388;
wire v_5389;
wire v_5390;
wire v_5391;
wire v_5392;
wire v_5393;
wire v_5395;
wire v_5396;
wire v_5397;
wire v_5398;
wire v_5399;
wire v_5400;
wire v_5401;
wire v_5402;
wire v_5403;
wire v_5404;
wire v_5405;
wire v_5406;
wire v_5407;
wire v_5408;
wire v_5409;
wire v_5410;
wire v_5411;
wire v_5412;
wire v_5413;
wire v_5414;
wire v_5415;
wire v_5416;
wire v_5417;
wire v_5418;
wire v_5419;
wire v_5420;
wire v_5421;
wire v_5422;
wire v_5423;
wire v_5424;
wire v_5425;
wire v_5426;
wire v_5427;
wire v_5428;
wire v_5429;
wire v_5430;
wire v_5431;
wire v_5432;
wire v_5433;
wire v_5434;
wire v_5435;
wire v_5436;
wire v_5437;
wire v_5438;
wire v_5439;
wire v_5440;
wire v_5441;
wire v_5442;
wire v_5443;
wire v_5444;
wire v_5445;
wire v_5446;
wire v_5447;
wire v_5448;
wire v_5449;
wire v_5450;
wire v_5451;
wire v_5452;
wire v_5453;
wire v_5454;
wire v_5455;
wire v_5456;
wire v_5457;
wire v_5458;
wire v_5459;
wire v_5460;
wire v_5461;
wire v_5462;
wire v_5463;
wire v_5464;
wire v_5465;
wire v_5466;
wire v_5467;
wire v_5468;
wire v_5469;
wire v_5470;
wire v_5471;
wire v_5472;
wire v_5473;
wire v_5474;
wire v_5475;
wire v_5476;
wire v_5477;
wire v_5478;
wire v_5479;
wire v_5480;
wire v_5481;
wire v_5482;
wire v_5483;
wire v_5484;
wire v_5485;
wire v_5486;
wire v_5487;
wire v_5488;
wire v_5489;
wire v_5490;
wire v_5491;
wire v_5492;
wire v_5493;
wire v_5494;
wire v_5495;
wire v_5496;
wire v_5497;
wire v_5498;
wire v_5499;
wire v_5500;
wire v_5501;
wire v_5502;
wire v_5503;
wire v_5504;
wire v_5505;
wire v_5506;
wire v_5507;
wire v_5508;
wire v_5509;
wire v_5510;
wire v_5511;
wire v_5512;
wire v_5513;
wire v_5514;
wire v_5515;
wire v_5516;
wire v_5517;
wire v_5518;
wire v_5519;
wire v_5520;
wire v_5521;
wire v_5522;
wire v_5523;
wire v_5524;
wire v_5525;
wire v_5526;
wire v_5527;
wire v_5528;
wire v_5529;
wire v_5530;
wire v_5531;
wire v_5532;
wire v_5533;
wire v_5534;
wire v_5535;
wire v_5536;
wire v_5537;
wire v_5538;
wire v_5539;
wire v_5540;
wire v_5541;
wire v_5542;
wire v_5543;
wire v_5544;
wire v_5545;
wire v_5546;
wire v_5547;
wire v_5548;
wire v_5549;
wire v_5550;
wire v_5551;
wire v_5552;
wire v_5553;
wire v_5554;
wire v_5555;
wire v_5556;
wire v_5557;
wire v_5558;
wire v_5559;
wire v_5560;
wire v_5561;
wire v_5562;
wire v_5563;
wire v_5564;
wire v_5565;
wire v_5566;
wire v_5567;
wire v_5568;
wire v_5569;
wire v_5570;
wire v_5571;
wire v_5572;
wire v_5573;
wire v_5574;
wire v_5575;
wire v_5576;
wire v_5577;
wire v_5578;
wire v_5579;
wire v_5580;
wire v_5581;
wire v_5582;
wire v_5583;
wire v_5584;
wire v_5585;
wire v_5586;
wire v_5587;
wire v_5588;
wire v_5589;
wire v_5590;
wire v_5591;
wire v_5592;
wire v_5593;
wire v_5594;
wire v_5595;
wire v_5596;
wire v_5597;
wire v_5598;
wire v_5599;
wire v_5600;
wire v_5601;
wire v_5602;
wire v_5603;
wire v_5604;
wire v_5606;
wire v_5607;
wire v_5608;
wire v_5609;
wire v_5610;
wire v_5611;
wire v_5612;
wire v_5613;
wire v_5614;
wire v_5615;
wire v_5616;
wire v_5617;
wire v_5618;
wire v_5619;
wire v_5620;
wire v_5621;
wire v_5622;
wire v_5623;
wire v_5624;
wire v_5626;
wire v_5627;
wire v_5628;
wire v_5629;
wire v_5630;
wire v_5631;
wire v_5632;
wire v_5633;
wire v_5634;
wire v_5635;
wire v_5636;
wire v_5637;
wire v_5638;
wire v_5639;
wire v_5640;
wire v_5641;
wire v_5642;
wire v_5643;
wire v_5644;
wire v_5645;
wire v_5646;
wire v_5647;
wire v_5648;
wire v_5649;
wire v_5650;
wire v_5651;
wire v_5652;
wire v_5653;
wire v_5654;
wire v_5655;
wire v_5656;
wire v_5657;
wire v_5658;
wire v_5659;
wire v_5660;
wire v_5661;
wire v_5662;
wire v_5663;
wire v_5664;
wire v_5665;
wire v_5666;
wire v_5667;
wire v_5668;
wire v_5669;
wire v_5670;
wire v_5671;
wire v_5672;
wire v_5673;
wire v_5674;
wire v_5675;
wire v_5677;
wire v_5678;
wire v_5679;
wire v_5680;
wire v_5681;
wire v_5682;
wire v_5683;
wire v_5684;
wire v_5685;
wire v_5686;
wire v_5687;
wire v_5688;
wire v_5689;
wire v_5690;
wire v_5691;
wire v_5692;
wire v_5693;
wire v_5695;
wire v_5696;
wire v_5697;
wire v_5698;
wire v_5699;
wire v_5700;
wire v_5701;
wire v_5702;
wire v_5703;
wire v_5704;
wire v_5705;
wire v_5706;
wire v_5707;
wire v_5708;
wire v_5709;
wire v_5710;
wire v_5711;
wire v_5712;
wire v_5713;
wire v_5714;
wire v_5715;
wire v_5716;
wire v_5717;
wire v_5718;
wire v_5719;
wire v_5720;
wire v_5721;
wire v_5722;
wire v_5723;
wire v_5724;
wire v_5725;
wire v_5726;
wire v_5727;
wire v_5728;
wire v_5729;
wire v_5730;
wire v_5731;
wire v_5732;
wire v_5733;
wire v_5734;
wire v_5735;
wire v_5736;
wire v_5737;
wire v_5738;
wire v_5739;
wire v_5740;
wire v_5741;
wire v_5742;
wire v_5743;
wire v_5744;
wire v_5745;
wire v_5746;
wire v_5747;
wire v_5748;
wire v_5749;
wire v_5750;
wire v_5751;
wire v_5752;
wire v_5753;
wire v_5754;
wire v_5755;
wire v_5756;
wire v_5757;
wire v_5758;
wire v_5759;
wire v_5760;
wire v_5761;
wire v_5762;
wire v_5763;
wire v_5764;
wire v_5765;
wire v_5766;
wire v_5767;
wire v_5768;
wire v_5769;
wire v_5770;
wire v_5771;
wire v_5772;
wire v_5773;
wire v_5774;
wire v_5775;
wire v_5776;
wire v_5777;
wire v_5778;
wire v_5779;
wire v_5780;
wire v_5781;
wire v_5782;
wire v_5783;
wire v_5784;
wire v_5785;
wire v_5786;
wire v_5787;
wire v_5788;
wire v_5789;
wire v_5790;
wire v_5791;
wire v_5792;
wire v_5793;
wire v_5794;
wire v_5795;
wire v_5796;
wire v_5797;
wire v_5798;
wire v_5799;
wire v_5800;
wire v_5801;
wire v_5802;
wire v_5803;
wire v_5804;
wire v_5805;
wire v_5806;
wire v_5807;
wire v_5808;
wire v_5809;
wire v_5810;
wire v_5811;
wire v_5812;
wire v_5813;
wire v_5814;
wire v_5815;
wire v_5816;
wire v_5817;
wire v_5818;
wire v_5819;
wire v_5820;
wire v_5821;
wire v_5822;
wire v_5824;
wire v_5825;
wire v_5826;
wire v_5827;
wire v_5828;
wire v_5829;
wire v_5830;
wire v_5831;
wire v_5832;
wire v_5833;
wire v_5834;
wire v_5835;
wire v_5836;
wire v_5837;
wire v_5838;
wire v_5839;
wire v_5840;
wire v_5841;
wire v_5842;
wire v_5844;
wire v_5845;
wire v_5846;
wire v_5847;
wire v_5848;
wire v_5849;
wire v_5850;
wire v_5851;
wire v_5852;
wire v_5853;
wire v_5854;
wire v_5855;
wire v_5856;
wire v_5857;
wire v_5858;
wire v_5859;
wire v_5860;
wire v_5861;
wire v_5862;
wire v_5863;
wire v_5864;
wire v_5865;
wire v_5866;
wire v_5867;
wire v_5868;
wire v_5869;
wire v_5870;
wire v_5871;
wire v_5872;
wire v_5873;
wire v_5874;
wire v_5875;
wire v_5876;
wire v_5877;
wire v_5878;
wire v_5879;
wire v_5880;
wire v_5881;
wire v_5882;
wire v_5883;
wire v_5884;
wire v_5885;
wire v_5886;
wire v_5887;
wire v_5888;
wire v_5889;
wire v_5890;
wire v_5891;
wire v_5892;
wire v_5893;
wire v_5895;
wire v_5896;
wire v_5897;
wire v_5898;
wire v_5899;
wire v_5900;
wire v_5901;
wire v_5902;
wire v_5903;
wire v_5904;
wire v_5905;
wire v_5906;
wire v_5907;
wire v_5908;
wire v_5909;
wire v_5910;
wire v_5911;
wire v_5913;
wire v_5914;
wire v_5915;
wire v_5916;
wire v_5917;
wire v_5918;
wire v_5920;
wire v_5921;
wire v_5922;
wire v_5923;
wire v_5924;
wire v_5925;
wire v_5926;
wire v_5927;
wire v_5928;
wire v_5929;
wire v_5930;
wire v_5931;
wire v_5932;
wire v_5933;
wire v_5934;
wire v_5935;
wire v_5936;
wire v_5937;
wire v_5938;
wire v_5939;
wire v_5940;
wire v_5941;
wire v_5942;
wire v_5943;
wire v_5944;
wire v_5945;
wire v_5946;
wire v_5947;
wire v_5948;
wire v_5949;
wire v_5950;
wire v_5951;
wire v_5952;
wire v_5953;
wire v_5954;
wire v_5955;
wire v_5956;
wire v_5957;
wire v_5958;
wire v_5959;
wire v_5960;
wire v_5961;
wire v_5962;
wire v_5963;
wire v_5964;
wire v_5965;
wire v_5966;
wire v_5967;
wire v_5968;
wire v_5969;
wire v_5970;
wire v_5971;
wire v_5972;
wire v_5973;
wire v_5974;
wire v_5975;
wire v_5976;
wire v_5977;
wire v_5978;
wire v_5979;
wire v_5980;
wire v_5981;
wire v_5982;
wire v_5983;
wire v_5984;
wire v_5985;
wire v_5986;
wire v_5987;
wire v_5988;
wire v_5989;
wire v_5990;
wire v_5991;
wire v_5992;
wire v_5993;
wire v_5994;
wire v_5995;
wire v_5996;
wire v_5997;
wire v_5998;
wire v_5999;
wire v_6000;
wire v_6001;
wire v_6002;
wire v_6003;
wire v_6004;
wire v_6005;
wire v_6006;
wire v_6007;
wire v_6008;
wire v_6009;
wire v_6010;
wire v_6011;
wire v_6012;
wire v_6013;
wire v_6014;
wire v_6015;
wire v_6016;
wire v_6017;
wire v_6018;
wire v_6019;
wire v_6020;
wire v_6021;
wire v_6022;
wire v_6023;
wire v_6024;
wire v_6025;
wire v_6026;
wire v_6027;
wire v_6028;
wire v_6029;
wire v_6030;
wire v_6031;
wire v_6032;
wire v_6033;
wire v_6034;
wire v_6035;
wire v_6036;
wire v_6037;
wire v_6038;
wire v_6039;
wire v_6040;
wire v_6041;
wire v_6042;
wire v_6043;
wire v_6045;
wire v_6046;
wire v_6047;
wire v_6048;
wire v_6049;
wire v_6050;
wire v_6051;
wire v_6052;
wire v_6053;
wire v_6054;
wire v_6055;
wire v_6056;
wire v_6057;
wire v_6058;
wire v_6059;
wire v_6060;
wire v_6061;
wire v_6062;
wire v_6063;
wire v_6065;
wire v_6066;
wire v_6067;
wire v_6068;
wire v_6069;
wire v_6070;
wire v_6071;
wire v_6072;
wire v_6073;
wire v_6074;
wire v_6075;
wire v_6076;
wire v_6077;
wire v_6078;
wire v_6079;
wire v_6080;
wire v_6081;
wire v_6082;
wire v_6083;
wire v_6084;
wire v_6085;
wire v_6086;
wire v_6087;
wire v_6088;
wire v_6089;
wire v_6090;
wire v_6091;
wire v_6092;
wire v_6093;
wire v_6094;
wire v_6095;
wire v_6096;
wire v_6097;
wire v_6098;
wire v_6099;
wire v_6100;
wire v_6101;
wire v_6102;
wire v_6103;
wire v_6104;
wire v_6105;
wire v_6106;
wire v_6107;
wire v_6108;
wire v_6109;
wire v_6110;
wire v_6111;
wire v_6112;
wire v_6113;
wire v_6114;
wire v_6116;
wire v_6117;
wire v_6118;
wire v_6119;
wire v_6120;
wire v_6121;
wire v_6122;
wire v_6123;
wire v_6124;
wire v_6125;
wire v_6126;
wire v_6127;
wire v_6128;
wire v_6129;
wire v_6130;
wire v_6131;
wire v_6132;
wire v_6134;
wire v_6135;
wire v_6136;
wire v_6137;
wire v_6138;
wire v_6139;
wire v_6141;
wire v_6142;
wire v_6143;
wire v_6144;
wire v_6145;
wire v_6146;
wire v_6147;
wire v_6148;
wire v_6149;
wire v_6150;
wire v_6151;
wire v_6152;
wire v_6153;
wire v_6154;
wire v_6155;
wire v_6156;
wire v_6157;
wire v_6158;
wire v_6159;
wire v_6160;
wire v_6161;
wire v_6162;
wire v_6163;
wire v_6164;
wire v_6165;
wire v_6166;
wire v_6167;
wire v_6168;
wire v_6169;
wire v_6170;
wire v_6171;
wire v_6172;
wire v_6173;
wire v_6174;
wire v_6175;
wire v_6176;
wire v_6177;
wire v_6178;
wire v_6179;
wire v_6180;
wire v_6181;
wire v_6182;
wire v_6183;
wire v_6184;
wire v_6185;
wire v_6186;
wire v_6187;
wire v_6188;
wire v_6189;
wire v_6190;
wire v_6191;
wire v_6192;
wire v_6193;
wire v_6194;
wire v_6195;
wire v_6196;
wire v_6197;
wire v_6198;
wire v_6199;
wire v_6200;
wire v_6201;
wire v_6202;
wire v_6203;
wire v_6204;
wire v_6205;
wire v_6206;
wire v_6207;
wire v_6208;
wire v_6209;
wire v_6210;
wire v_6211;
wire v_6212;
wire v_6213;
wire v_6214;
wire v_6215;
wire v_6216;
wire v_6217;
wire v_6218;
wire v_6219;
wire v_6220;
wire v_6221;
wire v_6222;
wire v_6223;
wire v_6224;
wire v_6225;
wire v_6226;
wire v_6227;
wire v_6228;
wire v_6229;
wire v_6230;
wire v_6231;
wire v_6232;
wire v_6233;
wire v_6234;
wire v_6235;
wire v_6236;
wire v_6237;
wire v_6238;
wire v_6239;
wire v_6240;
wire v_6241;
wire v_6242;
wire v_6243;
wire v_6244;
wire v_6245;
wire v_6246;
wire v_6247;
wire v_6248;
wire v_6249;
wire v_6250;
wire v_6251;
wire v_6252;
wire v_6253;
wire v_6254;
wire v_6255;
wire v_6256;
wire v_6257;
wire v_6258;
wire v_6259;
wire v_6260;
wire v_6261;
wire v_6262;
wire v_6263;
wire v_6264;
wire v_6266;
wire v_6267;
wire v_6268;
wire v_6269;
wire v_6270;
wire v_6271;
wire v_6272;
wire v_6273;
wire v_6274;
wire v_6275;
wire v_6276;
wire v_6277;
wire v_6278;
wire v_6279;
wire v_6280;
wire v_6281;
wire v_6282;
wire v_6283;
wire v_6284;
wire v_6286;
wire v_6287;
wire v_6288;
wire v_6289;
wire v_6290;
wire v_6291;
wire v_6292;
wire v_6293;
wire v_6294;
wire v_6295;
wire v_6296;
wire v_6297;
wire v_6298;
wire v_6299;
wire v_6300;
wire v_6301;
wire v_6302;
wire v_6303;
wire v_6304;
wire v_6305;
wire v_6306;
wire v_6307;
wire v_6308;
wire v_6309;
wire v_6310;
wire v_6311;
wire v_6312;
wire v_6313;
wire v_6314;
wire v_6315;
wire v_6316;
wire v_6317;
wire v_6318;
wire v_6319;
wire v_6320;
wire v_6321;
wire v_6322;
wire v_6323;
wire v_6324;
wire v_6325;
wire v_6326;
wire v_6327;
wire v_6328;
wire v_6329;
wire v_6330;
wire v_6331;
wire v_6332;
wire v_6333;
wire v_6334;
wire v_6335;
wire v_6337;
wire v_6338;
wire v_6339;
wire v_6340;
wire v_6341;
wire v_6342;
wire v_6343;
wire v_6344;
wire v_6345;
wire v_6346;
wire v_6347;
wire v_6348;
wire v_6349;
wire v_6350;
wire v_6351;
wire v_6352;
wire v_6353;
wire v_6355;
wire v_6356;
wire v_6357;
wire v_6358;
wire v_6359;
wire v_6360;
wire v_6361;
wire v_6362;
wire v_6363;
wire v_6364;
wire v_6365;
wire v_6366;
wire v_6367;
wire v_6368;
wire v_6369;
wire v_6370;
wire v_6371;
wire v_6372;
wire v_6373;
wire v_6374;
wire v_6375;
wire v_6376;
wire v_6377;
wire v_6378;
wire v_6379;
wire v_6380;
wire v_6381;
wire v_6382;
wire v_6383;
wire v_6384;
wire v_6385;
wire v_6386;
wire v_6387;
wire v_6388;
wire v_6389;
wire v_6390;
wire v_6391;
wire v_6392;
wire v_6393;
wire v_6394;
wire v_6395;
wire v_6396;
wire v_6397;
wire v_6398;
wire v_6399;
wire v_6400;
wire v_6401;
wire v_6402;
wire v_6403;
wire v_6404;
wire v_6405;
wire v_6406;
wire v_6407;
wire v_6408;
wire v_6409;
wire v_6410;
wire v_6411;
wire v_6412;
wire v_6413;
wire v_6414;
wire v_6415;
wire v_6416;
wire v_6417;
wire v_6418;
wire v_6419;
wire v_6420;
wire v_6421;
wire v_6422;
wire v_6423;
wire v_6424;
wire v_6425;
wire v_6426;
wire v_6427;
wire v_6428;
wire v_6429;
wire v_6430;
wire v_6431;
wire v_6432;
wire v_6433;
wire v_6434;
wire v_6435;
wire v_6436;
wire v_6437;
wire v_6438;
wire v_6439;
wire v_6440;
wire v_6441;
wire v_6442;
wire v_6443;
wire v_6444;
wire v_6445;
wire v_6446;
wire v_6447;
wire v_6448;
wire v_6449;
wire v_6450;
wire v_6451;
wire v_6452;
wire v_6453;
wire v_6454;
wire v_6455;
wire v_6456;
wire v_6457;
wire v_6458;
wire v_6459;
wire v_6460;
wire v_6461;
wire v_6462;
wire v_6463;
wire v_6464;
wire v_6465;
wire v_6466;
wire v_6467;
wire v_6468;
wire v_6469;
wire v_6470;
wire v_6471;
wire v_6472;
wire v_6473;
wire v_6474;
wire v_6475;
wire v_6476;
wire v_6477;
wire v_6478;
wire v_6479;
wire v_6480;
wire v_6481;
wire v_6482;
wire v_6483;
wire v_6484;
wire v_6486;
wire v_6487;
wire v_6488;
wire v_6489;
wire v_6490;
wire v_6491;
wire v_6492;
wire v_6493;
wire v_6494;
wire v_6495;
wire v_6496;
wire v_6497;
wire v_6498;
wire v_6499;
wire v_6500;
wire v_6501;
wire v_6502;
wire v_6503;
wire v_6504;
wire v_6506;
wire v_6507;
wire v_6508;
wire v_6509;
wire v_6510;
wire v_6511;
wire v_6512;
wire v_6513;
wire v_6514;
wire v_6515;
wire v_6516;
wire v_6517;
wire v_6518;
wire v_6519;
wire v_6520;
wire v_6521;
wire v_6522;
wire v_6523;
wire v_6524;
wire v_6525;
wire v_6526;
wire v_6527;
wire v_6528;
wire v_6529;
wire v_6530;
wire v_6531;
wire v_6532;
wire v_6533;
wire v_6534;
wire v_6535;
wire v_6536;
wire v_6537;
wire v_6538;
wire v_6539;
wire v_6540;
wire v_6541;
wire v_6542;
wire v_6543;
wire v_6544;
wire v_6545;
wire v_6546;
wire v_6547;
wire v_6548;
wire v_6549;
wire v_6550;
wire v_6551;
wire v_6552;
wire v_6553;
wire v_6554;
wire v_6555;
wire v_6557;
wire v_6558;
wire v_6559;
wire v_6560;
wire v_6561;
wire v_6562;
wire v_6563;
wire v_6564;
wire v_6565;
wire v_6566;
wire v_6567;
wire v_6568;
wire v_6569;
wire v_6570;
wire v_6571;
wire v_6572;
wire v_6573;
wire v_6575;
wire v_6576;
wire v_6577;
wire v_6578;
wire v_6579;
wire v_6580;
wire v_6582;
wire v_6583;
wire v_6584;
wire v_6585;
wire v_6586;
wire v_6587;
wire v_6588;
wire v_6589;
wire v_6590;
wire v_6591;
wire v_6592;
wire v_6593;
wire v_6594;
wire v_6595;
wire v_6596;
wire v_6597;
wire v_6598;
wire v_6599;
wire v_6600;
wire v_6601;
wire v_6602;
wire v_6603;
wire v_6604;
wire v_6605;
wire v_6606;
wire v_6607;
wire v_6608;
wire v_6609;
wire v_6610;
wire v_6611;
wire v_6612;
wire v_6613;
wire v_6614;
wire v_6615;
wire v_6616;
wire v_6617;
wire v_6618;
wire v_6619;
wire v_6620;
wire v_6621;
wire v_6622;
wire v_6623;
wire v_6624;
wire v_6625;
wire v_6626;
wire v_6627;
wire v_6628;
wire v_6629;
wire v_6630;
wire v_6631;
wire v_6632;
wire v_6633;
wire v_6634;
wire v_6635;
wire v_6636;
wire v_6637;
wire v_6638;
wire v_6639;
wire v_6640;
wire v_6641;
wire v_6642;
wire v_6643;
wire v_6644;
wire v_6645;
wire v_6646;
wire v_6647;
wire v_6648;
wire v_6649;
wire v_6650;
wire v_6651;
wire v_6652;
wire v_6653;
wire v_6654;
wire v_6655;
wire v_6656;
wire v_6657;
wire v_6658;
wire v_6659;
wire v_6660;
wire v_6661;
wire v_6662;
wire v_6663;
wire v_6664;
wire v_6665;
wire v_6666;
wire v_6667;
wire v_6668;
wire v_6669;
wire v_6670;
wire v_6671;
wire v_6672;
wire v_6673;
wire v_6674;
wire v_6675;
wire v_6676;
wire v_6677;
wire v_6678;
wire v_6679;
wire v_6680;
wire v_6681;
wire v_6682;
wire v_6683;
wire v_6684;
wire v_6685;
wire v_6686;
wire v_6687;
wire v_6688;
wire v_6689;
wire v_6690;
wire v_6691;
wire v_6692;
wire v_6693;
wire v_6694;
wire v_6695;
wire v_6696;
wire v_6697;
wire v_6698;
wire v_6699;
wire v_6700;
wire v_6701;
wire v_6702;
wire v_6703;
wire v_6704;
wire v_6705;
wire v_6707;
wire v_6708;
wire v_6709;
wire v_6710;
wire v_6711;
wire v_6712;
wire v_6713;
wire v_6714;
wire v_6715;
wire v_6716;
wire v_6717;
wire v_6718;
wire v_6719;
wire v_6720;
wire v_6721;
wire v_6722;
wire v_6723;
wire v_6724;
wire v_6725;
wire v_6727;
wire v_6728;
wire v_6729;
wire v_6730;
wire v_6731;
wire v_6732;
wire v_6733;
wire v_6734;
wire v_6735;
wire v_6736;
wire v_6737;
wire v_6738;
wire v_6739;
wire v_6740;
wire v_6741;
wire v_6742;
wire v_6743;
wire v_6744;
wire v_6745;
wire v_6746;
wire v_6747;
wire v_6748;
wire v_6749;
wire v_6750;
wire v_6751;
wire v_6752;
wire v_6753;
wire v_6754;
wire v_6755;
wire v_6756;
wire v_6757;
wire v_6758;
wire v_6759;
wire v_6760;
wire v_6761;
wire v_6762;
wire v_6763;
wire v_6764;
wire v_6765;
wire v_6766;
wire v_6767;
wire v_6768;
wire v_6769;
wire v_6770;
wire v_6771;
wire v_6772;
wire v_6773;
wire v_6774;
wire v_6775;
wire v_6776;
wire v_6778;
wire v_6779;
wire v_6780;
wire v_6781;
wire v_6782;
wire v_6783;
wire v_6784;
wire v_6785;
wire v_6786;
wire v_6787;
wire v_6788;
wire v_6789;
wire v_6790;
wire v_6791;
wire v_6792;
wire v_6793;
wire v_6794;
wire v_6796;
wire v_6797;
wire v_6798;
wire v_6799;
wire v_6800;
wire v_6801;
wire v_6803;
wire v_6804;
wire v_6805;
wire v_6806;
wire v_6808;
wire v_6809;
wire v_6810;
wire v_6811;
wire v_6812;
wire v_6813;
wire v_6814;
wire v_6815;
wire v_6816;
wire v_6817;
wire v_6818;
wire v_6819;
wire v_6820;
wire v_6821;
wire v_6822;
wire v_6823;
wire v_6824;
wire v_6825;
wire v_6826;
wire v_6827;
wire v_6828;
wire v_6829;
wire v_6830;
wire v_6831;
wire v_6832;
wire v_6833;
wire v_6834;
wire v_6835;
wire v_6836;
wire v_6837;
wire v_6838;
wire v_6839;
wire v_6840;
wire v_6841;
wire v_6842;
wire v_6843;
wire v_6844;
wire v_6845;
wire v_6846;
wire v_6847;
wire v_6848;
wire v_6849;
wire v_6850;
wire v_6851;
wire v_6852;
wire v_6853;
wire v_6854;
wire v_6855;
wire v_6856;
wire v_6857;
wire v_6858;
wire v_6859;
wire v_6860;
wire v_6861;
wire v_6862;
wire v_6863;
wire v_6864;
wire v_6865;
wire v_6866;
wire v_6867;
wire v_6868;
wire v_6869;
wire v_6870;
wire v_6871;
wire v_6872;
wire v_6873;
wire v_6874;
wire v_6875;
wire v_6876;
wire v_6877;
wire v_6878;
wire v_6879;
wire v_6880;
wire v_6881;
wire v_6882;
wire v_6883;
wire v_6884;
wire v_6885;
wire v_6886;
wire v_6887;
wire v_6888;
wire v_6889;
wire v_6890;
wire v_6891;
wire v_6892;
wire v_6893;
wire v_6894;
wire v_6895;
wire v_6896;
wire v_6897;
wire v_6898;
wire v_6899;
wire v_6900;
wire v_6901;
wire v_6903;
wire v_6904;
wire v_6905;
wire v_6906;
wire v_6907;
wire v_6908;
wire v_6909;
wire v_6910;
wire v_6911;
wire v_6912;
wire v_6913;
wire v_6914;
wire v_6915;
wire v_6916;
wire v_6917;
wire v_6918;
wire v_6919;
wire v_6920;
wire v_6921;
wire v_6922;
wire v_6923;
wire v_6924;
wire v_6925;
wire v_6926;
wire v_6927;
wire v_6928;
wire v_6929;
wire v_6930;
wire v_6931;
wire v_6932;
wire v_6933;
wire v_6934;
wire v_6935;
wire v_6936;
wire v_6937;
wire v_6938;
wire v_6939;
wire v_6940;
wire v_6941;
wire v_6942;
wire v_6943;
wire v_6944;
wire v_6945;
wire v_6946;
wire v_6947;
wire v_6948;
wire v_6949;
wire v_6950;
wire v_6951;
wire v_6952;
wire v_6953;
wire v_6954;
wire v_6955;
wire v_6956;
wire v_6957;
wire v_6958;
wire v_6959;
wire v_6960;
wire v_6961;
wire v_6962;
wire v_6963;
wire v_6964;
wire v_6965;
wire v_6966;
wire v_6967;
wire v_6968;
wire v_6969;
wire v_6970;
wire v_6971;
wire v_6972;
wire v_6973;
wire v_6974;
wire v_6975;
wire v_6976;
wire v_6977;
wire v_6978;
wire v_6979;
wire v_6980;
wire v_6981;
wire v_6982;
wire v_6983;
wire v_6984;
wire v_6985;
wire v_6986;
wire v_6987;
wire v_6989;
wire v_6990;
wire v_6991;
wire v_6992;
wire v_6993;
wire v_6994;
wire v_6995;
wire v_6996;
wire v_6997;
wire v_6998;
wire v_6999;
wire v_7000;
wire v_7001;
wire v_7002;
wire v_7003;
wire v_7004;
wire v_7005;
wire v_7006;
wire v_7007;
wire v_7008;
wire v_7009;
wire v_7010;
wire v_7011;
wire v_7012;
wire v_7013;
wire v_7014;
wire v_7015;
wire v_7016;
wire v_7017;
wire v_7018;
wire v_7019;
wire v_7020;
wire v_7021;
wire v_7022;
wire v_7023;
wire v_7024;
wire v_7025;
wire v_7026;
wire v_7027;
wire v_7028;
wire v_7029;
wire v_7030;
wire v_7031;
wire v_7032;
wire v_7033;
wire v_7034;
wire v_7035;
wire v_7036;
wire v_7037;
wire v_7038;
wire v_7039;
wire v_7040;
wire v_7041;
wire v_7042;
wire v_7043;
wire v_7044;
wire v_7045;
wire v_7046;
wire v_7047;
wire v_7048;
wire v_7049;
wire v_7050;
wire v_7051;
wire v_7052;
wire v_7053;
wire v_7054;
wire v_7055;
wire v_7056;
wire v_7057;
wire v_7058;
wire v_7059;
wire v_7060;
wire v_7061;
wire v_7062;
wire v_7063;
wire v_7064;
wire v_7065;
wire v_7066;
wire v_7067;
wire v_7068;
wire v_7069;
wire v_7070;
wire v_7071;
wire v_7072;
wire v_7073;
wire v_7074;
wire v_7075;
wire v_7076;
wire v_7077;
wire v_7078;
wire v_7079;
wire v_7080;
wire v_7081;
wire v_7082;
wire v_7083;
wire v_7084;
wire v_7085;
wire v_7086;
wire v_7087;
wire v_7088;
wire v_7089;
wire v_7090;
wire v_7091;
wire v_7092;
wire v_7093;
wire v_7094;
wire v_7095;
wire v_7096;
wire v_7097;
wire v_7098;
wire v_7099;
wire v_7100;
wire v_7101;
wire v_7102;
wire v_7103;
wire v_7104;
wire v_7105;
wire v_7106;
wire v_7107;
wire v_7108;
wire v_7109;
wire v_7110;
wire v_7111;
wire v_7112;
wire v_7114;
wire v_7115;
wire v_7116;
wire v_7117;
wire v_7118;
wire v_7119;
wire v_7120;
wire v_7121;
wire v_7122;
wire v_7123;
wire v_7124;
wire v_7125;
wire v_7126;
wire v_7127;
wire v_7128;
wire v_7129;
wire v_7130;
wire v_7131;
wire v_7132;
wire v_7134;
wire v_7135;
wire v_7136;
wire v_7137;
wire v_7138;
wire v_7139;
wire v_7140;
wire v_7141;
wire v_7142;
wire v_7143;
wire v_7144;
wire v_7145;
wire v_7146;
wire v_7147;
wire v_7148;
wire v_7149;
wire v_7150;
wire v_7151;
wire v_7152;
wire v_7153;
wire v_7154;
wire v_7155;
wire v_7156;
wire v_7157;
wire v_7158;
wire v_7159;
wire v_7160;
wire v_7161;
wire v_7162;
wire v_7163;
wire v_7164;
wire v_7165;
wire v_7166;
wire v_7167;
wire v_7168;
wire v_7169;
wire v_7170;
wire v_7171;
wire v_7172;
wire v_7173;
wire v_7174;
wire v_7175;
wire v_7176;
wire v_7177;
wire v_7178;
wire v_7179;
wire v_7180;
wire v_7181;
wire v_7182;
wire v_7183;
wire v_7185;
wire v_7186;
wire v_7187;
wire v_7188;
wire v_7189;
wire v_7190;
wire v_7191;
wire v_7192;
wire v_7193;
wire v_7194;
wire v_7195;
wire v_7196;
wire v_7197;
wire v_7198;
wire v_7199;
wire v_7200;
wire v_7201;
wire v_7203;
wire v_7204;
wire v_7205;
wire v_7206;
wire v_7207;
wire v_7208;
wire v_7209;
wire v_7210;
wire v_7211;
wire v_7212;
wire v_7213;
wire v_7214;
wire v_7215;
wire v_7216;
wire v_7217;
wire v_7218;
wire v_7219;
wire v_7220;
wire v_7221;
wire v_7222;
wire v_7223;
wire v_7224;
wire v_7225;
wire v_7226;
wire v_7227;
wire v_7228;
wire v_7229;
wire v_7230;
wire v_7231;
wire v_7232;
wire v_7233;
wire v_7234;
wire v_7235;
wire v_7236;
wire v_7237;
wire v_7238;
wire v_7239;
wire v_7240;
wire v_7241;
wire v_7242;
wire v_7243;
wire v_7244;
wire v_7245;
wire v_7246;
wire v_7247;
wire v_7248;
wire v_7249;
wire v_7250;
wire v_7251;
wire v_7252;
wire v_7253;
wire v_7254;
wire v_7255;
wire v_7256;
wire v_7257;
wire v_7258;
wire v_7259;
wire v_7260;
wire v_7261;
wire v_7262;
wire v_7263;
wire v_7264;
wire v_7265;
wire v_7266;
wire v_7267;
wire v_7268;
wire v_7269;
wire v_7270;
wire v_7271;
wire v_7272;
wire v_7273;
wire v_7274;
wire v_7275;
wire v_7276;
wire v_7277;
wire v_7278;
wire v_7279;
wire v_7280;
wire v_7281;
wire v_7282;
wire v_7283;
wire v_7284;
wire v_7285;
wire v_7286;
wire v_7287;
wire v_7288;
wire v_7289;
wire v_7290;
wire v_7291;
wire v_7292;
wire v_7293;
wire v_7294;
wire v_7295;
wire v_7296;
wire v_7297;
wire v_7298;
wire v_7299;
wire v_7300;
wire v_7301;
wire v_7302;
wire v_7303;
wire v_7304;
wire v_7305;
wire v_7306;
wire v_7307;
wire v_7308;
wire v_7309;
wire v_7310;
wire v_7311;
wire v_7312;
wire v_7313;
wire v_7314;
wire v_7315;
wire v_7316;
wire v_7317;
wire v_7318;
wire v_7319;
wire v_7320;
wire v_7321;
wire v_7322;
wire v_7323;
wire v_7324;
wire v_7325;
wire v_7326;
wire v_7327;
wire v_7328;
wire v_7329;
wire v_7330;
wire v_7331;
wire v_7332;
wire v_7333;
wire v_7334;
wire v_7335;
wire v_7336;
wire v_7337;
wire v_7338;
wire v_7339;
wire v_7340;
wire v_7341;
wire v_7342;
wire v_7343;
wire v_7344;
wire v_7345;
wire v_7346;
wire v_7347;
wire v_7348;
wire v_7349;
wire v_7350;
wire v_7351;
wire v_7352;
wire v_7353;
wire v_7354;
wire v_7355;
wire v_7356;
wire v_7357;
wire v_7358;
wire v_7359;
wire v_7360;
wire v_7361;
wire v_7362;
wire v_7363;
wire v_7364;
wire v_7365;
wire v_7366;
wire v_7367;
wire v_7368;
wire v_7369;
wire v_7370;
wire v_7371;
wire v_7372;
wire v_7373;
wire v_7374;
wire v_7375;
wire v_7376;
wire v_7377;
wire v_7378;
wire v_7379;
wire v_7380;
wire v_7381;
wire v_7382;
wire v_7383;
wire v_7384;
wire v_7385;
wire v_7386;
wire v_7387;
wire v_7388;
wire v_7389;
wire v_7390;
wire v_7391;
wire v_7392;
wire v_7393;
wire v_7394;
wire v_7395;
wire v_7396;
wire v_7397;
wire v_7398;
wire v_7399;
wire v_7400;
wire v_7401;
wire v_7402;
wire v_7403;
wire v_7404;
wire v_7405;
wire v_7406;
wire v_7407;
wire v_7408;
wire v_7409;
wire v_7410;
wire v_7411;
wire v_7412;
wire v_7413;
wire v_7414;
wire v_7415;
wire v_7416;
wire v_7417;
wire v_7418;
wire v_7419;
wire v_7420;
wire v_7421;
wire v_7422;
wire v_7423;
wire v_7424;
wire v_7425;
wire v_7426;
wire v_7427;
wire v_7428;
wire v_7429;
wire v_7430;
wire v_7431;
wire v_7432;
wire v_7433;
wire v_7434;
wire v_7435;
wire v_7436;
wire v_7437;
wire v_7438;
wire v_7439;
wire v_7440;
wire v_7441;
wire v_7442;
wire v_7443;
wire v_7444;
wire v_7445;
wire v_7446;
wire v_7447;
wire v_7448;
wire v_7449;
wire v_7450;
wire v_7451;
wire v_7452;
wire v_7453;
wire v_7454;
wire v_7455;
wire v_7456;
wire v_7457;
wire v_7458;
wire v_7459;
wire v_7460;
wire v_7461;
wire v_7462;
wire v_7463;
wire v_7464;
wire v_7465;
wire v_7466;
wire v_7467;
wire v_7468;
wire v_7469;
wire v_7470;
wire v_7471;
wire v_7472;
wire v_7473;
wire v_7474;
wire v_7475;
wire v_7476;
wire v_7477;
wire v_7478;
wire v_7479;
wire v_7480;
wire v_7481;
wire v_7482;
wire v_7483;
wire v_7484;
wire v_7485;
wire v_7486;
wire v_7487;
wire v_7488;
wire v_7489;
wire v_7490;
wire v_7491;
wire v_7492;
wire v_7493;
wire v_7494;
wire v_7495;
wire v_7496;
wire v_7497;
wire v_7498;
wire v_7499;
wire v_7500;
wire v_7501;
wire v_7502;
wire v_7503;
wire v_7504;
wire v_7505;
wire v_7506;
wire v_7507;
wire v_7508;
wire v_7509;
wire v_7510;
wire v_7511;
wire v_7512;
wire v_7513;
wire v_7514;
wire v_7515;
wire v_7516;
wire v_7517;
wire v_7518;
wire v_7519;
wire v_7520;
wire v_7521;
wire v_7522;
wire v_7523;
wire v_7524;
wire v_7525;
wire v_7526;
wire v_7527;
wire v_7528;
wire v_7529;
wire v_7530;
wire v_7531;
wire v_7532;
wire v_7533;
wire v_7534;
wire v_7535;
wire v_7536;
wire v_7537;
wire v_7538;
wire v_7539;
wire v_7540;
wire v_7541;
wire v_7542;
wire v_7543;
wire v_7544;
wire v_7545;
wire v_7546;
wire v_7547;
wire v_7548;
wire v_7549;
wire v_7550;
wire v_7551;
wire v_7552;
wire v_7553;
wire v_7554;
wire v_7555;
wire v_7556;
wire v_7557;
wire v_7558;
wire v_7559;
wire v_7560;
wire v_7561;
wire v_7562;
wire v_7563;
wire v_7564;
wire v_7565;
wire v_7566;
wire v_7567;
wire v_7568;
wire v_7569;
wire v_7570;
wire v_7571;
wire v_7572;
wire v_7573;
wire v_7574;
wire v_7575;
wire v_7576;
wire v_7577;
wire v_7578;
wire v_7579;
wire v_7580;
wire v_7581;
wire v_7582;
wire v_7583;
wire v_7584;
wire v_7585;
wire v_7586;
wire v_7587;
wire v_7588;
wire v_7589;
wire v_7590;
wire v_7591;
wire v_7592;
wire v_7593;
wire v_7594;
wire v_7595;
wire v_7596;
wire v_7597;
wire v_7598;
wire v_7599;
wire v_7600;
wire v_7601;
wire v_7602;
wire v_7603;
wire v_7604;
wire v_7605;
wire v_7606;
wire v_7607;
wire v_7608;
wire v_7609;
wire v_7610;
wire v_7611;
wire v_7612;
wire v_7613;
wire v_7614;
wire v_7615;
wire v_7616;
wire v_7617;
wire v_7618;
wire v_7619;
wire v_7620;
wire v_7621;
wire v_7622;
wire v_7623;
wire v_7624;
wire v_7625;
wire v_7626;
wire v_7627;
wire v_7628;
wire v_7629;
wire v_7630;
wire v_7631;
wire v_7632;
wire v_7633;
wire v_7634;
wire v_7635;
wire v_7636;
wire v_7637;
wire v_7638;
wire v_7639;
wire v_7640;
wire v_7641;
wire v_7642;
wire v_7643;
wire v_7644;
wire v_7645;
wire v_7646;
wire v_7647;
wire v_7648;
wire v_7649;
wire v_7650;
wire v_7651;
wire v_7652;
wire v_7653;
wire v_7654;
wire v_7655;
wire v_7656;
wire v_7657;
wire v_7658;
wire v_7659;
wire v_7660;
wire v_7661;
wire v_7662;
wire v_7663;
wire v_7664;
wire v_7665;
wire v_7666;
wire v_7667;
wire v_7668;
wire v_7669;
wire v_7670;
wire v_7671;
wire v_7672;
wire v_7673;
wire v_7674;
wire v_7675;
wire v_7676;
wire v_7677;
wire v_7678;
wire v_7679;
wire v_7680;
wire v_7681;
wire v_7682;
wire v_7683;
wire v_7684;
wire v_7685;
wire v_7686;
wire v_7687;
wire v_7688;
wire v_7689;
wire v_7690;
wire v_7691;
wire v_7692;
wire v_7693;
wire v_7694;
wire v_7695;
wire v_7696;
wire v_7697;
wire v_7698;
wire v_7699;
wire v_7700;
wire v_7701;
wire v_7702;
wire v_7703;
wire v_7704;
wire v_7705;
wire v_7706;
wire v_7707;
wire v_7708;
wire v_7709;
wire v_7710;
wire v_7711;
wire v_7712;
wire v_7713;
wire v_7714;
wire v_7715;
wire v_7716;
wire v_7717;
wire v_7718;
wire v_7719;
wire v_7720;
wire v_7721;
wire v_7722;
wire v_7723;
wire v_7724;
wire v_7725;
wire v_7726;
wire v_7727;
wire v_7728;
wire v_7729;
wire v_7730;
wire v_7731;
wire v_7732;
wire v_7733;
wire v_7734;
wire v_7735;
wire v_7736;
wire v_7737;
wire v_7738;
wire v_7739;
wire v_7740;
wire v_7741;
wire v_7742;
wire v_7743;
wire v_7744;
wire v_7745;
wire v_7746;
wire v_7747;
wire v_7748;
wire v_7749;
wire v_7750;
wire v_7751;
wire v_7752;
wire v_7753;
wire v_7754;
wire v_7755;
wire v_7756;
wire v_7757;
wire v_7758;
wire v_7759;
wire v_7760;
wire v_7761;
wire v_7762;
wire v_7763;
wire v_7764;
wire v_7765;
wire v_7766;
wire v_7767;
wire v_7768;
wire v_7769;
wire v_7770;
wire v_7771;
wire v_7772;
wire v_7773;
wire v_7774;
wire v_7775;
wire v_7776;
wire v_7777;
wire v_7778;
wire v_7779;
wire v_7780;
wire v_7781;
wire v_7782;
wire v_7783;
wire v_7784;
wire v_7785;
wire v_7786;
wire v_7787;
wire v_7788;
wire v_7789;
wire v_7790;
wire v_7791;
wire v_7792;
wire v_7793;
wire v_7794;
wire v_7795;
wire v_7796;
wire v_7797;
wire v_7798;
wire v_7799;
wire v_7800;
wire v_7801;
wire v_7802;
wire v_7803;
wire v_7804;
wire v_7805;
wire v_7806;
wire v_7807;
wire v_7808;
wire v_7809;
wire v_7810;
wire v_7811;
wire v_7812;
wire v_7813;
wire v_7814;
wire v_7815;
wire v_7816;
wire v_7817;
wire v_7818;
wire v_7819;
wire v_7820;
wire v_7821;
wire v_7822;
wire v_7823;
wire v_7824;
wire v_7825;
wire v_7826;
wire v_7827;
wire v_7828;
wire v_7829;
wire v_7830;
wire v_7831;
wire v_7832;
wire v_7833;
wire v_7834;
wire v_7835;
wire v_7836;
wire v_7837;
wire v_7838;
wire v_7839;
wire v_7840;
wire v_7841;
wire v_7842;
wire v_7843;
wire v_7844;
wire v_7845;
wire v_7846;
wire v_7847;
wire v_7848;
wire v_7849;
wire v_7850;
wire v_7851;
wire v_7852;
wire v_7853;
wire v_7854;
wire v_7855;
wire v_7856;
wire v_7857;
wire v_7858;
wire v_7859;
wire v_7860;
wire v_7861;
wire v_7862;
wire v_7863;
wire v_7864;
wire v_7865;
wire v_7866;
wire v_7867;
wire v_7868;
wire v_7869;
wire v_7870;
wire v_7871;
wire v_7872;
wire v_7873;
wire v_7874;
wire v_7875;
wire v_7876;
wire v_7877;
wire v_7878;
wire v_7879;
wire v_7880;
wire v_7881;
wire v_7882;
wire v_7883;
wire v_7884;
wire v_7885;
wire v_7886;
wire v_7887;
wire v_7888;
wire v_7889;
wire v_7890;
wire v_7891;
wire v_7892;
wire v_7893;
wire v_7894;
wire v_7895;
wire v_7896;
wire v_7897;
wire v_7898;
wire v_7899;
wire v_7900;
wire v_7901;
wire v_7902;
wire v_7903;
wire v_7904;
wire v_7905;
wire v_7906;
wire v_7907;
wire v_7908;
wire v_7909;
wire v_7910;
wire v_7911;
wire v_7912;
wire v_7913;
wire v_7914;
wire v_7915;
wire v_7916;
wire v_7917;
wire v_7918;
wire v_7919;
wire v_7920;
wire v_7921;
wire v_7922;
wire v_7923;
wire v_7924;
wire v_7925;
wire v_7926;
wire v_7927;
wire v_7928;
wire v_7929;
wire v_7930;
wire v_7931;
wire v_7932;
wire v_7933;
wire v_7934;
wire v_7935;
wire v_7936;
wire v_7937;
wire v_7938;
wire v_7939;
wire v_7940;
wire v_7941;
wire v_7942;
wire v_7943;
wire v_7944;
wire v_7945;
wire v_7946;
wire v_7947;
wire v_7948;
wire v_7949;
wire v_7950;
wire v_7951;
wire v_7952;
wire v_7953;
wire v_7954;
wire v_7955;
wire v_7956;
wire v_7957;
wire v_7958;
wire v_7959;
wire v_7960;
wire v_7961;
wire v_7962;
wire v_7963;
wire v_7964;
wire v_7965;
wire v_7966;
wire v_7967;
wire x_1;
assign v_1 = 1;
assign v_220 = 1;
assign v_226 = 1;
assign v_231 = 1;
assign v_250 = 1;
assign v_273 = 1;
assign v_339 = 1;
assign v_487 = 1;
assign v_490 = 1;
assign v_495 = 1;
assign v_514 = 1;
assign v_538 = 1;
assign v_550 = 1;
assign v_556 = 1;
assign v_564 = 1;
assign v_608 = 1;
assign v_614 = 1;
assign v_622 = 1;
assign v_664 = 1;
assign v_667 = 1;
assign v_714 = 1;
assign v_720 = 1;
assign v_728 = 1;
assign v_754 = 1;
assign v_756 = 1;
assign v_767 = 1;
assign v_769 = 1;
assign v_773 = 1;
assign v_783 = 1;
assign v_789 = 1;
assign v_1051 = 1;
assign v_2019 = 1;
assign v_4476 = 1;
assign v_4482 = 1;
assign v_4487 = 1;
assign v_4506 = 1;
assign v_4529 = 1;
assign v_4595 = 1;
assign v_4743 = 1;
assign v_4746 = 1;
assign v_4751 = 1;
assign v_4770 = 1;
assign v_4794 = 1;
assign v_4806 = 1;
assign v_4812 = 1;
assign v_4820 = 1;
assign v_4864 = 1;
assign v_4870 = 1;
assign v_4878 = 1;
assign v_4920 = 1;
assign v_4923 = 1;
assign v_4970 = 1;
assign v_4976 = 1;
assign v_4984 = 1;
assign v_5010 = 1;
assign v_5012 = 1;
assign v_5023 = 1;
assign v_5025 = 1;
assign v_5029 = 1;
assign v_5039 = 1;
assign v_5045 = 1;
assign v_5064 = 1;
assign v_5705 = 1;
assign v_6 = ~v_4 & ~v_5;
assign v_9 = ~v_7 & v_8;
assign v_10 = ~v_6 & ~v_9;
assign v_11 = ~v_4 & ~v_5;
assign v_12 = ~v_7 & v_8;
assign v_13 = ~v_11 & ~v_12;
assign v_14 = v_10 & v_13;
assign v_15 = ~v_4 & ~v_5;
assign v_16 = ~v_7 & v_8;
assign v_17 = ~v_15 & ~v_16;
assign v_18 = v_14 & v_17;
assign v_19 = ~v_4 & ~v_5;
assign v_20 = ~v_7 & v_8;
assign v_21 = ~v_19 & ~v_20;
assign v_22 = v_18 & v_21;
assign v_23 = ~v_4 & ~v_5;
assign v_24 = ~v_7 & v_8;
assign v_25 = ~v_23 & ~v_24;
assign v_26 = v_22 & v_25;
assign v_27 = ~v_4 & ~v_5;
assign v_28 = ~v_7 & v_8;
assign v_29 = ~v_27 & ~v_28;
assign v_30 = v_26 & v_29;
assign v_31 = ~v_4 & ~v_5;
assign v_32 = ~v_7 & v_8;
assign v_33 = ~v_31 & ~v_32;
assign v_34 = v_30 & v_33;
assign v_35 = ~v_4 & ~v_5;
assign v_36 = ~v_7 & v_8;
assign v_37 = ~v_35 & ~v_36;
assign v_38 = v_34 & v_37;
assign v_39 = ~v_4 & ~v_5;
assign v_40 = ~v_7 & v_8;
assign v_41 = ~v_39 & ~v_40;
assign v_42 = v_38 & v_41;
assign v_43 = ~v_4 & ~v_5;
assign v_44 = ~v_7 & v_8;
assign v_45 = ~v_43 & ~v_44;
assign v_46 = v_42 & v_45;
assign v_47 = ~v_4 & ~v_5;
assign v_48 = ~v_7 & v_8;
assign v_49 = ~v_47 & ~v_48;
assign v_50 = v_46 & v_49;
assign v_51 = ~v_4 & ~v_5;
assign v_52 = ~v_7 & v_8;
assign v_53 = ~v_51 & ~v_52;
assign v_54 = v_50 & v_53;
assign v_55 = ~v_4 & ~v_5;
assign v_56 = ~v_7 & v_8;
assign v_57 = ~v_55 & ~v_56;
assign v_58 = v_54 & v_57;
assign v_59 = ~v_4 & ~v_5;
assign v_60 = ~v_7 & v_8;
assign v_61 = ~v_59 & ~v_60;
assign v_62 = v_58 & v_61;
assign v_63 = ~v_4 & ~v_5;
assign v_64 = ~v_7 & v_8;
assign v_65 = ~v_63 & ~v_64;
assign v_66 = v_62 & v_65;
assign v_67 = ~v_4 & ~v_5;
assign v_68 = ~v_7 & v_8;
assign v_69 = ~v_67 & ~v_68;
assign v_70 = v_66 & v_69;
assign v_71 = ~v_4 & ~v_5;
assign v_72 = ~v_7 & v_8;
assign v_73 = ~v_71 & ~v_72;
assign v_74 = v_70 & v_73;
assign v_75 = ~v_4 & ~v_5;
assign v_76 = ~v_7 & v_8;
assign v_77 = ~v_75 & ~v_76;
assign v_78 = v_74 & v_77;
assign v_79 = ~v_4 & ~v_5;
assign v_80 = ~v_7 & v_8;
assign v_81 = ~v_79 & ~v_80;
assign v_82 = v_78 & v_81;
assign v_83 = ~v_4 & ~v_5;
assign v_84 = ~v_7 & v_8;
assign v_85 = ~v_83 & ~v_84;
assign v_86 = v_82 & v_85;
assign v_87 = ~v_4 & ~v_5;
assign v_88 = ~v_7 & v_8;
assign v_89 = ~v_87 & ~v_88;
assign v_90 = v_86 & v_89;
assign v_91 = ~v_4 & ~v_5;
assign v_92 = ~v_7 & v_8;
assign v_93 = ~v_91 & ~v_92;
assign v_94 = v_90 & v_93;
assign v_95 = ~v_4 & ~v_5;
assign v_96 = ~v_7 & v_8;
assign v_97 = ~v_95 & ~v_96;
assign v_98 = v_94 & v_97;
assign v_99 = ~v_4 & ~v_5;
assign v_100 = ~v_7 & v_8;
assign v_101 = ~v_99 & ~v_100;
assign v_102 = v_98 & v_101;
assign v_103 = ~v_4 & ~v_5;
assign v_104 = ~v_7 & v_8;
assign v_105 = ~v_103 & ~v_104;
assign v_106 = v_102 & v_105;
assign v_107 = ~v_4 & ~v_5;
assign v_108 = ~v_7 & v_8;
assign v_109 = ~v_107 & ~v_108;
assign v_110 = v_106 & v_109;
assign v_111 = ~v_4 & ~v_5;
assign v_112 = ~v_7 & v_8;
assign v_113 = ~v_111 & ~v_112;
assign v_114 = v_110 & v_113;
assign v_115 = ~v_4 & ~v_5;
assign v_116 = ~v_7 & v_8;
assign v_117 = ~v_115 & ~v_116;
assign v_118 = v_114 & v_117;
assign v_119 = ~v_4 & ~v_5;
assign v_120 = ~v_7 & v_8;
assign v_121 = ~v_119 & ~v_120;
assign v_122 = v_118 & v_121;
assign v_123 = ~v_4 & ~v_5;
assign v_124 = ~v_7 & v_8;
assign v_125 = ~v_123 & ~v_124;
assign v_126 = v_122 & v_125;
assign v_127 = ~v_4 & ~v_5;
assign v_128 = ~v_7 & v_8;
assign v_129 = ~v_127 & ~v_128;
assign v_130 = v_126 & v_129;
assign v_131 = ~v_4 & ~v_5;
assign v_132 = ~v_7 & v_8;
assign v_133 = ~v_131 & ~v_132;
assign v_134 = v_130 & v_133;
assign v_135 = ~v_4 & ~v_5;
assign v_136 = ~v_7 & v_8;
assign v_137 = ~v_135 & ~v_136;
assign v_138 = v_134 & v_137;
assign v_139 = ~v_4 & ~v_5;
assign v_140 = ~v_7 & v_8;
assign v_141 = ~v_139 & ~v_140;
assign v_142 = v_138 & v_141;
assign v_143 = ~v_4 & ~v_5;
assign v_144 = ~v_7 & v_8;
assign v_145 = ~v_143 & ~v_144;
assign v_146 = v_142 & v_145;
assign v_147 = ~v_4 & ~v_5;
assign v_148 = ~v_7 & v_8;
assign v_149 = ~v_147 & ~v_148;
assign v_150 = v_146 & v_149;
assign v_151 = ~v_4 & ~v_5;
assign v_152 = ~v_7 & v_8;
assign v_153 = ~v_151 & ~v_152;
assign v_154 = v_150 & v_153;
assign v_155 = ~v_4 & ~v_5;
assign v_156 = ~v_7 & v_8;
assign v_157 = ~v_155 & ~v_156;
assign v_158 = v_154 & v_157;
assign v_159 = ~v_4 & ~v_5;
assign v_160 = ~v_7 & v_8;
assign v_161 = ~v_159 & ~v_160;
assign v_162 = v_158 & v_161;
assign v_163 = ~v_4 & ~v_5;
assign v_164 = ~v_7 & v_8;
assign v_165 = ~v_163 & ~v_164;
assign v_166 = v_162 & v_165;
assign v_167 = ~v_4 & ~v_5;
assign v_168 = ~v_7 & v_8;
assign v_169 = ~v_167 & ~v_168;
assign v_170 = v_166 & v_169;
assign v_171 = ~v_4 & ~v_5;
assign v_172 = ~v_7 & v_8;
assign v_173 = ~v_171 & ~v_172;
assign v_174 = v_170 & v_173;
assign v_175 = ~v_4 & ~v_5;
assign v_176 = ~v_7 & v_8;
assign v_177 = ~v_175 & ~v_176;
assign v_178 = v_174 & v_177;
assign v_179 = ~v_4 & ~v_5;
assign v_180 = ~v_7 & v_8;
assign v_181 = ~v_179 & ~v_180;
assign v_182 = v_178 & v_181;
assign v_183 = ~v_4 & ~v_5;
assign v_184 = ~v_7 & v_8;
assign v_185 = ~v_183 & ~v_184;
assign v_186 = v_182 & v_185;
assign v_187 = ~v_4 & ~v_5;
assign v_188 = ~v_7 & v_8;
assign v_189 = ~v_187 & ~v_188;
assign v_190 = v_186 & v_189;
assign v_191 = ~v_4 & ~v_5;
assign v_192 = ~v_7 & v_8;
assign v_193 = ~v_191 & ~v_192;
assign v_194 = v_190 & v_193;
assign v_195 = ~v_4 & ~v_5;
assign v_196 = ~v_7 & v_8;
assign v_197 = ~v_195 & ~v_196;
assign v_198 = v_194 & v_197;
assign v_199 = ~v_4 & ~v_5;
assign v_200 = ~v_7 & v_8;
assign v_201 = ~v_199 & ~v_200;
assign v_202 = v_198 & v_201;
assign v_203 = ~v_7 & v_8;
assign v_204 = v_202 & ~v_203;
assign v_205 = ~v_7 & v_8;
assign v_206 = v_204 & ~v_205;
assign v_207 = ~v_7 & v_8;
assign v_208 = v_206 & ~v_207;
assign v_209 = ~v_7 & v_8;
assign v_210 = v_208 & ~v_209;
assign v_211 = ~v_7 & v_8;
assign v_212 = v_210 & ~v_211;
assign v_215 = v_213 & v_214;
assign v_216 = v_213 & ~v_214;
assign v_218 = v_212 & v_217;
assign v_222 = v_221;
assign v_223 = ~v_221;
assign v_228 = v_227;
assign v_233 = ~v_232;
assign v_235 = v_232 & v_234;
assign v_238 = v_232 & ~v_234 & v_236 & v_237;
assign v_240 = v_232 & ~v_234 & v_236 & ~v_237 & ~v_239;
assign v_242 = v_232 & ~v_234 & ~v_236 & ~v_241;
assign v_244 = v_232 & ~v_234 & ~v_236 & v_241 & v_243;
assign v_246 = v_7220 & v_7221;
assign v_248 = v_7222 & v_7223;
assign v_252 = v_7224 & v_7225;
assign v_253 = v_7226 & v_7227;
assign v_256 = v_254 & v_255;
assign v_257 = v_254 & ~v_255;
assign v_259 = v_7228 & v_7229;
assign v_261 = ~v_227 & ~v_229 & v_260;
assign v_263 = ~v_227 & v_229 & ~v_262;
assign v_265 = ~v_227 & v_229 & v_262 & ~v_264;
assign v_266 = ~v_227 & v_229 & v_262 & v_264;
assign v_269 = v_267 & v_268;
assign v_270 = v_267 & ~v_268;
assign v_275 = v_224 & v_271 & v_274;
assign v_276 = v_224 & v_271 & ~v_274;
assign v_278 = v_218 & v_277;
assign v_282 = v_280 & v_281;
assign v_284 = v_280 & ~v_281 & v_283;
assign v_287 = v_285 & ~v_286;
assign v_289 = v_285 & v_286 & v_288;
assign v_290 = v_285 & v_286 & ~v_288;
assign v_294 = v_279 & v_291 & v_292 & v_293;
assign v_296 = v_279 & v_291 & v_292 & ~v_293 & v_295;
assign v_299 = ~v_297 & v_298;
assign v_301 = v_279 & v_291 & ~v_292 & v_300;
assign v_304 = v_302 & v_303;
assign v_305 = v_302 & ~v_303;
assign v_307 = v_278 & v_306;
assign v_310 = ~v_308 & ~v_309;
assign v_313 = v_311 & v_312;
assign v_314 = v_311 & ~v_312;
assign v_317 = v_315 & ~v_316;
assign v_319 = v_315 & v_316 & v_318;
assign v_320 = v_315 & v_316 & ~v_318;
assign v_323 = v_321 & v_322;
assign v_325 = v_321 & ~v_322 & v_324;
assign v_327 = v_321 & ~v_322 & ~v_324 & v_326;
assign v_328 = v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_330 = ~v_308 & v_309 & v_329;
assign v_332 = v_307 & v_331;
assign v_335 = v_333 & ~v_334;
assign v_337 = v_333 & v_334 & ~v_336;
assign v_341 = v_333 & v_334 & v_336 & v_340;
assign v_342 = v_333 & v_334 & v_336 & ~v_340;
assign v_344 = v_332 & v_343;
assign v_347 = v_345 & v_346;
assign v_349 = v_345 & ~v_346 & v_348;
assign v_351 = v_345 & ~v_346 & ~v_348 & v_350;
assign v_353 = v_345 & ~v_346 & ~v_348 & ~v_350 & v_352;
assign v_355 = v_7230 & v_7231;
assign v_358 = v_356 & v_357;
assign v_361 = v_359 & v_360;
assign v_363 = v_359 & ~v_360 & v_362;
assign v_365 = v_359 & ~v_360 & ~v_362 & v_364;
assign v_367 = v_359 & ~v_360 & ~v_362 & ~v_364 & v_366;
assign v_368 = v_359 & ~v_360 & ~v_362 & ~v_364 & ~v_366;
assign v_371 = v_356 & ~v_357 & v_369 & v_370;
assign v_374 = v_372 & v_373;
assign v_376 = v_372 & ~v_373 & v_375;
assign v_378 = v_372 & ~v_373 & ~v_375 & v_377;
assign v_380 = v_372 & ~v_373 & ~v_375 & ~v_377 & v_379;
assign v_382 = v_7232 & v_7233;
assign v_383 = v_7234 & v_7235;
assign v_386 = v_384 & v_385;
assign v_387 = v_384 & ~v_385;
assign v_390 = v_7236 & v_7237;
assign v_393 = v_391 & v_392;
assign v_395 = v_391 & ~v_392 & v_394;
assign v_397 = v_391 & ~v_392 & ~v_394 & v_396;
assign v_399 = v_391 & ~v_392 & ~v_394 & ~v_396 & ~v_398;
assign v_401 = v_7238 & v_7239;
assign v_402 = v_7240 & v_7241;
assign v_404 = v_7242 & v_7243;
assign v_407 = v_405 & v_406;
assign v_408 = v_405 & ~v_406;
assign v_412 = v_410 & v_411;
assign v_414 = v_410 & ~v_411 & v_413;
assign v_416 = v_410 & ~v_411 & ~v_413 & v_415;
assign v_418 = v_410 & ~v_411 & ~v_413 & ~v_415 & v_417;
assign v_420 = v_7244 & v_7245;
assign v_423 = v_421 & v_422;
assign v_426 = v_424 & v_425;
assign v_428 = v_424 & ~v_425 & v_427;
assign v_430 = v_424 & ~v_425 & ~v_427 & v_429;
assign v_432 = v_424 & ~v_425 & ~v_427 & ~v_429 & v_431;
assign v_433 = v_424 & ~v_425 & ~v_427 & ~v_429 & ~v_431;
assign v_436 = v_421 & ~v_422 & v_434 & v_435;
assign v_439 = v_437 & v_438;
assign v_441 = v_437 & ~v_438 & v_440;
assign v_443 = v_437 & ~v_438 & ~v_440 & v_442;
assign v_445 = v_437 & ~v_438 & ~v_440 & ~v_442 & v_444;
assign v_447 = v_7246 & v_7247;
assign v_448 = v_7248 & v_7249;
assign v_451 = v_449 & v_450;
assign v_452 = v_449 & ~v_450;
assign v_455 = v_7250 & v_7251;
assign v_458 = v_456 & v_457;
assign v_460 = v_456 & ~v_457 & v_459;
assign v_462 = v_456 & ~v_457 & ~v_459 & v_461;
assign v_464 = v_456 & ~v_457 & ~v_459 & ~v_461 & ~v_463;
assign v_466 = v_7252 & v_7253;
assign v_467 = v_7254 & v_7255;
assign v_469 = v_7256 & v_7257;
assign v_472 = v_470 & v_471;
assign v_473 = v_470 & ~v_471;
assign v_476 = v_409 & v_474 & v_475;
assign v_478 = v_409 & v_474 & ~v_475 & v_477;
assign v_479 = v_409 & v_474 & ~v_475 & ~v_477;
assign v_482 = v_480 & v_481;
assign v_483 = v_480 & ~v_481;
assign v_485 = v_344 & v_484;
assign v_488 = v_485;
assign v_492 = v_491;
assign v_497 = ~v_496;
assign v_499 = v_496 & v_498;
assign v_502 = v_496 & ~v_498 & v_500 & v_501;
assign v_504 = v_496 & ~v_498 & v_500 & ~v_501 & ~v_503;
assign v_506 = v_496 & ~v_498 & ~v_500 & ~v_505;
assign v_508 = v_496 & ~v_498 & ~v_500 & v_505 & v_507;
assign v_510 = v_7258 & v_7259;
assign v_512 = v_7260 & v_7261;
assign v_516 = v_7262 & v_7263;
assign v_517 = v_7264 & v_7265;
assign v_520 = v_518 & v_519;
assign v_521 = v_518 & ~v_519;
assign v_523 = v_7266 & v_7267;
assign v_525 = ~v_491 & ~v_493 & v_524;
assign v_527 = ~v_491 & v_493 & ~v_526;
assign v_529 = ~v_491 & v_493 & v_526 & ~v_528;
assign v_530 = ~v_491 & v_493 & v_526 & v_528;
assign v_533 = v_531 & v_532;
assign v_534 = v_531 & ~v_532;
assign v_536 = v_488 & v_535;
assign v_539 = v_3 & v_536;
assign v_540 = ~v_3 & v_488 & v_535;
assign v_544 = v_542 & v_543;
assign v_545 = v_542 & ~v_543;
assign v_548 = v_546 & v_547;
assign v_552 = v_546 & ~v_547 & ~v_551;
assign v_553 = v_546 & ~v_547 & v_551;
assign v_557 = v_554;
assign v_560 = v_558 & v_559;
assign v_562 = v_558 & ~v_559 & v_561;
assign v_566 = v_558 & ~v_559 & ~v_561 & v_565;
assign v_567 = v_558 & ~v_559 & ~v_561 & ~v_565;
assign v_570 = v_568 & v_569;
assign v_572 = v_568 & ~v_569 & v_571;
assign v_575 = v_573 & v_574;
assign v_576 = v_573 & ~v_574;
assign v_579 = v_568 & ~v_569 & ~v_571 & v_577 & v_578;
assign v_580 = v_568 & ~v_569 & ~v_571 & v_577 & ~v_578;
assign v_582 = v_541 & v_581;
assign v_585 = ~v_583 & v_584;
assign v_587 = ~v_583 & ~v_584 & v_586;
assign v_590 = v_588 & v_589;
assign v_592 = v_588 & ~v_589 & v_591;
assign v_595 = v_593 & ~v_594;
assign v_596 = v_588 & ~v_589 & ~v_591;
assign v_597 = v_593 & v_594;
assign v_599 = v_582 & v_598;
assign v_602 = v_600 & v_601;
assign v_603 = v_600 & ~v_601;
assign v_606 = v_604 & v_605;
assign v_610 = v_604 & ~v_605 & ~v_609;
assign v_611 = v_604 & ~v_605 & v_609;
assign v_615 = v_612;
assign v_618 = v_616 & v_617;
assign v_620 = v_616 & ~v_617 & v_619;
assign v_624 = v_616 & ~v_617 & ~v_619 & v_623;
assign v_625 = v_616 & ~v_617 & ~v_619 & ~v_623;
assign v_628 = v_626 & v_627;
assign v_630 = v_626 & ~v_627 & v_629;
assign v_633 = v_631 & v_632;
assign v_634 = v_631 & ~v_632;
assign v_637 = v_626 & ~v_627 & ~v_629 & v_635 & v_636;
assign v_638 = v_626 & ~v_627 & ~v_629 & v_635 & ~v_636;
assign v_640 = v_2 & v_599 & v_639;
assign v_642 = v_641 & v_541 & v_581;
assign v_644 = v_643 & v_536;
assign v_646 = v_645 & v_536;
assign v_648 = v_647 & v_488 & v_535;
assign v_650 = v_649 & v_488 & v_535;
assign v_651 = ~v_649 & v_485;
assign v_653 = ~v_647 & v_652;
assign v_655 = ~v_645 & v_654;
assign v_657 = ~v_643 & v_656;
assign v_659 = ~v_641 & v_658;
assign v_661 = ~v_2 & v_660;
assign v_665 = v_662;
assign v_668 = v_665;
assign v_671 = v_669 & ~v_670;
assign v_673 = v_669 & v_670 & ~v_672;
assign v_676 = v_669 & v_670 & v_672 & ~v_674 & ~v_675;
assign v_677 = v_669 & v_670 & v_672 & v_674;
assign v_678 = v_669 & v_670 & v_672 & ~v_674 & v_675;
assign v_681 = v_679 & v_680;
assign v_683 = v_679 & ~v_680 & v_682;
assign v_686 = ~v_684 & v_685;
assign v_688 = ~v_684 & ~v_685 & v_687;
assign v_691 = v_689 & v_690;
assign v_693 = v_689 & ~v_690 & v_692;
assign v_696 = v_694 & ~v_695;
assign v_697 = v_689 & ~v_690 & ~v_692;
assign v_698 = v_694 & v_695;
assign v_701 = v_679 & ~v_680 & ~v_682 & v_699 & v_700;
assign v_702 = v_679 & ~v_680 & ~v_682 & v_699 & ~v_700;
assign v_704 = v_668 & v_703;
assign v_708 = v_706 & v_707;
assign v_709 = v_706 & ~v_707;
assign v_712 = v_710 & v_711;
assign v_716 = v_710 & ~v_711 & ~v_715;
assign v_717 = v_710 & ~v_711 & v_715;
assign v_721 = v_718;
assign v_725 = v_705 & v_722 & v_723 & ~v_724;
assign v_730 = v_7268 & v_7269;
assign v_732 = v_7270 & v_7271;
assign v_734 = v_7272 & v_7273;
assign v_736 = v_7274 & v_7275;
assign v_740 = v_737 & ~v_738 & v_739;
assign v_741 = v_737 & ~v_738 & ~v_739;
assign v_743 = v_737 & v_738 & v_742;
assign v_744 = v_737 & v_738 & ~v_742;
assign v_748 = v_746 & v_747;
assign v_749 = v_746 & ~v_747;
assign v_752 = v_750 & v_751;
assign v_757 = v_750 & ~v_751;
assign v_761 = v_759 & v_760;
assign v_762 = v_759 & ~v_760;
assign v_765 = v_763 & v_764;
assign v_770 = v_763 & ~v_764;
assign v_774 = v_745 & v_758 & v_771;
assign v_777 = v_775 & v_776;
assign v_778 = v_775 & ~v_776;
assign v_781 = v_779 & v_780;
assign v_785 = v_779 & ~v_780 & ~v_784;
assign v_786 = v_779 & ~v_780 & v_784;
assign v_790 = v_787;
assign v_793 = v_705 & v_722 & ~v_723 & v_791 & v_792;
assign v_794 = v_705 & v_722 & ~v_723 & v_791 & ~v_792;
assign v_795 = v_705 & v_722 & v_723 & v_724 & v_726;
assign v_797 = v_704 & v_796;
assign v_802 = v_800 & v_801;
assign v_803 = v_800 & ~v_801;
assign v_806 = v_804 & v_805;
assign v_807 = v_804 & ~v_805;
assign v_810 = v_808 & ~v_809;
assign v_812 = v_808 & v_809 & v_811;
assign v_813 = v_808 & v_809 & ~v_811;
assign v_816 = v_798 & v_799 & v_814 & v_815;
assign v_818 = v_798 & ~v_799 & v_817;
assign v_819 = v_798 & v_799 & v_814 & ~v_815;
assign v_820 = v_798 & ~v_799 & ~v_817;
assign v_825 = v_823 & v_824;
assign v_826 = v_823 & ~v_824;
assign v_829 = v_827 & v_828;
assign v_830 = v_827 & ~v_828;
assign v_833 = v_831 & ~v_832;
assign v_835 = v_831 & v_832 & v_834;
assign v_836 = v_831 & v_832 & ~v_834;
assign v_839 = v_821 & v_822 & v_837 & v_838;
assign v_841 = v_821 & ~v_822 & v_840;
assign v_842 = v_821 & v_822 & v_837 & ~v_838;
assign v_843 = v_821 & ~v_822 & ~v_840;
assign v_848 = v_846 & v_847;
assign v_849 = v_846 & ~v_847;
assign v_852 = v_850 & v_851;
assign v_853 = v_850 & ~v_851;
assign v_856 = v_854 & ~v_855;
assign v_858 = v_854 & v_855 & v_857;
assign v_859 = v_854 & v_855 & ~v_857;
assign v_862 = v_844 & v_845 & v_860 & v_861;
assign v_864 = v_844 & ~v_845 & v_863;
assign v_865 = v_844 & v_845 & v_860 & ~v_861;
assign v_866 = v_844 & ~v_845 & ~v_863;
assign v_871 = v_867 & v_868 & ~v_869 & v_870;
assign v_873 = v_867 & ~v_868 & v_872;
assign v_874 = v_867 & ~v_868 & ~v_872;
assign v_875 = v_867 & v_868 & ~v_869 & ~v_870;
assign v_876 = v_867 & v_868 & v_869;
assign v_878 = v_797 & v_877;
assign v_883 = v_881 & v_882;
assign v_884 = v_881 & ~v_882;
assign v_887 = v_885 & v_886;
assign v_888 = v_885 & ~v_886;
assign v_891 = v_889 & ~v_890;
assign v_893 = v_889 & v_890 & v_892;
assign v_894 = v_889 & v_890 & ~v_892;
assign v_897 = v_879 & v_880 & v_895 & v_896;
assign v_899 = v_879 & ~v_880 & v_898;
assign v_900 = v_879 & v_880 & v_895 & ~v_896;
assign v_901 = v_879 & ~v_880 & ~v_898;
assign v_906 = v_904 & v_905;
assign v_907 = v_904 & ~v_905;
assign v_910 = v_908 & v_909;
assign v_911 = v_908 & ~v_909;
assign v_914 = v_912 & ~v_913;
assign v_916 = v_912 & v_913 & v_915;
assign v_917 = v_912 & v_913 & ~v_915;
assign v_920 = v_902 & v_903 & v_918 & v_919;
assign v_922 = v_902 & ~v_903 & v_921;
assign v_923 = v_902 & v_903 & v_918 & ~v_919;
assign v_924 = v_902 & ~v_903 & ~v_921;
assign v_929 = v_927 & v_928;
assign v_930 = v_927 & ~v_928;
assign v_933 = v_931 & v_932;
assign v_934 = v_931 & ~v_932;
assign v_937 = v_935 & ~v_936;
assign v_939 = v_935 & v_936 & v_938;
assign v_940 = v_935 & v_936 & ~v_938;
assign v_943 = v_925 & v_926 & v_941 & v_942;
assign v_945 = v_925 & ~v_926 & v_944;
assign v_946 = v_925 & v_926 & v_941 & ~v_942;
assign v_947 = v_925 & ~v_926 & ~v_944;
assign v_952 = v_948 & v_949 & ~v_950 & v_951;
assign v_954 = v_948 & ~v_949 & v_953;
assign v_955 = v_948 & ~v_949 & ~v_953;
assign v_956 = v_948 & v_949 & ~v_950 & ~v_951;
assign v_957 = v_948 & v_949 & v_950;
assign v_959 = v_878 & v_958;
assign v_964 = v_962 & v_963;
assign v_965 = v_962 & ~v_963;
assign v_968 = v_966 & v_967;
assign v_969 = v_966 & ~v_967;
assign v_972 = v_970 & ~v_971;
assign v_974 = v_970 & v_971 & v_973;
assign v_975 = v_970 & v_971 & ~v_973;
assign v_978 = v_960 & v_961 & v_976 & v_977;
assign v_980 = v_960 & ~v_961 & v_979;
assign v_981 = v_960 & v_961 & v_976 & ~v_977;
assign v_982 = v_960 & ~v_961 & ~v_979;
assign v_987 = v_985 & v_986;
assign v_988 = v_985 & ~v_986;
assign v_991 = v_989 & v_990;
assign v_992 = v_989 & ~v_990;
assign v_995 = v_993 & ~v_994;
assign v_997 = v_993 & v_994 & v_996;
assign v_998 = v_993 & v_994 & ~v_996;
assign v_1001 = v_983 & v_984 & v_999 & v_1000;
assign v_1003 = v_983 & ~v_984 & v_1002;
assign v_1004 = v_983 & v_984 & v_999 & ~v_1000;
assign v_1005 = v_983 & ~v_984 & ~v_1002;
assign v_1010 = v_1008 & v_1009;
assign v_1011 = v_1008 & ~v_1009;
assign v_1014 = v_1012 & v_1013;
assign v_1015 = v_1012 & ~v_1013;
assign v_1018 = v_1016 & ~v_1017;
assign v_1020 = v_1016 & v_1017 & v_1019;
assign v_1021 = v_1016 & v_1017 & ~v_1019;
assign v_1024 = v_1006 & v_1007 & v_1022 & v_1023;
assign v_1026 = v_1006 & ~v_1007 & v_1025;
assign v_1027 = v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_1028 = v_1006 & ~v_1007 & ~v_1025;
assign v_1033 = v_1029 & v_1030 & ~v_1031 & v_1032;
assign v_1035 = v_1029 & ~v_1030 & v_1034;
assign v_1036 = v_1029 & ~v_1030 & ~v_1034;
assign v_1037 = v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_1038 = v_1029 & v_1030 & v_1031;
assign v_1040 = v_959 & v_1039;
assign v_1044 = v_1042 & ~v_1043;
assign v_1046 = v_1041 & v_1045;
assign v_1048 = ~v_227 & v_229 & v_262 & ~v_264;
assign v_1049 = ~v_227 & v_229 & v_262 & v_264;
assign v_1050 = ~v_227 & v_229 & ~v_262;
assign v_1053 = v_1052;
assign v_1055 = v_1054;
assign v_1056 = v_7276 & v_7277;
assign v_1058 = v_1057 & ~v_227 & ~v_229 & v_260;
assign v_1060 = v_1047 & ~v_1059;
assign v_1062 = v_1061 & v_267 & v_268;
assign v_1063 = v_1061 & v_267 & ~v_268;
assign v_1065 = v_1064 & ~v_279;
assign v_1067 = v_1064 & v_1066;
assign v_1068 = v_1064 & v_279 & v_291 & ~v_292 & v_300;
assign v_1071 = v_1069 & v_1070;
assign v_1072 = v_1069 & v_321 & v_322;
assign v_1073 = v_1069 & v_321 & ~v_322 & v_324;
assign v_1074 = v_1069 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_1075 = v_1069 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_1078 = v_1076 & v_1077;
assign v_1080 = v_1079 & ~v_308 & v_309 & v_329;
assign v_1083 = v_1081 & v_1082;
assign v_1085 = v_1081 & v_1084;
assign v_1087 = ~v_1041 & v_1086;
assign v_1089 = v_1088 & v_345 & v_346;
assign v_1090 = v_1088 & v_345 & ~v_346 & v_348;
assign v_1091 = v_1088 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_1092 = v_1088 & v_356 & v_357;
assign v_1093 = v_1088 & v_359 & v_360;
assign v_1094 = v_1088 & v_359 & ~v_360 & v_362;
assign v_1095 = v_1088 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_1097 = v_1088 & v_1096;
assign v_1100 = v_1098 & v_1099;
assign v_1102 = v_1101 & v_356 & ~v_357 & v_369 & v_370;
assign v_1103 = v_1101 & v_372 & v_373;
assign v_1104 = v_1101 & v_372 & ~v_373 & v_375;
assign v_1105 = v_1101 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_1107 = v_1101 & v_1106;
assign v_1108 = v_7278 & v_7279;
assign v_1110 = v_1109 & v_384 & v_385;
assign v_1111 = v_1109 & v_384 & ~v_385;
assign v_1114 = v_1112 & v_1113;
assign v_1116 = v_7280 & v_7281;
assign v_1117 = v_1115 & v_391 & v_392;
assign v_1118 = v_1115 & v_391 & ~v_392 & v_394;
assign v_1119 = v_1115 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_1121 = v_1115 & v_1120;
assign v_1123 = v_7282 & v_7283;
assign v_1126 = v_1124 & v_1125;
assign v_1128 = v_1127 & v_410 & v_411;
assign v_1129 = v_1127 & v_410 & ~v_411 & v_413;
assign v_1130 = v_1127 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_1131 = v_1127 & v_421 & v_422;
assign v_1132 = v_1127 & v_424 & v_425;
assign v_1133 = v_1127 & v_424 & ~v_425 & v_427;
assign v_1134 = v_1127 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_1136 = v_1127 & v_1135;
assign v_1139 = v_1137 & v_1138;
assign v_1141 = v_1140 & v_421 & ~v_422 & v_434 & v_435;
assign v_1142 = v_1140 & v_437 & v_438;
assign v_1143 = v_1140 & v_437 & ~v_438 & v_440;
assign v_1144 = v_1140 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_1146 = v_1140 & v_1145;
assign v_1147 = v_7284 & v_7285;
assign v_1149 = v_1148 & v_449 & v_450;
assign v_1150 = v_1148 & v_449 & ~v_450;
assign v_1153 = v_1151 & v_1152;
assign v_1155 = v_7286 & v_7287;
assign v_1156 = v_1154 & v_456 & v_457;
assign v_1157 = v_1154 & v_456 & ~v_457 & v_459;
assign v_1158 = v_1154 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_1160 = v_1154 & v_1159;
assign v_1162 = v_7288 & v_7289;
assign v_1165 = v_1163 & v_1164;
assign v_1167 = v_1166 & v_491;
assign v_1170 = v_1169 & ~v_1166;
assign v_1172 = v_1171 & ~v_491 & v_493 & v_526 & ~v_528;
assign v_1173 = v_1171 & ~v_491 & v_493 & v_526 & v_528;
assign v_1174 = v_1171 & ~v_491 & v_493 & ~v_526;
assign v_1175 = v_1171 & v_494;
assign v_1176 = v_1171 & ~v_494;
assign v_1179 = v_1177 & v_1178;
assign v_1181 = v_1177 & v_1180;
assign v_1182 = v_7290 & v_7291;
assign v_1184 = v_1183 & ~v_491 & ~v_493 & v_524;
assign v_1186 = v_1168 & ~v_1185;
assign v_1188 = v_1187 & v_531 & v_532;
assign v_1189 = v_1187 & v_531 & ~v_532;
assign v_1191 = v_1190 & v_546 & v_547;
assign v_1192 = v_1190 & v_554;
assign v_1194 = v_1193 & v_558 & v_559;
assign v_1195 = v_1193 & v_558 & ~v_559 & v_561;
assign v_1197 = v_1193 & v_1196;
assign v_1200 = v_1198 & v_1199;
assign v_1202 = v_1198 & v_1201;
assign v_1204 = v_1203 & v_588 & ~v_589 & ~v_591;
assign v_1205 = v_1203 & v_593 & ~v_594;
assign v_1206 = v_1203 & v_593 & v_594;
assign v_1207 = v_1203 & v_583;
assign v_1209 = v_1208 & v_604 & v_605;
assign v_1210 = v_1208 & v_612;
assign v_1212 = v_1211 & v_616 & v_617;
assign v_1213 = v_1211 & v_616 & ~v_617 & v_619;
assign v_1215 = v_1211 & v_1214;
assign v_1218 = v_1216 & v_1217;
assign v_1220 = v_1216 & v_1219;
assign v_1222 = v_2 & v_1221;
assign v_1223 = v_641 & v_1203;
assign v_1224 = v_643 & v_1190;
assign v_1225 = v_645 & v_1190;
assign v_1226 = v_647 & v_1190;
assign v_1227 = v_649 & v_1190;
assign v_1228 = ~v_649 & v_1166;
assign v_1230 = ~v_647 & v_1229;
assign v_1232 = ~v_645 & v_1231;
assign v_1234 = ~v_643 & v_1233;
assign v_1236 = ~v_641 & v_1235;
assign v_1238 = ~v_2 & v_1237;
assign v_1240 = v_1239 & ~v_669;
assign v_1241 = v_7292 & v_7293;
assign v_1242 = v_1239 & v_669 & v_670 & v_672 & v_674;
assign v_1243 = v_7294 & v_7295;
assign v_1245 = v_1244 & v_679 & ~v_680 & v_682;
assign v_1246 = v_1244 & v_689 & ~v_690 & ~v_692;
assign v_1247 = v_1244 & v_694 & ~v_695;
assign v_1248 = v_1244 & v_694 & v_695;
assign v_1249 = v_1244 & v_684;
assign v_1252 = v_1250 & v_1251;
assign v_1255 = v_1253 & v_1254;
assign v_1256 = v_1244 & v_679 & v_680;
assign v_1258 = v_1239 & v_1257;
assign v_1260 = v_1259 & ~v_705;
assign v_1261 = v_1259 & v_710 & v_711;
assign v_1262 = v_1259 & v_718;
assign v_1264 = v_1263 & v_705 & v_722 & v_723 & ~v_724;
assign v_1266 = v_1263 & v_1265;
assign v_1267 = v_1263 & v_750 & v_751;
assign v_1268 = v_1263 & v_750 & ~v_751;
assign v_1270 = v_1269 & v_763 & v_764;
assign v_1271 = v_1269 & v_763 & ~v_764;
assign v_1273 = v_1272 & v_745 & v_758 & v_771;
assign v_1274 = v_7296 & v_7297;
assign v_1275 = v_1263 & v_779 & v_780;
assign v_1276 = v_1263 & v_787;
assign v_1279 = v_1277 & v_1278;
assign v_1281 = v_1280 & v_798 & ~v_799 & v_817;
assign v_1282 = v_1280 & v_798 & ~v_799 & ~v_817;
assign v_1283 = v_1280 & ~v_800;
assign v_1284 = v_1280 & v_808 & ~v_809;
assign v_1286 = v_1280 & v_1285;
assign v_1288 = v_1287 & v_798 & v_799 & v_814 & ~v_815;
assign v_1290 = v_1289 & v_821 & ~v_822 & v_840;
assign v_1291 = v_1289 & v_821 & ~v_822 & ~v_840;
assign v_1292 = v_1289 & ~v_823;
assign v_1293 = v_1289 & v_831 & ~v_832;
assign v_1295 = v_1289 & v_1294;
assign v_1297 = v_1296 & v_821 & v_822 & v_837 & ~v_838;
assign v_1299 = v_1298 & v_844 & ~v_845 & v_863;
assign v_1300 = v_1298 & ~v_846;
assign v_1301 = v_1298 & v_854 & ~v_855;
assign v_1303 = v_1298 & v_1302;
assign v_1305 = v_1304 & v_844 & v_845 & v_860 & v_861;
assign v_1306 = v_1298 & v_844 & ~v_845 & ~v_863;
assign v_1307 = v_1304 & v_844 & v_845 & v_860 & ~v_861;
assign v_1310 = v_1308 & v_1309;
assign v_1311 = v_1308 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_1312 = v_1308 & v_867 & v_868 & v_869;
assign v_1313 = v_1308 & v_867 & ~v_868 & ~v_872;
assign v_1316 = v_1314 & v_1315;
assign v_1317 = v_1296 & v_821 & v_822 & v_837 & v_838;
assign v_1318 = v_1287 & v_798 & v_799 & v_814 & v_815;
assign v_1320 = v_1319 & v_879 & ~v_880 & v_898;
assign v_1321 = v_1319 & v_879 & ~v_880 & ~v_898;
assign v_1322 = v_1319 & ~v_881;
assign v_1323 = v_1319 & v_889 & ~v_890;
assign v_1325 = v_1319 & v_1324;
assign v_1327 = v_1326 & v_879 & v_880 & v_895 & ~v_896;
assign v_1329 = v_1328 & v_902 & ~v_903 & v_921;
assign v_1330 = v_1328 & v_902 & ~v_903 & ~v_921;
assign v_1331 = v_1328 & ~v_904;
assign v_1332 = v_1328 & v_912 & ~v_913;
assign v_1334 = v_1328 & v_1333;
assign v_1336 = v_1335 & v_902 & v_903 & v_918 & ~v_919;
assign v_1338 = v_1337 & v_925 & ~v_926 & v_944;
assign v_1339 = v_1337 & ~v_927;
assign v_1340 = v_1337 & v_935 & ~v_936;
assign v_1342 = v_1337 & v_1341;
assign v_1344 = v_1343 & v_925 & v_926 & v_941 & v_942;
assign v_1345 = v_1337 & v_925 & ~v_926 & ~v_944;
assign v_1346 = v_1343 & v_925 & v_926 & v_941 & ~v_942;
assign v_1349 = v_1347 & v_1348;
assign v_1350 = v_1347 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_1351 = v_1347 & v_948 & v_949 & v_950;
assign v_1352 = v_1347 & v_948 & ~v_949 & ~v_953;
assign v_1355 = v_1353 & v_1354;
assign v_1356 = v_1335 & v_902 & v_903 & v_918 & v_919;
assign v_1357 = v_1326 & v_879 & v_880 & v_895 & v_896;
assign v_1359 = v_1358 & v_960 & ~v_961 & v_979;
assign v_1360 = v_1358 & v_960 & ~v_961 & ~v_979;
assign v_1361 = v_1358 & ~v_962;
assign v_1362 = v_1358 & v_970 & ~v_971;
assign v_1364 = v_1358 & v_1363;
assign v_1366 = v_1365 & v_960 & v_961 & v_976 & ~v_977;
assign v_1368 = v_1367 & v_983 & ~v_984 & v_1002;
assign v_1369 = v_1367 & v_983 & ~v_984 & ~v_1002;
assign v_1370 = v_1367 & ~v_985;
assign v_1371 = v_1367 & v_993 & ~v_994;
assign v_1373 = v_1367 & v_1372;
assign v_1375 = v_1374 & v_983 & v_984 & v_999 & ~v_1000;
assign v_1377 = v_1376 & v_1006 & ~v_1007 & v_1025;
assign v_1378 = v_1376 & ~v_1008;
assign v_1379 = v_1376 & v_1016 & ~v_1017;
assign v_1381 = v_1376 & v_1380;
assign v_1383 = v_1382 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_1384 = v_1376 & v_1006 & ~v_1007 & ~v_1025;
assign v_1385 = v_1382 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_1388 = v_1386 & v_1387;
assign v_1389 = v_1386 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_1390 = v_1386 & v_1029 & v_1030 & v_1031;
assign v_1391 = v_1386 & v_1029 & ~v_1030 & ~v_1034;
assign v_1394 = v_1392 & v_1393;
assign v_1395 = v_1374 & v_983 & v_984 & v_999 & v_1000;
assign v_1396 = v_1365 & v_960 & v_961 & v_976 & v_977;
assign v_1400 = v_1041 & v_1399;
assign v_1401 = v_227;
assign v_1404 = v_1403 & v_267 & v_268;
assign v_1405 = v_1403 & v_267 & ~v_268;
assign v_1407 = v_1406 & ~v_279;
assign v_1409 = v_1406 & v_1408;
assign v_1410 = v_1406 & v_279 & v_291 & ~v_292 & v_300;
assign v_1413 = v_1411 & v_1412;
assign v_1414 = v_1411 & v_321 & v_322;
assign v_1415 = v_1411 & v_321 & ~v_322 & v_324;
assign v_1416 = v_1411 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_1417 = v_1411 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_1419 = v_1418 & v_1077;
assign v_1421 = v_1420 & ~v_308 & v_309 & v_329;
assign v_1424 = v_1422 & v_1423;
assign v_1425 = v_1422 & v_1084;
assign v_1427 = ~v_1041 & v_1426;
assign v_1429 = v_1428 & v_345 & v_346;
assign v_1430 = v_1428 & v_345 & ~v_346 & v_348;
assign v_1431 = v_1428 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_1432 = v_1428 & v_356 & v_357;
assign v_1433 = v_1428 & v_359 & v_360;
assign v_1434 = v_1428 & v_359 & ~v_360 & v_362;
assign v_1435 = v_1428 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_1436 = v_1428 & v_1096;
assign v_1438 = v_1437 & v_1099;
assign v_1440 = v_1439 & v_356 & ~v_357 & v_369 & v_370;
assign v_1441 = v_1439 & v_372 & v_373;
assign v_1442 = v_1439 & v_372 & ~v_373 & v_375;
assign v_1443 = v_1439 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_1445 = v_1439 & v_1444;
assign v_1446 = v_7298 & v_7299;
assign v_1448 = v_1447 & v_384 & v_385;
assign v_1449 = v_1447 & v_384 & ~v_385;
assign v_1451 = v_1450 & v_1113;
assign v_1453 = v_7300 & v_7301;
assign v_1454 = v_1452 & v_391 & v_392;
assign v_1455 = v_1452 & v_391 & ~v_392 & v_394;
assign v_1456 = v_1452 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_1457 = v_1452 & v_1120;
assign v_1459 = v_7302 & v_7303;
assign v_1461 = v_1460 & v_1125;
assign v_1463 = v_1462 & v_410 & v_411;
assign v_1464 = v_1462 & v_410 & ~v_411 & v_413;
assign v_1465 = v_1462 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_1466 = v_1462 & v_421 & v_422;
assign v_1467 = v_1462 & v_424 & v_425;
assign v_1468 = v_1462 & v_424 & ~v_425 & v_427;
assign v_1469 = v_1462 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_1470 = v_1462 & v_1135;
assign v_1472 = v_1471 & v_1138;
assign v_1474 = v_1473 & v_421 & ~v_422 & v_434 & v_435;
assign v_1475 = v_1473 & v_437 & v_438;
assign v_1476 = v_1473 & v_437 & ~v_438 & v_440;
assign v_1477 = v_1473 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_1479 = v_1473 & v_1478;
assign v_1480 = v_7304 & v_7305;
assign v_1482 = v_1481 & v_449 & v_450;
assign v_1483 = v_1481 & v_449 & ~v_450;
assign v_1485 = v_1484 & v_1152;
assign v_1487 = v_7306 & v_7307;
assign v_1488 = v_1486 & v_456 & v_457;
assign v_1489 = v_1486 & v_456 & ~v_457 & v_459;
assign v_1490 = v_1486 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_1491 = v_1486 & v_1159;
assign v_1493 = v_7308 & v_7309;
assign v_1495 = v_1494 & v_1164;
assign v_1497 = v_1496 & v_491;
assign v_1500 = v_1499 & v_531 & v_532;
assign v_1501 = v_1499 & v_531 & ~v_532;
assign v_1503 = v_1502 & v_546 & v_547;
assign v_1504 = v_1502 & v_554;
assign v_1506 = v_1505 & v_558 & v_559;
assign v_1507 = v_1505 & v_558 & ~v_559 & v_561;
assign v_1508 = v_1505 & v_1196;
assign v_1511 = v_1509 & v_1510;
assign v_1512 = v_1509 & v_1201;
assign v_1514 = v_1513 & v_588 & ~v_589 & ~v_591;
assign v_1515 = v_1513 & v_593 & ~v_594;
assign v_1516 = v_1513 & v_593 & v_594;
assign v_1517 = v_1513 & v_583;
assign v_1519 = v_1518 & v_604 & v_605;
assign v_1520 = v_1518 & v_612;
assign v_1522 = v_1521 & v_616 & v_617;
assign v_1523 = v_1521 & v_616 & ~v_617 & v_619;
assign v_1524 = v_1521 & v_1214;
assign v_1527 = v_1525 & v_1526;
assign v_1528 = v_1525 & v_1219;
assign v_1530 = v_2 & v_1529;
assign v_1531 = v_641 & v_1513;
assign v_1532 = v_643 & v_1502;
assign v_1533 = v_645 & v_1502;
assign v_1534 = v_647 & v_1502;
assign v_1535 = v_649 & v_1502;
assign v_1536 = ~v_649 & v_1496;
assign v_1538 = ~v_647 & v_1537;
assign v_1540 = ~v_645 & v_1539;
assign v_1542 = ~v_643 & v_1541;
assign v_1544 = ~v_641 & v_1543;
assign v_1546 = ~v_2 & v_1545;
assign v_1548 = v_1547 & ~v_669;
assign v_1549 = v_7310 & v_7311;
assign v_1550 = v_1547 & v_669 & v_670 & v_672 & v_674;
assign v_1551 = v_7312 & v_7313;
assign v_1553 = v_1552 & v_679 & ~v_680 & v_682;
assign v_1554 = v_1552 & v_689 & ~v_690 & ~v_692;
assign v_1555 = v_1552 & v_694 & ~v_695;
assign v_1556 = v_1552 & v_694 & v_695;
assign v_1557 = v_1552 & v_684;
assign v_1559 = v_1558 & v_1251;
assign v_1561 = v_1560 & v_1254;
assign v_1562 = v_1552 & v_679 & v_680;
assign v_1563 = v_1547 & v_1257;
assign v_1565 = v_1564 & ~v_705;
assign v_1566 = v_1564 & v_710 & v_711;
assign v_1567 = v_1564 & v_718;
assign v_1569 = v_1568 & v_705 & v_722 & v_723 & ~v_724;
assign v_1571 = v_1568 & v_1570;
assign v_1572 = v_1568 & v_750 & v_751;
assign v_1573 = v_1568 & v_750 & ~v_751;
assign v_1575 = v_1574 & v_763 & v_764;
assign v_1576 = v_1574 & v_763 & ~v_764;
assign v_1578 = v_1577 & v_745 & v_758 & v_771;
assign v_1579 = v_7314 & v_7315;
assign v_1580 = v_1568 & v_779 & v_780;
assign v_1581 = v_1568 & v_787;
assign v_1583 = v_1582 & v_1278;
assign v_1585 = v_1584 & v_798 & ~v_799 & v_817;
assign v_1586 = v_1584 & v_798 & ~v_799 & ~v_817;
assign v_1587 = v_1584 & ~v_800;
assign v_1588 = v_1584 & v_808 & ~v_809;
assign v_1589 = v_1584 & v_1285;
assign v_1591 = v_1590 & v_798 & v_799 & v_814 & ~v_815;
assign v_1593 = v_1592 & v_821 & ~v_822 & v_840;
assign v_1594 = v_1592 & v_821 & ~v_822 & ~v_840;
assign v_1595 = v_1592 & ~v_823;
assign v_1596 = v_1592 & v_831 & ~v_832;
assign v_1597 = v_1592 & v_1294;
assign v_1599 = v_1598 & v_821 & v_822 & v_837 & ~v_838;
assign v_1601 = v_1600 & v_844 & ~v_845 & v_863;
assign v_1602 = v_1600 & ~v_846;
assign v_1603 = v_1600 & v_854 & ~v_855;
assign v_1604 = v_1600 & v_1302;
assign v_1606 = v_1605 & v_844 & v_845 & v_860 & v_861;
assign v_1607 = v_1600 & v_844 & ~v_845 & ~v_863;
assign v_1608 = v_1605 & v_844 & v_845 & v_860 & ~v_861;
assign v_1611 = v_1609 & v_1610;
assign v_1612 = v_1609 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_1613 = v_1609 & v_867 & v_868 & v_869;
assign v_1614 = v_1609 & v_867 & ~v_868 & ~v_872;
assign v_1616 = v_1615 & v_1315;
assign v_1617 = v_1598 & v_821 & v_822 & v_837 & v_838;
assign v_1618 = v_1590 & v_798 & v_799 & v_814 & v_815;
assign v_1620 = v_1619 & v_879 & ~v_880 & v_898;
assign v_1621 = v_1619 & v_879 & ~v_880 & ~v_898;
assign v_1622 = v_1619 & ~v_881;
assign v_1623 = v_1619 & v_889 & ~v_890;
assign v_1624 = v_1619 & v_1324;
assign v_1626 = v_1625 & v_879 & v_880 & v_895 & ~v_896;
assign v_1628 = v_1627 & v_902 & ~v_903 & v_921;
assign v_1629 = v_1627 & v_902 & ~v_903 & ~v_921;
assign v_1630 = v_1627 & ~v_904;
assign v_1631 = v_1627 & v_912 & ~v_913;
assign v_1632 = v_1627 & v_1333;
assign v_1634 = v_1633 & v_902 & v_903 & v_918 & ~v_919;
assign v_1636 = v_1635 & v_925 & ~v_926 & v_944;
assign v_1637 = v_1635 & ~v_927;
assign v_1638 = v_1635 & v_935 & ~v_936;
assign v_1639 = v_1635 & v_1341;
assign v_1641 = v_1640 & v_925 & v_926 & v_941 & v_942;
assign v_1642 = v_1635 & v_925 & ~v_926 & ~v_944;
assign v_1643 = v_1640 & v_925 & v_926 & v_941 & ~v_942;
assign v_1646 = v_1644 & v_1645;
assign v_1647 = v_1644 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_1648 = v_1644 & v_948 & v_949 & v_950;
assign v_1649 = v_1644 & v_948 & ~v_949 & ~v_953;
assign v_1651 = v_1650 & v_1354;
assign v_1652 = v_1633 & v_902 & v_903 & v_918 & v_919;
assign v_1653 = v_1625 & v_879 & v_880 & v_895 & v_896;
assign v_1655 = v_1654 & v_960 & ~v_961 & v_979;
assign v_1656 = v_1654 & v_960 & ~v_961 & ~v_979;
assign v_1657 = v_1654 & ~v_962;
assign v_1658 = v_1654 & v_970 & ~v_971;
assign v_1659 = v_1654 & v_1363;
assign v_1661 = v_1660 & v_960 & v_961 & v_976 & ~v_977;
assign v_1663 = v_1662 & v_983 & ~v_984 & v_1002;
assign v_1664 = v_1662 & v_983 & ~v_984 & ~v_1002;
assign v_1665 = v_1662 & ~v_985;
assign v_1666 = v_1662 & v_993 & ~v_994;
assign v_1667 = v_1662 & v_1372;
assign v_1669 = v_1668 & v_983 & v_984 & v_999 & ~v_1000;
assign v_1671 = v_1670 & v_1006 & ~v_1007 & v_1025;
assign v_1672 = v_1670 & ~v_1008;
assign v_1673 = v_1670 & v_1016 & ~v_1017;
assign v_1674 = v_1670 & v_1380;
assign v_1676 = v_1675 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_1677 = v_1670 & v_1006 & ~v_1007 & ~v_1025;
assign v_1678 = v_1675 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_1681 = v_1679 & v_1680;
assign v_1682 = v_1679 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_1683 = v_1679 & v_1029 & v_1030 & v_1031;
assign v_1684 = v_1679 & v_1029 & ~v_1030 & ~v_1034;
assign v_1686 = v_1685 & v_1393;
assign v_1687 = v_1668 & v_983 & v_984 & v_999 & v_1000;
assign v_1688 = v_1660 & v_960 & v_961 & v_976 & v_977;
assign v_1690 = v_8 & v_227;
assign v_1691 = v_8 & ~v_227 & v_229 & v_262 & ~v_264;
assign v_1692 = v_8 & ~v_227 & v_229 & v_262 & v_264;
assign v_1693 = v_8 & ~v_227 & v_229 & ~v_262;
assign v_1694 = v_8 & v_230;
assign v_1695 = v_8 & ~v_230;
assign v_1698 = v_1696 & v_1697;
assign v_1699 = v_1696 & v_1054;
assign v_1700 = v_7316 & v_7317;
assign v_1702 = v_1701 & ~v_227 & ~v_229 & v_260;
assign v_1704 = v_1703 & v_267 & v_268;
assign v_1705 = v_1703 & v_267 & ~v_268;
assign v_1707 = v_1706 & ~v_279;
assign v_1709 = v_1706 & v_1708;
assign v_1710 = v_1706 & v_279 & v_291 & ~v_292 & v_300;
assign v_1713 = v_1711 & v_1712;
assign v_1714 = v_1711 & v_321 & v_322;
assign v_1715 = v_1711 & v_321 & ~v_322 & v_324;
assign v_1716 = v_1711 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_1717 = v_1711 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_1719 = v_1718 & v_1077;
assign v_1721 = v_1720 & ~v_308 & v_309 & v_329;
assign v_1724 = v_1722 & v_1723;
assign v_1725 = v_1722 & v_1084;
assign v_1727 = v_1726 & v_345 & v_346;
assign v_1728 = v_1726 & v_345 & ~v_346 & v_348;
assign v_1729 = v_1726 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_1730 = v_1726 & v_356 & v_357;
assign v_1731 = v_1726 & v_359 & v_360;
assign v_1732 = v_1726 & v_359 & ~v_360 & v_362;
assign v_1733 = v_1726 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_1734 = v_1726 & v_1096;
assign v_1736 = v_1735 & v_1099;
assign v_1738 = v_1737 & v_356 & ~v_357 & v_369 & v_370;
assign v_1739 = v_1737 & v_372 & v_373;
assign v_1740 = v_1737 & v_372 & ~v_373 & v_375;
assign v_1741 = v_1737 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_1743 = v_1737 & v_1742;
assign v_1744 = v_7318 & v_7319;
assign v_1746 = v_1745 & v_384 & v_385;
assign v_1747 = v_1745 & v_384 & ~v_385;
assign v_1749 = v_1748 & v_1113;
assign v_1751 = v_7320 & v_7321;
assign v_1752 = v_1750 & v_391 & v_392;
assign v_1753 = v_1750 & v_391 & ~v_392 & v_394;
assign v_1754 = v_1750 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_1755 = v_1750 & v_1120;
assign v_1757 = v_7322 & v_7323;
assign v_1759 = v_1758 & v_1125;
assign v_1761 = v_1760 & v_410 & v_411;
assign v_1762 = v_1760 & v_410 & ~v_411 & v_413;
assign v_1763 = v_1760 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_1764 = v_1760 & v_421 & v_422;
assign v_1765 = v_1760 & v_424 & v_425;
assign v_1766 = v_1760 & v_424 & ~v_425 & v_427;
assign v_1767 = v_1760 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_1768 = v_1760 & v_1135;
assign v_1770 = v_1769 & v_1138;
assign v_1772 = v_1771 & v_421 & ~v_422 & v_434 & v_435;
assign v_1773 = v_1771 & v_437 & v_438;
assign v_1774 = v_1771 & v_437 & ~v_438 & v_440;
assign v_1775 = v_1771 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_1777 = v_1771 & v_1776;
assign v_1778 = v_7324 & v_7325;
assign v_1780 = v_1779 & v_449 & v_450;
assign v_1781 = v_1779 & v_449 & ~v_450;
assign v_1783 = v_1782 & v_1152;
assign v_1785 = v_7326 & v_7327;
assign v_1786 = v_1784 & v_456 & v_457;
assign v_1787 = v_1784 & v_456 & ~v_457 & v_459;
assign v_1788 = v_1784 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_1789 = v_1784 & v_1159;
assign v_1791 = v_7328 & v_7329;
assign v_1793 = v_1792 & v_1164;
assign v_1795 = v_1794 & v_491;
assign v_1796 = v_1794 & ~v_491 & v_493 & v_526 & ~v_528;
assign v_1797 = v_1794 & ~v_491 & v_493 & v_526 & v_528;
assign v_1798 = v_1794 & ~v_491 & v_493 & ~v_526;
assign v_1799 = v_1794 & v_494;
assign v_1800 = v_1794 & ~v_494;
assign v_1803 = v_1801 & v_1802;
assign v_1804 = v_1801 & v_1180;
assign v_1805 = v_7330 & v_7331;
assign v_1807 = v_1806 & ~v_491 & ~v_493 & v_524;
assign v_1809 = v_1808 & v_531 & v_532;
assign v_1810 = v_1808 & v_531 & ~v_532;
assign v_1812 = v_1811 & v_546 & v_547;
assign v_1813 = v_1811 & v_546 & ~v_547 & ~v_551;
assign v_1815 = v_1814 & v_546 & ~v_547 & v_551;
assign v_1817 = v_1816 & v_554;
assign v_1819 = v_1818 & v_558 & v_559;
assign v_1820 = v_1818 & v_558 & ~v_559 & v_561;
assign v_1821 = v_1818 & v_1196;
assign v_1824 = v_1822 & v_1823;
assign v_1825 = v_1822 & v_1201;
assign v_1827 = v_1826 & v_588 & ~v_589 & ~v_591;
assign v_1828 = v_1826 & v_593 & ~v_594;
assign v_1829 = v_1826 & v_593 & v_594;
assign v_1830 = v_1826 & v_583;
assign v_1832 = v_1831 & v_604 & v_605;
assign v_1833 = v_1831 & v_604 & ~v_605 & ~v_609;
assign v_1835 = v_1834 & v_604 & ~v_605 & v_609;
assign v_1837 = v_1836 & v_612;
assign v_1839 = v_1838 & v_616 & v_617;
assign v_1840 = v_1838 & v_616 & ~v_617 & v_619;
assign v_1841 = v_1838 & v_1214;
assign v_1844 = v_1842 & v_1843;
assign v_1845 = v_1842 & v_1219;
assign v_1847 = v_2 & v_1846;
assign v_1848 = v_641 & v_1826;
assign v_1849 = v_643 & v_1811;
assign v_1850 = v_645 & v_1811;
assign v_1851 = v_647 & v_1811;
assign v_1852 = v_649 & v_1811;
assign v_1853 = ~v_649 & v_1794;
assign v_1855 = ~v_647 & v_1854;
assign v_1857 = ~v_645 & v_1856;
assign v_1859 = ~v_643 & v_1858;
assign v_1861 = ~v_641 & v_1860;
assign v_1863 = ~v_2 & v_1862;
assign v_1865 = v_1864 & ~v_669;
assign v_1866 = v_7332 & v_7333;
assign v_1867 = v_1864 & v_669 & v_670 & v_672 & v_674;
assign v_1868 = v_7334 & v_7335;
assign v_1870 = v_1869 & v_679 & ~v_680 & v_682;
assign v_1871 = v_1869 & v_689 & ~v_690 & ~v_692;
assign v_1872 = v_1869 & v_694 & ~v_695;
assign v_1873 = v_1869 & v_694 & v_695;
assign v_1874 = v_1869 & v_684;
assign v_1876 = v_1875 & v_1251;
assign v_1878 = v_1877 & v_1254;
assign v_1879 = v_1869 & v_679 & v_680;
assign v_1880 = v_1864 & v_1257;
assign v_1882 = v_1881 & ~v_705;
assign v_1883 = v_1881 & v_710 & v_711;
assign v_1884 = v_1881 & v_710 & ~v_711 & ~v_715;
assign v_1886 = v_1885 & v_710 & ~v_711 & v_715;
assign v_1888 = v_1887 & v_718;
assign v_1890 = v_1889 & v_705 & v_722 & v_723 & ~v_724;
assign v_1892 = v_1889 & v_1891;
assign v_1893 = v_1889 & v_750 & v_751;
assign v_1894 = v_1889 & v_750 & ~v_751;
assign v_1896 = v_1895 & v_763 & v_764;
assign v_1897 = v_1895 & v_763 & ~v_764;
assign v_1899 = v_1898 & v_745 & v_758 & v_771;
assign v_1900 = v_7336 & v_7337;
assign v_1901 = v_1889 & v_779 & v_780;
assign v_1902 = v_1889 & v_779 & ~v_780 & ~v_784;
assign v_1904 = v_1903 & v_779 & ~v_780 & v_784;
assign v_1906 = v_1905 & v_787;
assign v_1908 = v_1907 & v_1278;
assign v_1910 = v_1909 & v_798 & ~v_799 & v_817;
assign v_1911 = v_1909 & v_798 & ~v_799 & ~v_817;
assign v_1912 = v_1909 & ~v_800;
assign v_1913 = v_1909 & v_808 & ~v_809;
assign v_1914 = v_1909 & v_1285;
assign v_1916 = v_1915 & v_798 & v_799 & v_814 & ~v_815;
assign v_1918 = v_1917 & v_821 & ~v_822 & v_840;
assign v_1919 = v_1917 & v_821 & ~v_822 & ~v_840;
assign v_1920 = v_1917 & ~v_823;
assign v_1921 = v_1917 & v_831 & ~v_832;
assign v_1922 = v_1917 & v_1294;
assign v_1924 = v_1923 & v_821 & v_822 & v_837 & ~v_838;
assign v_1926 = v_1925 & v_844 & ~v_845 & v_863;
assign v_1927 = v_1925 & ~v_846;
assign v_1928 = v_1925 & v_854 & ~v_855;
assign v_1929 = v_1925 & v_1302;
assign v_1931 = v_1930 & v_844 & v_845 & v_860 & v_861;
assign v_1932 = v_1925 & v_844 & ~v_845 & ~v_863;
assign v_1933 = v_1930 & v_844 & v_845 & v_860 & ~v_861;
assign v_1936 = v_1934 & v_1935;
assign v_1937 = v_1934 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_1938 = v_1934 & v_867 & v_868 & v_869;
assign v_1939 = v_1934 & v_867 & ~v_868 & ~v_872;
assign v_1941 = v_1940 & v_1315;
assign v_1942 = v_1923 & v_821 & v_822 & v_837 & v_838;
assign v_1943 = v_1915 & v_798 & v_799 & v_814 & v_815;
assign v_1945 = v_1944 & v_879 & ~v_880 & v_898;
assign v_1946 = v_1944 & v_879 & ~v_880 & ~v_898;
assign v_1947 = v_1944 & ~v_881;
assign v_1948 = v_1944 & v_889 & ~v_890;
assign v_1949 = v_1944 & v_1324;
assign v_1951 = v_1950 & v_879 & v_880 & v_895 & ~v_896;
assign v_1953 = v_1952 & v_902 & ~v_903 & v_921;
assign v_1954 = v_1952 & v_902 & ~v_903 & ~v_921;
assign v_1955 = v_1952 & ~v_904;
assign v_1956 = v_1952 & v_912 & ~v_913;
assign v_1957 = v_1952 & v_1333;
assign v_1959 = v_1958 & v_902 & v_903 & v_918 & ~v_919;
assign v_1961 = v_1960 & v_925 & ~v_926 & v_944;
assign v_1962 = v_1960 & ~v_927;
assign v_1963 = v_1960 & v_935 & ~v_936;
assign v_1964 = v_1960 & v_1341;
assign v_1966 = v_1965 & v_925 & v_926 & v_941 & v_942;
assign v_1967 = v_1960 & v_925 & ~v_926 & ~v_944;
assign v_1968 = v_1965 & v_925 & v_926 & v_941 & ~v_942;
assign v_1971 = v_1969 & v_1970;
assign v_1972 = v_1969 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_1973 = v_1969 & v_948 & v_949 & v_950;
assign v_1974 = v_1969 & v_948 & ~v_949 & ~v_953;
assign v_1976 = v_1975 & v_1354;
assign v_1977 = v_1958 & v_902 & v_903 & v_918 & v_919;
assign v_1978 = v_1950 & v_879 & v_880 & v_895 & v_896;
assign v_1980 = v_1979 & v_960 & ~v_961 & v_979;
assign v_1981 = v_1979 & v_960 & ~v_961 & ~v_979;
assign v_1982 = v_1979 & ~v_962;
assign v_1983 = v_1979 & v_970 & ~v_971;
assign v_1984 = v_1979 & v_1363;
assign v_1986 = v_1985 & v_960 & v_961 & v_976 & ~v_977;
assign v_1988 = v_1987 & v_983 & ~v_984 & v_1002;
assign v_1989 = v_1987 & v_983 & ~v_984 & ~v_1002;
assign v_1990 = v_1987 & ~v_985;
assign v_1991 = v_1987 & v_993 & ~v_994;
assign v_1992 = v_1987 & v_1372;
assign v_1994 = v_1993 & v_983 & v_984 & v_999 & ~v_1000;
assign v_1996 = v_1995 & v_1006 & ~v_1007 & v_1025;
assign v_1997 = v_1995 & ~v_1008;
assign v_1998 = v_1995 & v_1016 & ~v_1017;
assign v_1999 = v_1995 & v_1380;
assign v_2001 = v_2000 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_2002 = v_1995 & v_1006 & ~v_1007 & ~v_1025;
assign v_2003 = v_2000 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_2006 = v_2004 & v_2005;
assign v_2007 = v_2004 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_2008 = v_2004 & v_1029 & v_1030 & v_1031;
assign v_2009 = v_2004 & v_1029 & ~v_1030 & ~v_1034;
assign v_2011 = v_2010 & v_1393;
assign v_2012 = v_1993 & v_983 & v_984 & v_999 & v_1000;
assign v_2013 = v_1985 & v_960 & v_961 & v_976 & v_977;
assign v_2015 = v_227;
assign v_2016 = ~v_227 & v_229 & v_262 & ~v_264;
assign v_2017 = ~v_227 & v_229 & v_262 & v_264;
assign v_2018 = ~v_227 & v_229 & ~v_262;
assign v_2021 = v_2020;
assign v_2022 = v_1054;
assign v_2023 = v_7338 & v_7339;
assign v_2025 = v_2024 & ~v_227 & ~v_229 & v_260;
assign v_2027 = v_2026 & v_267 & v_268;
assign v_2028 = v_2026 & v_267 & ~v_268;
assign v_2030 = v_2029 & ~v_279;
assign v_2032 = v_2029 & v_2031;
assign v_2033 = v_2029 & v_279 & v_291 & ~v_292 & v_300;
assign v_2036 = v_2034 & v_2035;
assign v_2037 = v_2034 & v_321 & v_322;
assign v_2038 = v_2034 & v_321 & ~v_322 & v_324;
assign v_2039 = v_2034 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_2040 = v_2034 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_2042 = v_2041 & v_1077;
assign v_2044 = v_2043 & ~v_308 & v_309 & v_329;
assign v_2047 = v_2045 & v_2046;
assign v_2048 = v_2045 & v_1084;
assign v_2050 = v_2049 & v_345 & v_346;
assign v_2051 = v_2049 & v_345 & ~v_346 & v_348;
assign v_2052 = v_2049 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_2053 = v_2049 & v_356 & v_357;
assign v_2054 = v_2049 & v_359 & v_360;
assign v_2055 = v_2049 & v_359 & ~v_360 & v_362;
assign v_2056 = v_2049 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_2057 = v_2049 & v_1096;
assign v_2059 = v_2058 & v_1099;
assign v_2061 = v_2060 & v_356 & ~v_357 & v_369 & v_370;
assign v_2062 = v_2060 & v_372 & v_373;
assign v_2063 = v_2060 & v_372 & ~v_373 & v_375;
assign v_2064 = v_2060 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_2066 = v_2060 & v_2065;
assign v_2067 = v_7340 & v_7341;
assign v_2069 = v_2068 & v_384 & v_385;
assign v_2070 = v_2068 & v_384 & ~v_385;
assign v_2072 = v_2071 & v_1113;
assign v_2074 = v_7342 & v_7343;
assign v_2075 = v_2073 & v_391 & v_392;
assign v_2076 = v_2073 & v_391 & ~v_392 & v_394;
assign v_2077 = v_2073 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_2078 = v_2073 & v_1120;
assign v_2080 = v_7344 & v_7345;
assign v_2082 = v_2081 & v_1125;
assign v_2084 = v_2083 & v_410 & v_411;
assign v_2085 = v_2083 & v_410 & ~v_411 & v_413;
assign v_2086 = v_2083 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_2087 = v_2083 & v_421 & v_422;
assign v_2088 = v_2083 & v_424 & v_425;
assign v_2089 = v_2083 & v_424 & ~v_425 & v_427;
assign v_2090 = v_2083 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_2091 = v_2083 & v_1135;
assign v_2093 = v_2092 & v_1138;
assign v_2095 = v_2094 & v_421 & ~v_422 & v_434 & v_435;
assign v_2096 = v_2094 & v_437 & v_438;
assign v_2097 = v_2094 & v_437 & ~v_438 & v_440;
assign v_2098 = v_2094 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_2100 = v_2094 & v_2099;
assign v_2101 = v_7346 & v_7347;
assign v_2103 = v_2102 & v_449 & v_450;
assign v_2104 = v_2102 & v_449 & ~v_450;
assign v_2106 = v_2105 & v_1152;
assign v_2108 = v_7348 & v_7349;
assign v_2109 = v_2107 & v_456 & v_457;
assign v_2110 = v_2107 & v_456 & ~v_457 & v_459;
assign v_2111 = v_2107 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_2112 = v_2107 & v_1159;
assign v_2114 = v_7350 & v_7351;
assign v_2116 = v_2115 & v_1164;
assign v_2118 = v_2117 & v_491;
assign v_2119 = v_2117 & ~v_491 & v_493 & v_526 & ~v_528;
assign v_2120 = v_2117 & ~v_491 & v_493 & v_526 & v_528;
assign v_2121 = v_2117 & ~v_491 & v_493 & ~v_526;
assign v_2122 = v_2117 & v_494;
assign v_2123 = v_2117 & ~v_494;
assign v_2126 = v_2124 & v_2125;
assign v_2127 = v_2124 & v_1180;
assign v_2128 = v_7352 & v_7353;
assign v_2130 = v_2129 & ~v_491 & ~v_493 & v_524;
assign v_2132 = v_2131 & v_531 & v_532;
assign v_2133 = v_2131 & v_531 & ~v_532;
assign v_2135 = v_2134 & v_546 & v_547;
assign v_2136 = v_2134 & v_546 & ~v_547 & ~v_551;
assign v_2138 = v_2137 & v_546 & ~v_547 & v_551;
assign v_2140 = v_2139 & v_554;
assign v_2142 = v_2141 & v_558 & v_559;
assign v_2143 = v_2141 & v_558 & ~v_559 & v_561;
assign v_2144 = v_2141 & v_1196;
assign v_2147 = v_2145 & v_2146;
assign v_2148 = v_2145 & v_1201;
assign v_2150 = v_2149 & v_588 & ~v_589 & ~v_591;
assign v_2151 = v_2149 & v_593 & ~v_594;
assign v_2152 = v_2149 & v_593 & v_594;
assign v_2153 = v_2149 & v_583;
assign v_2155 = v_2154 & v_604 & v_605;
assign v_2156 = v_2154 & v_604 & ~v_605 & ~v_609;
assign v_2158 = v_2157 & v_604 & ~v_605 & v_609;
assign v_2160 = v_2159 & v_612;
assign v_2162 = v_2161 & v_616 & v_617;
assign v_2163 = v_2161 & v_616 & ~v_617 & v_619;
assign v_2164 = v_2161 & v_1214;
assign v_2167 = v_2165 & v_2166;
assign v_2168 = v_2165 & v_1219;
assign v_2170 = v_2 & v_2169;
assign v_2171 = v_641 & v_2149;
assign v_2172 = v_643 & v_2134;
assign v_2173 = v_645 & v_2134;
assign v_2174 = v_647 & v_2134;
assign v_2175 = v_649 & v_2134;
assign v_2176 = ~v_649 & v_2117;
assign v_2178 = ~v_647 & v_2177;
assign v_2180 = ~v_645 & v_2179;
assign v_2182 = ~v_643 & v_2181;
assign v_2184 = ~v_641 & v_2183;
assign v_2186 = ~v_2 & v_2185;
assign v_2188 = v_2187 & ~v_669;
assign v_2189 = v_7354 & v_7355;
assign v_2190 = v_2187 & v_669 & v_670 & v_672 & v_674;
assign v_2191 = v_7356 & v_7357;
assign v_2193 = v_2192 & v_679 & ~v_680 & v_682;
assign v_2194 = v_2192 & v_689 & ~v_690 & ~v_692;
assign v_2195 = v_2192 & v_694 & ~v_695;
assign v_2196 = v_2192 & v_694 & v_695;
assign v_2197 = v_2192 & v_684;
assign v_2199 = v_2198 & v_1251;
assign v_2201 = v_2200 & v_1254;
assign v_2202 = v_2192 & v_679 & v_680;
assign v_2203 = v_2187 & v_1257;
assign v_2205 = v_2204 & ~v_705;
assign v_2206 = v_2204 & v_710 & v_711;
assign v_2207 = v_2204 & v_710 & ~v_711 & ~v_715;
assign v_2209 = v_2208 & v_710 & ~v_711 & v_715;
assign v_2211 = v_2210 & v_718;
assign v_2213 = v_2212 & v_705 & v_722 & v_723 & ~v_724;
assign v_2215 = v_2212 & v_2214;
assign v_2216 = v_2212 & v_750 & v_751;
assign v_2217 = v_2212 & v_750 & ~v_751;
assign v_2219 = v_2218 & v_763 & v_764;
assign v_2220 = v_2218 & v_763 & ~v_764;
assign v_2222 = v_2221 & v_745 & v_758 & v_771;
assign v_2223 = v_7358 & v_7359;
assign v_2224 = v_2212 & v_779 & v_780;
assign v_2225 = v_2212 & v_779 & ~v_780 & ~v_784;
assign v_2227 = v_2226 & v_779 & ~v_780 & v_784;
assign v_2229 = v_2228 & v_787;
assign v_2231 = v_2230 & v_1278;
assign v_2233 = v_2232 & v_798 & ~v_799 & v_817;
assign v_2234 = v_2232 & v_798 & ~v_799 & ~v_817;
assign v_2235 = v_2232 & ~v_800;
assign v_2236 = v_2232 & v_808 & ~v_809;
assign v_2237 = v_2232 & v_1285;
assign v_2239 = v_2238 & v_798 & v_799 & v_814 & ~v_815;
assign v_2241 = v_2240 & v_821 & ~v_822 & v_840;
assign v_2242 = v_2240 & v_821 & ~v_822 & ~v_840;
assign v_2243 = v_2240 & ~v_823;
assign v_2244 = v_2240 & v_831 & ~v_832;
assign v_2245 = v_2240 & v_1294;
assign v_2247 = v_2246 & v_821 & v_822 & v_837 & ~v_838;
assign v_2249 = v_2248 & v_844 & ~v_845 & v_863;
assign v_2250 = v_2248 & ~v_846;
assign v_2251 = v_2248 & v_854 & ~v_855;
assign v_2252 = v_2248 & v_1302;
assign v_2254 = v_2253 & v_844 & v_845 & v_860 & v_861;
assign v_2255 = v_2248 & v_844 & ~v_845 & ~v_863;
assign v_2256 = v_2253 & v_844 & v_845 & v_860 & ~v_861;
assign v_2259 = v_2257 & v_2258;
assign v_2260 = v_2257 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_2261 = v_2257 & v_867 & v_868 & v_869;
assign v_2262 = v_2257 & v_867 & ~v_868 & ~v_872;
assign v_2264 = v_2263 & v_1315;
assign v_2265 = v_2246 & v_821 & v_822 & v_837 & v_838;
assign v_2266 = v_2238 & v_798 & v_799 & v_814 & v_815;
assign v_2268 = v_2267 & v_879 & ~v_880 & v_898;
assign v_2269 = v_2267 & v_879 & ~v_880 & ~v_898;
assign v_2270 = v_2267 & ~v_881;
assign v_2271 = v_2267 & v_889 & ~v_890;
assign v_2272 = v_2267 & v_1324;
assign v_2274 = v_2273 & v_879 & v_880 & v_895 & ~v_896;
assign v_2276 = v_2275 & v_902 & ~v_903 & v_921;
assign v_2277 = v_2275 & v_902 & ~v_903 & ~v_921;
assign v_2278 = v_2275 & ~v_904;
assign v_2279 = v_2275 & v_912 & ~v_913;
assign v_2280 = v_2275 & v_1333;
assign v_2282 = v_2281 & v_902 & v_903 & v_918 & ~v_919;
assign v_2284 = v_2283 & v_925 & ~v_926 & v_944;
assign v_2285 = v_2283 & ~v_927;
assign v_2286 = v_2283 & v_935 & ~v_936;
assign v_2287 = v_2283 & v_1341;
assign v_2289 = v_2288 & v_925 & v_926 & v_941 & v_942;
assign v_2290 = v_2283 & v_925 & ~v_926 & ~v_944;
assign v_2291 = v_2288 & v_925 & v_926 & v_941 & ~v_942;
assign v_2294 = v_2292 & v_2293;
assign v_2295 = v_2292 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_2296 = v_2292 & v_948 & v_949 & v_950;
assign v_2297 = v_2292 & v_948 & ~v_949 & ~v_953;
assign v_2299 = v_2298 & v_1354;
assign v_2300 = v_2281 & v_902 & v_903 & v_918 & v_919;
assign v_2301 = v_2273 & v_879 & v_880 & v_895 & v_896;
assign v_2303 = v_2302 & v_960 & ~v_961 & v_979;
assign v_2304 = v_2302 & v_960 & ~v_961 & ~v_979;
assign v_2305 = v_2302 & ~v_962;
assign v_2306 = v_2302 & v_970 & ~v_971;
assign v_2307 = v_2302 & v_1363;
assign v_2309 = v_2308 & v_960 & v_961 & v_976 & ~v_977;
assign v_2311 = v_2310 & v_983 & ~v_984 & v_1002;
assign v_2312 = v_2310 & v_983 & ~v_984 & ~v_1002;
assign v_2313 = v_2310 & ~v_985;
assign v_2314 = v_2310 & v_993 & ~v_994;
assign v_2315 = v_2310 & v_1372;
assign v_2317 = v_2316 & v_983 & v_984 & v_999 & ~v_1000;
assign v_2319 = v_2318 & v_1006 & ~v_1007 & v_1025;
assign v_2320 = v_2318 & ~v_1008;
assign v_2321 = v_2318 & v_1016 & ~v_1017;
assign v_2322 = v_2318 & v_1380;
assign v_2324 = v_2323 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_2325 = v_2318 & v_1006 & ~v_1007 & ~v_1025;
assign v_2326 = v_2323 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_2329 = v_2327 & v_2328;
assign v_2330 = v_2327 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_2331 = v_2327 & v_1029 & v_1030 & v_1031;
assign v_2332 = v_2327 & v_1029 & ~v_1030 & ~v_1034;
assign v_2334 = v_2333 & v_1393;
assign v_2335 = v_2316 & v_983 & v_984 & v_999 & v_1000;
assign v_2336 = v_2308 & v_960 & v_961 & v_976 & v_977;
assign v_2339 = v_2338 & v_227;
assign v_2340 = v_2338 & ~v_227 & v_229 & v_262 & ~v_264;
assign v_2341 = v_2338 & ~v_227 & v_229 & v_262 & v_264;
assign v_2342 = v_2338 & ~v_227 & v_229 & ~v_262;
assign v_2343 = v_2338 & v_230;
assign v_2344 = v_2338 & ~v_230;
assign v_2347 = v_2345 & v_2346;
assign v_2348 = v_2345 & v_1054;
assign v_2349 = v_7360 & v_7361;
assign v_2351 = v_2350 & ~v_227 & ~v_229 & v_260;
assign v_2353 = v_2352 & v_267 & v_268;
assign v_2354 = v_2352 & v_267 & ~v_268;
assign v_2356 = v_2355 & ~v_279;
assign v_2358 = v_2355 & v_2357;
assign v_2359 = v_2355 & v_279 & v_291 & ~v_292 & v_300;
assign v_2362 = v_2360 & v_2361;
assign v_2363 = v_2360 & v_321 & v_322;
assign v_2364 = v_2360 & v_321 & ~v_322 & v_324;
assign v_2365 = v_2360 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_2366 = v_2360 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_2368 = v_2367 & v_1077;
assign v_2370 = v_2369 & ~v_308 & v_309 & v_329;
assign v_2373 = v_2371 & v_2372;
assign v_2374 = v_2371 & v_1084;
assign v_2376 = v_2375 & v_345 & v_346;
assign v_2377 = v_2375 & v_345 & ~v_346 & v_348;
assign v_2378 = v_2375 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_2379 = v_2375 & v_356 & v_357;
assign v_2380 = v_2375 & v_359 & v_360;
assign v_2381 = v_2375 & v_359 & ~v_360 & v_362;
assign v_2382 = v_2375 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_2383 = v_2375 & v_1096;
assign v_2385 = v_2384 & v_1099;
assign v_2387 = v_2386 & v_356 & ~v_357 & v_369 & v_370;
assign v_2388 = v_2386 & v_372 & v_373;
assign v_2389 = v_2386 & v_372 & ~v_373 & v_375;
assign v_2390 = v_2386 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_2392 = v_2386 & v_2391;
assign v_2393 = v_7362 & v_7363;
assign v_2395 = v_2394 & v_384 & v_385;
assign v_2396 = v_2394 & v_384 & ~v_385;
assign v_2398 = v_2397 & v_1113;
assign v_2400 = v_7364 & v_7365;
assign v_2401 = v_2399 & v_391 & v_392;
assign v_2402 = v_2399 & v_391 & ~v_392 & v_394;
assign v_2403 = v_2399 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_2404 = v_2399 & v_1120;
assign v_2406 = v_7366 & v_7367;
assign v_2408 = v_2407 & v_1125;
assign v_2410 = v_2409 & v_410 & v_411;
assign v_2411 = v_2409 & v_410 & ~v_411 & v_413;
assign v_2412 = v_2409 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_2413 = v_2409 & v_421 & v_422;
assign v_2414 = v_2409 & v_424 & v_425;
assign v_2415 = v_2409 & v_424 & ~v_425 & v_427;
assign v_2416 = v_2409 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_2417 = v_2409 & v_1135;
assign v_2419 = v_2418 & v_1138;
assign v_2421 = v_2420 & v_421 & ~v_422 & v_434 & v_435;
assign v_2422 = v_2420 & v_437 & v_438;
assign v_2423 = v_2420 & v_437 & ~v_438 & v_440;
assign v_2424 = v_2420 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_2426 = v_2420 & v_2425;
assign v_2427 = v_7368 & v_7369;
assign v_2429 = v_2428 & v_449 & v_450;
assign v_2430 = v_2428 & v_449 & ~v_450;
assign v_2432 = v_2431 & v_1152;
assign v_2434 = v_7370 & v_7371;
assign v_2435 = v_2433 & v_456 & v_457;
assign v_2436 = v_2433 & v_456 & ~v_457 & v_459;
assign v_2437 = v_2433 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_2438 = v_2433 & v_1159;
assign v_2440 = v_7372 & v_7373;
assign v_2442 = v_2441 & v_1164;
assign v_2444 = v_2443 & v_491;
assign v_2445 = v_2443 & ~v_491 & v_493 & v_526 & ~v_528;
assign v_2446 = v_2443 & ~v_491 & v_493 & v_526 & v_528;
assign v_2447 = v_2443 & ~v_491 & v_493 & ~v_526;
assign v_2448 = v_2443 & v_494;
assign v_2449 = v_2443 & ~v_494;
assign v_2452 = v_2450 & v_2451;
assign v_2453 = v_2450 & v_1180;
assign v_2454 = v_7374 & v_7375;
assign v_2456 = v_2455 & ~v_491 & ~v_493 & v_524;
assign v_2458 = v_2457 & v_531 & v_532;
assign v_2459 = v_2457 & v_531 & ~v_532;
assign v_2461 = v_2460 & v_546 & v_547;
assign v_2462 = v_2460 & v_546 & ~v_547 & ~v_551;
assign v_2464 = v_2463 & v_546 & ~v_547 & v_551;
assign v_2466 = v_2465 & v_554;
assign v_2468 = v_2467 & v_558 & v_559;
assign v_2469 = v_2467 & v_558 & ~v_559 & v_561;
assign v_2470 = v_2467 & v_1196;
assign v_2473 = v_2471 & v_2472;
assign v_2474 = v_2471 & v_1201;
assign v_2476 = v_2475 & v_588 & ~v_589 & ~v_591;
assign v_2477 = v_2475 & v_593 & ~v_594;
assign v_2478 = v_2475 & v_593 & v_594;
assign v_2479 = v_2475 & v_583;
assign v_2481 = v_2480 & v_604 & v_605;
assign v_2482 = v_2480 & v_604 & ~v_605 & ~v_609;
assign v_2484 = v_2483 & v_604 & ~v_605 & v_609;
assign v_2486 = v_2485 & v_612;
assign v_2488 = v_2487 & v_616 & v_617;
assign v_2489 = v_2487 & v_616 & ~v_617 & v_619;
assign v_2490 = v_2487 & v_1214;
assign v_2493 = v_2491 & v_2492;
assign v_2494 = v_2491 & v_1219;
assign v_2496 = v_2 & v_2495;
assign v_2497 = v_641 & v_2475;
assign v_2498 = v_643 & v_2460;
assign v_2499 = v_645 & v_2460;
assign v_2500 = v_647 & v_2460;
assign v_2501 = v_649 & v_2460;
assign v_2502 = ~v_649 & v_2443;
assign v_2504 = ~v_647 & v_2503;
assign v_2506 = ~v_645 & v_2505;
assign v_2508 = ~v_643 & v_2507;
assign v_2510 = ~v_641 & v_2509;
assign v_2512 = ~v_2 & v_2511;
assign v_2514 = v_2513 & ~v_669;
assign v_2515 = v_7376 & v_7377;
assign v_2516 = v_2513 & v_669 & v_670 & v_672 & v_674;
assign v_2517 = v_7378 & v_7379;
assign v_2519 = v_2518 & v_679 & ~v_680 & v_682;
assign v_2520 = v_2518 & v_689 & ~v_690 & ~v_692;
assign v_2521 = v_2518 & v_694 & ~v_695;
assign v_2522 = v_2518 & v_694 & v_695;
assign v_2523 = v_2518 & v_684;
assign v_2525 = v_2524 & v_1251;
assign v_2527 = v_2526 & v_1254;
assign v_2528 = v_2518 & v_679 & v_680;
assign v_2529 = v_2513 & v_1257;
assign v_2531 = v_2530 & ~v_705;
assign v_2532 = v_2530 & v_710 & v_711;
assign v_2533 = v_2530 & v_710 & ~v_711 & ~v_715;
assign v_2535 = v_2534 & v_710 & ~v_711 & v_715;
assign v_2537 = v_2536 & v_718;
assign v_2539 = v_2538 & v_705 & v_722 & v_723 & ~v_724;
assign v_2541 = v_2538 & v_2540;
assign v_2542 = v_2538 & v_750 & v_751;
assign v_2543 = v_2538 & v_750 & ~v_751;
assign v_2545 = v_2544 & v_763 & v_764;
assign v_2546 = v_2544 & v_763 & ~v_764;
assign v_2548 = v_2547 & v_745 & v_758 & v_771;
assign v_2549 = v_7380 & v_7381;
assign v_2550 = v_2538 & v_779 & v_780;
assign v_2551 = v_2538 & v_779 & ~v_780 & ~v_784;
assign v_2553 = v_2552 & v_779 & ~v_780 & v_784;
assign v_2555 = v_2554 & v_787;
assign v_2557 = v_2556 & v_1278;
assign v_2559 = v_2558 & v_798 & ~v_799 & v_817;
assign v_2560 = v_2558 & v_798 & ~v_799 & ~v_817;
assign v_2561 = v_2558 & ~v_800;
assign v_2562 = v_2558 & v_808 & ~v_809;
assign v_2563 = v_2558 & v_1285;
assign v_2565 = v_2564 & v_798 & v_799 & v_814 & ~v_815;
assign v_2567 = v_2566 & v_821 & ~v_822 & v_840;
assign v_2568 = v_2566 & v_821 & ~v_822 & ~v_840;
assign v_2569 = v_2566 & ~v_823;
assign v_2570 = v_2566 & v_831 & ~v_832;
assign v_2571 = v_2566 & v_1294;
assign v_2573 = v_2572 & v_821 & v_822 & v_837 & ~v_838;
assign v_2575 = v_2574 & v_844 & ~v_845 & v_863;
assign v_2576 = v_2574 & ~v_846;
assign v_2577 = v_2574 & v_854 & ~v_855;
assign v_2578 = v_2574 & v_1302;
assign v_2580 = v_2579 & v_844 & v_845 & v_860 & v_861;
assign v_2581 = v_2574 & v_844 & ~v_845 & ~v_863;
assign v_2582 = v_2579 & v_844 & v_845 & v_860 & ~v_861;
assign v_2585 = v_2583 & v_2584;
assign v_2586 = v_2583 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_2587 = v_2583 & v_867 & v_868 & v_869;
assign v_2588 = v_2583 & v_867 & ~v_868 & ~v_872;
assign v_2590 = v_2589 & v_1315;
assign v_2591 = v_2572 & v_821 & v_822 & v_837 & v_838;
assign v_2592 = v_2564 & v_798 & v_799 & v_814 & v_815;
assign v_2594 = v_2593 & v_879 & ~v_880 & v_898;
assign v_2595 = v_2593 & v_879 & ~v_880 & ~v_898;
assign v_2596 = v_2593 & ~v_881;
assign v_2597 = v_2593 & v_889 & ~v_890;
assign v_2598 = v_2593 & v_1324;
assign v_2600 = v_2599 & v_879 & v_880 & v_895 & ~v_896;
assign v_2602 = v_2601 & v_902 & ~v_903 & v_921;
assign v_2603 = v_2601 & v_902 & ~v_903 & ~v_921;
assign v_2604 = v_2601 & ~v_904;
assign v_2605 = v_2601 & v_912 & ~v_913;
assign v_2606 = v_2601 & v_1333;
assign v_2608 = v_2607 & v_902 & v_903 & v_918 & ~v_919;
assign v_2610 = v_2609 & v_925 & ~v_926 & v_944;
assign v_2611 = v_2609 & ~v_927;
assign v_2612 = v_2609 & v_935 & ~v_936;
assign v_2613 = v_2609 & v_1341;
assign v_2615 = v_2614 & v_925 & v_926 & v_941 & v_942;
assign v_2616 = v_2609 & v_925 & ~v_926 & ~v_944;
assign v_2617 = v_2614 & v_925 & v_926 & v_941 & ~v_942;
assign v_2620 = v_2618 & v_2619;
assign v_2621 = v_2618 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_2622 = v_2618 & v_948 & v_949 & v_950;
assign v_2623 = v_2618 & v_948 & ~v_949 & ~v_953;
assign v_2625 = v_2624 & v_1354;
assign v_2626 = v_2607 & v_902 & v_903 & v_918 & v_919;
assign v_2627 = v_2599 & v_879 & v_880 & v_895 & v_896;
assign v_2629 = v_2628 & v_960 & ~v_961 & v_979;
assign v_2630 = v_2628 & v_960 & ~v_961 & ~v_979;
assign v_2631 = v_2628 & ~v_962;
assign v_2632 = v_2628 & v_970 & ~v_971;
assign v_2633 = v_2628 & v_1363;
assign v_2635 = v_2634 & v_960 & v_961 & v_976 & ~v_977;
assign v_2637 = v_2636 & v_983 & ~v_984 & v_1002;
assign v_2638 = v_2636 & v_983 & ~v_984 & ~v_1002;
assign v_2639 = v_2636 & ~v_985;
assign v_2640 = v_2636 & v_993 & ~v_994;
assign v_2641 = v_2636 & v_1372;
assign v_2643 = v_2642 & v_983 & v_984 & v_999 & ~v_1000;
assign v_2645 = v_2644 & v_1006 & ~v_1007 & v_1025;
assign v_2646 = v_2644 & ~v_1008;
assign v_2647 = v_2644 & v_1016 & ~v_1017;
assign v_2648 = v_2644 & v_1380;
assign v_2650 = v_2649 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_2651 = v_2644 & v_1006 & ~v_1007 & ~v_1025;
assign v_2652 = v_2649 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_2655 = v_2653 & v_2654;
assign v_2656 = v_2653 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_2657 = v_2653 & v_1029 & v_1030 & v_1031;
assign v_2658 = v_2653 & v_1029 & ~v_1030 & ~v_1034;
assign v_2660 = v_2659 & v_1393;
assign v_2661 = v_2642 & v_983 & v_984 & v_999 & v_1000;
assign v_2662 = v_2634 & v_960 & v_961 & v_976 & v_977;
assign v_2665 = v_2664 & v_227;
assign v_2666 = v_2664 & ~v_227 & v_229 & v_262 & ~v_264;
assign v_2667 = v_2664 & ~v_227 & v_229 & v_262 & v_264;
assign v_2668 = v_2664 & ~v_227 & v_229 & ~v_262;
assign v_2669 = v_2664 & v_230;
assign v_2670 = v_2664 & ~v_230;
assign v_2673 = v_2671 & v_2672;
assign v_2674 = v_2671 & v_1054;
assign v_2675 = v_7382 & v_7383;
assign v_2677 = v_2676 & ~v_227 & ~v_229 & v_260;
assign v_2679 = v_2678 & v_267 & v_268;
assign v_2680 = v_2678 & v_267 & ~v_268;
assign v_2682 = v_2681 & ~v_279;
assign v_2684 = v_2681 & v_2683;
assign v_2685 = v_2681 & v_279 & v_291 & ~v_292 & v_300;
assign v_2688 = v_2686 & v_2687;
assign v_2689 = v_2686 & v_321 & v_322;
assign v_2690 = v_2686 & v_321 & ~v_322 & v_324;
assign v_2691 = v_2686 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_2692 = v_2686 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_2694 = v_2693 & v_1077;
assign v_2696 = v_2695 & ~v_308 & v_309 & v_329;
assign v_2699 = v_2697 & v_2698;
assign v_2700 = v_2697 & v_1084;
assign v_2702 = v_2701 & v_345 & v_346;
assign v_2703 = v_2701 & v_345 & ~v_346 & v_348;
assign v_2704 = v_2701 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_2705 = v_2701 & v_356 & v_357;
assign v_2706 = v_2701 & v_359 & v_360;
assign v_2707 = v_2701 & v_359 & ~v_360 & v_362;
assign v_2708 = v_2701 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_2709 = v_2701 & v_1096;
assign v_2711 = v_2710 & v_1099;
assign v_2713 = v_2712 & v_356 & ~v_357 & v_369 & v_370;
assign v_2714 = v_2712 & v_372 & v_373;
assign v_2715 = v_2712 & v_372 & ~v_373 & v_375;
assign v_2716 = v_2712 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_2718 = v_2712 & v_2717;
assign v_2719 = v_7384 & v_7385;
assign v_2721 = v_2720 & v_384 & v_385;
assign v_2722 = v_2720 & v_384 & ~v_385;
assign v_2724 = v_2723 & v_1113;
assign v_2726 = v_7386 & v_7387;
assign v_2727 = v_2725 & v_391 & v_392;
assign v_2728 = v_2725 & v_391 & ~v_392 & v_394;
assign v_2729 = v_2725 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_2730 = v_2725 & v_1120;
assign v_2732 = v_7388 & v_7389;
assign v_2734 = v_2733 & v_1125;
assign v_2736 = v_2735 & v_410 & v_411;
assign v_2737 = v_2735 & v_410 & ~v_411 & v_413;
assign v_2738 = v_2735 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_2739 = v_2735 & v_421 & v_422;
assign v_2740 = v_2735 & v_424 & v_425;
assign v_2741 = v_2735 & v_424 & ~v_425 & v_427;
assign v_2742 = v_2735 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_2743 = v_2735 & v_1135;
assign v_2745 = v_2744 & v_1138;
assign v_2747 = v_2746 & v_421 & ~v_422 & v_434 & v_435;
assign v_2748 = v_2746 & v_437 & v_438;
assign v_2749 = v_2746 & v_437 & ~v_438 & v_440;
assign v_2750 = v_2746 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_2752 = v_2746 & v_2751;
assign v_2753 = v_7390 & v_7391;
assign v_2755 = v_2754 & v_449 & v_450;
assign v_2756 = v_2754 & v_449 & ~v_450;
assign v_2758 = v_2757 & v_1152;
assign v_2760 = v_7392 & v_7393;
assign v_2761 = v_2759 & v_456 & v_457;
assign v_2762 = v_2759 & v_456 & ~v_457 & v_459;
assign v_2763 = v_2759 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_2764 = v_2759 & v_1159;
assign v_2766 = v_7394 & v_7395;
assign v_2768 = v_2767 & v_1164;
assign v_2770 = v_2769 & v_491;
assign v_2771 = v_2769 & ~v_491 & v_493 & v_526 & ~v_528;
assign v_2772 = v_2769 & ~v_491 & v_493 & v_526 & v_528;
assign v_2773 = v_2769 & ~v_491 & v_493 & ~v_526;
assign v_2774 = v_2769 & v_494;
assign v_2775 = v_2769 & ~v_494;
assign v_2778 = v_2776 & v_2777;
assign v_2779 = v_2776 & v_1180;
assign v_2780 = v_7396 & v_7397;
assign v_2782 = v_2781 & ~v_491 & ~v_493 & v_524;
assign v_2784 = v_2783 & v_531 & v_532;
assign v_2785 = v_2783 & v_531 & ~v_532;
assign v_2787 = v_2786 & v_546 & v_547;
assign v_2788 = v_2786 & v_546 & ~v_547 & ~v_551;
assign v_2790 = v_2789 & v_546 & ~v_547 & v_551;
assign v_2792 = v_2791 & v_554;
assign v_2794 = v_2793 & v_558 & v_559;
assign v_2795 = v_2793 & v_558 & ~v_559 & v_561;
assign v_2796 = v_2793 & v_1196;
assign v_2799 = v_2797 & v_2798;
assign v_2800 = v_2797 & v_1201;
assign v_2802 = v_2801 & v_588 & ~v_589 & ~v_591;
assign v_2803 = v_2801 & v_593 & ~v_594;
assign v_2804 = v_2801 & v_593 & v_594;
assign v_2805 = v_2801 & v_583;
assign v_2807 = v_2806 & v_604 & v_605;
assign v_2808 = v_2806 & v_604 & ~v_605 & ~v_609;
assign v_2810 = v_2809 & v_604 & ~v_605 & v_609;
assign v_2812 = v_2811 & v_612;
assign v_2814 = v_2813 & v_616 & v_617;
assign v_2815 = v_2813 & v_616 & ~v_617 & v_619;
assign v_2816 = v_2813 & v_1214;
assign v_2819 = v_2817 & v_2818;
assign v_2820 = v_2817 & v_1219;
assign v_2822 = v_2 & v_2821;
assign v_2823 = v_641 & v_2801;
assign v_2824 = v_643 & v_2786;
assign v_2825 = v_645 & v_2786;
assign v_2826 = v_647 & v_2786;
assign v_2827 = v_649 & v_2786;
assign v_2828 = ~v_649 & v_2769;
assign v_2830 = ~v_647 & v_2829;
assign v_2832 = ~v_645 & v_2831;
assign v_2834 = ~v_643 & v_2833;
assign v_2836 = ~v_641 & v_2835;
assign v_2838 = ~v_2 & v_2837;
assign v_2840 = v_2839 & ~v_669;
assign v_2841 = v_7398 & v_7399;
assign v_2842 = v_2839 & v_669 & v_670 & v_672 & v_674;
assign v_2843 = v_7400 & v_7401;
assign v_2845 = v_2844 & v_679 & ~v_680 & v_682;
assign v_2846 = v_2844 & v_689 & ~v_690 & ~v_692;
assign v_2847 = v_2844 & v_694 & ~v_695;
assign v_2848 = v_2844 & v_694 & v_695;
assign v_2849 = v_2844 & v_684;
assign v_2851 = v_2850 & v_1251;
assign v_2853 = v_2852 & v_1254;
assign v_2854 = v_2844 & v_679 & v_680;
assign v_2855 = v_2839 & v_1257;
assign v_2857 = v_2856 & ~v_705;
assign v_2858 = v_2856 & v_710 & v_711;
assign v_2859 = v_2856 & v_710 & ~v_711 & ~v_715;
assign v_2861 = v_2860 & v_710 & ~v_711 & v_715;
assign v_2863 = v_2862 & v_718;
assign v_2865 = v_2864 & v_705 & v_722 & v_723 & ~v_724;
assign v_2867 = v_2864 & v_2866;
assign v_2868 = v_2864 & v_750 & v_751;
assign v_2869 = v_2864 & v_750 & ~v_751;
assign v_2871 = v_2870 & v_763 & v_764;
assign v_2872 = v_2870 & v_763 & ~v_764;
assign v_2874 = v_2873 & v_745 & v_758 & v_771;
assign v_2875 = v_7402 & v_7403;
assign v_2876 = v_2864 & v_779 & v_780;
assign v_2877 = v_2864 & v_779 & ~v_780 & ~v_784;
assign v_2879 = v_2878 & v_779 & ~v_780 & v_784;
assign v_2881 = v_2880 & v_787;
assign v_2883 = v_2882 & v_1278;
assign v_2885 = v_2884 & v_798 & ~v_799 & v_817;
assign v_2886 = v_2884 & v_798 & ~v_799 & ~v_817;
assign v_2887 = v_2884 & ~v_800;
assign v_2888 = v_2884 & v_808 & ~v_809;
assign v_2889 = v_2884 & v_1285;
assign v_2891 = v_2890 & v_798 & v_799 & v_814 & ~v_815;
assign v_2893 = v_2892 & v_821 & ~v_822 & v_840;
assign v_2894 = v_2892 & v_821 & ~v_822 & ~v_840;
assign v_2895 = v_2892 & ~v_823;
assign v_2896 = v_2892 & v_831 & ~v_832;
assign v_2897 = v_2892 & v_1294;
assign v_2899 = v_2898 & v_821 & v_822 & v_837 & ~v_838;
assign v_2901 = v_2900 & v_844 & ~v_845 & v_863;
assign v_2902 = v_2900 & ~v_846;
assign v_2903 = v_2900 & v_854 & ~v_855;
assign v_2904 = v_2900 & v_1302;
assign v_2906 = v_2905 & v_844 & v_845 & v_860 & v_861;
assign v_2907 = v_2900 & v_844 & ~v_845 & ~v_863;
assign v_2908 = v_2905 & v_844 & v_845 & v_860 & ~v_861;
assign v_2911 = v_2909 & v_2910;
assign v_2912 = v_2909 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_2913 = v_2909 & v_867 & v_868 & v_869;
assign v_2914 = v_2909 & v_867 & ~v_868 & ~v_872;
assign v_2916 = v_2915 & v_1315;
assign v_2917 = v_2898 & v_821 & v_822 & v_837 & v_838;
assign v_2918 = v_2890 & v_798 & v_799 & v_814 & v_815;
assign v_2920 = v_2919 & v_879 & ~v_880 & v_898;
assign v_2921 = v_2919 & v_879 & ~v_880 & ~v_898;
assign v_2922 = v_2919 & ~v_881;
assign v_2923 = v_2919 & v_889 & ~v_890;
assign v_2924 = v_2919 & v_1324;
assign v_2926 = v_2925 & v_879 & v_880 & v_895 & ~v_896;
assign v_2928 = v_2927 & v_902 & ~v_903 & v_921;
assign v_2929 = v_2927 & v_902 & ~v_903 & ~v_921;
assign v_2930 = v_2927 & ~v_904;
assign v_2931 = v_2927 & v_912 & ~v_913;
assign v_2932 = v_2927 & v_1333;
assign v_2934 = v_2933 & v_902 & v_903 & v_918 & ~v_919;
assign v_2936 = v_2935 & v_925 & ~v_926 & v_944;
assign v_2937 = v_2935 & ~v_927;
assign v_2938 = v_2935 & v_935 & ~v_936;
assign v_2939 = v_2935 & v_1341;
assign v_2941 = v_2940 & v_925 & v_926 & v_941 & v_942;
assign v_2942 = v_2935 & v_925 & ~v_926 & ~v_944;
assign v_2943 = v_2940 & v_925 & v_926 & v_941 & ~v_942;
assign v_2946 = v_2944 & v_2945;
assign v_2947 = v_2944 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_2948 = v_2944 & v_948 & v_949 & v_950;
assign v_2949 = v_2944 & v_948 & ~v_949 & ~v_953;
assign v_2951 = v_2950 & v_1354;
assign v_2952 = v_2933 & v_902 & v_903 & v_918 & v_919;
assign v_2953 = v_2925 & v_879 & v_880 & v_895 & v_896;
assign v_2955 = v_2954 & v_960 & ~v_961 & v_979;
assign v_2956 = v_2954 & v_960 & ~v_961 & ~v_979;
assign v_2957 = v_2954 & ~v_962;
assign v_2958 = v_2954 & v_970 & ~v_971;
assign v_2959 = v_2954 & v_1363;
assign v_2961 = v_2960 & v_960 & v_961 & v_976 & ~v_977;
assign v_2963 = v_2962 & v_983 & ~v_984 & v_1002;
assign v_2964 = v_2962 & v_983 & ~v_984 & ~v_1002;
assign v_2965 = v_2962 & ~v_985;
assign v_2966 = v_2962 & v_993 & ~v_994;
assign v_2967 = v_2962 & v_1372;
assign v_2969 = v_2968 & v_983 & v_984 & v_999 & ~v_1000;
assign v_2971 = v_2970 & v_1006 & ~v_1007 & v_1025;
assign v_2972 = v_2970 & ~v_1008;
assign v_2973 = v_2970 & v_1016 & ~v_1017;
assign v_2974 = v_2970 & v_1380;
assign v_2976 = v_2975 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_2977 = v_2970 & v_1006 & ~v_1007 & ~v_1025;
assign v_2978 = v_2975 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_2981 = v_2979 & v_2980;
assign v_2982 = v_2979 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_2983 = v_2979 & v_1029 & v_1030 & v_1031;
assign v_2984 = v_2979 & v_1029 & ~v_1030 & ~v_1034;
assign v_2986 = v_2985 & v_1393;
assign v_2987 = v_2968 & v_983 & v_984 & v_999 & v_1000;
assign v_2988 = v_2960 & v_960 & v_961 & v_976 & v_977;
assign v_2990 = v_7 & v_227;
assign v_2991 = v_7 & ~v_227 & v_229 & v_262 & ~v_264;
assign v_2992 = v_7 & ~v_227 & v_229 & v_262 & v_264;
assign v_2993 = v_7 & ~v_227 & v_229 & ~v_262;
assign v_2994 = v_7 & v_230;
assign v_2995 = v_7 & ~v_230;
assign v_2998 = v_2996 & v_2997;
assign v_2999 = v_2996 & v_1054;
assign v_3000 = v_7404 & v_7405;
assign v_3002 = v_3001 & ~v_227 & ~v_229 & v_260;
assign v_3004 = v_3003 & v_267 & v_268;
assign v_3005 = v_3003 & v_267 & ~v_268;
assign v_3007 = v_3006 & ~v_279;
assign v_3009 = v_3006 & v_3008;
assign v_3010 = v_3006 & v_279 & v_291 & ~v_292 & v_300;
assign v_3013 = v_3011 & v_3012;
assign v_3014 = v_3011 & v_321 & v_322;
assign v_3015 = v_3011 & v_321 & ~v_322 & v_324;
assign v_3016 = v_3011 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_3017 = v_3011 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_3019 = v_3018 & v_1077;
assign v_3021 = v_3020 & ~v_308 & v_309 & v_329;
assign v_3024 = v_3022 & v_3023;
assign v_3025 = v_3022 & v_1084;
assign v_3027 = v_3026 & v_345 & v_346;
assign v_3028 = v_3026 & v_345 & ~v_346 & v_348;
assign v_3029 = v_3026 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_3030 = v_3026 & v_356 & v_357;
assign v_3031 = v_3026 & v_359 & v_360;
assign v_3032 = v_3026 & v_359 & ~v_360 & v_362;
assign v_3033 = v_3026 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_3034 = v_3026 & v_1096;
assign v_3036 = v_3035 & v_1099;
assign v_3038 = v_3037 & v_356 & ~v_357 & v_369 & v_370;
assign v_3039 = v_3037 & v_372 & v_373;
assign v_3040 = v_3037 & v_372 & ~v_373 & v_375;
assign v_3041 = v_3037 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_3043 = v_3037 & v_3042;
assign v_3044 = v_7406 & v_7407;
assign v_3046 = v_3045 & v_384 & v_385;
assign v_3047 = v_3045 & v_384 & ~v_385;
assign v_3049 = v_3048 & v_1113;
assign v_3051 = v_7408 & v_7409;
assign v_3052 = v_3050 & v_391 & v_392;
assign v_3053 = v_3050 & v_391 & ~v_392 & v_394;
assign v_3054 = v_3050 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_3055 = v_3050 & v_1120;
assign v_3057 = v_7410 & v_7411;
assign v_3059 = v_3058 & v_1125;
assign v_3061 = v_3060 & v_410 & v_411;
assign v_3062 = v_3060 & v_410 & ~v_411 & v_413;
assign v_3063 = v_3060 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_3064 = v_3060 & v_421 & v_422;
assign v_3065 = v_3060 & v_424 & v_425;
assign v_3066 = v_3060 & v_424 & ~v_425 & v_427;
assign v_3067 = v_3060 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_3068 = v_3060 & v_1135;
assign v_3070 = v_3069 & v_1138;
assign v_3072 = v_3071 & v_421 & ~v_422 & v_434 & v_435;
assign v_3073 = v_3071 & v_437 & v_438;
assign v_3074 = v_3071 & v_437 & ~v_438 & v_440;
assign v_3075 = v_3071 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_3077 = v_3071 & v_3076;
assign v_3078 = v_7412 & v_7413;
assign v_3080 = v_3079 & v_449 & v_450;
assign v_3081 = v_3079 & v_449 & ~v_450;
assign v_3083 = v_3082 & v_1152;
assign v_3085 = v_7414 & v_7415;
assign v_3086 = v_3084 & v_456 & v_457;
assign v_3087 = v_3084 & v_456 & ~v_457 & v_459;
assign v_3088 = v_3084 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_3089 = v_3084 & v_1159;
assign v_3091 = v_7416 & v_7417;
assign v_3093 = v_3092 & v_1164;
assign v_3095 = v_3094 & v_491;
assign v_3096 = v_3094 & ~v_491 & v_493 & v_526 & ~v_528;
assign v_3097 = v_3094 & ~v_491 & v_493 & v_526 & v_528;
assign v_3098 = v_3094 & ~v_491 & v_493 & ~v_526;
assign v_3099 = v_3094 & v_494;
assign v_3100 = v_3094 & ~v_494;
assign v_3103 = v_3101 & v_3102;
assign v_3104 = v_3101 & v_1180;
assign v_3105 = v_7418 & v_7419;
assign v_3107 = v_3106 & ~v_491 & ~v_493 & v_524;
assign v_3109 = v_3108 & v_531 & v_532;
assign v_3110 = v_3108 & v_531 & ~v_532;
assign v_3112 = v_3111 & v_546 & v_547;
assign v_3113 = v_3111 & v_546 & ~v_547 & ~v_551;
assign v_3115 = v_3114 & v_546 & ~v_547 & v_551;
assign v_3117 = v_3116 & v_554;
assign v_3119 = v_3118 & v_558 & v_559;
assign v_3120 = v_3118 & v_558 & ~v_559 & v_561;
assign v_3121 = v_3118 & v_1196;
assign v_3124 = v_3122 & v_3123;
assign v_3125 = v_3122 & v_1201;
assign v_3127 = v_3126 & v_588 & ~v_589 & ~v_591;
assign v_3128 = v_3126 & v_593 & ~v_594;
assign v_3129 = v_3126 & v_593 & v_594;
assign v_3130 = v_3126 & v_583;
assign v_3132 = v_3131 & v_604 & v_605;
assign v_3133 = v_3131 & v_604 & ~v_605 & ~v_609;
assign v_3135 = v_3134 & v_604 & ~v_605 & v_609;
assign v_3137 = v_3136 & v_612;
assign v_3139 = v_3138 & v_616 & v_617;
assign v_3140 = v_3138 & v_616 & ~v_617 & v_619;
assign v_3141 = v_3138 & v_1214;
assign v_3144 = v_3142 & v_3143;
assign v_3145 = v_3142 & v_1219;
assign v_3147 = v_2 & v_3146;
assign v_3148 = v_641 & v_3126;
assign v_3149 = v_643 & v_3111;
assign v_3150 = v_645 & v_3111;
assign v_3151 = v_647 & v_3111;
assign v_3152 = v_649 & v_3111;
assign v_3153 = ~v_649 & v_3094;
assign v_3155 = ~v_647 & v_3154;
assign v_3157 = ~v_645 & v_3156;
assign v_3159 = ~v_643 & v_3158;
assign v_3161 = ~v_641 & v_3160;
assign v_3163 = ~v_2 & v_3162;
assign v_3165 = v_3164 & ~v_669;
assign v_3166 = v_7420 & v_7421;
assign v_3167 = v_3164 & v_669 & v_670 & v_672 & v_674;
assign v_3168 = v_7422 & v_7423;
assign v_3170 = v_3169 & v_679 & ~v_680 & v_682;
assign v_3171 = v_3169 & v_689 & ~v_690 & ~v_692;
assign v_3172 = v_3169 & v_694 & ~v_695;
assign v_3173 = v_3169 & v_694 & v_695;
assign v_3174 = v_3169 & v_684;
assign v_3176 = v_3175 & v_1251;
assign v_3178 = v_3177 & v_1254;
assign v_3179 = v_3169 & v_679 & v_680;
assign v_3180 = v_3164 & v_1257;
assign v_3182 = v_3181 & ~v_705;
assign v_3183 = v_3181 & v_710 & v_711;
assign v_3184 = v_3181 & v_710 & ~v_711 & ~v_715;
assign v_3186 = v_3185 & v_710 & ~v_711 & v_715;
assign v_3188 = v_3187 & v_718;
assign v_3190 = v_3189 & v_705 & v_722 & v_723 & ~v_724;
assign v_3192 = v_3189 & v_3191;
assign v_3193 = v_3189 & v_750 & v_751;
assign v_3194 = v_3189 & v_750 & ~v_751;
assign v_3196 = v_3195 & v_763 & v_764;
assign v_3197 = v_3195 & v_763 & ~v_764;
assign v_3199 = v_3198 & v_745 & v_758 & v_771;
assign v_3200 = v_7424 & v_7425;
assign v_3201 = v_3189 & v_779 & v_780;
assign v_3202 = v_3189 & v_779 & ~v_780 & ~v_784;
assign v_3204 = v_3203 & v_779 & ~v_780 & v_784;
assign v_3206 = v_3205 & v_787;
assign v_3208 = v_3207 & v_1278;
assign v_3210 = v_3209 & v_798 & ~v_799 & v_817;
assign v_3211 = v_3209 & v_798 & ~v_799 & ~v_817;
assign v_3212 = v_3209 & ~v_800;
assign v_3213 = v_3209 & v_808 & ~v_809;
assign v_3214 = v_3209 & v_1285;
assign v_3216 = v_3215 & v_798 & v_799 & v_814 & ~v_815;
assign v_3218 = v_3217 & v_821 & ~v_822 & v_840;
assign v_3219 = v_3217 & v_821 & ~v_822 & ~v_840;
assign v_3220 = v_3217 & ~v_823;
assign v_3221 = v_3217 & v_831 & ~v_832;
assign v_3222 = v_3217 & v_1294;
assign v_3224 = v_3223 & v_821 & v_822 & v_837 & ~v_838;
assign v_3226 = v_3225 & v_844 & ~v_845 & v_863;
assign v_3227 = v_3225 & ~v_846;
assign v_3228 = v_3225 & v_854 & ~v_855;
assign v_3229 = v_3225 & v_1302;
assign v_3231 = v_3230 & v_844 & v_845 & v_860 & v_861;
assign v_3232 = v_3225 & v_844 & ~v_845 & ~v_863;
assign v_3233 = v_3230 & v_844 & v_845 & v_860 & ~v_861;
assign v_3236 = v_3234 & v_3235;
assign v_3237 = v_3234 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_3238 = v_3234 & v_867 & v_868 & v_869;
assign v_3239 = v_3234 & v_867 & ~v_868 & ~v_872;
assign v_3241 = v_3240 & v_1315;
assign v_3242 = v_3223 & v_821 & v_822 & v_837 & v_838;
assign v_3243 = v_3215 & v_798 & v_799 & v_814 & v_815;
assign v_3245 = v_3244 & v_879 & ~v_880 & v_898;
assign v_3246 = v_3244 & v_879 & ~v_880 & ~v_898;
assign v_3247 = v_3244 & ~v_881;
assign v_3248 = v_3244 & v_889 & ~v_890;
assign v_3249 = v_3244 & v_1324;
assign v_3251 = v_3250 & v_879 & v_880 & v_895 & ~v_896;
assign v_3253 = v_3252 & v_902 & ~v_903 & v_921;
assign v_3254 = v_3252 & v_902 & ~v_903 & ~v_921;
assign v_3255 = v_3252 & ~v_904;
assign v_3256 = v_3252 & v_912 & ~v_913;
assign v_3257 = v_3252 & v_1333;
assign v_3259 = v_3258 & v_902 & v_903 & v_918 & ~v_919;
assign v_3261 = v_3260 & v_925 & ~v_926 & v_944;
assign v_3262 = v_3260 & ~v_927;
assign v_3263 = v_3260 & v_935 & ~v_936;
assign v_3264 = v_3260 & v_1341;
assign v_3266 = v_3265 & v_925 & v_926 & v_941 & v_942;
assign v_3267 = v_3260 & v_925 & ~v_926 & ~v_944;
assign v_3268 = v_3265 & v_925 & v_926 & v_941 & ~v_942;
assign v_3271 = v_3269 & v_3270;
assign v_3272 = v_3269 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_3273 = v_3269 & v_948 & v_949 & v_950;
assign v_3274 = v_3269 & v_948 & ~v_949 & ~v_953;
assign v_3276 = v_3275 & v_1354;
assign v_3277 = v_3258 & v_902 & v_903 & v_918 & v_919;
assign v_3278 = v_3250 & v_879 & v_880 & v_895 & v_896;
assign v_3280 = v_3279 & v_960 & ~v_961 & v_979;
assign v_3281 = v_3279 & v_960 & ~v_961 & ~v_979;
assign v_3282 = v_3279 & ~v_962;
assign v_3283 = v_3279 & v_970 & ~v_971;
assign v_3284 = v_3279 & v_1363;
assign v_3286 = v_3285 & v_960 & v_961 & v_976 & ~v_977;
assign v_3288 = v_3287 & v_983 & ~v_984 & v_1002;
assign v_3289 = v_3287 & v_983 & ~v_984 & ~v_1002;
assign v_3290 = v_3287 & ~v_985;
assign v_3291 = v_3287 & v_993 & ~v_994;
assign v_3292 = v_3287 & v_1372;
assign v_3294 = v_3293 & v_983 & v_984 & v_999 & ~v_1000;
assign v_3296 = v_3295 & v_1006 & ~v_1007 & v_1025;
assign v_3297 = v_3295 & ~v_1008;
assign v_3298 = v_3295 & v_1016 & ~v_1017;
assign v_3299 = v_3295 & v_1380;
assign v_3301 = v_3300 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_3302 = v_3295 & v_1006 & ~v_1007 & ~v_1025;
assign v_3303 = v_3300 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_3306 = v_3304 & v_3305;
assign v_3307 = v_3304 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_3308 = v_3304 & v_1029 & v_1030 & v_1031;
assign v_3309 = v_3304 & v_1029 & ~v_1030 & ~v_1034;
assign v_3311 = v_3310 & v_1393;
assign v_3312 = v_3293 & v_983 & v_984 & v_999 & v_1000;
assign v_3313 = v_3285 & v_960 & v_961 & v_976 & v_977;
assign v_3316 = v_3315 & v_227;
assign v_3317 = v_3315 & ~v_227 & v_229 & v_262 & ~v_264;
assign v_3318 = v_3315 & ~v_227 & v_229 & v_262 & v_264;
assign v_3319 = v_3315 & ~v_227 & v_229 & ~v_262;
assign v_3320 = v_3315 & v_230;
assign v_3321 = v_3315 & ~v_230;
assign v_3324 = v_3322 & v_3323;
assign v_3325 = v_3322 & v_1054;
assign v_3326 = v_7426 & v_7427;
assign v_3328 = v_3327 & ~v_227 & ~v_229 & v_260;
assign v_3330 = v_3329 & v_267 & v_268;
assign v_3331 = v_3329 & v_267 & ~v_268;
assign v_3333 = v_3332 & ~v_279;
assign v_3335 = v_3332 & v_3334;
assign v_3336 = v_3332 & v_279 & v_291 & ~v_292 & v_300;
assign v_3339 = v_3337 & v_3338;
assign v_3340 = v_3337 & v_321 & v_322;
assign v_3341 = v_3337 & v_321 & ~v_322 & v_324;
assign v_3342 = v_3337 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_3343 = v_3337 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_3345 = v_3344 & v_1077;
assign v_3347 = v_3346 & ~v_308 & v_309 & v_329;
assign v_3350 = v_3348 & v_3349;
assign v_3351 = v_3348 & v_1084;
assign v_3353 = v_3352 & v_345 & v_346;
assign v_3354 = v_3352 & v_345 & ~v_346 & v_348;
assign v_3355 = v_3352 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_3356 = v_3352 & v_356 & v_357;
assign v_3357 = v_3352 & v_359 & v_360;
assign v_3358 = v_3352 & v_359 & ~v_360 & v_362;
assign v_3359 = v_3352 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_3360 = v_3352 & v_1096;
assign v_3362 = v_3361 & v_1099;
assign v_3364 = v_3363 & v_356 & ~v_357 & v_369 & v_370;
assign v_3365 = v_3363 & v_372 & v_373;
assign v_3366 = v_3363 & v_372 & ~v_373 & v_375;
assign v_3367 = v_3363 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_3369 = v_3363 & v_3368;
assign v_3370 = v_7428 & v_7429;
assign v_3372 = v_3371 & v_384 & v_385;
assign v_3373 = v_3371 & v_384 & ~v_385;
assign v_3375 = v_3374 & v_1113;
assign v_3377 = v_7430 & v_7431;
assign v_3378 = v_3376 & v_391 & v_392;
assign v_3379 = v_3376 & v_391 & ~v_392 & v_394;
assign v_3380 = v_3376 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_3381 = v_3376 & v_1120;
assign v_3383 = v_7432 & v_7433;
assign v_3385 = v_3384 & v_1125;
assign v_3387 = v_3386 & v_410 & v_411;
assign v_3388 = v_3386 & v_410 & ~v_411 & v_413;
assign v_3389 = v_3386 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_3390 = v_3386 & v_421 & v_422;
assign v_3391 = v_3386 & v_424 & v_425;
assign v_3392 = v_3386 & v_424 & ~v_425 & v_427;
assign v_3393 = v_3386 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_3394 = v_3386 & v_1135;
assign v_3396 = v_3395 & v_1138;
assign v_3398 = v_3397 & v_421 & ~v_422 & v_434 & v_435;
assign v_3399 = v_3397 & v_437 & v_438;
assign v_3400 = v_3397 & v_437 & ~v_438 & v_440;
assign v_3401 = v_3397 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_3403 = v_3397 & v_3402;
assign v_3404 = v_7434 & v_7435;
assign v_3406 = v_3405 & v_449 & v_450;
assign v_3407 = v_3405 & v_449 & ~v_450;
assign v_3409 = v_3408 & v_1152;
assign v_3411 = v_7436 & v_7437;
assign v_3412 = v_3410 & v_456 & v_457;
assign v_3413 = v_3410 & v_456 & ~v_457 & v_459;
assign v_3414 = v_3410 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_3415 = v_3410 & v_1159;
assign v_3417 = v_7438 & v_7439;
assign v_3419 = v_3418 & v_1164;
assign v_3421 = v_3420 & v_491;
assign v_3422 = v_3420 & ~v_491 & v_493 & v_526 & ~v_528;
assign v_3423 = v_3420 & ~v_491 & v_493 & v_526 & v_528;
assign v_3424 = v_3420 & ~v_491 & v_493 & ~v_526;
assign v_3425 = v_3420 & v_494;
assign v_3426 = v_3420 & ~v_494;
assign v_3429 = v_3427 & v_3428;
assign v_3430 = v_3427 & v_1180;
assign v_3431 = v_7440 & v_7441;
assign v_3433 = v_3432 & ~v_491 & ~v_493 & v_524;
assign v_3435 = v_3434 & v_531 & v_532;
assign v_3436 = v_3434 & v_531 & ~v_532;
assign v_3438 = v_3437 & v_546 & v_547;
assign v_3439 = v_3437 & v_546 & ~v_547 & ~v_551;
assign v_3441 = v_3440 & v_546 & ~v_547 & v_551;
assign v_3443 = v_3442 & v_554;
assign v_3445 = v_3444 & v_558 & v_559;
assign v_3446 = v_3444 & v_558 & ~v_559 & v_561;
assign v_3447 = v_3444 & v_1196;
assign v_3450 = v_3448 & v_3449;
assign v_3451 = v_3448 & v_1201;
assign v_3453 = v_3452 & v_588 & ~v_589 & ~v_591;
assign v_3454 = v_3452 & v_593 & ~v_594;
assign v_3455 = v_3452 & v_593 & v_594;
assign v_3456 = v_3452 & v_583;
assign v_3458 = v_3457 & v_604 & v_605;
assign v_3459 = v_3457 & v_604 & ~v_605 & ~v_609;
assign v_3461 = v_3460 & v_604 & ~v_605 & v_609;
assign v_3463 = v_3462 & v_612;
assign v_3465 = v_3464 & v_616 & v_617;
assign v_3466 = v_3464 & v_616 & ~v_617 & v_619;
assign v_3467 = v_3464 & v_1214;
assign v_3470 = v_3468 & v_3469;
assign v_3471 = v_3468 & v_1219;
assign v_3473 = v_2 & v_3472;
assign v_3474 = v_641 & v_3452;
assign v_3475 = v_643 & v_3437;
assign v_3476 = v_645 & v_3437;
assign v_3477 = v_647 & v_3437;
assign v_3478 = v_649 & v_3437;
assign v_3479 = ~v_649 & v_3420;
assign v_3481 = ~v_647 & v_3480;
assign v_3483 = ~v_645 & v_3482;
assign v_3485 = ~v_643 & v_3484;
assign v_3487 = ~v_641 & v_3486;
assign v_3489 = ~v_2 & v_3488;
assign v_3491 = v_3490 & ~v_669;
assign v_3492 = v_7442 & v_7443;
assign v_3493 = v_3490 & v_669 & v_670 & v_672 & v_674;
assign v_3494 = v_7444 & v_7445;
assign v_3496 = v_3495 & v_679 & ~v_680 & v_682;
assign v_3497 = v_3495 & v_689 & ~v_690 & ~v_692;
assign v_3498 = v_3495 & v_694 & ~v_695;
assign v_3499 = v_3495 & v_694 & v_695;
assign v_3500 = v_3495 & v_684;
assign v_3502 = v_3501 & v_1251;
assign v_3504 = v_3503 & v_1254;
assign v_3505 = v_3495 & v_679 & v_680;
assign v_3506 = v_3490 & v_1257;
assign v_3508 = v_3507 & ~v_705;
assign v_3509 = v_3507 & v_710 & v_711;
assign v_3510 = v_3507 & v_710 & ~v_711 & ~v_715;
assign v_3512 = v_3511 & v_710 & ~v_711 & v_715;
assign v_3514 = v_3513 & v_718;
assign v_3516 = v_3515 & v_705 & v_722 & v_723 & ~v_724;
assign v_3518 = v_3515 & v_3517;
assign v_3519 = v_3515 & v_750 & v_751;
assign v_3520 = v_3515 & v_750 & ~v_751;
assign v_3522 = v_3521 & v_763 & v_764;
assign v_3523 = v_3521 & v_763 & ~v_764;
assign v_3525 = v_3524 & v_745 & v_758 & v_771;
assign v_3526 = v_7446 & v_7447;
assign v_3527 = v_3515 & v_779 & v_780;
assign v_3528 = v_3515 & v_779 & ~v_780 & ~v_784;
assign v_3530 = v_3529 & v_779 & ~v_780 & v_784;
assign v_3532 = v_3531 & v_787;
assign v_3534 = v_3533 & v_1278;
assign v_3536 = v_3535 & v_798 & ~v_799 & v_817;
assign v_3537 = v_3535 & v_798 & ~v_799 & ~v_817;
assign v_3538 = v_3535 & ~v_800;
assign v_3539 = v_3535 & v_808 & ~v_809;
assign v_3540 = v_3535 & v_1285;
assign v_3542 = v_3541 & v_798 & v_799 & v_814 & ~v_815;
assign v_3544 = v_3543 & v_821 & ~v_822 & v_840;
assign v_3545 = v_3543 & v_821 & ~v_822 & ~v_840;
assign v_3546 = v_3543 & ~v_823;
assign v_3547 = v_3543 & v_831 & ~v_832;
assign v_3548 = v_3543 & v_1294;
assign v_3550 = v_3549 & v_821 & v_822 & v_837 & ~v_838;
assign v_3552 = v_3551 & v_844 & ~v_845 & v_863;
assign v_3553 = v_3551 & ~v_846;
assign v_3554 = v_3551 & v_854 & ~v_855;
assign v_3555 = v_3551 & v_1302;
assign v_3557 = v_3556 & v_844 & v_845 & v_860 & v_861;
assign v_3558 = v_3551 & v_844 & ~v_845 & ~v_863;
assign v_3559 = v_3556 & v_844 & v_845 & v_860 & ~v_861;
assign v_3562 = v_3560 & v_3561;
assign v_3563 = v_3560 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_3564 = v_3560 & v_867 & v_868 & v_869;
assign v_3565 = v_3560 & v_867 & ~v_868 & ~v_872;
assign v_3567 = v_3566 & v_1315;
assign v_3568 = v_3549 & v_821 & v_822 & v_837 & v_838;
assign v_3569 = v_3541 & v_798 & v_799 & v_814 & v_815;
assign v_3571 = v_3570 & v_879 & ~v_880 & v_898;
assign v_3572 = v_3570 & v_879 & ~v_880 & ~v_898;
assign v_3573 = v_3570 & ~v_881;
assign v_3574 = v_3570 & v_889 & ~v_890;
assign v_3575 = v_3570 & v_1324;
assign v_3577 = v_3576 & v_879 & v_880 & v_895 & ~v_896;
assign v_3579 = v_3578 & v_902 & ~v_903 & v_921;
assign v_3580 = v_3578 & v_902 & ~v_903 & ~v_921;
assign v_3581 = v_3578 & ~v_904;
assign v_3582 = v_3578 & v_912 & ~v_913;
assign v_3583 = v_3578 & v_1333;
assign v_3585 = v_3584 & v_902 & v_903 & v_918 & ~v_919;
assign v_3587 = v_3586 & v_925 & ~v_926 & v_944;
assign v_3588 = v_3586 & ~v_927;
assign v_3589 = v_3586 & v_935 & ~v_936;
assign v_3590 = v_3586 & v_1341;
assign v_3592 = v_3591 & v_925 & v_926 & v_941 & v_942;
assign v_3593 = v_3586 & v_925 & ~v_926 & ~v_944;
assign v_3594 = v_3591 & v_925 & v_926 & v_941 & ~v_942;
assign v_3597 = v_3595 & v_3596;
assign v_3598 = v_3595 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_3599 = v_3595 & v_948 & v_949 & v_950;
assign v_3600 = v_3595 & v_948 & ~v_949 & ~v_953;
assign v_3602 = v_3601 & v_1354;
assign v_3603 = v_3584 & v_902 & v_903 & v_918 & v_919;
assign v_3604 = v_3576 & v_879 & v_880 & v_895 & v_896;
assign v_3606 = v_3605 & v_960 & ~v_961 & v_979;
assign v_3607 = v_3605 & v_960 & ~v_961 & ~v_979;
assign v_3608 = v_3605 & ~v_962;
assign v_3609 = v_3605 & v_970 & ~v_971;
assign v_3610 = v_3605 & v_1363;
assign v_3612 = v_3611 & v_960 & v_961 & v_976 & ~v_977;
assign v_3614 = v_3613 & v_983 & ~v_984 & v_1002;
assign v_3615 = v_3613 & v_983 & ~v_984 & ~v_1002;
assign v_3616 = v_3613 & ~v_985;
assign v_3617 = v_3613 & v_993 & ~v_994;
assign v_3618 = v_3613 & v_1372;
assign v_3620 = v_3619 & v_983 & v_984 & v_999 & ~v_1000;
assign v_3622 = v_3621 & v_1006 & ~v_1007 & v_1025;
assign v_3623 = v_3621 & ~v_1008;
assign v_3624 = v_3621 & v_1016 & ~v_1017;
assign v_3625 = v_3621 & v_1380;
assign v_3627 = v_3626 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_3628 = v_3621 & v_1006 & ~v_1007 & ~v_1025;
assign v_3629 = v_3626 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_3632 = v_3630 & v_3631;
assign v_3633 = v_3630 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_3634 = v_3630 & v_1029 & v_1030 & v_1031;
assign v_3635 = v_3630 & v_1029 & ~v_1030 & ~v_1034;
assign v_3637 = v_3636 & v_1393;
assign v_3638 = v_3619 & v_983 & v_984 & v_999 & v_1000;
assign v_3639 = v_3611 & v_960 & v_961 & v_976 & v_977;
assign v_3642 = v_3641 & ~v_1086;
assign v_3644 = v_1041 & v_3643;
assign v_3645 = v_227;
assign v_3647 = v_3646 & v_267 & v_268;
assign v_3648 = v_3646 & v_267 & ~v_268;
assign v_3650 = v_3649 & ~v_279;
assign v_3652 = v_3649 & v_3651;
assign v_3653 = v_3649 & v_279 & v_291 & ~v_292 & v_300;
assign v_3656 = v_3654 & v_3655;
assign v_3657 = v_3654 & v_321 & v_322;
assign v_3658 = v_3654 & v_321 & ~v_322 & v_324;
assign v_3659 = v_3654 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_3660 = v_3654 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_3662 = v_3661 & v_1077;
assign v_3664 = v_3663 & ~v_308 & v_309 & v_329;
assign v_3667 = v_3665 & v_3666;
assign v_3668 = v_3665 & v_1084;
assign v_3670 = ~v_1041 & v_3669;
assign v_3672 = v_3671 & v_345 & v_346;
assign v_3673 = v_3671 & v_345 & ~v_346 & v_348;
assign v_3674 = v_3671 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_3675 = v_3671 & v_356 & v_357;
assign v_3676 = v_3671 & v_359 & v_360;
assign v_3677 = v_3671 & v_359 & ~v_360 & v_362;
assign v_3678 = v_3671 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_3679 = v_3671 & v_1096;
assign v_3681 = v_3680 & v_1099;
assign v_3683 = v_3682 & v_356 & ~v_357 & v_369 & v_370;
assign v_3684 = v_3682 & v_372 & v_373;
assign v_3685 = v_3682 & v_372 & ~v_373 & v_375;
assign v_3686 = v_3682 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_3688 = v_3682 & v_3687;
assign v_3689 = v_7448 & v_7449;
assign v_3691 = v_3690 & v_384 & v_385;
assign v_3692 = v_3690 & v_384 & ~v_385;
assign v_3694 = v_3693 & v_1113;
assign v_3696 = v_7450 & v_7451;
assign v_3697 = v_3695 & v_391 & v_392;
assign v_3698 = v_3695 & v_391 & ~v_392 & v_394;
assign v_3699 = v_3695 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_3700 = v_3695 & v_1120;
assign v_3702 = v_7452 & v_7453;
assign v_3704 = v_3703 & v_1125;
assign v_3706 = v_3705 & v_410 & v_411;
assign v_3707 = v_3705 & v_410 & ~v_411 & v_413;
assign v_3708 = v_3705 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_3709 = v_3705 & v_421 & v_422;
assign v_3710 = v_3705 & v_424 & v_425;
assign v_3711 = v_3705 & v_424 & ~v_425 & v_427;
assign v_3712 = v_3705 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_3713 = v_3705 & v_1135;
assign v_3715 = v_3714 & v_1138;
assign v_3717 = v_3716 & v_421 & ~v_422 & v_434 & v_435;
assign v_3718 = v_3716 & v_437 & v_438;
assign v_3719 = v_3716 & v_437 & ~v_438 & v_440;
assign v_3720 = v_3716 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_3722 = v_3716 & v_3721;
assign v_3723 = v_7454 & v_7455;
assign v_3725 = v_3724 & v_449 & v_450;
assign v_3726 = v_3724 & v_449 & ~v_450;
assign v_3728 = v_3727 & v_1152;
assign v_3730 = v_7456 & v_7457;
assign v_3731 = v_3729 & v_456 & v_457;
assign v_3732 = v_3729 & v_456 & ~v_457 & v_459;
assign v_3733 = v_3729 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_3734 = v_3729 & v_1159;
assign v_3736 = v_7458 & v_7459;
assign v_3738 = v_3737 & v_1164;
assign v_3740 = v_3739 & v_491;
assign v_3742 = v_3741 & v_531 & v_532;
assign v_3743 = v_3741 & v_531 & ~v_532;
assign v_3745 = v_3744 & v_546 & v_547;
assign v_3746 = v_3744 & v_554;
assign v_3748 = v_3747 & v_558 & v_559;
assign v_3749 = v_3747 & v_558 & ~v_559 & v_561;
assign v_3750 = v_3747 & v_1196;
assign v_3753 = v_3751 & v_3752;
assign v_3754 = v_3751 & v_1201;
assign v_3756 = v_3755 & v_588 & ~v_589 & ~v_591;
assign v_3757 = v_3755 & v_593 & ~v_594;
assign v_3758 = v_3755 & v_593 & v_594;
assign v_3759 = v_3755 & v_583;
assign v_3761 = v_3760 & v_604 & v_605;
assign v_3762 = v_3760 & v_612;
assign v_3764 = v_3763 & v_616 & v_617;
assign v_3765 = v_3763 & v_616 & ~v_617 & v_619;
assign v_3766 = v_3763 & v_1214;
assign v_3769 = v_3767 & v_3768;
assign v_3770 = v_3767 & v_1219;
assign v_3772 = v_2 & v_3771;
assign v_3773 = v_641 & v_3755;
assign v_3774 = v_643 & v_3744;
assign v_3775 = v_645 & v_3744;
assign v_3776 = v_647 & v_3744;
assign v_3777 = v_649 & v_3744;
assign v_3778 = ~v_649 & v_3739;
assign v_3780 = ~v_647 & v_3779;
assign v_3782 = ~v_645 & v_3781;
assign v_3784 = ~v_643 & v_3783;
assign v_3786 = ~v_641 & v_3785;
assign v_3788 = ~v_2 & v_3787;
assign v_3790 = v_3789 & ~v_669;
assign v_3791 = v_7460 & v_7461;
assign v_3792 = v_3789 & v_669 & v_670 & v_672 & v_674;
assign v_3793 = v_7462 & v_7463;
assign v_3795 = v_3794 & v_679 & ~v_680 & v_682;
assign v_3796 = v_3794 & v_689 & ~v_690 & ~v_692;
assign v_3797 = v_3794 & v_694 & ~v_695;
assign v_3798 = v_3794 & v_694 & v_695;
assign v_3799 = v_3794 & v_684;
assign v_3801 = v_3800 & v_1251;
assign v_3803 = v_3802 & v_1254;
assign v_3804 = v_3794 & v_679 & v_680;
assign v_3805 = v_3789 & v_1257;
assign v_3807 = v_3806 & ~v_705;
assign v_3808 = v_3806 & v_710 & v_711;
assign v_3809 = v_3806 & v_718;
assign v_3811 = v_3810 & v_705 & v_722 & v_723 & ~v_724;
assign v_3813 = v_3810 & v_3812;
assign v_3814 = v_3810 & v_750 & v_751;
assign v_3815 = v_3810 & v_750 & ~v_751;
assign v_3817 = v_3816 & v_763 & v_764;
assign v_3818 = v_3816 & v_763 & ~v_764;
assign v_3820 = v_3819 & v_745 & v_758 & v_771;
assign v_3821 = v_7464 & v_7465;
assign v_3822 = v_3810 & v_779 & v_780;
assign v_3823 = v_3810 & v_787;
assign v_3825 = v_3824 & v_1278;
assign v_3827 = v_3826 & v_798 & ~v_799 & v_817;
assign v_3828 = v_3826 & v_798 & ~v_799 & ~v_817;
assign v_3829 = v_3826 & ~v_800;
assign v_3830 = v_3826 & v_808 & ~v_809;
assign v_3831 = v_3826 & v_1285;
assign v_3833 = v_3832 & v_798 & v_799 & v_814 & ~v_815;
assign v_3835 = v_3834 & v_821 & ~v_822 & v_840;
assign v_3836 = v_3834 & v_821 & ~v_822 & ~v_840;
assign v_3837 = v_3834 & ~v_823;
assign v_3838 = v_3834 & v_831 & ~v_832;
assign v_3839 = v_3834 & v_1294;
assign v_3841 = v_3840 & v_821 & v_822 & v_837 & ~v_838;
assign v_3843 = v_3842 & v_844 & ~v_845 & v_863;
assign v_3844 = v_3842 & ~v_846;
assign v_3845 = v_3842 & v_854 & ~v_855;
assign v_3846 = v_3842 & v_1302;
assign v_3848 = v_3847 & v_844 & v_845 & v_860 & v_861;
assign v_3849 = v_3842 & v_844 & ~v_845 & ~v_863;
assign v_3850 = v_3847 & v_844 & v_845 & v_860 & ~v_861;
assign v_3853 = v_3851 & v_3852;
assign v_3854 = v_3851 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_3855 = v_3851 & v_867 & v_868 & v_869;
assign v_3856 = v_3851 & v_867 & ~v_868 & ~v_872;
assign v_3858 = v_3857 & v_1315;
assign v_3859 = v_3840 & v_821 & v_822 & v_837 & v_838;
assign v_3860 = v_3832 & v_798 & v_799 & v_814 & v_815;
assign v_3862 = v_3861 & v_879 & ~v_880 & v_898;
assign v_3863 = v_3861 & v_879 & ~v_880 & ~v_898;
assign v_3864 = v_3861 & ~v_881;
assign v_3865 = v_3861 & v_889 & ~v_890;
assign v_3866 = v_3861 & v_1324;
assign v_3868 = v_3867 & v_879 & v_880 & v_895 & ~v_896;
assign v_3870 = v_3869 & v_902 & ~v_903 & v_921;
assign v_3871 = v_3869 & v_902 & ~v_903 & ~v_921;
assign v_3872 = v_3869 & ~v_904;
assign v_3873 = v_3869 & v_912 & ~v_913;
assign v_3874 = v_3869 & v_1333;
assign v_3876 = v_3875 & v_902 & v_903 & v_918 & ~v_919;
assign v_3878 = v_3877 & v_925 & ~v_926 & v_944;
assign v_3879 = v_3877 & ~v_927;
assign v_3880 = v_3877 & v_935 & ~v_936;
assign v_3881 = v_3877 & v_1341;
assign v_3883 = v_3882 & v_925 & v_926 & v_941 & v_942;
assign v_3884 = v_3877 & v_925 & ~v_926 & ~v_944;
assign v_3885 = v_3882 & v_925 & v_926 & v_941 & ~v_942;
assign v_3888 = v_3886 & v_3887;
assign v_3889 = v_3886 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_3890 = v_3886 & v_948 & v_949 & v_950;
assign v_3891 = v_3886 & v_948 & ~v_949 & ~v_953;
assign v_3893 = v_3892 & v_1354;
assign v_3894 = v_3875 & v_902 & v_903 & v_918 & v_919;
assign v_3895 = v_3867 & v_879 & v_880 & v_895 & v_896;
assign v_3897 = v_3896 & v_960 & ~v_961 & v_979;
assign v_3898 = v_3896 & v_960 & ~v_961 & ~v_979;
assign v_3899 = v_3896 & ~v_962;
assign v_3900 = v_3896 & v_970 & ~v_971;
assign v_3901 = v_3896 & v_1363;
assign v_3903 = v_3902 & v_960 & v_961 & v_976 & ~v_977;
assign v_3905 = v_3904 & v_983 & ~v_984 & v_1002;
assign v_3906 = v_3904 & v_983 & ~v_984 & ~v_1002;
assign v_3907 = v_3904 & ~v_985;
assign v_3908 = v_3904 & v_993 & ~v_994;
assign v_3909 = v_3904 & v_1372;
assign v_3911 = v_3910 & v_983 & v_984 & v_999 & ~v_1000;
assign v_3913 = v_3912 & v_1006 & ~v_1007 & v_1025;
assign v_3914 = v_3912 & ~v_1008;
assign v_3915 = v_3912 & v_1016 & ~v_1017;
assign v_3916 = v_3912 & v_1380;
assign v_3918 = v_3917 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_3919 = v_3912 & v_1006 & ~v_1007 & ~v_1025;
assign v_3920 = v_3917 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_3923 = v_3921 & v_3922;
assign v_3924 = v_3921 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_3925 = v_3921 & v_1029 & v_1030 & v_1031;
assign v_3926 = v_3921 & v_1029 & ~v_1030 & ~v_1034;
assign v_3928 = v_3927 & v_1393;
assign v_3929 = v_3910 & v_983 & v_984 & v_999 & v_1000;
assign v_3930 = v_3902 & v_960 & v_961 & v_976 & v_977;
assign v_3933 = v_3932 & v_227;
assign v_3934 = v_3932 & ~v_227 & v_229 & v_262 & ~v_264;
assign v_3935 = v_3932 & ~v_227 & v_229 & v_262 & v_264;
assign v_3936 = v_3932 & ~v_227 & v_229 & ~v_262;
assign v_3937 = v_3932 & v_230;
assign v_3938 = v_3932 & ~v_230;
assign v_3941 = v_3939 & v_3940;
assign v_3942 = v_3939 & v_1054;
assign v_3943 = v_7466 & v_7467;
assign v_3945 = v_3944 & ~v_227 & ~v_229 & v_260;
assign v_3947 = v_3946 & v_267 & v_268;
assign v_3948 = v_3946 & v_267 & ~v_268;
assign v_3950 = v_3949 & ~v_279;
assign v_3952 = v_3949 & v_3951;
assign v_3953 = v_3949 & v_279 & v_291 & ~v_292 & v_300;
assign v_3956 = v_3954 & v_3955;
assign v_3957 = v_3954 & v_321 & v_322;
assign v_3958 = v_3954 & v_321 & ~v_322 & v_324;
assign v_3959 = v_3954 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_3960 = v_3954 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_3962 = v_3961 & v_1077;
assign v_3964 = v_3963 & ~v_308 & v_309 & v_329;
assign v_3967 = v_3965 & v_3966;
assign v_3968 = v_3965 & v_1084;
assign v_3970 = v_3969 & v_345 & v_346;
assign v_3971 = v_3969 & v_345 & ~v_346 & v_348;
assign v_3972 = v_3969 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_3973 = v_3969 & v_356 & v_357;
assign v_3974 = v_3969 & v_359 & v_360;
assign v_3975 = v_3969 & v_359 & ~v_360 & v_362;
assign v_3976 = v_3969 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_3977 = v_3969 & v_1096;
assign v_3979 = v_3978 & v_1099;
assign v_3981 = v_3980 & v_356 & ~v_357 & v_369 & v_370;
assign v_3982 = v_3980 & v_372 & v_373;
assign v_3983 = v_3980 & v_372 & ~v_373 & v_375;
assign v_3984 = v_3980 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_3986 = v_3980 & v_3985;
assign v_3987 = v_7468 & v_7469;
assign v_3989 = v_3988 & v_384 & v_385;
assign v_3990 = v_3988 & v_384 & ~v_385;
assign v_3992 = v_3991 & v_1113;
assign v_3994 = v_7470 & v_7471;
assign v_3995 = v_3993 & v_391 & v_392;
assign v_3996 = v_3993 & v_391 & ~v_392 & v_394;
assign v_3997 = v_3993 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_3998 = v_3993 & v_1120;
assign v_4000 = v_7472 & v_7473;
assign v_4002 = v_4001 & v_1125;
assign v_4004 = v_4003 & v_410 & v_411;
assign v_4005 = v_4003 & v_410 & ~v_411 & v_413;
assign v_4006 = v_4003 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_4007 = v_4003 & v_421 & v_422;
assign v_4008 = v_4003 & v_424 & v_425;
assign v_4009 = v_4003 & v_424 & ~v_425 & v_427;
assign v_4010 = v_4003 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_4011 = v_4003 & v_1135;
assign v_4013 = v_4012 & v_1138;
assign v_4015 = v_4014 & v_421 & ~v_422 & v_434 & v_435;
assign v_4016 = v_4014 & v_437 & v_438;
assign v_4017 = v_4014 & v_437 & ~v_438 & v_440;
assign v_4018 = v_4014 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_4020 = v_4014 & v_4019;
assign v_4021 = v_7474 & v_7475;
assign v_4023 = v_4022 & v_449 & v_450;
assign v_4024 = v_4022 & v_449 & ~v_450;
assign v_4026 = v_4025 & v_1152;
assign v_4028 = v_7476 & v_7477;
assign v_4029 = v_4027 & v_456 & v_457;
assign v_4030 = v_4027 & v_456 & ~v_457 & v_459;
assign v_4031 = v_4027 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_4032 = v_4027 & v_1159;
assign v_4034 = v_7478 & v_7479;
assign v_4036 = v_4035 & v_1164;
assign v_4038 = v_4037 & v_491;
assign v_4039 = v_4037 & ~v_491 & v_493 & v_526 & ~v_528;
assign v_4040 = v_4037 & ~v_491 & v_493 & v_526 & v_528;
assign v_4041 = v_4037 & ~v_491 & v_493 & ~v_526;
assign v_4042 = v_4037 & v_494;
assign v_4043 = v_4037 & ~v_494;
assign v_4046 = v_4044 & v_4045;
assign v_4047 = v_4044 & v_1180;
assign v_4048 = v_7480 & v_7481;
assign v_4050 = v_4049 & ~v_491 & ~v_493 & v_524;
assign v_4052 = v_4051 & v_531 & v_532;
assign v_4053 = v_4051 & v_531 & ~v_532;
assign v_4055 = v_4054 & v_546 & v_547;
assign v_4056 = v_4054 & v_546 & ~v_547 & ~v_551;
assign v_4058 = v_4057 & v_546 & ~v_547 & v_551;
assign v_4060 = v_4059 & v_554;
assign v_4062 = v_4061 & v_558 & v_559;
assign v_4063 = v_4061 & v_558 & ~v_559 & v_561;
assign v_4064 = v_4061 & v_1196;
assign v_4067 = v_4065 & v_4066;
assign v_4068 = v_4065 & v_1201;
assign v_4070 = v_4069 & v_588 & ~v_589 & ~v_591;
assign v_4071 = v_4069 & v_593 & ~v_594;
assign v_4072 = v_4069 & v_593 & v_594;
assign v_4073 = v_4069 & v_583;
assign v_4075 = v_4074 & v_604 & v_605;
assign v_4076 = v_4074 & v_604 & ~v_605 & ~v_609;
assign v_4078 = v_4077 & v_604 & ~v_605 & v_609;
assign v_4080 = v_4079 & v_612;
assign v_4082 = v_4081 & v_616 & v_617;
assign v_4083 = v_4081 & v_616 & ~v_617 & v_619;
assign v_4084 = v_4081 & v_1214;
assign v_4087 = v_4085 & v_4086;
assign v_4088 = v_4085 & v_1219;
assign v_4090 = v_2 & v_4089;
assign v_4091 = v_641 & v_4069;
assign v_4092 = v_643 & v_4054;
assign v_4093 = v_645 & v_4054;
assign v_4094 = v_647 & v_4054;
assign v_4095 = v_649 & v_4054;
assign v_4096 = ~v_649 & v_4037;
assign v_4098 = ~v_647 & v_4097;
assign v_4100 = ~v_645 & v_4099;
assign v_4102 = ~v_643 & v_4101;
assign v_4104 = ~v_641 & v_4103;
assign v_4106 = ~v_2 & v_4105;
assign v_4108 = v_4107 & ~v_669;
assign v_4109 = v_7482 & v_7483;
assign v_4110 = v_4107 & v_669 & v_670 & v_672 & v_674;
assign v_4111 = v_7484 & v_7485;
assign v_4113 = v_4112 & v_679 & ~v_680 & v_682;
assign v_4114 = v_4112 & v_689 & ~v_690 & ~v_692;
assign v_4115 = v_4112 & v_694 & ~v_695;
assign v_4116 = v_4112 & v_694 & v_695;
assign v_4117 = v_4112 & v_684;
assign v_4119 = v_4118 & v_1251;
assign v_4121 = v_4120 & v_1254;
assign v_4122 = v_4112 & v_679 & v_680;
assign v_4123 = v_4107 & v_1257;
assign v_4125 = v_4124 & ~v_705;
assign v_4126 = v_4124 & v_710 & v_711;
assign v_4127 = v_4124 & v_710 & ~v_711 & ~v_715;
assign v_4129 = v_4128 & v_710 & ~v_711 & v_715;
assign v_4131 = v_4130 & v_718;
assign v_4133 = v_4132 & v_705 & v_722 & v_723 & ~v_724;
assign v_4135 = v_4132 & v_4134;
assign v_4136 = v_4132 & v_750 & v_751;
assign v_4137 = v_4132 & v_750 & ~v_751;
assign v_4139 = v_4138 & v_763 & v_764;
assign v_4140 = v_4138 & v_763 & ~v_764;
assign v_4142 = v_4141 & v_745 & v_758 & v_771;
assign v_4143 = v_7486 & v_7487;
assign v_4144 = v_4132 & v_779 & v_780;
assign v_4145 = v_4132 & v_779 & ~v_780 & ~v_784;
assign v_4147 = v_4146 & v_779 & ~v_780 & v_784;
assign v_4149 = v_4148 & v_787;
assign v_4151 = v_4150 & v_1278;
assign v_4153 = v_4152 & v_798 & ~v_799 & v_817;
assign v_4154 = v_4152 & v_798 & ~v_799 & ~v_817;
assign v_4155 = v_4152 & ~v_800;
assign v_4156 = v_4152 & v_808 & ~v_809;
assign v_4157 = v_4152 & v_1285;
assign v_4159 = v_4158 & v_798 & v_799 & v_814 & ~v_815;
assign v_4161 = v_4160 & v_821 & ~v_822 & v_840;
assign v_4162 = v_4160 & v_821 & ~v_822 & ~v_840;
assign v_4163 = v_4160 & ~v_823;
assign v_4164 = v_4160 & v_831 & ~v_832;
assign v_4165 = v_4160 & v_1294;
assign v_4167 = v_4166 & v_821 & v_822 & v_837 & ~v_838;
assign v_4169 = v_4168 & v_844 & ~v_845 & v_863;
assign v_4170 = v_4168 & ~v_846;
assign v_4171 = v_4168 & v_854 & ~v_855;
assign v_4172 = v_4168 & v_1302;
assign v_4174 = v_4173 & v_844 & v_845 & v_860 & v_861;
assign v_4175 = v_4168 & v_844 & ~v_845 & ~v_863;
assign v_4176 = v_4173 & v_844 & v_845 & v_860 & ~v_861;
assign v_4179 = v_4177 & v_4178;
assign v_4180 = v_4177 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_4181 = v_4177 & v_867 & v_868 & v_869;
assign v_4182 = v_4177 & v_867 & ~v_868 & ~v_872;
assign v_4184 = v_4183 & v_1315;
assign v_4185 = v_4166 & v_821 & v_822 & v_837 & v_838;
assign v_4186 = v_4158 & v_798 & v_799 & v_814 & v_815;
assign v_4188 = v_4187 & v_879 & ~v_880 & v_898;
assign v_4189 = v_4187 & v_879 & ~v_880 & ~v_898;
assign v_4190 = v_4187 & ~v_881;
assign v_4191 = v_4187 & v_889 & ~v_890;
assign v_4192 = v_4187 & v_1324;
assign v_4194 = v_4193 & v_879 & v_880 & v_895 & ~v_896;
assign v_4196 = v_4195 & v_902 & ~v_903 & v_921;
assign v_4197 = v_4195 & v_902 & ~v_903 & ~v_921;
assign v_4198 = v_4195 & ~v_904;
assign v_4199 = v_4195 & v_912 & ~v_913;
assign v_4200 = v_4195 & v_1333;
assign v_4202 = v_4201 & v_902 & v_903 & v_918 & ~v_919;
assign v_4204 = v_4203 & v_925 & ~v_926 & v_944;
assign v_4205 = v_4203 & ~v_927;
assign v_4206 = v_4203 & v_935 & ~v_936;
assign v_4207 = v_4203 & v_1341;
assign v_4209 = v_4208 & v_925 & v_926 & v_941 & v_942;
assign v_4210 = v_4203 & v_925 & ~v_926 & ~v_944;
assign v_4211 = v_4208 & v_925 & v_926 & v_941 & ~v_942;
assign v_4214 = v_4212 & v_4213;
assign v_4215 = v_4212 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_4216 = v_4212 & v_948 & v_949 & v_950;
assign v_4217 = v_4212 & v_948 & ~v_949 & ~v_953;
assign v_4219 = v_4218 & v_1354;
assign v_4220 = v_4201 & v_902 & v_903 & v_918 & v_919;
assign v_4221 = v_4193 & v_879 & v_880 & v_895 & v_896;
assign v_4223 = v_4222 & v_960 & ~v_961 & v_979;
assign v_4224 = v_4222 & v_960 & ~v_961 & ~v_979;
assign v_4225 = v_4222 & ~v_962;
assign v_4226 = v_4222 & v_970 & ~v_971;
assign v_4227 = v_4222 & v_1363;
assign v_4229 = v_4228 & v_960 & v_961 & v_976 & ~v_977;
assign v_4231 = v_4230 & v_983 & ~v_984 & v_1002;
assign v_4232 = v_4230 & v_983 & ~v_984 & ~v_1002;
assign v_4233 = v_4230 & ~v_985;
assign v_4234 = v_4230 & v_993 & ~v_994;
assign v_4235 = v_4230 & v_1372;
assign v_4237 = v_4236 & v_983 & v_984 & v_999 & ~v_1000;
assign v_4239 = v_4238 & v_1006 & ~v_1007 & v_1025;
assign v_4240 = v_4238 & ~v_1008;
assign v_4241 = v_4238 & v_1016 & ~v_1017;
assign v_4242 = v_4238 & v_1380;
assign v_4244 = v_4243 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_4245 = v_4238 & v_1006 & ~v_1007 & ~v_1025;
assign v_4246 = v_4243 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_4249 = v_4247 & v_4248;
assign v_4250 = v_4247 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_4251 = v_4247 & v_1029 & v_1030 & v_1031;
assign v_4252 = v_4247 & v_1029 & ~v_1030 & ~v_1034;
assign v_4254 = v_4253 & v_1393;
assign v_4255 = v_4236 & v_983 & v_984 & v_999 & v_1000;
assign v_4256 = v_4228 & v_960 & v_961 & v_976 & v_977;
assign v_4262 = ~v_4260 & ~v_4261;
assign v_4265 = ~v_4263 & v_4264;
assign v_4266 = ~v_4262 & ~v_4265;
assign v_4267 = ~v_4260 & ~v_4261;
assign v_4268 = ~v_4263 & v_4264;
assign v_4269 = ~v_4267 & ~v_4268;
assign v_4270 = v_4266 & v_4269;
assign v_4271 = ~v_4260 & ~v_4261;
assign v_4272 = ~v_4263 & v_4264;
assign v_4273 = ~v_4271 & ~v_4272;
assign v_4274 = v_4270 & v_4273;
assign v_4275 = ~v_4260 & ~v_4261;
assign v_4276 = ~v_4263 & v_4264;
assign v_4277 = ~v_4275 & ~v_4276;
assign v_4278 = v_4274 & v_4277;
assign v_4279 = ~v_4260 & ~v_4261;
assign v_4280 = ~v_4263 & v_4264;
assign v_4281 = ~v_4279 & ~v_4280;
assign v_4282 = v_4278 & v_4281;
assign v_4283 = ~v_4260 & ~v_4261;
assign v_4284 = ~v_4263 & v_4264;
assign v_4285 = ~v_4283 & ~v_4284;
assign v_4286 = v_4282 & v_4285;
assign v_4287 = ~v_4260 & ~v_4261;
assign v_4288 = ~v_4263 & v_4264;
assign v_4289 = ~v_4287 & ~v_4288;
assign v_4290 = v_4286 & v_4289;
assign v_4291 = ~v_4260 & ~v_4261;
assign v_4292 = ~v_4263 & v_4264;
assign v_4293 = ~v_4291 & ~v_4292;
assign v_4294 = v_4290 & v_4293;
assign v_4295 = ~v_4260 & ~v_4261;
assign v_4296 = ~v_4263 & v_4264;
assign v_4297 = ~v_4295 & ~v_4296;
assign v_4298 = v_4294 & v_4297;
assign v_4299 = ~v_4260 & ~v_4261;
assign v_4300 = ~v_4263 & v_4264;
assign v_4301 = ~v_4299 & ~v_4300;
assign v_4302 = v_4298 & v_4301;
assign v_4303 = ~v_4260 & ~v_4261;
assign v_4304 = ~v_4263 & v_4264;
assign v_4305 = ~v_4303 & ~v_4304;
assign v_4306 = v_4302 & v_4305;
assign v_4307 = ~v_4260 & ~v_4261;
assign v_4308 = ~v_4263 & v_4264;
assign v_4309 = ~v_4307 & ~v_4308;
assign v_4310 = v_4306 & v_4309;
assign v_4311 = ~v_4260 & ~v_4261;
assign v_4312 = ~v_4263 & v_4264;
assign v_4313 = ~v_4311 & ~v_4312;
assign v_4314 = v_4310 & v_4313;
assign v_4315 = ~v_4260 & ~v_4261;
assign v_4316 = ~v_4263 & v_4264;
assign v_4317 = ~v_4315 & ~v_4316;
assign v_4318 = v_4314 & v_4317;
assign v_4319 = ~v_4260 & ~v_4261;
assign v_4320 = ~v_4263 & v_4264;
assign v_4321 = ~v_4319 & ~v_4320;
assign v_4322 = v_4318 & v_4321;
assign v_4323 = ~v_4260 & ~v_4261;
assign v_4324 = ~v_4263 & v_4264;
assign v_4325 = ~v_4323 & ~v_4324;
assign v_4326 = v_4322 & v_4325;
assign v_4327 = ~v_4260 & ~v_4261;
assign v_4328 = ~v_4263 & v_4264;
assign v_4329 = ~v_4327 & ~v_4328;
assign v_4330 = v_4326 & v_4329;
assign v_4331 = ~v_4260 & ~v_4261;
assign v_4332 = ~v_4263 & v_4264;
assign v_4333 = ~v_4331 & ~v_4332;
assign v_4334 = v_4330 & v_4333;
assign v_4335 = ~v_4260 & ~v_4261;
assign v_4336 = ~v_4263 & v_4264;
assign v_4337 = ~v_4335 & ~v_4336;
assign v_4338 = v_4334 & v_4337;
assign v_4339 = ~v_4260 & ~v_4261;
assign v_4340 = ~v_4263 & v_4264;
assign v_4341 = ~v_4339 & ~v_4340;
assign v_4342 = v_4338 & v_4341;
assign v_4343 = ~v_4260 & ~v_4261;
assign v_4344 = ~v_4263 & v_4264;
assign v_4345 = ~v_4343 & ~v_4344;
assign v_4346 = v_4342 & v_4345;
assign v_4347 = ~v_4260 & ~v_4261;
assign v_4348 = ~v_4263 & v_4264;
assign v_4349 = ~v_4347 & ~v_4348;
assign v_4350 = v_4346 & v_4349;
assign v_4351 = ~v_4260 & ~v_4261;
assign v_4352 = ~v_4263 & v_4264;
assign v_4353 = ~v_4351 & ~v_4352;
assign v_4354 = v_4350 & v_4353;
assign v_4355 = ~v_4260 & ~v_4261;
assign v_4356 = ~v_4263 & v_4264;
assign v_4357 = ~v_4355 & ~v_4356;
assign v_4358 = v_4354 & v_4357;
assign v_4359 = ~v_4260 & ~v_4261;
assign v_4360 = ~v_4263 & v_4264;
assign v_4361 = ~v_4359 & ~v_4360;
assign v_4362 = v_4358 & v_4361;
assign v_4363 = ~v_4260 & ~v_4261;
assign v_4364 = ~v_4263 & v_4264;
assign v_4365 = ~v_4363 & ~v_4364;
assign v_4366 = v_4362 & v_4365;
assign v_4367 = ~v_4260 & ~v_4261;
assign v_4368 = ~v_4263 & v_4264;
assign v_4369 = ~v_4367 & ~v_4368;
assign v_4370 = v_4366 & v_4369;
assign v_4371 = ~v_4260 & ~v_4261;
assign v_4372 = ~v_4263 & v_4264;
assign v_4373 = ~v_4371 & ~v_4372;
assign v_4374 = v_4370 & v_4373;
assign v_4375 = ~v_4260 & ~v_4261;
assign v_4376 = ~v_4263 & v_4264;
assign v_4377 = ~v_4375 & ~v_4376;
assign v_4378 = v_4374 & v_4377;
assign v_4379 = ~v_4260 & ~v_4261;
assign v_4380 = ~v_4263 & v_4264;
assign v_4381 = ~v_4379 & ~v_4380;
assign v_4382 = v_4378 & v_4381;
assign v_4383 = ~v_4260 & ~v_4261;
assign v_4384 = ~v_4263 & v_4264;
assign v_4385 = ~v_4383 & ~v_4384;
assign v_4386 = v_4382 & v_4385;
assign v_4387 = ~v_4260 & ~v_4261;
assign v_4388 = ~v_4263 & v_4264;
assign v_4389 = ~v_4387 & ~v_4388;
assign v_4390 = v_4386 & v_4389;
assign v_4391 = ~v_4260 & ~v_4261;
assign v_4392 = ~v_4263 & v_4264;
assign v_4393 = ~v_4391 & ~v_4392;
assign v_4394 = v_4390 & v_4393;
assign v_4395 = ~v_4260 & ~v_4261;
assign v_4396 = ~v_4263 & v_4264;
assign v_4397 = ~v_4395 & ~v_4396;
assign v_4398 = v_4394 & v_4397;
assign v_4399 = ~v_4260 & ~v_4261;
assign v_4400 = ~v_4263 & v_4264;
assign v_4401 = ~v_4399 & ~v_4400;
assign v_4402 = v_4398 & v_4401;
assign v_4403 = ~v_4260 & ~v_4261;
assign v_4404 = ~v_4263 & v_4264;
assign v_4405 = ~v_4403 & ~v_4404;
assign v_4406 = v_4402 & v_4405;
assign v_4407 = ~v_4260 & ~v_4261;
assign v_4408 = ~v_4263 & v_4264;
assign v_4409 = ~v_4407 & ~v_4408;
assign v_4410 = v_4406 & v_4409;
assign v_4411 = ~v_4260 & ~v_4261;
assign v_4412 = ~v_4263 & v_4264;
assign v_4413 = ~v_4411 & ~v_4412;
assign v_4414 = v_4410 & v_4413;
assign v_4415 = ~v_4260 & ~v_4261;
assign v_4416 = ~v_4263 & v_4264;
assign v_4417 = ~v_4415 & ~v_4416;
assign v_4418 = v_4414 & v_4417;
assign v_4419 = ~v_4260 & ~v_4261;
assign v_4420 = ~v_4263 & v_4264;
assign v_4421 = ~v_4419 & ~v_4420;
assign v_4422 = v_4418 & v_4421;
assign v_4423 = ~v_4260 & ~v_4261;
assign v_4424 = ~v_4263 & v_4264;
assign v_4425 = ~v_4423 & ~v_4424;
assign v_4426 = v_4422 & v_4425;
assign v_4427 = ~v_4260 & ~v_4261;
assign v_4428 = ~v_4263 & v_4264;
assign v_4429 = ~v_4427 & ~v_4428;
assign v_4430 = v_4426 & v_4429;
assign v_4431 = ~v_4260 & ~v_4261;
assign v_4432 = ~v_4263 & v_4264;
assign v_4433 = ~v_4431 & ~v_4432;
assign v_4434 = v_4430 & v_4433;
assign v_4435 = ~v_4260 & ~v_4261;
assign v_4436 = ~v_4263 & v_4264;
assign v_4437 = ~v_4435 & ~v_4436;
assign v_4438 = v_4434 & v_4437;
assign v_4439 = ~v_4260 & ~v_4261;
assign v_4440 = ~v_4263 & v_4264;
assign v_4441 = ~v_4439 & ~v_4440;
assign v_4442 = v_4438 & v_4441;
assign v_4443 = ~v_4260 & ~v_4261;
assign v_4444 = ~v_4263 & v_4264;
assign v_4445 = ~v_4443 & ~v_4444;
assign v_4446 = v_4442 & v_4445;
assign v_4447 = ~v_4260 & ~v_4261;
assign v_4448 = ~v_4263 & v_4264;
assign v_4449 = ~v_4447 & ~v_4448;
assign v_4450 = v_4446 & v_4449;
assign v_4451 = ~v_4260 & ~v_4261;
assign v_4452 = ~v_4263 & v_4264;
assign v_4453 = ~v_4451 & ~v_4452;
assign v_4454 = v_4450 & v_4453;
assign v_4455 = ~v_4260 & ~v_4261;
assign v_4456 = ~v_4263 & v_4264;
assign v_4457 = ~v_4455 & ~v_4456;
assign v_4458 = v_4454 & v_4457;
assign v_4459 = ~v_4263 & v_4264;
assign v_4460 = v_4458 & ~v_4459;
assign v_4461 = ~v_4263 & v_4264;
assign v_4462 = v_4460 & ~v_4461;
assign v_4463 = ~v_4263 & v_4264;
assign v_4464 = v_4462 & ~v_4463;
assign v_4465 = ~v_4263 & v_4264;
assign v_4466 = v_4464 & ~v_4465;
assign v_4467 = ~v_4263 & v_4264;
assign v_4468 = v_4466 & ~v_4467;
assign v_4471 = v_4469 & v_4470;
assign v_4472 = v_4469 & ~v_4470;
assign v_4474 = v_4468 & v_4473;
assign v_4478 = v_4477;
assign v_4479 = ~v_4477;
assign v_4484 = v_4483;
assign v_4489 = ~v_4488;
assign v_4491 = v_4488 & v_4490;
assign v_4494 = v_4488 & ~v_4490 & v_4492 & v_4493;
assign v_4496 = v_4488 & ~v_4490 & v_4492 & ~v_4493 & ~v_4495;
assign v_4498 = v_4488 & ~v_4490 & ~v_4492 & ~v_4497;
assign v_4500 = v_4488 & ~v_4490 & ~v_4492 & v_4497 & v_4499;
assign v_4502 = v_7488 & v_7489;
assign v_4504 = v_7490 & v_7491;
assign v_4508 = v_7492 & v_7493;
assign v_4509 = v_7494 & v_7495;
assign v_4512 = v_4510 & v_4511;
assign v_4513 = v_4510 & ~v_4511;
assign v_4515 = v_7496 & v_7497;
assign v_4517 = ~v_4483 & ~v_4485 & v_4516;
assign v_4519 = ~v_4483 & v_4485 & ~v_4518;
assign v_4521 = ~v_4483 & v_4485 & v_4518 & ~v_4520;
assign v_4522 = ~v_4483 & v_4485 & v_4518 & v_4520;
assign v_4525 = v_4523 & v_4524;
assign v_4526 = v_4523 & ~v_4524;
assign v_4531 = v_4480 & v_4527 & v_4530;
assign v_4532 = v_4480 & v_4527 & ~v_4530;
assign v_4534 = v_4474 & v_4533;
assign v_4538 = v_4536 & v_4537;
assign v_4540 = v_4536 & ~v_4537 & v_4539;
assign v_4543 = v_4541 & ~v_4542;
assign v_4545 = v_4541 & v_4542 & v_4544;
assign v_4546 = v_4541 & v_4542 & ~v_4544;
assign v_4550 = v_4535 & v_4547 & v_4548 & v_4549;
assign v_4552 = v_4535 & v_4547 & v_4548 & ~v_4549 & v_4551;
assign v_4555 = ~v_4553 & v_4554;
assign v_4557 = v_4535 & v_4547 & ~v_4548 & v_4556;
assign v_4560 = v_4558 & v_4559;
assign v_4561 = v_4558 & ~v_4559;
assign v_4563 = v_4534 & v_4562;
assign v_4566 = ~v_4564 & ~v_4565;
assign v_4569 = v_4567 & v_4568;
assign v_4570 = v_4567 & ~v_4568;
assign v_4573 = v_4571 & ~v_4572;
assign v_4575 = v_4571 & v_4572 & v_4574;
assign v_4576 = v_4571 & v_4572 & ~v_4574;
assign v_4579 = v_4577 & v_4578;
assign v_4581 = v_4577 & ~v_4578 & v_4580;
assign v_4583 = v_4577 & ~v_4578 & ~v_4580 & v_4582;
assign v_4584 = v_4577 & ~v_4578 & ~v_4580 & ~v_4582;
assign v_4586 = ~v_4564 & v_4565 & v_4585;
assign v_4588 = v_4563 & v_4587;
assign v_4591 = v_4589 & ~v_4590;
assign v_4593 = v_4589 & v_4590 & ~v_4592;
assign v_4597 = v_4589 & v_4590 & v_4592 & v_4596;
assign v_4598 = v_4589 & v_4590 & v_4592 & ~v_4596;
assign v_4600 = v_4588 & v_4599;
assign v_4603 = v_4601 & v_4602;
assign v_4605 = v_4601 & ~v_4602 & v_4604;
assign v_4607 = v_4601 & ~v_4602 & ~v_4604 & v_4606;
assign v_4609 = v_4601 & ~v_4602 & ~v_4604 & ~v_4606 & v_4608;
assign v_4611 = v_7498 & v_7499;
assign v_4614 = v_4612 & v_4613;
assign v_4617 = v_4615 & v_4616;
assign v_4619 = v_4615 & ~v_4616 & v_4618;
assign v_4621 = v_4615 & ~v_4616 & ~v_4618 & v_4620;
assign v_4623 = v_4615 & ~v_4616 & ~v_4618 & ~v_4620 & v_4622;
assign v_4624 = v_4615 & ~v_4616 & ~v_4618 & ~v_4620 & ~v_4622;
assign v_4627 = v_4612 & ~v_4613 & v_4625 & v_4626;
assign v_4630 = v_4628 & v_4629;
assign v_4632 = v_4628 & ~v_4629 & v_4631;
assign v_4634 = v_4628 & ~v_4629 & ~v_4631 & v_4633;
assign v_4636 = v_4628 & ~v_4629 & ~v_4631 & ~v_4633 & v_4635;
assign v_4638 = v_7500 & v_7501;
assign v_4639 = v_7502 & v_7503;
assign v_4642 = v_4640 & v_4641;
assign v_4643 = v_4640 & ~v_4641;
assign v_4646 = v_7504 & v_7505;
assign v_4649 = v_4647 & v_4648;
assign v_4651 = v_4647 & ~v_4648 & v_4650;
assign v_4653 = v_4647 & ~v_4648 & ~v_4650 & v_4652;
assign v_4655 = v_4647 & ~v_4648 & ~v_4650 & ~v_4652 & ~v_4654;
assign v_4657 = v_7506 & v_7507;
assign v_4658 = v_7508 & v_7509;
assign v_4660 = v_7510 & v_7511;
assign v_4663 = v_4661 & v_4662;
assign v_4664 = v_4661 & ~v_4662;
assign v_4668 = v_4666 & v_4667;
assign v_4670 = v_4666 & ~v_4667 & v_4669;
assign v_4672 = v_4666 & ~v_4667 & ~v_4669 & v_4671;
assign v_4674 = v_4666 & ~v_4667 & ~v_4669 & ~v_4671 & v_4673;
assign v_4676 = v_7512 & v_7513;
assign v_4679 = v_4677 & v_4678;
assign v_4682 = v_4680 & v_4681;
assign v_4684 = v_4680 & ~v_4681 & v_4683;
assign v_4686 = v_4680 & ~v_4681 & ~v_4683 & v_4685;
assign v_4688 = v_4680 & ~v_4681 & ~v_4683 & ~v_4685 & v_4687;
assign v_4689 = v_4680 & ~v_4681 & ~v_4683 & ~v_4685 & ~v_4687;
assign v_4692 = v_4677 & ~v_4678 & v_4690 & v_4691;
assign v_4695 = v_4693 & v_4694;
assign v_4697 = v_4693 & ~v_4694 & v_4696;
assign v_4699 = v_4693 & ~v_4694 & ~v_4696 & v_4698;
assign v_4701 = v_4693 & ~v_4694 & ~v_4696 & ~v_4698 & v_4700;
assign v_4703 = v_7514 & v_7515;
assign v_4704 = v_7516 & v_7517;
assign v_4707 = v_4705 & v_4706;
assign v_4708 = v_4705 & ~v_4706;
assign v_4711 = v_7518 & v_7519;
assign v_4714 = v_4712 & v_4713;
assign v_4716 = v_4712 & ~v_4713 & v_4715;
assign v_4718 = v_4712 & ~v_4713 & ~v_4715 & v_4717;
assign v_4720 = v_4712 & ~v_4713 & ~v_4715 & ~v_4717 & ~v_4719;
assign v_4722 = v_7520 & v_7521;
assign v_4723 = v_7522 & v_7523;
assign v_4725 = v_7524 & v_7525;
assign v_4728 = v_4726 & v_4727;
assign v_4729 = v_4726 & ~v_4727;
assign v_4732 = v_4665 & v_4730 & v_4731;
assign v_4734 = v_4665 & v_4730 & ~v_4731 & v_4733;
assign v_4735 = v_4665 & v_4730 & ~v_4731 & ~v_4733;
assign v_4738 = v_4736 & v_4737;
assign v_4739 = v_4736 & ~v_4737;
assign v_4741 = v_4600 & v_4740;
assign v_4744 = v_4741;
assign v_4748 = v_4747;
assign v_4753 = ~v_4752;
assign v_4755 = v_4752 & v_4754;
assign v_4758 = v_4752 & ~v_4754 & v_4756 & v_4757;
assign v_4760 = v_4752 & ~v_4754 & v_4756 & ~v_4757 & ~v_4759;
assign v_4762 = v_4752 & ~v_4754 & ~v_4756 & ~v_4761;
assign v_4764 = v_4752 & ~v_4754 & ~v_4756 & v_4761 & v_4763;
assign v_4766 = v_7526 & v_7527;
assign v_4768 = v_7528 & v_7529;
assign v_4772 = v_7530 & v_7531;
assign v_4773 = v_7532 & v_7533;
assign v_4776 = v_4774 & v_4775;
assign v_4777 = v_4774 & ~v_4775;
assign v_4779 = v_7534 & v_7535;
assign v_4781 = ~v_4747 & ~v_4749 & v_4780;
assign v_4783 = ~v_4747 & v_4749 & ~v_4782;
assign v_4785 = ~v_4747 & v_4749 & v_4782 & ~v_4784;
assign v_4786 = ~v_4747 & v_4749 & v_4782 & v_4784;
assign v_4789 = v_4787 & v_4788;
assign v_4790 = v_4787 & ~v_4788;
assign v_4792 = v_4744 & v_4791;
assign v_4795 = v_4259 & v_4792;
assign v_4796 = ~v_4259 & v_4744 & v_4791;
assign v_4800 = v_4798 & v_4799;
assign v_4801 = v_4798 & ~v_4799;
assign v_4804 = v_4802 & v_4803;
assign v_4808 = v_4802 & ~v_4803 & ~v_4807;
assign v_4809 = v_4802 & ~v_4803 & v_4807;
assign v_4813 = v_4810;
assign v_4816 = v_4814 & v_4815;
assign v_4818 = v_4814 & ~v_4815 & v_4817;
assign v_4822 = v_4814 & ~v_4815 & ~v_4817 & v_4821;
assign v_4823 = v_4814 & ~v_4815 & ~v_4817 & ~v_4821;
assign v_4826 = v_4824 & v_4825;
assign v_4828 = v_4824 & ~v_4825 & v_4827;
assign v_4831 = v_4829 & v_4830;
assign v_4832 = v_4829 & ~v_4830;
assign v_4835 = v_4824 & ~v_4825 & ~v_4827 & v_4833 & v_4834;
assign v_4836 = v_4824 & ~v_4825 & ~v_4827 & v_4833 & ~v_4834;
assign v_4838 = v_4797 & v_4837;
assign v_4841 = ~v_4839 & v_4840;
assign v_4843 = ~v_4839 & ~v_4840 & v_4842;
assign v_4846 = v_4844 & v_4845;
assign v_4848 = v_4844 & ~v_4845 & v_4847;
assign v_4851 = v_4849 & ~v_4850;
assign v_4852 = v_4844 & ~v_4845 & ~v_4847;
assign v_4853 = v_4849 & v_4850;
assign v_4855 = v_4838 & v_4854;
assign v_4858 = v_4856 & v_4857;
assign v_4859 = v_4856 & ~v_4857;
assign v_4862 = v_4860 & v_4861;
assign v_4866 = v_4860 & ~v_4861 & ~v_4865;
assign v_4867 = v_4860 & ~v_4861 & v_4865;
assign v_4871 = v_4868;
assign v_4874 = v_4872 & v_4873;
assign v_4876 = v_4872 & ~v_4873 & v_4875;
assign v_4880 = v_4872 & ~v_4873 & ~v_4875 & v_4879;
assign v_4881 = v_4872 & ~v_4873 & ~v_4875 & ~v_4879;
assign v_4884 = v_4882 & v_4883;
assign v_4886 = v_4882 & ~v_4883 & v_4885;
assign v_4889 = v_4887 & v_4888;
assign v_4890 = v_4887 & ~v_4888;
assign v_4893 = v_4882 & ~v_4883 & ~v_4885 & v_4891 & v_4892;
assign v_4894 = v_4882 & ~v_4883 & ~v_4885 & v_4891 & ~v_4892;
assign v_4896 = v_4258 & v_4855 & v_4895;
assign v_4898 = v_4897 & v_4797 & v_4837;
assign v_4900 = v_4899 & v_4792;
assign v_4902 = v_4901 & v_4792;
assign v_4904 = v_4903 & v_4744 & v_4791;
assign v_4906 = v_4905 & v_4744 & v_4791;
assign v_4907 = ~v_4905 & v_4741;
assign v_4909 = ~v_4903 & v_4908;
assign v_4911 = ~v_4901 & v_4910;
assign v_4913 = ~v_4899 & v_4912;
assign v_4915 = ~v_4897 & v_4914;
assign v_4917 = ~v_4258 & v_4916;
assign v_4921 = v_4918;
assign v_4924 = v_4921;
assign v_4927 = v_4925 & ~v_4926;
assign v_4929 = v_4925 & v_4926 & ~v_4928;
assign v_4932 = v_4925 & v_4926 & v_4928 & ~v_4930 & ~v_4931;
assign v_4933 = v_4925 & v_4926 & v_4928 & v_4930;
assign v_4934 = v_4925 & v_4926 & v_4928 & ~v_4930 & v_4931;
assign v_4937 = v_4935 & v_4936;
assign v_4939 = v_4935 & ~v_4936 & v_4938;
assign v_4942 = ~v_4940 & v_4941;
assign v_4944 = ~v_4940 & ~v_4941 & v_4943;
assign v_4947 = v_4945 & v_4946;
assign v_4949 = v_4945 & ~v_4946 & v_4948;
assign v_4952 = v_4950 & ~v_4951;
assign v_4953 = v_4945 & ~v_4946 & ~v_4948;
assign v_4954 = v_4950 & v_4951;
assign v_4957 = v_4935 & ~v_4936 & ~v_4938 & v_4955 & v_4956;
assign v_4958 = v_4935 & ~v_4936 & ~v_4938 & v_4955 & ~v_4956;
assign v_4960 = v_4924 & v_4959;
assign v_4964 = v_4962 & v_4963;
assign v_4965 = v_4962 & ~v_4963;
assign v_4968 = v_4966 & v_4967;
assign v_4972 = v_4966 & ~v_4967 & ~v_4971;
assign v_4973 = v_4966 & ~v_4967 & v_4971;
assign v_4977 = v_4974;
assign v_4981 = v_4961 & v_4978 & v_4979 & ~v_4980;
assign v_4986 = v_7536 & v_7537;
assign v_4988 = v_7538 & v_7539;
assign v_4990 = v_7540 & v_7541;
assign v_4992 = v_7542 & v_7543;
assign v_4996 = v_4993 & ~v_4994 & v_4995;
assign v_4997 = v_4993 & ~v_4994 & ~v_4995;
assign v_4999 = v_4993 & v_4994 & v_4998;
assign v_5000 = v_4993 & v_4994 & ~v_4998;
assign v_5004 = v_5002 & v_5003;
assign v_5005 = v_5002 & ~v_5003;
assign v_5008 = v_5006 & v_5007;
assign v_5013 = v_5006 & ~v_5007;
assign v_5017 = v_5015 & v_5016;
assign v_5018 = v_5015 & ~v_5016;
assign v_5021 = v_5019 & v_5020;
assign v_5026 = v_5019 & ~v_5020;
assign v_5030 = v_5001 & v_5014 & v_5027;
assign v_5033 = v_5031 & v_5032;
assign v_5034 = v_5031 & ~v_5032;
assign v_5037 = v_5035 & v_5036;
assign v_5041 = v_5035 & ~v_5036 & ~v_5040;
assign v_5042 = v_5035 & ~v_5036 & v_5040;
assign v_5046 = v_5043;
assign v_5049 = v_4961 & v_4978 & ~v_4979 & v_5047 & v_5048;
assign v_5050 = v_4961 & v_4978 & ~v_4979 & v_5047 & ~v_5048;
assign v_5051 = v_4961 & v_4978 & v_4979 & v_4980 & v_4982;
assign v_5053 = v_4960 & v_5052;
assign v_5057 = v_5055 & ~v_5056;
assign v_5059 = v_5054 & v_5058;
assign v_5061 = ~v_4483 & v_4485 & v_4518 & ~v_4520;
assign v_5062 = ~v_4483 & v_4485 & v_4518 & v_4520;
assign v_5063 = ~v_4483 & v_4485 & ~v_4518;
assign v_5066 = v_5065;
assign v_5068 = v_5067;
assign v_5069 = v_7544 & v_7545;
assign v_5071 = v_5070 & ~v_4483 & ~v_4485 & v_4516;
assign v_5073 = v_5060 & ~v_5072;
assign v_5075 = v_5074 & v_4523 & v_4524;
assign v_5076 = v_5074 & v_4523 & ~v_4524;
assign v_5078 = v_5077 & ~v_4535;
assign v_5080 = v_5077 & v_5079;
assign v_5081 = v_5077 & v_4535 & v_4547 & ~v_4548 & v_4556;
assign v_5084 = v_5082 & v_5083;
assign v_5085 = v_5082 & v_4577 & v_4578;
assign v_5086 = v_5082 & v_4577 & ~v_4578 & v_4580;
assign v_5087 = v_5082 & v_4577 & ~v_4578 & ~v_4580 & v_4582;
assign v_5088 = v_5082 & v_4577 & ~v_4578 & ~v_4580 & ~v_4582;
assign v_5091 = v_5089 & v_5090;
assign v_5093 = v_5092 & ~v_4564 & v_4565 & v_4585;
assign v_5096 = v_5094 & v_5095;
assign v_5098 = v_5094 & v_5097;
assign v_5100 = ~v_5054 & v_5099;
assign v_5102 = v_5101 & v_4601 & v_4602;
assign v_5103 = v_5101 & v_4601 & ~v_4602 & v_4604;
assign v_5104 = v_5101 & v_4601 & ~v_4602 & ~v_4604 & v_4606;
assign v_5105 = v_5101 & v_4612 & v_4613;
assign v_5106 = v_5101 & v_4615 & v_4616;
assign v_5107 = v_5101 & v_4615 & ~v_4616 & v_4618;
assign v_5108 = v_5101 & v_4615 & ~v_4616 & ~v_4618 & v_4620;
assign v_5110 = v_5101 & v_5109;
assign v_5113 = v_5111 & v_5112;
assign v_5115 = v_5114 & v_4612 & ~v_4613 & v_4625 & v_4626;
assign v_5116 = v_5114 & v_4628 & v_4629;
assign v_5117 = v_5114 & v_4628 & ~v_4629 & v_4631;
assign v_5118 = v_5114 & v_4628 & ~v_4629 & ~v_4631 & v_4633;
assign v_5120 = v_5114 & v_5119;
assign v_5121 = v_7546 & v_7547;
assign v_5123 = v_5122 & v_4640 & v_4641;
assign v_5124 = v_5122 & v_4640 & ~v_4641;
assign v_5127 = v_5125 & v_5126;
assign v_5129 = v_7548 & v_7549;
assign v_5130 = v_5128 & v_4647 & v_4648;
assign v_5131 = v_5128 & v_4647 & ~v_4648 & v_4650;
assign v_5132 = v_5128 & v_4647 & ~v_4648 & ~v_4650 & v_4652;
assign v_5134 = v_5128 & v_5133;
assign v_5136 = v_7550 & v_7551;
assign v_5139 = v_5137 & v_5138;
assign v_5141 = v_5140 & v_4666 & v_4667;
assign v_5142 = v_5140 & v_4666 & ~v_4667 & v_4669;
assign v_5143 = v_5140 & v_4666 & ~v_4667 & ~v_4669 & v_4671;
assign v_5144 = v_5140 & v_4677 & v_4678;
assign v_5145 = v_5140 & v_4680 & v_4681;
assign v_5146 = v_5140 & v_4680 & ~v_4681 & v_4683;
assign v_5147 = v_5140 & v_4680 & ~v_4681 & ~v_4683 & v_4685;
assign v_5149 = v_5140 & v_5148;
assign v_5152 = v_5150 & v_5151;
assign v_5154 = v_5153 & v_4677 & ~v_4678 & v_4690 & v_4691;
assign v_5155 = v_5153 & v_4693 & v_4694;
assign v_5156 = v_5153 & v_4693 & ~v_4694 & v_4696;
assign v_5157 = v_5153 & v_4693 & ~v_4694 & ~v_4696 & v_4698;
assign v_5159 = v_5153 & v_5158;
assign v_5160 = v_7552 & v_7553;
assign v_5162 = v_5161 & v_4705 & v_4706;
assign v_5163 = v_5161 & v_4705 & ~v_4706;
assign v_5166 = v_5164 & v_5165;
assign v_5168 = v_7554 & v_7555;
assign v_5169 = v_5167 & v_4712 & v_4713;
assign v_5170 = v_5167 & v_4712 & ~v_4713 & v_4715;
assign v_5171 = v_5167 & v_4712 & ~v_4713 & ~v_4715 & v_4717;
assign v_5173 = v_5167 & v_5172;
assign v_5175 = v_7556 & v_7557;
assign v_5178 = v_5176 & v_5177;
assign v_5180 = v_5179 & v_4747;
assign v_5183 = v_5182 & ~v_5179;
assign v_5185 = v_5184 & ~v_4747 & v_4749 & v_4782 & ~v_4784;
assign v_5186 = v_5184 & ~v_4747 & v_4749 & v_4782 & v_4784;
assign v_5187 = v_5184 & ~v_4747 & v_4749 & ~v_4782;
assign v_5188 = v_5184 & v_4750;
assign v_5189 = v_5184 & ~v_4750;
assign v_5192 = v_5190 & v_5191;
assign v_5194 = v_5190 & v_5193;
assign v_5195 = v_7558 & v_7559;
assign v_5197 = v_5196 & ~v_4747 & ~v_4749 & v_4780;
assign v_5199 = v_5181 & ~v_5198;
assign v_5201 = v_5200 & v_4787 & v_4788;
assign v_5202 = v_5200 & v_4787 & ~v_4788;
assign v_5204 = v_5203 & v_4802 & v_4803;
assign v_5205 = v_5203 & v_4810;
assign v_5207 = v_5206 & v_4814 & v_4815;
assign v_5208 = v_5206 & v_4814 & ~v_4815 & v_4817;
assign v_5210 = v_5206 & v_5209;
assign v_5213 = v_5211 & v_5212;
assign v_5215 = v_5211 & v_5214;
assign v_5217 = v_5216 & v_4844 & ~v_4845 & ~v_4847;
assign v_5218 = v_5216 & v_4849 & ~v_4850;
assign v_5219 = v_5216 & v_4849 & v_4850;
assign v_5220 = v_5216 & v_4839;
assign v_5222 = v_5221 & v_4860 & v_4861;
assign v_5223 = v_5221 & v_4868;
assign v_5225 = v_5224 & v_4872 & v_4873;
assign v_5226 = v_5224 & v_4872 & ~v_4873 & v_4875;
assign v_5228 = v_5224 & v_5227;
assign v_5231 = v_5229 & v_5230;
assign v_5233 = v_5229 & v_5232;
assign v_5235 = v_4258 & v_5234;
assign v_5236 = v_4897 & v_5216;
assign v_5237 = v_4899 & v_5203;
assign v_5238 = v_4901 & v_5203;
assign v_5239 = v_4903 & v_5203;
assign v_5240 = v_4905 & v_5203;
assign v_5241 = ~v_4905 & v_5179;
assign v_5243 = ~v_4903 & v_5242;
assign v_5245 = ~v_4901 & v_5244;
assign v_5247 = ~v_4899 & v_5246;
assign v_5249 = ~v_4897 & v_5248;
assign v_5251 = ~v_4258 & v_5250;
assign v_5253 = v_5252 & ~v_4925;
assign v_5254 = v_7560 & v_7561;
assign v_5255 = v_5252 & v_4925 & v_4926 & v_4928 & v_4930;
assign v_5256 = v_7562 & v_7563;
assign v_5258 = v_5257 & v_4935 & ~v_4936 & v_4938;
assign v_5259 = v_5257 & v_4945 & ~v_4946 & ~v_4948;
assign v_5260 = v_5257 & v_4950 & ~v_4951;
assign v_5261 = v_5257 & v_4950 & v_4951;
assign v_5262 = v_5257 & v_4940;
assign v_5265 = v_5263 & v_5264;
assign v_5268 = v_5266 & v_5267;
assign v_5269 = v_5257 & v_4935 & v_4936;
assign v_5271 = v_5252 & v_5270;
assign v_5273 = v_5272 & ~v_4961;
assign v_5274 = v_5272 & v_4966 & v_4967;
assign v_5275 = v_5272 & v_4974;
assign v_5277 = v_5276 & v_4961 & v_4978 & v_4979 & ~v_4980;
assign v_5279 = v_5276 & v_5278;
assign v_5280 = v_5276 & v_5006 & v_5007;
assign v_5281 = v_5276 & v_5006 & ~v_5007;
assign v_5283 = v_5282 & v_5019 & v_5020;
assign v_5284 = v_5282 & v_5019 & ~v_5020;
assign v_5286 = v_5285 & v_5001 & v_5014 & v_5027;
assign v_5287 = v_7564 & v_7565;
assign v_5288 = v_5276 & v_5035 & v_5036;
assign v_5289 = v_5276 & v_5043;
assign v_5292 = v_5290 & v_5291;
assign v_5296 = v_5054 & v_5295;
assign v_5297 = v_4483;
assign v_5300 = v_5299 & v_4523 & v_4524;
assign v_5301 = v_5299 & v_4523 & ~v_4524;
assign v_5303 = v_5302 & ~v_4535;
assign v_5305 = v_5302 & v_5304;
assign v_5306 = v_5302 & v_4535 & v_4547 & ~v_4548 & v_4556;
assign v_5309 = v_5307 & v_5308;
assign v_5310 = v_5307 & v_4577 & v_4578;
assign v_5311 = v_5307 & v_4577 & ~v_4578 & v_4580;
assign v_5312 = v_5307 & v_4577 & ~v_4578 & ~v_4580 & v_4582;
assign v_5313 = v_5307 & v_4577 & ~v_4578 & ~v_4580 & ~v_4582;
assign v_5315 = v_5314 & v_5090;
assign v_5317 = v_5316 & ~v_4564 & v_4565 & v_4585;
assign v_5320 = v_5318 & v_5319;
assign v_5321 = v_5318 & v_5097;
assign v_5323 = ~v_5054 & v_5322;
assign v_5325 = v_5324 & v_4601 & v_4602;
assign v_5326 = v_5324 & v_4601 & ~v_4602 & v_4604;
assign v_5327 = v_5324 & v_4601 & ~v_4602 & ~v_4604 & v_4606;
assign v_5328 = v_5324 & v_4612 & v_4613;
assign v_5329 = v_5324 & v_4615 & v_4616;
assign v_5330 = v_5324 & v_4615 & ~v_4616 & v_4618;
assign v_5331 = v_5324 & v_4615 & ~v_4616 & ~v_4618 & v_4620;
assign v_5332 = v_5324 & v_5109;
assign v_5334 = v_5333 & v_5112;
assign v_5336 = v_5335 & v_4612 & ~v_4613 & v_4625 & v_4626;
assign v_5337 = v_5335 & v_4628 & v_4629;
assign v_5338 = v_5335 & v_4628 & ~v_4629 & v_4631;
assign v_5339 = v_5335 & v_4628 & ~v_4629 & ~v_4631 & v_4633;
assign v_5341 = v_5335 & v_5340;
assign v_5342 = v_7566 & v_7567;
assign v_5344 = v_5343 & v_4640 & v_4641;
assign v_5345 = v_5343 & v_4640 & ~v_4641;
assign v_5347 = v_5346 & v_5126;
assign v_5349 = v_7568 & v_7569;
assign v_5350 = v_5348 & v_4647 & v_4648;
assign v_5351 = v_5348 & v_4647 & ~v_4648 & v_4650;
assign v_5352 = v_5348 & v_4647 & ~v_4648 & ~v_4650 & v_4652;
assign v_5353 = v_5348 & v_5133;
assign v_5355 = v_7570 & v_7571;
assign v_5357 = v_5356 & v_5138;
assign v_5359 = v_5358 & v_4666 & v_4667;
assign v_5360 = v_5358 & v_4666 & ~v_4667 & v_4669;
assign v_5361 = v_5358 & v_4666 & ~v_4667 & ~v_4669 & v_4671;
assign v_5362 = v_5358 & v_4677 & v_4678;
assign v_5363 = v_5358 & v_4680 & v_4681;
assign v_5364 = v_5358 & v_4680 & ~v_4681 & v_4683;
assign v_5365 = v_5358 & v_4680 & ~v_4681 & ~v_4683 & v_4685;
assign v_5366 = v_5358 & v_5148;
assign v_5368 = v_5367 & v_5151;
assign v_5370 = v_5369 & v_4677 & ~v_4678 & v_4690 & v_4691;
assign v_5371 = v_5369 & v_4693 & v_4694;
assign v_5372 = v_5369 & v_4693 & ~v_4694 & v_4696;
assign v_5373 = v_5369 & v_4693 & ~v_4694 & ~v_4696 & v_4698;
assign v_5375 = v_5369 & v_5374;
assign v_5376 = v_7572 & v_7573;
assign v_5378 = v_5377 & v_4705 & v_4706;
assign v_5379 = v_5377 & v_4705 & ~v_4706;
assign v_5381 = v_5380 & v_5165;
assign v_5383 = v_7574 & v_7575;
assign v_5384 = v_5382 & v_4712 & v_4713;
assign v_5385 = v_5382 & v_4712 & ~v_4713 & v_4715;
assign v_5386 = v_5382 & v_4712 & ~v_4713 & ~v_4715 & v_4717;
assign v_5387 = v_5382 & v_5172;
assign v_5389 = v_7576 & v_7577;
assign v_5391 = v_5390 & v_5177;
assign v_5393 = v_5392 & v_4747;
assign v_5396 = v_5395 & v_4787 & v_4788;
assign v_5397 = v_5395 & v_4787 & ~v_4788;
assign v_5399 = v_5398 & v_4802 & v_4803;
assign v_5400 = v_5398 & v_4810;
assign v_5402 = v_5401 & v_4814 & v_4815;
assign v_5403 = v_5401 & v_4814 & ~v_4815 & v_4817;
assign v_5404 = v_5401 & v_5209;
assign v_5407 = v_5405 & v_5406;
assign v_5408 = v_5405 & v_5214;
assign v_5410 = v_5409 & v_4844 & ~v_4845 & ~v_4847;
assign v_5411 = v_5409 & v_4849 & ~v_4850;
assign v_5412 = v_5409 & v_4849 & v_4850;
assign v_5413 = v_5409 & v_4839;
assign v_5415 = v_5414 & v_4860 & v_4861;
assign v_5416 = v_5414 & v_4868;
assign v_5418 = v_5417 & v_4872 & v_4873;
assign v_5419 = v_5417 & v_4872 & ~v_4873 & v_4875;
assign v_5420 = v_5417 & v_5227;
assign v_5423 = v_5421 & v_5422;
assign v_5424 = v_5421 & v_5232;
assign v_5426 = v_4258 & v_5425;
assign v_5427 = v_4897 & v_5409;
assign v_5428 = v_4899 & v_5398;
assign v_5429 = v_4901 & v_5398;
assign v_5430 = v_4903 & v_5398;
assign v_5431 = v_4905 & v_5398;
assign v_5432 = ~v_4905 & v_5392;
assign v_5434 = ~v_4903 & v_5433;
assign v_5436 = ~v_4901 & v_5435;
assign v_5438 = ~v_4899 & v_5437;
assign v_5440 = ~v_4897 & v_5439;
assign v_5442 = ~v_4258 & v_5441;
assign v_5444 = v_5443 & ~v_4925;
assign v_5445 = v_7578 & v_7579;
assign v_5446 = v_5443 & v_4925 & v_4926 & v_4928 & v_4930;
assign v_5447 = v_7580 & v_7581;
assign v_5449 = v_5448 & v_4935 & ~v_4936 & v_4938;
assign v_5450 = v_5448 & v_4945 & ~v_4946 & ~v_4948;
assign v_5451 = v_5448 & v_4950 & ~v_4951;
assign v_5452 = v_5448 & v_4950 & v_4951;
assign v_5453 = v_5448 & v_4940;
assign v_5455 = v_5454 & v_5264;
assign v_5457 = v_5456 & v_5267;
assign v_5458 = v_5448 & v_4935 & v_4936;
assign v_5459 = v_5443 & v_5270;
assign v_5461 = v_5460 & ~v_4961;
assign v_5462 = v_5460 & v_4966 & v_4967;
assign v_5463 = v_5460 & v_4974;
assign v_5465 = v_5464 & v_4961 & v_4978 & v_4979 & ~v_4980;
assign v_5467 = v_5464 & v_5466;
assign v_5468 = v_5464 & v_5006 & v_5007;
assign v_5469 = v_5464 & v_5006 & ~v_5007;
assign v_5471 = v_5470 & v_5019 & v_5020;
assign v_5472 = v_5470 & v_5019 & ~v_5020;
assign v_5474 = v_5473 & v_5001 & v_5014 & v_5027;
assign v_5475 = v_7582 & v_7583;
assign v_5476 = v_5464 & v_5035 & v_5036;
assign v_5477 = v_5464 & v_5043;
assign v_5479 = v_5478 & v_5291;
assign v_5481 = v_4264 & v_4483;
assign v_5482 = v_4264 & ~v_4483 & v_4485 & v_4518 & ~v_4520;
assign v_5483 = v_4264 & ~v_4483 & v_4485 & v_4518 & v_4520;
assign v_5484 = v_4264 & ~v_4483 & v_4485 & ~v_4518;
assign v_5485 = v_4264 & v_4486;
assign v_5486 = v_4264 & ~v_4486;
assign v_5489 = v_5487 & v_5488;
assign v_5490 = v_5487 & v_5067;
assign v_5491 = v_7584 & v_7585;
assign v_5493 = v_5492 & ~v_4483 & ~v_4485 & v_4516;
assign v_5495 = v_5494 & v_4523 & v_4524;
assign v_5496 = v_5494 & v_4523 & ~v_4524;
assign v_5498 = v_5497 & ~v_4535;
assign v_5500 = v_5497 & v_5499;
assign v_5501 = v_5497 & v_4535 & v_4547 & ~v_4548 & v_4556;
assign v_5504 = v_5502 & v_5503;
assign v_5505 = v_5502 & v_4577 & v_4578;
assign v_5506 = v_5502 & v_4577 & ~v_4578 & v_4580;
assign v_5507 = v_5502 & v_4577 & ~v_4578 & ~v_4580 & v_4582;
assign v_5508 = v_5502 & v_4577 & ~v_4578 & ~v_4580 & ~v_4582;
assign v_5510 = v_5509 & v_5090;
assign v_5512 = v_5511 & ~v_4564 & v_4565 & v_4585;
assign v_5515 = v_5513 & v_5514;
assign v_5516 = v_5513 & v_5097;
assign v_5518 = v_5517 & v_4601 & v_4602;
assign v_5519 = v_5517 & v_4601 & ~v_4602 & v_4604;
assign v_5520 = v_5517 & v_4601 & ~v_4602 & ~v_4604 & v_4606;
assign v_5521 = v_5517 & v_4612 & v_4613;
assign v_5522 = v_5517 & v_4615 & v_4616;
assign v_5523 = v_5517 & v_4615 & ~v_4616 & v_4618;
assign v_5524 = v_5517 & v_4615 & ~v_4616 & ~v_4618 & v_4620;
assign v_5525 = v_5517 & v_5109;
assign v_5527 = v_5526 & v_5112;
assign v_5529 = v_5528 & v_4612 & ~v_4613 & v_4625 & v_4626;
assign v_5530 = v_5528 & v_4628 & v_4629;
assign v_5531 = v_5528 & v_4628 & ~v_4629 & v_4631;
assign v_5532 = v_5528 & v_4628 & ~v_4629 & ~v_4631 & v_4633;
assign v_5534 = v_5528 & v_5533;
assign v_5535 = v_7586 & v_7587;
assign v_5537 = v_5536 & v_4640 & v_4641;
assign v_5538 = v_5536 & v_4640 & ~v_4641;
assign v_5540 = v_5539 & v_5126;
assign v_5542 = v_7588 & v_7589;
assign v_5543 = v_5541 & v_4647 & v_4648;
assign v_5544 = v_5541 & v_4647 & ~v_4648 & v_4650;
assign v_5545 = v_5541 & v_4647 & ~v_4648 & ~v_4650 & v_4652;
assign v_5546 = v_5541 & v_5133;
assign v_5548 = v_7590 & v_7591;
assign v_5550 = v_5549 & v_5138;
assign v_5552 = v_5551 & v_4666 & v_4667;
assign v_5553 = v_5551 & v_4666 & ~v_4667 & v_4669;
assign v_5554 = v_5551 & v_4666 & ~v_4667 & ~v_4669 & v_4671;
assign v_5555 = v_5551 & v_4677 & v_4678;
assign v_5556 = v_5551 & v_4680 & v_4681;
assign v_5557 = v_5551 & v_4680 & ~v_4681 & v_4683;
assign v_5558 = v_5551 & v_4680 & ~v_4681 & ~v_4683 & v_4685;
assign v_5559 = v_5551 & v_5148;
assign v_5561 = v_5560 & v_5151;
assign v_5563 = v_5562 & v_4677 & ~v_4678 & v_4690 & v_4691;
assign v_5564 = v_5562 & v_4693 & v_4694;
assign v_5565 = v_5562 & v_4693 & ~v_4694 & v_4696;
assign v_5566 = v_5562 & v_4693 & ~v_4694 & ~v_4696 & v_4698;
assign v_5568 = v_5562 & v_5567;
assign v_5569 = v_7592 & v_7593;
assign v_5571 = v_5570 & v_4705 & v_4706;
assign v_5572 = v_5570 & v_4705 & ~v_4706;
assign v_5574 = v_5573 & v_5165;
assign v_5576 = v_7594 & v_7595;
assign v_5577 = v_5575 & v_4712 & v_4713;
assign v_5578 = v_5575 & v_4712 & ~v_4713 & v_4715;
assign v_5579 = v_5575 & v_4712 & ~v_4713 & ~v_4715 & v_4717;
assign v_5580 = v_5575 & v_5172;
assign v_5582 = v_7596 & v_7597;
assign v_5584 = v_5583 & v_5177;
assign v_5586 = v_5585 & v_4747;
assign v_5587 = v_5585 & ~v_4747 & v_4749 & v_4782 & ~v_4784;
assign v_5588 = v_5585 & ~v_4747 & v_4749 & v_4782 & v_4784;
assign v_5589 = v_5585 & ~v_4747 & v_4749 & ~v_4782;
assign v_5590 = v_5585 & v_4750;
assign v_5591 = v_5585 & ~v_4750;
assign v_5594 = v_5592 & v_5593;
assign v_5595 = v_5592 & v_5193;
assign v_5596 = v_7598 & v_7599;
assign v_5598 = v_5597 & ~v_4747 & ~v_4749 & v_4780;
assign v_5600 = v_5599 & v_4787 & v_4788;
assign v_5601 = v_5599 & v_4787 & ~v_4788;
assign v_5603 = v_5602 & v_4802 & v_4803;
assign v_5604 = v_5602 & v_4802 & ~v_4803 & ~v_4807;
assign v_5606 = v_5605 & v_4802 & ~v_4803 & v_4807;
assign v_5608 = v_5607 & v_4810;
assign v_5610 = v_5609 & v_4814 & v_4815;
assign v_5611 = v_5609 & v_4814 & ~v_4815 & v_4817;
assign v_5612 = v_5609 & v_5209;
assign v_5615 = v_5613 & v_5614;
assign v_5616 = v_5613 & v_5214;
assign v_5618 = v_5617 & v_4844 & ~v_4845 & ~v_4847;
assign v_5619 = v_5617 & v_4849 & ~v_4850;
assign v_5620 = v_5617 & v_4849 & v_4850;
assign v_5621 = v_5617 & v_4839;
assign v_5623 = v_5622 & v_4860 & v_4861;
assign v_5624 = v_5622 & v_4860 & ~v_4861 & ~v_4865;
assign v_5626 = v_5625 & v_4860 & ~v_4861 & v_4865;
assign v_5628 = v_5627 & v_4868;
assign v_5630 = v_5629 & v_4872 & v_4873;
assign v_5631 = v_5629 & v_4872 & ~v_4873 & v_4875;
assign v_5632 = v_5629 & v_5227;
assign v_5635 = v_5633 & v_5634;
assign v_5636 = v_5633 & v_5232;
assign v_5638 = v_4258 & v_5637;
assign v_5639 = v_4897 & v_5617;
assign v_5640 = v_4899 & v_5602;
assign v_5641 = v_4901 & v_5602;
assign v_5642 = v_4903 & v_5602;
assign v_5643 = v_4905 & v_5602;
assign v_5644 = ~v_4905 & v_5585;
assign v_5646 = ~v_4903 & v_5645;
assign v_5648 = ~v_4901 & v_5647;
assign v_5650 = ~v_4899 & v_5649;
assign v_5652 = ~v_4897 & v_5651;
assign v_5654 = ~v_4258 & v_5653;
assign v_5656 = v_5655 & ~v_4925;
assign v_5657 = v_7600 & v_7601;
assign v_5658 = v_5655 & v_4925 & v_4926 & v_4928 & v_4930;
assign v_5659 = v_7602 & v_7603;
assign v_5661 = v_5660 & v_4935 & ~v_4936 & v_4938;
assign v_5662 = v_5660 & v_4945 & ~v_4946 & ~v_4948;
assign v_5663 = v_5660 & v_4950 & ~v_4951;
assign v_5664 = v_5660 & v_4950 & v_4951;
assign v_5665 = v_5660 & v_4940;
assign v_5667 = v_5666 & v_5264;
assign v_5669 = v_5668 & v_5267;
assign v_5670 = v_5660 & v_4935 & v_4936;
assign v_5671 = v_5655 & v_5270;
assign v_5673 = v_5672 & ~v_4961;
assign v_5674 = v_5672 & v_4966 & v_4967;
assign v_5675 = v_5672 & v_4966 & ~v_4967 & ~v_4971;
assign v_5677 = v_5676 & v_4966 & ~v_4967 & v_4971;
assign v_5679 = v_5678 & v_4974;
assign v_5681 = v_5680 & v_4961 & v_4978 & v_4979 & ~v_4980;
assign v_5683 = v_5680 & v_5682;
assign v_5684 = v_5680 & v_5006 & v_5007;
assign v_5685 = v_5680 & v_5006 & ~v_5007;
assign v_5687 = v_5686 & v_5019 & v_5020;
assign v_5688 = v_5686 & v_5019 & ~v_5020;
assign v_5690 = v_5689 & v_5001 & v_5014 & v_5027;
assign v_5691 = v_7604 & v_7605;
assign v_5692 = v_5680 & v_5035 & v_5036;
assign v_5693 = v_5680 & v_5035 & ~v_5036 & ~v_5040;
assign v_5695 = v_5694 & v_5035 & ~v_5036 & v_5040;
assign v_5697 = v_5696 & v_5043;
assign v_5699 = v_5698 & v_5291;
assign v_5701 = v_4483;
assign v_5702 = ~v_4483 & v_4485 & v_4518 & ~v_4520;
assign v_5703 = ~v_4483 & v_4485 & v_4518 & v_4520;
assign v_5704 = ~v_4483 & v_4485 & ~v_4518;
assign v_5707 = v_5706;
assign v_5708 = v_5067;
assign v_5709 = v_7606 & v_7607;
assign v_5711 = v_5710 & ~v_4483 & ~v_4485 & v_4516;
assign v_5713 = v_5712 & v_4523 & v_4524;
assign v_5714 = v_5712 & v_4523 & ~v_4524;
assign v_5716 = v_5715 & ~v_4535;
assign v_5718 = v_5715 & v_5717;
assign v_5719 = v_5715 & v_4535 & v_4547 & ~v_4548 & v_4556;
assign v_5722 = v_5720 & v_5721;
assign v_5723 = v_5720 & v_4577 & v_4578;
assign v_5724 = v_5720 & v_4577 & ~v_4578 & v_4580;
assign v_5725 = v_5720 & v_4577 & ~v_4578 & ~v_4580 & v_4582;
assign v_5726 = v_5720 & v_4577 & ~v_4578 & ~v_4580 & ~v_4582;
assign v_5728 = v_5727 & v_5090;
assign v_5730 = v_5729 & ~v_4564 & v_4565 & v_4585;
assign v_5733 = v_5731 & v_5732;
assign v_5734 = v_5731 & v_5097;
assign v_5736 = v_5735 & v_4601 & v_4602;
assign v_5737 = v_5735 & v_4601 & ~v_4602 & v_4604;
assign v_5738 = v_5735 & v_4601 & ~v_4602 & ~v_4604 & v_4606;
assign v_5739 = v_5735 & v_4612 & v_4613;
assign v_5740 = v_5735 & v_4615 & v_4616;
assign v_5741 = v_5735 & v_4615 & ~v_4616 & v_4618;
assign v_5742 = v_5735 & v_4615 & ~v_4616 & ~v_4618 & v_4620;
assign v_5743 = v_5735 & v_5109;
assign v_5745 = v_5744 & v_5112;
assign v_5747 = v_5746 & v_4612 & ~v_4613 & v_4625 & v_4626;
assign v_5748 = v_5746 & v_4628 & v_4629;
assign v_5749 = v_5746 & v_4628 & ~v_4629 & v_4631;
assign v_5750 = v_5746 & v_4628 & ~v_4629 & ~v_4631 & v_4633;
assign v_5752 = v_5746 & v_5751;
assign v_5753 = v_7608 & v_7609;
assign v_5755 = v_5754 & v_4640 & v_4641;
assign v_5756 = v_5754 & v_4640 & ~v_4641;
assign v_5758 = v_5757 & v_5126;
assign v_5760 = v_7610 & v_7611;
assign v_5761 = v_5759 & v_4647 & v_4648;
assign v_5762 = v_5759 & v_4647 & ~v_4648 & v_4650;
assign v_5763 = v_5759 & v_4647 & ~v_4648 & ~v_4650 & v_4652;
assign v_5764 = v_5759 & v_5133;
assign v_5766 = v_7612 & v_7613;
assign v_5768 = v_5767 & v_5138;
assign v_5770 = v_5769 & v_4666 & v_4667;
assign v_5771 = v_5769 & v_4666 & ~v_4667 & v_4669;
assign v_5772 = v_5769 & v_4666 & ~v_4667 & ~v_4669 & v_4671;
assign v_5773 = v_5769 & v_4677 & v_4678;
assign v_5774 = v_5769 & v_4680 & v_4681;
assign v_5775 = v_5769 & v_4680 & ~v_4681 & v_4683;
assign v_5776 = v_5769 & v_4680 & ~v_4681 & ~v_4683 & v_4685;
assign v_5777 = v_5769 & v_5148;
assign v_5779 = v_5778 & v_5151;
assign v_5781 = v_5780 & v_4677 & ~v_4678 & v_4690 & v_4691;
assign v_5782 = v_5780 & v_4693 & v_4694;
assign v_5783 = v_5780 & v_4693 & ~v_4694 & v_4696;
assign v_5784 = v_5780 & v_4693 & ~v_4694 & ~v_4696 & v_4698;
assign v_5786 = v_5780 & v_5785;
assign v_5787 = v_7614 & v_7615;
assign v_5789 = v_5788 & v_4705 & v_4706;
assign v_5790 = v_5788 & v_4705 & ~v_4706;
assign v_5792 = v_5791 & v_5165;
assign v_5794 = v_7616 & v_7617;
assign v_5795 = v_5793 & v_4712 & v_4713;
assign v_5796 = v_5793 & v_4712 & ~v_4713 & v_4715;
assign v_5797 = v_5793 & v_4712 & ~v_4713 & ~v_4715 & v_4717;
assign v_5798 = v_5793 & v_5172;
assign v_5800 = v_7618 & v_7619;
assign v_5802 = v_5801 & v_5177;
assign v_5804 = v_5803 & v_4747;
assign v_5805 = v_5803 & ~v_4747 & v_4749 & v_4782 & ~v_4784;
assign v_5806 = v_5803 & ~v_4747 & v_4749 & v_4782 & v_4784;
assign v_5807 = v_5803 & ~v_4747 & v_4749 & ~v_4782;
assign v_5808 = v_5803 & v_4750;
assign v_5809 = v_5803 & ~v_4750;
assign v_5812 = v_5810 & v_5811;
assign v_5813 = v_5810 & v_5193;
assign v_5814 = v_7620 & v_7621;
assign v_5816 = v_5815 & ~v_4747 & ~v_4749 & v_4780;
assign v_5818 = v_5817 & v_4787 & v_4788;
assign v_5819 = v_5817 & v_4787 & ~v_4788;
assign v_5821 = v_5820 & v_4802 & v_4803;
assign v_5822 = v_5820 & v_4802 & ~v_4803 & ~v_4807;
assign v_5824 = v_5823 & v_4802 & ~v_4803 & v_4807;
assign v_5826 = v_5825 & v_4810;
assign v_5828 = v_5827 & v_4814 & v_4815;
assign v_5829 = v_5827 & v_4814 & ~v_4815 & v_4817;
assign v_5830 = v_5827 & v_5209;
assign v_5833 = v_5831 & v_5832;
assign v_5834 = v_5831 & v_5214;
assign v_5836 = v_5835 & v_4844 & ~v_4845 & ~v_4847;
assign v_5837 = v_5835 & v_4849 & ~v_4850;
assign v_5838 = v_5835 & v_4849 & v_4850;
assign v_5839 = v_5835 & v_4839;
assign v_5841 = v_5840 & v_4860 & v_4861;
assign v_5842 = v_5840 & v_4860 & ~v_4861 & ~v_4865;
assign v_5844 = v_5843 & v_4860 & ~v_4861 & v_4865;
assign v_5846 = v_5845 & v_4868;
assign v_5848 = v_5847 & v_4872 & v_4873;
assign v_5849 = v_5847 & v_4872 & ~v_4873 & v_4875;
assign v_5850 = v_5847 & v_5227;
assign v_5853 = v_5851 & v_5852;
assign v_5854 = v_5851 & v_5232;
assign v_5856 = v_4258 & v_5855;
assign v_5857 = v_4897 & v_5835;
assign v_5858 = v_4899 & v_5820;
assign v_5859 = v_4901 & v_5820;
assign v_5860 = v_4903 & v_5820;
assign v_5861 = v_4905 & v_5820;
assign v_5862 = ~v_4905 & v_5803;
assign v_5864 = ~v_4903 & v_5863;
assign v_5866 = ~v_4901 & v_5865;
assign v_5868 = ~v_4899 & v_5867;
assign v_5870 = ~v_4897 & v_5869;
assign v_5872 = ~v_4258 & v_5871;
assign v_5874 = v_5873 & ~v_4925;
assign v_5875 = v_7622 & v_7623;
assign v_5876 = v_5873 & v_4925 & v_4926 & v_4928 & v_4930;
assign v_5877 = v_7624 & v_7625;
assign v_5879 = v_5878 & v_4935 & ~v_4936 & v_4938;
assign v_5880 = v_5878 & v_4945 & ~v_4946 & ~v_4948;
assign v_5881 = v_5878 & v_4950 & ~v_4951;
assign v_5882 = v_5878 & v_4950 & v_4951;
assign v_5883 = v_5878 & v_4940;
assign v_5885 = v_5884 & v_5264;
assign v_5887 = v_5886 & v_5267;
assign v_5888 = v_5878 & v_4935 & v_4936;
assign v_5889 = v_5873 & v_5270;
assign v_5891 = v_5890 & ~v_4961;
assign v_5892 = v_5890 & v_4966 & v_4967;
assign v_5893 = v_5890 & v_4966 & ~v_4967 & ~v_4971;
assign v_5895 = v_5894 & v_4966 & ~v_4967 & v_4971;
assign v_5897 = v_5896 & v_4974;
assign v_5899 = v_5898 & v_4961 & v_4978 & v_4979 & ~v_4980;
assign v_5901 = v_5898 & v_5900;
assign v_5902 = v_5898 & v_5006 & v_5007;
assign v_5903 = v_5898 & v_5006 & ~v_5007;
assign v_5905 = v_5904 & v_5019 & v_5020;
assign v_5906 = v_5904 & v_5019 & ~v_5020;
assign v_5908 = v_5907 & v_5001 & v_5014 & v_5027;
assign v_5909 = v_7626 & v_7627;
assign v_5910 = v_5898 & v_5035 & v_5036;
assign v_5911 = v_5898 & v_5035 & ~v_5036 & ~v_5040;
assign v_5913 = v_5912 & v_5035 & ~v_5036 & v_5040;
assign v_5915 = v_5914 & v_5043;
assign v_5917 = v_5916 & v_5291;
assign v_5920 = v_5919 & v_4483;
assign v_5921 = v_5919 & ~v_4483 & v_4485 & v_4518 & ~v_4520;
assign v_5922 = v_5919 & ~v_4483 & v_4485 & v_4518 & v_4520;
assign v_5923 = v_5919 & ~v_4483 & v_4485 & ~v_4518;
assign v_5924 = v_5919 & v_4486;
assign v_5925 = v_5919 & ~v_4486;
assign v_5928 = v_5926 & v_5927;
assign v_5929 = v_5926 & v_5067;
assign v_5930 = v_7628 & v_7629;
assign v_5932 = v_5931 & ~v_4483 & ~v_4485 & v_4516;
assign v_5934 = v_5933 & v_4523 & v_4524;
assign v_5935 = v_5933 & v_4523 & ~v_4524;
assign v_5937 = v_5936 & ~v_4535;
assign v_5939 = v_5936 & v_5938;
assign v_5940 = v_5936 & v_4535 & v_4547 & ~v_4548 & v_4556;
assign v_5943 = v_5941 & v_5942;
assign v_5944 = v_5941 & v_4577 & v_4578;
assign v_5945 = v_5941 & v_4577 & ~v_4578 & v_4580;
assign v_5946 = v_5941 & v_4577 & ~v_4578 & ~v_4580 & v_4582;
assign v_5947 = v_5941 & v_4577 & ~v_4578 & ~v_4580 & ~v_4582;
assign v_5949 = v_5948 & v_5090;
assign v_5951 = v_5950 & ~v_4564 & v_4565 & v_4585;
assign v_5954 = v_5952 & v_5953;
assign v_5955 = v_5952 & v_5097;
assign v_5957 = v_5956 & v_4601 & v_4602;
assign v_5958 = v_5956 & v_4601 & ~v_4602 & v_4604;
assign v_5959 = v_5956 & v_4601 & ~v_4602 & ~v_4604 & v_4606;
assign v_5960 = v_5956 & v_4612 & v_4613;
assign v_5961 = v_5956 & v_4615 & v_4616;
assign v_5962 = v_5956 & v_4615 & ~v_4616 & v_4618;
assign v_5963 = v_5956 & v_4615 & ~v_4616 & ~v_4618 & v_4620;
assign v_5964 = v_5956 & v_5109;
assign v_5966 = v_5965 & v_5112;
assign v_5968 = v_5967 & v_4612 & ~v_4613 & v_4625 & v_4626;
assign v_5969 = v_5967 & v_4628 & v_4629;
assign v_5970 = v_5967 & v_4628 & ~v_4629 & v_4631;
assign v_5971 = v_5967 & v_4628 & ~v_4629 & ~v_4631 & v_4633;
assign v_5973 = v_5967 & v_5972;
assign v_5974 = v_7630 & v_7631;
assign v_5976 = v_5975 & v_4640 & v_4641;
assign v_5977 = v_5975 & v_4640 & ~v_4641;
assign v_5979 = v_5978 & v_5126;
assign v_5981 = v_7632 & v_7633;
assign v_5982 = v_5980 & v_4647 & v_4648;
assign v_5983 = v_5980 & v_4647 & ~v_4648 & v_4650;
assign v_5984 = v_5980 & v_4647 & ~v_4648 & ~v_4650 & v_4652;
assign v_5985 = v_5980 & v_5133;
assign v_5987 = v_7634 & v_7635;
assign v_5989 = v_5988 & v_5138;
assign v_5991 = v_5990 & v_4666 & v_4667;
assign v_5992 = v_5990 & v_4666 & ~v_4667 & v_4669;
assign v_5993 = v_5990 & v_4666 & ~v_4667 & ~v_4669 & v_4671;
assign v_5994 = v_5990 & v_4677 & v_4678;
assign v_5995 = v_5990 & v_4680 & v_4681;
assign v_5996 = v_5990 & v_4680 & ~v_4681 & v_4683;
assign v_5997 = v_5990 & v_4680 & ~v_4681 & ~v_4683 & v_4685;
assign v_5998 = v_5990 & v_5148;
assign v_6000 = v_5999 & v_5151;
assign v_6002 = v_6001 & v_4677 & ~v_4678 & v_4690 & v_4691;
assign v_6003 = v_6001 & v_4693 & v_4694;
assign v_6004 = v_6001 & v_4693 & ~v_4694 & v_4696;
assign v_6005 = v_6001 & v_4693 & ~v_4694 & ~v_4696 & v_4698;
assign v_6007 = v_6001 & v_6006;
assign v_6008 = v_7636 & v_7637;
assign v_6010 = v_6009 & v_4705 & v_4706;
assign v_6011 = v_6009 & v_4705 & ~v_4706;
assign v_6013 = v_6012 & v_5165;
assign v_6015 = v_7638 & v_7639;
assign v_6016 = v_6014 & v_4712 & v_4713;
assign v_6017 = v_6014 & v_4712 & ~v_4713 & v_4715;
assign v_6018 = v_6014 & v_4712 & ~v_4713 & ~v_4715 & v_4717;
assign v_6019 = v_6014 & v_5172;
assign v_6021 = v_7640 & v_7641;
assign v_6023 = v_6022 & v_5177;
assign v_6025 = v_6024 & v_4747;
assign v_6026 = v_6024 & ~v_4747 & v_4749 & v_4782 & ~v_4784;
assign v_6027 = v_6024 & ~v_4747 & v_4749 & v_4782 & v_4784;
assign v_6028 = v_6024 & ~v_4747 & v_4749 & ~v_4782;
assign v_6029 = v_6024 & v_4750;
assign v_6030 = v_6024 & ~v_4750;
assign v_6033 = v_6031 & v_6032;
assign v_6034 = v_6031 & v_5193;
assign v_6035 = v_7642 & v_7643;
assign v_6037 = v_6036 & ~v_4747 & ~v_4749 & v_4780;
assign v_6039 = v_6038 & v_4787 & v_4788;
assign v_6040 = v_6038 & v_4787 & ~v_4788;
assign v_6042 = v_6041 & v_4802 & v_4803;
assign v_6043 = v_6041 & v_4802 & ~v_4803 & ~v_4807;
assign v_6045 = v_6044 & v_4802 & ~v_4803 & v_4807;
assign v_6047 = v_6046 & v_4810;
assign v_6049 = v_6048 & v_4814 & v_4815;
assign v_6050 = v_6048 & v_4814 & ~v_4815 & v_4817;
assign v_6051 = v_6048 & v_5209;
assign v_6054 = v_6052 & v_6053;
assign v_6055 = v_6052 & v_5214;
assign v_6057 = v_6056 & v_4844 & ~v_4845 & ~v_4847;
assign v_6058 = v_6056 & v_4849 & ~v_4850;
assign v_6059 = v_6056 & v_4849 & v_4850;
assign v_6060 = v_6056 & v_4839;
assign v_6062 = v_6061 & v_4860 & v_4861;
assign v_6063 = v_6061 & v_4860 & ~v_4861 & ~v_4865;
assign v_6065 = v_6064 & v_4860 & ~v_4861 & v_4865;
assign v_6067 = v_6066 & v_4868;
assign v_6069 = v_6068 & v_4872 & v_4873;
assign v_6070 = v_6068 & v_4872 & ~v_4873 & v_4875;
assign v_6071 = v_6068 & v_5227;
assign v_6074 = v_6072 & v_6073;
assign v_6075 = v_6072 & v_5232;
assign v_6077 = v_4258 & v_6076;
assign v_6078 = v_4897 & v_6056;
assign v_6079 = v_4899 & v_6041;
assign v_6080 = v_4901 & v_6041;
assign v_6081 = v_4903 & v_6041;
assign v_6082 = v_4905 & v_6041;
assign v_6083 = ~v_4905 & v_6024;
assign v_6085 = ~v_4903 & v_6084;
assign v_6087 = ~v_4901 & v_6086;
assign v_6089 = ~v_4899 & v_6088;
assign v_6091 = ~v_4897 & v_6090;
assign v_6093 = ~v_4258 & v_6092;
assign v_6095 = v_6094 & ~v_4925;
assign v_6096 = v_7644 & v_7645;
assign v_6097 = v_6094 & v_4925 & v_4926 & v_4928 & v_4930;
assign v_6098 = v_7646 & v_7647;
assign v_6100 = v_6099 & v_4935 & ~v_4936 & v_4938;
assign v_6101 = v_6099 & v_4945 & ~v_4946 & ~v_4948;
assign v_6102 = v_6099 & v_4950 & ~v_4951;
assign v_6103 = v_6099 & v_4950 & v_4951;
assign v_6104 = v_6099 & v_4940;
assign v_6106 = v_6105 & v_5264;
assign v_6108 = v_6107 & v_5267;
assign v_6109 = v_6099 & v_4935 & v_4936;
assign v_6110 = v_6094 & v_5270;
assign v_6112 = v_6111 & ~v_4961;
assign v_6113 = v_6111 & v_4966 & v_4967;
assign v_6114 = v_6111 & v_4966 & ~v_4967 & ~v_4971;
assign v_6116 = v_6115 & v_4966 & ~v_4967 & v_4971;
assign v_6118 = v_6117 & v_4974;
assign v_6120 = v_6119 & v_4961 & v_4978 & v_4979 & ~v_4980;
assign v_6122 = v_6119 & v_6121;
assign v_6123 = v_6119 & v_5006 & v_5007;
assign v_6124 = v_6119 & v_5006 & ~v_5007;
assign v_6126 = v_6125 & v_5019 & v_5020;
assign v_6127 = v_6125 & v_5019 & ~v_5020;
assign v_6129 = v_6128 & v_5001 & v_5014 & v_5027;
assign v_6130 = v_7648 & v_7649;
assign v_6131 = v_6119 & v_5035 & v_5036;
assign v_6132 = v_6119 & v_5035 & ~v_5036 & ~v_5040;
assign v_6134 = v_6133 & v_5035 & ~v_5036 & v_5040;
assign v_6136 = v_6135 & v_5043;
assign v_6138 = v_6137 & v_5291;
assign v_6141 = v_6140 & v_4483;
assign v_6142 = v_6140 & ~v_4483 & v_4485 & v_4518 & ~v_4520;
assign v_6143 = v_6140 & ~v_4483 & v_4485 & v_4518 & v_4520;
assign v_6144 = v_6140 & ~v_4483 & v_4485 & ~v_4518;
assign v_6145 = v_6140 & v_4486;
assign v_6146 = v_6140 & ~v_4486;
assign v_6149 = v_6147 & v_6148;
assign v_6150 = v_6147 & v_5067;
assign v_6151 = v_7650 & v_7651;
assign v_6153 = v_6152 & ~v_4483 & ~v_4485 & v_4516;
assign v_6155 = v_6154 & v_4523 & v_4524;
assign v_6156 = v_6154 & v_4523 & ~v_4524;
assign v_6158 = v_6157 & ~v_4535;
assign v_6160 = v_6157 & v_6159;
assign v_6161 = v_6157 & v_4535 & v_4547 & ~v_4548 & v_4556;
assign v_6164 = v_6162 & v_6163;
assign v_6165 = v_6162 & v_4577 & v_4578;
assign v_6166 = v_6162 & v_4577 & ~v_4578 & v_4580;
assign v_6167 = v_6162 & v_4577 & ~v_4578 & ~v_4580 & v_4582;
assign v_6168 = v_6162 & v_4577 & ~v_4578 & ~v_4580 & ~v_4582;
assign v_6170 = v_6169 & v_5090;
assign v_6172 = v_6171 & ~v_4564 & v_4565 & v_4585;
assign v_6175 = v_6173 & v_6174;
assign v_6176 = v_6173 & v_5097;
assign v_6178 = v_6177 & v_4601 & v_4602;
assign v_6179 = v_6177 & v_4601 & ~v_4602 & v_4604;
assign v_6180 = v_6177 & v_4601 & ~v_4602 & ~v_4604 & v_4606;
assign v_6181 = v_6177 & v_4612 & v_4613;
assign v_6182 = v_6177 & v_4615 & v_4616;
assign v_6183 = v_6177 & v_4615 & ~v_4616 & v_4618;
assign v_6184 = v_6177 & v_4615 & ~v_4616 & ~v_4618 & v_4620;
assign v_6185 = v_6177 & v_5109;
assign v_6187 = v_6186 & v_5112;
assign v_6189 = v_6188 & v_4612 & ~v_4613 & v_4625 & v_4626;
assign v_6190 = v_6188 & v_4628 & v_4629;
assign v_6191 = v_6188 & v_4628 & ~v_4629 & v_4631;
assign v_6192 = v_6188 & v_4628 & ~v_4629 & ~v_4631 & v_4633;
assign v_6194 = v_6188 & v_6193;
assign v_6195 = v_7652 & v_7653;
assign v_6197 = v_6196 & v_4640 & v_4641;
assign v_6198 = v_6196 & v_4640 & ~v_4641;
assign v_6200 = v_6199 & v_5126;
assign v_6202 = v_7654 & v_7655;
assign v_6203 = v_6201 & v_4647 & v_4648;
assign v_6204 = v_6201 & v_4647 & ~v_4648 & v_4650;
assign v_6205 = v_6201 & v_4647 & ~v_4648 & ~v_4650 & v_4652;
assign v_6206 = v_6201 & v_5133;
assign v_6208 = v_7656 & v_7657;
assign v_6210 = v_6209 & v_5138;
assign v_6212 = v_6211 & v_4666 & v_4667;
assign v_6213 = v_6211 & v_4666 & ~v_4667 & v_4669;
assign v_6214 = v_6211 & v_4666 & ~v_4667 & ~v_4669 & v_4671;
assign v_6215 = v_6211 & v_4677 & v_4678;
assign v_6216 = v_6211 & v_4680 & v_4681;
assign v_6217 = v_6211 & v_4680 & ~v_4681 & v_4683;
assign v_6218 = v_6211 & v_4680 & ~v_4681 & ~v_4683 & v_4685;
assign v_6219 = v_6211 & v_5148;
assign v_6221 = v_6220 & v_5151;
assign v_6223 = v_6222 & v_4677 & ~v_4678 & v_4690 & v_4691;
assign v_6224 = v_6222 & v_4693 & v_4694;
assign v_6225 = v_6222 & v_4693 & ~v_4694 & v_4696;
assign v_6226 = v_6222 & v_4693 & ~v_4694 & ~v_4696 & v_4698;
assign v_6228 = v_6222 & v_6227;
assign v_6229 = v_7658 & v_7659;
assign v_6231 = v_6230 & v_4705 & v_4706;
assign v_6232 = v_6230 & v_4705 & ~v_4706;
assign v_6234 = v_6233 & v_5165;
assign v_6236 = v_7660 & v_7661;
assign v_6237 = v_6235 & v_4712 & v_4713;
assign v_6238 = v_6235 & v_4712 & ~v_4713 & v_4715;
assign v_6239 = v_6235 & v_4712 & ~v_4713 & ~v_4715 & v_4717;
assign v_6240 = v_6235 & v_5172;
assign v_6242 = v_7662 & v_7663;
assign v_6244 = v_6243 & v_5177;
assign v_6246 = v_6245 & v_4747;
assign v_6247 = v_6245 & ~v_4747 & v_4749 & v_4782 & ~v_4784;
assign v_6248 = v_6245 & ~v_4747 & v_4749 & v_4782 & v_4784;
assign v_6249 = v_6245 & ~v_4747 & v_4749 & ~v_4782;
assign v_6250 = v_6245 & v_4750;
assign v_6251 = v_6245 & ~v_4750;
assign v_6254 = v_6252 & v_6253;
assign v_6255 = v_6252 & v_5193;
assign v_6256 = v_7664 & v_7665;
assign v_6258 = v_6257 & ~v_4747 & ~v_4749 & v_4780;
assign v_6260 = v_6259 & v_4787 & v_4788;
assign v_6261 = v_6259 & v_4787 & ~v_4788;
assign v_6263 = v_6262 & v_4802 & v_4803;
assign v_6264 = v_6262 & v_4802 & ~v_4803 & ~v_4807;
assign v_6266 = v_6265 & v_4802 & ~v_4803 & v_4807;
assign v_6268 = v_6267 & v_4810;
assign v_6270 = v_6269 & v_4814 & v_4815;
assign v_6271 = v_6269 & v_4814 & ~v_4815 & v_4817;
assign v_6272 = v_6269 & v_5209;
assign v_6275 = v_6273 & v_6274;
assign v_6276 = v_6273 & v_5214;
assign v_6278 = v_6277 & v_4844 & ~v_4845 & ~v_4847;
assign v_6279 = v_6277 & v_4849 & ~v_4850;
assign v_6280 = v_6277 & v_4849 & v_4850;
assign v_6281 = v_6277 & v_4839;
assign v_6283 = v_6282 & v_4860 & v_4861;
assign v_6284 = v_6282 & v_4860 & ~v_4861 & ~v_4865;
assign v_6286 = v_6285 & v_4860 & ~v_4861 & v_4865;
assign v_6288 = v_6287 & v_4868;
assign v_6290 = v_6289 & v_4872 & v_4873;
assign v_6291 = v_6289 & v_4872 & ~v_4873 & v_4875;
assign v_6292 = v_6289 & v_5227;
assign v_6295 = v_6293 & v_6294;
assign v_6296 = v_6293 & v_5232;
assign v_6298 = v_4258 & v_6297;
assign v_6299 = v_4897 & v_6277;
assign v_6300 = v_4899 & v_6262;
assign v_6301 = v_4901 & v_6262;
assign v_6302 = v_4903 & v_6262;
assign v_6303 = v_4905 & v_6262;
assign v_6304 = ~v_4905 & v_6245;
assign v_6306 = ~v_4903 & v_6305;
assign v_6308 = ~v_4901 & v_6307;
assign v_6310 = ~v_4899 & v_6309;
assign v_6312 = ~v_4897 & v_6311;
assign v_6314 = ~v_4258 & v_6313;
assign v_6316 = v_6315 & ~v_4925;
assign v_6317 = v_7666 & v_7667;
assign v_6318 = v_6315 & v_4925 & v_4926 & v_4928 & v_4930;
assign v_6319 = v_7668 & v_7669;
assign v_6321 = v_6320 & v_4935 & ~v_4936 & v_4938;
assign v_6322 = v_6320 & v_4945 & ~v_4946 & ~v_4948;
assign v_6323 = v_6320 & v_4950 & ~v_4951;
assign v_6324 = v_6320 & v_4950 & v_4951;
assign v_6325 = v_6320 & v_4940;
assign v_6327 = v_6326 & v_5264;
assign v_6329 = v_6328 & v_5267;
assign v_6330 = v_6320 & v_4935 & v_4936;
assign v_6331 = v_6315 & v_5270;
assign v_6333 = v_6332 & ~v_4961;
assign v_6334 = v_6332 & v_4966 & v_4967;
assign v_6335 = v_6332 & v_4966 & ~v_4967 & ~v_4971;
assign v_6337 = v_6336 & v_4966 & ~v_4967 & v_4971;
assign v_6339 = v_6338 & v_4974;
assign v_6341 = v_6340 & v_4961 & v_4978 & v_4979 & ~v_4980;
assign v_6343 = v_6340 & v_6342;
assign v_6344 = v_6340 & v_5006 & v_5007;
assign v_6345 = v_6340 & v_5006 & ~v_5007;
assign v_6347 = v_6346 & v_5019 & v_5020;
assign v_6348 = v_6346 & v_5019 & ~v_5020;
assign v_6350 = v_6349 & v_5001 & v_5014 & v_5027;
assign v_6351 = v_7670 & v_7671;
assign v_6352 = v_6340 & v_5035 & v_5036;
assign v_6353 = v_6340 & v_5035 & ~v_5036 & ~v_5040;
assign v_6355 = v_6354 & v_5035 & ~v_5036 & v_5040;
assign v_6357 = v_6356 & v_5043;
assign v_6359 = v_6358 & v_5291;
assign v_6361 = v_4263 & v_4483;
assign v_6362 = v_4263 & ~v_4483 & v_4485 & v_4518 & ~v_4520;
assign v_6363 = v_4263 & ~v_4483 & v_4485 & v_4518 & v_4520;
assign v_6364 = v_4263 & ~v_4483 & v_4485 & ~v_4518;
assign v_6365 = v_4263 & v_4486;
assign v_6366 = v_4263 & ~v_4486;
assign v_6369 = v_6367 & v_6368;
assign v_6370 = v_6367 & v_5067;
assign v_6371 = v_7672 & v_7673;
assign v_6373 = v_6372 & ~v_4483 & ~v_4485 & v_4516;
assign v_6375 = v_6374 & v_4523 & v_4524;
assign v_6376 = v_6374 & v_4523 & ~v_4524;
assign v_6378 = v_6377 & ~v_4535;
assign v_6380 = v_6377 & v_6379;
assign v_6381 = v_6377 & v_4535 & v_4547 & ~v_4548 & v_4556;
assign v_6384 = v_6382 & v_6383;
assign v_6385 = v_6382 & v_4577 & v_4578;
assign v_6386 = v_6382 & v_4577 & ~v_4578 & v_4580;
assign v_6387 = v_6382 & v_4577 & ~v_4578 & ~v_4580 & v_4582;
assign v_6388 = v_6382 & v_4577 & ~v_4578 & ~v_4580 & ~v_4582;
assign v_6390 = v_6389 & v_5090;
assign v_6392 = v_6391 & ~v_4564 & v_4565 & v_4585;
assign v_6395 = v_6393 & v_6394;
assign v_6396 = v_6393 & v_5097;
assign v_6398 = v_6397 & v_4601 & v_4602;
assign v_6399 = v_6397 & v_4601 & ~v_4602 & v_4604;
assign v_6400 = v_6397 & v_4601 & ~v_4602 & ~v_4604 & v_4606;
assign v_6401 = v_6397 & v_4612 & v_4613;
assign v_6402 = v_6397 & v_4615 & v_4616;
assign v_6403 = v_6397 & v_4615 & ~v_4616 & v_4618;
assign v_6404 = v_6397 & v_4615 & ~v_4616 & ~v_4618 & v_4620;
assign v_6405 = v_6397 & v_5109;
assign v_6407 = v_6406 & v_5112;
assign v_6409 = v_6408 & v_4612 & ~v_4613 & v_4625 & v_4626;
assign v_6410 = v_6408 & v_4628 & v_4629;
assign v_6411 = v_6408 & v_4628 & ~v_4629 & v_4631;
assign v_6412 = v_6408 & v_4628 & ~v_4629 & ~v_4631 & v_4633;
assign v_6414 = v_6408 & v_6413;
assign v_6415 = v_7674 & v_7675;
assign v_6417 = v_6416 & v_4640 & v_4641;
assign v_6418 = v_6416 & v_4640 & ~v_4641;
assign v_6420 = v_6419 & v_5126;
assign v_6422 = v_7676 & v_7677;
assign v_6423 = v_6421 & v_4647 & v_4648;
assign v_6424 = v_6421 & v_4647 & ~v_4648 & v_4650;
assign v_6425 = v_6421 & v_4647 & ~v_4648 & ~v_4650 & v_4652;
assign v_6426 = v_6421 & v_5133;
assign v_6428 = v_7678 & v_7679;
assign v_6430 = v_6429 & v_5138;
assign v_6432 = v_6431 & v_4666 & v_4667;
assign v_6433 = v_6431 & v_4666 & ~v_4667 & v_4669;
assign v_6434 = v_6431 & v_4666 & ~v_4667 & ~v_4669 & v_4671;
assign v_6435 = v_6431 & v_4677 & v_4678;
assign v_6436 = v_6431 & v_4680 & v_4681;
assign v_6437 = v_6431 & v_4680 & ~v_4681 & v_4683;
assign v_6438 = v_6431 & v_4680 & ~v_4681 & ~v_4683 & v_4685;
assign v_6439 = v_6431 & v_5148;
assign v_6441 = v_6440 & v_5151;
assign v_6443 = v_6442 & v_4677 & ~v_4678 & v_4690 & v_4691;
assign v_6444 = v_6442 & v_4693 & v_4694;
assign v_6445 = v_6442 & v_4693 & ~v_4694 & v_4696;
assign v_6446 = v_6442 & v_4693 & ~v_4694 & ~v_4696 & v_4698;
assign v_6448 = v_6442 & v_6447;
assign v_6449 = v_7680 & v_7681;
assign v_6451 = v_6450 & v_4705 & v_4706;
assign v_6452 = v_6450 & v_4705 & ~v_4706;
assign v_6454 = v_6453 & v_5165;
assign v_6456 = v_7682 & v_7683;
assign v_6457 = v_6455 & v_4712 & v_4713;
assign v_6458 = v_6455 & v_4712 & ~v_4713 & v_4715;
assign v_6459 = v_6455 & v_4712 & ~v_4713 & ~v_4715 & v_4717;
assign v_6460 = v_6455 & v_5172;
assign v_6462 = v_7684 & v_7685;
assign v_6464 = v_6463 & v_5177;
assign v_6466 = v_6465 & v_4747;
assign v_6467 = v_6465 & ~v_4747 & v_4749 & v_4782 & ~v_4784;
assign v_6468 = v_6465 & ~v_4747 & v_4749 & v_4782 & v_4784;
assign v_6469 = v_6465 & ~v_4747 & v_4749 & ~v_4782;
assign v_6470 = v_6465 & v_4750;
assign v_6471 = v_6465 & ~v_4750;
assign v_6474 = v_6472 & v_6473;
assign v_6475 = v_6472 & v_5193;
assign v_6476 = v_7686 & v_7687;
assign v_6478 = v_6477 & ~v_4747 & ~v_4749 & v_4780;
assign v_6480 = v_6479 & v_4787 & v_4788;
assign v_6481 = v_6479 & v_4787 & ~v_4788;
assign v_6483 = v_6482 & v_4802 & v_4803;
assign v_6484 = v_6482 & v_4802 & ~v_4803 & ~v_4807;
assign v_6486 = v_6485 & v_4802 & ~v_4803 & v_4807;
assign v_6488 = v_6487 & v_4810;
assign v_6490 = v_6489 & v_4814 & v_4815;
assign v_6491 = v_6489 & v_4814 & ~v_4815 & v_4817;
assign v_6492 = v_6489 & v_5209;
assign v_6495 = v_6493 & v_6494;
assign v_6496 = v_6493 & v_5214;
assign v_6498 = v_6497 & v_4844 & ~v_4845 & ~v_4847;
assign v_6499 = v_6497 & v_4849 & ~v_4850;
assign v_6500 = v_6497 & v_4849 & v_4850;
assign v_6501 = v_6497 & v_4839;
assign v_6503 = v_6502 & v_4860 & v_4861;
assign v_6504 = v_6502 & v_4860 & ~v_4861 & ~v_4865;
assign v_6506 = v_6505 & v_4860 & ~v_4861 & v_4865;
assign v_6508 = v_6507 & v_4868;
assign v_6510 = v_6509 & v_4872 & v_4873;
assign v_6511 = v_6509 & v_4872 & ~v_4873 & v_4875;
assign v_6512 = v_6509 & v_5227;
assign v_6515 = v_6513 & v_6514;
assign v_6516 = v_6513 & v_5232;
assign v_6518 = v_4258 & v_6517;
assign v_6519 = v_4897 & v_6497;
assign v_6520 = v_4899 & v_6482;
assign v_6521 = v_4901 & v_6482;
assign v_6522 = v_4903 & v_6482;
assign v_6523 = v_4905 & v_6482;
assign v_6524 = ~v_4905 & v_6465;
assign v_6526 = ~v_4903 & v_6525;
assign v_6528 = ~v_4901 & v_6527;
assign v_6530 = ~v_4899 & v_6529;
assign v_6532 = ~v_4897 & v_6531;
assign v_6534 = ~v_4258 & v_6533;
assign v_6536 = v_6535 & ~v_4925;
assign v_6537 = v_7688 & v_7689;
assign v_6538 = v_6535 & v_4925 & v_4926 & v_4928 & v_4930;
assign v_6539 = v_7690 & v_7691;
assign v_6541 = v_6540 & v_4935 & ~v_4936 & v_4938;
assign v_6542 = v_6540 & v_4945 & ~v_4946 & ~v_4948;
assign v_6543 = v_6540 & v_4950 & ~v_4951;
assign v_6544 = v_6540 & v_4950 & v_4951;
assign v_6545 = v_6540 & v_4940;
assign v_6547 = v_6546 & v_5264;
assign v_6549 = v_6548 & v_5267;
assign v_6550 = v_6540 & v_4935 & v_4936;
assign v_6551 = v_6535 & v_5270;
assign v_6553 = v_6552 & ~v_4961;
assign v_6554 = v_6552 & v_4966 & v_4967;
assign v_6555 = v_6552 & v_4966 & ~v_4967 & ~v_4971;
assign v_6557 = v_6556 & v_4966 & ~v_4967 & v_4971;
assign v_6559 = v_6558 & v_4974;
assign v_6561 = v_6560 & v_4961 & v_4978 & v_4979 & ~v_4980;
assign v_6563 = v_6560 & v_6562;
assign v_6564 = v_6560 & v_5006 & v_5007;
assign v_6565 = v_6560 & v_5006 & ~v_5007;
assign v_6567 = v_6566 & v_5019 & v_5020;
assign v_6568 = v_6566 & v_5019 & ~v_5020;
assign v_6570 = v_6569 & v_5001 & v_5014 & v_5027;
assign v_6571 = v_7692 & v_7693;
assign v_6572 = v_6560 & v_5035 & v_5036;
assign v_6573 = v_6560 & v_5035 & ~v_5036 & ~v_5040;
assign v_6575 = v_6574 & v_5035 & ~v_5036 & v_5040;
assign v_6577 = v_6576 & v_5043;
assign v_6579 = v_6578 & v_5291;
assign v_6582 = v_6581 & v_4483;
assign v_6583 = v_6581 & ~v_4483 & v_4485 & v_4518 & ~v_4520;
assign v_6584 = v_6581 & ~v_4483 & v_4485 & v_4518 & v_4520;
assign v_6585 = v_6581 & ~v_4483 & v_4485 & ~v_4518;
assign v_6586 = v_6581 & v_4486;
assign v_6587 = v_6581 & ~v_4486;
assign v_6590 = v_6588 & v_6589;
assign v_6591 = v_6588 & v_5067;
assign v_6592 = v_7694 & v_7695;
assign v_6594 = v_6593 & ~v_4483 & ~v_4485 & v_4516;
assign v_6596 = v_6595 & v_4523 & v_4524;
assign v_6597 = v_6595 & v_4523 & ~v_4524;
assign v_6599 = v_6598 & ~v_4535;
assign v_6601 = v_6598 & v_6600;
assign v_6602 = v_6598 & v_4535 & v_4547 & ~v_4548 & v_4556;
assign v_6605 = v_6603 & v_6604;
assign v_6606 = v_6603 & v_4577 & v_4578;
assign v_6607 = v_6603 & v_4577 & ~v_4578 & v_4580;
assign v_6608 = v_6603 & v_4577 & ~v_4578 & ~v_4580 & v_4582;
assign v_6609 = v_6603 & v_4577 & ~v_4578 & ~v_4580 & ~v_4582;
assign v_6611 = v_6610 & v_5090;
assign v_6613 = v_6612 & ~v_4564 & v_4565 & v_4585;
assign v_6616 = v_6614 & v_6615;
assign v_6617 = v_6614 & v_5097;
assign v_6619 = v_6618 & v_4601 & v_4602;
assign v_6620 = v_6618 & v_4601 & ~v_4602 & v_4604;
assign v_6621 = v_6618 & v_4601 & ~v_4602 & ~v_4604 & v_4606;
assign v_6622 = v_6618 & v_4612 & v_4613;
assign v_6623 = v_6618 & v_4615 & v_4616;
assign v_6624 = v_6618 & v_4615 & ~v_4616 & v_4618;
assign v_6625 = v_6618 & v_4615 & ~v_4616 & ~v_4618 & v_4620;
assign v_6626 = v_6618 & v_5109;
assign v_6628 = v_6627 & v_5112;
assign v_6630 = v_6629 & v_4612 & ~v_4613 & v_4625 & v_4626;
assign v_6631 = v_6629 & v_4628 & v_4629;
assign v_6632 = v_6629 & v_4628 & ~v_4629 & v_4631;
assign v_6633 = v_6629 & v_4628 & ~v_4629 & ~v_4631 & v_4633;
assign v_6635 = v_6629 & v_6634;
assign v_6636 = v_7696 & v_7697;
assign v_6638 = v_6637 & v_4640 & v_4641;
assign v_6639 = v_6637 & v_4640 & ~v_4641;
assign v_6641 = v_6640 & v_5126;
assign v_6643 = v_7698 & v_7699;
assign v_6644 = v_6642 & v_4647 & v_4648;
assign v_6645 = v_6642 & v_4647 & ~v_4648 & v_4650;
assign v_6646 = v_6642 & v_4647 & ~v_4648 & ~v_4650 & v_4652;
assign v_6647 = v_6642 & v_5133;
assign v_6649 = v_7700 & v_7701;
assign v_6651 = v_6650 & v_5138;
assign v_6653 = v_6652 & v_4666 & v_4667;
assign v_6654 = v_6652 & v_4666 & ~v_4667 & v_4669;
assign v_6655 = v_6652 & v_4666 & ~v_4667 & ~v_4669 & v_4671;
assign v_6656 = v_6652 & v_4677 & v_4678;
assign v_6657 = v_6652 & v_4680 & v_4681;
assign v_6658 = v_6652 & v_4680 & ~v_4681 & v_4683;
assign v_6659 = v_6652 & v_4680 & ~v_4681 & ~v_4683 & v_4685;
assign v_6660 = v_6652 & v_5148;
assign v_6662 = v_6661 & v_5151;
assign v_6664 = v_6663 & v_4677 & ~v_4678 & v_4690 & v_4691;
assign v_6665 = v_6663 & v_4693 & v_4694;
assign v_6666 = v_6663 & v_4693 & ~v_4694 & v_4696;
assign v_6667 = v_6663 & v_4693 & ~v_4694 & ~v_4696 & v_4698;
assign v_6669 = v_6663 & v_6668;
assign v_6670 = v_7702 & v_7703;
assign v_6672 = v_6671 & v_4705 & v_4706;
assign v_6673 = v_6671 & v_4705 & ~v_4706;
assign v_6675 = v_6674 & v_5165;
assign v_6677 = v_7704 & v_7705;
assign v_6678 = v_6676 & v_4712 & v_4713;
assign v_6679 = v_6676 & v_4712 & ~v_4713 & v_4715;
assign v_6680 = v_6676 & v_4712 & ~v_4713 & ~v_4715 & v_4717;
assign v_6681 = v_6676 & v_5172;
assign v_6683 = v_7706 & v_7707;
assign v_6685 = v_6684 & v_5177;
assign v_6687 = v_6686 & v_4747;
assign v_6688 = v_6686 & ~v_4747 & v_4749 & v_4782 & ~v_4784;
assign v_6689 = v_6686 & ~v_4747 & v_4749 & v_4782 & v_4784;
assign v_6690 = v_6686 & ~v_4747 & v_4749 & ~v_4782;
assign v_6691 = v_6686 & v_4750;
assign v_6692 = v_6686 & ~v_4750;
assign v_6695 = v_6693 & v_6694;
assign v_6696 = v_6693 & v_5193;
assign v_6697 = v_7708 & v_7709;
assign v_6699 = v_6698 & ~v_4747 & ~v_4749 & v_4780;
assign v_6701 = v_6700 & v_4787 & v_4788;
assign v_6702 = v_6700 & v_4787 & ~v_4788;
assign v_6704 = v_6703 & v_4802 & v_4803;
assign v_6705 = v_6703 & v_4802 & ~v_4803 & ~v_4807;
assign v_6707 = v_6706 & v_4802 & ~v_4803 & v_4807;
assign v_6709 = v_6708 & v_4810;
assign v_6711 = v_6710 & v_4814 & v_4815;
assign v_6712 = v_6710 & v_4814 & ~v_4815 & v_4817;
assign v_6713 = v_6710 & v_5209;
assign v_6716 = v_6714 & v_6715;
assign v_6717 = v_6714 & v_5214;
assign v_6719 = v_6718 & v_4844 & ~v_4845 & ~v_4847;
assign v_6720 = v_6718 & v_4849 & ~v_4850;
assign v_6721 = v_6718 & v_4849 & v_4850;
assign v_6722 = v_6718 & v_4839;
assign v_6724 = v_6723 & v_4860 & v_4861;
assign v_6725 = v_6723 & v_4860 & ~v_4861 & ~v_4865;
assign v_6727 = v_6726 & v_4860 & ~v_4861 & v_4865;
assign v_6729 = v_6728 & v_4868;
assign v_6731 = v_6730 & v_4872 & v_4873;
assign v_6732 = v_6730 & v_4872 & ~v_4873 & v_4875;
assign v_6733 = v_6730 & v_5227;
assign v_6736 = v_6734 & v_6735;
assign v_6737 = v_6734 & v_5232;
assign v_6739 = v_4258 & v_6738;
assign v_6740 = v_4897 & v_6718;
assign v_6741 = v_4899 & v_6703;
assign v_6742 = v_4901 & v_6703;
assign v_6743 = v_4903 & v_6703;
assign v_6744 = v_4905 & v_6703;
assign v_6745 = ~v_4905 & v_6686;
assign v_6747 = ~v_4903 & v_6746;
assign v_6749 = ~v_4901 & v_6748;
assign v_6751 = ~v_4899 & v_6750;
assign v_6753 = ~v_4897 & v_6752;
assign v_6755 = ~v_4258 & v_6754;
assign v_6757 = v_6756 & ~v_4925;
assign v_6758 = v_7710 & v_7711;
assign v_6759 = v_6756 & v_4925 & v_4926 & v_4928 & v_4930;
assign v_6760 = v_7712 & v_7713;
assign v_6762 = v_6761 & v_4935 & ~v_4936 & v_4938;
assign v_6763 = v_6761 & v_4945 & ~v_4946 & ~v_4948;
assign v_6764 = v_6761 & v_4950 & ~v_4951;
assign v_6765 = v_6761 & v_4950 & v_4951;
assign v_6766 = v_6761 & v_4940;
assign v_6768 = v_6767 & v_5264;
assign v_6770 = v_6769 & v_5267;
assign v_6771 = v_6761 & v_4935 & v_4936;
assign v_6772 = v_6756 & v_5270;
assign v_6774 = v_6773 & ~v_4961;
assign v_6775 = v_6773 & v_4966 & v_4967;
assign v_6776 = v_6773 & v_4966 & ~v_4967 & ~v_4971;
assign v_6778 = v_6777 & v_4966 & ~v_4967 & v_4971;
assign v_6780 = v_6779 & v_4974;
assign v_6782 = v_6781 & v_4961 & v_4978 & v_4979 & ~v_4980;
assign v_6784 = v_6781 & v_6783;
assign v_6785 = v_6781 & v_5006 & v_5007;
assign v_6786 = v_6781 & v_5006 & ~v_5007;
assign v_6788 = v_6787 & v_5019 & v_5020;
assign v_6789 = v_6787 & v_5019 & ~v_5020;
assign v_6791 = v_6790 & v_5001 & v_5014 & v_5027;
assign v_6792 = v_7714 & v_7715;
assign v_6793 = v_6781 & v_5035 & v_5036;
assign v_6794 = v_6781 & v_5035 & ~v_5036 & ~v_5040;
assign v_6796 = v_6795 & v_5035 & ~v_5036 & v_5040;
assign v_6798 = v_6797 & v_5043;
assign v_6800 = v_6799 & v_5291;
assign v_6803 = v_6802 & ~v_5099;
assign v_6805 = v_5054 & v_6804;
assign v_6806 = v_4483;
assign v_6808 = v_6807 & v_4523 & v_4524;
assign v_6809 = v_6807 & v_4523 & ~v_4524;
assign v_6811 = v_6810 & ~v_4535;
assign v_6813 = v_6810 & v_6812;
assign v_6814 = v_6810 & v_4535 & v_4547 & ~v_4548 & v_4556;
assign v_6817 = v_6815 & v_6816;
assign v_6818 = v_6815 & v_4577 & v_4578;
assign v_6819 = v_6815 & v_4577 & ~v_4578 & v_4580;
assign v_6820 = v_6815 & v_4577 & ~v_4578 & ~v_4580 & v_4582;
assign v_6821 = v_6815 & v_4577 & ~v_4578 & ~v_4580 & ~v_4582;
assign v_6823 = v_6822 & v_5090;
assign v_6825 = v_6824 & ~v_4564 & v_4565 & v_4585;
assign v_6828 = v_6826 & v_6827;
assign v_6829 = v_6826 & v_5097;
assign v_6831 = ~v_5054 & v_6830;
assign v_6833 = v_6832 & v_4601 & v_4602;
assign v_6834 = v_6832 & v_4601 & ~v_4602 & v_4604;
assign v_6835 = v_6832 & v_4601 & ~v_4602 & ~v_4604 & v_4606;
assign v_6836 = v_6832 & v_4612 & v_4613;
assign v_6837 = v_6832 & v_4615 & v_4616;
assign v_6838 = v_6832 & v_4615 & ~v_4616 & v_4618;
assign v_6839 = v_6832 & v_4615 & ~v_4616 & ~v_4618 & v_4620;
assign v_6840 = v_6832 & v_5109;
assign v_6842 = v_6841 & v_5112;
assign v_6844 = v_6843 & v_4612 & ~v_4613 & v_4625 & v_4626;
assign v_6845 = v_6843 & v_4628 & v_4629;
assign v_6846 = v_6843 & v_4628 & ~v_4629 & v_4631;
assign v_6847 = v_6843 & v_4628 & ~v_4629 & ~v_4631 & v_4633;
assign v_6849 = v_6843 & v_6848;
assign v_6850 = v_7716 & v_7717;
assign v_6852 = v_6851 & v_4640 & v_4641;
assign v_6853 = v_6851 & v_4640 & ~v_4641;
assign v_6855 = v_6854 & v_5126;
assign v_6857 = v_7718 & v_7719;
assign v_6858 = v_6856 & v_4647 & v_4648;
assign v_6859 = v_6856 & v_4647 & ~v_4648 & v_4650;
assign v_6860 = v_6856 & v_4647 & ~v_4648 & ~v_4650 & v_4652;
assign v_6861 = v_6856 & v_5133;
assign v_6863 = v_7720 & v_7721;
assign v_6865 = v_6864 & v_5138;
assign v_6867 = v_6866 & v_4666 & v_4667;
assign v_6868 = v_6866 & v_4666 & ~v_4667 & v_4669;
assign v_6869 = v_6866 & v_4666 & ~v_4667 & ~v_4669 & v_4671;
assign v_6870 = v_6866 & v_4677 & v_4678;
assign v_6871 = v_6866 & v_4680 & v_4681;
assign v_6872 = v_6866 & v_4680 & ~v_4681 & v_4683;
assign v_6873 = v_6866 & v_4680 & ~v_4681 & ~v_4683 & v_4685;
assign v_6874 = v_6866 & v_5148;
assign v_6876 = v_6875 & v_5151;
assign v_6878 = v_6877 & v_4677 & ~v_4678 & v_4690 & v_4691;
assign v_6879 = v_6877 & v_4693 & v_4694;
assign v_6880 = v_6877 & v_4693 & ~v_4694 & v_4696;
assign v_6881 = v_6877 & v_4693 & ~v_4694 & ~v_4696 & v_4698;
assign v_6883 = v_6877 & v_6882;
assign v_6884 = v_7722 & v_7723;
assign v_6886 = v_6885 & v_4705 & v_4706;
assign v_6887 = v_6885 & v_4705 & ~v_4706;
assign v_6889 = v_6888 & v_5165;
assign v_6891 = v_7724 & v_7725;
assign v_6892 = v_6890 & v_4712 & v_4713;
assign v_6893 = v_6890 & v_4712 & ~v_4713 & v_4715;
assign v_6894 = v_6890 & v_4712 & ~v_4713 & ~v_4715 & v_4717;
assign v_6895 = v_6890 & v_5172;
assign v_6897 = v_7726 & v_7727;
assign v_6899 = v_6898 & v_5177;
assign v_6901 = v_6900 & v_4747;
assign v_6903 = v_6902 & v_4787 & v_4788;
assign v_6904 = v_6902 & v_4787 & ~v_4788;
assign v_6906 = v_6905 & v_4802 & v_4803;
assign v_6907 = v_6905 & v_4810;
assign v_6909 = v_6908 & v_4814 & v_4815;
assign v_6910 = v_6908 & v_4814 & ~v_4815 & v_4817;
assign v_6911 = v_6908 & v_5209;
assign v_6914 = v_6912 & v_6913;
assign v_6915 = v_6912 & v_5214;
assign v_6917 = v_6916 & v_4844 & ~v_4845 & ~v_4847;
assign v_6918 = v_6916 & v_4849 & ~v_4850;
assign v_6919 = v_6916 & v_4849 & v_4850;
assign v_6920 = v_6916 & v_4839;
assign v_6922 = v_6921 & v_4860 & v_4861;
assign v_6923 = v_6921 & v_4868;
assign v_6925 = v_6924 & v_4872 & v_4873;
assign v_6926 = v_6924 & v_4872 & ~v_4873 & v_4875;
assign v_6927 = v_6924 & v_5227;
assign v_6930 = v_6928 & v_6929;
assign v_6931 = v_6928 & v_5232;
assign v_6933 = v_4258 & v_6932;
assign v_6934 = v_4897 & v_6916;
assign v_6935 = v_4899 & v_6905;
assign v_6936 = v_4901 & v_6905;
assign v_6937 = v_4903 & v_6905;
assign v_6938 = v_4905 & v_6905;
assign v_6939 = ~v_4905 & v_6900;
assign v_6941 = ~v_4903 & v_6940;
assign v_6943 = ~v_4901 & v_6942;
assign v_6945 = ~v_4899 & v_6944;
assign v_6947 = ~v_4897 & v_6946;
assign v_6949 = ~v_4258 & v_6948;
assign v_6951 = v_6950 & ~v_4925;
assign v_6952 = v_7728 & v_7729;
assign v_6953 = v_6950 & v_4925 & v_4926 & v_4928 & v_4930;
assign v_6954 = v_7730 & v_7731;
assign v_6956 = v_6955 & v_4935 & ~v_4936 & v_4938;
assign v_6957 = v_6955 & v_4945 & ~v_4946 & ~v_4948;
assign v_6958 = v_6955 & v_4950 & ~v_4951;
assign v_6959 = v_6955 & v_4950 & v_4951;
assign v_6960 = v_6955 & v_4940;
assign v_6962 = v_6961 & v_5264;
assign v_6964 = v_6963 & v_5267;
assign v_6965 = v_6955 & v_4935 & v_4936;
assign v_6966 = v_6950 & v_5270;
assign v_6968 = v_6967 & ~v_4961;
assign v_6969 = v_6967 & v_4966 & v_4967;
assign v_6970 = v_6967 & v_4974;
assign v_6972 = v_6971 & v_4961 & v_4978 & v_4979 & ~v_4980;
assign v_6974 = v_6971 & v_6973;
assign v_6975 = v_6971 & v_5006 & v_5007;
assign v_6976 = v_6971 & v_5006 & ~v_5007;
assign v_6978 = v_6977 & v_5019 & v_5020;
assign v_6979 = v_6977 & v_5019 & ~v_5020;
assign v_6981 = v_6980 & v_5001 & v_5014 & v_5027;
assign v_6982 = v_7732 & v_7733;
assign v_6983 = v_6971 & v_5035 & v_5036;
assign v_6984 = v_6971 & v_5043;
assign v_6986 = v_6985 & v_5291;
assign v_6989 = v_6988 & v_4483;
assign v_6990 = v_6988 & ~v_4483 & v_4485 & v_4518 & ~v_4520;
assign v_6991 = v_6988 & ~v_4483 & v_4485 & v_4518 & v_4520;
assign v_6992 = v_6988 & ~v_4483 & v_4485 & ~v_4518;
assign v_6993 = v_6988 & v_4486;
assign v_6994 = v_6988 & ~v_4486;
assign v_6997 = v_6995 & v_6996;
assign v_6998 = v_6995 & v_5067;
assign v_6999 = v_7734 & v_7735;
assign v_7001 = v_7000 & ~v_4483 & ~v_4485 & v_4516;
assign v_7003 = v_7002 & v_4523 & v_4524;
assign v_7004 = v_7002 & v_4523 & ~v_4524;
assign v_7006 = v_7005 & ~v_4535;
assign v_7008 = v_7005 & v_7007;
assign v_7009 = v_7005 & v_4535 & v_4547 & ~v_4548 & v_4556;
assign v_7012 = v_7010 & v_7011;
assign v_7013 = v_7010 & v_4577 & v_4578;
assign v_7014 = v_7010 & v_4577 & ~v_4578 & v_4580;
assign v_7015 = v_7010 & v_4577 & ~v_4578 & ~v_4580 & v_4582;
assign v_7016 = v_7010 & v_4577 & ~v_4578 & ~v_4580 & ~v_4582;
assign v_7018 = v_7017 & v_5090;
assign v_7020 = v_7019 & ~v_4564 & v_4565 & v_4585;
assign v_7023 = v_7021 & v_7022;
assign v_7024 = v_7021 & v_5097;
assign v_7026 = v_7025 & v_4601 & v_4602;
assign v_7027 = v_7025 & v_4601 & ~v_4602 & v_4604;
assign v_7028 = v_7025 & v_4601 & ~v_4602 & ~v_4604 & v_4606;
assign v_7029 = v_7025 & v_4612 & v_4613;
assign v_7030 = v_7025 & v_4615 & v_4616;
assign v_7031 = v_7025 & v_4615 & ~v_4616 & v_4618;
assign v_7032 = v_7025 & v_4615 & ~v_4616 & ~v_4618 & v_4620;
assign v_7033 = v_7025 & v_5109;
assign v_7035 = v_7034 & v_5112;
assign v_7037 = v_7036 & v_4612 & ~v_4613 & v_4625 & v_4626;
assign v_7038 = v_7036 & v_4628 & v_4629;
assign v_7039 = v_7036 & v_4628 & ~v_4629 & v_4631;
assign v_7040 = v_7036 & v_4628 & ~v_4629 & ~v_4631 & v_4633;
assign v_7042 = v_7036 & v_7041;
assign v_7043 = v_7736 & v_7737;
assign v_7045 = v_7044 & v_4640 & v_4641;
assign v_7046 = v_7044 & v_4640 & ~v_4641;
assign v_7048 = v_7047 & v_5126;
assign v_7050 = v_7738 & v_7739;
assign v_7051 = v_7049 & v_4647 & v_4648;
assign v_7052 = v_7049 & v_4647 & ~v_4648 & v_4650;
assign v_7053 = v_7049 & v_4647 & ~v_4648 & ~v_4650 & v_4652;
assign v_7054 = v_7049 & v_5133;
assign v_7056 = v_7740 & v_7741;
assign v_7058 = v_7057 & v_5138;
assign v_7060 = v_7059 & v_4666 & v_4667;
assign v_7061 = v_7059 & v_4666 & ~v_4667 & v_4669;
assign v_7062 = v_7059 & v_4666 & ~v_4667 & ~v_4669 & v_4671;
assign v_7063 = v_7059 & v_4677 & v_4678;
assign v_7064 = v_7059 & v_4680 & v_4681;
assign v_7065 = v_7059 & v_4680 & ~v_4681 & v_4683;
assign v_7066 = v_7059 & v_4680 & ~v_4681 & ~v_4683 & v_4685;
assign v_7067 = v_7059 & v_5148;
assign v_7069 = v_7068 & v_5151;
assign v_7071 = v_7070 & v_4677 & ~v_4678 & v_4690 & v_4691;
assign v_7072 = v_7070 & v_4693 & v_4694;
assign v_7073 = v_7070 & v_4693 & ~v_4694 & v_4696;
assign v_7074 = v_7070 & v_4693 & ~v_4694 & ~v_4696 & v_4698;
assign v_7076 = v_7070 & v_7075;
assign v_7077 = v_7742 & v_7743;
assign v_7079 = v_7078 & v_4705 & v_4706;
assign v_7080 = v_7078 & v_4705 & ~v_4706;
assign v_7082 = v_7081 & v_5165;
assign v_7084 = v_7744 & v_7745;
assign v_7085 = v_7083 & v_4712 & v_4713;
assign v_7086 = v_7083 & v_4712 & ~v_4713 & v_4715;
assign v_7087 = v_7083 & v_4712 & ~v_4713 & ~v_4715 & v_4717;
assign v_7088 = v_7083 & v_5172;
assign v_7090 = v_7746 & v_7747;
assign v_7092 = v_7091 & v_5177;
assign v_7094 = v_7093 & v_4747;
assign v_7095 = v_7093 & ~v_4747 & v_4749 & v_4782 & ~v_4784;
assign v_7096 = v_7093 & ~v_4747 & v_4749 & v_4782 & v_4784;
assign v_7097 = v_7093 & ~v_4747 & v_4749 & ~v_4782;
assign v_7098 = v_7093 & v_4750;
assign v_7099 = v_7093 & ~v_4750;
assign v_7102 = v_7100 & v_7101;
assign v_7103 = v_7100 & v_5193;
assign v_7104 = v_7748 & v_7749;
assign v_7106 = v_7105 & ~v_4747 & ~v_4749 & v_4780;
assign v_7108 = v_7107 & v_4787 & v_4788;
assign v_7109 = v_7107 & v_4787 & ~v_4788;
assign v_7111 = v_7110 & v_4802 & v_4803;
assign v_7112 = v_7110 & v_4802 & ~v_4803 & ~v_4807;
assign v_7114 = v_7113 & v_4802 & ~v_4803 & v_4807;
assign v_7116 = v_7115 & v_4810;
assign v_7118 = v_7117 & v_4814 & v_4815;
assign v_7119 = v_7117 & v_4814 & ~v_4815 & v_4817;
assign v_7120 = v_7117 & v_5209;
assign v_7123 = v_7121 & v_7122;
assign v_7124 = v_7121 & v_5214;
assign v_7126 = v_7125 & v_4844 & ~v_4845 & ~v_4847;
assign v_7127 = v_7125 & v_4849 & ~v_4850;
assign v_7128 = v_7125 & v_4849 & v_4850;
assign v_7129 = v_7125 & v_4839;
assign v_7131 = v_7130 & v_4860 & v_4861;
assign v_7132 = v_7130 & v_4860 & ~v_4861 & ~v_4865;
assign v_7134 = v_7133 & v_4860 & ~v_4861 & v_4865;
assign v_7136 = v_7135 & v_4868;
assign v_7138 = v_7137 & v_4872 & v_4873;
assign v_7139 = v_7137 & v_4872 & ~v_4873 & v_4875;
assign v_7140 = v_7137 & v_5227;
assign v_7143 = v_7141 & v_7142;
assign v_7144 = v_7141 & v_5232;
assign v_7146 = v_4258 & v_7145;
assign v_7147 = v_4897 & v_7125;
assign v_7148 = v_4899 & v_7110;
assign v_7149 = v_4901 & v_7110;
assign v_7150 = v_4903 & v_7110;
assign v_7151 = v_4905 & v_7110;
assign v_7152 = ~v_4905 & v_7093;
assign v_7154 = ~v_4903 & v_7153;
assign v_7156 = ~v_4901 & v_7155;
assign v_7158 = ~v_4899 & v_7157;
assign v_7160 = ~v_4897 & v_7159;
assign v_7162 = ~v_4258 & v_7161;
assign v_7164 = v_7163 & ~v_4925;
assign v_7165 = v_7750 & v_7751;
assign v_7166 = v_7163 & v_4925 & v_4926 & v_4928 & v_4930;
assign v_7167 = v_7752 & v_7753;
assign v_7169 = v_7168 & v_4935 & ~v_4936 & v_4938;
assign v_7170 = v_7168 & v_4945 & ~v_4946 & ~v_4948;
assign v_7171 = v_7168 & v_4950 & ~v_4951;
assign v_7172 = v_7168 & v_4950 & v_4951;
assign v_7173 = v_7168 & v_4940;
assign v_7175 = v_7174 & v_5264;
assign v_7177 = v_7176 & v_5267;
assign v_7178 = v_7168 & v_4935 & v_4936;
assign v_7179 = v_7163 & v_5270;
assign v_7181 = v_7180 & ~v_4961;
assign v_7182 = v_7180 & v_4966 & v_4967;
assign v_7183 = v_7180 & v_4966 & ~v_4967 & ~v_4971;
assign v_7185 = v_7184 & v_4966 & ~v_4967 & v_4971;
assign v_7187 = v_7186 & v_4974;
assign v_7189 = v_7188 & v_4961 & v_4978 & v_4979 & ~v_4980;
assign v_7191 = v_7188 & v_7190;
assign v_7192 = v_7188 & v_5006 & v_5007;
assign v_7193 = v_7188 & v_5006 & ~v_5007;
assign v_7195 = v_7194 & v_5019 & v_5020;
assign v_7196 = v_7194 & v_5019 & ~v_5020;
assign v_7198 = v_7197 & v_5001 & v_5014 & v_5027;
assign v_7199 = v_7754 & v_7755;
assign v_7200 = v_7188 & v_5035 & v_5036;
assign v_7201 = v_7188 & v_5035 & ~v_5036 & ~v_5040;
assign v_7203 = v_7202 & v_5035 & ~v_5036 & v_5040;
assign v_7205 = v_7204 & v_5043;
assign v_7207 = v_7206 & v_5291;
assign v_7219 = v_7756 & v_7757 & v_7758;
assign v_7220 = v_232 & ~v_234 & v_236 & ~v_237 & v_239;
assign v_7221 = v_245;
assign v_7222 = v_232 & ~v_234 & v_236 & ~v_237 & v_239;
assign v_7223 = ~v_245 & v_247;
assign v_7224 = v_232 & ~v_234 & ~v_236 & v_241 & ~v_243;
assign v_7225 = v_251;
assign v_7226 = v_232 & ~v_234 & ~v_236 & v_241 & ~v_243;
assign v_7227 = ~v_251;
assign v_7228 = v_232 & ~v_234 & v_236 & ~v_237 & v_239;
assign v_7229 = ~v_245 & ~v_247 & v_258;
assign v_7230 = v_345 & ~v_346 & ~v_348 & ~v_350 & ~v_352;
assign v_7231 = ~v_354;
assign v_7232 = v_372 & ~v_373 & ~v_375 & ~v_377 & ~v_379;
assign v_7233 = v_381;
assign v_7234 = v_372 & ~v_373 & ~v_375 & ~v_377 & ~v_379;
assign v_7235 = ~v_381;
assign v_7236 = v_356 & ~v_357 & v_369 & ~v_370 & v_388;
assign v_7237 = v_389;
assign v_7238 = v_391 & ~v_392 & ~v_394 & ~v_396 & v_398;
assign v_7239 = v_400;
assign v_7240 = v_391 & ~v_392 & ~v_394 & ~v_396 & v_398;
assign v_7241 = ~v_400;
assign v_7242 = v_356 & ~v_357 & v_369 & ~v_370 & v_388;
assign v_7243 = ~v_389 & v_403;
assign v_7244 = v_410 & ~v_411 & ~v_413 & ~v_415 & ~v_417;
assign v_7245 = ~v_419;
assign v_7246 = v_437 & ~v_438 & ~v_440 & ~v_442 & ~v_444;
assign v_7247 = v_446;
assign v_7248 = v_437 & ~v_438 & ~v_440 & ~v_442 & ~v_444;
assign v_7249 = ~v_446;
assign v_7250 = v_421 & ~v_422 & v_434 & ~v_435 & v_453;
assign v_7251 = v_454;
assign v_7252 = v_456 & ~v_457 & ~v_459 & ~v_461 & v_463;
assign v_7253 = v_465;
assign v_7254 = v_456 & ~v_457 & ~v_459 & ~v_461 & v_463;
assign v_7255 = ~v_465;
assign v_7256 = v_421 & ~v_422 & v_434 & ~v_435 & v_453;
assign v_7257 = ~v_454 & v_468;
assign v_7258 = v_496 & ~v_498 & v_500 & ~v_501 & v_503;
assign v_7259 = v_509;
assign v_7260 = v_496 & ~v_498 & v_500 & ~v_501 & v_503;
assign v_7261 = ~v_509 & v_511;
assign v_7262 = v_496 & ~v_498 & ~v_500 & v_505 & ~v_507;
assign v_7263 = v_515;
assign v_7264 = v_496 & ~v_498 & ~v_500 & v_505 & ~v_507;
assign v_7265 = ~v_515;
assign v_7266 = v_496 & ~v_498 & v_500 & ~v_501 & v_503;
assign v_7267 = ~v_509 & ~v_511 & v_522;
assign v_7268 = v_705 & v_722 & v_723 & v_724 & ~v_726;
assign v_7269 = v_729;
assign v_7270 = v_705 & v_722 & v_723 & v_724 & ~v_726;
assign v_7271 = ~v_729 & ~v_731;
assign v_7272 = v_705 & v_722 & v_723 & v_724 & ~v_726;
assign v_7273 = ~v_729 & v_731 & ~v_733;
assign v_7274 = v_705 & v_722 & v_723 & v_724 & ~v_726;
assign v_7275 = ~v_729 & v_731 & v_733 & v_735;
assign v_7276 = v_258 & v_232 & ~v_234 & v_236 & ~v_237;
assign v_7277 = v_239 & ~v_245 & ~v_247;
assign v_7278 = v_1101 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_7279 = ~v_379 & ~v_381;
assign v_7280 = v_1115 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7281 = v_388 & v_389;
assign v_7282 = v_1122 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7283 = v_388 & ~v_389 & v_403;
assign v_7284 = v_1140 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_7285 = ~v_444 & ~v_446;
assign v_7286 = v_1154 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7287 = v_453 & v_454;
assign v_7288 = v_1161 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7289 = v_453 & ~v_454 & v_468;
assign v_7290 = v_1177 & v_496 & ~v_498 & v_500 & ~v_501;
assign v_7291 = v_503 & ~v_509 & ~v_511 & v_522;
assign v_7292 = v_1239 & v_669 & v_670 & v_672 & ~v_674;
assign v_7293 = ~v_675;
assign v_7294 = v_1239 & v_669 & v_670 & v_672 & ~v_674;
assign v_7295 = v_675;
assign v_7296 = v_1263 & v_705 & v_722 & v_723 & v_724;
assign v_7297 = v_726;
assign v_7298 = v_1439 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_7299 = ~v_379 & ~v_381;
assign v_7300 = v_1452 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7301 = v_388 & v_389;
assign v_7302 = v_1458 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7303 = v_388 & ~v_389 & v_403;
assign v_7304 = v_1473 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_7305 = ~v_444 & ~v_446;
assign v_7306 = v_1486 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7307 = v_453 & v_454;
assign v_7308 = v_1492 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7309 = v_453 & ~v_454 & v_468;
assign v_7310 = v_1547 & v_669 & v_670 & v_672 & ~v_674;
assign v_7311 = ~v_675;
assign v_7312 = v_1547 & v_669 & v_670 & v_672 & ~v_674;
assign v_7313 = v_675;
assign v_7314 = v_1568 & v_705 & v_722 & v_723 & v_724;
assign v_7315 = v_726;
assign v_7316 = v_1696 & v_232 & ~v_234 & v_236 & ~v_237;
assign v_7317 = v_239 & ~v_245 & ~v_247 & v_258;
assign v_7318 = v_1737 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_7319 = ~v_379 & ~v_381;
assign v_7320 = v_1750 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7321 = v_388 & v_389;
assign v_7322 = v_1756 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7323 = v_388 & ~v_389 & v_403;
assign v_7324 = v_1771 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_7325 = ~v_444 & ~v_446;
assign v_7326 = v_1784 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7327 = v_453 & v_454;
assign v_7328 = v_1790 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7329 = v_453 & ~v_454 & v_468;
assign v_7330 = v_1801 & v_496 & ~v_498 & v_500 & ~v_501;
assign v_7331 = v_503 & ~v_509 & ~v_511 & v_522;
assign v_7332 = v_1864 & v_669 & v_670 & v_672 & ~v_674;
assign v_7333 = ~v_675;
assign v_7334 = v_1864 & v_669 & v_670 & v_672 & ~v_674;
assign v_7335 = v_675;
assign v_7336 = v_1889 & v_705 & v_722 & v_723 & v_724;
assign v_7337 = v_726;
assign v_7338 = v_258 & v_232 & ~v_234 & v_236 & ~v_237;
assign v_7339 = v_239 & ~v_245 & ~v_247;
assign v_7340 = v_2060 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_7341 = ~v_379 & ~v_381;
assign v_7342 = v_2073 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7343 = v_388 & v_389;
assign v_7344 = v_2079 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7345 = v_388 & ~v_389 & v_403;
assign v_7346 = v_2094 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_7347 = ~v_444 & ~v_446;
assign v_7348 = v_2107 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7349 = v_453 & v_454;
assign v_7350 = v_2113 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7351 = v_453 & ~v_454 & v_468;
assign v_7352 = v_2124 & v_496 & ~v_498 & v_500 & ~v_501;
assign v_7353 = v_503 & ~v_509 & ~v_511 & v_522;
assign v_7354 = v_2187 & v_669 & v_670 & v_672 & ~v_674;
assign v_7355 = ~v_675;
assign v_7356 = v_2187 & v_669 & v_670 & v_672 & ~v_674;
assign v_7357 = v_675;
assign v_7358 = v_2212 & v_705 & v_722 & v_723 & v_724;
assign v_7359 = v_726;
assign v_7360 = v_2345 & v_232 & ~v_234 & v_236 & ~v_237;
assign v_7361 = v_239 & ~v_245 & ~v_247 & v_258;
assign v_7362 = v_2386 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_7363 = ~v_379 & ~v_381;
assign v_7364 = v_2399 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7365 = v_388 & v_389;
assign v_7366 = v_2405 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7367 = v_388 & ~v_389 & v_403;
assign v_7368 = v_2420 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_7369 = ~v_444 & ~v_446;
assign v_7370 = v_2433 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7371 = v_453 & v_454;
assign v_7372 = v_2439 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7373 = v_453 & ~v_454 & v_468;
assign v_7374 = v_2450 & v_496 & ~v_498 & v_500 & ~v_501;
assign v_7375 = v_503 & ~v_509 & ~v_511 & v_522;
assign v_7376 = v_2513 & v_669 & v_670 & v_672 & ~v_674;
assign v_7377 = ~v_675;
assign v_7378 = v_2513 & v_669 & v_670 & v_672 & ~v_674;
assign v_7379 = v_675;
assign v_7380 = v_2538 & v_705 & v_722 & v_723 & v_724;
assign v_7381 = v_726;
assign v_7382 = v_2671 & v_232 & ~v_234 & v_236 & ~v_237;
assign v_7383 = v_239 & ~v_245 & ~v_247 & v_258;
assign v_7384 = v_2712 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_7385 = ~v_379 & ~v_381;
assign v_7386 = v_2725 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7387 = v_388 & v_389;
assign v_7388 = v_2731 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7389 = v_388 & ~v_389 & v_403;
assign v_7390 = v_2746 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_7391 = ~v_444 & ~v_446;
assign v_7392 = v_2759 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7393 = v_453 & v_454;
assign v_7394 = v_2765 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7395 = v_453 & ~v_454 & v_468;
assign v_7396 = v_2776 & v_496 & ~v_498 & v_500 & ~v_501;
assign v_7397 = v_503 & ~v_509 & ~v_511 & v_522;
assign v_7398 = v_2839 & v_669 & v_670 & v_672 & ~v_674;
assign v_7399 = ~v_675;
assign v_7400 = v_2839 & v_669 & v_670 & v_672 & ~v_674;
assign v_7401 = v_675;
assign v_7402 = v_2864 & v_705 & v_722 & v_723 & v_724;
assign v_7403 = v_726;
assign v_7404 = v_2996 & v_232 & ~v_234 & v_236 & ~v_237;
assign v_7405 = v_239 & ~v_245 & ~v_247 & v_258;
assign v_7406 = v_3037 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_7407 = ~v_379 & ~v_381;
assign v_7408 = v_3050 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7409 = v_388 & v_389;
assign v_7410 = v_3056 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7411 = v_388 & ~v_389 & v_403;
assign v_7412 = v_3071 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_7413 = ~v_444 & ~v_446;
assign v_7414 = v_3084 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7415 = v_453 & v_454;
assign v_7416 = v_3090 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7417 = v_453 & ~v_454 & v_468;
assign v_7418 = v_3101 & v_496 & ~v_498 & v_500 & ~v_501;
assign v_7419 = v_503 & ~v_509 & ~v_511 & v_522;
assign v_7420 = v_3164 & v_669 & v_670 & v_672 & ~v_674;
assign v_7421 = ~v_675;
assign v_7422 = v_3164 & v_669 & v_670 & v_672 & ~v_674;
assign v_7423 = v_675;
assign v_7424 = v_3189 & v_705 & v_722 & v_723 & v_724;
assign v_7425 = v_726;
assign v_7426 = v_3322 & v_232 & ~v_234 & v_236 & ~v_237;
assign v_7427 = v_239 & ~v_245 & ~v_247 & v_258;
assign v_7428 = v_3363 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_7429 = ~v_379 & ~v_381;
assign v_7430 = v_3376 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7431 = v_388 & v_389;
assign v_7432 = v_3382 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7433 = v_388 & ~v_389 & v_403;
assign v_7434 = v_3397 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_7435 = ~v_444 & ~v_446;
assign v_7436 = v_3410 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7437 = v_453 & v_454;
assign v_7438 = v_3416 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7439 = v_453 & ~v_454 & v_468;
assign v_7440 = v_3427 & v_496 & ~v_498 & v_500 & ~v_501;
assign v_7441 = v_503 & ~v_509 & ~v_511 & v_522;
assign v_7442 = v_3490 & v_669 & v_670 & v_672 & ~v_674;
assign v_7443 = ~v_675;
assign v_7444 = v_3490 & v_669 & v_670 & v_672 & ~v_674;
assign v_7445 = v_675;
assign v_7446 = v_3515 & v_705 & v_722 & v_723 & v_724;
assign v_7447 = v_726;
assign v_7448 = v_3682 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_7449 = ~v_379 & ~v_381;
assign v_7450 = v_3695 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7451 = v_388 & v_389;
assign v_7452 = v_3701 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7453 = v_388 & ~v_389 & v_403;
assign v_7454 = v_3716 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_7455 = ~v_444 & ~v_446;
assign v_7456 = v_3729 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7457 = v_453 & v_454;
assign v_7458 = v_3735 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7459 = v_453 & ~v_454 & v_468;
assign v_7460 = v_3789 & v_669 & v_670 & v_672 & ~v_674;
assign v_7461 = ~v_675;
assign v_7462 = v_3789 & v_669 & v_670 & v_672 & ~v_674;
assign v_7463 = v_675;
assign v_7464 = v_3810 & v_705 & v_722 & v_723 & v_724;
assign v_7465 = v_726;
assign v_7466 = v_3939 & v_232 & ~v_234 & v_236 & ~v_237;
assign v_7467 = v_239 & ~v_245 & ~v_247 & v_258;
assign v_7468 = v_3980 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_7469 = ~v_379 & ~v_381;
assign v_7470 = v_3993 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7471 = v_388 & v_389;
assign v_7472 = v_3999 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_7473 = v_388 & ~v_389 & v_403;
assign v_7474 = v_4014 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_7475 = ~v_444 & ~v_446;
assign v_7476 = v_4027 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7477 = v_453 & v_454;
assign v_7478 = v_4033 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_7479 = v_453 & ~v_454 & v_468;
assign v_7480 = v_4044 & v_496 & ~v_498 & v_500 & ~v_501;
assign v_7481 = v_503 & ~v_509 & ~v_511 & v_522;
assign v_7482 = v_4107 & v_669 & v_670 & v_672 & ~v_674;
assign v_7483 = ~v_675;
assign v_7484 = v_4107 & v_669 & v_670 & v_672 & ~v_674;
assign v_7485 = v_675;
assign v_7486 = v_4132 & v_705 & v_722 & v_723 & v_724;
assign v_7487 = v_726;
assign v_7488 = v_4488 & ~v_4490 & v_4492 & ~v_4493 & v_4495;
assign v_7489 = v_4501;
assign v_7490 = v_4488 & ~v_4490 & v_4492 & ~v_4493 & v_4495;
assign v_7491 = ~v_4501 & v_4503;
assign v_7492 = v_4488 & ~v_4490 & ~v_4492 & v_4497 & ~v_4499;
assign v_7493 = v_4507;
assign v_7494 = v_4488 & ~v_4490 & ~v_4492 & v_4497 & ~v_4499;
assign v_7495 = ~v_4507;
assign v_7496 = v_4488 & ~v_4490 & v_4492 & ~v_4493 & v_4495;
assign v_7497 = ~v_4501 & ~v_4503 & v_4514;
assign v_7498 = v_4601 & ~v_4602 & ~v_4604 & ~v_4606 & ~v_4608;
assign v_7499 = ~v_4610;
assign v_7500 = v_4628 & ~v_4629 & ~v_4631 & ~v_4633 & ~v_4635;
assign v_7501 = v_4637;
assign v_7502 = v_4628 & ~v_4629 & ~v_4631 & ~v_4633 & ~v_4635;
assign v_7503 = ~v_4637;
assign v_7504 = v_4612 & ~v_4613 & v_4625 & ~v_4626 & v_4644;
assign v_7505 = v_4645;
assign v_7506 = v_4647 & ~v_4648 & ~v_4650 & ~v_4652 & v_4654;
assign v_7507 = v_4656;
assign v_7508 = v_4647 & ~v_4648 & ~v_4650 & ~v_4652 & v_4654;
assign v_7509 = ~v_4656;
assign v_7510 = v_4612 & ~v_4613 & v_4625 & ~v_4626 & v_4644;
assign v_7511 = ~v_4645 & v_4659;
assign v_7512 = v_4666 & ~v_4667 & ~v_4669 & ~v_4671 & ~v_4673;
assign v_7513 = ~v_4675;
assign v_7514 = v_4693 & ~v_4694 & ~v_4696 & ~v_4698 & ~v_4700;
assign v_7515 = v_4702;
assign v_7516 = v_4693 & ~v_4694 & ~v_4696 & ~v_4698 & ~v_4700;
assign v_7517 = ~v_4702;
assign v_7518 = v_4677 & ~v_4678 & v_4690 & ~v_4691 & v_4709;
assign v_7519 = v_4710;
assign v_7520 = v_4712 & ~v_4713 & ~v_4715 & ~v_4717 & v_4719;
assign v_7521 = v_4721;
assign v_7522 = v_4712 & ~v_4713 & ~v_4715 & ~v_4717 & v_4719;
assign v_7523 = ~v_4721;
assign v_7524 = v_4677 & ~v_4678 & v_4690 & ~v_4691 & v_4709;
assign v_7525 = ~v_4710 & v_4724;
assign v_7526 = v_4752 & ~v_4754 & v_4756 & ~v_4757 & v_4759;
assign v_7527 = v_4765;
assign v_7528 = v_4752 & ~v_4754 & v_4756 & ~v_4757 & v_4759;
assign v_7529 = ~v_4765 & v_4767;
assign v_7530 = v_4752 & ~v_4754 & ~v_4756 & v_4761 & ~v_4763;
assign v_7531 = v_4771;
assign v_7532 = v_4752 & ~v_4754 & ~v_4756 & v_4761 & ~v_4763;
assign v_7533 = ~v_4771;
assign v_7534 = v_4752 & ~v_4754 & v_4756 & ~v_4757 & v_4759;
assign v_7535 = ~v_4765 & ~v_4767 & v_4778;
assign v_7536 = v_4961 & v_4978 & v_4979 & v_4980 & ~v_4982;
assign v_7537 = v_4985;
assign v_7538 = v_4961 & v_4978 & v_4979 & v_4980 & ~v_4982;
assign v_7539 = ~v_4985 & ~v_4987;
assign v_7540 = v_4961 & v_4978 & v_4979 & v_4980 & ~v_4982;
assign v_7541 = ~v_4985 & v_4987 & ~v_4989;
assign v_7542 = v_4961 & v_4978 & v_4979 & v_4980 & ~v_4982;
assign v_7543 = ~v_4985 & v_4987 & v_4989 & v_4991;
assign v_7544 = v_4514 & v_4488 & ~v_4490 & v_4492 & ~v_4493;
assign v_7545 = v_4495 & ~v_4501 & ~v_4503;
assign v_7546 = v_5114 & v_4628 & ~v_4629 & ~v_4631 & ~v_4633;
assign v_7547 = ~v_4635 & ~v_4637;
assign v_7548 = v_5128 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7549 = v_4644 & v_4645;
assign v_7550 = v_5135 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7551 = v_4644 & ~v_4645 & v_4659;
assign v_7552 = v_5153 & v_4693 & ~v_4694 & ~v_4696 & ~v_4698;
assign v_7553 = ~v_4700 & ~v_4702;
assign v_7554 = v_5167 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7555 = v_4709 & v_4710;
assign v_7556 = v_5174 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7557 = v_4709 & ~v_4710 & v_4724;
assign v_7558 = v_5190 & v_4752 & ~v_4754 & v_4756 & ~v_4757;
assign v_7559 = v_4759 & ~v_4765 & ~v_4767 & v_4778;
assign v_7560 = v_5252 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7561 = ~v_4931;
assign v_7562 = v_5252 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7563 = v_4931;
assign v_7564 = v_5276 & v_4961 & v_4978 & v_4979 & v_4980;
assign v_7565 = v_4982;
assign v_7566 = v_5335 & v_4628 & ~v_4629 & ~v_4631 & ~v_4633;
assign v_7567 = ~v_4635 & ~v_4637;
assign v_7568 = v_5348 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7569 = v_4644 & v_4645;
assign v_7570 = v_5354 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7571 = v_4644 & ~v_4645 & v_4659;
assign v_7572 = v_5369 & v_4693 & ~v_4694 & ~v_4696 & ~v_4698;
assign v_7573 = ~v_4700 & ~v_4702;
assign v_7574 = v_5382 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7575 = v_4709 & v_4710;
assign v_7576 = v_5388 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7577 = v_4709 & ~v_4710 & v_4724;
assign v_7578 = v_5443 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7579 = ~v_4931;
assign v_7580 = v_5443 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7581 = v_4931;
assign v_7582 = v_5464 & v_4961 & v_4978 & v_4979 & v_4980;
assign v_7583 = v_4982;
assign v_7584 = v_5487 & v_4488 & ~v_4490 & v_4492 & ~v_4493;
assign v_7585 = v_4495 & ~v_4501 & ~v_4503 & v_4514;
assign v_7586 = v_5528 & v_4628 & ~v_4629 & ~v_4631 & ~v_4633;
assign v_7587 = ~v_4635 & ~v_4637;
assign v_7588 = v_5541 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7589 = v_4644 & v_4645;
assign v_7590 = v_5547 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7591 = v_4644 & ~v_4645 & v_4659;
assign v_7592 = v_5562 & v_4693 & ~v_4694 & ~v_4696 & ~v_4698;
assign v_7593 = ~v_4700 & ~v_4702;
assign v_7594 = v_5575 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7595 = v_4709 & v_4710;
assign v_7596 = v_5581 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7597 = v_4709 & ~v_4710 & v_4724;
assign v_7598 = v_5592 & v_4752 & ~v_4754 & v_4756 & ~v_4757;
assign v_7599 = v_4759 & ~v_4765 & ~v_4767 & v_4778;
assign v_7600 = v_5655 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7601 = ~v_4931;
assign v_7602 = v_5655 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7603 = v_4931;
assign v_7604 = v_5680 & v_4961 & v_4978 & v_4979 & v_4980;
assign v_7605 = v_4982;
assign v_7606 = v_4514 & v_4488 & ~v_4490 & v_4492 & ~v_4493;
assign v_7607 = v_4495 & ~v_4501 & ~v_4503;
assign v_7608 = v_5746 & v_4628 & ~v_4629 & ~v_4631 & ~v_4633;
assign v_7609 = ~v_4635 & ~v_4637;
assign v_7610 = v_5759 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7611 = v_4644 & v_4645;
assign v_7612 = v_5765 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7613 = v_4644 & ~v_4645 & v_4659;
assign v_7614 = v_5780 & v_4693 & ~v_4694 & ~v_4696 & ~v_4698;
assign v_7615 = ~v_4700 & ~v_4702;
assign v_7616 = v_5793 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7617 = v_4709 & v_4710;
assign v_7618 = v_5799 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7619 = v_4709 & ~v_4710 & v_4724;
assign v_7620 = v_5810 & v_4752 & ~v_4754 & v_4756 & ~v_4757;
assign v_7621 = v_4759 & ~v_4765 & ~v_4767 & v_4778;
assign v_7622 = v_5873 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7623 = ~v_4931;
assign v_7624 = v_5873 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7625 = v_4931;
assign v_7626 = v_5898 & v_4961 & v_4978 & v_4979 & v_4980;
assign v_7627 = v_4982;
assign v_7628 = v_5926 & v_4488 & ~v_4490 & v_4492 & ~v_4493;
assign v_7629 = v_4495 & ~v_4501 & ~v_4503 & v_4514;
assign v_7630 = v_5967 & v_4628 & ~v_4629 & ~v_4631 & ~v_4633;
assign v_7631 = ~v_4635 & ~v_4637;
assign v_7632 = v_5980 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7633 = v_4644 & v_4645;
assign v_7634 = v_5986 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7635 = v_4644 & ~v_4645 & v_4659;
assign v_7636 = v_6001 & v_4693 & ~v_4694 & ~v_4696 & ~v_4698;
assign v_7637 = ~v_4700 & ~v_4702;
assign v_7638 = v_6014 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7639 = v_4709 & v_4710;
assign v_7640 = v_6020 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7641 = v_4709 & ~v_4710 & v_4724;
assign v_7642 = v_6031 & v_4752 & ~v_4754 & v_4756 & ~v_4757;
assign v_7643 = v_4759 & ~v_4765 & ~v_4767 & v_4778;
assign v_7644 = v_6094 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7645 = ~v_4931;
assign v_7646 = v_6094 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7647 = v_4931;
assign v_7648 = v_6119 & v_4961 & v_4978 & v_4979 & v_4980;
assign v_7649 = v_4982;
assign v_7650 = v_6147 & v_4488 & ~v_4490 & v_4492 & ~v_4493;
assign v_7651 = v_4495 & ~v_4501 & ~v_4503 & v_4514;
assign v_7652 = v_6188 & v_4628 & ~v_4629 & ~v_4631 & ~v_4633;
assign v_7653 = ~v_4635 & ~v_4637;
assign v_7654 = v_6201 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7655 = v_4644 & v_4645;
assign v_7656 = v_6207 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7657 = v_4644 & ~v_4645 & v_4659;
assign v_7658 = v_6222 & v_4693 & ~v_4694 & ~v_4696 & ~v_4698;
assign v_7659 = ~v_4700 & ~v_4702;
assign v_7660 = v_6235 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7661 = v_4709 & v_4710;
assign v_7662 = v_6241 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7663 = v_4709 & ~v_4710 & v_4724;
assign v_7664 = v_6252 & v_4752 & ~v_4754 & v_4756 & ~v_4757;
assign v_7665 = v_4759 & ~v_4765 & ~v_4767 & v_4778;
assign v_7666 = v_6315 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7667 = ~v_4931;
assign v_7668 = v_6315 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7669 = v_4931;
assign v_7670 = v_6340 & v_4961 & v_4978 & v_4979 & v_4980;
assign v_7671 = v_4982;
assign v_7672 = v_6367 & v_4488 & ~v_4490 & v_4492 & ~v_4493;
assign v_7673 = v_4495 & ~v_4501 & ~v_4503 & v_4514;
assign v_7674 = v_6408 & v_4628 & ~v_4629 & ~v_4631 & ~v_4633;
assign v_7675 = ~v_4635 & ~v_4637;
assign v_7676 = v_6421 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7677 = v_4644 & v_4645;
assign v_7678 = v_6427 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7679 = v_4644 & ~v_4645 & v_4659;
assign v_7680 = v_6442 & v_4693 & ~v_4694 & ~v_4696 & ~v_4698;
assign v_7681 = ~v_4700 & ~v_4702;
assign v_7682 = v_6455 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7683 = v_4709 & v_4710;
assign v_7684 = v_6461 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7685 = v_4709 & ~v_4710 & v_4724;
assign v_7686 = v_6472 & v_4752 & ~v_4754 & v_4756 & ~v_4757;
assign v_7687 = v_4759 & ~v_4765 & ~v_4767 & v_4778;
assign v_7688 = v_6535 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7689 = ~v_4931;
assign v_7690 = v_6535 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7691 = v_4931;
assign v_7692 = v_6560 & v_4961 & v_4978 & v_4979 & v_4980;
assign v_7693 = v_4982;
assign v_7694 = v_6588 & v_4488 & ~v_4490 & v_4492 & ~v_4493;
assign v_7695 = v_4495 & ~v_4501 & ~v_4503 & v_4514;
assign v_7696 = v_6629 & v_4628 & ~v_4629 & ~v_4631 & ~v_4633;
assign v_7697 = ~v_4635 & ~v_4637;
assign v_7698 = v_6642 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7699 = v_4644 & v_4645;
assign v_7700 = v_6648 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7701 = v_4644 & ~v_4645 & v_4659;
assign v_7702 = v_6663 & v_4693 & ~v_4694 & ~v_4696 & ~v_4698;
assign v_7703 = ~v_4700 & ~v_4702;
assign v_7704 = v_6676 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7705 = v_4709 & v_4710;
assign v_7706 = v_6682 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7707 = v_4709 & ~v_4710 & v_4724;
assign v_7708 = v_6693 & v_4752 & ~v_4754 & v_4756 & ~v_4757;
assign v_7709 = v_4759 & ~v_4765 & ~v_4767 & v_4778;
assign v_7710 = v_6756 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7711 = ~v_4931;
assign v_7712 = v_6756 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7713 = v_4931;
assign v_7714 = v_6781 & v_4961 & v_4978 & v_4979 & v_4980;
assign v_7715 = v_4982;
assign v_7716 = v_6843 & v_4628 & ~v_4629 & ~v_4631 & ~v_4633;
assign v_7717 = ~v_4635 & ~v_4637;
assign v_7718 = v_6856 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7719 = v_4644 & v_4645;
assign v_7720 = v_6862 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7721 = v_4644 & ~v_4645 & v_4659;
assign v_7722 = v_6877 & v_4693 & ~v_4694 & ~v_4696 & ~v_4698;
assign v_7723 = ~v_4700 & ~v_4702;
assign v_7724 = v_6890 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7725 = v_4709 & v_4710;
assign v_7726 = v_6896 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7727 = v_4709 & ~v_4710 & v_4724;
assign v_7728 = v_6950 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7729 = ~v_4931;
assign v_7730 = v_6950 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7731 = v_4931;
assign v_7732 = v_6971 & v_4961 & v_4978 & v_4979 & v_4980;
assign v_7733 = v_4982;
assign v_7734 = v_6995 & v_4488 & ~v_4490 & v_4492 & ~v_4493;
assign v_7735 = v_4495 & ~v_4501 & ~v_4503 & v_4514;
assign v_7736 = v_7036 & v_4628 & ~v_4629 & ~v_4631 & ~v_4633;
assign v_7737 = ~v_4635 & ~v_4637;
assign v_7738 = v_7049 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7739 = v_4644 & v_4645;
assign v_7740 = v_7055 & v_4612 & ~v_4613 & v_4625 & ~v_4626;
assign v_7741 = v_4644 & ~v_4645 & v_4659;
assign v_7742 = v_7070 & v_4693 & ~v_4694 & ~v_4696 & ~v_4698;
assign v_7743 = ~v_4700 & ~v_4702;
assign v_7744 = v_7083 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7745 = v_4709 & v_4710;
assign v_7746 = v_7089 & v_4677 & ~v_4678 & v_4690 & ~v_4691;
assign v_7747 = v_4709 & ~v_4710 & v_4724;
assign v_7748 = v_7100 & v_4752 & ~v_4754 & v_4756 & ~v_4757;
assign v_7749 = v_4759 & ~v_4765 & ~v_4767 & v_4778;
assign v_7750 = v_7163 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7751 = ~v_4931;
assign v_7752 = v_7163 & v_4925 & v_4926 & v_4928 & ~v_4930;
assign v_7753 = v_4931;
assign v_7754 = v_7188 & v_4961 & v_4978 & v_4979 & v_4980;
assign v_7755 = v_4982;
assign v_7756 = ~v_7209 & ~v_7210 & ~v_7211 & ~v_7212 & ~v_7213;
assign v_7757 = ~v_7214 & ~v_7215 & ~v_7216 & ~v_7217 & ~v_7218;
assign v_7758 = v_5053;
assign v_217 = ~v_213 | v_215 | v_216;
assign v_224 = v_222 | v_223;
assign v_258 = ~v_254 | v_256 | v_257;
assign v_260 = v_7759 | v_7760 | v_7761;
assign v_267 = v_261 | v_263 | v_265 | v_266;
assign v_271 = v_228 | v_269 | v_270;
assign v_277 = v_275 | v_276;
assign v_285 = v_282 | v_284;
assign v_291 = ~v_280 | v_287 | v_289 | v_290;
assign v_300 = v_297 | v_299;
assign v_302 = ~v_279 | v_294 | v_296 | v_301;
assign v_306 = v_304 | v_305;
assign v_315 = ~v_311 | v_313 | v_314;
assign v_321 = v_317 | v_319 | v_320;
assign v_329 = v_323 | v_325 | v_327 | v_328;
assign v_331 = v_308 | v_310 | v_330;
assign v_343 = ~v_333 | v_335 | v_337 | v_341 | v_342;
assign v_356 = v_353 | v_355;
assign v_369 = v_361 | v_363 | v_365 | v_367 | v_368;
assign v_384 = v_380 | v_382 | v_383;
assign v_388 = v_374 | v_376 | v_378 | v_386 | v_387;
assign v_403 = v_7762 | v_7763;
assign v_405 = v_371 | v_390 | v_404;
assign v_409 = v_7764 | v_7765;
assign v_421 = v_418 | v_420;
assign v_434 = v_426 | v_428 | v_430 | v_432 | v_433;
assign v_449 = v_445 | v_447 | v_448;
assign v_453 = v_439 | v_441 | v_443 | v_451 | v_452;
assign v_468 = v_7766 | v_7767;
assign v_470 = v_436 | v_455 | v_469;
assign v_474 = v_7768 | v_7769;
assign v_480 = v_476 | v_478 | v_479;
assign v_484 = v_482 | v_483;
assign v_522 = ~v_518 | v_520 | v_521;
assign v_524 = v_7770 | v_7771 | v_7772;
assign v_531 = v_525 | v_527 | v_529 | v_530;
assign v_535 = v_492 | v_533 | v_534;
assign v_541 = v_539 | v_540;
assign v_546 = ~v_542 | v_544 | v_545;
assign v_554 = v_552 | v_553;
assign v_558 = v_548 | v_557;
assign v_568 = v_562 | v_566 | v_567;
assign v_577 = ~v_573 | v_575 | v_576;
assign v_581 = v_560 | v_570 | v_572 | v_579 | v_580;
assign v_588 = v_585 | v_587;
assign v_593 = v_590 | v_592;
assign v_598 = v_595 | v_583 | v_596 | v_597;
assign v_604 = ~v_600 | v_602 | v_603;
assign v_612 = v_610 | v_611;
assign v_616 = v_606 | v_615;
assign v_626 = v_620 | v_624 | v_625;
assign v_635 = ~v_631 | v_633 | v_634;
assign v_639 = v_618 | v_628 | v_630 | v_637 | v_638;
assign v_652 = v_650 | v_651;
assign v_654 = v_648 | v_653;
assign v_656 = v_646 | v_655;
assign v_658 = v_644 | v_657;
assign v_660 = v_642 | v_659;
assign v_662 = v_640 | v_661;
assign v_679 = v_677 | v_678;
assign v_689 = v_686 | v_688;
assign v_694 = v_691 | v_693;
assign v_699 = v_696 | v_684 | v_697 | v_698;
assign v_703 = v_7773 | v_7774;
assign v_710 = ~v_706 | v_708 | v_709;
assign v_718 = v_716 | v_717;
assign v_722 = v_712 | v_721;
assign v_737 = v_734 | v_736;
assign v_745 = v_740 | v_741 | v_743 | v_744;
assign v_750 = ~v_746 | v_748 | v_749;
assign v_758 = v_752 | v_757;
assign v_763 = ~v_759 | v_761 | v_762;
assign v_771 = v_765 | v_770;
assign v_779 = ~v_775 | v_777 | v_778;
assign v_787 = v_785 | v_786;
assign v_791 = v_781 | v_790;
assign v_796 = v_7775 | v_7776;
assign v_804 = v_802 | v_803;
assign v_808 = v_806 | v_807;
assign v_814 = ~v_800 | v_810 | v_812 | v_813;
assign v_821 = v_819 | v_820;
assign v_827 = v_825 | v_826;
assign v_831 = v_829 | v_830;
assign v_837 = ~v_823 | v_833 | v_835 | v_836;
assign v_844 = v_842 | v_843;
assign v_850 = v_848 | v_849;
assign v_854 = v_852 | v_853;
assign v_860 = ~v_846 | v_856 | v_858 | v_859;
assign v_867 = v_865 | v_866;
assign v_877 = v_7777 | v_7778 | v_7779;
assign v_885 = v_883 | v_884;
assign v_889 = v_887 | v_888;
assign v_895 = ~v_881 | v_891 | v_893 | v_894;
assign v_902 = v_900 | v_901;
assign v_908 = v_906 | v_907;
assign v_912 = v_910 | v_911;
assign v_918 = ~v_904 | v_914 | v_916 | v_917;
assign v_925 = v_923 | v_924;
assign v_931 = v_929 | v_930;
assign v_935 = v_933 | v_934;
assign v_941 = ~v_927 | v_937 | v_939 | v_940;
assign v_948 = v_946 | v_947;
assign v_958 = v_7780 | v_7781 | v_7782;
assign v_966 = v_964 | v_965;
assign v_970 = v_968 | v_969;
assign v_976 = ~v_962 | v_972 | v_974 | v_975;
assign v_983 = v_981 | v_982;
assign v_989 = v_987 | v_988;
assign v_993 = v_991 | v_992;
assign v_999 = ~v_985 | v_995 | v_997 | v_998;
assign v_1006 = v_1004 | v_1005;
assign v_1012 = v_1010 | v_1011;
assign v_1016 = v_1014 | v_1015;
assign v_1022 = ~v_1008 | v_1018 | v_1020 | v_1021;
assign v_1029 = v_1027 | v_1028;
assign v_1039 = v_7783 | v_7784 | v_7785;
assign v_1045 = v_1044 | ~v_1043;
assign v_1052 = v_7786 | v_7787;
assign v_1054 = v_252 | v_253;
assign v_1057 = v_1053 | v_1055 | v_1056;
assign v_1059 = v_1048 | v_1049 | v_1050 | v_1058;
assign v_1061 = v_1060 | ~v_1059;
assign v_1064 = v_1062 | v_1063;
assign v_1066 = v_294 | v_296;
assign v_1069 = v_1065 | v_1067 | v_1068;
assign v_1070 = v_308 | v_310;
assign v_1076 = v_1073 | v_1074 | v_1075;
assign v_1077 = v_325 | v_327 | v_328;
assign v_1079 = v_1072 | v_1078;
assign v_1081 = v_1071 | v_1080;
assign v_1082 = ~v_333 | v_335 | v_337;
assign v_1084 = v_341 | v_342;
assign v_1086 = v_1083 | v_1085;
assign v_1088 = v_1046 | v_1087;
assign v_1096 = v_367 | v_368;
assign v_1098 = v_1095 | v_1097;
assign v_1099 = v_365 | v_367 | v_368;
assign v_1101 = v_1093 | v_1094 | v_1100;
assign v_1106 = v_380 | v_382;
assign v_1109 = v_1107 | v_1108;
assign v_1112 = v_1110 | v_1111;
assign v_1113 = v_386 | v_387;
assign v_1115 = v_1103 | v_1104 | v_1105 | v_1114;
assign v_1120 = v_399 | v_401 | v_402;
assign v_1122 = v_1117 | v_1118 | v_1119 | v_1121;
assign v_1124 = v_1102 | v_1116 | v_1123;
assign v_1125 = v_407 | v_408;
assign v_1127 = v_1089 | v_1090 | v_1091 | v_1092 | v_1126;
assign v_1135 = v_432 | v_433;
assign v_1137 = v_1134 | v_1136;
assign v_1138 = v_430 | v_432 | v_433;
assign v_1140 = v_1132 | v_1133 | v_1139;
assign v_1145 = v_445 | v_447;
assign v_1148 = v_1146 | v_1147;
assign v_1151 = v_1149 | v_1150;
assign v_1152 = v_451 | v_452;
assign v_1154 = v_1142 | v_1143 | v_1144 | v_1153;
assign v_1159 = v_464 | v_466 | v_467;
assign v_1161 = v_1156 | v_1157 | v_1158 | v_1160;
assign v_1163 = v_1141 | v_1155 | v_1162;
assign v_1164 = v_472 | v_473;
assign v_1166 = v_1128 | v_1129 | v_1130 | v_1131 | v_1165;
assign v_1171 = v_1170 | ~v_1166;
assign v_1177 = v_1175 | v_1176;
assign v_1178 = v_7788 | v_7789;
assign v_1180 = v_516 | v_517;
assign v_1183 = v_1179 | v_1181 | v_1182;
assign v_1185 = v_1172 | v_1173 | v_1174 | v_1184;
assign v_1187 = v_1186 | ~v_1185;
assign v_1190 = v_1167 | v_1188 | v_1189;
assign v_1193 = v_1191 | v_1192;
assign v_1196 = v_566 | v_567;
assign v_1198 = v_1195 | v_1197;
assign v_1199 = v_570 | v_572;
assign v_1201 = v_579 | v_580;
assign v_1203 = v_1194 | v_1200 | v_1202;
assign v_1208 = v_1204 | v_1205 | v_1206 | v_1207;
assign v_1211 = v_1209 | v_1210;
assign v_1214 = v_624 | v_625;
assign v_1216 = v_1213 | v_1215;
assign v_1217 = v_628 | v_630;
assign v_1219 = v_637 | v_638;
assign v_1221 = v_1212 | v_1218 | v_1220;
assign v_1229 = v_1227 | v_1228;
assign v_1231 = v_1226 | v_1230;
assign v_1233 = v_1225 | v_1232;
assign v_1235 = v_1224 | v_1234;
assign v_1237 = v_1223 | v_1236;
assign v_1239 = v_1222 | v_1238;
assign v_1244 = v_1242 | v_1243;
assign v_1250 = v_1246 | v_1247 | v_1248 | v_1249;
assign v_1251 = v_701 | v_702;
assign v_1253 = v_1245 | v_1252;
assign v_1254 = v_683 | v_701 | v_702;
assign v_1257 = v_671 | v_673;
assign v_1259 = v_1240 | v_1241 | v_1255 | v_1256 | v_1258;
assign v_1263 = v_1261 | v_1262;
assign v_1265 = v_730 | v_732;
assign v_1269 = v_1267 | v_1268;
assign v_1272 = v_1270 | v_1271;
assign v_1277 = v_1275 | v_1276;
assign v_1278 = v_793 | v_794;
assign v_1280 = v_7790 | v_7791;
assign v_1285 = v_812 | v_813;
assign v_1287 = v_1283 | v_1284 | v_1286;
assign v_1289 = v_1282 | v_1288;
assign v_1294 = v_835 | v_836;
assign v_1296 = v_1292 | v_1293 | v_1295;
assign v_1298 = v_1291 | v_1297;
assign v_1302 = v_858 | v_859;
assign v_1304 = v_1300 | v_1301 | v_1303;
assign v_1308 = v_1306 | v_1307;
assign v_1309 = v_873 | v_871;
assign v_1314 = v_1310 | v_1311 | v_1312 | v_1313;
assign v_1315 = v_871 | v_873 | v_874 | v_875 | v_876;
assign v_1319 = v_7792 | v_7793;
assign v_1324 = v_893 | v_894;
assign v_1326 = v_1322 | v_1323 | v_1325;
assign v_1328 = v_1321 | v_1327;
assign v_1333 = v_916 | v_917;
assign v_1335 = v_1331 | v_1332 | v_1334;
assign v_1337 = v_1330 | v_1336;
assign v_1341 = v_939 | v_940;
assign v_1343 = v_1339 | v_1340 | v_1342;
assign v_1347 = v_1345 | v_1346;
assign v_1348 = v_954 | v_952;
assign v_1353 = v_1349 | v_1350 | v_1351 | v_1352;
assign v_1354 = v_952 | v_954 | v_955 | v_956 | v_957;
assign v_1358 = v_7794 | v_7795;
assign v_1363 = v_974 | v_975;
assign v_1365 = v_1361 | v_1362 | v_1364;
assign v_1367 = v_1360 | v_1366;
assign v_1372 = v_997 | v_998;
assign v_1374 = v_1370 | v_1371 | v_1373;
assign v_1376 = v_1369 | v_1375;
assign v_1380 = v_1020 | v_1021;
assign v_1382 = v_1378 | v_1379 | v_1381;
assign v_1386 = v_1384 | v_1385;
assign v_1387 = v_1035 | v_1033;
assign v_1392 = v_1388 | v_1389 | v_1390 | v_1391;
assign v_1393 = v_1033 | v_1035 | v_1036 | v_1037 | v_1038;
assign v_1397 = v_7796 | v_7797;
assign v_1399 = v_1398 | v_1043;
assign v_1403 = v_1402 | v_1059;
assign v_1406 = v_1401 | v_1404 | v_1405;
assign v_1408 = v_294 | v_296;
assign v_1411 = v_1407 | v_1409 | v_1410;
assign v_1412 = v_308 | v_310;
assign v_1418 = v_1415 | v_1416 | v_1417;
assign v_1420 = v_1414 | v_1419;
assign v_1422 = v_1413 | v_1421;
assign v_1423 = ~v_333 | v_335 | v_337;
assign v_1426 = v_1424 | v_1425;
assign v_1428 = v_1400 | v_1427;
assign v_1437 = v_1435 | v_1436;
assign v_1439 = v_1433 | v_1434 | v_1438;
assign v_1444 = v_380 | v_382;
assign v_1447 = v_1445 | v_1446;
assign v_1450 = v_1448 | v_1449;
assign v_1452 = v_1441 | v_1442 | v_1443 | v_1451;
assign v_1458 = v_1454 | v_1455 | v_1456 | v_1457;
assign v_1460 = v_1440 | v_1453 | v_1459;
assign v_1462 = v_1429 | v_1430 | v_1431 | v_1432 | v_1461;
assign v_1471 = v_1469 | v_1470;
assign v_1473 = v_1467 | v_1468 | v_1472;
assign v_1478 = v_445 | v_447;
assign v_1481 = v_1479 | v_1480;
assign v_1484 = v_1482 | v_1483;
assign v_1486 = v_1475 | v_1476 | v_1477 | v_1485;
assign v_1492 = v_1488 | v_1489 | v_1490 | v_1491;
assign v_1494 = v_1474 | v_1487 | v_1493;
assign v_1496 = v_1463 | v_1464 | v_1465 | v_1466 | v_1495;
assign v_1499 = v_1498 | v_1185;
assign v_1502 = v_1497 | v_1500 | v_1501;
assign v_1505 = v_1503 | v_1504;
assign v_1509 = v_1507 | v_1508;
assign v_1510 = v_570 | v_572;
assign v_1513 = v_1506 | v_1511 | v_1512;
assign v_1518 = v_1514 | v_1515 | v_1516 | v_1517;
assign v_1521 = v_1519 | v_1520;
assign v_1525 = v_1523 | v_1524;
assign v_1526 = v_628 | v_630;
assign v_1529 = v_1522 | v_1527 | v_1528;
assign v_1537 = v_1535 | v_1536;
assign v_1539 = v_1534 | v_1538;
assign v_1541 = v_1533 | v_1540;
assign v_1543 = v_1532 | v_1542;
assign v_1545 = v_1531 | v_1544;
assign v_1547 = v_1530 | v_1546;
assign v_1552 = v_1550 | v_1551;
assign v_1558 = v_1554 | v_1555 | v_1556 | v_1557;
assign v_1560 = v_1553 | v_1559;
assign v_1564 = v_1548 | v_1549 | v_1561 | v_1562 | v_1563;
assign v_1568 = v_1566 | v_1567;
assign v_1570 = v_730 | v_732;
assign v_1574 = v_1572 | v_1573;
assign v_1577 = v_1575 | v_1576;
assign v_1582 = v_1580 | v_1581;
assign v_1584 = v_7798 | v_7799;
assign v_1590 = v_1587 | v_1588 | v_1589;
assign v_1592 = v_1586 | v_1591;
assign v_1598 = v_1595 | v_1596 | v_1597;
assign v_1600 = v_1594 | v_1599;
assign v_1605 = v_1602 | v_1603 | v_1604;
assign v_1609 = v_1607 | v_1608;
assign v_1610 = v_873 | v_871;
assign v_1615 = v_1611 | v_1612 | v_1613 | v_1614;
assign v_1619 = v_7800 | v_7801;
assign v_1625 = v_1622 | v_1623 | v_1624;
assign v_1627 = v_1621 | v_1626;
assign v_1633 = v_1630 | v_1631 | v_1632;
assign v_1635 = v_1629 | v_1634;
assign v_1640 = v_1637 | v_1638 | v_1639;
assign v_1644 = v_1642 | v_1643;
assign v_1645 = v_954 | v_952;
assign v_1650 = v_1646 | v_1647 | v_1648 | v_1649;
assign v_1654 = v_7802 | v_7803;
assign v_1660 = v_1657 | v_1658 | v_1659;
assign v_1662 = v_1656 | v_1661;
assign v_1668 = v_1665 | v_1666 | v_1667;
assign v_1670 = v_1664 | v_1669;
assign v_1675 = v_1672 | v_1673 | v_1674;
assign v_1679 = v_1677 | v_1678;
assign v_1680 = v_1035 | v_1033;
assign v_1685 = v_1681 | v_1682 | v_1683 | v_1684;
assign v_1689 = v_7804 | v_7805;
assign v_1696 = v_1694 | v_1695;
assign v_1697 = v_7806 | v_7807;
assign v_1701 = v_1698 | v_1699 | v_1700;
assign v_1703 = v_1691 | v_1692 | v_1693 | v_1702;
assign v_1706 = v_1690 | v_1704 | v_1705;
assign v_1708 = v_294 | v_296;
assign v_1711 = v_1707 | v_1709 | v_1710;
assign v_1712 = v_308 | v_310;
assign v_1718 = v_1715 | v_1716 | v_1717;
assign v_1720 = v_1714 | v_1719;
assign v_1722 = v_1713 | v_1721;
assign v_1723 = ~v_333 | v_335 | v_337;
assign v_1726 = v_1724 | v_1725;
assign v_1735 = v_1733 | v_1734;
assign v_1737 = v_1731 | v_1732 | v_1736;
assign v_1742 = v_380 | v_382;
assign v_1745 = v_1743 | v_1744;
assign v_1748 = v_1746 | v_1747;
assign v_1750 = v_1739 | v_1740 | v_1741 | v_1749;
assign v_1756 = v_1752 | v_1753 | v_1754 | v_1755;
assign v_1758 = v_1738 | v_1751 | v_1757;
assign v_1760 = v_1727 | v_1728 | v_1729 | v_1730 | v_1759;
assign v_1769 = v_1767 | v_1768;
assign v_1771 = v_1765 | v_1766 | v_1770;
assign v_1776 = v_445 | v_447;
assign v_1779 = v_1777 | v_1778;
assign v_1782 = v_1780 | v_1781;
assign v_1784 = v_1773 | v_1774 | v_1775 | v_1783;
assign v_1790 = v_1786 | v_1787 | v_1788 | v_1789;
assign v_1792 = v_1772 | v_1785 | v_1791;
assign v_1794 = v_1761 | v_1762 | v_1763 | v_1764 | v_1793;
assign v_1801 = v_1799 | v_1800;
assign v_1802 = v_7808 | v_7809;
assign v_1806 = v_1803 | v_1804 | v_1805;
assign v_1808 = v_1796 | v_1797 | v_1798 | v_1807;
assign v_1811 = v_1795 | v_1809 | v_1810;
assign v_1816 = v_1813 | v_1815;
assign v_1818 = v_1812 | v_1817;
assign v_1822 = v_1820 | v_1821;
assign v_1823 = v_570 | v_572;
assign v_1826 = v_1819 | v_1824 | v_1825;
assign v_1831 = v_1827 | v_1828 | v_1829 | v_1830;
assign v_1836 = v_1833 | v_1835;
assign v_1838 = v_1832 | v_1837;
assign v_1842 = v_1840 | v_1841;
assign v_1843 = v_628 | v_630;
assign v_1846 = v_1839 | v_1844 | v_1845;
assign v_1854 = v_1852 | v_1853;
assign v_1856 = v_1851 | v_1855;
assign v_1858 = v_1850 | v_1857;
assign v_1860 = v_1849 | v_1859;
assign v_1862 = v_1848 | v_1861;
assign v_1864 = v_1847 | v_1863;
assign v_1869 = v_1867 | v_1868;
assign v_1875 = v_1871 | v_1872 | v_1873 | v_1874;
assign v_1877 = v_1870 | v_1876;
assign v_1881 = v_1865 | v_1866 | v_1878 | v_1879 | v_1880;
assign v_1887 = v_1884 | v_1886;
assign v_1889 = v_1883 | v_1888;
assign v_1891 = v_730 | v_732;
assign v_1895 = v_1893 | v_1894;
assign v_1898 = v_1896 | v_1897;
assign v_1905 = v_1902 | v_1904;
assign v_1907 = v_1901 | v_1906;
assign v_1909 = v_7810 | v_7811;
assign v_1915 = v_1912 | v_1913 | v_1914;
assign v_1917 = v_1911 | v_1916;
assign v_1923 = v_1920 | v_1921 | v_1922;
assign v_1925 = v_1919 | v_1924;
assign v_1930 = v_1927 | v_1928 | v_1929;
assign v_1934 = v_1932 | v_1933;
assign v_1935 = v_873 | v_871;
assign v_1940 = v_1936 | v_1937 | v_1938 | v_1939;
assign v_1944 = v_7812 | v_7813;
assign v_1950 = v_1947 | v_1948 | v_1949;
assign v_1952 = v_1946 | v_1951;
assign v_1958 = v_1955 | v_1956 | v_1957;
assign v_1960 = v_1954 | v_1959;
assign v_1965 = v_1962 | v_1963 | v_1964;
assign v_1969 = v_1967 | v_1968;
assign v_1970 = v_954 | v_952;
assign v_1975 = v_1971 | v_1972 | v_1973 | v_1974;
assign v_1979 = v_7814 | v_7815;
assign v_1985 = v_1982 | v_1983 | v_1984;
assign v_1987 = v_1981 | v_1986;
assign v_1993 = v_1990 | v_1991 | v_1992;
assign v_1995 = v_1989 | v_1994;
assign v_2000 = v_1997 | v_1998 | v_1999;
assign v_2004 = v_2002 | v_2003;
assign v_2005 = v_1035 | v_1033;
assign v_2010 = v_2006 | v_2007 | v_2008 | v_2009;
assign v_2014 = v_7816 | v_7817;
assign v_2020 = v_7818 | v_7819;
assign v_2024 = v_2021 | v_2022 | v_2023;
assign v_2026 = v_2016 | v_2017 | v_2018 | v_2025;
assign v_2029 = v_2015 | v_2027 | v_2028;
assign v_2031 = v_294 | v_296;
assign v_2034 = v_2030 | v_2032 | v_2033;
assign v_2035 = v_308 | v_310;
assign v_2041 = v_2038 | v_2039 | v_2040;
assign v_2043 = v_2037 | v_2042;
assign v_2045 = v_2036 | v_2044;
assign v_2046 = ~v_333 | v_335 | v_337;
assign v_2049 = v_2047 | v_2048;
assign v_2058 = v_2056 | v_2057;
assign v_2060 = v_2054 | v_2055 | v_2059;
assign v_2065 = v_380 | v_382;
assign v_2068 = v_2066 | v_2067;
assign v_2071 = v_2069 | v_2070;
assign v_2073 = v_2062 | v_2063 | v_2064 | v_2072;
assign v_2079 = v_2075 | v_2076 | v_2077 | v_2078;
assign v_2081 = v_2061 | v_2074 | v_2080;
assign v_2083 = v_2050 | v_2051 | v_2052 | v_2053 | v_2082;
assign v_2092 = v_2090 | v_2091;
assign v_2094 = v_2088 | v_2089 | v_2093;
assign v_2099 = v_445 | v_447;
assign v_2102 = v_2100 | v_2101;
assign v_2105 = v_2103 | v_2104;
assign v_2107 = v_2096 | v_2097 | v_2098 | v_2106;
assign v_2113 = v_2109 | v_2110 | v_2111 | v_2112;
assign v_2115 = v_2095 | v_2108 | v_2114;
assign v_2117 = v_2084 | v_2085 | v_2086 | v_2087 | v_2116;
assign v_2124 = v_2122 | v_2123;
assign v_2125 = v_7820 | v_7821;
assign v_2129 = v_2126 | v_2127 | v_2128;
assign v_2131 = v_2119 | v_2120 | v_2121 | v_2130;
assign v_2134 = v_2118 | v_2132 | v_2133;
assign v_2139 = v_2136 | v_2138;
assign v_2141 = v_2135 | v_2140;
assign v_2145 = v_2143 | v_2144;
assign v_2146 = v_570 | v_572;
assign v_2149 = v_2142 | v_2147 | v_2148;
assign v_2154 = v_2150 | v_2151 | v_2152 | v_2153;
assign v_2159 = v_2156 | v_2158;
assign v_2161 = v_2155 | v_2160;
assign v_2165 = v_2163 | v_2164;
assign v_2166 = v_628 | v_630;
assign v_2169 = v_2162 | v_2167 | v_2168;
assign v_2177 = v_2175 | v_2176;
assign v_2179 = v_2174 | v_2178;
assign v_2181 = v_2173 | v_2180;
assign v_2183 = v_2172 | v_2182;
assign v_2185 = v_2171 | v_2184;
assign v_2187 = v_2170 | v_2186;
assign v_2192 = v_2190 | v_2191;
assign v_2198 = v_2194 | v_2195 | v_2196 | v_2197;
assign v_2200 = v_2193 | v_2199;
assign v_2204 = v_2188 | v_2189 | v_2201 | v_2202 | v_2203;
assign v_2210 = v_2207 | v_2209;
assign v_2212 = v_2206 | v_2211;
assign v_2214 = v_730 | v_732;
assign v_2218 = v_2216 | v_2217;
assign v_2221 = v_2219 | v_2220;
assign v_2228 = v_2225 | v_2227;
assign v_2230 = v_2224 | v_2229;
assign v_2232 = v_7822 | v_7823;
assign v_2238 = v_2235 | v_2236 | v_2237;
assign v_2240 = v_2234 | v_2239;
assign v_2246 = v_2243 | v_2244 | v_2245;
assign v_2248 = v_2242 | v_2247;
assign v_2253 = v_2250 | v_2251 | v_2252;
assign v_2257 = v_2255 | v_2256;
assign v_2258 = v_873 | v_871;
assign v_2263 = v_2259 | v_2260 | v_2261 | v_2262;
assign v_2267 = v_7824 | v_7825;
assign v_2273 = v_2270 | v_2271 | v_2272;
assign v_2275 = v_2269 | v_2274;
assign v_2281 = v_2278 | v_2279 | v_2280;
assign v_2283 = v_2277 | v_2282;
assign v_2288 = v_2285 | v_2286 | v_2287;
assign v_2292 = v_2290 | v_2291;
assign v_2293 = v_954 | v_952;
assign v_2298 = v_2294 | v_2295 | v_2296 | v_2297;
assign v_2302 = v_7826 | v_7827;
assign v_2308 = v_2305 | v_2306 | v_2307;
assign v_2310 = v_2304 | v_2309;
assign v_2316 = v_2313 | v_2314 | v_2315;
assign v_2318 = v_2312 | v_2317;
assign v_2323 = v_2320 | v_2321 | v_2322;
assign v_2327 = v_2325 | v_2326;
assign v_2328 = v_1035 | v_1033;
assign v_2333 = v_2329 | v_2330 | v_2331 | v_2332;
assign v_2337 = v_7828 | v_7829;
assign v_2345 = v_2343 | v_2344;
assign v_2346 = v_7830 | v_7831;
assign v_2350 = v_2347 | v_2348 | v_2349;
assign v_2352 = v_2340 | v_2341 | v_2342 | v_2351;
assign v_2355 = v_2339 | v_2353 | v_2354;
assign v_2357 = v_294 | v_296;
assign v_2360 = v_2356 | v_2358 | v_2359;
assign v_2361 = v_308 | v_310;
assign v_2367 = v_2364 | v_2365 | v_2366;
assign v_2369 = v_2363 | v_2368;
assign v_2371 = v_2362 | v_2370;
assign v_2372 = ~v_333 | v_335 | v_337;
assign v_2375 = v_2373 | v_2374;
assign v_2384 = v_2382 | v_2383;
assign v_2386 = v_2380 | v_2381 | v_2385;
assign v_2391 = v_380 | v_382;
assign v_2394 = v_2392 | v_2393;
assign v_2397 = v_2395 | v_2396;
assign v_2399 = v_2388 | v_2389 | v_2390 | v_2398;
assign v_2405 = v_2401 | v_2402 | v_2403 | v_2404;
assign v_2407 = v_2387 | v_2400 | v_2406;
assign v_2409 = v_2376 | v_2377 | v_2378 | v_2379 | v_2408;
assign v_2418 = v_2416 | v_2417;
assign v_2420 = v_2414 | v_2415 | v_2419;
assign v_2425 = v_445 | v_447;
assign v_2428 = v_2426 | v_2427;
assign v_2431 = v_2429 | v_2430;
assign v_2433 = v_2422 | v_2423 | v_2424 | v_2432;
assign v_2439 = v_2435 | v_2436 | v_2437 | v_2438;
assign v_2441 = v_2421 | v_2434 | v_2440;
assign v_2443 = v_2410 | v_2411 | v_2412 | v_2413 | v_2442;
assign v_2450 = v_2448 | v_2449;
assign v_2451 = v_7832 | v_7833;
assign v_2455 = v_2452 | v_2453 | v_2454;
assign v_2457 = v_2445 | v_2446 | v_2447 | v_2456;
assign v_2460 = v_2444 | v_2458 | v_2459;
assign v_2465 = v_2462 | v_2464;
assign v_2467 = v_2461 | v_2466;
assign v_2471 = v_2469 | v_2470;
assign v_2472 = v_570 | v_572;
assign v_2475 = v_2468 | v_2473 | v_2474;
assign v_2480 = v_2476 | v_2477 | v_2478 | v_2479;
assign v_2485 = v_2482 | v_2484;
assign v_2487 = v_2481 | v_2486;
assign v_2491 = v_2489 | v_2490;
assign v_2492 = v_628 | v_630;
assign v_2495 = v_2488 | v_2493 | v_2494;
assign v_2503 = v_2501 | v_2502;
assign v_2505 = v_2500 | v_2504;
assign v_2507 = v_2499 | v_2506;
assign v_2509 = v_2498 | v_2508;
assign v_2511 = v_2497 | v_2510;
assign v_2513 = v_2496 | v_2512;
assign v_2518 = v_2516 | v_2517;
assign v_2524 = v_2520 | v_2521 | v_2522 | v_2523;
assign v_2526 = v_2519 | v_2525;
assign v_2530 = v_2514 | v_2515 | v_2527 | v_2528 | v_2529;
assign v_2536 = v_2533 | v_2535;
assign v_2538 = v_2532 | v_2537;
assign v_2540 = v_730 | v_732;
assign v_2544 = v_2542 | v_2543;
assign v_2547 = v_2545 | v_2546;
assign v_2554 = v_2551 | v_2553;
assign v_2556 = v_2550 | v_2555;
assign v_2558 = v_7834 | v_7835;
assign v_2564 = v_2561 | v_2562 | v_2563;
assign v_2566 = v_2560 | v_2565;
assign v_2572 = v_2569 | v_2570 | v_2571;
assign v_2574 = v_2568 | v_2573;
assign v_2579 = v_2576 | v_2577 | v_2578;
assign v_2583 = v_2581 | v_2582;
assign v_2584 = v_873 | v_871;
assign v_2589 = v_2585 | v_2586 | v_2587 | v_2588;
assign v_2593 = v_7836 | v_7837;
assign v_2599 = v_2596 | v_2597 | v_2598;
assign v_2601 = v_2595 | v_2600;
assign v_2607 = v_2604 | v_2605 | v_2606;
assign v_2609 = v_2603 | v_2608;
assign v_2614 = v_2611 | v_2612 | v_2613;
assign v_2618 = v_2616 | v_2617;
assign v_2619 = v_954 | v_952;
assign v_2624 = v_2620 | v_2621 | v_2622 | v_2623;
assign v_2628 = v_7838 | v_7839;
assign v_2634 = v_2631 | v_2632 | v_2633;
assign v_2636 = v_2630 | v_2635;
assign v_2642 = v_2639 | v_2640 | v_2641;
assign v_2644 = v_2638 | v_2643;
assign v_2649 = v_2646 | v_2647 | v_2648;
assign v_2653 = v_2651 | v_2652;
assign v_2654 = v_1035 | v_1033;
assign v_2659 = v_2655 | v_2656 | v_2657 | v_2658;
assign v_2663 = v_7840 | v_7841;
assign v_2671 = v_2669 | v_2670;
assign v_2672 = v_7842 | v_7843;
assign v_2676 = v_2673 | v_2674 | v_2675;
assign v_2678 = v_2666 | v_2667 | v_2668 | v_2677;
assign v_2681 = v_2665 | v_2679 | v_2680;
assign v_2683 = v_294 | v_296;
assign v_2686 = v_2682 | v_2684 | v_2685;
assign v_2687 = v_308 | v_310;
assign v_2693 = v_2690 | v_2691 | v_2692;
assign v_2695 = v_2689 | v_2694;
assign v_2697 = v_2688 | v_2696;
assign v_2698 = ~v_333 | v_335 | v_337;
assign v_2701 = v_2699 | v_2700;
assign v_2710 = v_2708 | v_2709;
assign v_2712 = v_2706 | v_2707 | v_2711;
assign v_2717 = v_380 | v_382;
assign v_2720 = v_2718 | v_2719;
assign v_2723 = v_2721 | v_2722;
assign v_2725 = v_2714 | v_2715 | v_2716 | v_2724;
assign v_2731 = v_2727 | v_2728 | v_2729 | v_2730;
assign v_2733 = v_2713 | v_2726 | v_2732;
assign v_2735 = v_2702 | v_2703 | v_2704 | v_2705 | v_2734;
assign v_2744 = v_2742 | v_2743;
assign v_2746 = v_2740 | v_2741 | v_2745;
assign v_2751 = v_445 | v_447;
assign v_2754 = v_2752 | v_2753;
assign v_2757 = v_2755 | v_2756;
assign v_2759 = v_2748 | v_2749 | v_2750 | v_2758;
assign v_2765 = v_2761 | v_2762 | v_2763 | v_2764;
assign v_2767 = v_2747 | v_2760 | v_2766;
assign v_2769 = v_2736 | v_2737 | v_2738 | v_2739 | v_2768;
assign v_2776 = v_2774 | v_2775;
assign v_2777 = v_7844 | v_7845;
assign v_2781 = v_2778 | v_2779 | v_2780;
assign v_2783 = v_2771 | v_2772 | v_2773 | v_2782;
assign v_2786 = v_2770 | v_2784 | v_2785;
assign v_2791 = v_2788 | v_2790;
assign v_2793 = v_2787 | v_2792;
assign v_2797 = v_2795 | v_2796;
assign v_2798 = v_570 | v_572;
assign v_2801 = v_2794 | v_2799 | v_2800;
assign v_2806 = v_2802 | v_2803 | v_2804 | v_2805;
assign v_2811 = v_2808 | v_2810;
assign v_2813 = v_2807 | v_2812;
assign v_2817 = v_2815 | v_2816;
assign v_2818 = v_628 | v_630;
assign v_2821 = v_2814 | v_2819 | v_2820;
assign v_2829 = v_2827 | v_2828;
assign v_2831 = v_2826 | v_2830;
assign v_2833 = v_2825 | v_2832;
assign v_2835 = v_2824 | v_2834;
assign v_2837 = v_2823 | v_2836;
assign v_2839 = v_2822 | v_2838;
assign v_2844 = v_2842 | v_2843;
assign v_2850 = v_2846 | v_2847 | v_2848 | v_2849;
assign v_2852 = v_2845 | v_2851;
assign v_2856 = v_2840 | v_2841 | v_2853 | v_2854 | v_2855;
assign v_2862 = v_2859 | v_2861;
assign v_2864 = v_2858 | v_2863;
assign v_2866 = v_730 | v_732;
assign v_2870 = v_2868 | v_2869;
assign v_2873 = v_2871 | v_2872;
assign v_2880 = v_2877 | v_2879;
assign v_2882 = v_2876 | v_2881;
assign v_2884 = v_7846 | v_7847;
assign v_2890 = v_2887 | v_2888 | v_2889;
assign v_2892 = v_2886 | v_2891;
assign v_2898 = v_2895 | v_2896 | v_2897;
assign v_2900 = v_2894 | v_2899;
assign v_2905 = v_2902 | v_2903 | v_2904;
assign v_2909 = v_2907 | v_2908;
assign v_2910 = v_873 | v_871;
assign v_2915 = v_2911 | v_2912 | v_2913 | v_2914;
assign v_2919 = v_7848 | v_7849;
assign v_2925 = v_2922 | v_2923 | v_2924;
assign v_2927 = v_2921 | v_2926;
assign v_2933 = v_2930 | v_2931 | v_2932;
assign v_2935 = v_2929 | v_2934;
assign v_2940 = v_2937 | v_2938 | v_2939;
assign v_2944 = v_2942 | v_2943;
assign v_2945 = v_954 | v_952;
assign v_2950 = v_2946 | v_2947 | v_2948 | v_2949;
assign v_2954 = v_7850 | v_7851;
assign v_2960 = v_2957 | v_2958 | v_2959;
assign v_2962 = v_2956 | v_2961;
assign v_2968 = v_2965 | v_2966 | v_2967;
assign v_2970 = v_2964 | v_2969;
assign v_2975 = v_2972 | v_2973 | v_2974;
assign v_2979 = v_2977 | v_2978;
assign v_2980 = v_1035 | v_1033;
assign v_2985 = v_2981 | v_2982 | v_2983 | v_2984;
assign v_2989 = v_7852 | v_7853;
assign v_2996 = v_2994 | v_2995;
assign v_2997 = v_7854 | v_7855;
assign v_3001 = v_2998 | v_2999 | v_3000;
assign v_3003 = v_2991 | v_2992 | v_2993 | v_3002;
assign v_3006 = v_2990 | v_3004 | v_3005;
assign v_3008 = v_294 | v_296;
assign v_3011 = v_3007 | v_3009 | v_3010;
assign v_3012 = v_308 | v_310;
assign v_3018 = v_3015 | v_3016 | v_3017;
assign v_3020 = v_3014 | v_3019;
assign v_3022 = v_3013 | v_3021;
assign v_3023 = ~v_333 | v_335 | v_337;
assign v_3026 = v_3024 | v_3025;
assign v_3035 = v_3033 | v_3034;
assign v_3037 = v_3031 | v_3032 | v_3036;
assign v_3042 = v_380 | v_382;
assign v_3045 = v_3043 | v_3044;
assign v_3048 = v_3046 | v_3047;
assign v_3050 = v_3039 | v_3040 | v_3041 | v_3049;
assign v_3056 = v_3052 | v_3053 | v_3054 | v_3055;
assign v_3058 = v_3038 | v_3051 | v_3057;
assign v_3060 = v_3027 | v_3028 | v_3029 | v_3030 | v_3059;
assign v_3069 = v_3067 | v_3068;
assign v_3071 = v_3065 | v_3066 | v_3070;
assign v_3076 = v_445 | v_447;
assign v_3079 = v_3077 | v_3078;
assign v_3082 = v_3080 | v_3081;
assign v_3084 = v_3073 | v_3074 | v_3075 | v_3083;
assign v_3090 = v_3086 | v_3087 | v_3088 | v_3089;
assign v_3092 = v_3072 | v_3085 | v_3091;
assign v_3094 = v_3061 | v_3062 | v_3063 | v_3064 | v_3093;
assign v_3101 = v_3099 | v_3100;
assign v_3102 = v_7856 | v_7857;
assign v_3106 = v_3103 | v_3104 | v_3105;
assign v_3108 = v_3096 | v_3097 | v_3098 | v_3107;
assign v_3111 = v_3095 | v_3109 | v_3110;
assign v_3116 = v_3113 | v_3115;
assign v_3118 = v_3112 | v_3117;
assign v_3122 = v_3120 | v_3121;
assign v_3123 = v_570 | v_572;
assign v_3126 = v_3119 | v_3124 | v_3125;
assign v_3131 = v_3127 | v_3128 | v_3129 | v_3130;
assign v_3136 = v_3133 | v_3135;
assign v_3138 = v_3132 | v_3137;
assign v_3142 = v_3140 | v_3141;
assign v_3143 = v_628 | v_630;
assign v_3146 = v_3139 | v_3144 | v_3145;
assign v_3154 = v_3152 | v_3153;
assign v_3156 = v_3151 | v_3155;
assign v_3158 = v_3150 | v_3157;
assign v_3160 = v_3149 | v_3159;
assign v_3162 = v_3148 | v_3161;
assign v_3164 = v_3147 | v_3163;
assign v_3169 = v_3167 | v_3168;
assign v_3175 = v_3171 | v_3172 | v_3173 | v_3174;
assign v_3177 = v_3170 | v_3176;
assign v_3181 = v_3165 | v_3166 | v_3178 | v_3179 | v_3180;
assign v_3187 = v_3184 | v_3186;
assign v_3189 = v_3183 | v_3188;
assign v_3191 = v_730 | v_732;
assign v_3195 = v_3193 | v_3194;
assign v_3198 = v_3196 | v_3197;
assign v_3205 = v_3202 | v_3204;
assign v_3207 = v_3201 | v_3206;
assign v_3209 = v_7858 | v_7859;
assign v_3215 = v_3212 | v_3213 | v_3214;
assign v_3217 = v_3211 | v_3216;
assign v_3223 = v_3220 | v_3221 | v_3222;
assign v_3225 = v_3219 | v_3224;
assign v_3230 = v_3227 | v_3228 | v_3229;
assign v_3234 = v_3232 | v_3233;
assign v_3235 = v_873 | v_871;
assign v_3240 = v_3236 | v_3237 | v_3238 | v_3239;
assign v_3244 = v_7860 | v_7861;
assign v_3250 = v_3247 | v_3248 | v_3249;
assign v_3252 = v_3246 | v_3251;
assign v_3258 = v_3255 | v_3256 | v_3257;
assign v_3260 = v_3254 | v_3259;
assign v_3265 = v_3262 | v_3263 | v_3264;
assign v_3269 = v_3267 | v_3268;
assign v_3270 = v_954 | v_952;
assign v_3275 = v_3271 | v_3272 | v_3273 | v_3274;
assign v_3279 = v_7862 | v_7863;
assign v_3285 = v_3282 | v_3283 | v_3284;
assign v_3287 = v_3281 | v_3286;
assign v_3293 = v_3290 | v_3291 | v_3292;
assign v_3295 = v_3289 | v_3294;
assign v_3300 = v_3297 | v_3298 | v_3299;
assign v_3304 = v_3302 | v_3303;
assign v_3305 = v_1035 | v_1033;
assign v_3310 = v_3306 | v_3307 | v_3308 | v_3309;
assign v_3314 = v_7864 | v_7865;
assign v_3322 = v_3320 | v_3321;
assign v_3323 = v_7866 | v_7867;
assign v_3327 = v_3324 | v_3325 | v_3326;
assign v_3329 = v_3317 | v_3318 | v_3319 | v_3328;
assign v_3332 = v_3316 | v_3330 | v_3331;
assign v_3334 = v_294 | v_296;
assign v_3337 = v_3333 | v_3335 | v_3336;
assign v_3338 = v_308 | v_310;
assign v_3344 = v_3341 | v_3342 | v_3343;
assign v_3346 = v_3340 | v_3345;
assign v_3348 = v_3339 | v_3347;
assign v_3349 = ~v_333 | v_335 | v_337;
assign v_3352 = v_3350 | v_3351;
assign v_3361 = v_3359 | v_3360;
assign v_3363 = v_3357 | v_3358 | v_3362;
assign v_3368 = v_380 | v_382;
assign v_3371 = v_3369 | v_3370;
assign v_3374 = v_3372 | v_3373;
assign v_3376 = v_3365 | v_3366 | v_3367 | v_3375;
assign v_3382 = v_3378 | v_3379 | v_3380 | v_3381;
assign v_3384 = v_3364 | v_3377 | v_3383;
assign v_3386 = v_3353 | v_3354 | v_3355 | v_3356 | v_3385;
assign v_3395 = v_3393 | v_3394;
assign v_3397 = v_3391 | v_3392 | v_3396;
assign v_3402 = v_445 | v_447;
assign v_3405 = v_3403 | v_3404;
assign v_3408 = v_3406 | v_3407;
assign v_3410 = v_3399 | v_3400 | v_3401 | v_3409;
assign v_3416 = v_3412 | v_3413 | v_3414 | v_3415;
assign v_3418 = v_3398 | v_3411 | v_3417;
assign v_3420 = v_3387 | v_3388 | v_3389 | v_3390 | v_3419;
assign v_3427 = v_3425 | v_3426;
assign v_3428 = v_7868 | v_7869;
assign v_3432 = v_3429 | v_3430 | v_3431;
assign v_3434 = v_3422 | v_3423 | v_3424 | v_3433;
assign v_3437 = v_3421 | v_3435 | v_3436;
assign v_3442 = v_3439 | v_3441;
assign v_3444 = v_3438 | v_3443;
assign v_3448 = v_3446 | v_3447;
assign v_3449 = v_570 | v_572;
assign v_3452 = v_3445 | v_3450 | v_3451;
assign v_3457 = v_3453 | v_3454 | v_3455 | v_3456;
assign v_3462 = v_3459 | v_3461;
assign v_3464 = v_3458 | v_3463;
assign v_3468 = v_3466 | v_3467;
assign v_3469 = v_628 | v_630;
assign v_3472 = v_3465 | v_3470 | v_3471;
assign v_3480 = v_3478 | v_3479;
assign v_3482 = v_3477 | v_3481;
assign v_3484 = v_3476 | v_3483;
assign v_3486 = v_3475 | v_3485;
assign v_3488 = v_3474 | v_3487;
assign v_3490 = v_3473 | v_3489;
assign v_3495 = v_3493 | v_3494;
assign v_3501 = v_3497 | v_3498 | v_3499 | v_3500;
assign v_3503 = v_3496 | v_3502;
assign v_3507 = v_3491 | v_3492 | v_3504 | v_3505 | v_3506;
assign v_3513 = v_3510 | v_3512;
assign v_3515 = v_3509 | v_3514;
assign v_3517 = v_730 | v_732;
assign v_3521 = v_3519 | v_3520;
assign v_3524 = v_3522 | v_3523;
assign v_3531 = v_3528 | v_3530;
assign v_3533 = v_3527 | v_3532;
assign v_3535 = v_7870 | v_7871;
assign v_3541 = v_3538 | v_3539 | v_3540;
assign v_3543 = v_3537 | v_3542;
assign v_3549 = v_3546 | v_3547 | v_3548;
assign v_3551 = v_3545 | v_3550;
assign v_3556 = v_3553 | v_3554 | v_3555;
assign v_3560 = v_3558 | v_3559;
assign v_3561 = v_873 | v_871;
assign v_3566 = v_3562 | v_3563 | v_3564 | v_3565;
assign v_3570 = v_7872 | v_7873;
assign v_3576 = v_3573 | v_3574 | v_3575;
assign v_3578 = v_3572 | v_3577;
assign v_3584 = v_3581 | v_3582 | v_3583;
assign v_3586 = v_3580 | v_3585;
assign v_3591 = v_3588 | v_3589 | v_3590;
assign v_3595 = v_3593 | v_3594;
assign v_3596 = v_954 | v_952;
assign v_3601 = v_3597 | v_3598 | v_3599 | v_3600;
assign v_3605 = v_7874 | v_7875;
assign v_3611 = v_3608 | v_3609 | v_3610;
assign v_3613 = v_3607 | v_3612;
assign v_3619 = v_3616 | v_3617 | v_3618;
assign v_3621 = v_3615 | v_3620;
assign v_3626 = v_3623 | v_3624 | v_3625;
assign v_3630 = v_3628 | v_3629;
assign v_3631 = v_1035 | v_1033;
assign v_3636 = v_3632 | v_3633 | v_3634 | v_3635;
assign v_3640 = v_7876 | v_7877;
assign v_3643 = v_3642 | ~v_1086;
assign v_3649 = v_3645 | v_3647 | v_3648;
assign v_3651 = v_294 | v_296;
assign v_3654 = v_3650 | v_3652 | v_3653;
assign v_3655 = v_308 | v_310;
assign v_3661 = v_3658 | v_3659 | v_3660;
assign v_3663 = v_3657 | v_3662;
assign v_3665 = v_3656 | v_3664;
assign v_3666 = ~v_333 | v_335 | v_337;
assign v_3669 = v_3667 | v_3668;
assign v_3671 = v_3644 | v_3670;
assign v_3680 = v_3678 | v_3679;
assign v_3682 = v_3676 | v_3677 | v_3681;
assign v_3687 = v_380 | v_382;
assign v_3690 = v_3688 | v_3689;
assign v_3693 = v_3691 | v_3692;
assign v_3695 = v_3684 | v_3685 | v_3686 | v_3694;
assign v_3701 = v_3697 | v_3698 | v_3699 | v_3700;
assign v_3703 = v_3683 | v_3696 | v_3702;
assign v_3705 = v_3672 | v_3673 | v_3674 | v_3675 | v_3704;
assign v_3714 = v_3712 | v_3713;
assign v_3716 = v_3710 | v_3711 | v_3715;
assign v_3721 = v_445 | v_447;
assign v_3724 = v_3722 | v_3723;
assign v_3727 = v_3725 | v_3726;
assign v_3729 = v_3718 | v_3719 | v_3720 | v_3728;
assign v_3735 = v_3731 | v_3732 | v_3733 | v_3734;
assign v_3737 = v_3717 | v_3730 | v_3736;
assign v_3739 = v_3706 | v_3707 | v_3708 | v_3709 | v_3738;
assign v_3744 = v_3740 | v_3742 | v_3743;
assign v_3747 = v_3745 | v_3746;
assign v_3751 = v_3749 | v_3750;
assign v_3752 = v_570 | v_572;
assign v_3755 = v_3748 | v_3753 | v_3754;
assign v_3760 = v_3756 | v_3757 | v_3758 | v_3759;
assign v_3763 = v_3761 | v_3762;
assign v_3767 = v_3765 | v_3766;
assign v_3768 = v_628 | v_630;
assign v_3771 = v_3764 | v_3769 | v_3770;
assign v_3779 = v_3777 | v_3778;
assign v_3781 = v_3776 | v_3780;
assign v_3783 = v_3775 | v_3782;
assign v_3785 = v_3774 | v_3784;
assign v_3787 = v_3773 | v_3786;
assign v_3789 = v_3772 | v_3788;
assign v_3794 = v_3792 | v_3793;
assign v_3800 = v_3796 | v_3797 | v_3798 | v_3799;
assign v_3802 = v_3795 | v_3801;
assign v_3806 = v_3790 | v_3791 | v_3803 | v_3804 | v_3805;
assign v_3810 = v_3808 | v_3809;
assign v_3812 = v_730 | v_732;
assign v_3816 = v_3814 | v_3815;
assign v_3819 = v_3817 | v_3818;
assign v_3824 = v_3822 | v_3823;
assign v_3826 = v_7878 | v_7879;
assign v_3832 = v_3829 | v_3830 | v_3831;
assign v_3834 = v_3828 | v_3833;
assign v_3840 = v_3837 | v_3838 | v_3839;
assign v_3842 = v_3836 | v_3841;
assign v_3847 = v_3844 | v_3845 | v_3846;
assign v_3851 = v_3849 | v_3850;
assign v_3852 = v_873 | v_871;
assign v_3857 = v_3853 | v_3854 | v_3855 | v_3856;
assign v_3861 = v_7880 | v_7881;
assign v_3867 = v_3864 | v_3865 | v_3866;
assign v_3869 = v_3863 | v_3868;
assign v_3875 = v_3872 | v_3873 | v_3874;
assign v_3877 = v_3871 | v_3876;
assign v_3882 = v_3879 | v_3880 | v_3881;
assign v_3886 = v_3884 | v_3885;
assign v_3887 = v_954 | v_952;
assign v_3892 = v_3888 | v_3889 | v_3890 | v_3891;
assign v_3896 = v_7882 | v_7883;
assign v_3902 = v_3899 | v_3900 | v_3901;
assign v_3904 = v_3898 | v_3903;
assign v_3910 = v_3907 | v_3908 | v_3909;
assign v_3912 = v_3906 | v_3911;
assign v_3917 = v_3914 | v_3915 | v_3916;
assign v_3921 = v_3919 | v_3920;
assign v_3922 = v_1035 | v_1033;
assign v_3927 = v_3923 | v_3924 | v_3925 | v_3926;
assign v_3931 = v_7884 | v_7885;
assign v_3939 = v_3937 | v_3938;
assign v_3940 = v_7886 | v_7887;
assign v_3944 = v_3941 | v_3942 | v_3943;
assign v_3946 = v_3934 | v_3935 | v_3936 | v_3945;
assign v_3949 = v_3933 | v_3947 | v_3948;
assign v_3951 = v_294 | v_296;
assign v_3954 = v_3950 | v_3952 | v_3953;
assign v_3955 = v_308 | v_310;
assign v_3961 = v_3958 | v_3959 | v_3960;
assign v_3963 = v_3957 | v_3962;
assign v_3965 = v_3956 | v_3964;
assign v_3966 = ~v_333 | v_335 | v_337;
assign v_3969 = v_3967 | v_3968;
assign v_3978 = v_3976 | v_3977;
assign v_3980 = v_3974 | v_3975 | v_3979;
assign v_3985 = v_380 | v_382;
assign v_3988 = v_3986 | v_3987;
assign v_3991 = v_3989 | v_3990;
assign v_3993 = v_3982 | v_3983 | v_3984 | v_3992;
assign v_3999 = v_3995 | v_3996 | v_3997 | v_3998;
assign v_4001 = v_3981 | v_3994 | v_4000;
assign v_4003 = v_3970 | v_3971 | v_3972 | v_3973 | v_4002;
assign v_4012 = v_4010 | v_4011;
assign v_4014 = v_4008 | v_4009 | v_4013;
assign v_4019 = v_445 | v_447;
assign v_4022 = v_4020 | v_4021;
assign v_4025 = v_4023 | v_4024;
assign v_4027 = v_4016 | v_4017 | v_4018 | v_4026;
assign v_4033 = v_4029 | v_4030 | v_4031 | v_4032;
assign v_4035 = v_4015 | v_4028 | v_4034;
assign v_4037 = v_4004 | v_4005 | v_4006 | v_4007 | v_4036;
assign v_4044 = v_4042 | v_4043;
assign v_4045 = v_7888 | v_7889;
assign v_4049 = v_4046 | v_4047 | v_4048;
assign v_4051 = v_4039 | v_4040 | v_4041 | v_4050;
assign v_4054 = v_4038 | v_4052 | v_4053;
assign v_4059 = v_4056 | v_4058;
assign v_4061 = v_4055 | v_4060;
assign v_4065 = v_4063 | v_4064;
assign v_4066 = v_570 | v_572;
assign v_4069 = v_4062 | v_4067 | v_4068;
assign v_4074 = v_4070 | v_4071 | v_4072 | v_4073;
assign v_4079 = v_4076 | v_4078;
assign v_4081 = v_4075 | v_4080;
assign v_4085 = v_4083 | v_4084;
assign v_4086 = v_628 | v_630;
assign v_4089 = v_4082 | v_4087 | v_4088;
assign v_4097 = v_4095 | v_4096;
assign v_4099 = v_4094 | v_4098;
assign v_4101 = v_4093 | v_4100;
assign v_4103 = v_4092 | v_4102;
assign v_4105 = v_4091 | v_4104;
assign v_4107 = v_4090 | v_4106;
assign v_4112 = v_4110 | v_4111;
assign v_4118 = v_4114 | v_4115 | v_4116 | v_4117;
assign v_4120 = v_4113 | v_4119;
assign v_4124 = v_4108 | v_4109 | v_4121 | v_4122 | v_4123;
assign v_4130 = v_4127 | v_4129;
assign v_4132 = v_4126 | v_4131;
assign v_4134 = v_730 | v_732;
assign v_4138 = v_4136 | v_4137;
assign v_4141 = v_4139 | v_4140;
assign v_4148 = v_4145 | v_4147;
assign v_4150 = v_4144 | v_4149;
assign v_4152 = v_7890 | v_7891;
assign v_4158 = v_4155 | v_4156 | v_4157;
assign v_4160 = v_4154 | v_4159;
assign v_4166 = v_4163 | v_4164 | v_4165;
assign v_4168 = v_4162 | v_4167;
assign v_4173 = v_4170 | v_4171 | v_4172;
assign v_4177 = v_4175 | v_4176;
assign v_4178 = v_873 | v_871;
assign v_4183 = v_4179 | v_4180 | v_4181 | v_4182;
assign v_4187 = v_7892 | v_7893;
assign v_4193 = v_4190 | v_4191 | v_4192;
assign v_4195 = v_4189 | v_4194;
assign v_4201 = v_4198 | v_4199 | v_4200;
assign v_4203 = v_4197 | v_4202;
assign v_4208 = v_4205 | v_4206 | v_4207;
assign v_4212 = v_4210 | v_4211;
assign v_4213 = v_954 | v_952;
assign v_4218 = v_4214 | v_4215 | v_4216 | v_4217;
assign v_4222 = v_7894 | v_7895;
assign v_4228 = v_4225 | v_4226 | v_4227;
assign v_4230 = v_4224 | v_4229;
assign v_4236 = v_4233 | v_4234 | v_4235;
assign v_4238 = v_4232 | v_4237;
assign v_4243 = v_4240 | v_4241 | v_4242;
assign v_4247 = v_4245 | v_4246;
assign v_4248 = v_1035 | v_1033;
assign v_4253 = v_4249 | v_4250 | v_4251 | v_4252;
assign v_4257 = v_7896 | v_7897;
assign v_4473 = ~v_4469 | v_4471 | v_4472;
assign v_4480 = v_4478 | v_4479;
assign v_4514 = ~v_4510 | v_4512 | v_4513;
assign v_4516 = v_7898 | v_7899 | v_7900;
assign v_4523 = v_4517 | v_4519 | v_4521 | v_4522;
assign v_4527 = v_4484 | v_4525 | v_4526;
assign v_4533 = v_4531 | v_4532;
assign v_4541 = v_4538 | v_4540;
assign v_4547 = ~v_4536 | v_4543 | v_4545 | v_4546;
assign v_4556 = v_4553 | v_4555;
assign v_4558 = ~v_4535 | v_4550 | v_4552 | v_4557;
assign v_4562 = v_4560 | v_4561;
assign v_4571 = ~v_4567 | v_4569 | v_4570;
assign v_4577 = v_4573 | v_4575 | v_4576;
assign v_4585 = v_4579 | v_4581 | v_4583 | v_4584;
assign v_4587 = v_4564 | v_4566 | v_4586;
assign v_4599 = ~v_4589 | v_4591 | v_4593 | v_4597 | v_4598;
assign v_4612 = v_4609 | v_4611;
assign v_4625 = v_4617 | v_4619 | v_4621 | v_4623 | v_4624;
assign v_4640 = v_4636 | v_4638 | v_4639;
assign v_4644 = v_4630 | v_4632 | v_4634 | v_4642 | v_4643;
assign v_4659 = v_7901 | v_7902;
assign v_4661 = v_4627 | v_4646 | v_4660;
assign v_4665 = v_7903 | v_7904;
assign v_4677 = v_4674 | v_4676;
assign v_4690 = v_4682 | v_4684 | v_4686 | v_4688 | v_4689;
assign v_4705 = v_4701 | v_4703 | v_4704;
assign v_4709 = v_4695 | v_4697 | v_4699 | v_4707 | v_4708;
assign v_4724 = v_7905 | v_7906;
assign v_4726 = v_4692 | v_4711 | v_4725;
assign v_4730 = v_7907 | v_7908;
assign v_4736 = v_4732 | v_4734 | v_4735;
assign v_4740 = v_4738 | v_4739;
assign v_4778 = ~v_4774 | v_4776 | v_4777;
assign v_4780 = v_7909 | v_7910 | v_7911;
assign v_4787 = v_4781 | v_4783 | v_4785 | v_4786;
assign v_4791 = v_4748 | v_4789 | v_4790;
assign v_4797 = v_4795 | v_4796;
assign v_4802 = ~v_4798 | v_4800 | v_4801;
assign v_4810 = v_4808 | v_4809;
assign v_4814 = v_4804 | v_4813;
assign v_4824 = v_4818 | v_4822 | v_4823;
assign v_4833 = ~v_4829 | v_4831 | v_4832;
assign v_4837 = v_4816 | v_4826 | v_4828 | v_4835 | v_4836;
assign v_4844 = v_4841 | v_4843;
assign v_4849 = v_4846 | v_4848;
assign v_4854 = v_4851 | v_4839 | v_4852 | v_4853;
assign v_4860 = ~v_4856 | v_4858 | v_4859;
assign v_4868 = v_4866 | v_4867;
assign v_4872 = v_4862 | v_4871;
assign v_4882 = v_4876 | v_4880 | v_4881;
assign v_4891 = ~v_4887 | v_4889 | v_4890;
assign v_4895 = v_4874 | v_4884 | v_4886 | v_4893 | v_4894;
assign v_4908 = v_4906 | v_4907;
assign v_4910 = v_4904 | v_4909;
assign v_4912 = v_4902 | v_4911;
assign v_4914 = v_4900 | v_4913;
assign v_4916 = v_4898 | v_4915;
assign v_4918 = v_4896 | v_4917;
assign v_4935 = v_4933 | v_4934;
assign v_4945 = v_4942 | v_4944;
assign v_4950 = v_4947 | v_4949;
assign v_4955 = v_4952 | v_4940 | v_4953 | v_4954;
assign v_4959 = v_7912 | v_7913;
assign v_4966 = ~v_4962 | v_4964 | v_4965;
assign v_4974 = v_4972 | v_4973;
assign v_4978 = v_4968 | v_4977;
assign v_4993 = v_4990 | v_4992;
assign v_5001 = v_4996 | v_4997 | v_4999 | v_5000;
assign v_5006 = ~v_5002 | v_5004 | v_5005;
assign v_5014 = v_5008 | v_5013;
assign v_5019 = ~v_5015 | v_5017 | v_5018;
assign v_5027 = v_5021 | v_5026;
assign v_5035 = ~v_5031 | v_5033 | v_5034;
assign v_5043 = v_5041 | v_5042;
assign v_5047 = v_5037 | v_5046;
assign v_5052 = v_7914 | v_7915;
assign v_5058 = v_5057 | ~v_5056;
assign v_5065 = v_7916 | v_7917;
assign v_5067 = v_4508 | v_4509;
assign v_5070 = v_5066 | v_5068 | v_5069;
assign v_5072 = v_5061 | v_5062 | v_5063 | v_5071;
assign v_5074 = v_5073 | ~v_5072;
assign v_5077 = v_5075 | v_5076;
assign v_5079 = v_4550 | v_4552;
assign v_5082 = v_5078 | v_5080 | v_5081;
assign v_5083 = v_4564 | v_4566;
assign v_5089 = v_5086 | v_5087 | v_5088;
assign v_5090 = v_4581 | v_4583 | v_4584;
assign v_5092 = v_5085 | v_5091;
assign v_5094 = v_5084 | v_5093;
assign v_5095 = ~v_4589 | v_4591 | v_4593;
assign v_5097 = v_4597 | v_4598;
assign v_5099 = v_5096 | v_5098;
assign v_5101 = v_5059 | v_5100;
assign v_5109 = v_4623 | v_4624;
assign v_5111 = v_5108 | v_5110;
assign v_5112 = v_4621 | v_4623 | v_4624;
assign v_5114 = v_5106 | v_5107 | v_5113;
assign v_5119 = v_4636 | v_4638;
assign v_5122 = v_5120 | v_5121;
assign v_5125 = v_5123 | v_5124;
assign v_5126 = v_4642 | v_4643;
assign v_5128 = v_5116 | v_5117 | v_5118 | v_5127;
assign v_5133 = v_4655 | v_4657 | v_4658;
assign v_5135 = v_5130 | v_5131 | v_5132 | v_5134;
assign v_5137 = v_5115 | v_5129 | v_5136;
assign v_5138 = v_4663 | v_4664;
assign v_5140 = v_5102 | v_5103 | v_5104 | v_5105 | v_5139;
assign v_5148 = v_4688 | v_4689;
assign v_5150 = v_5147 | v_5149;
assign v_5151 = v_4686 | v_4688 | v_4689;
assign v_5153 = v_5145 | v_5146 | v_5152;
assign v_5158 = v_4701 | v_4703;
assign v_5161 = v_5159 | v_5160;
assign v_5164 = v_5162 | v_5163;
assign v_5165 = v_4707 | v_4708;
assign v_5167 = v_5155 | v_5156 | v_5157 | v_5166;
assign v_5172 = v_4720 | v_4722 | v_4723;
assign v_5174 = v_5169 | v_5170 | v_5171 | v_5173;
assign v_5176 = v_5154 | v_5168 | v_5175;
assign v_5177 = v_4728 | v_4729;
assign v_5179 = v_5141 | v_5142 | v_5143 | v_5144 | v_5178;
assign v_5184 = v_5183 | ~v_5179;
assign v_5190 = v_5188 | v_5189;
assign v_5191 = v_7918 | v_7919;
assign v_5193 = v_4772 | v_4773;
assign v_5196 = v_5192 | v_5194 | v_5195;
assign v_5198 = v_5185 | v_5186 | v_5187 | v_5197;
assign v_5200 = v_5199 | ~v_5198;
assign v_5203 = v_5180 | v_5201 | v_5202;
assign v_5206 = v_5204 | v_5205;
assign v_5209 = v_4822 | v_4823;
assign v_5211 = v_5208 | v_5210;
assign v_5212 = v_4826 | v_4828;
assign v_5214 = v_4835 | v_4836;
assign v_5216 = v_5207 | v_5213 | v_5215;
assign v_5221 = v_5217 | v_5218 | v_5219 | v_5220;
assign v_5224 = v_5222 | v_5223;
assign v_5227 = v_4880 | v_4881;
assign v_5229 = v_5226 | v_5228;
assign v_5230 = v_4884 | v_4886;
assign v_5232 = v_4893 | v_4894;
assign v_5234 = v_5225 | v_5231 | v_5233;
assign v_5242 = v_5240 | v_5241;
assign v_5244 = v_5239 | v_5243;
assign v_5246 = v_5238 | v_5245;
assign v_5248 = v_5237 | v_5247;
assign v_5250 = v_5236 | v_5249;
assign v_5252 = v_5235 | v_5251;
assign v_5257 = v_5255 | v_5256;
assign v_5263 = v_5259 | v_5260 | v_5261 | v_5262;
assign v_5264 = v_4957 | v_4958;
assign v_5266 = v_5258 | v_5265;
assign v_5267 = v_4939 | v_4957 | v_4958;
assign v_5270 = v_4927 | v_4929;
assign v_5272 = v_5253 | v_5254 | v_5268 | v_5269 | v_5271;
assign v_5276 = v_5274 | v_5275;
assign v_5278 = v_4986 | v_4988;
assign v_5282 = v_5280 | v_5281;
assign v_5285 = v_5283 | v_5284;
assign v_5290 = v_5288 | v_5289;
assign v_5291 = v_5049 | v_5050;
assign v_5293 = v_7920 | v_7921;
assign v_5295 = v_5294 | v_5056;
assign v_5299 = v_5298 | v_5072;
assign v_5302 = v_5297 | v_5300 | v_5301;
assign v_5304 = v_4550 | v_4552;
assign v_5307 = v_5303 | v_5305 | v_5306;
assign v_5308 = v_4564 | v_4566;
assign v_5314 = v_5311 | v_5312 | v_5313;
assign v_5316 = v_5310 | v_5315;
assign v_5318 = v_5309 | v_5317;
assign v_5319 = ~v_4589 | v_4591 | v_4593;
assign v_5322 = v_5320 | v_5321;
assign v_5324 = v_5296 | v_5323;
assign v_5333 = v_5331 | v_5332;
assign v_5335 = v_5329 | v_5330 | v_5334;
assign v_5340 = v_4636 | v_4638;
assign v_5343 = v_5341 | v_5342;
assign v_5346 = v_5344 | v_5345;
assign v_5348 = v_5337 | v_5338 | v_5339 | v_5347;
assign v_5354 = v_5350 | v_5351 | v_5352 | v_5353;
assign v_5356 = v_5336 | v_5349 | v_5355;
assign v_5358 = v_5325 | v_5326 | v_5327 | v_5328 | v_5357;
assign v_5367 = v_5365 | v_5366;
assign v_5369 = v_5363 | v_5364 | v_5368;
assign v_5374 = v_4701 | v_4703;
assign v_5377 = v_5375 | v_5376;
assign v_5380 = v_5378 | v_5379;
assign v_5382 = v_5371 | v_5372 | v_5373 | v_5381;
assign v_5388 = v_5384 | v_5385 | v_5386 | v_5387;
assign v_5390 = v_5370 | v_5383 | v_5389;
assign v_5392 = v_5359 | v_5360 | v_5361 | v_5362 | v_5391;
assign v_5395 = v_5394 | v_5198;
assign v_5398 = v_5393 | v_5396 | v_5397;
assign v_5401 = v_5399 | v_5400;
assign v_5405 = v_5403 | v_5404;
assign v_5406 = v_4826 | v_4828;
assign v_5409 = v_5402 | v_5407 | v_5408;
assign v_5414 = v_5410 | v_5411 | v_5412 | v_5413;
assign v_5417 = v_5415 | v_5416;
assign v_5421 = v_5419 | v_5420;
assign v_5422 = v_4884 | v_4886;
assign v_5425 = v_5418 | v_5423 | v_5424;
assign v_5433 = v_5431 | v_5432;
assign v_5435 = v_5430 | v_5434;
assign v_5437 = v_5429 | v_5436;
assign v_5439 = v_5428 | v_5438;
assign v_5441 = v_5427 | v_5440;
assign v_5443 = v_5426 | v_5442;
assign v_5448 = v_5446 | v_5447;
assign v_5454 = v_5450 | v_5451 | v_5452 | v_5453;
assign v_5456 = v_5449 | v_5455;
assign v_5460 = v_5444 | v_5445 | v_5457 | v_5458 | v_5459;
assign v_5464 = v_5462 | v_5463;
assign v_5466 = v_4986 | v_4988;
assign v_5470 = v_5468 | v_5469;
assign v_5473 = v_5471 | v_5472;
assign v_5478 = v_5476 | v_5477;
assign v_5480 = v_7922 | v_7923;
assign v_5487 = v_5485 | v_5486;
assign v_5488 = v_7924 | v_7925;
assign v_5492 = v_5489 | v_5490 | v_5491;
assign v_5494 = v_5482 | v_5483 | v_5484 | v_5493;
assign v_5497 = v_5481 | v_5495 | v_5496;
assign v_5499 = v_4550 | v_4552;
assign v_5502 = v_5498 | v_5500 | v_5501;
assign v_5503 = v_4564 | v_4566;
assign v_5509 = v_5506 | v_5507 | v_5508;
assign v_5511 = v_5505 | v_5510;
assign v_5513 = v_5504 | v_5512;
assign v_5514 = ~v_4589 | v_4591 | v_4593;
assign v_5517 = v_5515 | v_5516;
assign v_5526 = v_5524 | v_5525;
assign v_5528 = v_5522 | v_5523 | v_5527;
assign v_5533 = v_4636 | v_4638;
assign v_5536 = v_5534 | v_5535;
assign v_5539 = v_5537 | v_5538;
assign v_5541 = v_5530 | v_5531 | v_5532 | v_5540;
assign v_5547 = v_5543 | v_5544 | v_5545 | v_5546;
assign v_5549 = v_5529 | v_5542 | v_5548;
assign v_5551 = v_5518 | v_5519 | v_5520 | v_5521 | v_5550;
assign v_5560 = v_5558 | v_5559;
assign v_5562 = v_5556 | v_5557 | v_5561;
assign v_5567 = v_4701 | v_4703;
assign v_5570 = v_5568 | v_5569;
assign v_5573 = v_5571 | v_5572;
assign v_5575 = v_5564 | v_5565 | v_5566 | v_5574;
assign v_5581 = v_5577 | v_5578 | v_5579 | v_5580;
assign v_5583 = v_5563 | v_5576 | v_5582;
assign v_5585 = v_5552 | v_5553 | v_5554 | v_5555 | v_5584;
assign v_5592 = v_5590 | v_5591;
assign v_5593 = v_7926 | v_7927;
assign v_5597 = v_5594 | v_5595 | v_5596;
assign v_5599 = v_5587 | v_5588 | v_5589 | v_5598;
assign v_5602 = v_5586 | v_5600 | v_5601;
assign v_5607 = v_5604 | v_5606;
assign v_5609 = v_5603 | v_5608;
assign v_5613 = v_5611 | v_5612;
assign v_5614 = v_4826 | v_4828;
assign v_5617 = v_5610 | v_5615 | v_5616;
assign v_5622 = v_5618 | v_5619 | v_5620 | v_5621;
assign v_5627 = v_5624 | v_5626;
assign v_5629 = v_5623 | v_5628;
assign v_5633 = v_5631 | v_5632;
assign v_5634 = v_4884 | v_4886;
assign v_5637 = v_5630 | v_5635 | v_5636;
assign v_5645 = v_5643 | v_5644;
assign v_5647 = v_5642 | v_5646;
assign v_5649 = v_5641 | v_5648;
assign v_5651 = v_5640 | v_5650;
assign v_5653 = v_5639 | v_5652;
assign v_5655 = v_5638 | v_5654;
assign v_5660 = v_5658 | v_5659;
assign v_5666 = v_5662 | v_5663 | v_5664 | v_5665;
assign v_5668 = v_5661 | v_5667;
assign v_5672 = v_5656 | v_5657 | v_5669 | v_5670 | v_5671;
assign v_5678 = v_5675 | v_5677;
assign v_5680 = v_5674 | v_5679;
assign v_5682 = v_4986 | v_4988;
assign v_5686 = v_5684 | v_5685;
assign v_5689 = v_5687 | v_5688;
assign v_5696 = v_5693 | v_5695;
assign v_5698 = v_5692 | v_5697;
assign v_5700 = v_7928 | v_7929;
assign v_5706 = v_7930 | v_7931;
assign v_5710 = v_5707 | v_5708 | v_5709;
assign v_5712 = v_5702 | v_5703 | v_5704 | v_5711;
assign v_5715 = v_5701 | v_5713 | v_5714;
assign v_5717 = v_4550 | v_4552;
assign v_5720 = v_5716 | v_5718 | v_5719;
assign v_5721 = v_4564 | v_4566;
assign v_5727 = v_5724 | v_5725 | v_5726;
assign v_5729 = v_5723 | v_5728;
assign v_5731 = v_5722 | v_5730;
assign v_5732 = ~v_4589 | v_4591 | v_4593;
assign v_5735 = v_5733 | v_5734;
assign v_5744 = v_5742 | v_5743;
assign v_5746 = v_5740 | v_5741 | v_5745;
assign v_5751 = v_4636 | v_4638;
assign v_5754 = v_5752 | v_5753;
assign v_5757 = v_5755 | v_5756;
assign v_5759 = v_5748 | v_5749 | v_5750 | v_5758;
assign v_5765 = v_5761 | v_5762 | v_5763 | v_5764;
assign v_5767 = v_5747 | v_5760 | v_5766;
assign v_5769 = v_5736 | v_5737 | v_5738 | v_5739 | v_5768;
assign v_5778 = v_5776 | v_5777;
assign v_5780 = v_5774 | v_5775 | v_5779;
assign v_5785 = v_4701 | v_4703;
assign v_5788 = v_5786 | v_5787;
assign v_5791 = v_5789 | v_5790;
assign v_5793 = v_5782 | v_5783 | v_5784 | v_5792;
assign v_5799 = v_5795 | v_5796 | v_5797 | v_5798;
assign v_5801 = v_5781 | v_5794 | v_5800;
assign v_5803 = v_5770 | v_5771 | v_5772 | v_5773 | v_5802;
assign v_5810 = v_5808 | v_5809;
assign v_5811 = v_7932 | v_7933;
assign v_5815 = v_5812 | v_5813 | v_5814;
assign v_5817 = v_5805 | v_5806 | v_5807 | v_5816;
assign v_5820 = v_5804 | v_5818 | v_5819;
assign v_5825 = v_5822 | v_5824;
assign v_5827 = v_5821 | v_5826;
assign v_5831 = v_5829 | v_5830;
assign v_5832 = v_4826 | v_4828;
assign v_5835 = v_5828 | v_5833 | v_5834;
assign v_5840 = v_5836 | v_5837 | v_5838 | v_5839;
assign v_5845 = v_5842 | v_5844;
assign v_5847 = v_5841 | v_5846;
assign v_5851 = v_5849 | v_5850;
assign v_5852 = v_4884 | v_4886;
assign v_5855 = v_5848 | v_5853 | v_5854;
assign v_5863 = v_5861 | v_5862;
assign v_5865 = v_5860 | v_5864;
assign v_5867 = v_5859 | v_5866;
assign v_5869 = v_5858 | v_5868;
assign v_5871 = v_5857 | v_5870;
assign v_5873 = v_5856 | v_5872;
assign v_5878 = v_5876 | v_5877;
assign v_5884 = v_5880 | v_5881 | v_5882 | v_5883;
assign v_5886 = v_5879 | v_5885;
assign v_5890 = v_5874 | v_5875 | v_5887 | v_5888 | v_5889;
assign v_5896 = v_5893 | v_5895;
assign v_5898 = v_5892 | v_5897;
assign v_5900 = v_4986 | v_4988;
assign v_5904 = v_5902 | v_5903;
assign v_5907 = v_5905 | v_5906;
assign v_5914 = v_5911 | v_5913;
assign v_5916 = v_5910 | v_5915;
assign v_5918 = v_7934 | v_7935;
assign v_5926 = v_5924 | v_5925;
assign v_5927 = v_7936 | v_7937;
assign v_5931 = v_5928 | v_5929 | v_5930;
assign v_5933 = v_5921 | v_5922 | v_5923 | v_5932;
assign v_5936 = v_5920 | v_5934 | v_5935;
assign v_5938 = v_4550 | v_4552;
assign v_5941 = v_5937 | v_5939 | v_5940;
assign v_5942 = v_4564 | v_4566;
assign v_5948 = v_5945 | v_5946 | v_5947;
assign v_5950 = v_5944 | v_5949;
assign v_5952 = v_5943 | v_5951;
assign v_5953 = ~v_4589 | v_4591 | v_4593;
assign v_5956 = v_5954 | v_5955;
assign v_5965 = v_5963 | v_5964;
assign v_5967 = v_5961 | v_5962 | v_5966;
assign v_5972 = v_4636 | v_4638;
assign v_5975 = v_5973 | v_5974;
assign v_5978 = v_5976 | v_5977;
assign v_5980 = v_5969 | v_5970 | v_5971 | v_5979;
assign v_5986 = v_5982 | v_5983 | v_5984 | v_5985;
assign v_5988 = v_5968 | v_5981 | v_5987;
assign v_5990 = v_5957 | v_5958 | v_5959 | v_5960 | v_5989;
assign v_5999 = v_5997 | v_5998;
assign v_6001 = v_5995 | v_5996 | v_6000;
assign v_6006 = v_4701 | v_4703;
assign v_6009 = v_6007 | v_6008;
assign v_6012 = v_6010 | v_6011;
assign v_6014 = v_6003 | v_6004 | v_6005 | v_6013;
assign v_6020 = v_6016 | v_6017 | v_6018 | v_6019;
assign v_6022 = v_6002 | v_6015 | v_6021;
assign v_6024 = v_5991 | v_5992 | v_5993 | v_5994 | v_6023;
assign v_6031 = v_6029 | v_6030;
assign v_6032 = v_7938 | v_7939;
assign v_6036 = v_6033 | v_6034 | v_6035;
assign v_6038 = v_6026 | v_6027 | v_6028 | v_6037;
assign v_6041 = v_6025 | v_6039 | v_6040;
assign v_6046 = v_6043 | v_6045;
assign v_6048 = v_6042 | v_6047;
assign v_6052 = v_6050 | v_6051;
assign v_6053 = v_4826 | v_4828;
assign v_6056 = v_6049 | v_6054 | v_6055;
assign v_6061 = v_6057 | v_6058 | v_6059 | v_6060;
assign v_6066 = v_6063 | v_6065;
assign v_6068 = v_6062 | v_6067;
assign v_6072 = v_6070 | v_6071;
assign v_6073 = v_4884 | v_4886;
assign v_6076 = v_6069 | v_6074 | v_6075;
assign v_6084 = v_6082 | v_6083;
assign v_6086 = v_6081 | v_6085;
assign v_6088 = v_6080 | v_6087;
assign v_6090 = v_6079 | v_6089;
assign v_6092 = v_6078 | v_6091;
assign v_6094 = v_6077 | v_6093;
assign v_6099 = v_6097 | v_6098;
assign v_6105 = v_6101 | v_6102 | v_6103 | v_6104;
assign v_6107 = v_6100 | v_6106;
assign v_6111 = v_6095 | v_6096 | v_6108 | v_6109 | v_6110;
assign v_6117 = v_6114 | v_6116;
assign v_6119 = v_6113 | v_6118;
assign v_6121 = v_4986 | v_4988;
assign v_6125 = v_6123 | v_6124;
assign v_6128 = v_6126 | v_6127;
assign v_6135 = v_6132 | v_6134;
assign v_6137 = v_6131 | v_6136;
assign v_6139 = v_7940 | v_7941;
assign v_6147 = v_6145 | v_6146;
assign v_6148 = v_7942 | v_7943;
assign v_6152 = v_6149 | v_6150 | v_6151;
assign v_6154 = v_6142 | v_6143 | v_6144 | v_6153;
assign v_6157 = v_6141 | v_6155 | v_6156;
assign v_6159 = v_4550 | v_4552;
assign v_6162 = v_6158 | v_6160 | v_6161;
assign v_6163 = v_4564 | v_4566;
assign v_6169 = v_6166 | v_6167 | v_6168;
assign v_6171 = v_6165 | v_6170;
assign v_6173 = v_6164 | v_6172;
assign v_6174 = ~v_4589 | v_4591 | v_4593;
assign v_6177 = v_6175 | v_6176;
assign v_6186 = v_6184 | v_6185;
assign v_6188 = v_6182 | v_6183 | v_6187;
assign v_6193 = v_4636 | v_4638;
assign v_6196 = v_6194 | v_6195;
assign v_6199 = v_6197 | v_6198;
assign v_6201 = v_6190 | v_6191 | v_6192 | v_6200;
assign v_6207 = v_6203 | v_6204 | v_6205 | v_6206;
assign v_6209 = v_6189 | v_6202 | v_6208;
assign v_6211 = v_6178 | v_6179 | v_6180 | v_6181 | v_6210;
assign v_6220 = v_6218 | v_6219;
assign v_6222 = v_6216 | v_6217 | v_6221;
assign v_6227 = v_4701 | v_4703;
assign v_6230 = v_6228 | v_6229;
assign v_6233 = v_6231 | v_6232;
assign v_6235 = v_6224 | v_6225 | v_6226 | v_6234;
assign v_6241 = v_6237 | v_6238 | v_6239 | v_6240;
assign v_6243 = v_6223 | v_6236 | v_6242;
assign v_6245 = v_6212 | v_6213 | v_6214 | v_6215 | v_6244;
assign v_6252 = v_6250 | v_6251;
assign v_6253 = v_7944 | v_7945;
assign v_6257 = v_6254 | v_6255 | v_6256;
assign v_6259 = v_6247 | v_6248 | v_6249 | v_6258;
assign v_6262 = v_6246 | v_6260 | v_6261;
assign v_6267 = v_6264 | v_6266;
assign v_6269 = v_6263 | v_6268;
assign v_6273 = v_6271 | v_6272;
assign v_6274 = v_4826 | v_4828;
assign v_6277 = v_6270 | v_6275 | v_6276;
assign v_6282 = v_6278 | v_6279 | v_6280 | v_6281;
assign v_6287 = v_6284 | v_6286;
assign v_6289 = v_6283 | v_6288;
assign v_6293 = v_6291 | v_6292;
assign v_6294 = v_4884 | v_4886;
assign v_6297 = v_6290 | v_6295 | v_6296;
assign v_6305 = v_6303 | v_6304;
assign v_6307 = v_6302 | v_6306;
assign v_6309 = v_6301 | v_6308;
assign v_6311 = v_6300 | v_6310;
assign v_6313 = v_6299 | v_6312;
assign v_6315 = v_6298 | v_6314;
assign v_6320 = v_6318 | v_6319;
assign v_6326 = v_6322 | v_6323 | v_6324 | v_6325;
assign v_6328 = v_6321 | v_6327;
assign v_6332 = v_6316 | v_6317 | v_6329 | v_6330 | v_6331;
assign v_6338 = v_6335 | v_6337;
assign v_6340 = v_6334 | v_6339;
assign v_6342 = v_4986 | v_4988;
assign v_6346 = v_6344 | v_6345;
assign v_6349 = v_6347 | v_6348;
assign v_6356 = v_6353 | v_6355;
assign v_6358 = v_6352 | v_6357;
assign v_6360 = v_7946 | v_7947;
assign v_6367 = v_6365 | v_6366;
assign v_6368 = v_7948 | v_7949;
assign v_6372 = v_6369 | v_6370 | v_6371;
assign v_6374 = v_6362 | v_6363 | v_6364 | v_6373;
assign v_6377 = v_6361 | v_6375 | v_6376;
assign v_6379 = v_4550 | v_4552;
assign v_6382 = v_6378 | v_6380 | v_6381;
assign v_6383 = v_4564 | v_4566;
assign v_6389 = v_6386 | v_6387 | v_6388;
assign v_6391 = v_6385 | v_6390;
assign v_6393 = v_6384 | v_6392;
assign v_6394 = ~v_4589 | v_4591 | v_4593;
assign v_6397 = v_6395 | v_6396;
assign v_6406 = v_6404 | v_6405;
assign v_6408 = v_6402 | v_6403 | v_6407;
assign v_6413 = v_4636 | v_4638;
assign v_6416 = v_6414 | v_6415;
assign v_6419 = v_6417 | v_6418;
assign v_6421 = v_6410 | v_6411 | v_6412 | v_6420;
assign v_6427 = v_6423 | v_6424 | v_6425 | v_6426;
assign v_6429 = v_6409 | v_6422 | v_6428;
assign v_6431 = v_6398 | v_6399 | v_6400 | v_6401 | v_6430;
assign v_6440 = v_6438 | v_6439;
assign v_6442 = v_6436 | v_6437 | v_6441;
assign v_6447 = v_4701 | v_4703;
assign v_6450 = v_6448 | v_6449;
assign v_6453 = v_6451 | v_6452;
assign v_6455 = v_6444 | v_6445 | v_6446 | v_6454;
assign v_6461 = v_6457 | v_6458 | v_6459 | v_6460;
assign v_6463 = v_6443 | v_6456 | v_6462;
assign v_6465 = v_6432 | v_6433 | v_6434 | v_6435 | v_6464;
assign v_6472 = v_6470 | v_6471;
assign v_6473 = v_7950 | v_7951;
assign v_6477 = v_6474 | v_6475 | v_6476;
assign v_6479 = v_6467 | v_6468 | v_6469 | v_6478;
assign v_6482 = v_6466 | v_6480 | v_6481;
assign v_6487 = v_6484 | v_6486;
assign v_6489 = v_6483 | v_6488;
assign v_6493 = v_6491 | v_6492;
assign v_6494 = v_4826 | v_4828;
assign v_6497 = v_6490 | v_6495 | v_6496;
assign v_6502 = v_6498 | v_6499 | v_6500 | v_6501;
assign v_6507 = v_6504 | v_6506;
assign v_6509 = v_6503 | v_6508;
assign v_6513 = v_6511 | v_6512;
assign v_6514 = v_4884 | v_4886;
assign v_6517 = v_6510 | v_6515 | v_6516;
assign v_6525 = v_6523 | v_6524;
assign v_6527 = v_6522 | v_6526;
assign v_6529 = v_6521 | v_6528;
assign v_6531 = v_6520 | v_6530;
assign v_6533 = v_6519 | v_6532;
assign v_6535 = v_6518 | v_6534;
assign v_6540 = v_6538 | v_6539;
assign v_6546 = v_6542 | v_6543 | v_6544 | v_6545;
assign v_6548 = v_6541 | v_6547;
assign v_6552 = v_6536 | v_6537 | v_6549 | v_6550 | v_6551;
assign v_6558 = v_6555 | v_6557;
assign v_6560 = v_6554 | v_6559;
assign v_6562 = v_4986 | v_4988;
assign v_6566 = v_6564 | v_6565;
assign v_6569 = v_6567 | v_6568;
assign v_6576 = v_6573 | v_6575;
assign v_6578 = v_6572 | v_6577;
assign v_6580 = v_7952 | v_7953;
assign v_6588 = v_6586 | v_6587;
assign v_6589 = v_7954 | v_7955;
assign v_6593 = v_6590 | v_6591 | v_6592;
assign v_6595 = v_6583 | v_6584 | v_6585 | v_6594;
assign v_6598 = v_6582 | v_6596 | v_6597;
assign v_6600 = v_4550 | v_4552;
assign v_6603 = v_6599 | v_6601 | v_6602;
assign v_6604 = v_4564 | v_4566;
assign v_6610 = v_6607 | v_6608 | v_6609;
assign v_6612 = v_6606 | v_6611;
assign v_6614 = v_6605 | v_6613;
assign v_6615 = ~v_4589 | v_4591 | v_4593;
assign v_6618 = v_6616 | v_6617;
assign v_6627 = v_6625 | v_6626;
assign v_6629 = v_6623 | v_6624 | v_6628;
assign v_6634 = v_4636 | v_4638;
assign v_6637 = v_6635 | v_6636;
assign v_6640 = v_6638 | v_6639;
assign v_6642 = v_6631 | v_6632 | v_6633 | v_6641;
assign v_6648 = v_6644 | v_6645 | v_6646 | v_6647;
assign v_6650 = v_6630 | v_6643 | v_6649;
assign v_6652 = v_6619 | v_6620 | v_6621 | v_6622 | v_6651;
assign v_6661 = v_6659 | v_6660;
assign v_6663 = v_6657 | v_6658 | v_6662;
assign v_6668 = v_4701 | v_4703;
assign v_6671 = v_6669 | v_6670;
assign v_6674 = v_6672 | v_6673;
assign v_6676 = v_6665 | v_6666 | v_6667 | v_6675;
assign v_6682 = v_6678 | v_6679 | v_6680 | v_6681;
assign v_6684 = v_6664 | v_6677 | v_6683;
assign v_6686 = v_6653 | v_6654 | v_6655 | v_6656 | v_6685;
assign v_6693 = v_6691 | v_6692;
assign v_6694 = v_7956 | v_7957;
assign v_6698 = v_6695 | v_6696 | v_6697;
assign v_6700 = v_6688 | v_6689 | v_6690 | v_6699;
assign v_6703 = v_6687 | v_6701 | v_6702;
assign v_6708 = v_6705 | v_6707;
assign v_6710 = v_6704 | v_6709;
assign v_6714 = v_6712 | v_6713;
assign v_6715 = v_4826 | v_4828;
assign v_6718 = v_6711 | v_6716 | v_6717;
assign v_6723 = v_6719 | v_6720 | v_6721 | v_6722;
assign v_6728 = v_6725 | v_6727;
assign v_6730 = v_6724 | v_6729;
assign v_6734 = v_6732 | v_6733;
assign v_6735 = v_4884 | v_4886;
assign v_6738 = v_6731 | v_6736 | v_6737;
assign v_6746 = v_6744 | v_6745;
assign v_6748 = v_6743 | v_6747;
assign v_6750 = v_6742 | v_6749;
assign v_6752 = v_6741 | v_6751;
assign v_6754 = v_6740 | v_6753;
assign v_6756 = v_6739 | v_6755;
assign v_6761 = v_6759 | v_6760;
assign v_6767 = v_6763 | v_6764 | v_6765 | v_6766;
assign v_6769 = v_6762 | v_6768;
assign v_6773 = v_6757 | v_6758 | v_6770 | v_6771 | v_6772;
assign v_6779 = v_6776 | v_6778;
assign v_6781 = v_6775 | v_6780;
assign v_6783 = v_4986 | v_4988;
assign v_6787 = v_6785 | v_6786;
assign v_6790 = v_6788 | v_6789;
assign v_6797 = v_6794 | v_6796;
assign v_6799 = v_6793 | v_6798;
assign v_6801 = v_7958 | v_7959;
assign v_6804 = v_6803 | ~v_5099;
assign v_6810 = v_6806 | v_6808 | v_6809;
assign v_6812 = v_4550 | v_4552;
assign v_6815 = v_6811 | v_6813 | v_6814;
assign v_6816 = v_4564 | v_4566;
assign v_6822 = v_6819 | v_6820 | v_6821;
assign v_6824 = v_6818 | v_6823;
assign v_6826 = v_6817 | v_6825;
assign v_6827 = ~v_4589 | v_4591 | v_4593;
assign v_6830 = v_6828 | v_6829;
assign v_6832 = v_6805 | v_6831;
assign v_6841 = v_6839 | v_6840;
assign v_6843 = v_6837 | v_6838 | v_6842;
assign v_6848 = v_4636 | v_4638;
assign v_6851 = v_6849 | v_6850;
assign v_6854 = v_6852 | v_6853;
assign v_6856 = v_6845 | v_6846 | v_6847 | v_6855;
assign v_6862 = v_6858 | v_6859 | v_6860 | v_6861;
assign v_6864 = v_6844 | v_6857 | v_6863;
assign v_6866 = v_6833 | v_6834 | v_6835 | v_6836 | v_6865;
assign v_6875 = v_6873 | v_6874;
assign v_6877 = v_6871 | v_6872 | v_6876;
assign v_6882 = v_4701 | v_4703;
assign v_6885 = v_6883 | v_6884;
assign v_6888 = v_6886 | v_6887;
assign v_6890 = v_6879 | v_6880 | v_6881 | v_6889;
assign v_6896 = v_6892 | v_6893 | v_6894 | v_6895;
assign v_6898 = v_6878 | v_6891 | v_6897;
assign v_6900 = v_6867 | v_6868 | v_6869 | v_6870 | v_6899;
assign v_6905 = v_6901 | v_6903 | v_6904;
assign v_6908 = v_6906 | v_6907;
assign v_6912 = v_6910 | v_6911;
assign v_6913 = v_4826 | v_4828;
assign v_6916 = v_6909 | v_6914 | v_6915;
assign v_6921 = v_6917 | v_6918 | v_6919 | v_6920;
assign v_6924 = v_6922 | v_6923;
assign v_6928 = v_6926 | v_6927;
assign v_6929 = v_4884 | v_4886;
assign v_6932 = v_6925 | v_6930 | v_6931;
assign v_6940 = v_6938 | v_6939;
assign v_6942 = v_6937 | v_6941;
assign v_6944 = v_6936 | v_6943;
assign v_6946 = v_6935 | v_6945;
assign v_6948 = v_6934 | v_6947;
assign v_6950 = v_6933 | v_6949;
assign v_6955 = v_6953 | v_6954;
assign v_6961 = v_6957 | v_6958 | v_6959 | v_6960;
assign v_6963 = v_6956 | v_6962;
assign v_6967 = v_6951 | v_6952 | v_6964 | v_6965 | v_6966;
assign v_6971 = v_6969 | v_6970;
assign v_6973 = v_4986 | v_4988;
assign v_6977 = v_6975 | v_6976;
assign v_6980 = v_6978 | v_6979;
assign v_6985 = v_6983 | v_6984;
assign v_6987 = v_7960 | v_7961;
assign v_6995 = v_6993 | v_6994;
assign v_6996 = v_7962 | v_7963;
assign v_7000 = v_6997 | v_6998 | v_6999;
assign v_7002 = v_6990 | v_6991 | v_6992 | v_7001;
assign v_7005 = v_6989 | v_7003 | v_7004;
assign v_7007 = v_4550 | v_4552;
assign v_7010 = v_7006 | v_7008 | v_7009;
assign v_7011 = v_4564 | v_4566;
assign v_7017 = v_7014 | v_7015 | v_7016;
assign v_7019 = v_7013 | v_7018;
assign v_7021 = v_7012 | v_7020;
assign v_7022 = ~v_4589 | v_4591 | v_4593;
assign v_7025 = v_7023 | v_7024;
assign v_7034 = v_7032 | v_7033;
assign v_7036 = v_7030 | v_7031 | v_7035;
assign v_7041 = v_4636 | v_4638;
assign v_7044 = v_7042 | v_7043;
assign v_7047 = v_7045 | v_7046;
assign v_7049 = v_7038 | v_7039 | v_7040 | v_7048;
assign v_7055 = v_7051 | v_7052 | v_7053 | v_7054;
assign v_7057 = v_7037 | v_7050 | v_7056;
assign v_7059 = v_7026 | v_7027 | v_7028 | v_7029 | v_7058;
assign v_7068 = v_7066 | v_7067;
assign v_7070 = v_7064 | v_7065 | v_7069;
assign v_7075 = v_4701 | v_4703;
assign v_7078 = v_7076 | v_7077;
assign v_7081 = v_7079 | v_7080;
assign v_7083 = v_7072 | v_7073 | v_7074 | v_7082;
assign v_7089 = v_7085 | v_7086 | v_7087 | v_7088;
assign v_7091 = v_7071 | v_7084 | v_7090;
assign v_7093 = v_7060 | v_7061 | v_7062 | v_7063 | v_7092;
assign v_7100 = v_7098 | v_7099;
assign v_7101 = v_7964 | v_7965;
assign v_7105 = v_7102 | v_7103 | v_7104;
assign v_7107 = v_7095 | v_7096 | v_7097 | v_7106;
assign v_7110 = v_7094 | v_7108 | v_7109;
assign v_7115 = v_7112 | v_7114;
assign v_7117 = v_7111 | v_7116;
assign v_7121 = v_7119 | v_7120;
assign v_7122 = v_4826 | v_4828;
assign v_7125 = v_7118 | v_7123 | v_7124;
assign v_7130 = v_7126 | v_7127 | v_7128 | v_7129;
assign v_7135 = v_7132 | v_7134;
assign v_7137 = v_7131 | v_7136;
assign v_7141 = v_7139 | v_7140;
assign v_7142 = v_4884 | v_4886;
assign v_7145 = v_7138 | v_7143 | v_7144;
assign v_7153 = v_7151 | v_7152;
assign v_7155 = v_7150 | v_7154;
assign v_7157 = v_7149 | v_7156;
assign v_7159 = v_7148 | v_7158;
assign v_7161 = v_7147 | v_7160;
assign v_7163 = v_7146 | v_7162;
assign v_7168 = v_7166 | v_7167;
assign v_7174 = v_7170 | v_7171 | v_7172 | v_7173;
assign v_7176 = v_7169 | v_7175;
assign v_7180 = v_7164 | v_7165 | v_7177 | v_7178 | v_7179;
assign v_7186 = v_7183 | v_7185;
assign v_7188 = v_7182 | v_7187;
assign v_7190 = v_4986 | v_4988;
assign v_7194 = v_7192 | v_7193;
assign v_7197 = v_7195 | v_7196;
assign v_7204 = v_7201 | v_7203;
assign v_7206 = v_7200 | v_7205;
assign v_7208 = v_7966 | v_7967;
assign v_7759 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_7760 = v_244 | v_246 | v_248 | v_252 | v_253;
assign v_7761 = v_259;
assign v_7762 = v_393 | v_395 | v_397 | v_399 | v_401;
assign v_7763 = v_402;
assign v_7764 = v_347 | v_349 | v_351 | v_358 | v_407;
assign v_7765 = v_408;
assign v_7766 = v_458 | v_460 | v_462 | v_464 | v_466;
assign v_7767 = v_467;
assign v_7768 = v_412 | v_414 | v_416 | v_423 | v_472;
assign v_7769 = v_473;
assign v_7770 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_7771 = v_508 | v_510 | v_512 | v_516 | v_517;
assign v_7772 = v_523;
assign v_7773 = ~v_669 | v_671 | v_673 | v_676 | v_681;
assign v_7774 = v_683 | v_701 | v_702;
assign v_7775 = ~v_705 | v_725 | v_730 | v_732 | v_774;
assign v_7776 = v_793 | v_794 | v_795;
assign v_7777 = v_816 | v_818 | v_839 | v_841 | v_862;
assign v_7778 = v_864 | v_871 | v_873 | v_874 | v_875;
assign v_7779 = v_876;
assign v_7780 = v_897 | v_899 | v_920 | v_922 | v_943;
assign v_7781 = v_945 | v_952 | v_954 | v_955 | v_956;
assign v_7782 = v_957;
assign v_7783 = v_978 | v_980 | v_1001 | v_1003 | v_1024;
assign v_7784 = v_1026 | v_1033 | v_1035 | v_1036 | v_1037;
assign v_7785 = v_1038;
assign v_7786 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_7787 = v_244 | v_246 | v_248;
assign v_7788 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_7789 = v_508 | v_510 | v_512;
assign v_7790 = v_1260 | v_1264 | v_1266 | v_1273 | v_1274;
assign v_7791 = v_1279;
assign v_7792 = v_1281 | v_1290 | v_1299 | v_1305 | v_1316;
assign v_7793 = v_1317 | v_1318;
assign v_7794 = v_1320 | v_1329 | v_1338 | v_1344 | v_1355;
assign v_7795 = v_1356 | v_1357;
assign v_7796 = v_1359 | v_1368 | v_1377 | v_1383 | v_1394;
assign v_7797 = v_1395 | v_1396;
assign v_7798 = v_1565 | v_1569 | v_1571 | v_1578 | v_1579;
assign v_7799 = v_1583;
assign v_7800 = v_1585 | v_1593 | v_1601 | v_1606 | v_1616;
assign v_7801 = v_1617 | v_1618;
assign v_7802 = v_1620 | v_1628 | v_1636 | v_1641 | v_1651;
assign v_7803 = v_1652 | v_1653;
assign v_7804 = v_1655 | v_1663 | v_1671 | v_1676 | v_1686;
assign v_7805 = v_1687 | v_1688;
assign v_7806 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_7807 = v_244 | v_246 | v_248;
assign v_7808 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_7809 = v_508 | v_510 | v_512;
assign v_7810 = v_1882 | v_1890 | v_1892 | v_1899 | v_1900;
assign v_7811 = v_1908;
assign v_7812 = v_1910 | v_1918 | v_1926 | v_1931 | v_1941;
assign v_7813 = v_1942 | v_1943;
assign v_7814 = v_1945 | v_1953 | v_1961 | v_1966 | v_1976;
assign v_7815 = v_1977 | v_1978;
assign v_7816 = v_1980 | v_1988 | v_1996 | v_2001 | v_2011;
assign v_7817 = v_2012 | v_2013;
assign v_7818 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_7819 = v_244 | v_246 | v_248;
assign v_7820 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_7821 = v_508 | v_510 | v_512;
assign v_7822 = v_2205 | v_2213 | v_2215 | v_2222 | v_2223;
assign v_7823 = v_2231;
assign v_7824 = v_2233 | v_2241 | v_2249 | v_2254 | v_2264;
assign v_7825 = v_2265 | v_2266;
assign v_7826 = v_2268 | v_2276 | v_2284 | v_2289 | v_2299;
assign v_7827 = v_2300 | v_2301;
assign v_7828 = v_2303 | v_2311 | v_2319 | v_2324 | v_2334;
assign v_7829 = v_2335 | v_2336;
assign v_7830 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_7831 = v_244 | v_246 | v_248;
assign v_7832 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_7833 = v_508 | v_510 | v_512;
assign v_7834 = v_2531 | v_2539 | v_2541 | v_2548 | v_2549;
assign v_7835 = v_2557;
assign v_7836 = v_2559 | v_2567 | v_2575 | v_2580 | v_2590;
assign v_7837 = v_2591 | v_2592;
assign v_7838 = v_2594 | v_2602 | v_2610 | v_2615 | v_2625;
assign v_7839 = v_2626 | v_2627;
assign v_7840 = v_2629 | v_2637 | v_2645 | v_2650 | v_2660;
assign v_7841 = v_2661 | v_2662;
assign v_7842 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_7843 = v_244 | v_246 | v_248;
assign v_7844 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_7845 = v_508 | v_510 | v_512;
assign v_7846 = v_2857 | v_2865 | v_2867 | v_2874 | v_2875;
assign v_7847 = v_2883;
assign v_7848 = v_2885 | v_2893 | v_2901 | v_2906 | v_2916;
assign v_7849 = v_2917 | v_2918;
assign v_7850 = v_2920 | v_2928 | v_2936 | v_2941 | v_2951;
assign v_7851 = v_2952 | v_2953;
assign v_7852 = v_2955 | v_2963 | v_2971 | v_2976 | v_2986;
assign v_7853 = v_2987 | v_2988;
assign v_7854 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_7855 = v_244 | v_246 | v_248;
assign v_7856 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_7857 = v_508 | v_510 | v_512;
assign v_7858 = v_3182 | v_3190 | v_3192 | v_3199 | v_3200;
assign v_7859 = v_3208;
assign v_7860 = v_3210 | v_3218 | v_3226 | v_3231 | v_3241;
assign v_7861 = v_3242 | v_3243;
assign v_7862 = v_3245 | v_3253 | v_3261 | v_3266 | v_3276;
assign v_7863 = v_3277 | v_3278;
assign v_7864 = v_3280 | v_3288 | v_3296 | v_3301 | v_3311;
assign v_7865 = v_3312 | v_3313;
assign v_7866 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_7867 = v_244 | v_246 | v_248;
assign v_7868 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_7869 = v_508 | v_510 | v_512;
assign v_7870 = v_3508 | v_3516 | v_3518 | v_3525 | v_3526;
assign v_7871 = v_3534;
assign v_7872 = v_3536 | v_3544 | v_3552 | v_3557 | v_3567;
assign v_7873 = v_3568 | v_3569;
assign v_7874 = v_3571 | v_3579 | v_3587 | v_3592 | v_3602;
assign v_7875 = v_3603 | v_3604;
assign v_7876 = v_3606 | v_3614 | v_3622 | v_3627 | v_3637;
assign v_7877 = v_3638 | v_3639;
assign v_7878 = v_3807 | v_3811 | v_3813 | v_3820 | v_3821;
assign v_7879 = v_3825;
assign v_7880 = v_3827 | v_3835 | v_3843 | v_3848 | v_3858;
assign v_7881 = v_3859 | v_3860;
assign v_7882 = v_3862 | v_3870 | v_3878 | v_3883 | v_3893;
assign v_7883 = v_3894 | v_3895;
assign v_7884 = v_3897 | v_3905 | v_3913 | v_3918 | v_3928;
assign v_7885 = v_3929 | v_3930;
assign v_7886 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_7887 = v_244 | v_246 | v_248;
assign v_7888 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_7889 = v_508 | v_510 | v_512;
assign v_7890 = v_4125 | v_4133 | v_4135 | v_4142 | v_4143;
assign v_7891 = v_4151;
assign v_7892 = v_4153 | v_4161 | v_4169 | v_4174 | v_4184;
assign v_7893 = v_4185 | v_4186;
assign v_7894 = v_4188 | v_4196 | v_4204 | v_4209 | v_4219;
assign v_7895 = v_4220 | v_4221;
assign v_7896 = v_4223 | v_4231 | v_4239 | v_4244 | v_4254;
assign v_7897 = v_4255 | v_4256;
assign v_7898 = v_4489 | v_4491 | v_4494 | v_4496 | v_4498;
assign v_7899 = v_4500 | v_4502 | v_4504 | v_4508 | v_4509;
assign v_7900 = v_4515;
assign v_7901 = v_4649 | v_4651 | v_4653 | v_4655 | v_4657;
assign v_7902 = v_4658;
assign v_7903 = v_4603 | v_4605 | v_4607 | v_4614 | v_4663;
assign v_7904 = v_4664;
assign v_7905 = v_4714 | v_4716 | v_4718 | v_4720 | v_4722;
assign v_7906 = v_4723;
assign v_7907 = v_4668 | v_4670 | v_4672 | v_4679 | v_4728;
assign v_7908 = v_4729;
assign v_7909 = v_4753 | v_4755 | v_4758 | v_4760 | v_4762;
assign v_7910 = v_4764 | v_4766 | v_4768 | v_4772 | v_4773;
assign v_7911 = v_4779;
assign v_7912 = ~v_4925 | v_4927 | v_4929 | v_4932 | v_4937;
assign v_7913 = v_4939 | v_4957 | v_4958;
assign v_7914 = ~v_4961 | v_4981 | v_4986 | v_4988 | v_5030;
assign v_7915 = v_5049 | v_5050 | v_5051;
assign v_7916 = v_4489 | v_4491 | v_4494 | v_4496 | v_4498;
assign v_7917 = v_4500 | v_4502 | v_4504;
assign v_7918 = v_4753 | v_4755 | v_4758 | v_4760 | v_4762;
assign v_7919 = v_4764 | v_4766 | v_4768;
assign v_7920 = v_5273 | v_5277 | v_5279 | v_5286 | v_5287;
assign v_7921 = v_5292;
assign v_7922 = v_5461 | v_5465 | v_5467 | v_5474 | v_5475;
assign v_7923 = v_5479;
assign v_7924 = v_4489 | v_4491 | v_4494 | v_4496 | v_4498;
assign v_7925 = v_4500 | v_4502 | v_4504;
assign v_7926 = v_4753 | v_4755 | v_4758 | v_4760 | v_4762;
assign v_7927 = v_4764 | v_4766 | v_4768;
assign v_7928 = v_5673 | v_5681 | v_5683 | v_5690 | v_5691;
assign v_7929 = v_5699;
assign v_7930 = v_4489 | v_4491 | v_4494 | v_4496 | v_4498;
assign v_7931 = v_4500 | v_4502 | v_4504;
assign v_7932 = v_4753 | v_4755 | v_4758 | v_4760 | v_4762;
assign v_7933 = v_4764 | v_4766 | v_4768;
assign v_7934 = v_5891 | v_5899 | v_5901 | v_5908 | v_5909;
assign v_7935 = v_5917;
assign v_7936 = v_4489 | v_4491 | v_4494 | v_4496 | v_4498;
assign v_7937 = v_4500 | v_4502 | v_4504;
assign v_7938 = v_4753 | v_4755 | v_4758 | v_4760 | v_4762;
assign v_7939 = v_4764 | v_4766 | v_4768;
assign v_7940 = v_6112 | v_6120 | v_6122 | v_6129 | v_6130;
assign v_7941 = v_6138;
assign v_7942 = v_4489 | v_4491 | v_4494 | v_4496 | v_4498;
assign v_7943 = v_4500 | v_4502 | v_4504;
assign v_7944 = v_4753 | v_4755 | v_4758 | v_4760 | v_4762;
assign v_7945 = v_4764 | v_4766 | v_4768;
assign v_7946 = v_6333 | v_6341 | v_6343 | v_6350 | v_6351;
assign v_7947 = v_6359;
assign v_7948 = v_4489 | v_4491 | v_4494 | v_4496 | v_4498;
assign v_7949 = v_4500 | v_4502 | v_4504;
assign v_7950 = v_4753 | v_4755 | v_4758 | v_4760 | v_4762;
assign v_7951 = v_4764 | v_4766 | v_4768;
assign v_7952 = v_6553 | v_6561 | v_6563 | v_6570 | v_6571;
assign v_7953 = v_6579;
assign v_7954 = v_4489 | v_4491 | v_4494 | v_4496 | v_4498;
assign v_7955 = v_4500 | v_4502 | v_4504;
assign v_7956 = v_4753 | v_4755 | v_4758 | v_4760 | v_4762;
assign v_7957 = v_4764 | v_4766 | v_4768;
assign v_7958 = v_6774 | v_6782 | v_6784 | v_6791 | v_6792;
assign v_7959 = v_6800;
assign v_7960 = v_6968 | v_6972 | v_6974 | v_6981 | v_6982;
assign v_7961 = v_6986;
assign v_7962 = v_4489 | v_4491 | v_4494 | v_4496 | v_4498;
assign v_7963 = v_4500 | v_4502 | v_4504;
assign v_7964 = v_4753 | v_4755 | v_4758 | v_4760 | v_4762;
assign v_7965 = v_4764 | v_4766 | v_4768;
assign v_7966 = v_7181 | v_7189 | v_7191 | v_7198 | v_7199;
assign v_7967 = v_7207;
assign v_7209 = ~v_5293 ^ ~v_1397;
assign v_7210 = ~v_5480 ^ ~v_1689;
assign v_7211 = ~v_5700 ^ ~v_2014;
assign v_7212 = ~v_5918 ^ ~v_2337;
assign v_7213 = ~v_6139 ^ ~v_2663;
assign v_7214 = ~v_6360 ^ ~v_2989;
assign v_7215 = ~v_6580 ^ ~v_3314;
assign v_7216 = ~v_6801 ^ ~v_3640;
assign v_7217 = ~v_6987 ^ ~v_3931;
assign v_7218 = ~v_7208 ^ ~v_4257;
assign x_1 = ~v_1040 | v_7219;
assign o_1 = x_1;
endmodule
