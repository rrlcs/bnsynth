// Benchmark "SKOLEMFORMULA" written by ABC on Tue May 17 15:13:17 2022

module SKOLEMFORMULA ( 
    i0,
    i1  );
  input  i0;
  output i1;
  assign i1 = ~i0;
endmodule


