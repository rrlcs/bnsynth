// skolem function for order file variables
// Generated using findDep.cpp 
module small-pipeline-fixpoint-1 (v_1, v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_12, v_13, v_14, v_15, v_16, v_17, v_18, v_19, v_20, v_21, v_22, v_23, v_24, v_25, v_26, v_27, v_28, v_29, v_30, v_31, v_32, v_33, v_34, v_35, v_36, v_37, v_38, v_39, v_40, v_41, v_42, v_43, v_44, v_45, v_46, v_47, v_48, v_49, v_50, v_51, v_52, v_53, v_54, v_55, v_56, v_57, v_58, v_59, v_60, v_61, v_62, v_63, v_64, v_65, v_66, v_67, v_68, v_69, v_70, v_71, v_72, v_73, v_74, v_75, v_76, v_77, v_78, v_79, v_80, v_81, v_82, v_83, v_84, v_85, v_86, v_87, v_88, v_89, v_90, v_91, v_92, v_93, v_94, v_95, v_96, v_97, v_98, v_99, v_100, v_101, v_102, v_103, v_104, v_105, v_106, v_107, v_108, v_109, v_110, v_111, v_112, v_113, v_114, v_115, v_116, v_117, v_118, v_119, v_120, v_121, v_122, v_123, v_124, v_125, v_126, v_127, v_128, v_129, v_130, v_131, v_132, v_133, v_134, v_135, v_136, v_137, v_138, v_139, v_140, v_141, v_142, v_143, v_144, v_145, v_146, v_147, v_148, v_149, v_150, v_151, v_152, v_153, v_154, v_155, v_156, v_157, v_158, v_159, v_160, v_161, v_162, v_163, v_164, v_165, v_166, v_167, v_168, v_169, v_170, v_171, v_172, v_173, v_174, v_175, v_176, v_177, v_178, v_179, v_180, v_181, v_182, v_183, v_184, v_185, v_186, v_187, v_188, v_189, v_190, v_191, v_192, v_193, v_194, v_195, v_196, v_197, v_198, v_199, v_200, v_201, v_202, v_203, v_204, v_205, v_206, v_207, v_208, v_209, v_210, v_211, v_212, v_213, v_214, v_215, v_216, v_217, v_218, v_219, v_220, v_221, v_222, v_223, v_224, v_225, v_226, v_227, v_228, v_229, v_230, v_231, v_232, v_233, v_234, v_235, v_236, v_237, v_238, v_239, v_240, v_241, v_242, v_243, v_244, v_245, v_246, v_247, v_248, v_249, v_250, v_251, v_252, v_253, v_254, v_255, v_256, v_257, v_258, v_259, v_260, v_261, v_262, v_263, v_264, v_265, v_266, v_267, v_268, v_269, v_270, v_271, v_272, v_273, v_274, v_275, v_276, v_277, v_278, v_279, v_280, v_281, v_282, v_283, v_284, v_285, v_286, v_287, v_288, v_289, v_290, v_291, v_292, v_293, v_294, v_295, v_296, v_297, v_298, v_299, v_300, v_301, v_302, v_303, v_304, v_305, v_306, v_307, v_308, v_309, v_310, v_311, v_312, v_313, v_314, v_315, v_316, v_317, v_318, v_319, v_320, v_321, v_322, v_323, v_324, v_325, v_326, v_327, v_328, v_329, v_330, v_331, v_332, v_333, v_334, v_335, v_336, v_337, v_338, v_339, v_340, v_341, v_342, v_343, v_344, v_345, v_346, v_347, v_348, v_349, v_350, v_351, v_352, v_353, v_354, v_355, v_356, v_357, v_358, v_359, v_360, v_361, v_362, v_363, v_364, v_365, v_366, v_367, v_368, v_369, v_370, v_371, v_372, v_373, v_374, v_375, v_376, v_377, v_378, v_379, v_380, v_381, v_382, v_383, v_384, v_385, v_386, v_387, v_388, v_389, v_390, v_391, v_392, v_393, v_394, v_395, v_396, v_397, v_398, v_399, v_400, v_401, v_402, v_403, v_404, v_405, v_406, v_407, v_408, v_409, v_410, v_411, v_412, v_413, v_414, v_415, v_416, v_417, v_418, v_419, v_420, v_421, v_422, v_423, v_424, v_425, v_426, v_427, v_428, v_429, v_430, v_431, v_432, v_433, v_434, v_435, v_436, v_437, v_438, v_439, v_440, v_441, v_442, v_443, v_444, v_445, v_446, v_447, v_448, v_449, v_450, v_451, v_452, v_453, v_454, v_455, v_456, v_457, v_458, v_459, v_460, v_461, v_462, v_463, v_464, v_465, v_466, v_467, v_468, v_469, v_470, v_471, v_472, v_473, v_474, v_475, v_476, v_477, v_478, v_479, v_480, v_481, v_482, v_483, v_484, v_485, v_486, v_487, v_488, v_489, v_490, v_491, v_492, v_493, v_494, v_495, v_496, v_497, v_498, v_499, v_500, v_501, v_502, v_503, v_504, v_505, v_506, v_507, v_508, v_509, v_510, v_511, v_512, v_513, v_514, v_515, v_516, v_517, v_518, v_519, v_520, v_521, v_522, v_523, v_524, v_525, v_526, v_527, v_528, v_529, v_530, v_531, v_532, v_533, v_534, v_535, v_536, v_537, v_538, v_539, v_540, v_541, v_542, v_543, v_544, v_545, v_546, v_547, v_548, v_549, v_550, v_551, v_552, v_553, v_554, v_555, v_556, v_557, v_558, v_559, v_560, v_561, v_562, v_563, v_564, v_565, v_566, v_567, v_568, v_569, v_570, v_571, v_572, v_573, v_574, v_575, v_576, v_577, o_1);
input v_1;
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_13;
input v_14;
input v_15;
input v_16;
input v_17;
input v_18;
input v_19;
input v_20;
input v_21;
input v_22;
input v_23;
input v_24;
input v_25;
input v_26;
input v_27;
input v_28;
input v_29;
input v_30;
input v_31;
input v_32;
input v_33;
input v_34;
input v_35;
input v_36;
input v_37;
input v_38;
input v_39;
input v_40;
input v_41;
input v_42;
input v_43;
input v_44;
input v_45;
input v_46;
input v_47;
input v_48;
input v_49;
input v_50;
input v_51;
input v_52;
input v_53;
input v_54;
input v_55;
input v_56;
input v_57;
input v_58;
input v_59;
input v_60;
input v_61;
input v_62;
input v_63;
input v_64;
input v_65;
input v_66;
input v_67;
input v_68;
input v_69;
input v_70;
input v_71;
input v_72;
input v_73;
input v_74;
input v_75;
input v_76;
input v_77;
input v_78;
input v_79;
input v_80;
input v_81;
input v_82;
input v_83;
input v_84;
input v_85;
input v_86;
input v_87;
input v_88;
input v_89;
input v_90;
input v_91;
input v_92;
input v_93;
input v_94;
input v_95;
input v_96;
input v_97;
input v_98;
input v_99;
input v_100;
input v_101;
input v_102;
input v_103;
input v_104;
input v_105;
input v_106;
input v_107;
input v_108;
input v_109;
input v_110;
input v_111;
input v_112;
input v_113;
input v_114;
input v_115;
input v_116;
input v_117;
input v_118;
input v_119;
input v_120;
input v_121;
input v_122;
input v_123;
input v_124;
input v_125;
input v_126;
input v_127;
input v_128;
input v_129;
input v_130;
input v_131;
input v_132;
input v_133;
input v_134;
input v_135;
input v_136;
input v_137;
input v_138;
input v_139;
input v_140;
input v_141;
input v_142;
input v_143;
input v_144;
input v_145;
input v_146;
input v_147;
input v_148;
input v_149;
input v_150;
input v_151;
input v_152;
input v_153;
input v_154;
input v_155;
input v_156;
input v_157;
input v_158;
input v_159;
input v_160;
input v_161;
input v_162;
input v_163;
input v_164;
input v_165;
input v_166;
input v_167;
input v_168;
input v_169;
input v_170;
input v_171;
input v_172;
input v_173;
input v_174;
input v_175;
input v_176;
input v_177;
input v_178;
input v_179;
input v_180;
input v_181;
input v_182;
input v_183;
input v_184;
input v_185;
input v_186;
input v_187;
input v_188;
input v_189;
input v_190;
input v_191;
input v_192;
input v_193;
input v_194;
input v_195;
input v_196;
input v_197;
input v_198;
input v_199;
input v_200;
input v_201;
input v_202;
input v_203;
input v_204;
input v_205;
input v_206;
input v_207;
input v_208;
input v_209;
input v_210;
input v_211;
input v_212;
input v_213;
input v_214;
input v_215;
input v_216;
input v_217;
input v_218;
input v_219;
input v_220;
input v_221;
input v_222;
input v_223;
input v_224;
input v_225;
input v_226;
input v_227;
input v_228;
input v_229;
input v_230;
input v_231;
input v_232;
input v_233;
input v_234;
input v_235;
input v_236;
input v_237;
input v_238;
input v_239;
input v_240;
input v_241;
input v_242;
input v_243;
input v_244;
input v_245;
input v_246;
input v_247;
input v_248;
input v_249;
input v_250;
input v_251;
input v_252;
input v_253;
input v_254;
input v_255;
input v_256;
input v_257;
input v_258;
input v_259;
input v_260;
input v_261;
input v_262;
input v_263;
input v_264;
input v_265;
input v_266;
input v_267;
input v_268;
input v_269;
input v_270;
input v_271;
input v_272;
input v_273;
input v_274;
input v_275;
input v_276;
input v_277;
input v_278;
input v_279;
input v_280;
input v_281;
input v_282;
input v_283;
input v_284;
input v_285;
input v_286;
input v_287;
input v_288;
input v_289;
input v_290;
input v_291;
input v_292;
input v_293;
input v_294;
input v_295;
input v_296;
input v_297;
input v_298;
input v_299;
input v_300;
input v_301;
input v_302;
input v_303;
input v_304;
input v_305;
input v_306;
input v_307;
input v_308;
input v_309;
input v_310;
input v_311;
input v_312;
input v_313;
input v_314;
input v_315;
input v_316;
input v_317;
input v_318;
input v_319;
input v_320;
input v_321;
input v_322;
input v_323;
input v_324;
input v_325;
input v_326;
input v_327;
input v_328;
input v_329;
input v_330;
input v_331;
input v_332;
input v_333;
input v_334;
input v_335;
input v_336;
input v_337;
input v_338;
input v_339;
input v_340;
input v_341;
input v_342;
input v_343;
input v_344;
input v_345;
input v_346;
input v_347;
input v_348;
input v_349;
input v_350;
input v_351;
input v_352;
input v_353;
input v_354;
input v_355;
input v_356;
input v_357;
input v_358;
input v_359;
input v_360;
input v_361;
input v_362;
input v_363;
input v_364;
input v_365;
input v_366;
input v_367;
input v_368;
input v_369;
input v_370;
input v_371;
input v_372;
input v_373;
input v_374;
input v_375;
input v_376;
input v_377;
input v_378;
input v_379;
input v_380;
input v_381;
input v_382;
input v_383;
input v_384;
input v_385;
input v_386;
input v_387;
input v_388;
input v_389;
input v_390;
input v_391;
input v_392;
input v_393;
input v_394;
input v_395;
input v_396;
input v_397;
input v_398;
input v_399;
input v_400;
input v_401;
input v_402;
input v_403;
input v_404;
input v_405;
input v_406;
input v_407;
input v_408;
input v_409;
input v_410;
input v_411;
input v_412;
input v_413;
input v_414;
input v_415;
input v_416;
input v_417;
input v_418;
input v_419;
input v_420;
input v_421;
input v_422;
input v_423;
input v_424;
input v_425;
input v_426;
input v_427;
input v_428;
input v_429;
input v_430;
input v_431;
input v_432;
input v_433;
input v_434;
input v_435;
input v_436;
input v_437;
input v_438;
input v_439;
input v_440;
input v_441;
input v_442;
input v_443;
input v_444;
input v_445;
input v_446;
input v_447;
input v_448;
input v_449;
input v_450;
input v_451;
input v_452;
input v_453;
input v_454;
input v_455;
input v_456;
input v_457;
input v_458;
input v_459;
input v_460;
input v_461;
input v_462;
input v_463;
input v_464;
input v_465;
input v_466;
input v_467;
input v_468;
input v_469;
input v_470;
input v_471;
input v_472;
input v_473;
input v_474;
input v_475;
input v_476;
input v_477;
input v_478;
input v_479;
input v_480;
input v_481;
input v_482;
input v_483;
input v_484;
input v_485;
input v_486;
input v_487;
input v_488;
input v_489;
input v_490;
input v_491;
input v_492;
input v_493;
input v_494;
input v_495;
input v_496;
input v_497;
input v_498;
input v_499;
input v_500;
input v_501;
input v_502;
input v_503;
input v_504;
input v_505;
input v_506;
input v_507;
input v_508;
input v_509;
input v_510;
input v_511;
input v_512;
input v_513;
input v_514;
input v_515;
input v_516;
input v_517;
input v_518;
input v_519;
input v_520;
input v_521;
input v_522;
input v_523;
input v_524;
input v_525;
input v_526;
input v_527;
input v_528;
input v_529;
input v_530;
input v_531;
input v_532;
input v_533;
input v_534;
input v_535;
input v_536;
input v_537;
input v_538;
input v_539;
input v_540;
input v_541;
input v_542;
input v_543;
input v_544;
input v_545;
input v_546;
input v_547;
input v_548;
input v_549;
input v_550;
input v_551;
input v_552;
input v_553;
input v_554;
input v_555;
input v_556;
input v_557;
input v_558;
input v_559;
input v_560;
input v_561;
input v_562;
input v_563;
input v_564;
input v_565;
input v_566;
input v_567;
input v_568;
input v_569;
input v_570;
input v_571;
input v_572;
input v_573;
input v_574;
input v_575;
input v_576;
input v_577;
output o_1;
wire v_578;
wire v_579;
wire v_580;
wire v_581;
wire v_582;
wire v_583;
wire v_584;
wire v_585;
wire v_586;
wire v_587;
wire v_588;
wire v_589;
wire v_590;
wire v_591;
wire v_592;
wire v_593;
wire v_594;
wire v_595;
wire v_596;
wire v_597;
wire v_598;
wire v_599;
wire v_600;
wire v_601;
wire v_602;
wire v_603;
wire v_604;
wire v_605;
wire v_606;
wire v_607;
wire v_608;
wire v_609;
wire v_610;
wire v_611;
wire v_612;
wire v_613;
wire v_614;
wire v_615;
wire v_616;
wire v_617;
wire v_618;
wire v_619;
wire v_620;
wire v_621;
wire v_622;
wire v_623;
wire v_624;
wire v_625;
wire v_626;
wire v_627;
wire v_628;
wire v_629;
wire v_630;
wire v_631;
wire v_632;
wire v_633;
wire v_634;
wire v_635;
wire v_636;
wire v_637;
wire v_638;
wire v_639;
wire v_640;
wire v_641;
wire v_642;
wire v_643;
wire v_644;
wire v_645;
wire v_646;
wire v_647;
wire v_648;
wire v_649;
wire v_650;
wire v_651;
wire v_652;
wire v_653;
wire v_654;
wire v_655;
wire v_656;
wire v_657;
wire v_658;
wire v_659;
wire v_660;
wire v_661;
wire v_662;
wire v_663;
wire v_664;
wire v_665;
wire v_666;
wire v_667;
wire v_668;
wire v_669;
wire v_670;
wire v_671;
wire v_672;
wire v_673;
wire v_674;
wire v_675;
wire v_676;
wire v_677;
wire v_678;
wire v_679;
wire v_680;
wire v_681;
wire v_682;
wire v_683;
wire v_684;
wire v_685;
wire v_686;
wire v_687;
wire v_688;
wire v_689;
wire v_690;
wire v_691;
wire v_692;
wire v_693;
wire v_694;
wire v_695;
wire v_696;
wire v_697;
wire v_698;
wire v_699;
wire v_700;
wire v_701;
wire v_702;
wire v_703;
wire v_704;
wire v_705;
wire v_706;
wire v_707;
wire v_708;
wire v_709;
wire v_710;
wire v_711;
wire v_712;
wire v_713;
wire v_714;
wire v_715;
wire v_716;
wire v_717;
wire v_718;
wire v_719;
wire v_720;
wire v_721;
wire v_722;
wire v_723;
wire v_724;
wire v_725;
wire v_726;
wire v_727;
wire v_728;
wire v_729;
wire v_730;
wire v_731;
wire v_732;
wire v_733;
wire v_734;
wire v_735;
wire v_736;
wire v_737;
wire v_738;
wire v_739;
wire v_740;
wire v_741;
wire v_742;
wire v_743;
wire v_744;
wire v_745;
wire v_746;
wire v_747;
wire v_748;
wire v_749;
wire v_750;
wire v_751;
wire v_752;
wire v_753;
wire v_754;
wire v_755;
wire v_756;
wire v_757;
wire v_758;
wire v_759;
wire v_760;
wire v_761;
wire v_762;
wire v_763;
wire v_764;
wire v_765;
wire v_766;
wire v_767;
wire v_768;
wire v_769;
wire v_770;
wire v_771;
wire v_772;
wire v_773;
wire v_774;
wire v_775;
wire v_776;
wire v_777;
wire v_778;
wire v_779;
wire v_780;
wire v_781;
wire v_782;
wire v_783;
wire v_784;
wire v_785;
wire v_786;
wire v_787;
wire v_788;
wire v_789;
wire v_790;
wire v_791;
wire v_792;
wire v_793;
wire v_794;
wire v_795;
wire v_796;
wire v_797;
wire v_798;
wire v_799;
wire v_800;
wire v_801;
wire v_802;
wire v_803;
wire v_804;
wire v_805;
wire v_806;
wire v_807;
wire v_808;
wire v_809;
wire v_810;
wire v_811;
wire v_812;
wire v_813;
wire v_814;
wire v_815;
wire v_816;
wire v_817;
wire v_818;
wire v_819;
wire v_820;
wire v_821;
wire v_822;
wire v_823;
wire v_824;
wire v_825;
wire v_826;
wire v_827;
wire v_828;
wire v_829;
wire v_830;
wire v_831;
wire v_832;
wire v_833;
wire v_834;
wire v_835;
wire v_836;
wire v_837;
wire v_838;
wire v_839;
wire v_840;
wire v_841;
wire v_842;
wire v_843;
wire v_844;
wire v_845;
wire v_846;
wire v_847;
wire v_848;
wire v_849;
wire v_850;
wire v_851;
wire v_852;
wire v_853;
wire v_854;
wire v_855;
wire v_856;
wire v_857;
wire v_858;
wire v_859;
wire v_860;
wire v_861;
wire v_862;
wire v_863;
wire v_864;
wire v_865;
wire v_866;
wire v_867;
wire v_868;
wire v_869;
wire v_870;
wire v_871;
wire v_872;
wire v_873;
wire v_874;
wire v_875;
wire v_876;
wire v_877;
wire v_878;
wire v_879;
wire v_880;
wire v_881;
wire v_882;
wire v_883;
wire v_884;
wire v_885;
wire v_886;
wire v_887;
wire v_888;
wire v_889;
wire v_890;
wire v_891;
wire v_892;
wire v_893;
wire v_894;
wire v_895;
wire v_896;
wire v_897;
wire v_898;
wire v_899;
wire v_900;
wire v_901;
wire v_902;
wire v_903;
wire v_904;
wire v_905;
wire v_906;
wire v_907;
wire v_908;
wire v_909;
wire v_910;
wire v_911;
wire v_912;
wire v_913;
wire v_914;
wire v_915;
wire v_916;
wire v_917;
wire v_918;
wire v_919;
wire v_920;
wire v_921;
wire v_922;
wire v_923;
wire v_924;
wire v_925;
wire v_926;
wire v_927;
wire v_928;
wire v_929;
wire v_930;
wire v_931;
wire v_932;
wire v_933;
wire v_934;
wire v_935;
wire v_936;
wire v_937;
wire v_938;
wire v_939;
wire v_940;
wire v_941;
wire v_942;
wire v_943;
wire v_944;
wire v_945;
wire v_946;
wire v_947;
wire v_948;
wire v_949;
wire v_950;
wire v_951;
wire v_952;
wire v_953;
wire v_954;
wire v_955;
wire v_956;
wire v_957;
wire v_958;
wire v_959;
wire v_960;
wire v_961;
wire v_962;
wire v_963;
wire v_964;
wire v_965;
wire v_966;
wire v_967;
wire v_968;
wire v_969;
wire v_970;
wire v_971;
wire v_972;
wire v_973;
wire v_974;
wire v_975;
wire v_976;
wire v_977;
wire v_978;
wire v_979;
wire v_980;
wire v_981;
wire v_982;
wire v_983;
wire v_984;
wire v_985;
wire v_986;
wire v_987;
wire v_988;
wire v_989;
wire v_990;
wire v_991;
wire v_992;
wire v_993;
wire v_994;
wire v_995;
wire v_996;
wire v_997;
wire v_998;
wire v_999;
wire v_1000;
wire v_1001;
wire v_1002;
wire v_1003;
wire v_1004;
wire v_1005;
wire v_1006;
wire v_1007;
wire v_1008;
wire v_1009;
wire v_1010;
wire v_1011;
wire v_1012;
wire v_1013;
wire v_1014;
wire v_1015;
wire v_1016;
wire v_1017;
wire v_1018;
wire v_1019;
wire v_1020;
wire v_1021;
wire v_1022;
wire v_1023;
wire v_1024;
wire v_1025;
wire v_1026;
wire v_1027;
wire v_1028;
wire v_1029;
wire v_1030;
wire v_1031;
wire v_1032;
wire v_1033;
wire v_1034;
wire v_1035;
wire v_1036;
wire v_1037;
wire v_1038;
wire v_1039;
wire v_1040;
wire v_1041;
wire v_1042;
wire v_1043;
wire v_1044;
wire v_1045;
wire v_1046;
wire v_1047;
wire v_1048;
wire v_1049;
wire v_1050;
wire v_1051;
wire v_1052;
wire v_1053;
wire v_1054;
wire v_1055;
wire v_1056;
wire v_1057;
wire v_1058;
wire v_1059;
wire v_1060;
wire v_1061;
wire v_1062;
wire v_1063;
wire v_1064;
wire v_1065;
wire v_1066;
wire v_1067;
wire v_1068;
wire v_1069;
wire v_1070;
wire v_1071;
wire v_1072;
wire v_1073;
wire v_1074;
wire v_1075;
wire v_1076;
wire v_1077;
wire v_1078;
wire v_1079;
wire v_1080;
wire v_1081;
wire v_1082;
wire v_1083;
wire v_1084;
wire v_1085;
wire v_1086;
wire v_1087;
wire v_1088;
wire v_1089;
wire v_1090;
wire v_1091;
wire v_1092;
wire v_1093;
wire v_1094;
wire v_1095;
wire v_1096;
wire v_1097;
wire v_1098;
wire v_1099;
wire v_1100;
wire v_1101;
wire v_1102;
wire v_1103;
wire v_1104;
wire v_1105;
wire v_1106;
wire v_1107;
wire v_1108;
wire v_1109;
wire v_1110;
wire v_1111;
wire v_1112;
wire v_1113;
wire v_1114;
wire v_1115;
wire v_1116;
wire v_1117;
wire v_1118;
wire v_1119;
wire v_1120;
wire v_1121;
wire v_1122;
wire v_1123;
wire v_1124;
wire v_1125;
wire v_1126;
wire v_1127;
wire v_1128;
wire v_1129;
wire v_1130;
wire v_1131;
wire v_1132;
wire v_1133;
wire v_1134;
wire v_1135;
wire v_1136;
wire v_1137;
wire v_1138;
wire v_1139;
wire v_1140;
wire v_1141;
wire v_1142;
wire v_1143;
wire v_1144;
wire v_1145;
wire v_1146;
wire v_1147;
wire v_1148;
wire v_1149;
wire v_1150;
wire v_1151;
wire v_1152;
wire v_1153;
wire v_1154;
wire v_1155;
wire v_1156;
wire v_1157;
wire v_1158;
wire v_1159;
wire v_1160;
wire v_1161;
wire v_1162;
wire v_1163;
wire v_1164;
wire v_1165;
wire v_1166;
wire v_1167;
wire v_1168;
wire v_1169;
wire v_1170;
wire v_1171;
wire v_1172;
wire v_1173;
wire v_1174;
wire v_1175;
wire v_1176;
wire v_1177;
wire v_1178;
wire v_1179;
wire v_1180;
wire v_1181;
wire v_1182;
wire v_1183;
wire v_1184;
wire v_1185;
wire v_1186;
wire v_1187;
wire v_1188;
wire v_1189;
wire v_1190;
wire v_1191;
wire v_1192;
wire v_1193;
wire v_1194;
wire v_1195;
wire v_1196;
wire v_1197;
wire v_1198;
wire v_1199;
wire v_1200;
wire v_1201;
wire v_1202;
wire v_1203;
wire v_1204;
wire v_1205;
wire v_1206;
wire v_1207;
wire v_1208;
wire v_1209;
wire v_1210;
wire v_1211;
wire v_1212;
wire v_1213;
wire v_1214;
wire v_1215;
wire v_1216;
wire v_1217;
wire v_1218;
wire v_1219;
wire v_1220;
wire v_1221;
wire v_1222;
wire v_1223;
wire v_1224;
wire v_1225;
wire v_1226;
wire v_1227;
wire v_1228;
wire v_1229;
wire v_1230;
wire v_1231;
wire v_1232;
wire v_1233;
wire v_1234;
wire v_1235;
wire v_1236;
wire v_1237;
wire v_1238;
wire v_1239;
wire v_1240;
wire v_1241;
wire v_1242;
wire v_1243;
wire v_1244;
wire v_1245;
wire v_1246;
wire v_1247;
wire v_1248;
wire v_1249;
wire v_1250;
wire v_1251;
wire v_1252;
wire v_1253;
wire v_1254;
wire v_1255;
wire v_1256;
wire v_1257;
wire v_1258;
wire v_1259;
wire v_1260;
wire v_1261;
wire v_1262;
wire v_1263;
wire v_1264;
wire v_1265;
wire v_1266;
wire v_1267;
wire v_1268;
wire v_1269;
wire v_1270;
wire v_1271;
wire v_1272;
wire v_1273;
wire v_1274;
wire v_1275;
wire v_1276;
wire v_1277;
wire v_1278;
wire v_1279;
wire v_1280;
wire v_1281;
wire v_1282;
wire v_1283;
wire v_1284;
wire v_1285;
wire v_1286;
wire v_1287;
wire v_1288;
wire v_1289;
wire v_1290;
wire v_1291;
wire v_1292;
wire v_1293;
wire v_1294;
wire v_1295;
wire v_1296;
wire v_1297;
wire v_1298;
wire v_1299;
wire v_1300;
wire v_1301;
wire v_1302;
wire v_1303;
wire v_1304;
wire v_1305;
wire v_1306;
wire v_1307;
wire v_1308;
wire v_1309;
wire v_1310;
wire v_1311;
wire v_1312;
wire v_1313;
wire v_1314;
wire v_1315;
wire v_1316;
wire v_1317;
wire v_1318;
wire v_1319;
wire v_1320;
wire v_1321;
wire v_1322;
wire v_1323;
wire v_1324;
wire v_1325;
wire v_1326;
wire v_1327;
wire v_1328;
wire v_1329;
wire v_1330;
wire v_1331;
wire v_1332;
wire v_1333;
wire v_1334;
wire v_1335;
wire v_1336;
wire v_1337;
wire v_1338;
wire v_1339;
wire v_1340;
wire v_1341;
wire v_1342;
wire v_1343;
wire v_1344;
wire v_1345;
wire v_1346;
wire v_1347;
wire v_1348;
wire v_1349;
wire v_1350;
wire v_1351;
wire v_1352;
wire v_1353;
wire v_1354;
wire v_1355;
wire v_1356;
wire v_1357;
wire v_1358;
wire v_1359;
wire v_1360;
wire v_1361;
wire v_1362;
wire v_1363;
wire v_1364;
wire v_1365;
wire v_1366;
wire v_1367;
wire v_1368;
wire v_1369;
wire v_1370;
wire v_1371;
wire v_1372;
wire v_1373;
wire v_1374;
wire v_1375;
wire v_1376;
wire v_1377;
wire v_1378;
wire v_1379;
wire v_1380;
wire v_1381;
wire v_1382;
wire v_1383;
wire v_1384;
wire v_1385;
wire v_1386;
wire v_1387;
wire v_1388;
wire v_1389;
wire v_1390;
wire v_1391;
wire v_1392;
wire v_1393;
wire v_1394;
wire v_1395;
wire v_1396;
wire v_1397;
wire v_1398;
wire v_1399;
wire v_1400;
wire v_1401;
wire v_1402;
wire v_1403;
wire v_1404;
wire v_1405;
wire v_1406;
wire v_1407;
wire v_1408;
wire v_1409;
wire v_1410;
wire v_1411;
wire v_1412;
wire v_1413;
wire v_1414;
wire v_1415;
wire v_1416;
wire v_1417;
wire v_1418;
wire v_1419;
wire v_1420;
wire v_1421;
wire v_1422;
wire v_1423;
wire v_1424;
wire v_1425;
wire v_1426;
wire v_1427;
wire v_1428;
wire v_1429;
wire v_1430;
wire v_1431;
wire v_1432;
wire v_1433;
wire v_1434;
wire v_1435;
wire v_1436;
wire v_1437;
wire v_1438;
wire v_1439;
wire v_1440;
wire v_1441;
wire v_1442;
wire v_1443;
wire v_1444;
wire v_1445;
wire v_1446;
wire v_1447;
wire v_1448;
wire v_1449;
wire v_1450;
wire v_1451;
wire v_1452;
wire v_1453;
wire v_1454;
wire v_1455;
wire v_1456;
wire v_1457;
wire v_1458;
wire v_1459;
wire v_1460;
wire v_1461;
wire v_1462;
wire v_1463;
wire v_1464;
wire v_1465;
wire v_1466;
wire v_1467;
wire v_1468;
wire v_1469;
wire v_1470;
wire v_1471;
wire v_1472;
wire v_1473;
wire v_1474;
wire v_1475;
wire v_1476;
wire v_1477;
wire v_1478;
wire v_1479;
wire v_1480;
wire v_1481;
wire v_1482;
wire v_1483;
wire v_1484;
wire v_1485;
wire v_1486;
wire v_1487;
wire v_1488;
wire v_1489;
wire v_1490;
wire v_1491;
wire v_1492;
wire v_1493;
wire v_1494;
wire v_1495;
wire v_1496;
wire v_1497;
wire v_1498;
wire v_1499;
wire v_1500;
wire v_1501;
wire v_1502;
wire v_1503;
wire v_1504;
wire v_1505;
wire v_1506;
wire v_1507;
wire v_1508;
wire v_1509;
wire v_1510;
wire v_1511;
wire v_1512;
wire v_1513;
wire v_1514;
wire v_1515;
wire v_1516;
wire v_1517;
wire v_1518;
wire v_1519;
wire v_1520;
wire v_1521;
wire v_1522;
wire v_1523;
wire v_1524;
wire v_1525;
wire v_1526;
wire v_1527;
wire v_1528;
wire v_1529;
wire v_1530;
wire v_1531;
wire v_1532;
wire v_1533;
wire v_1534;
wire v_1535;
wire v_1536;
wire v_1537;
wire v_1538;
wire v_1539;
wire v_1540;
wire v_1541;
wire v_1542;
wire v_1543;
wire v_1544;
wire v_1545;
wire x_1;
assign v_578 = v_1373 & v_1374;
assign v_579 = v_1382 & v_1383;
assign v_580 = v_1391 & v_1392;
assign v_581 = v_1400 & v_1401;
assign v_582 = v_1409 & v_1410;
assign v_583 = v_578 & v_579 & v_580 & v_581 & v_582;
assign v_585 = v_65 & v_33;
assign v_586 = v_585;
assign v_589 = v_66 & v_34;
assign v_590 = v_66 & v_586;
assign v_591 = v_34 & v_586;
assign v_595 = v_67 & v_35;
assign v_596 = v_67 & v_592;
assign v_597 = v_35 & v_592;
assign v_601 = v_68 & v_36;
assign v_602 = v_68 & v_598;
assign v_603 = v_36 & v_598;
assign v_607 = v_69 & v_37;
assign v_608 = v_69 & v_604;
assign v_609 = v_37 & v_604;
assign v_613 = v_70 & v_38;
assign v_614 = v_70 & v_610;
assign v_615 = v_38 & v_610;
assign v_619 = v_71 & v_39;
assign v_620 = v_71 & v_616;
assign v_621 = v_39 & v_616;
assign v_625 = v_72 & v_40;
assign v_626 = v_72 & v_622;
assign v_627 = v_40 & v_622;
assign v_631 = v_73 & v_41;
assign v_632 = v_73 & v_628;
assign v_633 = v_41 & v_628;
assign v_637 = v_74 & v_42;
assign v_638 = v_74 & v_634;
assign v_639 = v_42 & v_634;
assign v_643 = v_75 & v_43;
assign v_644 = v_75 & v_640;
assign v_645 = v_43 & v_640;
assign v_649 = v_76 & v_44;
assign v_650 = v_76 & v_646;
assign v_651 = v_44 & v_646;
assign v_655 = v_77 & v_45;
assign v_656 = v_77 & v_652;
assign v_657 = v_45 & v_652;
assign v_661 = v_78 & v_46;
assign v_662 = v_78 & v_658;
assign v_663 = v_46 & v_658;
assign v_667 = v_79 & v_47;
assign v_668 = v_79 & v_664;
assign v_669 = v_47 & v_664;
assign v_673 = v_80 & v_48;
assign v_674 = v_80 & v_670;
assign v_675 = v_48 & v_670;
assign v_679 = v_81 & v_49;
assign v_680 = v_81 & v_676;
assign v_681 = v_49 & v_676;
assign v_685 = v_82 & v_50;
assign v_686 = v_82 & v_682;
assign v_687 = v_50 & v_682;
assign v_691 = v_83 & v_51;
assign v_692 = v_83 & v_688;
assign v_693 = v_51 & v_688;
assign v_697 = v_84 & v_52;
assign v_698 = v_84 & v_694;
assign v_699 = v_52 & v_694;
assign v_703 = v_85 & v_53;
assign v_704 = v_85 & v_700;
assign v_705 = v_53 & v_700;
assign v_709 = v_86 & v_54;
assign v_710 = v_86 & v_706;
assign v_711 = v_54 & v_706;
assign v_715 = v_87 & v_55;
assign v_716 = v_87 & v_712;
assign v_717 = v_55 & v_712;
assign v_721 = v_88 & v_56;
assign v_722 = v_88 & v_718;
assign v_723 = v_56 & v_718;
assign v_727 = v_89 & v_57;
assign v_728 = v_89 & v_724;
assign v_729 = v_57 & v_724;
assign v_733 = v_90 & v_58;
assign v_734 = v_90 & v_730;
assign v_735 = v_58 & v_730;
assign v_739 = v_91 & v_59;
assign v_740 = v_91 & v_736;
assign v_741 = v_59 & v_736;
assign v_745 = v_92 & v_60;
assign v_746 = v_92 & v_742;
assign v_747 = v_60 & v_742;
assign v_751 = v_93 & v_61;
assign v_752 = v_93 & v_748;
assign v_753 = v_61 & v_748;
assign v_757 = v_94 & v_62;
assign v_758 = v_94 & v_754;
assign v_759 = v_62 & v_754;
assign v_763 = v_95 & v_63;
assign v_764 = v_95 & v_760;
assign v_765 = v_63 & v_760;
assign v_769 = v_96 & v_64;
assign v_770 = v_96 & v_766;
assign v_771 = v_64 & v_766;
assign v_773 = ~v_193 & v_584;
assign v_774 = ~v_193 & v_588;
assign v_775 = ~v_193 & v_594;
assign v_776 = ~v_193 & v_600;
assign v_777 = ~v_193 & v_606;
assign v_778 = ~v_193 & v_612;
assign v_779 = ~v_193 & v_618;
assign v_780 = ~v_193 & v_624;
assign v_781 = ~v_193 & v_630;
assign v_782 = ~v_193 & v_636;
assign v_783 = ~v_193 & v_642;
assign v_784 = ~v_193 & v_648;
assign v_785 = ~v_193 & v_654;
assign v_786 = ~v_193 & v_660;
assign v_787 = ~v_193 & v_666;
assign v_788 = ~v_193 & v_672;
assign v_789 = ~v_193 & v_678;
assign v_790 = ~v_193 & v_684;
assign v_791 = ~v_193 & v_690;
assign v_792 = ~v_193 & v_696;
assign v_793 = ~v_193 & v_702;
assign v_794 = ~v_193 & v_708;
assign v_795 = ~v_193 & v_714;
assign v_796 = ~v_193 & v_720;
assign v_797 = ~v_193 & v_726;
assign v_798 = ~v_193 & v_732;
assign v_799 = ~v_193 & v_738;
assign v_800 = ~v_193 & v_744;
assign v_801 = ~v_193 & v_750;
assign v_802 = ~v_193 & v_756;
assign v_803 = ~v_193 & v_762;
assign v_804 = ~v_193 & v_768;
assign v_837 = v_1418 & v_1419;
assign v_839 = v_226 & v_258;
assign v_840 = v_839;
assign v_843 = v_227 & v_259;
assign v_844 = v_227 & v_840;
assign v_845 = v_259 & v_840;
assign v_849 = v_228 & v_260;
assign v_850 = v_228 & v_846;
assign v_851 = v_260 & v_846;
assign v_855 = v_229 & v_261;
assign v_856 = v_229 & v_852;
assign v_857 = v_261 & v_852;
assign v_861 = v_230 & v_262;
assign v_862 = v_230 & v_858;
assign v_863 = v_262 & v_858;
assign v_867 = v_231 & v_263;
assign v_868 = v_231 & v_864;
assign v_869 = v_263 & v_864;
assign v_873 = v_232 & v_264;
assign v_874 = v_232 & v_870;
assign v_875 = v_264 & v_870;
assign v_879 = v_233 & v_265;
assign v_880 = v_233 & v_876;
assign v_881 = v_265 & v_876;
assign v_885 = v_234 & v_266;
assign v_886 = v_234 & v_882;
assign v_887 = v_266 & v_882;
assign v_891 = v_235 & v_267;
assign v_892 = v_235 & v_888;
assign v_893 = v_267 & v_888;
assign v_897 = v_236 & v_268;
assign v_898 = v_236 & v_894;
assign v_899 = v_268 & v_894;
assign v_903 = v_237 & v_269;
assign v_904 = v_237 & v_900;
assign v_905 = v_269 & v_900;
assign v_909 = v_238 & v_270;
assign v_910 = v_238 & v_906;
assign v_911 = v_270 & v_906;
assign v_915 = v_239 & v_271;
assign v_916 = v_239 & v_912;
assign v_917 = v_271 & v_912;
assign v_921 = v_240 & v_272;
assign v_922 = v_240 & v_918;
assign v_923 = v_272 & v_918;
assign v_927 = v_241 & v_273;
assign v_928 = v_241 & v_924;
assign v_929 = v_273 & v_924;
assign v_933 = v_242 & v_274;
assign v_934 = v_242 & v_930;
assign v_935 = v_274 & v_930;
assign v_939 = v_243 & v_275;
assign v_940 = v_243 & v_936;
assign v_941 = v_275 & v_936;
assign v_945 = v_244 & v_276;
assign v_946 = v_244 & v_942;
assign v_947 = v_276 & v_942;
assign v_951 = v_245 & v_277;
assign v_952 = v_245 & v_948;
assign v_953 = v_277 & v_948;
assign v_957 = v_246 & v_278;
assign v_958 = v_246 & v_954;
assign v_959 = v_278 & v_954;
assign v_963 = v_247 & v_279;
assign v_964 = v_247 & v_960;
assign v_965 = v_279 & v_960;
assign v_969 = v_248 & v_280;
assign v_970 = v_248 & v_966;
assign v_971 = v_280 & v_966;
assign v_975 = v_249 & v_281;
assign v_976 = v_249 & v_972;
assign v_977 = v_281 & v_972;
assign v_981 = v_250 & v_282;
assign v_982 = v_250 & v_978;
assign v_983 = v_282 & v_978;
assign v_987 = v_251 & v_283;
assign v_988 = v_251 & v_984;
assign v_989 = v_283 & v_984;
assign v_993 = v_252 & v_284;
assign v_994 = v_252 & v_990;
assign v_995 = v_284 & v_990;
assign v_999 = v_253 & v_285;
assign v_1000 = v_253 & v_996;
assign v_1001 = v_285 & v_996;
assign v_1005 = v_254 & v_286;
assign v_1006 = v_254 & v_1002;
assign v_1007 = v_286 & v_1002;
assign v_1011 = v_255 & v_287;
assign v_1012 = v_255 & v_1008;
assign v_1013 = v_287 & v_1008;
assign v_1017 = v_256 & v_288;
assign v_1018 = v_256 & v_1014;
assign v_1019 = v_288 & v_1014;
assign v_1023 = v_257 & v_289;
assign v_1024 = v_257 & v_1020;
assign v_1025 = v_289 & v_1020;
assign v_1059 = v_1427 & v_1428;
assign v_1060 = v_33 & v_322;
assign v_1061 = v_34 & v_323;
assign v_1062 = v_35 & v_324;
assign v_1063 = v_36 & v_325;
assign v_1064 = v_37 & v_326;
assign v_1065 = v_38 & v_327;
assign v_1066 = v_39 & v_328;
assign v_1067 = v_40 & v_329;
assign v_1068 = v_41 & v_330;
assign v_1069 = v_42 & v_331;
assign v_1070 = v_43 & v_332;
assign v_1071 = v_44 & v_333;
assign v_1072 = v_45 & v_334;
assign v_1073 = v_46 & v_335;
assign v_1074 = v_47 & v_336;
assign v_1075 = v_48 & v_337;
assign v_1076 = v_49 & v_338;
assign v_1077 = v_50 & v_339;
assign v_1078 = v_51 & v_340;
assign v_1079 = v_52 & v_341;
assign v_1080 = v_53 & v_342;
assign v_1081 = v_54 & v_343;
assign v_1082 = v_55 & v_344;
assign v_1083 = v_56 & v_345;
assign v_1084 = v_57 & v_346;
assign v_1085 = v_58 & v_347;
assign v_1086 = v_59 & v_348;
assign v_1087 = v_60 & v_349;
assign v_1088 = v_61 & v_350;
assign v_1089 = v_62 & v_351;
assign v_1090 = v_63 & v_352;
assign v_1091 = v_64 & v_353;
assign v_1124 = v_1436 & v_1437;
assign v_1157 = v_1445 & v_1446;
assign v_1190 = v_1454 & v_1455;
assign v_1191 = v_837 & v_1059 & v_1124 & v_1157 & v_1190;
assign v_1192 = v_583 & v_1191;
assign v_1193 = v_1463 & v_1464;
assign v_1194 = v_1472 & v_1473;
assign v_1195 = v_1481 & v_1482;
assign v_1196 = v_1490 & v_1491;
assign v_1197 = v_1499 & v_1500;
assign v_1198 = v_1193 & v_1194 & v_1195 & v_1196 & v_1197;
assign v_1231 = v_1508 & v_1509;
assign v_1264 = v_1517 & v_1518;
assign v_1297 = v_1526 & v_1527;
assign v_1330 = v_1535 & v_1536;
assign v_1363 = v_1544 & v_1545;
assign v_1364 = v_1231 & v_1264 & v_1297 & v_1330 & v_1363;
assign v_1365 = v_1198 & v_1364;
assign v_1366 = ~v_1 & ~v_2 & ~v_3 & ~v_4 & ~v_5;
assign v_1367 = ~v_6 & ~v_7 & ~v_8 & ~v_9 & ~v_10;
assign v_1368 = ~v_11 & ~v_12 & ~v_13 & ~v_14 & ~v_15;
assign v_1369 = ~v_16 & ~v_17 & ~v_18 & ~v_19 & ~v_20;
assign v_1370 = ~v_21 & ~v_22 & ~v_23 & ~v_24 & ~v_25;
assign v_1371 = ~v_26 & ~v_27 & ~v_28 & ~v_29 & ~v_30;
assign v_1372 = ~v_31 & ~v_32;
assign v_1373 = v_1366 & v_1367 & v_1368 & v_1369 & v_1370;
assign v_1374 = v_1371 & v_1372;
assign v_1375 = ~v_33 & ~v_34 & ~v_35 & ~v_36 & ~v_37;
assign v_1376 = ~v_38 & ~v_39 & ~v_40 & ~v_41 & ~v_42;
assign v_1377 = ~v_43 & ~v_44 & ~v_45 & ~v_46 & ~v_47;
assign v_1378 = ~v_48 & ~v_49 & ~v_50 & ~v_51 & ~v_52;
assign v_1379 = ~v_53 & ~v_54 & ~v_55 & ~v_56 & ~v_57;
assign v_1380 = ~v_58 & ~v_59 & ~v_60 & ~v_61 & ~v_62;
assign v_1381 = ~v_63 & ~v_64;
assign v_1382 = v_1375 & v_1376 & v_1377 & v_1378 & v_1379;
assign v_1383 = v_1380 & v_1381;
assign v_1384 = ~v_65 & ~v_66 & ~v_67 & ~v_68 & ~v_69;
assign v_1385 = ~v_70 & ~v_71 & ~v_72 & ~v_73 & ~v_74;
assign v_1386 = ~v_75 & ~v_76 & ~v_77 & ~v_78 & ~v_79;
assign v_1387 = ~v_80 & ~v_81 & ~v_82 & ~v_83 & ~v_84;
assign v_1388 = ~v_85 & ~v_86 & ~v_87 & ~v_88 & ~v_89;
assign v_1389 = ~v_90 & ~v_91 & ~v_92 & ~v_93 & ~v_94;
assign v_1390 = ~v_95 & ~v_96;
assign v_1391 = v_1384 & v_1385 & v_1386 & v_1387 & v_1388;
assign v_1392 = v_1389 & v_1390;
assign v_1393 = ~v_97 & ~v_98 & ~v_99 & ~v_100 & ~v_101;
assign v_1394 = ~v_102 & ~v_103 & ~v_104 & ~v_105 & ~v_106;
assign v_1395 = ~v_107 & ~v_108 & ~v_109 & ~v_110 & ~v_111;
assign v_1396 = ~v_112 & ~v_113 & ~v_114 & ~v_115 & ~v_116;
assign v_1397 = ~v_117 & ~v_118 & ~v_119 & ~v_120 & ~v_121;
assign v_1398 = ~v_122 & ~v_123 & ~v_124 & ~v_125 & ~v_126;
assign v_1399 = ~v_127 & ~v_128;
assign v_1400 = v_1393 & v_1394 & v_1395 & v_1396 & v_1397;
assign v_1401 = v_1398 & v_1399;
assign v_1402 = ~v_129 & ~v_130 & ~v_131 & ~v_132 & ~v_133;
assign v_1403 = ~v_134 & ~v_135 & ~v_136 & ~v_137 & ~v_138;
assign v_1404 = ~v_139 & ~v_140 & ~v_141 & ~v_142 & ~v_143;
assign v_1405 = ~v_144 & ~v_145 & ~v_146 & ~v_147 & ~v_148;
assign v_1406 = ~v_149 & ~v_150 & ~v_151 & ~v_152 & ~v_153;
assign v_1407 = ~v_154 & ~v_155 & ~v_156 & ~v_157 & ~v_158;
assign v_1408 = ~v_159 & ~v_160;
assign v_1409 = v_1402 & v_1403 & v_1404 & v_1405 & v_1406;
assign v_1410 = v_1407 & v_1408;
assign v_1411 = ~v_805 & ~v_806 & ~v_807 & ~v_808 & ~v_809;
assign v_1412 = ~v_810 & ~v_811 & ~v_812 & ~v_813 & ~v_814;
assign v_1413 = ~v_815 & ~v_816 & ~v_817 & ~v_818 & ~v_819;
assign v_1414 = ~v_820 & ~v_821 & ~v_822 & ~v_823 & ~v_824;
assign v_1415 = ~v_825 & ~v_826 & ~v_827 & ~v_828 & ~v_829;
assign v_1416 = ~v_830 & ~v_831 & ~v_832 & ~v_833 & ~v_834;
assign v_1417 = ~v_835 & ~v_836;
assign v_1418 = v_1411 & v_1412 & v_1413 & v_1414 & v_1415;
assign v_1419 = v_1416 & v_1417;
assign v_1420 = ~v_1027 & ~v_1028 & ~v_1029 & ~v_1030 & ~v_1031;
assign v_1421 = ~v_1032 & ~v_1033 & ~v_1034 & ~v_1035 & ~v_1036;
assign v_1422 = ~v_1037 & ~v_1038 & ~v_1039 & ~v_1040 & ~v_1041;
assign v_1423 = ~v_1042 & ~v_1043 & ~v_1044 & ~v_1045 & ~v_1046;
assign v_1424 = ~v_1047 & ~v_1048 & ~v_1049 & ~v_1050 & ~v_1051;
assign v_1425 = ~v_1052 & ~v_1053 & ~v_1054 & ~v_1055 & ~v_1056;
assign v_1426 = ~v_1057 & ~v_1058;
assign v_1427 = v_1420 & v_1421 & v_1422 & v_1423 & v_1424;
assign v_1428 = v_1425 & v_1426;
assign v_1429 = ~v_1092 & ~v_1093 & ~v_1094 & ~v_1095 & ~v_1096;
assign v_1430 = ~v_1097 & ~v_1098 & ~v_1099 & ~v_1100 & ~v_1101;
assign v_1431 = ~v_1102 & ~v_1103 & ~v_1104 & ~v_1105 & ~v_1106;
assign v_1432 = ~v_1107 & ~v_1108 & ~v_1109 & ~v_1110 & ~v_1111;
assign v_1433 = ~v_1112 & ~v_1113 & ~v_1114 & ~v_1115 & ~v_1116;
assign v_1434 = ~v_1117 & ~v_1118 & ~v_1119 & ~v_1120 & ~v_1121;
assign v_1435 = ~v_1122 & ~v_1123;
assign v_1436 = v_1429 & v_1430 & v_1431 & v_1432 & v_1433;
assign v_1437 = v_1434 & v_1435;
assign v_1438 = ~v_1125 & ~v_1126 & ~v_1127 & ~v_1128 & ~v_1129;
assign v_1439 = ~v_1130 & ~v_1131 & ~v_1132 & ~v_1133 & ~v_1134;
assign v_1440 = ~v_1135 & ~v_1136 & ~v_1137 & ~v_1138 & ~v_1139;
assign v_1441 = ~v_1140 & ~v_1141 & ~v_1142 & ~v_1143 & ~v_1144;
assign v_1442 = ~v_1145 & ~v_1146 & ~v_1147 & ~v_1148 & ~v_1149;
assign v_1443 = ~v_1150 & ~v_1151 & ~v_1152 & ~v_1153 & ~v_1154;
assign v_1444 = ~v_1155 & ~v_1156;
assign v_1445 = v_1438 & v_1439 & v_1440 & v_1441 & v_1442;
assign v_1446 = v_1443 & v_1444;
assign v_1447 = ~v_1158 & ~v_1159 & ~v_1160 & ~v_1161 & ~v_1162;
assign v_1448 = ~v_1163 & ~v_1164 & ~v_1165 & ~v_1166 & ~v_1167;
assign v_1449 = ~v_1168 & ~v_1169 & ~v_1170 & ~v_1171 & ~v_1172;
assign v_1450 = ~v_1173 & ~v_1174 & ~v_1175 & ~v_1176 & ~v_1177;
assign v_1451 = ~v_1178 & ~v_1179 & ~v_1180 & ~v_1181 & ~v_1182;
assign v_1452 = ~v_1183 & ~v_1184 & ~v_1185 & ~v_1186 & ~v_1187;
assign v_1453 = ~v_1188 & ~v_1189;
assign v_1454 = v_1447 & v_1448 & v_1449 & v_1450 & v_1451;
assign v_1455 = v_1452 & v_1453;
assign v_1456 = ~v_418 & ~v_419 & ~v_420 & ~v_421 & ~v_422;
assign v_1457 = ~v_423 & ~v_424 & ~v_425 & ~v_426 & ~v_427;
assign v_1458 = ~v_428 & ~v_429 & ~v_430 & ~v_431 & ~v_432;
assign v_1459 = ~v_433 & ~v_434 & ~v_435 & ~v_436 & ~v_437;
assign v_1460 = ~v_438 & ~v_439 & ~v_440 & ~v_441 & ~v_442;
assign v_1461 = ~v_443 & ~v_444 & ~v_445 & ~v_446 & ~v_447;
assign v_1462 = ~v_448 & ~v_449;
assign v_1463 = v_1456 & v_1457 & v_1458 & v_1459 & v_1460;
assign v_1464 = v_1461 & v_1462;
assign v_1465 = ~v_450 & ~v_451 & ~v_452 & ~v_453 & ~v_454;
assign v_1466 = ~v_455 & ~v_456 & ~v_457 & ~v_458 & ~v_459;
assign v_1467 = ~v_460 & ~v_461 & ~v_462 & ~v_463 & ~v_464;
assign v_1468 = ~v_465 & ~v_466 & ~v_467 & ~v_468 & ~v_469;
assign v_1469 = ~v_470 & ~v_471 & ~v_472 & ~v_473 & ~v_474;
assign v_1470 = ~v_475 & ~v_476 & ~v_477 & ~v_478 & ~v_479;
assign v_1471 = ~v_480 & ~v_481;
assign v_1472 = v_1465 & v_1466 & v_1467 & v_1468 & v_1469;
assign v_1473 = v_1470 & v_1471;
assign v_1474 = ~v_482 & ~v_483 & ~v_484 & ~v_485 & ~v_486;
assign v_1475 = ~v_487 & ~v_488 & ~v_489 & ~v_490 & ~v_491;
assign v_1476 = ~v_492 & ~v_493 & ~v_494 & ~v_495 & ~v_496;
assign v_1477 = ~v_497 & ~v_498 & ~v_499 & ~v_500 & ~v_501;
assign v_1478 = ~v_502 & ~v_503 & ~v_504 & ~v_505 & ~v_506;
assign v_1479 = ~v_507 & ~v_508 & ~v_509 & ~v_510 & ~v_511;
assign v_1480 = ~v_512 & ~v_513;
assign v_1481 = v_1474 & v_1475 & v_1476 & v_1477 & v_1478;
assign v_1482 = v_1479 & v_1480;
assign v_1483 = ~v_514 & ~v_515 & ~v_516 & ~v_517 & ~v_518;
assign v_1484 = ~v_519 & ~v_520 & ~v_521 & ~v_522 & ~v_523;
assign v_1485 = ~v_524 & ~v_525 & ~v_526 & ~v_527 & ~v_528;
assign v_1486 = ~v_529 & ~v_530 & ~v_531 & ~v_532 & ~v_533;
assign v_1487 = ~v_534 & ~v_535 & ~v_536 & ~v_537 & ~v_538;
assign v_1488 = ~v_539 & ~v_540 & ~v_541 & ~v_542 & ~v_543;
assign v_1489 = ~v_544 & ~v_545;
assign v_1490 = v_1483 & v_1484 & v_1485 & v_1486 & v_1487;
assign v_1491 = v_1488 & v_1489;
assign v_1492 = ~v_546 & ~v_547 & ~v_548 & ~v_549 & ~v_550;
assign v_1493 = ~v_551 & ~v_552 & ~v_553 & ~v_554 & ~v_555;
assign v_1494 = ~v_556 & ~v_557 & ~v_558 & ~v_559 & ~v_560;
assign v_1495 = ~v_561 & ~v_562 & ~v_563 & ~v_564 & ~v_565;
assign v_1496 = ~v_566 & ~v_567 & ~v_568 & ~v_569 & ~v_570;
assign v_1497 = ~v_571 & ~v_572 & ~v_573 & ~v_574 & ~v_575;
assign v_1498 = ~v_576 & ~v_577;
assign v_1499 = v_1492 & v_1493 & v_1494 & v_1495 & v_1496;
assign v_1500 = v_1497 & v_1498;
assign v_1501 = ~v_1199 & ~v_1200 & ~v_1201 & ~v_1202 & ~v_1203;
assign v_1502 = ~v_1204 & ~v_1205 & ~v_1206 & ~v_1207 & ~v_1208;
assign v_1503 = ~v_1209 & ~v_1210 & ~v_1211 & ~v_1212 & ~v_1213;
assign v_1504 = ~v_1214 & ~v_1215 & ~v_1216 & ~v_1217 & ~v_1218;
assign v_1505 = ~v_1219 & ~v_1220 & ~v_1221 & ~v_1222 & ~v_1223;
assign v_1506 = ~v_1224 & ~v_1225 & ~v_1226 & ~v_1227 & ~v_1228;
assign v_1507 = ~v_1229 & ~v_1230;
assign v_1508 = v_1501 & v_1502 & v_1503 & v_1504 & v_1505;
assign v_1509 = v_1506 & v_1507;
assign v_1510 = ~v_1232 & ~v_1233 & ~v_1234 & ~v_1235 & ~v_1236;
assign v_1511 = ~v_1237 & ~v_1238 & ~v_1239 & ~v_1240 & ~v_1241;
assign v_1512 = ~v_1242 & ~v_1243 & ~v_1244 & ~v_1245 & ~v_1246;
assign v_1513 = ~v_1247 & ~v_1248 & ~v_1249 & ~v_1250 & ~v_1251;
assign v_1514 = ~v_1252 & ~v_1253 & ~v_1254 & ~v_1255 & ~v_1256;
assign v_1515 = ~v_1257 & ~v_1258 & ~v_1259 & ~v_1260 & ~v_1261;
assign v_1516 = ~v_1262 & ~v_1263;
assign v_1517 = v_1510 & v_1511 & v_1512 & v_1513 & v_1514;
assign v_1518 = v_1515 & v_1516;
assign v_1519 = ~v_1265 & ~v_1266 & ~v_1267 & ~v_1268 & ~v_1269;
assign v_1520 = ~v_1270 & ~v_1271 & ~v_1272 & ~v_1273 & ~v_1274;
assign v_1521 = ~v_1275 & ~v_1276 & ~v_1277 & ~v_1278 & ~v_1279;
assign v_1522 = ~v_1280 & ~v_1281 & ~v_1282 & ~v_1283 & ~v_1284;
assign v_1523 = ~v_1285 & ~v_1286 & ~v_1287 & ~v_1288 & ~v_1289;
assign v_1524 = ~v_1290 & ~v_1291 & ~v_1292 & ~v_1293 & ~v_1294;
assign v_1525 = ~v_1295 & ~v_1296;
assign v_1526 = v_1519 & v_1520 & v_1521 & v_1522 & v_1523;
assign v_1527 = v_1524 & v_1525;
assign v_1528 = ~v_1298 & ~v_1299 & ~v_1300 & ~v_1301 & ~v_1302;
assign v_1529 = ~v_1303 & ~v_1304 & ~v_1305 & ~v_1306 & ~v_1307;
assign v_1530 = ~v_1308 & ~v_1309 & ~v_1310 & ~v_1311 & ~v_1312;
assign v_1531 = ~v_1313 & ~v_1314 & ~v_1315 & ~v_1316 & ~v_1317;
assign v_1532 = ~v_1318 & ~v_1319 & ~v_1320 & ~v_1321 & ~v_1322;
assign v_1533 = ~v_1323 & ~v_1324 & ~v_1325 & ~v_1326 & ~v_1327;
assign v_1534 = ~v_1328 & ~v_1329;
assign v_1535 = v_1528 & v_1529 & v_1530 & v_1531 & v_1532;
assign v_1536 = v_1533 & v_1534;
assign v_1537 = ~v_1331 & ~v_1332 & ~v_1333 & ~v_1334 & ~v_1335;
assign v_1538 = ~v_1336 & ~v_1337 & ~v_1338 & ~v_1339 & ~v_1340;
assign v_1539 = ~v_1341 & ~v_1342 & ~v_1343 & ~v_1344 & ~v_1345;
assign v_1540 = ~v_1346 & ~v_1347 & ~v_1348 & ~v_1349 & ~v_1350;
assign v_1541 = ~v_1351 & ~v_1352 & ~v_1353 & ~v_1354 & ~v_1355;
assign v_1542 = ~v_1356 & ~v_1357 & ~v_1358 & ~v_1359 & ~v_1360;
assign v_1543 = ~v_1361 & ~v_1362;
assign v_1544 = v_1537 & v_1538 & v_1539 & v_1540 & v_1541;
assign v_1545 = v_1542 & v_1543;
assign v_592 = v_589 | v_590 | v_591;
assign v_598 = v_595 | v_596 | v_597;
assign v_604 = v_601 | v_602 | v_603;
assign v_610 = v_607 | v_608 | v_609;
assign v_616 = v_613 | v_614 | v_615;
assign v_622 = v_619 | v_620 | v_621;
assign v_628 = v_625 | v_626 | v_627;
assign v_634 = v_631 | v_632 | v_633;
assign v_640 = v_637 | v_638 | v_639;
assign v_646 = v_643 | v_644 | v_645;
assign v_652 = v_649 | v_650 | v_651;
assign v_658 = v_655 | v_656 | v_657;
assign v_664 = v_661 | v_662 | v_663;
assign v_670 = v_667 | v_668 | v_669;
assign v_676 = v_673 | v_674 | v_675;
assign v_682 = v_679 | v_680 | v_681;
assign v_688 = v_685 | v_686 | v_687;
assign v_694 = v_691 | v_692 | v_693;
assign v_700 = v_697 | v_698 | v_699;
assign v_706 = v_703 | v_704 | v_705;
assign v_712 = v_709 | v_710 | v_711;
assign v_718 = v_715 | v_716 | v_717;
assign v_724 = v_721 | v_722 | v_723;
assign v_730 = v_727 | v_728 | v_729;
assign v_736 = v_733 | v_734 | v_735;
assign v_742 = v_739 | v_740 | v_741;
assign v_748 = v_745 | v_746 | v_747;
assign v_754 = v_751 | v_752 | v_753;
assign v_760 = v_757 | v_758 | v_759;
assign v_766 = v_763 | v_764 | v_765;
assign v_772 = v_769 | v_770 | v_771;
assign v_846 = v_843 | v_844 | v_845;
assign v_852 = v_849 | v_850 | v_851;
assign v_858 = v_855 | v_856 | v_857;
assign v_864 = v_861 | v_862 | v_863;
assign v_870 = v_867 | v_868 | v_869;
assign v_876 = v_873 | v_874 | v_875;
assign v_882 = v_879 | v_880 | v_881;
assign v_888 = v_885 | v_886 | v_887;
assign v_894 = v_891 | v_892 | v_893;
assign v_900 = v_897 | v_898 | v_899;
assign v_906 = v_903 | v_904 | v_905;
assign v_912 = v_909 | v_910 | v_911;
assign v_918 = v_915 | v_916 | v_917;
assign v_924 = v_921 | v_922 | v_923;
assign v_930 = v_927 | v_928 | v_929;
assign v_936 = v_933 | v_934 | v_935;
assign v_942 = v_939 | v_940 | v_941;
assign v_948 = v_945 | v_946 | v_947;
assign v_954 = v_951 | v_952 | v_953;
assign v_960 = v_957 | v_958 | v_959;
assign v_966 = v_963 | v_964 | v_965;
assign v_972 = v_969 | v_970 | v_971;
assign v_978 = v_975 | v_976 | v_977;
assign v_984 = v_981 | v_982 | v_983;
assign v_990 = v_987 | v_988 | v_989;
assign v_996 = v_993 | v_994 | v_995;
assign v_1002 = v_999 | v_1000 | v_1001;
assign v_1008 = v_1005 | v_1006 | v_1007;
assign v_1014 = v_1011 | v_1012 | v_1013;
assign v_1020 = v_1017 | v_1018 | v_1019;
assign v_1026 = v_1023 | v_1024 | v_1025;
assign v_584 = v_33 ^ v_65;
assign v_587 = v_34 ^ v_66;
assign v_588 = v_586 ^ v_587;
assign v_593 = v_35 ^ v_67;
assign v_594 = v_592 ^ v_593;
assign v_599 = v_36 ^ v_68;
assign v_600 = v_598 ^ v_599;
assign v_605 = v_37 ^ v_69;
assign v_606 = v_604 ^ v_605;
assign v_611 = v_38 ^ v_70;
assign v_612 = v_610 ^ v_611;
assign v_617 = v_39 ^ v_71;
assign v_618 = v_616 ^ v_617;
assign v_623 = v_40 ^ v_72;
assign v_624 = v_622 ^ v_623;
assign v_629 = v_41 ^ v_73;
assign v_630 = v_628 ^ v_629;
assign v_635 = v_42 ^ v_74;
assign v_636 = v_634 ^ v_635;
assign v_641 = v_43 ^ v_75;
assign v_642 = v_640 ^ v_641;
assign v_647 = v_44 ^ v_76;
assign v_648 = v_646 ^ v_647;
assign v_653 = v_45 ^ v_77;
assign v_654 = v_652 ^ v_653;
assign v_659 = v_46 ^ v_78;
assign v_660 = v_658 ^ v_659;
assign v_665 = v_47 ^ v_79;
assign v_666 = v_664 ^ v_665;
assign v_671 = v_48 ^ v_80;
assign v_672 = v_670 ^ v_671;
assign v_677 = v_49 ^ v_81;
assign v_678 = v_676 ^ v_677;
assign v_683 = v_50 ^ v_82;
assign v_684 = v_682 ^ v_683;
assign v_689 = v_51 ^ v_83;
assign v_690 = v_688 ^ v_689;
assign v_695 = v_52 ^ v_84;
assign v_696 = v_694 ^ v_695;
assign v_701 = v_53 ^ v_85;
assign v_702 = v_700 ^ v_701;
assign v_707 = v_54 ^ v_86;
assign v_708 = v_706 ^ v_707;
assign v_713 = v_55 ^ v_87;
assign v_714 = v_712 ^ v_713;
assign v_719 = v_56 ^ v_88;
assign v_720 = v_718 ^ v_719;
assign v_725 = v_57 ^ v_89;
assign v_726 = v_724 ^ v_725;
assign v_731 = v_58 ^ v_90;
assign v_732 = v_730 ^ v_731;
assign v_737 = v_59 ^ v_91;
assign v_738 = v_736 ^ v_737;
assign v_743 = v_60 ^ v_92;
assign v_744 = v_742 ^ v_743;
assign v_749 = v_61 ^ v_93;
assign v_750 = v_748 ^ v_749;
assign v_755 = v_62 ^ v_94;
assign v_756 = v_754 ^ v_755;
assign v_761 = v_63 ^ v_95;
assign v_762 = v_760 ^ v_761;
assign v_767 = v_64 ^ v_96;
assign v_768 = v_766 ^ v_767;
assign v_805 = v_773 ^ v_161;
assign v_806 = v_774 ^ v_162;
assign v_807 = v_775 ^ v_163;
assign v_808 = v_776 ^ v_164;
assign v_809 = v_777 ^ v_165;
assign v_810 = v_778 ^ v_166;
assign v_811 = v_779 ^ v_167;
assign v_812 = v_780 ^ v_168;
assign v_813 = v_781 ^ v_169;
assign v_814 = v_782 ^ v_170;
assign v_815 = v_783 ^ v_171;
assign v_816 = v_784 ^ v_172;
assign v_817 = v_785 ^ v_173;
assign v_818 = v_786 ^ v_174;
assign v_819 = v_787 ^ v_175;
assign v_820 = v_788 ^ v_176;
assign v_821 = v_789 ^ v_177;
assign v_822 = v_790 ^ v_178;
assign v_823 = v_791 ^ v_179;
assign v_824 = v_792 ^ v_180;
assign v_825 = v_793 ^ v_181;
assign v_826 = v_794 ^ v_182;
assign v_827 = v_795 ^ v_183;
assign v_828 = v_796 ^ v_184;
assign v_829 = v_797 ^ v_185;
assign v_830 = v_798 ^ v_186;
assign v_831 = v_799 ^ v_187;
assign v_832 = v_800 ^ v_188;
assign v_833 = v_801 ^ v_189;
assign v_834 = v_802 ^ v_190;
assign v_835 = v_803 ^ v_191;
assign v_836 = v_804 ^ v_192;
assign v_838 = v_258 ^ v_226;
assign v_841 = v_259 ^ v_227;
assign v_842 = v_840 ^ v_841;
assign v_847 = v_260 ^ v_228;
assign v_848 = v_846 ^ v_847;
assign v_853 = v_261 ^ v_229;
assign v_854 = v_852 ^ v_853;
assign v_859 = v_262 ^ v_230;
assign v_860 = v_858 ^ v_859;
assign v_865 = v_263 ^ v_231;
assign v_866 = v_864 ^ v_865;
assign v_871 = v_264 ^ v_232;
assign v_872 = v_870 ^ v_871;
assign v_877 = v_265 ^ v_233;
assign v_878 = v_876 ^ v_877;
assign v_883 = v_266 ^ v_234;
assign v_884 = v_882 ^ v_883;
assign v_889 = v_267 ^ v_235;
assign v_890 = v_888 ^ v_889;
assign v_895 = v_268 ^ v_236;
assign v_896 = v_894 ^ v_895;
assign v_901 = v_269 ^ v_237;
assign v_902 = v_900 ^ v_901;
assign v_907 = v_270 ^ v_238;
assign v_908 = v_906 ^ v_907;
assign v_913 = v_271 ^ v_239;
assign v_914 = v_912 ^ v_913;
assign v_919 = v_272 ^ v_240;
assign v_920 = v_918 ^ v_919;
assign v_925 = v_273 ^ v_241;
assign v_926 = v_924 ^ v_925;
assign v_931 = v_274 ^ v_242;
assign v_932 = v_930 ^ v_931;
assign v_937 = v_275 ^ v_243;
assign v_938 = v_936 ^ v_937;
assign v_943 = v_276 ^ v_244;
assign v_944 = v_942 ^ v_943;
assign v_949 = v_277 ^ v_245;
assign v_950 = v_948 ^ v_949;
assign v_955 = v_278 ^ v_246;
assign v_956 = v_954 ^ v_955;
assign v_961 = v_279 ^ v_247;
assign v_962 = v_960 ^ v_961;
assign v_967 = v_280 ^ v_248;
assign v_968 = v_966 ^ v_967;
assign v_973 = v_281 ^ v_249;
assign v_974 = v_972 ^ v_973;
assign v_979 = v_282 ^ v_250;
assign v_980 = v_978 ^ v_979;
assign v_985 = v_283 ^ v_251;
assign v_986 = v_984 ^ v_985;
assign v_991 = v_284 ^ v_252;
assign v_992 = v_990 ^ v_991;
assign v_997 = v_285 ^ v_253;
assign v_998 = v_996 ^ v_997;
assign v_1003 = v_286 ^ v_254;
assign v_1004 = v_1002 ^ v_1003;
assign v_1009 = v_287 ^ v_255;
assign v_1010 = v_1008 ^ v_1009;
assign v_1015 = v_288 ^ v_256;
assign v_1016 = v_1014 ^ v_1015;
assign v_1021 = v_289 ^ v_257;
assign v_1022 = v_1020 ^ v_1021;
assign v_1027 = v_838 ^ v_194;
assign v_1028 = v_842 ^ v_195;
assign v_1029 = v_848 ^ v_196;
assign v_1030 = v_854 ^ v_197;
assign v_1031 = v_860 ^ v_198;
assign v_1032 = v_866 ^ v_199;
assign v_1033 = v_872 ^ v_200;
assign v_1034 = v_878 ^ v_201;
assign v_1035 = v_884 ^ v_202;
assign v_1036 = v_890 ^ v_203;
assign v_1037 = v_896 ^ v_204;
assign v_1038 = v_902 ^ v_205;
assign v_1039 = v_908 ^ v_206;
assign v_1040 = v_914 ^ v_207;
assign v_1041 = v_920 ^ v_208;
assign v_1042 = v_926 ^ v_209;
assign v_1043 = v_932 ^ v_210;
assign v_1044 = v_938 ^ v_211;
assign v_1045 = v_944 ^ v_212;
assign v_1046 = v_950 ^ v_213;
assign v_1047 = v_956 ^ v_214;
assign v_1048 = v_962 ^ v_215;
assign v_1049 = v_968 ^ v_216;
assign v_1050 = v_974 ^ v_217;
assign v_1051 = v_980 ^ v_218;
assign v_1052 = v_986 ^ v_219;
assign v_1053 = v_992 ^ v_220;
assign v_1054 = v_998 ^ v_221;
assign v_1055 = v_1004 ^ v_222;
assign v_1056 = v_1010 ^ v_223;
assign v_1057 = v_1016 ^ v_224;
assign v_1058 = v_1022 ^ v_225;
assign v_1092 = v_1060 ^ v_290;
assign v_1093 = v_1061 ^ v_291;
assign v_1094 = v_1062 ^ v_292;
assign v_1095 = v_1063 ^ v_293;
assign v_1096 = v_1064 ^ v_294;
assign v_1097 = v_1065 ^ v_295;
assign v_1098 = v_1066 ^ v_296;
assign v_1099 = v_1067 ^ v_297;
assign v_1100 = v_1068 ^ v_298;
assign v_1101 = v_1069 ^ v_299;
assign v_1102 = v_1070 ^ v_300;
assign v_1103 = v_1071 ^ v_301;
assign v_1104 = v_1072 ^ v_302;
assign v_1105 = v_1073 ^ v_303;
assign v_1106 = v_1074 ^ v_304;
assign v_1107 = v_1075 ^ v_305;
assign v_1108 = v_1076 ^ v_306;
assign v_1109 = v_1077 ^ v_307;
assign v_1110 = v_1078 ^ v_308;
assign v_1111 = v_1079 ^ v_309;
assign v_1112 = v_1080 ^ v_310;
assign v_1113 = v_1081 ^ v_311;
assign v_1114 = v_1082 ^ v_312;
assign v_1115 = v_1083 ^ v_313;
assign v_1116 = v_1084 ^ v_314;
assign v_1117 = v_1085 ^ v_315;
assign v_1118 = v_1086 ^ v_316;
assign v_1119 = v_1087 ^ v_317;
assign v_1120 = v_1088 ^ v_318;
assign v_1121 = v_1089 ^ v_319;
assign v_1122 = v_1090 ^ v_320;
assign v_1123 = v_1091 ^ v_321;
assign v_1125 = v_33 ^ v_354;
assign v_1126 = v_34 ^ v_355;
assign v_1127 = v_35 ^ v_356;
assign v_1128 = v_36 ^ v_357;
assign v_1129 = v_37 ^ v_358;
assign v_1130 = v_38 ^ v_359;
assign v_1131 = v_39 ^ v_360;
assign v_1132 = v_40 ^ v_361;
assign v_1133 = v_41 ^ v_362;
assign v_1134 = v_42 ^ v_363;
assign v_1135 = v_43 ^ v_364;
assign v_1136 = v_44 ^ v_365;
assign v_1137 = v_45 ^ v_366;
assign v_1138 = v_46 ^ v_367;
assign v_1139 = v_47 ^ v_368;
assign v_1140 = v_48 ^ v_369;
assign v_1141 = v_49 ^ v_370;
assign v_1142 = v_50 ^ v_371;
assign v_1143 = v_51 ^ v_372;
assign v_1144 = v_52 ^ v_373;
assign v_1145 = v_53 ^ v_374;
assign v_1146 = v_54 ^ v_375;
assign v_1147 = v_55 ^ v_376;
assign v_1148 = v_56 ^ v_377;
assign v_1149 = v_57 ^ v_378;
assign v_1150 = v_58 ^ v_379;
assign v_1151 = v_59 ^ v_380;
assign v_1152 = v_60 ^ v_381;
assign v_1153 = v_61 ^ v_382;
assign v_1154 = v_62 ^ v_383;
assign v_1155 = v_63 ^ v_384;
assign v_1156 = v_64 ^ v_385;
assign v_1158 = v_65 ^ v_386;
assign v_1159 = v_66 ^ v_387;
assign v_1160 = v_67 ^ v_388;
assign v_1161 = v_68 ^ v_389;
assign v_1162 = v_69 ^ v_390;
assign v_1163 = v_70 ^ v_391;
assign v_1164 = v_71 ^ v_392;
assign v_1165 = v_72 ^ v_393;
assign v_1166 = v_73 ^ v_394;
assign v_1167 = v_74 ^ v_395;
assign v_1168 = v_75 ^ v_396;
assign v_1169 = v_76 ^ v_397;
assign v_1170 = v_77 ^ v_398;
assign v_1171 = v_78 ^ v_399;
assign v_1172 = v_79 ^ v_400;
assign v_1173 = v_80 ^ v_401;
assign v_1174 = v_81 ^ v_402;
assign v_1175 = v_82 ^ v_403;
assign v_1176 = v_83 ^ v_404;
assign v_1177 = v_84 ^ v_405;
assign v_1178 = v_85 ^ v_406;
assign v_1179 = v_86 ^ v_407;
assign v_1180 = v_87 ^ v_408;
assign v_1181 = v_88 ^ v_409;
assign v_1182 = v_89 ^ v_410;
assign v_1183 = v_90 ^ v_411;
assign v_1184 = v_91 ^ v_412;
assign v_1185 = v_92 ^ v_413;
assign v_1186 = v_93 ^ v_414;
assign v_1187 = v_94 ^ v_415;
assign v_1188 = v_95 ^ v_416;
assign v_1189 = v_96 ^ v_417;
assign v_1199 = v_418 ^ v_161;
assign v_1200 = v_419 ^ v_162;
assign v_1201 = v_420 ^ v_163;
assign v_1202 = v_421 ^ v_164;
assign v_1203 = v_422 ^ v_165;
assign v_1204 = v_423 ^ v_166;
assign v_1205 = v_424 ^ v_167;
assign v_1206 = v_425 ^ v_168;
assign v_1207 = v_426 ^ v_169;
assign v_1208 = v_427 ^ v_170;
assign v_1209 = v_428 ^ v_171;
assign v_1210 = v_429 ^ v_172;
assign v_1211 = v_430 ^ v_173;
assign v_1212 = v_431 ^ v_174;
assign v_1213 = v_432 ^ v_175;
assign v_1214 = v_433 ^ v_176;
assign v_1215 = v_434 ^ v_177;
assign v_1216 = v_435 ^ v_178;
assign v_1217 = v_436 ^ v_179;
assign v_1218 = v_437 ^ v_180;
assign v_1219 = v_438 ^ v_181;
assign v_1220 = v_439 ^ v_182;
assign v_1221 = v_440 ^ v_183;
assign v_1222 = v_441 ^ v_184;
assign v_1223 = v_442 ^ v_185;
assign v_1224 = v_443 ^ v_186;
assign v_1225 = v_444 ^ v_187;
assign v_1226 = v_445 ^ v_188;
assign v_1227 = v_446 ^ v_189;
assign v_1228 = v_447 ^ v_190;
assign v_1229 = v_448 ^ v_191;
assign v_1230 = v_449 ^ v_192;
assign v_1232 = v_450 ^ v_194;
assign v_1233 = v_451 ^ v_195;
assign v_1234 = v_452 ^ v_196;
assign v_1235 = v_453 ^ v_197;
assign v_1236 = v_454 ^ v_198;
assign v_1237 = v_455 ^ v_199;
assign v_1238 = v_456 ^ v_200;
assign v_1239 = v_457 ^ v_201;
assign v_1240 = v_458 ^ v_202;
assign v_1241 = v_459 ^ v_203;
assign v_1242 = v_460 ^ v_204;
assign v_1243 = v_461 ^ v_205;
assign v_1244 = v_462 ^ v_206;
assign v_1245 = v_463 ^ v_207;
assign v_1246 = v_464 ^ v_208;
assign v_1247 = v_465 ^ v_209;
assign v_1248 = v_466 ^ v_210;
assign v_1249 = v_467 ^ v_211;
assign v_1250 = v_468 ^ v_212;
assign v_1251 = v_469 ^ v_213;
assign v_1252 = v_470 ^ v_214;
assign v_1253 = v_471 ^ v_215;
assign v_1254 = v_472 ^ v_216;
assign v_1255 = v_473 ^ v_217;
assign v_1256 = v_474 ^ v_218;
assign v_1257 = v_475 ^ v_219;
assign v_1258 = v_476 ^ v_220;
assign v_1259 = v_477 ^ v_221;
assign v_1260 = v_478 ^ v_222;
assign v_1261 = v_479 ^ v_223;
assign v_1262 = v_480 ^ v_224;
assign v_1263 = v_481 ^ v_225;
assign v_1265 = v_482 ^ v_290;
assign v_1266 = v_483 ^ v_291;
assign v_1267 = v_484 ^ v_292;
assign v_1268 = v_485 ^ v_293;
assign v_1269 = v_486 ^ v_294;
assign v_1270 = v_487 ^ v_295;
assign v_1271 = v_488 ^ v_296;
assign v_1272 = v_489 ^ v_297;
assign v_1273 = v_490 ^ v_298;
assign v_1274 = v_491 ^ v_299;
assign v_1275 = v_492 ^ v_300;
assign v_1276 = v_493 ^ v_301;
assign v_1277 = v_494 ^ v_302;
assign v_1278 = v_495 ^ v_303;
assign v_1279 = v_496 ^ v_304;
assign v_1280 = v_497 ^ v_305;
assign v_1281 = v_498 ^ v_306;
assign v_1282 = v_499 ^ v_307;
assign v_1283 = v_500 ^ v_308;
assign v_1284 = v_501 ^ v_309;
assign v_1285 = v_502 ^ v_310;
assign v_1286 = v_503 ^ v_311;
assign v_1287 = v_504 ^ v_312;
assign v_1288 = v_505 ^ v_313;
assign v_1289 = v_506 ^ v_314;
assign v_1290 = v_507 ^ v_315;
assign v_1291 = v_508 ^ v_316;
assign v_1292 = v_509 ^ v_317;
assign v_1293 = v_510 ^ v_318;
assign v_1294 = v_511 ^ v_319;
assign v_1295 = v_512 ^ v_320;
assign v_1296 = v_513 ^ v_321;
assign v_1298 = v_514 ^ v_354;
assign v_1299 = v_515 ^ v_355;
assign v_1300 = v_516 ^ v_356;
assign v_1301 = v_517 ^ v_357;
assign v_1302 = v_518 ^ v_358;
assign v_1303 = v_519 ^ v_359;
assign v_1304 = v_520 ^ v_360;
assign v_1305 = v_521 ^ v_361;
assign v_1306 = v_522 ^ v_362;
assign v_1307 = v_523 ^ v_363;
assign v_1308 = v_524 ^ v_364;
assign v_1309 = v_525 ^ v_365;
assign v_1310 = v_526 ^ v_366;
assign v_1311 = v_527 ^ v_367;
assign v_1312 = v_528 ^ v_368;
assign v_1313 = v_529 ^ v_369;
assign v_1314 = v_530 ^ v_370;
assign v_1315 = v_531 ^ v_371;
assign v_1316 = v_532 ^ v_372;
assign v_1317 = v_533 ^ v_373;
assign v_1318 = v_534 ^ v_374;
assign v_1319 = v_535 ^ v_375;
assign v_1320 = v_536 ^ v_376;
assign v_1321 = v_537 ^ v_377;
assign v_1322 = v_538 ^ v_378;
assign v_1323 = v_539 ^ v_379;
assign v_1324 = v_540 ^ v_380;
assign v_1325 = v_541 ^ v_381;
assign v_1326 = v_542 ^ v_382;
assign v_1327 = v_543 ^ v_383;
assign v_1328 = v_544 ^ v_384;
assign v_1329 = v_545 ^ v_385;
assign v_1331 = v_546 ^ v_386;
assign v_1332 = v_547 ^ v_387;
assign v_1333 = v_548 ^ v_388;
assign v_1334 = v_549 ^ v_389;
assign v_1335 = v_550 ^ v_390;
assign v_1336 = v_551 ^ v_391;
assign v_1337 = v_552 ^ v_392;
assign v_1338 = v_553 ^ v_393;
assign v_1339 = v_554 ^ v_394;
assign v_1340 = v_555 ^ v_395;
assign v_1341 = v_556 ^ v_396;
assign v_1342 = v_557 ^ v_397;
assign v_1343 = v_558 ^ v_398;
assign v_1344 = v_559 ^ v_399;
assign v_1345 = v_560 ^ v_400;
assign v_1346 = v_561 ^ v_401;
assign v_1347 = v_562 ^ v_402;
assign v_1348 = v_563 ^ v_403;
assign v_1349 = v_564 ^ v_404;
assign v_1350 = v_565 ^ v_405;
assign v_1351 = v_566 ^ v_406;
assign v_1352 = v_567 ^ v_407;
assign v_1353 = v_568 ^ v_408;
assign v_1354 = v_569 ^ v_409;
assign v_1355 = v_570 ^ v_410;
assign v_1356 = v_571 ^ v_411;
assign v_1357 = v_572 ^ v_412;
assign v_1358 = v_573 ^ v_413;
assign v_1359 = v_574 ^ v_414;
assign v_1360 = v_575 ^ v_415;
assign v_1361 = v_576 ^ v_416;
assign v_1362 = v_577 ^ v_417;
assign x_1 = v_1365 | ~v_1192;
assign o_1 = x_1;
endmodule
