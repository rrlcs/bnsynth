// skolem function for order file variables
// Generated using findDep.cpp 
module small-dyn-partition-fixpoint-4 (v_1, v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_12, v_13, v_14, v_15, v_16, v_17, v_18, v_19, v_20, v_21, v_22, v_23, v_24, v_25, v_26, v_27, v_28, v_29, v_30, v_31, v_32, v_33, v_34, v_35, v_36, v_37, v_38, v_39, v_40, v_41, v_42, v_43, v_44, v_45, v_46, v_47, v_48, v_49, v_50, v_51, v_52, v_53, v_54, v_55, v_56, v_57, v_58, v_59, v_60, v_61, v_62, v_63, v_64, v_65, v_66, v_67, v_68, v_69, v_70, v_71, v_72, o_1);
input v_1;
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_13;
input v_14;
input v_15;
input v_16;
input v_17;
input v_18;
input v_19;
input v_20;
input v_21;
input v_22;
input v_23;
input v_24;
input v_25;
input v_26;
input v_27;
input v_28;
input v_29;
input v_30;
input v_31;
input v_32;
input v_33;
input v_34;
input v_35;
input v_36;
input v_37;
input v_38;
input v_39;
input v_40;
input v_41;
input v_42;
input v_43;
input v_44;
input v_45;
input v_46;
input v_47;
input v_48;
input v_49;
input v_50;
input v_51;
input v_52;
input v_53;
input v_54;
input v_55;
input v_56;
input v_57;
input v_58;
input v_59;
input v_60;
input v_61;
input v_62;
input v_63;
input v_64;
input v_65;
input v_66;
input v_67;
input v_68;
input v_69;
input v_70;
input v_71;
input v_72;
output o_1;
wire v_73;
wire v_74;
wire v_75;
wire v_76;
wire v_77;
wire v_78;
wire v_79;
wire v_80;
wire v_81;
wire v_82;
wire v_83;
wire v_84;
wire v_85;
wire v_86;
wire v_87;
wire v_88;
wire v_89;
wire v_90;
wire v_91;
wire v_92;
wire v_93;
wire v_94;
wire v_95;
wire v_96;
wire v_97;
wire v_98;
wire v_99;
wire v_100;
wire v_101;
wire v_102;
wire v_103;
wire v_104;
wire v_105;
wire v_106;
wire v_107;
wire v_108;
wire v_109;
wire v_110;
wire v_111;
wire v_112;
wire v_113;
wire v_114;
wire v_115;
wire v_116;
wire v_117;
wire v_118;
wire v_119;
wire v_120;
wire v_121;
wire v_122;
wire v_123;
wire v_124;
wire v_125;
wire v_126;
wire v_127;
wire v_128;
wire v_129;
wire v_130;
wire v_131;
wire v_132;
wire v_133;
wire v_134;
wire v_135;
wire v_136;
wire v_137;
wire v_138;
wire v_139;
wire v_140;
wire v_141;
wire v_142;
wire v_143;
wire v_144;
wire v_145;
wire v_146;
wire v_147;
wire v_148;
wire v_149;
wire v_150;
wire v_151;
wire v_152;
wire v_153;
wire v_154;
wire v_155;
wire v_156;
wire v_157;
wire v_158;
wire v_159;
wire v_160;
wire v_161;
wire v_162;
wire v_163;
wire v_164;
wire v_165;
wire v_166;
wire v_167;
wire v_168;
wire v_169;
wire v_170;
wire v_171;
wire v_172;
wire v_173;
wire v_174;
wire v_175;
wire v_176;
wire v_177;
wire v_178;
wire v_179;
wire v_180;
wire v_181;
wire v_182;
wire v_183;
wire v_184;
wire v_185;
wire v_186;
wire v_187;
wire v_188;
wire v_189;
wire v_190;
wire v_191;
wire v_192;
wire v_193;
wire v_194;
wire v_195;
wire v_196;
wire v_197;
wire v_198;
wire v_199;
wire v_200;
wire v_201;
wire v_202;
wire v_203;
wire v_204;
wire v_205;
wire v_206;
wire v_207;
wire v_208;
wire v_209;
wire v_210;
wire v_211;
wire v_212;
wire v_213;
wire v_214;
wire v_215;
wire v_216;
wire v_217;
wire v_218;
wire v_219;
wire v_220;
wire v_221;
wire v_222;
wire v_223;
wire v_224;
wire v_225;
wire v_226;
wire v_227;
wire v_228;
wire v_229;
wire v_230;
wire v_231;
wire v_232;
wire v_233;
wire v_234;
wire v_235;
wire v_236;
wire v_237;
wire v_238;
wire v_239;
wire v_240;
wire v_241;
wire v_242;
wire v_243;
wire v_244;
wire v_245;
wire v_246;
wire v_247;
wire v_248;
wire v_249;
wire v_250;
wire v_251;
wire v_252;
wire v_253;
wire v_254;
wire v_255;
wire v_256;
wire v_257;
wire v_258;
wire v_259;
wire v_260;
wire v_261;
wire v_262;
wire v_263;
wire v_264;
wire v_265;
wire v_266;
wire v_267;
wire v_268;
wire v_269;
wire v_270;
wire v_271;
wire v_272;
wire v_273;
wire v_274;
wire v_275;
wire v_276;
wire v_277;
wire v_278;
wire v_279;
wire v_280;
wire v_281;
wire v_282;
wire v_283;
wire v_284;
wire v_285;
wire v_286;
wire v_287;
wire v_288;
wire v_289;
wire v_290;
wire v_291;
wire v_292;
wire v_293;
wire v_294;
wire v_295;
wire v_296;
wire v_297;
wire v_298;
wire v_299;
wire v_300;
wire v_301;
wire v_302;
wire v_303;
wire v_304;
wire v_305;
wire v_306;
wire v_307;
wire v_308;
wire v_309;
wire v_310;
wire v_311;
wire v_312;
wire v_313;
wire v_314;
wire v_315;
wire v_316;
wire v_317;
wire v_318;
wire v_319;
wire v_320;
wire v_321;
wire v_322;
wire v_323;
wire v_324;
wire v_325;
wire v_326;
wire v_327;
wire v_328;
wire v_329;
wire v_330;
wire v_331;
wire v_332;
wire v_333;
wire v_334;
wire v_335;
wire v_336;
wire v_337;
wire v_338;
wire v_339;
wire v_340;
wire v_341;
wire v_342;
wire v_343;
wire v_344;
wire v_345;
wire v_346;
wire v_347;
wire v_348;
wire v_349;
wire v_350;
wire v_351;
wire v_352;
wire v_353;
wire v_354;
wire v_355;
wire v_356;
wire v_357;
wire v_358;
wire v_359;
wire v_360;
wire v_361;
wire v_362;
wire v_363;
wire v_364;
wire v_365;
wire v_366;
wire v_367;
wire v_368;
wire v_369;
wire v_370;
wire v_371;
wire v_372;
wire v_373;
wire v_374;
wire v_375;
wire v_376;
wire v_377;
wire v_378;
wire v_379;
wire v_380;
wire v_381;
wire v_382;
wire v_383;
wire v_384;
wire v_385;
wire v_386;
wire v_387;
wire v_388;
wire v_389;
wire v_390;
wire v_391;
wire v_392;
wire v_393;
wire v_394;
wire v_395;
wire v_396;
wire v_397;
wire v_398;
wire v_399;
wire v_400;
wire v_401;
wire v_402;
wire v_403;
wire v_404;
wire v_405;
wire v_406;
wire v_407;
wire v_408;
wire v_409;
wire v_410;
wire v_411;
wire v_412;
wire v_413;
wire v_414;
wire v_415;
wire v_416;
wire v_417;
wire v_418;
wire v_419;
wire v_420;
wire v_421;
wire v_422;
wire v_423;
wire v_424;
wire v_425;
wire v_426;
wire v_427;
wire v_428;
wire v_429;
wire v_430;
wire v_431;
wire v_432;
wire v_433;
wire v_434;
wire x_1;
assign v_73 = ~v_1 & ~v_2 & ~v_3;
assign v_74 = ~v_4 & ~v_5 & ~v_6;
assign v_75 = ~v_7 & ~v_8 & v_73 & v_74;
assign v_77 = v_1;
assign v_79 = v_2 & v_77;
assign v_80 = v_79;
assign v_82 = v_3 & v_80;
assign v_83 = v_82;
assign v_84 = ~v_76 & ~v_1;
assign v_85 = v_76 & v_1;
assign v_87 = ~v_76 & v_78;
assign v_88 = v_76 & v_2;
assign v_90 = ~v_76 & v_81;
assign v_91 = v_76 & v_3;
assign v_96 = ~v_93 & ~v_94 & ~v_95;
assign v_97 = v_4;
assign v_99 = v_5 & v_97;
assign v_100 = v_99;
assign v_102 = v_6 & v_100;
assign v_103 = v_102;
assign v_104 = ~v_76 & v_4;
assign v_105 = ~v_4 & v_76;
assign v_107 = ~v_76 & v_5;
assign v_108 = v_76 & v_98;
assign v_110 = ~v_76 & v_6;
assign v_111 = v_76 & v_101;
assign v_116 = ~v_113 & ~v_114 & ~v_115;
assign v_119 = ~v_117 & ~v_118 & v_96 & v_116;
assign v_121 = v_9;
assign v_123 = v_10 & v_121;
assign v_124 = v_123;
assign v_126 = v_11 & v_124;
assign v_127 = v_126;
assign v_128 = ~v_120 & ~v_9;
assign v_129 = v_120 & v_9;
assign v_131 = ~v_120 & v_122;
assign v_132 = v_120 & v_10;
assign v_134 = ~v_120 & v_125;
assign v_135 = v_120 & v_11;
assign v_140 = ~v_137 & ~v_138 & ~v_139;
assign v_141 = v_12;
assign v_143 = v_13 & v_141;
assign v_144 = v_143;
assign v_146 = v_14 & v_144;
assign v_147 = v_146;
assign v_148 = ~v_120 & v_12;
assign v_149 = ~v_12 & v_120;
assign v_151 = ~v_120 & v_13;
assign v_152 = v_120 & v_142;
assign v_154 = ~v_120 & v_14;
assign v_155 = v_120 & v_145;
assign v_160 = ~v_157 & ~v_158 & ~v_159;
assign v_163 = ~v_161 & ~v_162 & v_140 & v_160;
assign v_165 = v_17;
assign v_167 = v_18 & v_165;
assign v_168 = v_167;
assign v_170 = v_19 & v_168;
assign v_171 = v_170;
assign v_172 = ~v_164 & ~v_17;
assign v_173 = v_164 & v_17;
assign v_175 = ~v_164 & v_166;
assign v_176 = v_164 & v_18;
assign v_178 = ~v_164 & v_169;
assign v_179 = v_164 & v_19;
assign v_184 = ~v_181 & ~v_182 & ~v_183;
assign v_185 = v_20;
assign v_187 = v_21 & v_185;
assign v_188 = v_187;
assign v_190 = v_22 & v_188;
assign v_191 = v_190;
assign v_192 = ~v_164 & v_20;
assign v_193 = ~v_20 & v_164;
assign v_195 = ~v_164 & v_21;
assign v_196 = v_164 & v_186;
assign v_198 = ~v_164 & v_22;
assign v_199 = v_164 & v_189;
assign v_204 = ~v_201 & ~v_202 & ~v_203;
assign v_207 = ~v_205 & ~v_206 & v_184 & v_204;
assign v_209 = v_25;
assign v_211 = v_26 & v_209;
assign v_212 = v_211;
assign v_214 = v_27 & v_212;
assign v_215 = v_214;
assign v_216 = ~v_208 & ~v_25;
assign v_217 = v_208 & v_25;
assign v_219 = ~v_208 & v_210;
assign v_220 = v_208 & v_26;
assign v_222 = ~v_208 & v_213;
assign v_223 = v_208 & v_27;
assign v_228 = ~v_225 & ~v_226 & ~v_227;
assign v_229 = v_28;
assign v_231 = v_29 & v_229;
assign v_232 = v_231;
assign v_234 = v_30 & v_232;
assign v_235 = v_234;
assign v_236 = ~v_208 & v_28;
assign v_237 = ~v_28 & v_208;
assign v_239 = ~v_208 & v_29;
assign v_240 = v_208 & v_230;
assign v_242 = ~v_208 & v_30;
assign v_243 = v_208 & v_233;
assign v_248 = ~v_245 & ~v_246 & ~v_247;
assign v_251 = ~v_249 & ~v_250 & v_228 & v_248;
assign v_252 = v_75 & v_119 & v_163 & v_207 & v_251;
assign v_253 = ~v_41 & ~v_42 & ~v_43;
assign v_254 = ~v_44 & ~v_45 & ~v_46;
assign v_255 = ~v_47 & ~v_48 & v_253 & v_254;
assign v_257 = v_41;
assign v_259 = v_42 & v_257;
assign v_260 = v_259;
assign v_262 = v_43 & v_260;
assign v_263 = v_262;
assign v_264 = ~v_256 & ~v_41;
assign v_265 = v_256 & v_41;
assign v_267 = ~v_256 & v_258;
assign v_268 = v_256 & v_42;
assign v_270 = ~v_256 & v_261;
assign v_271 = v_256 & v_43;
assign v_276 = ~v_273 & ~v_274 & ~v_275;
assign v_277 = v_44;
assign v_279 = v_45 & v_277;
assign v_280 = v_279;
assign v_282 = v_46 & v_280;
assign v_283 = v_282;
assign v_284 = ~v_256 & v_44;
assign v_285 = ~v_44 & v_256;
assign v_287 = ~v_256 & v_45;
assign v_288 = v_256 & v_278;
assign v_290 = ~v_256 & v_46;
assign v_291 = v_256 & v_281;
assign v_296 = ~v_293 & ~v_294 & ~v_295;
assign v_299 = ~v_297 & ~v_298 & v_276 & v_296;
assign v_301 = v_49;
assign v_303 = v_50 & v_301;
assign v_304 = v_303;
assign v_306 = v_51 & v_304;
assign v_307 = v_306;
assign v_308 = ~v_300 & ~v_49;
assign v_309 = v_300 & v_49;
assign v_311 = ~v_300 & v_302;
assign v_312 = v_300 & v_50;
assign v_314 = ~v_300 & v_305;
assign v_315 = v_300 & v_51;
assign v_320 = ~v_317 & ~v_318 & ~v_319;
assign v_321 = v_52;
assign v_323 = v_53 & v_321;
assign v_324 = v_323;
assign v_326 = v_54 & v_324;
assign v_327 = v_326;
assign v_328 = ~v_300 & v_52;
assign v_329 = ~v_52 & v_300;
assign v_331 = ~v_300 & v_53;
assign v_332 = v_300 & v_322;
assign v_334 = ~v_300 & v_54;
assign v_335 = v_300 & v_325;
assign v_340 = ~v_337 & ~v_338 & ~v_339;
assign v_343 = ~v_341 & ~v_342 & v_320 & v_340;
assign v_345 = v_57;
assign v_347 = v_58 & v_345;
assign v_348 = v_347;
assign v_350 = v_59 & v_348;
assign v_351 = v_350;
assign v_352 = ~v_344 & ~v_57;
assign v_353 = v_344 & v_57;
assign v_355 = ~v_344 & v_346;
assign v_356 = v_344 & v_58;
assign v_358 = ~v_344 & v_349;
assign v_359 = v_344 & v_59;
assign v_364 = ~v_361 & ~v_362 & ~v_363;
assign v_365 = v_60;
assign v_367 = v_61 & v_365;
assign v_368 = v_367;
assign v_370 = v_62 & v_368;
assign v_371 = v_370;
assign v_372 = ~v_344 & v_60;
assign v_373 = ~v_60 & v_344;
assign v_375 = ~v_344 & v_61;
assign v_376 = v_344 & v_366;
assign v_378 = ~v_344 & v_62;
assign v_379 = v_344 & v_369;
assign v_384 = ~v_381 & ~v_382 & ~v_383;
assign v_387 = ~v_385 & ~v_386 & v_364 & v_384;
assign v_388 = v_255 & v_299 & v_343 & v_387;
assign v_392 = ~v_389 & ~v_390 & ~v_391;
assign v_396 = ~v_393 & ~v_394 & ~v_395;
assign v_399 = ~v_397 & ~v_398 & v_392 & v_396;
assign v_403 = ~v_400 & ~v_401 & ~v_402;
assign v_407 = ~v_404 & ~v_405 & ~v_406;
assign v_410 = ~v_408 & ~v_409 & v_403 & v_407;
assign v_414 = ~v_411 & ~v_412 & ~v_413;
assign v_418 = ~v_415 & ~v_416 & ~v_417;
assign v_421 = ~v_419 & ~v_420 & v_414 & v_418;
assign v_425 = ~v_422 & ~v_423 & ~v_424;
assign v_429 = ~v_426 & ~v_427 & ~v_428;
assign v_432 = ~v_430 & ~v_431 & v_425 & v_429;
assign v_434 = v_388 & v_433;
assign v_86 = v_84 | v_85;
assign v_89 = v_87 | v_88;
assign v_92 = v_90 | v_91;
assign v_106 = v_104 | v_105;
assign v_109 = v_107 | v_108;
assign v_112 = v_110 | v_111;
assign v_130 = v_128 | v_129;
assign v_133 = v_131 | v_132;
assign v_136 = v_134 | v_135;
assign v_150 = v_148 | v_149;
assign v_153 = v_151 | v_152;
assign v_156 = v_154 | v_155;
assign v_174 = v_172 | v_173;
assign v_177 = v_175 | v_176;
assign v_180 = v_178 | v_179;
assign v_194 = v_192 | v_193;
assign v_197 = v_195 | v_196;
assign v_200 = v_198 | v_199;
assign v_218 = v_216 | v_217;
assign v_221 = v_219 | v_220;
assign v_224 = v_222 | v_223;
assign v_238 = v_236 | v_237;
assign v_241 = v_239 | v_240;
assign v_244 = v_242 | v_243;
assign v_266 = v_264 | v_265;
assign v_269 = v_267 | v_268;
assign v_272 = v_270 | v_271;
assign v_286 = v_284 | v_285;
assign v_289 = v_287 | v_288;
assign v_292 = v_290 | v_291;
assign v_310 = v_308 | v_309;
assign v_313 = v_311 | v_312;
assign v_316 = v_314 | v_315;
assign v_330 = v_328 | v_329;
assign v_333 = v_331 | v_332;
assign v_336 = v_334 | v_335;
assign v_354 = v_352 | v_353;
assign v_357 = v_355 | v_356;
assign v_360 = v_358 | v_359;
assign v_374 = v_372 | v_373;
assign v_377 = v_375 | v_376;
assign v_380 = v_378 | v_379;
assign v_433 = v_399 | v_410 | v_421 | v_432;
assign v_76 = v_8 ^ v_7;
assign v_78 = v_77 ^ v_2;
assign v_81 = v_80 ^ v_3;
assign v_93 = v_86 ^ v_9;
assign v_94 = v_89 ^ v_10;
assign v_95 = v_92 ^ v_11;
assign v_98 = v_97 ^ v_5;
assign v_101 = v_100 ^ v_6;
assign v_113 = v_106 ^ v_12;
assign v_114 = v_109 ^ v_13;
assign v_115 = v_112 ^ v_14;
assign v_117 = ~v_15 ^ v_8;
assign v_118 = v_7 ^ v_16;
assign v_120 = v_16 ^ v_15;
assign v_122 = v_121 ^ v_10;
assign v_125 = v_124 ^ v_11;
assign v_137 = v_130 ^ v_17;
assign v_138 = v_133 ^ v_18;
assign v_139 = v_136 ^ v_19;
assign v_142 = v_141 ^ v_13;
assign v_145 = v_144 ^ v_14;
assign v_157 = v_150 ^ v_20;
assign v_158 = v_153 ^ v_21;
assign v_159 = v_156 ^ v_22;
assign v_161 = ~v_23 ^ v_16;
assign v_162 = v_15 ^ v_24;
assign v_164 = v_24 ^ v_23;
assign v_166 = v_165 ^ v_18;
assign v_169 = v_168 ^ v_19;
assign v_181 = v_174 ^ v_25;
assign v_182 = v_177 ^ v_26;
assign v_183 = v_180 ^ v_27;
assign v_186 = v_185 ^ v_21;
assign v_189 = v_188 ^ v_22;
assign v_201 = v_194 ^ v_28;
assign v_202 = v_197 ^ v_29;
assign v_203 = v_200 ^ v_30;
assign v_205 = ~v_31 ^ v_24;
assign v_206 = v_23 ^ v_32;
assign v_208 = v_32 ^ v_31;
assign v_210 = v_209 ^ v_26;
assign v_213 = v_212 ^ v_27;
assign v_225 = v_218 ^ v_33;
assign v_226 = v_221 ^ v_34;
assign v_227 = v_224 ^ v_35;
assign v_230 = v_229 ^ v_29;
assign v_233 = v_232 ^ v_30;
assign v_245 = v_238 ^ v_36;
assign v_246 = v_241 ^ v_37;
assign v_247 = v_244 ^ v_38;
assign v_249 = ~v_39 ^ v_32;
assign v_250 = v_31 ^ v_40;
assign v_256 = v_48 ^ v_47;
assign v_258 = v_257 ^ v_42;
assign v_261 = v_260 ^ v_43;
assign v_273 = v_266 ^ v_49;
assign v_274 = v_269 ^ v_50;
assign v_275 = v_272 ^ v_51;
assign v_278 = v_277 ^ v_45;
assign v_281 = v_280 ^ v_46;
assign v_293 = v_286 ^ v_52;
assign v_294 = v_289 ^ v_53;
assign v_295 = v_292 ^ v_54;
assign v_297 = ~v_55 ^ v_48;
assign v_298 = v_47 ^ v_56;
assign v_300 = v_56 ^ v_55;
assign v_302 = v_301 ^ v_50;
assign v_305 = v_304 ^ v_51;
assign v_317 = v_310 ^ v_57;
assign v_318 = v_313 ^ v_58;
assign v_319 = v_316 ^ v_59;
assign v_322 = v_321 ^ v_53;
assign v_325 = v_324 ^ v_54;
assign v_337 = v_330 ^ v_60;
assign v_338 = v_333 ^ v_61;
assign v_339 = v_336 ^ v_62;
assign v_341 = ~v_63 ^ v_56;
assign v_342 = v_55 ^ v_64;
assign v_344 = v_64 ^ v_63;
assign v_346 = v_345 ^ v_58;
assign v_349 = v_348 ^ v_59;
assign v_361 = v_354 ^ v_65;
assign v_362 = v_357 ^ v_66;
assign v_363 = v_360 ^ v_67;
assign v_366 = v_365 ^ v_61;
assign v_369 = v_368 ^ v_62;
assign v_381 = v_374 ^ v_68;
assign v_382 = v_377 ^ v_69;
assign v_383 = v_380 ^ v_70;
assign v_385 = ~v_71 ^ v_64;
assign v_386 = v_63 ^ v_72;
assign v_389 = v_41 ^ v_33;
assign v_390 = v_42 ^ v_34;
assign v_391 = v_43 ^ v_35;
assign v_393 = v_44 ^ v_36;
assign v_394 = v_45 ^ v_37;
assign v_395 = v_46 ^ v_38;
assign v_397 = v_47 ^ v_39;
assign v_398 = v_48 ^ v_40;
assign v_400 = v_49 ^ v_33;
assign v_401 = v_50 ^ v_34;
assign v_402 = v_51 ^ v_35;
assign v_404 = v_52 ^ v_36;
assign v_405 = v_53 ^ v_37;
assign v_406 = v_54 ^ v_38;
assign v_408 = v_55 ^ v_39;
assign v_409 = v_56 ^ v_40;
assign v_411 = v_57 ^ v_33;
assign v_412 = v_58 ^ v_34;
assign v_413 = v_59 ^ v_35;
assign v_415 = v_60 ^ v_36;
assign v_416 = v_61 ^ v_37;
assign v_417 = v_62 ^ v_38;
assign v_419 = v_63 ^ v_39;
assign v_420 = v_64 ^ v_40;
assign v_422 = v_65 ^ v_33;
assign v_423 = v_66 ^ v_34;
assign v_424 = v_67 ^ v_35;
assign v_426 = v_68 ^ v_36;
assign v_427 = v_69 ^ v_37;
assign v_428 = v_70 ^ v_38;
assign v_430 = v_71 ^ v_39;
assign v_431 = v_72 ^ v_40;
assign x_1 = v_434 | ~v_252;
assign o_1 = x_1;
endmodule
