module formula(v_117,v_119,v_121,v_123,v_125,v_127,v_129,v_131,v_133,v_135,v_137,v_139,v_141,v_143,v_145,v_147,v_149,v_151,v_153,v_155,v_157,v_159,v_161,v_163,v_165,v_167,v_169,v_171,v_173,v_175,v_177,v_179,v_180,v_181,v_182,v_183,v_184,v_185,v_186,v_187,v_188,v_189,v_190,v_191,v_192,v_193,v_194,v_195,v_196,v_197,v_198,v_199,v_200,v_201,v_202,v_203,v_204,v_205,v_206,v_207,v_208,v_209,v_210,v_211,v_116,v_118,v_120,v_122,v_124,v_126,v_128,v_130,v_132,v_134,v_136,v_138,v_140,v_142,v_144,v_146,v_148,v_150,v_152,v_154,v_156,v_158,v_160,v_162,v_164,v_166,v_168,v_170,v_172,v_174,v_176,v_178,v_7,v_8,v_9,v_10,v_11,v_12,v_13,v_14,v_15,v_16,v_17,v_18,v_19,v_20,v_21,v_22,v_23,v_24,v_25,v_26,v_27,v_28,v_29,v_30,v_31,v_32,v_33,v_34,v_35,v_36,v_37,v_38,v_39,v_40,v_41,v_42,v_43,v_44,v_45,v_46,v_49,v_50,v_51,v_52,v_53,v_54,v_55,v_56,v_57,v_58,v_59,v_60,v_61,v_62,v_63,v_64,v_65,v_66,v_67,v_68,v_69,v_70,v_71,v_72,v_73,v_74,v_75,v_76,v_77,v_78,v_79,v_80,v_81,v_82,v_83,v_84,v_85,v_86,v_87,v_88,v_99,v_110,o_1);
	input v_117;
	v_119;
	v_121;
	v_123;
	v_125;
	v_127;
	v_129;
	v_131;
	v_133;
	v_135;
	v_137;
	v_139;
	v_141;
	v_143;
	v_145;
	v_147;
	v_149;
	v_151;
	v_153;
	v_155;
	v_157;
	v_159;
	v_161;
	v_163;
	v_165;
	v_167;
	v_169;
	v_171;
	v_173;
	v_175;
	v_177;
	v_179;
	v_180;
	v_181;
	v_182;
	v_183;
	v_184;
	v_185;
	v_186;
	v_187;
	v_188;
	v_189;
	v_190;
	v_191;
	v_192;
	v_193;
	v_194;
	v_195;
	v_196;
	v_197;
	v_198;
	v_199;
	v_200;
	v_201;
	v_202;
	v_203;
	v_204;
	v_205;
	v_206;
	v_207;
	v_208;
	v_209;
	v_210;
	v_211;
	v_116;
	v_118;
	v_120;
	v_122;
	v_124;
	v_126;
	v_128;
	v_130;
	v_132;
	v_134;
	v_136;
	v_138;
	v_140;
	v_142;
	v_144;
	v_146;
	v_148;
	v_150;
	v_152;
	v_154;
	v_156;
	v_158;
	v_160;
	v_162;
	v_164;
	v_166;
	v_168;
	v_170;
	v_172;
	v_174;
	v_176;
	v_178;
	v_7;
	v_8;
	v_9;
	v_10;
	v_11;
	v_12;
	v_13;
	v_14;
	v_15;
	v_16;
	v_17;
	v_18;
	v_19;
	v_20;
	v_21;
	v_22;
	v_23;
	v_24;
	v_25;
	v_26;
	v_27;
	v_28;
	v_29;
	v_30;
	v_31;
	v_32;
	v_33;
	v_34;
	v_35;
	v_36;
	v_37;
	v_38;
	v_39;
	v_40;
	v_41;
	v_42;
	v_43;
	v_44;
	v_45;
	v_46;
	v_49;
	v_50;
	v_51;
	v_52;
	v_53;
	v_54;
	v_55;
	v_56;
	v_57;
	v_58;
	v_59;
	v_60;
	v_61;
	v_62;
	v_63;
	v_64;
	v_65;
	v_66;
	v_67;
	v_68;
	v_69;
	v_70;
	v_71;
	v_72;
	v_73;
	v_74;
	v_75;
	v_76;
	v_77;
	v_78;
	v_79;
	v_80;
	v_81;
	v_82;
	v_83;
	v_84;
	v_85;
	v_86;
	v_87;
	v_88;
	v_99;
	v_110;
	wire v_1;
	wire v_2;
	wire v_3;
	wire v_4;
	wire v_5;
	wire v_6;
	wire v_47;
	wire v_48;
	wire v_89;
	wire v_90;
	wire v_91;
	wire v_92;
	wire v_93;
	wire v_94;
	wire v_95;
	wire v_96;
	wire v_97;
	wire v_98;
	wire v_100;
	wire v_101;
	wire v_102;
	wire v_103;
	wire v_104;
	wire v_105;
	wire v_106;
	wire v_107;
	wire v_108;
	wire v_109;
	wire v_111;
	wire v_112;
	wire v_113;
	wire v_114;
	wire v_115;
	wire v_212;
	wire x_1;
	wire x_2;
	wire x_3;
	wire x_4;
	wire x_5;
	wire x_6;
	wire x_7;
	wire x_8;
	wire x_9;
	wire x_10;
	wire x_11;
	wire x_12;
	wire x_13;
	wire x_14;
	wire x_15;
	wire x_16;
	wire x_17;
	wire x_18;
	wire x_19;
	wire x_20;
	wire x_21;
	wire x_22;
	wire x_23;
	wire x_24;
	wire x_25;
	wire x_26;
	wire x_27;
	wire x_28;
	wire x_29;
	wire x_30;
	wire x_31;
	wire x_32;
	wire x_33;
	wire x_34;
	wire x_35;
	wire x_36;
	wire x_37;
	wire x_38;
	wire x_39;
	wire x_40;
	wire x_41;
	wire x_42;
	wire x_43;
	wire x_44;
	wire x_45;
	wire x_46;
	wire x_47;
	wire x_48;
	wire x_49;
	wire x_50;
	wire x_51;
	wire x_52;
	wire x_53;
	wire x_54;
	wire x_55;
	wire x_56;
	wire x_57;
	wire x_58;
	wire x_59;
	wire x_60;
	wire x_61;
	wire x_62;
	wire x_63;
	wire x_64;
	wire x_65;
	wire x_66;
	wire x_67;
	wire x_68;
	wire x_69;
	wire x_70;
	wire x_71;
	wire x_72;
	wire x_73;
	wire x_74;
	wire x_75;
	wire x_76;
	wire x_77;
	wire x_78;
	wire x_79;
	wire x_80;
	wire x_81;
	wire x_82;
	wire x_83;
	wire x_84;
	wire x_85;
	wire x_86;
	wire x_87;
	wire x_88;
	wire x_89;
	wire x_90;
	wire x_91;
	wire x_92;
	wire x_93;
	wire x_94;
	wire x_95;
	wire x_96;
	wire x_97;
	wire x_98;
	wire x_99;
	wire x_100;
	wire x_101;
	wire x_102;
	wire x_103;
	wire x_104;
	wire x_105;
	wire x_106;
	wire x_107;
	wire x_108;
	wire x_109;
	wire x_110;
	wire x_111;
	wire x_112;
	wire x_113;
	wire x_114;
	wire x_115;
	wire x_116;
	wire x_117;
	wire x_118;
	wire x_119;
	wire x_120;
	wire x_121;
	wire x_122;
	wire x_123;
	wire x_124;
	wire x_125;
	wire x_126;
	wire x_127;
	wire x_128;
	wire x_129;
	wire x_130;
	wire x_131;
	wire x_132;
	wire x_133;
	wire x_134;
	wire x_135;
	wire x_136;
	wire x_137;
	wire x_138;
	wire x_139;
	wire x_140;
	wire x_141;
	wire x_142;
	wire x_143;
	wire x_144;
	wire x_145;
	wire x_146;
	wire x_147;
	wire x_148;
	wire x_149;
	wire x_150;
	wire x_151;
	wire x_152;
	wire x_153;
	wire x_154;
	wire x_155;
	wire x_156;
	wire x_157;
	wire x_158;
	wire x_159;
	wire x_160;
	wire x_161;
	wire x_162;
	wire x_163;
	wire x_164;
	wire x_165;
	wire x_166;
	wire x_167;
	wire x_168;
	wire x_169;
	wire x_170;
	wire x_171;
	wire x_172;
	wire x_173;
	wire x_174;
	wire x_175;
	wire x_176;
	wire x_177;
	wire x_178;
	wire x_179;
	wire x_180;
	wire x_181;
	wire x_182;
	wire x_183;
	wire x_184;
	wire x_185;
	wire x_186;
	wire x_187;
	wire x_188;
	wire x_189;
	wire x_190;
	wire x_191;
	wire x_192;
	wire x_193;
	wire x_194;
	wire x_195;
	wire x_196;
	wire x_197;
	wire x_198;
	wire x_199;
	wire x_200;
	wire x_201;
	wire x_202;
	wire x_203;
	wire x_204;
	wire x_205;
	wire x_206;
	wire x_207;
	wire x_208;
	wire x_209;
	wire x_210;
	wire x_211;
	wire x_212;
	wire x_213;
	wire x_214;
	wire x_215;
	wire x_216;
	wire x_217;
	wire x_218;
	wire x_219;
	wire x_220;
	wire x_221;
	wire x_222;
	wire x_223;
	wire x_224;
	wire x_225;
	wire x_226;
	wire x_227;
	wire x_228;
	wire x_229;
	wire x_230;
	wire x_231;
	wire x_232;
	wire x_233;
	wire x_234;
	wire x_235;
	wire x_236;
	wire x_237;
	wire x_238;
	wire x_239;
	wire x_240;
	wire x_241;
	wire x_242;
	wire x_243;
	wire x_244;
	wire x_245;
	wire x_246;
	wire x_247;
	wire x_248;
	wire x_249;
	wire x_250;
	wire x_251;
	wire x_252;
	wire x_253;
	wire x_254;
	wire x_255;
	wire x_256;
	wire x_257;
	wire x_258;
	wire x_259;
	wire x_260;
	wire x_261;
	wire x_262;
	wire x_263;
	wire x_264;
	wire x_265;
	wire x_266;
	wire x_267;
	wire x_268;
	wire x_269;
	wire x_270;
	wire x_271;
	wire x_272;
	wire x_273;
	wire x_274;
	wire x_275;
	wire x_276;
	wire x_277;
	wire x_278;
	wire x_279;
	wire x_280;
	wire x_281;
	wire x_282;
	wire x_283;
	wire x_284;
	wire x_285;
	wire x_286;
	wire x_287;
	wire x_288;
	wire x_289;
	wire x_290;
	wire x_291;
	wire x_292;
	wire x_293;
	wire x_294;
	wire x_295;
	wire x_296;
	wire x_297;
	wire x_298;
	wire x_299;
	wire x_300;
	wire x_301;
	wire x_302;
	wire x_303;
	wire x_304;
	wire x_305;
	wire x_306;
	wire x_307;
	wire x_308;
	wire x_309;
	wire x_310;
	wire x_311;
	wire x_312;
	wire x_313;
	wire x_314;
	wire x_315;
	wire x_316;
	wire x_317;
	wire x_318;
	wire x_319;
	wire x_320;
	wire x_321;
	wire x_322;
	wire x_323;
	wire x_324;
	wire x_325;
	wire x_326;
	wire x_327;
	wire x_328;
	wire x_329;
	wire x_330;
	wire x_331;
	wire x_332;
	wire x_333;
	wire x_334;
	wire x_335;
	wire x_336;
	wire x_337;
	wire x_338;
	wire x_339;
	wire x_340;
	wire x_341;
	wire x_342;
	wire x_343;
	wire x_344;
	wire x_345;
	wire x_346;
	wire x_347;
	wire x_348;
	wire x_349;
	wire x_350;
	wire x_351;
	wire x_352;
	wire x_353;
	wire x_354;
	wire x_355;
	wire x_356;
	wire x_357;
	wire x_358;
	wire x_359;
	wire x_360;
	wire x_361;
	wire x_362;
	wire x_363;
	wire x_364;
	wire x_365;
	wire x_366;
	wire x_367;
	wire x_368;
	wire x_369;
	wire x_370;
	wire x_371;
	wire x_372;
	wire x_373;
	wire x_374;
	wire x_375;
	wire x_376;
	wire x_377;
	wire x_378;
	wire x_379;
	wire x_380;
	wire x_381;
	wire x_382;
	wire x_383;
	wire x_384;
	wire x_385;
	wire x_386;
	wire x_387;
	wire x_388;
	wire x_389;
	wire x_390;
	wire x_391;
	wire x_392;
	wire x_393;
	wire x_394;
	wire x_395;
	wire x_396;
	wire x_397;
	wire x_398;
	wire x_399;
	wire x_400;
	wire x_401;
	wire x_402;
	wire x_403;
	wire x_404;
	wire x_405;
	wire x_406;
	wire x_407;
	wire x_408;
	wire x_409;
	wire x_410;
	wire x_411;
	wire x_412;
	wire x_413;
	wire x_414;
	wire x_415;
	wire x_416;
	wire x_417;
	wire x_418;
	wire x_419;
	wire x_420;
	wire x_421;
	wire x_422;
	wire x_423;
	wire x_424;
	wire x_425;
	wire x_426;
	wire x_427;
	wire x_428;
	wire x_429;
	wire x_430;
	wire x_431;
	wire x_432;
	wire x_433;
	wire x_434;
	wire x_435;
	wire x_436;
	wire x_437;
	wire x_438;
	wire x_439;
	wire x_440;
	wire x_441;
	wire x_442;
	wire x_443;
	wire x_444;
	wire x_445;
	wire x_446;
	wire x_447;
	wire x_448;
	wire x_449;
	wire x_450;
	wire x_451;
	wire x_452;
	wire x_453;
	wire x_454;
	wire x_455;
	wire x_456;
	wire x_457;
	wire x_458;
	wire x_459;
	wire x_460;
	wire x_461;
	wire x_462;
	wire x_463;
	wire x_464;
	wire x_465;
	wire x_466;
	wire x_467;
	wire x_468;
	wire x_469;
	wire x_470;
	wire x_471;
	wire x_472;
	wire x_473;
	wire x_474;
	wire x_475;
	wire x_476;
	wire x_477;
	wire x_478;
	wire x_479;
	wire x_480;
	wire x_481;
	wire x_482;
	wire x_483;
	wire x_484;
	wire x_485;
	wire x_486;
	wire x_487;
	wire x_488;
	wire x_489;
	wire x_490;
	wire x_491;
	wire x_492;
	wire x_493;
	wire x_494;
	wire x_495;
	wire x_496;
	wire x_497;
	wire x_498;
	wire x_499;
	wire x_500;
	wire x_501;
	wire x_502;
	wire x_503;
	wire x_504;
	wire x_505;
	wire x_506;
	wire x_507;
	wire x_508;
	wire x_509;
	wire x_510;
	wire x_511;
	wire x_512;
	wire x_513;
	wire x_514;
	wire x_515;
	wire x_516;
	wire x_517;
	wire x_518;
	wire x_519;
	wire x_520;
	wire x_521;
	wire x_522;
	wire x_523;
	wire x_524;
	wire x_525;
	wire x_526;
	wire x_527;
	wire x_528;
	wire x_529;
	wire x_530;
	wire x_531;
	wire x_532;
	wire x_533;
	wire x_534;
	wire x_535;
	wire x_536;
	wire x_537;
	wire x_538;
	wire x_539;
	wire x_540;
	wire x_541;
	wire x_542;
	wire x_543;
	wire x_544;
	wire x_545;
	wire x_546;
	wire x_547;
	wire x_548;
	wire x_549;
	wire x_550;
	wire x_551;
	wire x_552;
	wire x_553;
	wire x_554;
	wire x_555;
	wire x_556;
	wire x_557;
	wire x_558;
	wire x_559;
	wire x_560;
	wire x_561;
	wire x_562;
	wire x_563;
	wire x_564;
	wire x_565;
	wire x_566;
	wire x_567;
	wire x_568;
	wire x_569;
	wire x_570;
	wire x_571;
	wire x_572;
	wire x_573;
	wire x_574;
	wire x_575;
	wire x_576;
	wire x_577;
	wire x_578;
	wire x_579;
	wire x_580;
	wire x_581;
	wire x_582;
	wire x_583;
	wire x_584;
	wire x_585;
	wire x_586;
	wire x_587;
	wire x_588;
	wire x_589;
	wire x_590;
	wire x_591;
	wire x_592;
	wire x_593;
	wire x_594;
	wire x_595;
	wire x_596;
	wire x_597;
	wire x_598;
	wire x_599;
	wire x_600;
	wire x_601;
	wire x_602;
	wire x_603;
	wire x_604;
	wire x_605;
	wire x_606;
	wire x_607;
	wire x_608;
	wire x_609;
	wire x_610;
	wire x_611;
	wire x_612;
	wire x_613;
	wire x_614;
	wire x_615;
	wire x_616;
	wire x_617;
	wire x_618;
	wire x_619;
	wire x_620;
	wire x_621;
	wire x_622;
	wire x_623;
	wire x_624;
	wire x_625;
	wire x_626;
	wire x_627;
	wire x_628;
	wire x_629;
	wire x_630;
	wire x_631;
	wire x_632;
	wire x_633;
	wire x_634;
	wire x_635;
	wire x_636;
	wire x_637;
	wire x_638;
	wire x_639;
	wire x_640;
	wire x_641;
	wire x_642;
	wire x_643;
	wire x_644;
	wire x_645;
	wire x_646;
	wire x_647;
	wire x_648;
	wire x_649;
	wire x_650;
	wire x_651;
	wire x_652;
	wire x_653;
	wire x_654;
	wire x_655;
	wire x_656;
	wire x_657;
	wire x_658;
	wire x_659;
	wire x_660;
	wire x_661;
	wire x_662;
	wire x_663;
	wire x_664;
	wire x_665;
	wire x_666;
	wire x_667;
	wire x_668;
	wire x_669;
	wire x_670;
	wire x_671;
	wire x_672;
	wire x_673;
	wire x_674;
	wire x_675;
	wire x_676;
	wire x_677;
	wire x_678;
	wire x_679;
	wire x_680;
	wire x_681;
	wire x_682;
	wire x_683;
	wire x_684;
	wire x_685;
	wire x_686;
	wire x_687;
	wire x_688;
	wire x_689;
	wire x_690;
	wire x_691;
	wire x_692;
	wire x_693;
	wire x_694;
	wire x_695;
	wire x_696;
	wire x_697;
	wire x_698;
	wire x_699;
	wire x_700;
	wire x_701;
	wire x_702;
	wire x_703;
	wire x_704;
	wire x_705;
	wire x_706;
	wire x_707;
	wire x_708;
	wire x_709;
	wire x_710;
	wire x_711;
	wire x_712;
	wire x_713;
	wire x_714;
	wire x_715;
	wire x_716;
	wire x_717;
	wire x_718;
	wire x_719;
	wire x_720;
	wire x_721;
	wire x_722;
	wire x_723;
	wire x_724;
	wire x_725;
	wire x_726;
	wire x_727;
	wire x_728;
	wire x_729;
	wire x_730;
	wire x_731;
	wire x_732;
	wire x_733;
	wire x_734;
	wire x_735;
	wire x_736;
	wire x_737;
	wire x_738;
	wire x_739;
	wire x_740;
	wire x_741;
	wire x_742;
	wire x_743;
	wire x_744;
	wire x_745;
	wire x_746;
	wire x_747;
	wire x_748;
	wire x_749;
	wire x_750;
	wire x_751;
	wire x_752;
	wire x_753;
	wire x_754;
	wire x_755;
	wire x_756;
	wire x_757;
	wire x_758;
	wire x_759;
	wire x_760;
	wire x_761;
	wire x_762;
	wire x_763;
	wire x_764;
	wire x_765;
	wire x_766;
	wire x_767;
	wire x_768;
	wire x_769;
	wire x_770;
	wire x_771;
	wire x_772;
	wire x_773;
	wire x_774;
	wire x_775;
	wire x_776;
	wire x_777;
	wire x_778;
	wire x_779;
	wire x_780;
	wire x_781;
	wire x_782;
	wire x_783;
	wire x_784;
	wire x_785;
	wire x_786;
	wire x_787;
	wire x_788;
	wire x_789;
	wire x_790;
	wire x_791;
	wire x_792;
	wire x_793;
	wire x_794;
	wire x_795;
	wire x_796;
	wire x_797;
	wire x_798;
	wire x_799;
	wire x_800;
	wire x_801;
	wire x_802;
	wire x_803;
	wire x_804;
	wire x_805;
	wire x_806;
	wire x_807;
	wire x_808;
	wire x_809;
	wire x_810;
	wire x_811;
	wire x_812;
	wire x_813;
	wire x_814;
	wire x_815;
	wire x_816;
	wire x_817;
	wire x_818;
	wire x_819;
	wire x_820;
	wire x_821;
	wire x_822;
	wire x_823;
	wire x_824;
	wire x_825;
	wire x_826;
	wire x_827;
	wire x_828;
	wire x_829;
	wire x_830;
	wire x_831;
	wire x_832;
	wire x_833;
	wire x_834;
	wire x_835;
	wire x_836;
	wire x_837;
	wire x_838;
	wire x_839;
	wire x_840;
	wire x_841;
	wire x_842;
	wire x_843;
	wire x_844;
	wire x_845;
	wire x_846;
	wire x_847;
	wire x_848;
	wire x_849;
	wire x_850;
	wire x_851;
	wire x_852;
	wire x_853;
	wire x_854;
	wire x_855;
	wire x_856;
	wire x_857;
	wire x_858;
	wire x_859;
	wire x_860;
	wire x_861;
	wire x_862;
	wire x_863;
	wire x_864;
	wire x_865;
	wire x_866;
	wire x_867;
	wire x_868;
	wire x_869;
	wire x_870;
	wire x_871;
	wire x_872;
	wire x_873;
	wire x_874;
	wire x_875;
	wire x_876;
	wire x_877;
	wire x_878;
	wire x_879;
	wire x_880;
	wire x_881;
	wire x_882;
	wire x_883;
	wire x_884;
	wire x_885;
	wire x_886;
	wire x_887;
	wire x_888;
	wire x_889;
	wire x_890;
	wire x_891;
	wire x_892;
	wire x_893;
	wire x_894;
	wire x_895;
	wire x_896;
	wire x_897;
	wire x_898;
	wire x_899;
	wire x_900;
	wire x_901;
	wire x_902;
	wire x_903;
	wire x_904;
	wire x_905;
	wire x_906;
	wire x_907;
	wire x_908;
	wire x_909;
	wire x_910;
	wire x_911;
	wire x_912;
	wire x_913;
	wire x_914;
	wire x_915;
	wire x_916;
	wire x_917;
	wire x_918;
	wire x_919;
	wire x_920;
	wire x_921;
	wire x_922;
	wire x_923;
	wire x_924;
	wire x_925;
	wire x_926;
	wire x_927;
	wire x_928;
	wire x_929;
	wire x_930;
	wire x_931;
	wire x_932;
	wire x_933;
	wire x_934;
	wire x_935;
	wire x_936;
	wire x_937;
	wire x_938;
	wire x_939;
	wire x_940;
	wire x_941;
	wire x_942;
	wire x_943;
	wire x_944;
	wire x_945;
	wire x_946;
	wire x_947;
	wire x_948;
	wire x_949;
	wire x_950;
	wire x_951;
	wire x_952;
	wire x_953;
	output o_1;
	assign v_6 = (v_116 & ~v_180);
	assign v_48 = (v_116 & ~v_117);
	assign x_464 = (~v_180 | v_116);
	assign x_463 = (~v_117 | v_116);
	assign v_111 = (~v_118 & v_181);
	assign v_100 = (~v_118 & v_119);
	assign x_57 = (((~v_17 | v_176)) | ~v_210);
	assign x_56 = (((~v_17 | v_178)) | ~v_211);
	assign x_55 = (((v_17 | v_210)) | v_211);
	assign x_54 = (((v_17 | ~v_176)) | ~v_178);
	assign x_53 = (((v_17 | ~v_176)) | v_211);
	assign x_52 = (((v_17 | ~v_178)) | v_210);
	assign x_63 = (((~v_18 | ~v_176)) | v_210);
	assign x_62 = (((~v_18 | ~v_174)) | v_209);
	assign x_61 = (((v_18 | v_176)) | ~v_209);
	assign x_59 = (((v_18 | ~v_209)) | ~v_210);
	assign x_58 = (((v_18 | v_174)) | v_176);
	assign x_51 = (((~v_16 | v_17)) | ~v_18);
	assign x_60 = (((v_18 | v_174)) | ~v_210);
	assign x_69 = (((~v_19 | v_172)) | ~v_208);
	assign x_68 = (((~v_19 | v_174)) | ~v_209);
	assign x_67 = (((v_19 | v_208)) | v_209);
	assign x_66 = (((v_19 | ~v_172)) | ~v_174);
	assign x_65 = (((v_19 | ~v_172)) | v_209);
	assign x_64 = (((v_19 | ~v_174)) | v_208);
	assign x_50 = (~v_16 | v_19);
	assign x_49 = (((v_16 | v_18)) | ~v_19);
	assign x_48 = (((v_16 | ~v_17)) | ~v_19);
	assign x_74 = (((~v_20 | ~v_170)) | v_207);
	assign x_73 = (((v_20 | v_172)) | ~v_207);
	assign x_72 = (((v_20 | v_170)) | ~v_208);
	assign x_71 = (((v_20 | ~v_207)) | ~v_208);
	assign x_70 = (((v_20 | v_170)) | v_172);
	assign x_75 = (((~v_20 | ~v_172)) | v_208);
	assign x_81 = (((~v_21 | v_168)) | ~v_206);
	assign x_80 = (((~v_21 | v_170)) | ~v_207);
	assign x_79 = (((v_21 | v_206)) | v_207);
	assign x_78 = (((v_21 | ~v_168)) | ~v_170);
	assign x_77 = (((v_21 | ~v_168)) | v_207);
	assign x_76 = (((v_21 | ~v_170)) | v_206);
	assign x_47 = (((~v_15 | v_20)) | ~v_21);
	assign x_46 = (((~v_15 | ~v_16)) | ~v_21);
	assign v_109 = (((((v_19 & v_20)) & v_21)) & v_22);
	assign x_87 = (((~v_22 | ~v_168)) | v_206);
	assign x_86 = (((~v_22 | ~v_166)) | v_205);
	assign x_85 = (((v_22 | v_168)) | ~v_205);
	assign x_84 = (((v_22 | v_166)) | ~v_206);
	assign x_83 = (((v_22 | ~v_205)) | ~v_206);
	assign x_82 = (((v_22 | v_166)) | v_168);
	assign x_44 = (((((v_15 | v_16)) | ~v_20)) | ~v_22);
	assign x_43 = (((v_15 | v_21)) | ~v_22);
	assign x_45 = (~v_15 | v_22);
	assign x_93 = (((~v_23 | v_164)) | ~v_204);
	assign x_92 = (((~v_23 | v_166)) | ~v_205);
	assign x_91 = (((v_23 | v_204)) | v_205);
	assign x_89 = (((v_23 | ~v_164)) | v_205);
	assign x_88 = (((v_23 | ~v_166)) | v_204);
	assign x_90 = (((v_23 | ~v_164)) | ~v_166);
	assign v_114 = (v_23 & v_24);
	assign x_99 = (((~v_24 | ~v_164)) | v_204);
	assign x_98 = (((~v_24 | ~v_162)) | v_203);
	assign x_97 = (((v_24 | v_164)) | ~v_203);
	assign x_96 = (((v_24 | v_162)) | ~v_204);
	assign x_95 = (((v_24 | ~v_203)) | ~v_204);
	assign x_94 = (((v_24 | v_162)) | v_164);
	assign x_42 = (((~v_14 | v_23)) | ~v_24);
	assign x_41 = (((~v_14 | ~v_15)) | ~v_24);
	assign x_104 = (((~v_25 | v_162)) | ~v_203);
	assign x_103 = (((v_25 | v_202)) | v_203);
	assign x_102 = (((v_25 | ~v_160)) | ~v_162);
	assign x_101 = (((v_25 | ~v_160)) | v_203);
	assign x_100 = (((v_25 | ~v_162)) | v_202);
	assign x_40 = (~v_14 | v_25);
	assign x_39 = (((((v_14 | v_15)) | ~v_23)) | ~v_25);
	assign x_38 = (((v_14 | v_24)) | ~v_25);
	assign x_105 = (((~v_25 | v_160)) | ~v_202);
	assign x_111 = (((~v_26 | ~v_160)) | v_202);
	assign x_110 = (((~v_26 | ~v_158)) | v_201);
	assign x_109 = (((v_26 | v_160)) | ~v_201);
	assign x_108 = (((v_26 | v_158)) | ~v_202);
	assign x_107 = (((v_26 | ~v_201)) | ~v_202);
	assign x_106 = (((v_26 | v_158)) | v_160);
	assign x_117 = (((~v_27 | v_156)) | ~v_200);
	assign x_116 = (((~v_27 | v_158)) | ~v_201);
	assign x_115 = (((v_27 | v_200)) | v_201);
	assign x_114 = (((v_27 | ~v_156)) | ~v_158);
	assign x_113 = (((v_27 | ~v_156)) | v_201);
	assign x_112 = (((v_27 | ~v_158)) | v_200);
	assign x_37 = (((~v_13 | v_26)) | ~v_27);
	assign x_36 = (((~v_13 | ~v_14)) | ~v_27);
	assign x_123 = (((~v_28 | ~v_156)) | v_200);
	assign x_122 = (((~v_28 | ~v_154)) | v_199);
	assign x_121 = (((v_28 | v_156)) | ~v_199);
	assign x_119 = (((v_28 | ~v_199)) | ~v_200);
	assign x_118 = (((v_28 | v_154)) | v_156);
	assign x_35 = (~v_13 | v_28);
	assign x_34 = (((((v_13 | v_14)) | ~v_26)) | ~v_28);
	assign x_33 = (((v_13 | v_27)) | ~v_28);
	assign x_120 = (((v_28 | v_154)) | ~v_200);
	assign x_129 = (((~v_29 | v_152)) | ~v_198);
	assign x_128 = (((~v_29 | v_154)) | ~v_199);
	assign x_126 = (((v_29 | ~v_152)) | ~v_154);
	assign x_125 = (((v_29 | ~v_152)) | v_199);
	assign x_124 = (((v_29 | ~v_154)) | v_198);
	assign x_127 = (((v_29 | v_198)) | v_199);
	assign v_113 = (((((v_27 & v_28)) & v_29)) & v_30);
	assign x_135 = (((~v_30 | ~v_152)) | v_198);
	assign x_133 = (((v_30 | v_152)) | ~v_197);
	assign x_132 = (((v_30 | v_150)) | ~v_198);
	assign x_131 = (((v_30 | ~v_197)) | ~v_198);
	assign x_130 = (((v_30 | v_150)) | v_152);
	assign x_32 = (((~v_12 | v_29)) | ~v_30);
	assign x_31 = (((~v_12 | ~v_13)) | ~v_30);
	assign x_134 = (((~v_30 | ~v_150)) | v_197);
	assign x_141 = (((~v_31 | v_148)) | ~v_196);
	assign x_140 = (((~v_31 | v_150)) | ~v_197);
	assign x_139 = (((v_31 | v_196)) | v_197);
	assign x_138 = (((v_31 | ~v_148)) | ~v_150);
	assign x_137 = (((v_31 | ~v_148)) | v_197);
	assign x_136 = (((v_31 | ~v_150)) | v_196);
	assign x_29 = (((((v_12 | v_13)) | ~v_29)) | ~v_31);
	assign x_28 = (((v_12 | v_30)) | ~v_31);
	assign x_30 = (~v_12 | v_31);
	assign x_147 = (((~v_32 | ~v_148)) | v_196);
	assign x_146 = (((~v_32 | ~v_146)) | v_195);
	assign x_145 = (((v_32 | v_148)) | ~v_195);
	assign x_144 = (((v_32 | v_146)) | ~v_196);
	assign x_143 = (((v_32 | ~v_195)) | ~v_196);
	assign x_142 = (((v_32 | v_146)) | v_148);
	assign x_153 = (((~v_33 | v_144)) | ~v_194);
	assign x_152 = (((~v_33 | v_146)) | ~v_195);
	assign x_151 = (((v_33 | v_194)) | v_195);
	assign x_150 = (((v_33 | ~v_144)) | ~v_146);
	assign x_148 = (((v_33 | ~v_146)) | v_194);
	assign x_27 = (((~v_11 | v_32)) | ~v_33);
	assign x_26 = (((~v_11 | ~v_12)) | ~v_33);
	assign x_149 = (((v_33 | ~v_144)) | v_195);
	assign v_105 = (((((v_31 & v_32)) & v_33)) & v_34);
	assign x_159 = (((~v_34 | ~v_144)) | v_194);
	assign x_158 = (((~v_34 | ~v_142)) | v_193);
	assign x_157 = (((v_34 | v_144)) | ~v_193);
	assign x_156 = (((v_34 | v_142)) | ~v_194);
	assign x_155 = (((v_34 | ~v_193)) | ~v_194);
	assign x_154 = (((v_34 | v_142)) | v_144);
	assign x_25 = (~v_11 | v_34);
	assign x_24 = (((((v_11 | v_12)) | ~v_32)) | ~v_34);
	assign x_23 = (((v_11 | v_33)) | ~v_34);
	assign x_165 = (((~v_35 | v_140)) | ~v_192);
	assign x_163 = (((v_35 | v_192)) | v_193);
	assign x_162 = (((v_35 | ~v_140)) | ~v_142);
	assign x_161 = (((v_35 | ~v_140)) | v_193);
	assign x_160 = (((v_35 | ~v_142)) | v_192);
	assign x_164 = (((~v_35 | v_142)) | ~v_193);
	assign x_171 = (((~v_36 | ~v_140)) | v_192);
	assign x_170 = (((~v_36 | ~v_138)) | v_191);
	assign x_169 = (((v_36 | v_140)) | ~v_191);
	assign x_168 = (((v_36 | v_138)) | ~v_192);
	assign x_167 = (((v_36 | ~v_191)) | ~v_192);
	assign x_166 = (((v_36 | v_138)) | v_140);
	assign x_22 = (((~v_10 | v_35)) | ~v_36);
	assign x_21 = (((~v_10 | ~v_11)) | ~v_36);
	assign x_177 = (((~v_37 | v_136)) | ~v_190);
	assign x_176 = (((~v_37 | v_138)) | ~v_191);
	assign x_175 = (((v_37 | v_190)) | v_191);
	assign x_174 = (((v_37 | ~v_136)) | ~v_138);
	assign x_173 = (((v_37 | ~v_136)) | v_191);
	assign x_172 = (((v_37 | ~v_138)) | v_190);
	assign x_20 = (~v_10 | v_37);
	assign x_19 = (((((v_10 | v_11)) | ~v_35)) | ~v_37);
	assign x_18 = (((v_10 | v_36)) | ~v_37);
	assign v_104 = (((((v_35 & v_36)) & v_37)) & v_38);
	assign x_183 = (((~v_38 | ~v_136)) | v_190);
	assign x_182 = (((~v_38 | ~v_134)) | v_189);
	assign x_181 = (((v_38 | v_136)) | ~v_189);
	assign x_180 = (((v_38 | v_134)) | ~v_190);
	assign x_178 = (((v_38 | v_134)) | v_136);
	assign x_179 = (((v_38 | ~v_189)) | ~v_190);
	assign x_189 = (((~v_39 | v_132)) | ~v_188);
	assign x_188 = (((~v_39 | v_134)) | ~v_189);
	assign x_187 = (((v_39 | v_188)) | v_189);
	assign x_186 = (((v_39 | ~v_132)) | ~v_134);
	assign x_185 = (((v_39 | ~v_132)) | v_189);
	assign x_184 = (((v_39 | ~v_134)) | v_188);
	assign x_17 = (((~v_9 | v_38)) | ~v_39);
	assign x_16 = (((~v_9 | ~v_10)) | ~v_39);
	assign x_195 = (((~v_40 | ~v_132)) | v_188);
	assign x_193 = (((v_40 | v_132)) | ~v_187);
	assign x_192 = (((v_40 | v_130)) | ~v_188);
	assign x_191 = (((v_40 | ~v_187)) | ~v_188);
	assign x_190 = (((v_40 | v_130)) | v_132);
	assign x_14 = (((((v_9 | v_10)) | ~v_38)) | ~v_40);
	assign x_13 = (((v_9 | v_39)) | ~v_40);
	assign x_194 = (((~v_40 | ~v_130)) | v_187);
	assign x_15 = (~v_9 | v_40);
	assign x_201 = (((~v_41 | v_128)) | ~v_186);
	assign x_200 = (((~v_41 | v_130)) | ~v_187);
	assign x_199 = (((v_41 | v_186)) | v_187);
	assign x_198 = (((v_41 | ~v_128)) | ~v_130);
	assign x_197 = (((v_41 | ~v_128)) | v_187);
	assign x_196 = (((v_41 | ~v_130)) | v_186);
	assign v_107 = (((((v_39 & v_40)) & v_41)) & v_42);
	assign x_207 = (((~v_42 | ~v_128)) | v_186);
	assign x_206 = (((~v_42 | ~v_126)) | v_185);
	assign x_205 = (((v_42 | v_128)) | ~v_185);
	assign x_204 = (((v_42 | v_126)) | ~v_186);
	assign x_203 = (((v_42 | ~v_185)) | ~v_186);
	assign x_202 = (((v_42 | v_126)) | v_128);
	assign x_12 = (((~v_8 | v_41)) | ~v_42);
	assign x_11 = (((~v_8 | ~v_9)) | ~v_42);
	assign x_213 = (((~v_43 | v_124)) | ~v_184);
	assign x_212 = (((~v_43 | v_126)) | ~v_185);
	assign x_211 = (((v_43 | v_184)) | v_185);
	assign x_210 = (((v_43 | ~v_124)) | ~v_126);
	assign x_208 = (((v_43 | ~v_126)) | v_184);
	assign x_10 = (~v_8 | v_43);
	assign x_9 = (((((v_8 | v_9)) | ~v_41)) | ~v_43);
	assign x_209 = (((v_43 | ~v_124)) | v_185);
	assign x_8 = (((v_8 | v_42)) | ~v_43);
	assign x_219 = (((~v_44 | ~v_124)) | v_184);
	assign x_218 = (((~v_44 | ~v_122)) | v_183);
	assign x_217 = (((v_44 | v_124)) | ~v_183);
	assign x_216 = (((v_44 | v_122)) | ~v_184);
	assign x_215 = (((v_44 | ~v_183)) | ~v_184);
	assign x_214 = (((v_44 | v_122)) | v_124);
	assign x_225 = (((~v_45 | v_120)) | ~v_182);
	assign x_223 = (((v_45 | v_182)) | v_183);
	assign x_222 = (((v_45 | ~v_120)) | ~v_122);
	assign x_221 = (((v_45 | ~v_120)) | v_183);
	assign x_220 = (((v_45 | ~v_122)) | v_182);
	assign x_7 = (((~v_7 | v_44)) | ~v_45);
	assign x_6 = (((~v_7 | ~v_8)) | ~v_45);
	assign x_224 = (((~v_45 | v_122)) | ~v_183);
	assign v_106 = (((((v_43 & v_44)) & v_45)) & v_46);
	assign x_231 = (((~v_46 | ~v_120)) | v_182);
	assign x_230 = (((~v_46 | ~v_118)) | v_181);
	assign x_229 = (((v_46 | v_120)) | ~v_181);
	assign x_228 = (((v_46 | v_118)) | ~v_182);
	assign x_227 = (((v_46 | ~v_181)) | ~v_182);
	assign x_226 = (((v_46 | v_118)) | v_120);
	assign x_5 = (~v_7 | v_46);
	assign x_4 = (((((v_7 | v_8)) | ~v_44)) | ~v_46);
	assign x_3 = (((v_7 | v_45)) | ~v_46);
	assign x_288 = (((~v_59 | v_178)) | ~v_179);
	assign x_287 = (((~v_59 | v_176)) | ~v_177);
	assign x_286 = (((v_59 | ~v_176)) | ~v_178);
	assign x_285 = (((v_59 | v_177)) | v_179);
	assign x_284 = (((v_59 | v_177)) | ~v_178);
	assign x_283 = (((v_59 | ~v_176)) | v_179);
	assign x_294 = (((~v_60 | ~v_176)) | v_177);
	assign x_293 = (((~v_60 | ~v_174)) | v_175);
	assign x_292 = (((v_60 | ~v_175)) | ~v_177);
	assign x_291 = (((v_60 | v_174)) | v_176);
	assign x_290 = (((v_60 | v_174)) | ~v_177);
	assign x_289 = (((v_60 | ~v_175)) | v_176);
	assign x_282 = (((~v_58 | v_59)) | ~v_60);
	assign x_300 = (((~v_61 | v_174)) | ~v_175);
	assign x_299 = (((~v_61 | v_172)) | ~v_173);
	assign x_297 = (((v_61 | v_173)) | v_175);
	assign x_296 = (((v_61 | v_173)) | ~v_174);
	assign x_295 = (((v_61 | ~v_172)) | v_175);
	assign x_281 = (~v_58 | v_61);
	assign x_280 = (((v_58 | v_60)) | ~v_61);
	assign x_279 = (((v_58 | ~v_59)) | ~v_61);
	assign x_298 = (((v_61 | ~v_172)) | ~v_174);
	assign x_306 = (((~v_62 | ~v_172)) | v_173);
	assign x_305 = (((~v_62 | ~v_170)) | v_171);
	assign x_304 = (((v_62 | ~v_171)) | ~v_173);
	assign x_303 = (((v_62 | v_170)) | v_172);
	assign x_302 = (((v_62 | v_170)) | ~v_173);
	assign x_301 = (((v_62 | ~v_171)) | v_172);
	assign x_312 = (((~v_63 | v_170)) | ~v_171);
	assign x_311 = (((~v_63 | v_168)) | ~v_169);
	assign x_310 = (((v_63 | ~v_168)) | ~v_170);
	assign x_309 = (((v_63 | v_169)) | v_171);
	assign x_308 = (((v_63 | v_169)) | ~v_170);
	assign x_307 = (((v_63 | ~v_168)) | v_171);
	assign x_278 = (((~v_57 | v_62)) | ~v_63);
	assign x_277 = (((~v_57 | ~v_58)) | ~v_63);
	assign v_98 = (((((v_61 & v_62)) & v_63)) & v_64);
	assign x_318 = (((~v_64 | ~v_168)) | v_169);
	assign x_317 = (((~v_64 | ~v_166)) | v_167);
	assign x_316 = (((v_64 | ~v_167)) | ~v_169);
	assign x_315 = (((v_64 | v_166)) | v_168);
	assign x_314 = (((v_64 | v_166)) | ~v_169);
	assign x_276 = (~v_57 | v_64);
	assign x_275 = (((((v_57 | v_58)) | ~v_62)) | ~v_64);
	assign x_274 = (((v_57 | v_63)) | ~v_64);
	assign x_313 = (((v_64 | ~v_167)) | v_168);
	assign x_324 = (((~v_65 | v_166)) | ~v_167);
	assign x_323 = (((~v_65 | v_164)) | ~v_165);
	assign x_322 = (((v_65 | ~v_164)) | ~v_166);
	assign x_321 = (((v_65 | v_165)) | v_167);
	assign x_320 = (((v_65 | v_165)) | ~v_166);
	assign x_319 = (((v_65 | ~v_164)) | v_167);
	assign x_330 = (((~v_66 | ~v_164)) | v_165);
	assign x_329 = (((~v_66 | ~v_162)) | v_163);
	assign x_327 = (((v_66 | v_162)) | v_164);
	assign x_326 = (((v_66 | v_162)) | ~v_165);
	assign x_325 = (((v_66 | ~v_163)) | v_164);
	assign x_273 = (((~v_56 | v_65)) | ~v_66);
	assign x_272 = (((~v_56 | ~v_57)) | ~v_66);
	assign x_328 = (((v_66 | ~v_163)) | ~v_165);
	assign x_336 = (((~v_67 | v_162)) | ~v_163);
	assign x_335 = (((~v_67 | v_160)) | ~v_161);
	assign x_334 = (((v_67 | ~v_160)) | ~v_162);
	assign x_333 = (((v_67 | v_161)) | v_163);
	assign x_332 = (((v_67 | v_161)) | ~v_162);
	assign x_331 = (((v_67 | ~v_160)) | v_163);
	assign x_271 = (~v_56 | v_67);
	assign x_270 = (((((v_56 | v_57)) | ~v_65)) | ~v_67);
	assign x_269 = (((v_56 | v_66)) | ~v_67);
	assign v_102 = (((((v_65 & v_66)) & v_67)) & v_68);
	assign x_342 = (((~v_68 | ~v_160)) | v_161);
	assign x_341 = (((~v_68 | ~v_158)) | v_159);
	assign x_340 = (((v_68 | ~v_159)) | ~v_161);
	assign x_339 = (((v_68 | v_158)) | v_160);
	assign x_338 = (((v_68 | v_158)) | ~v_161);
	assign x_337 = (((v_68 | ~v_159)) | v_160);
	assign x_348 = (((~v_69 | v_158)) | ~v_159);
	assign x_347 = (((~v_69 | v_156)) | ~v_157);
	assign x_346 = (((v_69 | ~v_156)) | ~v_158);
	assign x_345 = (((v_69 | v_157)) | v_159);
	assign x_344 = (((v_69 | v_157)) | ~v_158);
	assign x_267 = (((~v_55 | ~v_56)) | ~v_69);
	assign x_343 = (((v_69 | ~v_156)) | v_159);
	assign x_268 = (((~v_55 | v_68)) | ~v_69);
	assign x_354 = (((~v_70 | ~v_156)) | v_157);
	assign x_353 = (((~v_70 | ~v_154)) | v_155);
	assign x_352 = (((v_70 | ~v_155)) | ~v_157);
	assign x_351 = (((v_70 | v_154)) | v_156);
	assign x_350 = (((v_70 | v_154)) | ~v_157);
	assign x_349 = (((v_70 | ~v_155)) | v_156);
	assign x_266 = (~v_55 | v_70);
	assign x_265 = (((((v_55 | v_56)) | ~v_68)) | ~v_70);
	assign x_264 = (((v_55 | v_69)) | ~v_70);
	assign x_360 = (((~v_71 | v_154)) | ~v_155);
	assign x_359 = (((~v_71 | v_152)) | ~v_153);
	assign x_357 = (((v_71 | v_153)) | v_155);
	assign x_356 = (((v_71 | v_153)) | ~v_154);
	assign x_355 = (((v_71 | ~v_152)) | v_155);
	assign x_358 = (((v_71 | ~v_152)) | ~v_154);
	assign v_101 = (((((v_69 & v_70)) & v_71)) & v_72);
	assign x_366 = (((~v_72 | ~v_152)) | v_153);
	assign x_365 = (((~v_72 | ~v_150)) | v_151);
	assign x_364 = (((v_72 | ~v_151)) | ~v_153);
	assign x_363 = (((v_72 | v_150)) | v_152);
	assign x_362 = (((v_72 | v_150)) | ~v_153);
	assign x_361 = (((v_72 | ~v_151)) | v_152);
	assign x_263 = (((~v_54 | v_71)) | ~v_72);
	assign x_262 = (((~v_54 | ~v_55)) | ~v_72);
	assign x_372 = (((~v_73 | v_150)) | ~v_151);
	assign x_371 = (((~v_73 | v_148)) | ~v_149);
	assign x_370 = (((v_73 | ~v_148)) | ~v_150);
	assign x_369 = (((v_73 | v_149)) | v_151);
	assign x_368 = (((v_73 | v_149)) | ~v_150);
	assign x_367 = (((v_73 | ~v_148)) | v_151);
	assign x_261 = (~v_54 | v_73);
	assign x_260 = (((((v_54 | v_55)) | ~v_71)) | ~v_73);
	assign x_259 = (((v_54 | v_72)) | ~v_73);
	assign x_378 = (((~v_74 | ~v_148)) | v_149);
	assign x_377 = (((~v_74 | ~v_146)) | v_147);
	assign x_376 = (((v_74 | ~v_147)) | ~v_149);
	assign x_375 = (((v_74 | v_146)) | v_148);
	assign x_374 = (((v_74 | v_146)) | ~v_149);
	assign x_373 = (((v_74 | ~v_147)) | v_148);
	assign x_384 = (((~v_75 | v_146)) | ~v_147);
	assign x_383 = (((~v_75 | v_144)) | ~v_145);
	assign x_382 = (((v_75 | ~v_144)) | ~v_146);
	assign x_381 = (((v_75 | v_145)) | v_147);
	assign x_380 = (((v_75 | v_145)) | ~v_146);
	assign x_379 = (((v_75 | ~v_144)) | v_147);
	assign x_258 = (((~v_53 | v_74)) | ~v_75);
	assign x_257 = (((~v_53 | ~v_54)) | ~v_75);
	assign v_94 = (((((v_73 & v_74)) & v_75)) & v_76);
	assign x_390 = (((~v_76 | ~v_144)) | v_145);
	assign x_389 = (((~v_76 | ~v_142)) | v_143);
	assign x_387 = (((v_76 | v_142)) | v_144);
	assign x_386 = (((v_76 | v_142)) | ~v_145);
	assign x_385 = (((v_76 | ~v_143)) | v_144);
	assign x_256 = (~v_53 | v_76);
	assign x_255 = (((((v_53 | v_54)) | ~v_74)) | ~v_76);
	assign x_254 = (((v_53 | v_75)) | ~v_76);
	assign x_388 = (((v_76 | ~v_143)) | ~v_145);
	assign x_396 = (((~v_77 | v_142)) | ~v_143);
	assign x_395 = (((~v_77 | v_140)) | ~v_141);
	assign x_394 = (((v_77 | ~v_140)) | ~v_142);
	assign x_393 = (((v_77 | v_141)) | v_143);
	assign x_392 = (((v_77 | v_141)) | ~v_142);
	assign x_391 = (((v_77 | ~v_140)) | v_143);
	assign x_402 = (((~v_78 | ~v_140)) | v_141);
	assign x_401 = (((~v_78 | ~v_138)) | v_139);
	assign x_400 = (((v_78 | ~v_139)) | ~v_141);
	assign x_399 = (((v_78 | v_138)) | v_140);
	assign x_398 = (((v_78 | v_138)) | ~v_141);
	assign x_397 = (((v_78 | ~v_139)) | v_140);
	assign x_252 = (((~v_52 | ~v_53)) | ~v_78);
	assign x_253 = (((~v_52 | v_77)) | ~v_78);
	assign x_408 = (((~v_79 | v_138)) | ~v_139);
	assign x_407 = (((~v_79 | v_136)) | ~v_137);
	assign x_406 = (((v_79 | ~v_136)) | ~v_138);
	assign x_405 = (((v_79 | v_137)) | v_139);
	assign x_404 = (((v_79 | v_137)) | ~v_138);
	assign x_251 = (~v_52 | v_79);
	assign x_250 = (((((v_52 | v_53)) | ~v_77)) | ~v_79);
	assign x_249 = (((v_52 | v_78)) | ~v_79);
	assign x_403 = (((v_79 | ~v_136)) | v_139);
	assign v_93 = (((((v_77 & v_78)) & v_79)) & v_80);
	assign x_414 = (((~v_80 | ~v_136)) | v_137);
	assign x_413 = (((~v_80 | ~v_134)) | v_135);
	assign x_412 = (((v_80 | ~v_135)) | ~v_137);
	assign x_411 = (((v_80 | v_134)) | v_136);
	assign x_410 = (((v_80 | v_134)) | ~v_137);
	assign x_409 = (((v_80 | ~v_135)) | v_136);
	assign x_420 = (((~v_81 | v_134)) | ~v_135);
	assign x_419 = (((~v_81 | v_132)) | ~v_133);
	assign x_417 = (((v_81 | v_133)) | v_135);
	assign x_416 = (((v_81 | v_133)) | ~v_134);
	assign x_415 = (((v_81 | ~v_132)) | v_135);
	assign x_248 = (((~v_51 | v_80)) | ~v_81);
	assign x_247 = (((~v_51 | ~v_52)) | ~v_81);
	assign x_418 = (((v_81 | ~v_132)) | ~v_134);
	assign x_426 = (((~v_82 | ~v_132)) | v_133);
	assign x_425 = (((~v_82 | ~v_130)) | v_131);
	assign x_424 = (((v_82 | ~v_131)) | ~v_133);
	assign x_423 = (((v_82 | v_130)) | v_132);
	assign x_422 = (((v_82 | v_130)) | ~v_133);
	assign x_421 = (((v_82 | ~v_131)) | v_132);
	assign x_245 = (((((v_51 | v_52)) | ~v_80)) | ~v_82);
	assign x_244 = (((v_51 | v_81)) | ~v_82);
	assign x_246 = (~v_51 | v_82);
	assign x_432 = (((~v_83 | v_130)) | ~v_131);
	assign x_431 = (((~v_83 | v_128)) | ~v_129);
	assign x_430 = (((v_83 | ~v_128)) | ~v_130);
	assign x_429 = (((v_83 | v_129)) | v_131);
	assign x_428 = (((v_83 | v_129)) | ~v_130);
	assign x_427 = (((v_83 | ~v_128)) | v_131);
	assign v_96 = (((((v_81 & v_82)) & v_83)) & v_84);
	assign x_438 = (((~v_84 | ~v_128)) | v_129);
	assign x_437 = (((~v_84 | ~v_126)) | v_127);
	assign x_436 = (((v_84 | ~v_127)) | ~v_129);
	assign x_435 = (((v_84 | v_126)) | v_128);
	assign x_434 = (((v_84 | v_126)) | ~v_129);
	assign x_243 = (((~v_50 | v_83)) | ~v_84);
	assign x_242 = (((~v_50 | ~v_51)) | ~v_84);
	assign x_433 = (((v_84 | ~v_127)) | v_128);
	assign x_444 = (((~v_85 | v_126)) | ~v_127);
	assign x_443 = (((~v_85 | v_124)) | ~v_125);
	assign x_442 = (((v_85 | ~v_124)) | ~v_126);
	assign x_441 = (((v_85 | v_125)) | v_127);
	assign x_440 = (((v_85 | v_125)) | ~v_126);
	assign x_439 = (((v_85 | ~v_124)) | v_127);
	assign x_241 = (~v_50 | v_85);
	assign x_240 = (((((v_50 | v_51)) | ~v_83)) | ~v_85);
	assign x_239 = (((v_50 | v_84)) | ~v_85);
	assign x_450 = (((~v_86 | ~v_124)) | v_125);
	assign x_449 = (((~v_86 | ~v_122)) | v_123);
	assign x_447 = (((v_86 | v_122)) | v_124);
	assign x_446 = (((v_86 | v_122)) | ~v_125);
	assign x_445 = (((v_86 | ~v_123)) | v_124);
	assign x_448 = (((v_86 | ~v_123)) | ~v_125);
	assign x_456 = (((~v_87 | v_122)) | ~v_123);
	assign x_455 = (((~v_87 | v_120)) | ~v_121);
	assign x_454 = (((v_87 | ~v_120)) | ~v_122);
	assign x_453 = (((v_87 | v_121)) | v_123);
	assign x_452 = (((v_87 | v_121)) | ~v_122);
	assign x_451 = (((v_87 | ~v_120)) | v_123);
	assign x_238 = (((~v_49 | v_86)) | ~v_87);
	assign x_237 = (((~v_49 | ~v_50)) | ~v_87);
	assign v_95 = (((((v_85 & v_86)) & v_87)) & v_88);
	assign x_462 = (((~v_88 | ~v_120)) | v_121);
	assign x_461 = (((~v_88 | ~v_118)) | v_119);
	assign x_460 = (((v_88 | ~v_119)) | ~v_121);
	assign x_459 = (((v_88 | v_118)) | v_120);
	assign x_458 = (((v_88 | v_118)) | ~v_121);
	assign x_457 = (((v_88 | ~v_119)) | v_120);
	assign x_236 = (~v_49 | v_88);
	assign x_235 = (((((v_49 | v_50)) | ~v_86)) | ~v_88);
	assign x_234 = (((v_49 | v_87)) | ~v_88);
	assign x_472 = (((~v_99 | ~v_178)) | v_179);
	assign x_477 = (((~v_110 | ~v_178)) | v_211);
	assign x_476 = (~v_110 | ~v_6);
	assign x_2 = (((v_6 | v_118)) | ~v_181);
	assign x_1 = (~v_7 | v_6);
	assign x_471 = (~v_99 | ~v_48);
	assign x_233 = (((v_48 | v_118)) | ~v_119);
	assign x_232 = (~v_49 | v_48);
	assign x_475 = (~v_110 | ~v_111);
	assign x_474 = (((((v_110 | ~v_211)) | v_6)) | v_111);
	assign x_473 = (((((v_110 | v_178)) | v_6)) | v_111);
	assign x_470 = (~v_99 | ~v_100);
	assign x_469 = (((((v_99 | ~v_179)) | v_48)) | v_100);
	assign x_468 = (((((v_99 | v_178)) | v_48)) | v_100);
	assign x_529 = (x_56 & x_57);
	assign x_527 = (x_54 & x_55);
	assign x_526 = (x_52 & x_53);
	assign x_536 = (x_61 & x_62);
	assign x_530 = (x_58 & x_59);
	assign x_542 = (x_67 & x_68);
	assign x_539 = (x_65 & x_66);
	assign x_538 = (x_63 & x_64);
	assign x_523 = (x_50 & x_51);
	assign x_522 = (x_48 & x_49);
	assign x_546 = (x_73 & x_74);
	assign x_545 = (x_71 & x_72);
	assign x_543 = (x_69 & x_70);
	assign x_553 = (x_80 & x_81);
	assign x_552 = (x_78 & x_79);
	assign x_550 = (x_76 & x_77);
	assign x_520 = (x_46 & x_47);
	assign v_108 = (((((v_17 & v_18)) & v_109)) & v_110);
	assign x_559 = (x_86 & x_87);
	assign x_557 = (x_84 & x_85);
	assign x_556 = (x_82 & x_83);
	assign x_516 = (x_43 & x_44);
	assign x_565 = (x_91 & x_92);
	assign x_560 = (x_88 & x_89);
	assign x_571 = (x_97 & x_98);
	assign x_568 = (x_95 & x_96);
	assign x_567 = (x_93 & x_94);
	assign x_515 = (x_41 & x_42);
	assign x_575 = (x_103 & x_104);
	assign x_574 = (x_101 & x_102);
	assign x_572 = (x_99 & x_100);
	assign x_513 = (x_39 & x_40);
	assign x_582 = (x_110 & x_111);
	assign x_581 = (x_108 & x_109);
	assign x_579 = (x_106 & x_107);
	assign x_588 = (x_116 & x_117);
	assign x_586 = (x_114 & x_115);
	assign x_585 = (x_112 & x_113);
	assign x_512 = (x_37 & x_38);
	assign x_596 = (x_121 & x_122);
	assign x_589 = (x_118 & x_119);
	assign x_509 = (x_35 & x_36);
	assign x_508 = (x_33 & x_34);
	assign x_602 = (x_128 & x_129);
	assign x_599 = (x_125 & x_126);
	assign x_598 = (x_123 & x_124);
	assign v_112 = (((((v_25 & v_26)) & v_113)) & v_114);
	assign x_605 = (x_132 & x_133);
	assign x_604 = (x_130 & x_131);
	assign x_506 = (x_31 & x_32);
	assign x_612 = (x_139 & x_140);
	assign x_611 = (x_137 & x_138);
	assign x_609 = (x_135 & x_136);
	assign x_501 = (x_28 & x_29);
	assign x_618 = (x_145 & x_146);
	assign x_616 = (x_143 & x_144);
	assign x_615 = (x_141 & x_142);
	assign x_626 = (x_152 & x_153);
	assign x_624 = (x_150 & x_151);
	assign x_619 = (x_147 & x_148);
	assign x_500 = (x_26 & x_27);
	assign x_631 = (x_158 & x_159);
	assign x_630 = (x_156 & x_157);
	assign x_627 = (x_154 & x_155);
	assign x_498 = (x_24 & x_25);
	assign x_634 = (x_162 & x_163);
	assign x_633 = (x_160 & x_161);
	assign x_641 = (x_169 & x_170);
	assign x_640 = (x_167 & x_168);
	assign x_638 = (x_165 & x_166);
	assign x_497 = (x_22 & x_23);
	assign x_647 = (x_175 & x_176);
	assign x_645 = (x_173 & x_174);
	assign x_644 = (x_171 & x_172);
	assign x_494 = (x_20 & x_21);
	assign x_493 = (x_18 & x_19);
	assign x_656 = (x_182 & x_183);
	assign x_654 = (x_180 & x_181);
	assign x_648 = (x_177 & x_178);
	assign x_661 = (x_188 & x_189);
	assign x_660 = (x_186 & x_187);
	assign x_657 = (x_184 & x_185);
	assign x_491 = (x_16 & x_17);
	assign x_664 = (x_192 & x_193);
	assign x_663 = (x_190 & x_191);
	assign x_487 = (x_13 & x_14);
	assign x_671 = (x_199 & x_200);
	assign x_670 = (x_197 & x_198);
	assign x_668 = (x_195 & x_196);
	assign x_677 = (x_205 & x_206);
	assign x_675 = (x_203 & x_204);
	assign x_674 = (x_201 & x_202);
	assign x_486 = (x_11 & x_12);
	assign x_685 = (x_212 & x_213);
	assign x_683 = (x_210 & x_211);
	assign x_678 = (x_207 & x_208);
	assign x_484 = (x_9 & x_10);
	assign x_690 = (x_218 & x_219);
	assign x_689 = (x_216 & x_217);
	assign x_686 = (x_214 & x_215);
	assign x_693 = (x_222 & x_223);
	assign x_692 = (x_220 & x_221);
	assign x_481 = (x_6 & x_7);
	assign v_103 = (((((v_104 & v_105)) & v_106)) & v_107);
	assign x_700 = (x_229 & x_230);
	assign x_699 = (x_227 & x_228);
	assign x_697 = (x_225 & x_226);
	assign x_480 = (x_4 & x_5);
	assign x_759 = (x_286 & x_287);
	assign x_757 = (x_284 & x_285);
	assign x_764 = (x_292 & x_293);
	assign x_763 = (x_290 & x_291);
	assign x_760 = (x_288 & x_289);
	assign x_773 = (x_299 & x_300);
	assign x_767 = (x_296 & x_297);
	assign x_766 = (x_294 & x_295);
	assign x_753 = (x_281 & x_282);
	assign x_752 = (x_279 & x_280);
	assign x_779 = (x_305 & x_306);
	assign x_776 = (x_303 & x_304);
	assign x_775 = (x_301 & x_302);
	assign x_783 = (x_311 & x_312);
	assign x_782 = (x_309 & x_310);
	assign x_780 = (x_307 & x_308);
	assign x_750 = (x_277 & x_278);
	assign v_97 = (((((v_59 & v_60)) & v_98)) & v_99);
	assign x_789 = (x_316 & x_317);
	assign x_787 = (x_314 & x_315);
	assign x_749 = (x_275 & x_276);
	assign x_794 = (x_322 & x_323);
	assign x_793 = (x_320 & x_321);
	assign x_790 = (x_318 & x_319);
	assign x_802 = (x_329 & x_330);
	assign x_797 = (x_326 & x_327);
	assign x_796 = (x_324 & x_325);
	assign x_746 = (x_273 & x_274);
	assign x_808 = (x_335 & x_336);
	assign x_805 = (x_333 & x_334);
	assign x_804 = (x_331 & x_332);
	assign x_745 = (x_271 & x_272);
	assign x_743 = (x_269 & x_270);
	assign x_812 = (x_341 & x_342);
	assign x_811 = (x_339 & x_340);
	assign x_809 = (x_337 & x_338);
	assign x_818 = (x_346 & x_347);
	assign x_816 = (x_344 & x_345);
	assign x_823 = (x_352 & x_353);
	assign x_822 = (x_350 & x_351);
	assign x_819 = (x_348 & x_349);
	assign x_738 = (x_266 & x_267);
	assign x_737 = (x_264 & x_265);
	assign x_833 = (x_359 & x_360);
	assign x_826 = (x_356 & x_357);
	assign x_825 = (x_354 & x_355);
	assign x_839 = (x_365 & x_366);
	assign x_836 = (x_363 & x_364);
	assign x_835 = (x_361 & x_362);
	assign x_735 = (x_262 & x_263);
	assign x_843 = (x_371 & x_372);
	assign x_842 = (x_369 & x_370);
	assign x_840 = (x_367 & x_368);
	assign x_734 = (x_260 & x_261);
	assign x_849 = (x_376 & x_377);
	assign x_847 = (x_374 & x_375);
	assign x_854 = (x_382 & x_383);
	assign x_853 = (x_380 & x_381);
	assign x_850 = (x_378 & x_379);
	assign x_731 = (x_258 & x_259);
	assign x_862 = (x_389 & x_390);
	assign x_857 = (x_386 & x_387);
	assign x_856 = (x_384 & x_385);
	assign x_730 = (x_256 & x_257);
	assign x_728 = (x_254 & x_255);
	assign x_868 = (x_395 & x_396);
	assign x_865 = (x_393 & x_394);
	assign x_864 = (x_391 & x_392);
	assign x_872 = (x_401 & x_402);
	assign x_871 = (x_399 & x_400);
	assign x_869 = (x_397 & x_398);
	assign x_878 = (x_406 & x_407);
	assign x_876 = (x_404 & x_405);
	assign x_724 = (x_251 & x_252);
	assign x_723 = (x_249 & x_250);
	assign x_883 = (x_412 & x_413);
	assign x_882 = (x_410 & x_411);
	assign x_879 = (x_408 & x_409);
	assign x_892 = (x_419 & x_420);
	assign x_886 = (x_416 & x_417);
	assign x_885 = (x_414 & x_415);
	assign x_721 = (x_247 & x_248);
	assign x_898 = (x_425 & x_426);
	assign x_895 = (x_423 & x_424);
	assign x_894 = (x_421 & x_422);
	assign x_718 = (x_244 & x_245);
	assign x_902 = (x_431 & x_432);
	assign x_901 = (x_429 & x_430);
	assign x_899 = (x_427 & x_428);
	assign x_908 = (x_436 & x_437);
	assign x_906 = (x_434 & x_435);
	assign x_717 = (x_242 & x_243);
	assign x_913 = (x_442 & x_443);
	assign x_912 = (x_440 & x_441);
	assign x_909 = (x_438 & x_439);
	assign x_715 = (x_240 & x_241);
	assign x_921 = (x_449 & x_450);
	assign x_916 = (x_446 & x_447);
	assign x_915 = (x_444 & x_445);
	assign x_927 = (x_455 & x_456);
	assign x_924 = (x_453 & x_454);
	assign x_923 = (x_451 & x_452);
	assign x_707 = (x_237 & x_238);
	assign v_92 = (((((v_93 & v_94)) & v_95)) & v_96);
	assign x_931 = (x_461 & x_462);
	assign x_930 = (x_459 & x_460);
	assign x_928 = (x_457 & x_458);
	assign x_706 = (x_235 & x_236);
	assign x_945 = (x_476 & x_477);
	assign x_478 = (x_2 & x_3);
	assign x_704 = (x_233 & x_234);
	assign x_703 = (x_231 & x_232);
	assign x_944 = (x_474 & x_475);
	assign x_942 = (x_472 & x_473);
	assign x_941 = (x_470 & x_471);
	assign x_938 = (x_468 & x_469);
	assign x_528 = (x_526 & x_527);
	assign x_537 = (x_60 & x_536);
	assign x_531 = (x_529 & x_530);
	assign x_540 = (x_538 & x_539);
	assign x_524 = (x_522 & x_523);
	assign x_547 = (x_545 & x_546);
	assign x_544 = (x_542 & x_543);
	assign x_554 = (x_552 & x_553);
	assign x_551 = (x_75 & x_550);
	assign x_521 = (x_45 & x_520);
	assign x_558 = (x_556 & x_557);
	assign x_566 = (x_90 & x_565);
	assign x_561 = (x_559 & x_560);
	assign x_569 = (x_567 & x_568);
	assign x_517 = (x_515 & x_516);
	assign x_576 = (x_574 & x_575);
	assign x_573 = (x_571 & x_572);
	assign x_583 = (x_581 & x_582);
	assign x_580 = (x_105 & x_579);
	assign x_587 = (x_585 & x_586);
	assign x_514 = (x_512 & x_513);
	assign x_597 = (x_120 & x_596);
	assign x_590 = (x_588 & x_589);
	assign x_510 = (x_508 & x_509);
	assign x_603 = (x_127 & x_602);
	assign x_600 = (x_598 & x_599);
	assign x_606 = (x_604 & x_605);
	assign x_507 = (x_30 & x_506);
	assign x_613 = (x_611 & x_612);
	assign x_610 = (x_134 & x_609);
	assign x_617 = (x_615 & x_616);
	assign x_625 = (x_149 & x_624);
	assign x_620 = (x_618 & x_619);
	assign x_502 = (x_500 & x_501);
	assign x_632 = (x_630 & x_631);
	assign x_628 = (x_626 & x_627);
	assign x_635 = (x_633 & x_634);
	assign x_642 = (x_640 & x_641);
	assign x_639 = (x_164 & x_638);
	assign x_499 = (x_497 & x_498);
	assign x_646 = (x_644 & x_645);
	assign x_495 = (x_493 & x_494);
	assign x_655 = (x_179 & x_654);
	assign x_649 = (x_647 & x_648);
	assign x_662 = (x_660 & x_661);
	assign x_658 = (x_656 & x_657);
	assign x_492 = (x_15 & x_491);
	assign x_665 = (x_663 & x_664);
	assign x_672 = (x_670 & x_671);
	assign x_669 = (x_194 & x_668);
	assign x_676 = (x_674 & x_675);
	assign x_488 = (x_486 & x_487);
	assign x_684 = (x_209 & x_683);
	assign x_679 = (x_677 & x_678);
	assign x_485 = (x_8 & x_484);
	assign x_691 = (x_689 & x_690);
	assign x_687 = (x_685 & x_686);
	assign x_694 = (x_692 & x_693);
	assign x_701 = (x_699 & x_700);
	assign x_698 = (x_224 & x_697);
	assign x_482 = (x_480 & x_481);
	assign x_758 = (x_283 & x_757);
	assign x_765 = (x_763 & x_764);
	assign x_761 = (x_759 & x_760);
	assign x_774 = (x_298 & x_773);
	assign x_768 = (x_766 & x_767);
	assign x_754 = (x_752 & x_753);
	assign x_777 = (x_775 & x_776);
	assign x_784 = (x_782 & x_783);
	assign x_781 = (x_779 & x_780);
	assign x_788 = (x_313 & x_787);
	assign x_751 = (x_749 & x_750);
	assign x_795 = (x_793 & x_794);
	assign x_791 = (x_789 & x_790);
	assign x_803 = (x_328 & x_802);
	assign x_798 = (x_796 & x_797);
	assign x_806 = (x_804 & x_805);
	assign x_747 = (x_745 & x_746);
	assign x_744 = (x_268 & x_743);
	assign x_813 = (x_811 & x_812);
	assign x_810 = (x_808 & x_809);
	assign x_817 = (x_343 & x_816);
	assign x_824 = (x_822 & x_823);
	assign x_820 = (x_818 & x_819);
	assign x_739 = (x_737 & x_738);
	assign x_834 = (x_358 & x_833);
	assign x_827 = (x_825 & x_826);
	assign x_837 = (x_835 & x_836);
	assign x_844 = (x_842 & x_843);
	assign x_841 = (x_839 & x_840);
	assign x_736 = (x_734 & x_735);
	assign x_848 = (x_373 & x_847);
	assign x_855 = (x_853 & x_854);
	assign x_851 = (x_849 & x_850);
	assign x_863 = (x_388 & x_862);
	assign x_858 = (x_856 & x_857);
	assign x_732 = (x_730 & x_731);
	assign x_729 = (x_253 & x_728);
	assign x_866 = (x_864 & x_865);
	assign x_873 = (x_871 & x_872);
	assign x_870 = (x_868 & x_869);
	assign x_877 = (x_403 & x_876);
	assign x_725 = (x_723 & x_724);
	assign x_884 = (x_882 & x_883);
	assign x_880 = (x_878 & x_879);
	assign x_893 = (x_418 & x_892);
	assign x_887 = (x_885 & x_886);
	assign x_722 = (x_246 & x_721);
	assign x_896 = (x_894 & x_895);
	assign x_903 = (x_901 & x_902);
	assign x_900 = (x_898 & x_899);
	assign x_907 = (x_433 & x_906);
	assign x_719 = (x_717 & x_718);
	assign x_914 = (x_912 & x_913);
	assign x_910 = (x_908 & x_909);
	assign x_716 = (x_239 & x_715);
	assign x_922 = (x_448 & x_921);
	assign x_917 = (x_915 & x_916);
	assign x_925 = (x_923 & x_924);
	assign v_91 = (((((v_92 & v_97)) & v_101)) & v_102);
	assign x_932 = (x_930 & x_931);
	assign x_929 = (x_927 & x_928);
	assign x_708 = (x_706 & x_707);
	assign x_479 = (x_1 & x_478);
	assign x_705 = (x_703 & x_704);
	assign x_946 = (x_944 & x_945);
	assign x_943 = (x_941 & x_942);
	assign x_532 = (x_528 & x_531);
	assign x_541 = (x_537 & x_540);
	assign x_548 = (x_544 & x_547);
	assign x_555 = (x_551 & x_554);
	assign x_525 = (x_521 & x_524);
	assign x_562 = (x_558 & x_561);
	assign x_570 = (x_566 & x_569);
	assign x_577 = (x_573 & x_576);
	assign x_584 = (x_580 & x_583);
	assign x_518 = (x_514 & x_517);
	assign x_591 = (x_587 & x_590);
	assign x_601 = (x_597 & x_600);
	assign x_607 = (x_603 & x_606);
	assign x_511 = (x_507 & x_510);
	assign x_614 = (x_610 & x_613);
	assign x_621 = (x_617 & x_620);
	assign x_629 = (x_625 & x_628);
	assign x_636 = (x_632 & x_635);
	assign x_643 = (x_639 & x_642);
	assign x_503 = (x_499 & x_502);
	assign x_650 = (x_646 & x_649);
	assign x_659 = (x_655 & x_658);
	assign x_496 = (x_492 & x_495);
	assign x_666 = (x_662 & x_665);
	assign x_673 = (x_669 & x_672);
	assign x_680 = (x_676 & x_679);
	assign x_489 = (x_485 & x_488);
	assign x_688 = (x_684 & x_687);
	assign x_695 = (x_691 & x_694);
	assign x_702 = (x_698 & x_701);
	assign x_762 = (x_758 & x_761);
	assign x_769 = (x_765 & x_768);
	assign x_778 = (x_774 & x_777);
	assign x_785 = (x_781 & x_784);
	assign x_755 = (x_751 & x_754);
	assign x_792 = (x_788 & x_791);
	assign x_799 = (x_795 & x_798);
	assign x_807 = (x_803 & x_806);
	assign x_748 = (x_744 & x_747);
	assign x_814 = (x_810 & x_813);
	assign x_821 = (x_817 & x_820);
	assign x_828 = (x_824 & x_827);
	assign x_838 = (x_834 & x_837);
	assign x_845 = (x_841 & x_844);
	assign x_740 = (x_736 & x_739);
	assign x_852 = (x_848 & x_851);
	assign x_859 = (x_855 & x_858);
	assign x_733 = (x_729 & x_732);
	assign x_867 = (x_863 & x_866);
	assign x_874 = (x_870 & x_873);
	assign x_881 = (x_877 & x_880);
	assign x_888 = (x_884 & x_887);
	assign x_726 = (x_722 & x_725);
	assign x_897 = (x_893 & x_896);
	assign x_904 = (x_900 & x_903);
	assign x_911 = (x_907 & x_910);
	assign x_720 = (x_716 & x_719);
	assign x_918 = (x_914 & x_917);
	assign x_926 = (x_922 & x_925);
	assign x_467 = (v_112 | v_91);
	assign x_466 = (v_103 | v_91);
	assign x_465 = (v_108 | v_91);
	assign x_933 = (x_929 & x_932);
	assign x_483 = (x_479 & x_482);
	assign x_709 = (x_705 & x_708);
	assign x_947 = (x_943 & x_946);
	assign x_549 = (x_541 & x_548);
	assign x_533 = (x_525 & x_532);
	assign x_563 = (x_555 & x_562);
	assign x_578 = (x_570 & x_577);
	assign x_592 = (x_584 & x_591);
	assign x_608 = (x_601 & x_607);
	assign x_519 = (x_511 & x_518);
	assign x_622 = (x_614 & x_621);
	assign x_637 = (x_629 & x_636);
	assign x_651 = (x_643 & x_650);
	assign x_504 = (x_496 & x_503);
	assign x_667 = (x_659 & x_666);
	assign x_681 = (x_673 & x_680);
	assign x_696 = (x_688 & x_695);
	assign x_770 = (x_762 & x_769);
	assign x_786 = (x_778 & x_785);
	assign x_800 = (x_792 & x_799);
	assign x_756 = (x_748 & x_755);
	assign x_815 = (x_807 & x_814);
	assign x_829 = (x_821 & x_828);
	assign x_846 = (x_838 & x_845);
	assign x_860 = (x_852 & x_859);
	assign x_741 = (x_733 & x_740);
	assign x_875 = (x_867 & x_874);
	assign x_889 = (x_881 & x_888);
	assign x_905 = (x_897 & x_904);
	assign x_727 = (x_720 & x_726);
	assign x_919 = (x_911 & x_918);
	assign x_937 = (x_466 & x_467);
	assign x_935 = (x_464 & x_465);
	assign x_934 = (x_926 & x_933);
	assign x_490 = (x_483 & x_489);
	assign x_710 = (x_702 & x_709);
	assign x_564 = (x_549 & x_563);
	assign x_593 = (x_578 & x_592);
	assign x_534 = (x_519 & x_533);
	assign x_623 = (x_608 & x_622);
	assign x_652 = (x_637 & x_651);
	assign x_682 = (x_667 & x_681);
	assign x_801 = (x_786 & x_800);
	assign x_771 = (x_756 & x_770);
	assign x_830 = (x_815 & x_829);
	assign x_861 = (x_846 & x_860);
	assign x_890 = (x_875 & x_889);
	assign x_742 = (x_727 & x_741);
	assign x_920 = (x_905 & x_919);
	assign x_939 = (x_937 & x_938);
	assign x_936 = (x_463 & x_935);
	assign x_505 = (x_490 & x_504);
	assign x_711 = (x_696 & x_710);
	assign x_594 = (x_564 & x_593);
	assign x_653 = (x_623 & x_652);
	assign x_831 = (x_801 & x_830);
	assign x_891 = (x_861 & x_890);
	assign x_772 = (x_742 & x_771);
	assign x_940 = (x_936 & x_939);
	assign x_535 = (x_505 & x_534);
	assign x_712 = (x_682 & x_711);
	assign x_832 = (x_772 & x_831);
	assign x_948 = (x_940 & x_947);
	assign x_595 = (x_535 & x_594);
	assign x_713 = (x_653 & x_712);
	assign x_949 = (x_934 & x_948);
	assign x_714 = (x_595 & x_713);
	assign x_950 = (x_920 & x_949);
	assign x_951 = (x_891 & x_950);
	assign x_952 = (x_832 & x_951);
	assign x_953 = (x_714 & x_952);
	assign o_1 = x_95);
endmodule
