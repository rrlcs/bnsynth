// Benchmark "SKOLEMFORMULA" written by ABC on Wed May 18 01:29:28 2022

module SKOLEMFORMULA ( 
    i0,
    i1, i2, i3  );
  input  i0;
  output i1, i2, i3;
  assign i1 = 1'b1;
  assign i3 = 1'b1;
  assign i2 = ~i0;
endmodule


