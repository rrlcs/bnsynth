module formula(i_1,i_2,i_3,i_4,i_5,i_6,i_7,i_8,i_9,i_10,i_11,i_12,i_13,i_14,i_15,i_16,i_17,i_18,i_19,i_20,i_21,i_22,i_23,i_24,i_25,i_26,i_27,i_28,i_29,i_30,i_31,i_32,i_33,i_34,i_35,i_36,i_37,i_38,i_39,i_40,i_41,i_42,i_43,i_44,i_45,i_46,i_47,i_48,i_49,i_50,i_51,i_52,i_53,i_54,i_55,i_56,i_57,i_58,i_59,i_60,i_61,i_62,i_63,i_64,i_65,i_66,i_67,i_68,x_69,x_70,x_71,x_72,x_73,x_74,x_75,x_76,x_77,x_78,x_79,x_80,x_81,x_82,x_83,x_84,x_85,x_86,x_87,x_88,x_89,x_90,x_91,x_92,x_93,x_94,x_95,x_96,x_97,x_98,x_99,x_100,x_101,x_102,x_103,x_104,x_105,x_106,x_107,x_108,x_109,x_110,x_111,x_112,x_113,x_114,x_115,x_116,x_117,x_118,x_119,x_120,x_121,x_122,x_123,x_124,x_125,x_126,x_127,x_128,x_129,x_130,x_131,x_132,x_133,x_134,x_135,x_136,x_137,x_138,x_139,x_140,x_141,x_142,x_143,x_144,x_145,x_146,x_147,x_148,x_149,x_150,x_151,x_152,x_153,x_154,x_155,x_156,x_157,x_158,x_159,x_160,x_161,x_162,x_163,x_164,x_165,x_166,x_167,x_168,x_169,x_170,x_171,x_172,x_173,x_174,x_175,x_176,x_177,x_178,x_179,x_180,x_181,x_182,x_183,x_184,x_185,x_186,x_187,x_188,x_189,x_190,x_191,x_192,x_193,x_194,x_195,x_196,x_197,x_198,x_199,x_200,x_201,x_202,x_203,x_204,x_205,x_206,x_207,x_208,x_209,x_210,x_211,x_212,x_213,x_214,x_215,x_216,x_217,x_218,x_219,x_220,x_221,x_222,x_223,x_224,x_225,x_226,x_227,x_228,x_229,x_230,x_231,x_232,x_233,x_234,x_235,x_236,x_237,x_238,x_239,x_240,x_241,x_242,x_243,x_244,x_245,x_246,x_247,x_248,x_249,x_250,x_251,x_252,x_253,x_254,x_255,x_256,x_257,x_258,x_259,x_260,x_261,x_262,x_263,x_264,x_265,x_266,x_267,x_268,x_269,x_270,x_271,x_272,x_273,x_274,x_275,x_276,x_277,x_278,x_279,x_280,x_281,x_282,x_283,x_284,x_285,x_286,x_287,x_288,x_289,x_290,x_291,x_292,x_293,x_294,x_295,x_296,x_297,x_298,x_299,x_300,x_301,x_302,x_303,x_304,x_305,x_306,x_307,x_308,x_309,x_310,x_311,x_312,x_313,x_314,x_315,x_316,x_317,x_318,x_319,x_320,x_321,x_322,x_323,x_324,x_325,x_326,x_327,x_328,x_329,x_330,x_331,x_332,x_333,x_334,x_335,x_336,x_337,x_338,x_339,x_340,x_341,x_342,x_343,x_344,x_345,x_346,x_347,x_348,x_349,x_350,x_351,x_352,x_353,x_354,x_355,x_356,x_357,x_358,x_359,x_360,x_361,x_362,x_363,x_364,x_365,x_366,x_367,x_368,x_369,x_370,x_371,x_372,x_373,x_374,x_375,x_376,x_377,x_378,x_379,x_380,x_381,x_382,x_383,x_384,x_385,x_386,x_387,x_388,x_389,x_390,x_391,x_392,x_393,x_394,x_395,x_396,x_397,x_398,x_399,x_400,x_401,x_402,x_403,x_404,x_405,x_406,x_407,x_408,x_409,x_410,x_411,x_412,x_413,x_414,x_415,x_416,x_417,x_418,x_419,x_420,x_421,x_422,x_423,x_424,x_425,x_426,x_427,x_428,x_429,x_430,x_431,x_432,x_433,x_434,x_435,x_436,x_437,x_438,x_439,x_440,x_441,x_442,x_443,x_444,x_445,x_446,x_447,x_448,x_449,x_450,x_451,x_452,x_453,x_454,x_455,x_456,x_457,x_458,x_459,x_460,x_461,x_462,x_463,x_464,x_465,x_466,x_467,x_468,x_469,x_470,x_471,x_472,x_473,x_474,x_475,x_476,x_477,x_478,x_479,x_480,x_481,x_482,x_483,x_484,x_485,x_486,x_487,x_488,x_489,x_490,x_491,x_492,x_493,x_494,x_495,x_496,x_497,x_498,x_499,x_500,x_501,x_502,x_503,x_504,x_505,x_506,x_507,x_508,x_509,x_510,x_511,x_512,x_513,x_514,x_515,x_516,x_517,x_518,x_519,x_520,x_521,x_522,x_523,x_524,x_525,x_526,x_527,x_528,x_529,x_530,x_531,x_532,x_533,x_534,x_535,x_536,x_537,x_538,x_539,x_540,x_541,x_542,x_543,x_544,x_545,x_546,x_547,x_548,x_549,x_550,x_551,x_552,x_553,x_554,x_555,x_556,x_557,x_558,x_559,x_560,x_561,x_562,x_563,x_564,x_565,x_566,x_567,x_568,x_569,x_570,x_571,x_572,x_573,x_574,x_575,x_576,x_577,x_578,x_579,x_580,x_581,x_582,x_583,x_584,x_585,x_586,x_587,x_588,x_589,x_590,x_591,x_592,x_593,x_594,x_595,x_596,x_597,x_598,x_599,x_600,x_601,x_602,x_603,x_604,x_605,x_606,x_607,x_608,x_609,x_610,x_611,x_612,x_613,x_614,x_615,x_616,x_617,x_618,x_619,x_620,x_621,x_622,x_623,x_624,x_625,x_626,x_627,x_628,x_629,x_630,x_631,x_632,x_633,x_634,x_635,x_636,x_637,x_638,x_639,x_640,x_641,x_642,x_643,x_644,x_645,x_646,x_647,x_648,x_649,x_650,x_651,x_652,x_653,x_654,x_655,x_656,x_657,x_658,x_659,x_660,x_661,x_662,x_663,x_664,x_665,x_666,x_667,x_668,x_669,x_670,x_671,x_672,x_673,x_674,x_675,x_676,x_677,x_678,x_679,x_680,x_681,x_682,x_683,x_684,x_685,x_686,x_687,x_688,x_689,x_690,x_691,x_692,x_693,x_694,x_695,x_696,x_697,x_698,x_699,x_700,x_701,x_702,x_703,x_704,x_705,x_706,x_707,x_708,x_709,x_710,x_711,x_712,x_713,x_714,x_715,x_716,x_717,x_718,x_719,x_720,x_721,x_722,x_723,x_724,x_725,x_726,x_727,x_728,x_729,x_730,x_731,x_732,x_733,x_734,x_735,x_736,x_737,x_738,x_739,x_740,x_741,x_742,x_743,x_744,x_745,x_746,x_747,x_748,x_749,x_750,x_751,x_752,x_753,x_754,x_755,x_756,x_757,x_758,x_759,x_760,x_761,x_762,x_763,x_764,x_765,x_766,x_767,x_768,x_769,x_770,x_771,x_772,x_773,x_774,x_775,x_776,x_777,x_778,x_779,x_780,x_781,x_782,x_783,x_784,x_785,x_786,x_787,x_788,x_789,x_790,x_791,x_792,x_793,x_794,x_795,x_796,x_797,x_798,x_799,x_800,x_801,x_802,x_803,x_804,x_805,x_806,x_807,x_808,x_809,x_810,x_811,x_812,x_813,x_814,x_815,x_816,x_817,x_818,x_819,x_820,x_821,x_822,x_823,x_824,x_825,x_826,x_827,x_828,x_829,x_830,x_831,x_832,x_833,x_834,x_835,x_836,x_837,x_838,x_839,x_840,x_841,x_842,x_843,x_844,x_845,x_846,x_847,x_848,x_849,x_850,x_851,x_852,x_853,x_854,x_855,x_856,x_857,x_858,x_859,x_860,x_861,x_862,x_863,x_864,x_865,x_866,x_867,x_868,x_869,x_870,x_871,x_872,x_873,x_874,x_875,x_876,x_877,x_878,x_879,x_880,x_881,x_882,x_883,x_884,x_885,x_886,x_887,x_888,x_889,x_890,x_891,x_892,x_893,x_894,x_895,x_896,x_897,x_898,x_899,x_900,x_901,x_902,x_903,x_904,x_905,x_906,x_907,x_908,x_909,x_910,x_911,x_912,x_913,x_914,x_915,x_916,x_917,x_918,x_919,x_920,x_921,x_922,x_923,x_924,x_925,x_926,x_927,x_928,x_929,x_930,x_931,x_932,x_933,x_934,x_935,x_936,x_937,x_938,x_939,x_940,x_941,x_942,x_943,x_944,x_945,x_946,x_947,x_948,x_949,x_950,x_951,x_952,x_953,x_954,x_955,x_956,x_957,x_958,x_959,x_960,x_961,x_962,x_963,x_964,x_965,x_966,x_967,x_968,x_969,x_970,x_971,x_972,x_973,x_974,x_975,x_976,x_977,x_978,x_979,x_980,x_981,x_982,x_983,x_984,x_985,x_986,x_987,x_988,x_989,x_990,x_991,x_992,x_993,x_994,x_995,x_996,x_997,x_998,x_999,x_1000,x_1001,x_1002,x_1003,x_1004,x_1005,x_1006,x_1007,x_1008,x_1009,x_1010,x_1011,x_1012,x_1013,x_1014,x_1015,x_1016,x_1017,x_1018,x_1019,x_1020,x_1021,x_1022,x_1023,x_1024,x_1025,x_1026,x_1027,x_1028,x_1029,x_1030,x_1031,x_1032,x_1033,x_1034,x_1035,x_1036,x_1037,x_1038,x_1039,x_1040,x_1041,x_1042,x_1043,x_1044,x_1045,x_1046,x_1047,x_1048,x_1049,x_1050,x_1051,x_1052,x_1053,x_1054,x_1055,x_1056,x_1057,x_1058,x_1059,x_1060,x_1061,x_1062,x_1063,x_1064,x_1065,x_1066,x_1067,x_1068,x_1069,x_1070,x_1071,x_1072,x_1073,x_1074,x_1075,x_1076,x_1077,x_1078,x_1079,x_1080,x_1081,x_1082,x_1083,x_1084,x_1085,x_1086,x_1087,x_1088,x_1089,x_1090,x_1091,x_1092,x_1093,x_1094,x_1095,x_1096,x_1097,x_1098,x_1099,x_1100,x_1101,x_1102,x_1103,x_1104,x_1105,x_1106,x_1107,x_1108,x_1109,x_1110,x_1111,x_1112,x_1113,x_1114,x_1115,x_1116,x_1117,x_1118,x_1119,x_1120,x_1121,x_1122,x_1123,x_1124,x_1125,x_1126,x_1127,x_1128,x_1129,x_1130,x_1131,x_1132,x_1133,x_1134,x_1135,x_1136,x_1137,x_1138,x_1139,x_1140,x_1141,x_1142,x_1143,x_1144,x_1145,x_1146,x_1147,x_1148,x_1149,x_1150,x_1151,x_1152,x_1153,x_1154,x_1155,x_1156,x_1157,x_1158,x_1159,x_1160,x_1161,x_1162,x_1163,x_1164,x_1165,x_1166,x_1167,x_1168,x_1169,x_1170,x_1171,x_1172,x_1173,x_1174,x_1175,x_1176,x_1177,x_1178,x_1179,x_1180,x_1181,x_1182,x_1183,x_1184,x_1185,x_1186,x_1187,x_1188,x_1189,x_1190,x_1191,x_1192,x_1193,x_1194,x_1195,x_1196,x_1197,x_1198,x_1199,x_1200,x_1201,x_1202,x_1203,x_1204,x_1205,x_1206,x_1207,x_1208,x_1209,x_1210,x_1211,x_1212,x_1213,x_1214,x_1215,x_1216,x_1217,x_1218,x_1219,x_1220,x_1221,x_1222,x_1223,x_1224,x_1225,x_1226,x_1227,x_1228,x_1229,x_1230,x_1231,x_1232,x_1233,x_1234,x_1235,x_1236,x_1237,x_1238,x_1239,x_1240,x_1241,x_1242,x_1243,x_1244,x_1245,x_1246,x_1247,x_1248,x_1249,x_1250,x_1251,x_1252,x_1253,x_1254,x_1255,x_1256,x_1257,x_1258,x_1259,x_1260,x_1261,x_1262,x_1263,x_1264,x_1265,x_1266,x_1267,x_1268,x_1269,x_1270,x_1271,x_1272,x_1273,x_1274,x_1275,x_1276,x_1277,x_1278,x_1279,x_1280,x_1281,x_1282,x_1283,x_1284,x_1285,x_1286,x_1287,x_1288,x_1289,x_1290,x_1291,x_1292,x_1293,x_1294,x_1295,x_1296,x_1297,x_1298,x_1299,x_1300,x_1301,x_1302,x_1303,x_1304,x_1305,x_1306,x_1307,x_1308,x_1309,x_1310,x_1311,x_1312,x_1313,x_1314,x_1315,x_1316,x_1317,x_1318,x_1319,x_1320,x_1321,x_1322,x_1323,x_1324,x_1325,x_1326,x_1327,x_1328,x_1329,x_1330,x_1331,x_1332,x_1333,x_1334,x_1335,x_1336,x_1337,x_1338,x_1339,x_1340,x_1341,x_1342,x_1343,x_1344,x_1345,x_1346,x_1347,x_1348,x_1349,x_1350,x_1351,x_1352,x_1353,x_1354,x_1355,x_1356,x_1357,x_1358,x_1359,x_1360,x_1361,x_1362,x_1363,x_1364,x_1365,x_1366,x_1367,x_1368,x_1369,x_1370,x_1371,x_1372,x_1373,x_1374,x_1375,x_1376,x_1377,x_1378,x_1379,x_1380,x_1381,x_1382,x_1383,x_1384,x_1385,x_1386,x_1387,x_1388,x_1389,x_1390,x_1391,x_1392,x_1393,x_1394,x_1395,x_1396,x_1397,x_1398,x_1399,x_1400,x_1401,x_1402,x_1403,x_1404,x_1405,x_1406,x_1407,x_1408,x_1409,x_1410,x_1411,x_1412,x_1413,x_1414,x_1415,x_1416,x_1417,x_1418,x_1419,x_1420,x_1421,x_1422,x_1423,x_1424,x_1425,x_1426,x_1427,x_1428,x_1429,x_1430,x_1431,x_1432,x_1433,x_1434,x_1435,x_1436,x_1437,x_1438,x_1439,x_1440,x_1441,x_1442,x_1443,x_1444,x_1445,x_1446,x_1447,x_1448,x_1449,x_1450,x_1451,x_1452,x_1453,x_1454,x_1455,x_1456,x_1457,x_1458,x_1459,x_1460,x_1461,x_1462,x_1463,x_1464,x_1465,x_1466,x_1467,x_1468,x_1469,x_1470,x_1471,x_1472,x_1473,x_1474,x_1475,x_1476,x_1477,x_1478,x_1479,x_1480,x_1481,x_1482,x_1483,x_1484,x_1485,x_1486,x_1487,x_1488,x_1489,x_1490,x_1491,x_1492,x_1493,x_1494,x_1495,x_1496,x_1497,x_1498,x_1499,x_1500,x_1501,x_1502,x_1503,x_1504,x_1505,x_1506,x_1507,x_1508,x_1509,x_1510,x_1511,x_1512,x_1513,x_1514,x_1515,x_1516,x_1517,x_1518,x_1519,x_1520,x_1521,x_1522,x_1523,x_1524,x_1525,x_1526,x_1527,x_1528,x_1529,x_1530,x_1531,x_1532,x_1533,x_1534,x_1535,x_1536,x_1537,x_1538,x_1539,x_1540,x_1541,x_1542,x_1543,x_1544,x_1545,x_1546,x_1547,x_1548,x_1549,x_1550,x_1551,x_1552,x_1553,x_1554,x_1555,x_1556,x_1557,x_1558,x_1559,x_1560,x_1561,x_1562,x_1563,x_1564,x_1565,x_1566,x_1567,x_1568,x_1569,x_1570,x_1571,x_1572,x_1573,x_1574,x_1575,x_1576,x_1577,x_1578,o_1);
	input i_1;
	input i_2;
	input i_3;
	input i_4;
	input i_5;
	input i_6;
	input i_7;
	input i_8;
	input i_9;
	input i_10;
	input i_11;
	input i_12;
	input i_13;
	input i_14;
	input i_15;
	input i_16;
	input i_17;
	input i_18;
	input i_19;
	input i_20;
	input i_21;
	input i_22;
	input i_23;
	input i_24;
	input i_25;
	input i_26;
	input i_27;
	input i_28;
	input i_29;
	input i_30;
	input i_31;
	input i_32;
	input i_33;
	input i_34;
	input i_35;
	input i_36;
	input i_37;
	input i_38;
	input i_39;
	input i_40;
	input i_41;
	input i_42;
	input i_43;
	input i_44;
	input i_45;
	input i_46;
	input i_47;
	input i_48;
	input i_49;
	input i_50;
	input i_51;
	input i_52;
	input i_53;
	input i_54;
	input i_55;
	input i_56;
	input i_57;
	input i_58;
	input i_59;
	input i_60;
	input i_61;
	input i_62;
	input i_63;
	input i_64;
	input i_65;
	input i_66;
	input i_67;
	input i_68;
	input x_69;
	input x_70;
	input x_71;
	input x_72;
	input x_73;
	input x_74;
	input x_75;
	input x_76;
	input x_77;
	input x_78;
	input x_79;
	input x_80;
	input x_81;
	input x_82;
	input x_83;
	input x_84;
	input x_85;
	input x_86;
	input x_87;
	input x_88;
	input x_89;
	input x_90;
	input x_91;
	input x_92;
	input x_93;
	input x_94;
	input x_95;
	input x_96;
	input x_97;
	input x_98;
	input x_99;
	input x_100;
	input x_101;
	input x_102;
	input x_103;
	input x_104;
	input x_105;
	input x_106;
	input x_107;
	input x_108;
	input x_109;
	input x_110;
	input x_111;
	input x_112;
	input x_113;
	input x_114;
	input x_115;
	input x_116;
	input x_117;
	input x_118;
	input x_119;
	input x_120;
	input x_121;
	input x_122;
	input x_123;
	input x_124;
	input x_125;
	input x_126;
	input x_127;
	input x_128;
	input x_129;
	input x_130;
	input x_131;
	input x_132;
	input x_133;
	input x_134;
	input x_135;
	input x_136;
	input x_137;
	input x_138;
	input x_139;
	input x_140;
	input x_141;
	input x_142;
	input x_143;
	input x_144;
	input x_145;
	input x_146;
	input x_147;
	input x_148;
	input x_149;
	input x_150;
	input x_151;
	input x_152;
	input x_153;
	input x_154;
	input x_155;
	input x_156;
	input x_157;
	input x_158;
	input x_159;
	input x_160;
	input x_161;
	input x_162;
	input x_163;
	input x_164;
	input x_165;
	input x_166;
	input x_167;
	input x_168;
	input x_169;
	input x_170;
	input x_171;
	input x_172;
	input x_173;
	input x_174;
	input x_175;
	input x_176;
	input x_177;
	input x_178;
	input x_179;
	input x_180;
	input x_181;
	input x_182;
	input x_183;
	input x_184;
	input x_185;
	input x_186;
	input x_187;
	input x_188;
	input x_189;
	input x_190;
	input x_191;
	input x_192;
	input x_193;
	input x_194;
	input x_195;
	input x_196;
	input x_197;
	input x_198;
	input x_199;
	input x_200;
	input x_201;
	input x_202;
	input x_203;
	input x_204;
	input x_205;
	input x_206;
	input x_207;
	input x_208;
	input x_209;
	input x_210;
	input x_211;
	input x_212;
	input x_213;
	input x_214;
	input x_215;
	input x_216;
	input x_217;
	input x_218;
	input x_219;
	input x_220;
	input x_221;
	input x_222;
	input x_223;
	input x_224;
	input x_225;
	input x_226;
	input x_227;
	input x_228;
	input x_229;
	input x_230;
	input x_231;
	input x_232;
	input x_233;
	input x_234;
	input x_235;
	input x_236;
	input x_237;
	input x_238;
	input x_239;
	input x_240;
	input x_241;
	input x_242;
	input x_243;
	input x_244;
	input x_245;
	input x_246;
	input x_247;
	input x_248;
	input x_249;
	input x_250;
	input x_251;
	input x_252;
	input x_253;
	input x_254;
	input x_255;
	input x_256;
	input x_257;
	input x_258;
	input x_259;
	input x_260;
	input x_261;
	input x_262;
	input x_263;
	input x_264;
	input x_265;
	input x_266;
	input x_267;
	input x_268;
	input x_269;
	input x_270;
	input x_271;
	input x_272;
	input x_273;
	input x_274;
	input x_275;
	input x_276;
	input x_277;
	input x_278;
	input x_279;
	input x_280;
	input x_281;
	input x_282;
	input x_283;
	input x_284;
	input x_285;
	input x_286;
	input x_287;
	input x_288;
	input x_289;
	input x_290;
	input x_291;
	input x_292;
	input x_293;
	input x_294;
	input x_295;
	input x_296;
	input x_297;
	input x_298;
	input x_299;
	input x_300;
	input x_301;
	input x_302;
	input x_303;
	input x_304;
	input x_305;
	input x_306;
	input x_307;
	input x_308;
	input x_309;
	input x_310;
	input x_311;
	input x_312;
	input x_313;
	input x_314;
	input x_315;
	input x_316;
	input x_317;
	input x_318;
	input x_319;
	input x_320;
	input x_321;
	input x_322;
	input x_323;
	input x_324;
	input x_325;
	input x_326;
	input x_327;
	input x_328;
	input x_329;
	input x_330;
	input x_331;
	input x_332;
	input x_333;
	input x_334;
	input x_335;
	input x_336;
	input x_337;
	input x_338;
	input x_339;
	input x_340;
	input x_341;
	input x_342;
	input x_343;
	input x_344;
	input x_345;
	input x_346;
	input x_347;
	input x_348;
	input x_349;
	input x_350;
	input x_351;
	input x_352;
	input x_353;
	input x_354;
	input x_355;
	input x_356;
	input x_357;
	input x_358;
	input x_359;
	input x_360;
	input x_361;
	input x_362;
	input x_363;
	input x_364;
	input x_365;
	input x_366;
	input x_367;
	input x_368;
	input x_369;
	input x_370;
	input x_371;
	input x_372;
	input x_373;
	input x_374;
	input x_375;
	input x_376;
	input x_377;
	input x_378;
	input x_379;
	input x_380;
	input x_381;
	input x_382;
	input x_383;
	input x_384;
	input x_385;
	input x_386;
	input x_387;
	input x_388;
	input x_389;
	input x_390;
	input x_391;
	input x_392;
	input x_393;
	input x_394;
	input x_395;
	input x_396;
	input x_397;
	input x_398;
	input x_399;
	input x_400;
	input x_401;
	input x_402;
	input x_403;
	input x_404;
	input x_405;
	input x_406;
	input x_407;
	input x_408;
	input x_409;
	input x_410;
	input x_411;
	input x_412;
	input x_413;
	input x_414;
	input x_415;
	input x_416;
	input x_417;
	input x_418;
	input x_419;
	input x_420;
	input x_421;
	input x_422;
	input x_423;
	input x_424;
	input x_425;
	input x_426;
	input x_427;
	input x_428;
	input x_429;
	input x_430;
	input x_431;
	input x_432;
	input x_433;
	input x_434;
	input x_435;
	input x_436;
	input x_437;
	input x_438;
	input x_439;
	input x_440;
	input x_441;
	input x_442;
	input x_443;
	input x_444;
	input x_445;
	input x_446;
	input x_447;
	input x_448;
	input x_449;
	input x_450;
	input x_451;
	input x_452;
	input x_453;
	input x_454;
	input x_455;
	input x_456;
	input x_457;
	input x_458;
	input x_459;
	input x_460;
	input x_461;
	input x_462;
	input x_463;
	input x_464;
	input x_465;
	input x_466;
	input x_467;
	input x_468;
	input x_469;
	input x_470;
	input x_471;
	input x_472;
	input x_473;
	input x_474;
	input x_475;
	input x_476;
	input x_477;
	input x_478;
	input x_479;
	input x_480;
	input x_481;
	input x_482;
	input x_483;
	input x_484;
	input x_485;
	input x_486;
	input x_487;
	input x_488;
	input x_489;
	input x_490;
	input x_491;
	input x_492;
	input x_493;
	input x_494;
	input x_495;
	input x_496;
	input x_497;
	input x_498;
	input x_499;
	input x_500;
	input x_501;
	input x_502;
	input x_503;
	input x_504;
	input x_505;
	input x_506;
	input x_507;
	input x_508;
	input x_509;
	input x_510;
	input x_511;
	input x_512;
	input x_513;
	input x_514;
	input x_515;
	input x_516;
	input x_517;
	input x_518;
	input x_519;
	input x_520;
	input x_521;
	input x_522;
	input x_523;
	input x_524;
	input x_525;
	input x_526;
	input x_527;
	input x_528;
	input x_529;
	input x_530;
	input x_531;
	input x_532;
	input x_533;
	input x_534;
	input x_535;
	input x_536;
	input x_537;
	input x_538;
	input x_539;
	input x_540;
	input x_541;
	input x_542;
	input x_543;
	input x_544;
	input x_545;
	input x_546;
	input x_547;
	input x_548;
	input x_549;
	input x_550;
	input x_551;
	input x_552;
	input x_553;
	input x_554;
	input x_555;
	input x_556;
	input x_557;
	input x_558;
	input x_559;
	input x_560;
	input x_561;
	input x_562;
	input x_563;
	input x_564;
	input x_565;
	input x_566;
	input x_567;
	input x_568;
	input x_569;
	input x_570;
	input x_571;
	input x_572;
	input x_573;
	input x_574;
	input x_575;
	input x_576;
	input x_577;
	input x_578;
	input x_579;
	input x_580;
	input x_581;
	input x_582;
	input x_583;
	input x_584;
	input x_585;
	input x_586;
	input x_587;
	input x_588;
	input x_589;
	input x_590;
	input x_591;
	input x_592;
	input x_593;
	input x_594;
	input x_595;
	input x_596;
	input x_597;
	input x_598;
	input x_599;
	input x_600;
	input x_601;
	input x_602;
	input x_603;
	input x_604;
	input x_605;
	input x_606;
	input x_607;
	input x_608;
	input x_609;
	input x_610;
	input x_611;
	input x_612;
	input x_613;
	input x_614;
	input x_615;
	input x_616;
	input x_617;
	input x_618;
	input x_619;
	input x_620;
	input x_621;
	input x_622;
	input x_623;
	input x_624;
	input x_625;
	input x_626;
	input x_627;
	input x_628;
	input x_629;
	input x_630;
	input x_631;
	input x_632;
	input x_633;
	input x_634;
	input x_635;
	input x_636;
	input x_637;
	input x_638;
	input x_639;
	input x_640;
	input x_641;
	input x_642;
	input x_643;
	input x_644;
	input x_645;
	input x_646;
	input x_647;
	input x_648;
	input x_649;
	input x_650;
	input x_651;
	input x_652;
	input x_653;
	input x_654;
	input x_655;
	input x_656;
	input x_657;
	input x_658;
	input x_659;
	input x_660;
	input x_661;
	input x_662;
	input x_663;
	input x_664;
	input x_665;
	input x_666;
	input x_667;
	input x_668;
	input x_669;
	input x_670;
	input x_671;
	input x_672;
	input x_673;
	input x_674;
	input x_675;
	input x_676;
	input x_677;
	input x_678;
	input x_679;
	input x_680;
	input x_681;
	input x_682;
	input x_683;
	input x_684;
	input x_685;
	input x_686;
	input x_687;
	input x_688;
	input x_689;
	input x_690;
	input x_691;
	input x_692;
	input x_693;
	input x_694;
	input x_695;
	input x_696;
	input x_697;
	input x_698;
	input x_699;
	input x_700;
	input x_701;
	input x_702;
	input x_703;
	input x_704;
	input x_705;
	input x_706;
	input x_707;
	input x_708;
	input x_709;
	input x_710;
	input x_711;
	input x_712;
	input x_713;
	input x_714;
	input x_715;
	input x_716;
	input x_717;
	input x_718;
	input x_719;
	input x_720;
	input x_721;
	input x_722;
	input x_723;
	input x_724;
	input x_725;
	input x_726;
	input x_727;
	input x_728;
	input x_729;
	input x_730;
	input x_731;
	input x_732;
	input x_733;
	input x_734;
	input x_735;
	input x_736;
	input x_737;
	input x_738;
	input x_739;
	input x_740;
	input x_741;
	input x_742;
	input x_743;
	input x_744;
	input x_745;
	input x_746;
	input x_747;
	input x_748;
	input x_749;
	input x_750;
	input x_751;
	input x_752;
	input x_753;
	input x_754;
	input x_755;
	input x_756;
	input x_757;
	input x_758;
	input x_759;
	input x_760;
	input x_761;
	input x_762;
	input x_763;
	input x_764;
	input x_765;
	input x_766;
	input x_767;
	input x_768;
	input x_769;
	input x_770;
	input x_771;
	input x_772;
	input x_773;
	input x_774;
	input x_775;
	input x_776;
	input x_777;
	input x_778;
	input x_779;
	input x_780;
	input x_781;
	input x_782;
	input x_783;
	input x_784;
	input x_785;
	input x_786;
	input x_787;
	input x_788;
	input x_789;
	input x_790;
	input x_791;
	input x_792;
	input x_793;
	input x_794;
	input x_795;
	input x_796;
	input x_797;
	input x_798;
	input x_799;
	input x_800;
	input x_801;
	input x_802;
	input x_803;
	input x_804;
	input x_805;
	input x_806;
	input x_807;
	input x_808;
	input x_809;
	input x_810;
	input x_811;
	input x_812;
	input x_813;
	input x_814;
	input x_815;
	input x_816;
	input x_817;
	input x_818;
	input x_819;
	input x_820;
	input x_821;
	input x_822;
	input x_823;
	input x_824;
	input x_825;
	input x_826;
	input x_827;
	input x_828;
	input x_829;
	input x_830;
	input x_831;
	input x_832;
	input x_833;
	input x_834;
	input x_835;
	input x_836;
	input x_837;
	input x_838;
	input x_839;
	input x_840;
	input x_841;
	input x_842;
	input x_843;
	input x_844;
	input x_845;
	input x_846;
	input x_847;
	input x_848;
	input x_849;
	input x_850;
	input x_851;
	input x_852;
	input x_853;
	input x_854;
	input x_855;
	input x_856;
	input x_857;
	input x_858;
	input x_859;
	input x_860;
	input x_861;
	input x_862;
	input x_863;
	input x_864;
	input x_865;
	input x_866;
	input x_867;
	input x_868;
	input x_869;
	input x_870;
	input x_871;
	input x_872;
	input x_873;
	input x_874;
	input x_875;
	input x_876;
	input x_877;
	input x_878;
	input x_879;
	input x_880;
	input x_881;
	input x_882;
	input x_883;
	input x_884;
	input x_885;
	input x_886;
	input x_887;
	input x_888;
	input x_889;
	input x_890;
	input x_891;
	input x_892;
	input x_893;
	input x_894;
	input x_895;
	input x_896;
	input x_897;
	input x_898;
	input x_899;
	input x_900;
	input x_901;
	input x_902;
	input x_903;
	input x_904;
	input x_905;
	input x_906;
	input x_907;
	input x_908;
	input x_909;
	input x_910;
	input x_911;
	input x_912;
	input x_913;
	input x_914;
	input x_915;
	input x_916;
	input x_917;
	input x_918;
	input x_919;
	input x_920;
	input x_921;
	input x_922;
	input x_923;
	input x_924;
	input x_925;
	input x_926;
	input x_927;
	input x_928;
	input x_929;
	input x_930;
	input x_931;
	input x_932;
	input x_933;
	input x_934;
	input x_935;
	input x_936;
	input x_937;
	input x_938;
	input x_939;
	input x_940;
	input x_941;
	input x_942;
	input x_943;
	input x_944;
	input x_945;
	input x_946;
	input x_947;
	input x_948;
	input x_949;
	input x_950;
	input x_951;
	input x_952;
	input x_953;
	input x_954;
	input x_955;
	input x_956;
	input x_957;
	input x_958;
	input x_959;
	input x_960;
	input x_961;
	input x_962;
	input x_963;
	input x_964;
	input x_965;
	input x_966;
	input x_967;
	input x_968;
	input x_969;
	input x_970;
	input x_971;
	input x_972;
	input x_973;
	input x_974;
	input x_975;
	input x_976;
	input x_977;
	input x_978;
	input x_979;
	input x_980;
	input x_981;
	input x_982;
	input x_983;
	input x_984;
	input x_985;
	input x_986;
	input x_987;
	input x_988;
	input x_989;
	input x_990;
	input x_991;
	input x_992;
	input x_993;
	input x_994;
	input x_995;
	input x_996;
	input x_997;
	input x_998;
	input x_999;
	input x_1000;
	input x_1001;
	input x_1002;
	input x_1003;
	input x_1004;
	input x_1005;
	input x_1006;
	input x_1007;
	input x_1008;
	input x_1009;
	input x_1010;
	input x_1011;
	input x_1012;
	input x_1013;
	input x_1014;
	input x_1015;
	input x_1016;
	input x_1017;
	input x_1018;
	input x_1019;
	input x_1020;
	input x_1021;
	input x_1022;
	input x_1023;
	input x_1024;
	input x_1025;
	input x_1026;
	input x_1027;
	input x_1028;
	input x_1029;
	input x_1030;
	input x_1031;
	input x_1032;
	input x_1033;
	input x_1034;
	input x_1035;
	input x_1036;
	input x_1037;
	input x_1038;
	input x_1039;
	input x_1040;
	input x_1041;
	input x_1042;
	input x_1043;
	input x_1044;
	input x_1045;
	input x_1046;
	input x_1047;
	input x_1048;
	input x_1049;
	input x_1050;
	input x_1051;
	input x_1052;
	input x_1053;
	input x_1054;
	input x_1055;
	input x_1056;
	input x_1057;
	input x_1058;
	input x_1059;
	input x_1060;
	input x_1061;
	input x_1062;
	input x_1063;
	input x_1064;
	input x_1065;
	input x_1066;
	input x_1067;
	input x_1068;
	input x_1069;
	input x_1070;
	input x_1071;
	input x_1072;
	input x_1073;
	input x_1074;
	input x_1075;
	input x_1076;
	input x_1077;
	input x_1078;
	input x_1079;
	input x_1080;
	input x_1081;
	input x_1082;
	input x_1083;
	input x_1084;
	input x_1085;
	input x_1086;
	input x_1087;
	input x_1088;
	input x_1089;
	input x_1090;
	input x_1091;
	input x_1092;
	input x_1093;
	input x_1094;
	input x_1095;
	input x_1096;
	input x_1097;
	input x_1098;
	input x_1099;
	input x_1100;
	input x_1101;
	input x_1102;
	input x_1103;
	input x_1104;
	input x_1105;
	input x_1106;
	input x_1107;
	input x_1108;
	input x_1109;
	input x_1110;
	input x_1111;
	input x_1112;
	input x_1113;
	input x_1114;
	input x_1115;
	input x_1116;
	input x_1117;
	input x_1118;
	input x_1119;
	input x_1120;
	input x_1121;
	input x_1122;
	input x_1123;
	input x_1124;
	input x_1125;
	input x_1126;
	input x_1127;
	input x_1128;
	input x_1129;
	input x_1130;
	input x_1131;
	input x_1132;
	input x_1133;
	input x_1134;
	input x_1135;
	input x_1136;
	input x_1137;
	input x_1138;
	input x_1139;
	input x_1140;
	input x_1141;
	input x_1142;
	input x_1143;
	input x_1144;
	input x_1145;
	input x_1146;
	input x_1147;
	input x_1148;
	input x_1149;
	input x_1150;
	input x_1151;
	input x_1152;
	input x_1153;
	input x_1154;
	input x_1155;
	input x_1156;
	input x_1157;
	input x_1158;
	input x_1159;
	input x_1160;
	input x_1161;
	input x_1162;
	input x_1163;
	input x_1164;
	input x_1165;
	input x_1166;
	input x_1167;
	input x_1168;
	input x_1169;
	input x_1170;
	input x_1171;
	input x_1172;
	input x_1173;
	input x_1174;
	input x_1175;
	input x_1176;
	input x_1177;
	input x_1178;
	input x_1179;
	input x_1180;
	input x_1181;
	input x_1182;
	input x_1183;
	input x_1184;
	input x_1185;
	input x_1186;
	input x_1187;
	input x_1188;
	input x_1189;
	input x_1190;
	input x_1191;
	input x_1192;
	input x_1193;
	input x_1194;
	input x_1195;
	input x_1196;
	input x_1197;
	input x_1198;
	input x_1199;
	input x_1200;
	input x_1201;
	input x_1202;
	input x_1203;
	input x_1204;
	input x_1205;
	input x_1206;
	input x_1207;
	input x_1208;
	input x_1209;
	input x_1210;
	input x_1211;
	input x_1212;
	input x_1213;
	input x_1214;
	input x_1215;
	input x_1216;
	input x_1217;
	input x_1218;
	input x_1219;
	input x_1220;
	input x_1221;
	input x_1222;
	input x_1223;
	input x_1224;
	input x_1225;
	input x_1226;
	input x_1227;
	input x_1228;
	input x_1229;
	input x_1230;
	input x_1231;
	input x_1232;
	input x_1233;
	input x_1234;
	input x_1235;
	input x_1236;
	input x_1237;
	input x_1238;
	input x_1239;
	input x_1240;
	input x_1241;
	input x_1242;
	input x_1243;
	input x_1244;
	input x_1245;
	input x_1246;
	input x_1247;
	input x_1248;
	input x_1249;
	input x_1250;
	input x_1251;
	input x_1252;
	input x_1253;
	input x_1254;
	input x_1255;
	input x_1256;
	input x_1257;
	input x_1258;
	input x_1259;
	input x_1260;
	input x_1261;
	input x_1262;
	input x_1263;
	input x_1264;
	input x_1265;
	input x_1266;
	input x_1267;
	input x_1268;
	input x_1269;
	input x_1270;
	input x_1271;
	input x_1272;
	input x_1273;
	input x_1274;
	input x_1275;
	input x_1276;
	input x_1277;
	input x_1278;
	input x_1279;
	input x_1280;
	input x_1281;
	input x_1282;
	input x_1283;
	input x_1284;
	input x_1285;
	input x_1286;
	input x_1287;
	input x_1288;
	input x_1289;
	input x_1290;
	input x_1291;
	input x_1292;
	input x_1293;
	input x_1294;
	input x_1295;
	input x_1296;
	input x_1297;
	input x_1298;
	input x_1299;
	input x_1300;
	input x_1301;
	input x_1302;
	input x_1303;
	input x_1304;
	input x_1305;
	input x_1306;
	input x_1307;
	input x_1308;
	input x_1309;
	input x_1310;
	input x_1311;
	input x_1312;
	input x_1313;
	input x_1314;
	input x_1315;
	input x_1316;
	input x_1317;
	input x_1318;
	input x_1319;
	input x_1320;
	input x_1321;
	input x_1322;
	input x_1323;
	input x_1324;
	input x_1325;
	input x_1326;
	input x_1327;
	input x_1328;
	input x_1329;
	input x_1330;
	input x_1331;
	input x_1332;
	input x_1333;
	input x_1334;
	input x_1335;
	input x_1336;
	input x_1337;
	input x_1338;
	input x_1339;
	input x_1340;
	input x_1341;
	input x_1342;
	input x_1343;
	input x_1344;
	input x_1345;
	input x_1346;
	input x_1347;
	input x_1348;
	input x_1349;
	input x_1350;
	input x_1351;
	input x_1352;
	input x_1353;
	input x_1354;
	input x_1355;
	input x_1356;
	input x_1357;
	input x_1358;
	input x_1359;
	input x_1360;
	input x_1361;
	input x_1362;
	input x_1363;
	input x_1364;
	input x_1365;
	input x_1366;
	input x_1367;
	input x_1368;
	input x_1369;
	input x_1370;
	input x_1371;
	input x_1372;
	input x_1373;
	input x_1374;
	input x_1375;
	input x_1376;
	input x_1377;
	input x_1378;
	input x_1379;
	input x_1380;
	input x_1381;
	input x_1382;
	input x_1383;
	input x_1384;
	input x_1385;
	input x_1386;
	input x_1387;
	input x_1388;
	input x_1389;
	input x_1390;
	input x_1391;
	input x_1392;
	input x_1393;
	input x_1394;
	input x_1395;
	input x_1396;
	input x_1397;
	input x_1398;
	input x_1399;
	input x_1400;
	input x_1401;
	input x_1402;
	input x_1403;
	input x_1404;
	input x_1405;
	input x_1406;
	input x_1407;
	input x_1408;
	input x_1409;
	input x_1410;
	input x_1411;
	input x_1412;
	input x_1413;
	input x_1414;
	input x_1415;
	input x_1416;
	input x_1417;
	input x_1418;
	input x_1419;
	input x_1420;
	input x_1421;
	input x_1422;
	input x_1423;
	input x_1424;
	input x_1425;
	input x_1426;
	input x_1427;
	input x_1428;
	input x_1429;
	input x_1430;
	input x_1431;
	input x_1432;
	input x_1433;
	input x_1434;
	input x_1435;
	input x_1436;
	input x_1437;
	input x_1438;
	input x_1439;
	input x_1440;
	input x_1441;
	input x_1442;
	input x_1443;
	input x_1444;
	input x_1445;
	input x_1446;
	input x_1447;
	input x_1448;
	input x_1449;
	input x_1450;
	input x_1451;
	input x_1452;
	input x_1453;
	input x_1454;
	input x_1455;
	input x_1456;
	input x_1457;
	input x_1458;
	input x_1459;
	input x_1460;
	input x_1461;
	input x_1462;
	input x_1463;
	input x_1464;
	input x_1465;
	input x_1466;
	input x_1467;
	input x_1468;
	input x_1469;
	input x_1470;
	input x_1471;
	input x_1472;
	input x_1473;
	input x_1474;
	input x_1475;
	input x_1476;
	input x_1477;
	input x_1478;
	input x_1479;
	input x_1480;
	input x_1481;
	input x_1482;
	input x_1483;
	input x_1484;
	input x_1485;
	input x_1486;
	input x_1487;
	input x_1488;
	input x_1489;
	input x_1490;
	input x_1491;
	input x_1492;
	input x_1493;
	input x_1494;
	input x_1495;
	input x_1496;
	input x_1497;
	input x_1498;
	input x_1499;
	input x_1500;
	input x_1501;
	input x_1502;
	input x_1503;
	input x_1504;
	input x_1505;
	input x_1506;
	input x_1507;
	input x_1508;
	input x_1509;
	input x_1510;
	input x_1511;
	input x_1512;
	input x_1513;
	input x_1514;
	input x_1515;
	input x_1516;
	input x_1517;
	input x_1518;
	input x_1519;
	input x_1520;
	input x_1521;
	input x_1522;
	input x_1523;
	input x_1524;
	input x_1525;
	input x_1526;
	input x_1527;
	input x_1528;
	input x_1529;
	input x_1530;
	input x_1531;
	input x_1532;
	input x_1533;
	input x_1534;
	input x_1535;
	input x_1536;
	input x_1537;
	input x_1538;
	input x_1539;
	input x_1540;
	input x_1541;
	input x_1542;
	input x_1543;
	input x_1544;
	input x_1545;
	input x_1546;
	input x_1547;
	input x_1548;
	input x_1549;
	input x_1550;
	input x_1551;
	input x_1552;
	input x_1553;
	input x_1554;
	input x_1555;
	input x_1556;
	input x_1557;
	input x_1558;
	input x_1559;
	input x_1560;
	input x_1561;
	input x_1562;
	input x_1563;
	input x_1564;
	input x_1565;
	input x_1566;
	input x_1567;
	input x_1568;
	input x_1569;
	input x_1570;
	input x_1571;
	input x_1572;
	input x_1573;
	input x_1574;
	input x_1575;
	input x_1576;
	input x_1577;
	input x_1578;
	wire n_1;
	wire n_2;
	wire n_3;
	wire n_4;
	wire n_5;
	wire n_6;
	wire n_7;
	wire n_8;
	wire n_9;
	wire n_10;
	wire n_11;
	wire n_12;
	wire n_13;
	wire n_14;
	wire n_15;
	wire n_16;
	wire n_17;
	wire n_18;
	wire n_19;
	wire n_20;
	wire n_21;
	wire n_22;
	wire n_23;
	wire n_24;
	wire n_25;
	wire n_26;
	wire n_27;
	wire n_28;
	wire n_29;
	wire n_30;
	wire n_31;
	wire n_32;
	wire n_33;
	wire n_34;
	wire n_35;
	wire n_36;
	wire n_37;
	wire n_38;
	wire n_39;
	wire n_40;
	wire n_41;
	wire n_42;
	wire n_43;
	wire n_44;
	wire n_45;
	wire n_46;
	wire n_47;
	wire n_48;
	wire n_49;
	wire n_50;
	wire n_51;
	wire n_52;
	wire n_53;
	wire n_54;
	wire n_55;
	wire n_56;
	wire n_57;
	wire n_58;
	wire n_59;
	wire n_60;
	wire n_61;
	wire n_62;
	wire n_63;
	wire n_64;
	wire n_65;
	wire n_66;
	wire n_67;
	wire n_68;
	wire n_69;
	wire n_70;
	wire n_71;
	wire n_72;
	wire n_73;
	wire n_74;
	wire n_75;
	wire n_76;
	wire n_77;
	wire n_78;
	wire n_79;
	wire n_80;
	wire n_81;
	wire n_82;
	wire n_83;
	wire n_84;
	wire n_85;
	wire n_86;
	wire n_87;
	wire n_88;
	wire n_89;
	wire n_90;
	wire n_91;
	wire n_92;
	wire n_93;
	wire n_94;
	wire n_95;
	wire n_96;
	wire n_97;
	wire n_98;
	wire n_99;
	wire n_100;
	wire n_101;
	wire n_102;
	wire n_103;
	wire n_104;
	wire n_105;
	wire n_106;
	wire n_107;
	wire n_108;
	wire n_109;
	wire n_110;
	wire n_111;
	wire n_112;
	wire n_113;
	wire n_114;
	wire n_115;
	wire n_116;
	wire n_117;
	wire n_118;
	wire n_119;
	wire n_120;
	wire n_121;
	wire n_122;
	wire n_123;
	wire n_124;
	wire n_125;
	wire n_126;
	wire n_127;
	wire n_128;
	wire n_129;
	wire n_130;
	wire n_131;
	wire n_132;
	wire n_133;
	wire n_134;
	wire n_135;
	wire n_136;
	wire n_137;
	wire n_138;
	wire n_139;
	wire n_140;
	wire n_141;
	wire n_142;
	wire n_143;
	wire n_144;
	wire n_145;
	wire n_146;
	wire n_147;
	wire n_148;
	wire n_149;
	wire n_150;
	wire n_151;
	wire n_152;
	wire n_153;
	wire n_154;
	wire n_155;
	wire n_156;
	wire n_157;
	wire n_158;
	wire n_159;
	wire n_160;
	wire n_161;
	wire n_162;
	wire n_163;
	wire n_164;
	wire n_165;
	wire n_166;
	wire n_167;
	wire n_168;
	wire n_169;
	wire n_170;
	wire n_171;
	wire n_172;
	wire n_173;
	wire n_174;
	wire n_175;
	wire n_176;
	wire n_177;
	wire n_178;
	wire n_179;
	wire n_180;
	wire n_181;
	wire n_182;
	wire n_183;
	wire n_184;
	wire n_185;
	wire n_186;
	wire n_187;
	wire n_188;
	wire n_189;
	wire n_190;
	wire n_191;
	wire n_192;
	wire n_193;
	wire n_194;
	wire n_195;
	wire n_196;
	wire n_197;
	wire n_198;
	wire n_199;
	wire n_200;
	wire n_201;
	wire n_202;
	wire n_203;
	wire n_204;
	wire n_205;
	wire n_206;
	wire n_207;
	wire n_208;
	wire n_209;
	wire n_210;
	wire n_211;
	wire n_212;
	wire n_213;
	wire n_214;
	wire n_215;
	wire n_216;
	wire n_217;
	wire n_218;
	wire n_219;
	wire n_220;
	wire n_221;
	wire n_222;
	wire n_223;
	wire n_224;
	wire n_225;
	wire n_226;
	wire n_227;
	wire n_228;
	wire n_229;
	wire n_230;
	wire n_231;
	wire n_232;
	wire n_233;
	wire n_234;
	wire n_235;
	wire n_236;
	wire n_237;
	wire n_238;
	wire n_239;
	wire n_240;
	wire n_241;
	wire n_242;
	wire n_243;
	wire n_244;
	wire n_245;
	wire n_246;
	wire n_247;
	wire n_248;
	wire n_249;
	wire n_250;
	wire n_251;
	wire n_252;
	wire n_253;
	wire n_254;
	wire n_255;
	wire n_256;
	wire n_257;
	wire n_258;
	wire n_259;
	wire n_260;
	wire n_261;
	wire n_262;
	wire n_263;
	wire n_264;
	wire n_265;
	wire n_266;
	wire n_267;
	wire n_268;
	wire n_269;
	wire n_270;
	wire n_271;
	wire n_272;
	wire n_273;
	wire n_274;
	wire n_275;
	wire n_276;
	wire n_277;
	wire n_278;
	wire n_279;
	wire n_280;
	wire n_281;
	wire n_282;
	wire n_283;
	wire n_284;
	wire n_285;
	wire n_286;
	wire n_287;
	wire n_288;
	wire n_289;
	wire n_290;
	wire n_291;
	wire n_292;
	wire n_293;
	wire n_294;
	wire n_295;
	wire n_296;
	wire n_297;
	wire n_298;
	wire n_299;
	wire n_300;
	wire n_301;
	wire n_302;
	wire n_303;
	wire n_304;
	wire n_305;
	wire n_306;
	wire n_307;
	wire n_308;
	wire n_309;
	wire n_310;
	wire n_311;
	wire n_312;
	wire n_313;
	wire n_314;
	wire n_315;
	wire n_316;
	wire n_317;
	wire n_318;
	wire n_319;
	wire n_320;
	wire n_321;
	wire n_322;
	wire n_323;
	wire n_324;
	wire n_325;
	wire n_326;
	wire n_327;
	wire n_328;
	wire n_329;
	wire n_330;
	wire n_331;
	wire n_332;
	wire n_333;
	wire n_334;
	wire n_335;
	wire n_336;
	wire n_337;
	wire n_338;
	wire n_339;
	wire n_340;
	wire n_341;
	wire n_342;
	wire n_343;
	wire n_344;
	wire n_345;
	wire n_346;
	wire n_347;
	wire n_348;
	wire n_349;
	wire n_350;
	wire n_351;
	wire n_352;
	wire n_353;
	wire n_354;
	wire n_355;
	wire n_356;
	wire n_357;
	wire n_358;
	wire n_359;
	wire n_360;
	wire n_361;
	wire n_362;
	wire n_363;
	wire n_364;
	wire n_365;
	wire n_366;
	wire n_367;
	wire n_368;
	wire n_369;
	wire n_370;
	wire n_371;
	wire n_372;
	wire n_373;
	wire n_374;
	wire n_375;
	wire n_376;
	wire n_377;
	wire n_378;
	wire n_379;
	wire n_380;
	wire n_381;
	wire n_382;
	wire n_383;
	wire n_384;
	wire n_385;
	wire n_386;
	wire n_387;
	wire n_388;
	wire n_389;
	wire n_390;
	wire n_391;
	wire n_392;
	wire n_393;
	wire n_394;
	wire n_395;
	wire n_396;
	wire n_397;
	wire n_398;
	wire n_399;
	wire n_400;
	wire n_401;
	wire n_402;
	wire n_403;
	wire n_404;
	wire n_405;
	wire n_406;
	wire n_407;
	wire n_408;
	wire n_409;
	wire n_410;
	wire n_411;
	wire n_412;
	wire n_413;
	wire n_414;
	wire n_415;
	wire n_416;
	wire n_417;
	wire n_418;
	wire n_419;
	wire n_420;
	wire n_421;
	wire n_422;
	wire n_423;
	wire n_424;
	wire n_425;
	wire n_426;
	wire n_427;
	wire n_428;
	wire n_429;
	wire n_430;
	wire n_431;
	wire n_432;
	wire n_433;
	wire n_434;
	wire n_435;
	wire n_436;
	wire n_437;
	wire n_438;
	wire n_439;
	wire n_440;
	wire n_441;
	wire n_442;
	wire n_443;
	wire n_444;
	wire n_445;
	wire n_446;
	wire n_447;
	wire n_448;
	wire n_449;
	wire n_450;
	wire n_451;
	wire n_452;
	wire n_453;
	wire n_454;
	wire n_455;
	wire n_456;
	wire n_457;
	wire n_458;
	wire n_459;
	wire n_460;
	wire n_461;
	wire n_462;
	wire n_463;
	wire n_464;
	wire n_465;
	wire n_466;
	wire n_467;
	wire n_468;
	wire n_469;
	wire n_470;
	wire n_471;
	wire n_472;
	wire n_473;
	wire n_474;
	wire n_475;
	wire n_476;
	wire n_477;
	wire n_478;
	wire n_479;
	wire n_480;
	wire n_481;
	wire n_482;
	wire n_483;
	wire n_484;
	wire n_485;
	wire n_486;
	wire n_487;
	wire n_488;
	wire n_489;
	wire n_490;
	wire n_491;
	wire n_492;
	wire n_493;
	wire n_494;
	wire n_495;
	wire n_496;
	wire n_497;
	wire n_498;
	wire n_499;
	wire n_500;
	wire n_501;
	wire n_502;
	wire n_503;
	wire n_504;
	wire n_505;
	wire n_506;
	wire n_507;
	wire n_508;
	wire n_509;
	wire n_510;
	wire n_511;
	wire n_512;
	wire n_513;
	wire n_514;
	wire n_515;
	wire n_516;
	wire n_517;
	wire n_518;
	wire n_519;
	wire n_520;
	wire n_521;
	wire n_522;
	wire n_523;
	wire n_524;
	wire n_525;
	wire n_526;
	wire n_527;
	wire n_528;
	wire n_529;
	wire n_530;
	wire n_531;
	wire n_532;
	wire n_533;
	wire n_534;
	wire n_535;
	wire n_536;
	wire n_537;
	wire n_538;
	wire n_539;
	wire n_540;
	wire n_541;
	wire n_542;
	wire n_543;
	wire n_544;
	wire n_545;
	wire n_546;
	wire n_547;
	wire n_548;
	wire n_549;
	wire n_550;
	wire n_551;
	wire n_552;
	wire n_553;
	wire n_554;
	wire n_555;
	wire n_556;
	wire n_557;
	wire n_558;
	wire n_559;
	wire n_560;
	wire n_561;
	wire n_562;
	wire n_563;
	wire n_564;
	wire n_565;
	wire n_566;
	wire n_567;
	wire n_568;
	wire n_569;
	wire n_570;
	wire n_571;
	wire n_572;
	wire n_573;
	wire n_574;
	wire n_575;
	wire n_576;
	wire n_577;
	wire n_578;
	wire n_579;
	wire n_580;
	wire n_581;
	wire n_582;
	wire n_583;
	wire n_584;
	wire n_585;
	wire n_586;
	wire n_587;
	wire n_588;
	wire n_589;
	wire n_590;
	wire n_591;
	wire n_592;
	wire n_593;
	wire n_594;
	wire n_595;
	wire n_596;
	wire n_597;
	wire n_598;
	wire n_599;
	wire n_600;
	wire n_601;
	wire n_602;
	wire n_603;
	wire n_604;
	wire n_605;
	wire n_606;
	wire n_607;
	wire n_608;
	wire n_609;
	wire n_610;
	wire n_611;
	wire n_612;
	wire n_613;
	wire n_614;
	wire n_615;
	wire n_616;
	wire n_617;
	wire n_618;
	wire n_619;
	wire n_620;
	wire n_621;
	wire n_622;
	wire n_623;
	wire n_624;
	wire n_625;
	wire n_626;
	wire n_627;
	wire n_628;
	wire n_629;
	wire n_630;
	wire n_631;
	wire n_632;
	wire n_633;
	wire n_634;
	wire n_635;
	wire n_636;
	wire n_637;
	wire n_638;
	wire n_639;
	wire n_640;
	wire n_641;
	wire n_642;
	wire n_643;
	wire n_644;
	wire n_645;
	wire n_646;
	wire n_647;
	wire n_648;
	wire n_649;
	wire n_650;
	wire n_651;
	wire n_652;
	wire n_653;
	wire n_654;
	wire n_655;
	wire n_656;
	wire n_657;
	wire n_658;
	wire n_659;
	wire n_660;
	wire n_661;
	wire n_662;
	wire n_663;
	wire n_664;
	wire n_665;
	wire n_666;
	wire n_667;
	wire n_668;
	wire n_669;
	wire n_670;
	wire n_671;
	wire n_672;
	wire n_673;
	wire n_674;
	wire n_675;
	wire n_676;
	wire n_677;
	wire n_678;
	wire n_679;
	wire n_680;
	wire n_681;
	wire n_682;
	wire n_683;
	wire n_684;
	wire n_685;
	wire n_686;
	wire n_687;
	wire n_688;
	wire n_689;
	wire n_690;
	wire n_691;
	wire n_692;
	wire n_693;
	wire n_694;
	wire n_695;
	wire n_696;
	wire n_697;
	wire n_698;
	wire n_699;
	wire n_700;
	wire n_701;
	wire n_702;
	wire n_703;
	wire n_704;
	wire n_705;
	wire n_706;
	wire n_707;
	wire n_708;
	wire n_709;
	wire n_710;
	wire n_711;
	wire n_712;
	wire n_713;
	wire n_714;
	wire n_715;
	wire n_716;
	wire n_717;
	wire n_718;
	wire n_719;
	wire n_720;
	wire n_721;
	wire n_722;
	wire n_723;
	wire n_724;
	wire n_725;
	wire n_726;
	wire n_727;
	wire n_728;
	wire n_729;
	wire n_730;
	wire n_731;
	wire n_732;
	wire n_733;
	wire n_734;
	wire n_735;
	wire n_736;
	wire n_737;
	wire n_738;
	wire n_739;
	wire n_740;
	wire n_741;
	wire n_742;
	wire n_743;
	wire n_744;
	wire n_745;
	wire n_746;
	wire n_747;
	wire n_748;
	wire n_749;
	wire n_750;
	wire n_751;
	wire n_752;
	wire n_753;
	wire n_754;
	wire n_755;
	wire n_756;
	wire n_757;
	wire n_758;
	wire n_759;
	wire n_760;
	wire n_761;
	wire n_762;
	wire n_763;
	wire n_764;
	wire n_765;
	wire n_766;
	wire n_767;
	wire n_768;
	wire n_769;
	wire n_770;
	wire n_771;
	wire n_772;
	wire n_773;
	wire n_774;
	wire n_775;
	wire n_776;
	wire n_777;
	wire n_778;
	wire n_779;
	wire n_780;
	wire n_781;
	wire n_782;
	wire n_783;
	wire n_784;
	wire n_785;
	wire n_786;
	wire n_787;
	wire n_788;
	wire n_789;
	wire n_790;
	wire n_791;
	wire n_792;
	wire n_793;
	wire n_794;
	wire n_795;
	wire n_796;
	wire n_797;
	wire n_798;
	wire n_799;
	wire n_800;
	wire n_801;
	wire n_802;
	wire n_803;
	wire n_804;
	wire n_805;
	wire n_806;
	wire n_807;
	wire n_808;
	wire n_809;
	wire n_810;
	wire n_811;
	wire n_812;
	wire n_813;
	wire n_814;
	wire n_815;
	wire n_816;
	wire n_817;
	wire n_818;
	wire n_819;
	wire n_820;
	wire n_821;
	wire n_822;
	wire n_823;
	wire n_824;
	wire n_825;
	wire n_826;
	wire n_827;
	wire n_828;
	wire n_829;
	wire n_830;
	wire n_831;
	wire n_832;
	wire n_833;
	wire n_834;
	wire n_835;
	wire n_836;
	wire n_837;
	wire n_838;
	wire n_839;
	wire n_840;
	wire n_841;
	wire n_842;
	wire n_843;
	wire n_844;
	wire n_845;
	wire n_846;
	wire n_847;
	wire n_848;
	wire n_849;
	wire n_850;
	wire n_851;
	wire n_852;
	wire n_853;
	wire n_854;
	wire n_855;
	wire n_856;
	wire n_857;
	wire n_858;
	wire n_859;
	wire n_860;
	wire n_861;
	wire n_862;
	wire n_863;
	wire n_864;
	wire n_865;
	wire n_866;
	wire n_867;
	wire n_868;
	wire n_869;
	wire n_870;
	wire n_871;
	wire n_872;
	wire n_873;
	wire n_874;
	wire n_875;
	wire n_876;
	wire n_877;
	wire n_878;
	wire n_879;
	wire n_880;
	wire n_881;
	wire n_882;
	wire n_883;
	wire n_884;
	wire n_885;
	wire n_886;
	wire n_887;
	wire n_888;
	wire n_889;
	wire n_890;
	wire n_891;
	wire n_892;
	wire n_893;
	wire n_894;
	wire n_895;
	wire n_896;
	wire n_897;
	wire n_898;
	wire n_899;
	wire n_900;
	wire n_901;
	wire n_902;
	wire n_903;
	wire n_904;
	wire n_905;
	wire n_906;
	wire n_907;
	wire n_908;
	wire n_909;
	wire n_910;
	wire n_911;
	wire n_912;
	wire n_913;
	wire n_914;
	wire n_915;
	wire n_916;
	wire n_917;
	wire n_918;
	wire n_919;
	wire n_920;
	wire n_921;
	wire n_922;
	wire n_923;
	wire n_924;
	wire n_925;
	wire n_926;
	wire n_927;
	wire n_928;
	wire n_929;
	wire n_930;
	wire n_931;
	wire n_932;
	wire n_933;
	wire n_934;
	wire n_935;
	wire n_936;
	wire n_937;
	wire n_938;
	wire n_939;
	wire n_940;
	wire n_941;
	wire n_942;
	wire n_943;
	wire n_944;
	wire n_945;
	wire n_946;
	wire n_947;
	wire n_948;
	wire n_949;
	wire n_950;
	wire n_951;
	wire n_952;
	wire n_953;
	wire n_954;
	wire n_955;
	wire n_956;
	wire n_957;
	wire n_958;
	wire n_959;
	wire n_960;
	wire n_961;
	wire n_962;
	wire n_963;
	wire n_964;
	wire n_965;
	wire n_966;
	wire n_967;
	wire n_968;
	wire n_969;
	wire n_970;
	wire n_971;
	wire n_972;
	wire n_973;
	wire n_974;
	wire n_975;
	wire n_976;
	wire n_977;
	wire n_978;
	wire n_979;
	wire n_980;
	wire n_981;
	wire n_982;
	wire n_983;
	wire n_984;
	wire n_985;
	wire n_986;
	wire n_987;
	wire n_988;
	wire n_989;
	wire n_990;
	wire n_991;
	wire n_992;
	wire n_993;
	wire n_994;
	wire n_995;
	wire n_996;
	wire n_997;
	wire n_998;
	wire n_999;
	wire n_1000;
	wire n_1001;
	wire n_1002;
	wire n_1003;
	wire n_1004;
	wire n_1005;
	wire n_1006;
	wire n_1007;
	wire n_1008;
	wire n_1009;
	wire n_1010;
	wire n_1011;
	wire n_1012;
	wire n_1013;
	wire n_1014;
	wire n_1015;
	wire n_1016;
	wire n_1017;
	wire n_1018;
	wire n_1019;
	wire n_1020;
	wire n_1021;
	wire n_1022;
	wire n_1023;
	wire n_1024;
	wire n_1025;
	wire n_1026;
	wire n_1027;
	wire n_1028;
	wire n_1029;
	wire n_1030;
	wire n_1031;
	wire n_1032;
	wire n_1033;
	wire n_1034;
	wire n_1035;
	wire n_1036;
	wire n_1037;
	wire n_1038;
	wire n_1039;
	wire n_1040;
	wire n_1041;
	wire n_1042;
	wire n_1043;
	wire n_1044;
	wire n_1045;
	wire n_1046;
	wire n_1047;
	wire n_1048;
	wire n_1049;
	wire n_1050;
	wire n_1051;
	wire n_1052;
	wire n_1053;
	wire n_1054;
	wire n_1055;
	wire n_1056;
	wire n_1057;
	wire n_1058;
	wire n_1059;
	wire n_1060;
	wire n_1061;
	wire n_1062;
	wire n_1063;
	wire n_1064;
	wire n_1065;
	wire n_1066;
	wire n_1067;
	wire n_1068;
	wire n_1069;
	wire n_1070;
	wire n_1071;
	wire n_1072;
	wire n_1073;
	wire n_1074;
	wire n_1075;
	wire n_1076;
	wire n_1077;
	wire n_1078;
	wire n_1079;
	wire n_1080;
	wire n_1081;
	wire n_1082;
	wire n_1083;
	wire n_1084;
	wire n_1085;
	wire n_1086;
	wire n_1087;
	wire n_1088;
	wire n_1089;
	wire n_1090;
	wire n_1091;
	wire n_1092;
	wire n_1093;
	wire n_1094;
	wire n_1095;
	wire n_1096;
	wire n_1097;
	wire n_1098;
	wire n_1099;
	wire n_1100;
	wire n_1101;
	wire n_1102;
	wire n_1103;
	wire n_1104;
	wire n_1105;
	wire n_1106;
	wire n_1107;
	wire n_1108;
	wire n_1109;
	wire n_1110;
	wire n_1111;
	wire n_1112;
	wire n_1113;
	wire n_1114;
	wire n_1115;
	wire n_1116;
	wire n_1117;
	wire n_1118;
	wire n_1119;
	wire n_1120;
	wire n_1121;
	wire n_1122;
	wire n_1123;
	wire n_1124;
	wire n_1125;
	wire n_1126;
	wire n_1127;
	wire n_1128;
	wire n_1129;
	wire n_1130;
	wire n_1131;
	wire n_1132;
	wire n_1133;
	wire n_1134;
	wire n_1135;
	wire n_1136;
	wire n_1137;
	wire n_1138;
	wire n_1139;
	wire n_1140;
	wire n_1141;
	wire n_1142;
	wire n_1143;
	wire n_1144;
	wire n_1145;
	wire n_1146;
	wire n_1147;
	wire n_1148;
	wire n_1149;
	wire n_1150;
	wire n_1151;
	wire n_1152;
	wire n_1153;
	wire n_1154;
	wire n_1155;
	wire n_1156;
	wire n_1157;
	wire n_1158;
	wire n_1159;
	wire n_1160;
	wire n_1161;
	wire n_1162;
	wire n_1163;
	wire n_1164;
	wire n_1165;
	wire n_1166;
	wire n_1167;
	wire n_1168;
	wire n_1169;
	wire n_1170;
	wire n_1171;
	wire n_1172;
	wire n_1173;
	wire n_1174;
	wire n_1175;
	wire n_1176;
	wire n_1177;
	wire n_1178;
	wire n_1179;
	wire n_1180;
	wire n_1181;
	wire n_1182;
	wire n_1183;
	wire n_1184;
	wire n_1185;
	wire n_1186;
	wire n_1187;
	wire n_1188;
	wire n_1189;
	wire n_1190;
	wire n_1191;
	wire n_1192;
	wire n_1193;
	wire n_1194;
	wire n_1195;
	wire n_1196;
	wire n_1197;
	wire n_1198;
	wire n_1199;
	wire n_1200;
	wire n_1201;
	wire n_1202;
	wire n_1203;
	wire n_1204;
	wire n_1205;
	wire n_1206;
	wire n_1207;
	wire n_1208;
	wire n_1209;
	wire n_1210;
	wire n_1211;
	wire n_1212;
	wire n_1213;
	wire n_1214;
	wire n_1215;
	wire n_1216;
	wire n_1217;
	wire n_1218;
	wire n_1219;
	wire n_1220;
	wire n_1221;
	wire n_1222;
	wire n_1223;
	wire n_1224;
	wire n_1225;
	wire n_1226;
	wire n_1227;
	wire n_1228;
	wire n_1229;
	wire n_1230;
	wire n_1231;
	wire n_1232;
	wire n_1233;
	wire n_1234;
	wire n_1235;
	wire n_1236;
	wire n_1237;
	wire n_1238;
	wire n_1239;
	wire n_1240;
	wire n_1241;
	wire n_1242;
	wire n_1243;
	wire n_1244;
	wire n_1245;
	wire n_1246;
	wire n_1247;
	wire n_1248;
	wire n_1249;
	wire n_1250;
	wire n_1251;
	wire n_1252;
	wire n_1253;
	wire n_1254;
	wire n_1255;
	wire n_1256;
	wire n_1257;
	wire n_1258;
	wire n_1259;
	wire n_1260;
	wire n_1261;
	wire n_1262;
	wire n_1263;
	wire n_1264;
	wire n_1265;
	wire n_1266;
	wire n_1267;
	wire n_1268;
	wire n_1269;
	wire n_1270;
	wire n_1271;
	wire n_1272;
	wire n_1273;
	wire n_1274;
	wire n_1275;
	wire n_1276;
	wire n_1277;
	wire n_1278;
	wire n_1279;
	wire n_1280;
	wire n_1281;
	wire n_1282;
	wire n_1283;
	wire n_1284;
	wire n_1285;
	wire n_1286;
	wire n_1287;
	wire n_1288;
	wire n_1289;
	wire n_1290;
	wire n_1291;
	wire n_1292;
	wire n_1293;
	wire n_1294;
	wire n_1295;
	wire n_1296;
	wire n_1297;
	wire n_1298;
	wire n_1299;
	wire n_1300;
	wire n_1301;
	wire n_1302;
	wire n_1303;
	wire n_1304;
	wire n_1305;
	wire n_1306;
	wire n_1307;
	wire n_1308;
	wire n_1309;
	wire n_1310;
	wire n_1311;
	wire n_1312;
	wire n_1313;
	wire n_1314;
	wire n_1315;
	wire n_1316;
	wire n_1317;
	wire n_1318;
	wire n_1319;
	wire n_1320;
	wire n_1321;
	wire n_1322;
	wire n_1323;
	wire n_1324;
	wire n_1325;
	wire n_1326;
	wire n_1327;
	wire n_1328;
	wire n_1329;
	wire n_1330;
	wire n_1331;
	wire n_1332;
	wire n_1333;
	wire n_1334;
	wire n_1335;
	wire n_1336;
	wire n_1337;
	wire n_1338;
	wire n_1339;
	wire n_1340;
	wire n_1341;
	wire n_1342;
	wire n_1343;
	wire n_1344;
	wire n_1345;
	wire n_1346;
	wire n_1347;
	wire n_1348;
	wire n_1349;
	wire n_1350;
	wire n_1351;
	wire n_1352;
	wire n_1353;
	wire n_1354;
	wire n_1355;
	wire n_1356;
	wire n_1357;
	wire n_1358;
	wire n_1359;
	wire n_1360;
	wire n_1361;
	wire n_1362;
	wire n_1363;
	wire n_1364;
	wire n_1365;
	wire n_1366;
	wire n_1367;
	wire n_1368;
	wire n_1369;
	wire n_1370;
	wire n_1371;
	wire n_1372;
	wire n_1373;
	wire n_1374;
	wire n_1375;
	wire n_1376;
	wire n_1377;
	wire n_1378;
	wire n_1379;
	wire n_1380;
	wire n_1381;
	wire n_1382;
	wire n_1383;
	wire n_1384;
	wire n_1385;
	wire n_1386;
	wire n_1387;
	wire n_1388;
	wire n_1389;
	wire n_1390;
	wire n_1391;
	wire n_1392;
	wire n_1393;
	wire n_1394;
	wire n_1395;
	wire n_1396;
	wire n_1397;
	wire n_1398;
	wire n_1399;
	wire n_1400;
	wire n_1401;
	wire n_1402;
	wire n_1403;
	wire n_1404;
	wire n_1405;
	wire n_1406;
	wire n_1407;
	wire n_1408;
	wire n_1409;
	wire n_1410;
	wire n_1411;
	wire n_1412;
	wire n_1413;
	wire n_1414;
	wire n_1415;
	wire n_1416;
	wire n_1417;
	wire n_1418;
	wire n_1419;
	wire n_1420;
	wire n_1421;
	wire n_1422;
	wire n_1423;
	wire n_1424;
	wire n_1425;
	wire n_1426;
	wire n_1427;
	wire n_1428;
	wire n_1429;
	wire n_1430;
	wire n_1431;
	wire n_1432;
	wire n_1433;
	wire n_1434;
	wire n_1435;
	wire n_1436;
	wire n_1437;
	wire n_1438;
	wire n_1439;
	wire n_1440;
	wire n_1441;
	wire n_1442;
	wire n_1443;
	wire n_1444;
	wire n_1445;
	wire n_1446;
	wire n_1447;
	wire n_1448;
	wire n_1449;
	wire n_1450;
	wire n_1451;
	wire n_1452;
	wire n_1453;
	wire n_1454;
	wire n_1455;
	wire n_1456;
	wire n_1457;
	wire n_1458;
	wire n_1459;
	wire n_1460;
	wire n_1461;
	wire n_1462;
	wire n_1463;
	wire n_1464;
	wire n_1465;
	wire n_1466;
	wire n_1467;
	wire n_1468;
	wire n_1469;
	wire n_1470;
	wire n_1471;
	wire n_1472;
	wire n_1473;
	wire n_1474;
	wire n_1475;
	wire n_1476;
	wire n_1477;
	wire n_1478;
	wire n_1479;
	wire n_1480;
	wire n_1481;
	wire n_1482;
	wire n_1483;
	wire n_1484;
	wire n_1485;
	wire n_1486;
	wire n_1487;
	wire n_1488;
	wire n_1489;
	wire n_1490;
	wire n_1491;
	wire n_1492;
	wire n_1493;
	wire n_1494;
	wire n_1495;
	wire n_1496;
	wire n_1497;
	wire n_1498;
	wire n_1499;
	wire n_1500;
	wire n_1501;
	wire n_1502;
	wire n_1503;
	wire n_1504;
	wire n_1505;
	wire n_1506;
	wire n_1507;
	wire n_1508;
	wire n_1509;
	wire n_1510;
	wire n_1511;
	wire n_1512;
	wire n_1513;
	wire n_1514;
	wire n_1515;
	wire n_1516;
	wire n_1517;
	wire n_1518;
	wire n_1519;
	wire n_1520;
	wire n_1521;
	wire n_1522;
	wire n_1523;
	wire n_1524;
	wire n_1525;
	wire n_1526;
	wire n_1527;
	wire n_1528;
	wire n_1529;
	wire n_1530;
	wire n_1531;
	wire n_1532;
	wire n_1533;
	wire n_1534;
	wire n_1535;
	wire n_1536;
	wire n_1537;
	wire n_1538;
	wire n_1539;
	wire n_1540;
	wire n_1541;
	wire n_1542;
	wire n_1543;
	wire n_1544;
	wire n_1545;
	wire n_1546;
	wire n_1547;
	wire n_1548;
	wire n_1549;
	wire n_1550;
	wire n_1551;
	wire n_1552;
	wire n_1553;
	wire n_1554;
	wire n_1555;
	wire n_1556;
	wire n_1557;
	wire n_1558;
	wire n_1559;
	wire n_1560;
	wire n_1561;
	wire n_1562;
	wire n_1563;
	wire n_1564;
	wire n_1565;
	wire n_1566;
	wire n_1567;
	wire n_1568;
	wire n_1569;
	wire n_1570;
	wire n_1571;
	wire n_1572;
	wire n_1573;
	wire n_1574;
	wire n_1575;
	wire n_1576;
	wire n_1577;
	wire n_1578;
	wire n_1579;
	wire n_1580;
	wire n_1581;
	wire n_1582;
	wire n_1583;
	wire n_1584;
	wire n_1585;
	wire n_1586;
	wire n_1587;
	wire n_1588;
	wire n_1589;
	wire n_1590;
	wire n_1591;
	wire n_1592;
	wire n_1593;
	wire n_1594;
	wire n_1595;
	wire n_1596;
	wire n_1597;
	wire n_1598;
	wire n_1599;
	wire n_1600;
	wire n_1601;
	wire n_1602;
	wire n_1603;
	wire n_1604;
	wire n_1605;
	wire n_1606;
	wire n_1607;
	wire n_1608;
	wire n_1609;
	wire n_1610;
	wire n_1611;
	wire n_1612;
	wire n_1613;
	wire n_1614;
	wire n_1615;
	wire n_1616;
	wire n_1617;
	wire n_1618;
	wire n_1619;
	wire n_1620;
	wire n_1621;
	wire n_1622;
	wire n_1623;
	wire n_1624;
	wire n_1625;
	wire n_1626;
	wire n_1627;
	wire n_1628;
	wire n_1629;
	wire n_1630;
	wire n_1631;
	wire n_1632;
	wire n_1633;
	wire n_1634;
	wire n_1635;
	wire n_1636;
	wire n_1637;
	wire n_1638;
	wire n_1639;
	wire n_1640;
	wire n_1641;
	wire n_1642;
	wire n_1643;
	wire n_1644;
	wire n_1645;
	wire n_1646;
	wire n_1647;
	wire n_1648;
	wire n_1649;
	wire n_1650;
	wire n_1651;
	wire n_1652;
	wire n_1653;
	wire n_1654;
	wire n_1655;
	wire n_1656;
	wire n_1657;
	wire n_1658;
	wire n_1659;
	wire n_1660;
	wire n_1661;
	wire n_1662;
	wire n_1663;
	wire n_1664;
	wire n_1665;
	wire n_1666;
	wire n_1667;
	wire n_1668;
	wire n_1669;
	wire n_1670;
	wire n_1671;
	wire n_1672;
	wire n_1673;
	wire n_1674;
	wire n_1675;
	wire n_1676;
	wire n_1677;
	wire n_1678;
	wire n_1679;
	wire n_1680;
	wire n_1681;
	wire n_1682;
	wire n_1683;
	wire n_1684;
	wire n_1685;
	wire n_1686;
	wire n_1687;
	wire n_1688;
	wire n_1689;
	wire n_1690;
	wire n_1691;
	wire n_1692;
	wire n_1693;
	wire n_1694;
	wire n_1695;
	wire n_1696;
	wire n_1697;
	wire n_1698;
	wire n_1699;
	wire n_1700;
	wire n_1701;
	wire n_1702;
	wire n_1703;
	wire n_1704;
	wire n_1705;
	wire n_1706;
	wire n_1707;
	wire n_1708;
	wire n_1709;
	wire n_1710;
	wire n_1711;
	wire n_1712;
	wire n_1713;
	wire n_1714;
	wire n_1715;
	wire n_1716;
	wire n_1717;
	wire n_1718;
	wire n_1719;
	wire n_1720;
	wire n_1721;
	wire n_1722;
	wire n_1723;
	wire n_1724;
	wire n_1725;
	wire n_1726;
	wire n_1727;
	wire n_1728;
	wire n_1729;
	wire n_1730;
	wire n_1731;
	wire n_1732;
	wire n_1733;
	wire n_1734;
	wire n_1735;
	wire n_1736;
	wire n_1737;
	wire n_1738;
	wire n_1739;
	wire n_1740;
	wire n_1741;
	wire n_1742;
	wire n_1743;
	wire n_1744;
	wire n_1745;
	wire n_1746;
	wire n_1747;
	wire n_1748;
	wire n_1749;
	wire n_1750;
	wire n_1751;
	wire n_1752;
	wire n_1753;
	wire n_1754;
	wire n_1755;
	wire n_1756;
	wire n_1757;
	wire n_1758;
	wire n_1759;
	wire n_1760;
	wire n_1761;
	wire n_1762;
	wire n_1763;
	wire n_1764;
	wire n_1765;
	wire n_1766;
	wire n_1767;
	wire n_1768;
	wire n_1769;
	wire n_1770;
	wire n_1771;
	wire n_1772;
	wire n_1773;
	wire n_1774;
	wire n_1775;
	wire n_1776;
	wire n_1777;
	wire n_1778;
	wire n_1779;
	wire n_1780;
	wire n_1781;
	wire n_1782;
	wire n_1783;
	wire n_1784;
	wire n_1785;
	wire n_1786;
	wire n_1787;
	wire n_1788;
	wire n_1789;
	wire n_1790;
	wire n_1791;
	wire n_1792;
	wire n_1793;
	wire n_1794;
	wire n_1795;
	wire n_1796;
	wire n_1797;
	wire n_1798;
	wire n_1799;
	wire n_1800;
	wire n_1801;
	wire n_1802;
	wire n_1803;
	wire n_1804;
	wire n_1805;
	wire n_1806;
	wire n_1807;
	wire n_1808;
	wire n_1809;
	wire n_1810;
	wire n_1811;
	wire n_1812;
	wire n_1813;
	wire n_1814;
	wire n_1815;
	wire n_1816;
	wire n_1817;
	wire n_1818;
	wire n_1819;
	wire n_1820;
	wire n_1821;
	wire n_1822;
	wire n_1823;
	wire n_1824;
	wire n_1825;
	wire n_1826;
	wire n_1827;
	wire n_1828;
	wire n_1829;
	wire n_1830;
	wire n_1831;
	wire n_1832;
	wire n_1833;
	wire n_1834;
	wire n_1835;
	wire n_1836;
	wire n_1837;
	wire n_1838;
	wire n_1839;
	wire n_1840;
	wire n_1841;
	wire n_1842;
	wire n_1843;
	wire n_1844;
	wire n_1845;
	wire n_1846;
	wire n_1847;
	wire n_1848;
	wire n_1849;
	wire n_1850;
	wire n_1851;
	wire n_1852;
	wire n_1853;
	wire n_1854;
	wire n_1855;
	wire n_1856;
	wire n_1857;
	wire n_1858;
	wire n_1859;
	wire n_1860;
	wire n_1861;
	wire n_1862;
	wire n_1863;
	wire n_1864;
	wire n_1865;
	wire n_1866;
	wire n_1867;
	wire n_1868;
	wire n_1869;
	wire n_1870;
	wire n_1871;
	wire n_1872;
	wire n_1873;
	wire n_1874;
	wire n_1875;
	wire n_1876;
	wire n_1877;
	wire n_1878;
	wire n_1879;
	wire n_1880;
	wire n_1881;
	wire n_1882;
	wire n_1883;
	wire n_1884;
	wire n_1885;
	wire n_1886;
	wire n_1887;
	wire n_1888;
	wire n_1889;
	wire n_1890;
	wire n_1891;
	wire n_1892;
	wire n_1893;
	wire n_1894;
	wire n_1895;
	wire n_1896;
	wire n_1897;
	wire n_1898;
	wire n_1899;
	wire n_1900;
	wire n_1901;
	wire n_1902;
	wire n_1903;
	wire n_1904;
	wire n_1905;
	wire n_1906;
	wire n_1907;
	wire n_1908;
	wire n_1909;
	wire n_1910;
	wire n_1911;
	wire n_1912;
	wire n_1913;
	wire n_1914;
	wire n_1915;
	wire n_1916;
	wire n_1917;
	wire n_1918;
	wire n_1919;
	wire n_1920;
	wire n_1921;
	wire n_1922;
	wire n_1923;
	wire n_1924;
	wire n_1925;
	wire n_1926;
	wire n_1927;
	wire n_1928;
	wire n_1929;
	wire n_1930;
	wire n_1931;
	wire n_1932;
	wire n_1933;
	wire n_1934;
	wire n_1935;
	wire n_1936;
	wire n_1937;
	wire n_1938;
	wire n_1939;
	wire n_1940;
	wire n_1941;
	wire n_1942;
	wire n_1943;
	wire n_1944;
	wire n_1945;
	wire n_1946;
	wire n_1947;
	wire n_1948;
	wire n_1949;
	wire n_1950;
	wire n_1951;
	wire n_1952;
	wire n_1953;
	wire n_1954;
	wire n_1955;
	wire n_1956;
	wire n_1957;
	wire n_1958;
	wire n_1959;
	wire n_1960;
	wire n_1961;
	wire n_1962;
	wire n_1963;
	wire n_1964;
	wire n_1965;
	wire n_1966;
	wire n_1967;
	wire n_1968;
	wire n_1969;
	wire n_1970;
	wire n_1971;
	wire n_1972;
	wire n_1973;
	wire n_1974;
	wire n_1975;
	wire n_1976;
	wire n_1977;
	wire n_1978;
	wire n_1979;
	wire n_1980;
	wire n_1981;
	wire n_1982;
	wire n_1983;
	wire n_1984;
	wire n_1985;
	wire n_1986;
	wire n_1987;
	wire n_1988;
	wire n_1989;
	wire n_1990;
	wire n_1991;
	wire n_1992;
	wire n_1993;
	wire n_1994;
	wire n_1995;
	wire n_1996;
	wire n_1997;
	wire n_1998;
	wire n_1999;
	wire n_2000;
	wire n_2001;
	wire n_2002;
	wire n_2003;
	wire n_2004;
	wire n_2005;
	wire n_2006;
	wire n_2007;
	wire n_2008;
	wire n_2009;
	wire n_2010;
	wire n_2011;
	wire n_2012;
	wire n_2013;
	wire n_2014;
	wire n_2015;
	wire n_2016;
	wire n_2017;
	wire n_2018;
	wire n_2019;
	wire n_2020;
	wire n_2021;
	wire n_2022;
	wire n_2023;
	wire n_2024;
	wire n_2025;
	wire n_2026;
	wire n_2027;
	wire n_2028;
	wire n_2029;
	wire n_2030;
	wire n_2031;
	wire n_2032;
	wire n_2033;
	wire n_2034;
	wire n_2035;
	wire n_2036;
	wire n_2037;
	wire n_2038;
	wire n_2039;
	wire n_2040;
	wire n_2041;
	wire n_2042;
	wire n_2043;
	wire n_2044;
	wire n_2045;
	wire n_2046;
	wire n_2047;
	wire n_2048;
	wire n_2049;
	wire n_2050;
	wire n_2051;
	wire n_2052;
	wire n_2053;
	wire n_2054;
	wire n_2055;
	wire n_2056;
	wire n_2057;
	wire n_2058;
	wire n_2059;
	wire n_2060;
	wire n_2061;
	wire n_2062;
	wire n_2063;
	wire n_2064;
	wire n_2065;
	wire n_2066;
	wire n_2067;
	wire n_2068;
	wire n_2069;
	wire n_2070;
	wire n_2071;
	wire n_2072;
	wire n_2073;
	wire n_2074;
	wire n_2075;
	wire n_2076;
	wire n_2077;
	wire n_2078;
	wire n_2079;
	wire n_2080;
	wire n_2081;
	wire n_2082;
	wire n_2083;
	wire n_2084;
	wire n_2085;
	wire n_2086;
	wire n_2087;
	wire n_2088;
	wire n_2089;
	wire n_2090;
	wire n_2091;
	wire n_2092;
	wire n_2093;
	wire n_2094;
	wire n_2095;
	wire n_2096;
	wire n_2097;
	wire n_2098;
	wire n_2099;
	wire n_2100;
	wire n_2101;
	wire n_2102;
	wire n_2103;
	wire n_2104;
	wire n_2105;
	wire n_2106;
	wire n_2107;
	wire n_2108;
	wire n_2109;
	wire n_2110;
	wire n_2111;
	wire n_2112;
	wire n_2113;
	wire n_2114;
	wire n_2115;
	wire n_2116;
	wire n_2117;
	wire n_2118;
	wire n_2119;
	wire n_2120;
	wire n_2121;
	wire n_2122;
	wire n_2123;
	wire n_2124;
	wire n_2125;
	wire n_2126;
	wire n_2127;
	wire n_2128;
	wire n_2129;
	wire n_2130;
	wire n_2131;
	wire n_2132;
	wire n_2133;
	wire n_2134;
	wire n_2135;
	wire n_2136;
	wire n_2137;
	wire n_2138;
	wire n_2139;
	wire n_2140;
	wire n_2141;
	wire n_2142;
	wire n_2143;
	wire n_2144;
	wire n_2145;
	wire n_2146;
	wire n_2147;
	wire n_2148;
	wire n_2149;
	wire n_2150;
	wire n_2151;
	wire n_2152;
	wire n_2153;
	wire n_2154;
	wire n_2155;
	wire n_2156;
	wire n_2157;
	wire n_2158;
	wire n_2159;
	wire n_2160;
	wire n_2161;
	wire n_2162;
	wire n_2163;
	wire n_2164;
	wire n_2165;
	wire n_2166;
	wire n_2167;
	wire n_2168;
	wire n_2169;
	wire n_2170;
	wire n_2171;
	wire n_2172;
	wire n_2173;
	wire n_2174;
	wire n_2175;
	wire n_2176;
	wire n_2177;
	wire n_2178;
	wire n_2179;
	wire n_2180;
	wire n_2181;
	wire n_2182;
	wire n_2183;
	wire n_2184;
	wire n_2185;
	wire n_2186;
	wire n_2187;
	wire n_2188;
	wire n_2189;
	wire n_2190;
	wire n_2191;
	wire n_2192;
	wire n_2193;
	wire n_2194;
	wire n_2195;
	wire n_2196;
	wire n_2197;
	wire n_2198;
	wire n_2199;
	wire n_2200;
	wire n_2201;
	wire n_2202;
	wire n_2203;
	wire n_2204;
	wire n_2205;
	wire n_2206;
	wire n_2207;
	wire n_2208;
	wire n_2209;
	wire n_2210;
	wire n_2211;
	wire n_2212;
	wire n_2213;
	wire n_2214;
	wire n_2215;
	wire n_2216;
	wire n_2217;
	wire n_2218;
	wire n_2219;
	wire n_2220;
	wire n_2221;
	wire n_2222;
	wire n_2223;
	wire n_2224;
	wire n_2225;
	wire n_2226;
	wire n_2227;
	wire n_2228;
	wire n_2229;
	wire n_2230;
	wire n_2231;
	wire n_2232;
	wire n_2233;
	wire n_2234;
	wire n_2235;
	wire n_2236;
	wire n_2237;
	wire n_2238;
	wire n_2239;
	wire n_2240;
	wire n_2241;
	wire n_2242;
	wire n_2243;
	wire n_2244;
	wire n_2245;
	wire n_2246;
	wire n_2247;
	wire n_2248;
	wire n_2249;
	wire n_2250;
	wire n_2251;
	wire n_2252;
	wire n_2253;
	wire n_2254;
	wire n_2255;
	wire n_2256;
	wire n_2257;
	wire n_2258;
	wire n_2259;
	wire n_2260;
	wire n_2261;
	wire n_2262;
	wire n_2263;
	wire n_2264;
	wire n_2265;
	wire n_2266;
	wire n_2267;
	wire n_2268;
	wire n_2269;
	wire n_2270;
	wire n_2271;
	wire n_2272;
	wire n_2273;
	wire n_2274;
	wire n_2275;
	wire n_2276;
	wire n_2277;
	wire n_2278;
	wire n_2279;
	wire n_2280;
	wire n_2281;
	wire n_2282;
	wire n_2283;
	wire n_2284;
	wire n_2285;
	wire n_2286;
	wire n_2287;
	wire n_2288;
	wire n_2289;
	wire n_2290;
	wire n_2291;
	wire n_2292;
	wire n_2293;
	wire n_2294;
	wire n_2295;
	wire n_2296;
	wire n_2297;
	wire n_2298;
	wire n_2299;
	wire n_2300;
	wire n_2301;
	wire n_2302;
	wire n_2303;
	wire n_2304;
	wire n_2305;
	wire n_2306;
	wire n_2307;
	wire n_2308;
	wire n_2309;
	wire n_2310;
	wire n_2311;
	wire n_2312;
	wire n_2313;
	wire n_2314;
	wire n_2315;
	wire n_2316;
	wire n_2317;
	wire n_2318;
	wire n_2319;
	wire n_2320;
	wire n_2321;
	wire n_2322;
	wire n_2323;
	wire n_2324;
	wire n_2325;
	wire n_2326;
	wire n_2327;
	wire n_2328;
	wire n_2329;
	wire n_2330;
	wire n_2331;
	wire n_2332;
	wire n_2333;
	wire n_2334;
	wire n_2335;
	wire n_2336;
	wire n_2337;
	wire n_2338;
	wire n_2339;
	wire n_2340;
	wire n_2341;
	wire n_2342;
	wire n_2343;
	wire n_2344;
	wire n_2345;
	wire n_2346;
	wire n_2347;
	wire n_2348;
	wire n_2349;
	wire n_2350;
	wire n_2351;
	wire n_2352;
	wire n_2353;
	wire n_2354;
	wire n_2355;
	wire n_2356;
	wire n_2357;
	wire n_2358;
	wire n_2359;
	wire n_2360;
	wire n_2361;
	wire n_2362;
	wire n_2363;
	wire n_2364;
	wire n_2365;
	wire n_2366;
	wire n_2367;
	wire n_2368;
	wire n_2369;
	wire n_2370;
	wire n_2371;
	wire n_2372;
	wire n_2373;
	wire n_2374;
	wire n_2375;
	wire n_2376;
	wire n_2377;
	wire n_2378;
	wire n_2379;
	wire n_2380;
	wire n_2381;
	wire n_2382;
	wire n_2383;
	wire n_2384;
	wire n_2385;
	wire n_2386;
	wire n_2387;
	wire n_2388;
	wire n_2389;
	wire n_2390;
	wire n_2391;
	wire n_2392;
	wire n_2393;
	wire n_2394;
	wire n_2395;
	wire n_2396;
	wire n_2397;
	wire n_2398;
	wire n_2399;
	wire n_2400;
	wire n_2401;
	wire n_2402;
	wire n_2403;
	wire n_2404;
	wire n_2405;
	wire n_2406;
	wire n_2407;
	wire n_2408;
	wire n_2409;
	wire n_2410;
	wire n_2411;
	wire n_2412;
	wire n_2413;
	wire n_2414;
	wire n_2415;
	wire n_2416;
	wire n_2417;
	wire n_2418;
	wire n_2419;
	wire n_2420;
	wire n_2421;
	wire n_2422;
	wire n_2423;
	wire n_2424;
	wire n_2425;
	wire n_2426;
	wire n_2427;
	wire n_2428;
	wire n_2429;
	wire n_2430;
	wire n_2431;
	wire n_2432;
	wire n_2433;
	wire n_2434;
	wire n_2435;
	wire n_2436;
	wire n_2437;
	wire n_2438;
	wire n_2439;
	wire n_2440;
	wire n_2441;
	wire n_2442;
	wire n_2443;
	wire n_2444;
	wire n_2445;
	wire n_2446;
	wire n_2447;
	wire n_2448;
	wire n_2449;
	wire n_2450;
	wire n_2451;
	wire n_2452;
	wire n_2453;
	wire n_2454;
	wire n_2455;
	wire n_2456;
	wire n_2457;
	wire n_2458;
	wire n_2459;
	wire n_2460;
	wire n_2461;
	wire n_2462;
	wire n_2463;
	wire n_2464;
	wire n_2465;
	wire n_2466;
	wire n_2467;
	wire n_2468;
	wire n_2469;
	wire n_2470;
	wire n_2471;
	wire n_2472;
	wire n_2473;
	wire n_2474;
	wire n_2475;
	wire n_2476;
	wire n_2477;
	wire n_2478;
	wire n_2479;
	wire n_2480;
	wire n_2481;
	wire n_2482;
	wire n_2483;
	wire n_2484;
	wire n_2485;
	wire n_2486;
	wire n_2487;
	wire n_2488;
	wire n_2489;
	wire n_2490;
	wire n_2491;
	wire n_2492;
	wire n_2493;
	wire n_2494;
	wire n_2495;
	wire n_2496;
	wire n_2497;
	wire n_2498;
	wire n_2499;
	wire n_2500;
	wire n_2501;
	wire n_2502;
	wire n_2503;
	wire n_2504;
	wire n_2505;
	wire n_2506;
	wire n_2507;
	wire n_2508;
	wire n_2509;
	wire n_2510;
	wire n_2511;
	wire n_2512;
	wire n_2513;
	wire n_2514;
	wire n_2515;
	wire n_2516;
	wire n_2517;
	wire n_2518;
	wire n_2519;
	wire n_2520;
	wire n_2521;
	wire n_2522;
	wire n_2523;
	wire n_2524;
	wire n_2525;
	wire n_2526;
	wire n_2527;
	wire n_2528;
	wire n_2529;
	wire n_2530;
	wire n_2531;
	wire n_2532;
	wire n_2533;
	wire n_2534;
	wire n_2535;
	wire n_2536;
	wire n_2537;
	wire n_2538;
	wire n_2539;
	wire n_2540;
	wire n_2541;
	wire n_2542;
	wire n_2543;
	wire n_2544;
	wire n_2545;
	wire n_2546;
	wire n_2547;
	wire n_2548;
	wire n_2549;
	wire n_2550;
	wire n_2551;
	wire n_2552;
	wire n_2553;
	wire n_2554;
	wire n_2555;
	wire n_2556;
	wire n_2557;
	wire n_2558;
	wire n_2559;
	wire n_2560;
	wire n_2561;
	wire n_2562;
	wire n_2563;
	wire n_2564;
	wire n_2565;
	wire n_2566;
	wire n_2567;
	wire n_2568;
	wire n_2569;
	wire n_2570;
	wire n_2571;
	wire n_2572;
	wire n_2573;
	wire n_2574;
	wire n_2575;
	wire n_2576;
	wire n_2577;
	wire n_2578;
	wire n_2579;
	wire n_2580;
	wire n_2581;
	wire n_2582;
	wire n_2583;
	wire n_2584;
	wire n_2585;
	wire n_2586;
	wire n_2587;
	wire n_2588;
	wire n_2589;
	wire n_2590;
	wire n_2591;
	wire n_2592;
	wire n_2593;
	wire n_2594;
	wire n_2595;
	wire n_2596;
	wire n_2597;
	wire n_2598;
	wire n_2599;
	wire n_2600;
	wire n_2601;
	wire n_2602;
	wire n_2603;
	wire n_2604;
	wire n_2605;
	wire n_2606;
	wire n_2607;
	wire n_2608;
	wire n_2609;
	wire n_2610;
	wire n_2611;
	wire n_2612;
	wire n_2613;
	wire n_2614;
	wire n_2615;
	wire n_2616;
	wire n_2617;
	wire n_2618;
	wire n_2619;
	wire n_2620;
	wire n_2621;
	wire n_2622;
	wire n_2623;
	wire n_2624;
	wire n_2625;
	wire n_2626;
	wire n_2627;
	wire n_2628;
	wire n_2629;
	wire n_2630;
	wire n_2631;
	wire n_2632;
	wire n_2633;
	wire n_2634;
	wire n_2635;
	wire n_2636;
	wire n_2637;
	wire n_2638;
	wire n_2639;
	wire n_2640;
	wire n_2641;
	wire n_2642;
	wire n_2643;
	wire n_2644;
	wire n_2645;
	wire n_2646;
	wire n_2647;
	wire n_2648;
	wire n_2649;
	wire n_2650;
	wire n_2651;
	wire n_2652;
	wire n_2653;
	wire n_2654;
	wire n_2655;
	wire n_2656;
	wire n_2657;
	wire n_2658;
	wire n_2659;
	wire n_2660;
	wire n_2661;
	wire n_2662;
	wire n_2663;
	wire n_2664;
	wire n_2665;
	wire n_2666;
	wire n_2667;
	wire n_2668;
	wire n_2669;
	wire n_2670;
	wire n_2671;
	wire n_2672;
	wire n_2673;
	wire n_2674;
	wire n_2675;
	wire n_2676;
	wire n_2677;
	wire n_2678;
	wire n_2679;
	wire n_2680;
	wire n_2681;
	wire n_2682;
	wire n_2683;
	wire n_2684;
	wire n_2685;
	wire n_2686;
	wire n_2687;
	wire n_2688;
	wire n_2689;
	wire n_2690;
	wire n_2691;
	wire n_2692;
	wire n_2693;
	wire n_2694;
	wire n_2695;
	wire n_2696;
	wire n_2697;
	wire n_2698;
	wire n_2699;
	wire n_2700;
	wire n_2701;
	wire n_2702;
	wire n_2703;
	wire n_2704;
	wire n_2705;
	wire n_2706;
	wire n_2707;
	wire n_2708;
	wire n_2709;
	wire n_2710;
	wire n_2711;
	wire n_2712;
	wire n_2713;
	wire n_2714;
	wire n_2715;
	wire n_2716;
	wire n_2717;
	wire n_2718;
	wire n_2719;
	wire n_2720;
	wire n_2721;
	wire n_2722;
	wire n_2723;
	wire n_2724;
	wire n_2725;
	wire n_2726;
	wire n_2727;
	wire n_2728;
	wire n_2729;
	wire n_2730;
	wire n_2731;
	wire n_2732;
	wire n_2733;
	wire n_2734;
	wire n_2735;
	wire n_2736;
	wire n_2737;
	wire n_2738;
	wire n_2739;
	wire n_2740;
	wire n_2741;
	wire n_2742;
	wire n_2743;
	wire n_2744;
	wire n_2745;
	wire n_2746;
	wire n_2747;
	wire n_2748;
	wire n_2749;
	wire n_2750;
	wire n_2751;
	wire n_2752;
	wire n_2753;
	wire n_2754;
	wire n_2755;
	wire n_2756;
	wire n_2757;
	wire n_2758;
	wire n_2759;
	wire n_2760;
	wire n_2761;
	wire n_2762;
	wire n_2763;
	wire n_2764;
	wire n_2765;
	wire n_2766;
	wire n_2767;
	wire n_2768;
	wire n_2769;
	wire n_2770;
	wire n_2771;
	wire n_2772;
	wire n_2773;
	wire n_2774;
	wire n_2775;
	wire n_2776;
	wire n_2777;
	wire n_2778;
	wire n_2779;
	wire n_2780;
	wire n_2781;
	wire n_2782;
	wire n_2783;
	wire n_2784;
	wire n_2785;
	wire n_2786;
	wire n_2787;
	wire n_2788;
	wire n_2789;
	wire n_2790;
	wire n_2791;
	wire n_2792;
	wire n_2793;
	wire n_2794;
	wire n_2795;
	wire n_2796;
	wire n_2797;
	wire n_2798;
	wire n_2799;
	wire n_2800;
	wire n_2801;
	wire n_2802;
	wire n_2803;
	wire n_2804;
	wire n_2805;
	wire n_2806;
	wire n_2807;
	wire n_2808;
	wire n_2809;
	wire n_2810;
	wire n_2811;
	wire n_2812;
	wire n_2813;
	wire n_2814;
	wire n_2815;
	wire n_2816;
	wire n_2817;
	wire n_2818;
	wire n_2819;
	wire n_2820;
	wire n_2821;
	wire n_2822;
	wire n_2823;
	wire n_2824;
	wire n_2825;
	wire n_2826;
	wire n_2827;
	wire n_2828;
	wire n_2829;
	wire n_2830;
	wire n_2831;
	wire n_2832;
	wire n_2833;
	wire n_2834;
	wire n_2835;
	wire n_2836;
	wire n_2837;
	wire n_2838;
	wire n_2839;
	wire n_2840;
	wire n_2841;
	wire n_2842;
	wire n_2843;
	wire n_2844;
	wire n_2845;
	wire n_2846;
	wire n_2847;
	wire n_2848;
	wire n_2849;
	wire n_2850;
	wire n_2851;
	wire n_2852;
	wire n_2853;
	wire n_2854;
	wire n_2855;
	wire n_2856;
	wire n_2857;
	wire n_2858;
	wire n_2859;
	wire n_2860;
	wire n_2861;
	wire n_2862;
	wire n_2863;
	wire n_2864;
	wire n_2865;
	wire n_2866;
	wire n_2867;
	wire n_2868;
	wire n_2869;
	wire n_2870;
	wire n_2871;
	wire n_2872;
	wire n_2873;
	wire n_2874;
	wire n_2875;
	wire n_2876;
	wire n_2877;
	wire n_2878;
	wire n_2879;
	wire n_2880;
	wire n_2881;
	wire n_2882;
	wire n_2883;
	wire n_2884;
	wire n_2885;
	wire n_2886;
	wire n_2887;
	wire n_2888;
	wire n_2889;
	wire n_2890;
	wire n_2891;
	wire n_2892;
	wire n_2893;
	wire n_2894;
	wire n_2895;
	wire n_2896;
	wire n_2897;
	wire n_2898;
	wire n_2899;
	wire n_2900;
	wire n_2901;
	wire n_2902;
	wire n_2903;
	wire n_2904;
	wire n_2905;
	wire n_2906;
	wire n_2907;
	wire n_2908;
	wire n_2909;
	wire n_2910;
	wire n_2911;
	wire n_2912;
	wire n_2913;
	wire n_2914;
	wire n_2915;
	wire n_2916;
	wire n_2917;
	wire n_2918;
	wire n_2919;
	wire n_2920;
	wire n_2921;
	wire n_2922;
	wire n_2923;
	wire n_2924;
	wire n_2925;
	wire n_2926;
	wire n_2927;
	wire n_2928;
	wire n_2929;
	wire n_2930;
	wire n_2931;
	wire n_2932;
	wire n_2933;
	wire n_2934;
	wire n_2935;
	wire n_2936;
	wire n_2937;
	wire n_2938;
	wire n_2939;
	wire n_2940;
	wire n_2941;
	wire n_2942;
	wire n_2943;
	wire n_2944;
	wire n_2945;
	wire n_2946;
	wire n_2947;
	wire n_2948;
	wire n_2949;
	wire n_2950;
	wire n_2951;
	wire n_2952;
	wire n_2953;
	wire n_2954;
	wire n_2955;
	wire n_2956;
	wire n_2957;
	wire n_2958;
	wire n_2959;
	wire n_2960;
	wire n_2961;
	wire n_2962;
	wire n_2963;
	wire n_2964;
	wire n_2965;
	wire n_2966;
	wire n_2967;
	wire n_2968;
	wire n_2969;
	wire n_2970;
	wire n_2971;
	wire n_2972;
	wire n_2973;
	wire n_2974;
	wire n_2975;
	wire n_2976;
	wire n_2977;
	wire n_2978;
	wire n_2979;
	wire n_2980;
	wire n_2981;
	wire n_2982;
	wire n_2983;
	wire n_2984;
	wire n_2985;
	wire n_2986;
	wire n_2987;
	wire n_2988;
	wire n_2989;
	wire n_2990;
	wire n_2991;
	wire n_2992;
	wire n_2993;
	wire n_2994;
	wire n_2995;
	wire n_2996;
	wire n_2997;
	wire n_2998;
	wire n_2999;
	wire n_3000;
	wire n_3001;
	wire n_3002;
	wire n_3003;
	wire n_3004;
	wire n_3005;
	wire n_3006;
	wire n_3007;
	wire n_3008;
	wire n_3009;
	wire n_3010;
	wire n_3011;
	wire n_3012;
	wire n_3013;
	wire n_3014;
	wire n_3015;
	wire n_3016;
	wire n_3017;
	wire n_3018;
	wire n_3019;
	wire n_3020;
	wire n_3021;
	wire n_3022;
	wire n_3023;
	wire n_3024;
	wire n_3025;
	wire n_3026;
	wire n_3027;
	wire n_3028;
	wire n_3029;
	wire n_3030;
	wire n_3031;
	wire n_3032;
	wire n_3033;
	wire n_3034;
	wire n_3035;
	wire n_3036;
	wire n_3037;
	wire n_3038;
	wire n_3039;
	wire n_3040;
	wire n_3041;
	wire n_3042;
	wire n_3043;
	wire n_3044;
	wire n_3045;
	wire n_3046;
	wire n_3047;
	wire n_3048;
	wire n_3049;
	wire n_3050;
	wire n_3051;
	wire n_3052;
	wire n_3053;
	wire n_3054;
	wire n_3055;
	wire n_3056;
	wire n_3057;
	wire n_3058;
	wire n_3059;
	wire n_3060;
	wire n_3061;
	wire n_3062;
	wire n_3063;
	wire n_3064;
	wire n_3065;
	wire n_3066;
	wire n_3067;
	wire n_3068;
	wire n_3069;
	wire n_3070;
	wire n_3071;
	wire n_3072;
	wire n_3073;
	wire n_3074;
	wire n_3075;
	wire n_3076;
	wire n_3077;
	wire n_3078;
	wire n_3079;
	wire n_3080;
	wire n_3081;
	wire n_3082;
	wire n_3083;
	wire n_3084;
	wire n_3085;
	wire n_3086;
	wire n_3087;
	wire n_3088;
	wire n_3089;
	wire n_3090;
	wire n_3091;
	wire n_3092;
	wire n_3093;
	wire n_3094;
	wire n_3095;
	wire n_3096;
	wire n_3097;
	wire n_3098;
	wire n_3099;
	wire n_3100;
	wire n_3101;
	wire n_3102;
	wire n_3103;
	wire n_3104;
	wire n_3105;
	wire n_3106;
	wire n_3107;
	wire n_3108;
	wire n_3109;
	wire n_3110;
	wire n_3111;
	wire n_3112;
	wire n_3113;
	wire n_3114;
	wire n_3115;
	wire n_3116;
	wire n_3117;
	wire n_3118;
	wire n_3119;
	wire n_3120;
	wire n_3121;
	wire n_3122;
	wire n_3123;
	wire n_3124;
	wire n_3125;
	wire n_3126;
	wire n_3127;
	wire n_3128;
	wire n_3129;
	wire n_3130;
	wire n_3131;
	wire n_3132;
	wire n_3133;
	wire n_3134;
	wire n_3135;
	wire n_3136;
	wire n_3137;
	wire n_3138;
	wire n_3139;
	wire n_3140;
	wire n_3141;
	wire n_3142;
	wire n_3143;
	wire n_3144;
	wire n_3145;
	wire n_3146;
	wire n_3147;
	wire n_3148;
	wire n_3149;
	wire n_3150;
	wire n_3151;
	wire n_3152;
	wire n_3153;
	wire n_3154;
	wire n_3155;
	wire n_3156;
	wire n_3157;
	wire n_3158;
	wire n_3159;
	wire n_3160;
	wire n_3161;
	wire n_3162;
	wire n_3163;
	wire n_3164;
	wire n_3165;
	wire n_3166;
	wire n_3167;
	wire n_3168;
	wire n_3169;
	wire n_3170;
	wire n_3171;
	wire n_3172;
	wire n_3173;
	wire n_3174;
	wire n_3175;
	wire n_3176;
	wire n_3177;
	wire n_3178;
	wire n_3179;
	wire n_3180;
	wire n_3181;
	wire n_3182;
	wire n_3183;
	wire n_3184;
	wire n_3185;
	wire n_3186;
	wire n_3187;
	wire n_3188;
	wire n_3189;
	wire n_3190;
	wire n_3191;
	wire n_3192;
	wire n_3193;
	wire n_3194;
	wire n_3195;
	wire n_3196;
	wire n_3197;
	wire n_3198;
	wire n_3199;
	wire n_3200;
	wire n_3201;
	wire n_3202;
	wire n_3203;
	wire n_3204;
	wire n_3205;
	wire n_3206;
	wire n_3207;
	wire n_3208;
	wire n_3209;
	wire n_3210;
	wire n_3211;
	wire n_3212;
	wire n_3213;
	wire n_3214;
	wire n_3215;
	wire n_3216;
	wire n_3217;
	wire n_3218;
	wire n_3219;
	wire n_3220;
	wire n_3221;
	wire n_3222;
	wire n_3223;
	wire n_3224;
	wire n_3225;
	wire n_3226;
	wire n_3227;
	wire n_3228;
	wire n_3229;
	wire n_3230;
	wire n_3231;
	wire n_3232;
	wire n_3233;
	wire n_3234;
	wire n_3235;
	wire n_3236;
	wire n_3237;
	wire n_3238;
	wire n_3239;
	wire n_3240;
	wire n_3241;
	wire n_3242;
	wire n_3243;
	wire n_3244;
	wire n_3245;
	wire n_3246;
	wire n_3247;
	wire n_3248;
	wire n_3249;
	wire n_3250;
	wire n_3251;
	wire n_3252;
	wire n_3253;
	wire n_3254;
	wire n_3255;
	wire n_3256;
	wire n_3257;
	wire n_3258;
	wire n_3259;
	wire n_3260;
	wire n_3261;
	wire n_3262;
	wire n_3263;
	wire n_3264;
	wire n_3265;
	wire n_3266;
	wire n_3267;
	wire n_3268;
	wire n_3269;
	wire n_3270;
	wire n_3271;
	wire n_3272;
	wire n_3273;
	wire n_3274;
	wire n_3275;
	wire n_3276;
	wire n_3277;
	wire n_3278;
	wire n_3279;
	wire n_3280;
	wire n_3281;
	wire n_3282;
	wire n_3283;
	wire n_3284;
	wire n_3285;
	wire n_3286;
	wire n_3287;
	wire n_3288;
	wire n_3289;
	wire n_3290;
	wire n_3291;
	wire n_3292;
	wire n_3293;
	wire n_3294;
	wire n_3295;
	wire n_3296;
	wire n_3297;
	wire n_3298;
	wire n_3299;
	wire n_3300;
	wire n_3301;
	wire n_3302;
	wire n_3303;
	wire n_3304;
	wire n_3305;
	wire n_3306;
	wire n_3307;
	wire n_3308;
	wire n_3309;
	wire n_3310;
	wire n_3311;
	wire n_3312;
	wire n_3313;
	wire n_3314;
	wire n_3315;
	wire n_3316;
	wire n_3317;
	wire n_3318;
	wire n_3319;
	wire n_3320;
	wire n_3321;
	wire n_3322;
	wire n_3323;
	wire n_3324;
	wire n_3325;
	wire n_3326;
	wire n_3327;
	wire n_3328;
	wire n_3329;
	wire n_3330;
	wire n_3331;
	wire n_3332;
	wire n_3333;
	wire n_3334;
	wire n_3335;
	wire n_3336;
	wire n_3337;
	wire n_3338;
	wire n_3339;
	wire n_3340;
	wire n_3341;
	wire n_3342;
	wire n_3343;
	wire n_3344;
	wire n_3345;
	wire n_3346;
	wire n_3347;
	wire n_3348;
	wire n_3349;
	wire n_3350;
	wire n_3351;
	wire n_3352;
	wire n_3353;
	wire n_3354;
	wire n_3355;
	wire n_3356;
	wire n_3357;
	wire n_3358;
	wire n_3359;
	wire n_3360;
	wire n_3361;
	wire n_3362;
	wire n_3363;
	wire n_3364;
	wire n_3365;
	wire n_3366;
	wire n_3367;
	wire n_3368;
	wire n_3369;
	wire n_3370;
	wire n_3371;
	wire n_3372;
	wire n_3373;
	wire n_3374;
	wire n_3375;
	wire n_3376;
	wire n_3377;
	wire n_3378;
	wire n_3379;
	wire n_3380;
	wire n_3381;
	wire n_3382;
	wire n_3383;
	wire n_3384;
	wire n_3385;
	wire n_3386;
	wire n_3387;
	wire n_3388;
	wire n_3389;
	wire n_3390;
	wire n_3391;
	wire n_3392;
	wire n_3393;
	wire n_3394;
	wire n_3395;
	wire n_3396;
	wire n_3397;
	wire n_3398;
	wire n_3399;
	wire n_3400;
	wire n_3401;
	wire n_3402;
	wire n_3403;
	wire n_3404;
	wire n_3405;
	wire n_3406;
	wire n_3407;
	wire n_3408;
	wire n_3409;
	wire n_3410;
	wire n_3411;
	wire n_3412;
	wire n_3413;
	wire n_3414;
	wire n_3415;
	wire n_3416;
	wire n_3417;
	wire n_3418;
	wire n_3419;
	wire n_3420;
	wire n_3421;
	wire n_3422;
	wire n_3423;
	wire n_3424;
	wire n_3425;
	wire n_3426;
	wire n_3427;
	wire n_3428;
	wire n_3429;
	wire n_3430;
	wire n_3431;
	wire n_3432;
	wire n_3433;
	wire n_3434;
	wire n_3435;
	wire n_3436;
	wire n_3437;
	wire n_3438;
	wire n_3439;
	wire n_3440;
	wire n_3441;
	wire n_3442;
	wire n_3443;
	wire n_3444;
	wire n_3445;
	wire n_3446;
	wire n_3447;
	wire n_3448;
	wire n_3449;
	wire n_3450;
	wire n_3451;
	wire n_3452;
	wire n_3453;
	wire n_3454;
	wire n_3455;
	wire n_3456;
	wire n_3457;
	wire n_3458;
	wire n_3459;
	wire n_3460;
	wire n_3461;
	wire n_3462;
	wire n_3463;
	wire n_3464;
	wire n_3465;
	wire n_3466;
	wire n_3467;
	wire n_3468;
	wire n_3469;
	wire n_3470;
	wire n_3471;
	wire n_3472;
	wire n_3473;
	wire n_3474;
	wire n_3475;
	wire n_3476;
	wire n_3477;
	wire n_3478;
	wire n_3479;
	wire n_3480;
	wire n_3481;
	wire n_3482;
	wire n_3483;
	wire n_3484;
	wire n_3485;
	wire n_3486;
	wire n_3487;
	wire n_3488;
	wire n_3489;
	wire n_3490;
	wire n_3491;
	wire n_3492;
	wire n_3493;
	wire n_3494;
	wire n_3495;
	wire n_3496;
	wire n_3497;
	wire n_3498;
	wire n_3499;
	wire n_3500;
	wire n_3501;
	wire n_3502;
	wire n_3503;
	wire n_3504;
	wire n_3505;
	wire n_3506;
	wire n_3507;
	wire n_3508;
	wire n_3509;
	wire n_3510;
	wire n_3511;
	wire n_3512;
	wire n_3513;
	wire n_3514;
	wire n_3515;
	wire n_3516;
	wire n_3517;
	wire n_3518;
	wire n_3519;
	wire n_3520;
	wire n_3521;
	wire n_3522;
	wire n_3523;
	wire n_3524;
	wire n_3525;
	wire n_3526;
	wire n_3527;
	wire n_3528;
	wire n_3529;
	wire n_3530;
	wire n_3531;
	wire n_3532;
	wire n_3533;
	wire n_3534;
	wire n_3535;
	wire n_3536;
	wire n_3537;
	wire n_3538;
	wire n_3539;
	wire n_3540;
	wire n_3541;
	wire n_3542;
	wire n_3543;
	wire n_3544;
	wire n_3545;
	wire n_3546;
	wire n_3547;
	wire n_3548;
	wire n_3549;
	wire n_3550;
	wire n_3551;
	wire n_3552;
	wire n_3553;
	wire n_3554;
	wire n_3555;
	wire n_3556;
	wire n_3557;
	wire n_3558;
	wire n_3559;
	wire n_3560;
	wire n_3561;
	wire n_3562;
	wire n_3563;
	wire n_3564;
	wire n_3565;
	wire n_3566;
	wire n_3567;
	wire n_3568;
	wire n_3569;
	wire n_3570;
	wire n_3571;
	wire n_3572;
	wire n_3573;
	wire n_3574;
	wire n_3575;
	wire n_3576;
	wire n_3577;
	wire n_3578;
	wire n_3579;
	wire n_3580;
	wire n_3581;
	wire n_3582;
	wire n_3583;
	wire n_3584;
	wire n_3585;
	wire n_3586;
	wire n_3587;
	wire n_3588;
	wire n_3589;
	wire n_3590;
	wire n_3591;
	wire n_3592;
	wire n_3593;
	wire n_3594;
	wire n_3595;
	wire n_3596;
	wire n_3597;
	wire n_3598;
	wire n_3599;
	wire n_3600;
	wire n_3601;
	wire n_3602;
	wire n_3603;
	wire n_3604;
	wire n_3605;
	wire n_3606;
	wire n_3607;
	wire n_3608;
	wire n_3609;
	wire n_3610;
	wire n_3611;
	wire n_3612;
	wire n_3613;
	wire n_3614;
	wire n_3615;
	wire n_3616;
	wire n_3617;
	wire n_3618;
	wire n_3619;
	wire n_3620;
	wire n_3621;
	wire n_3622;
	wire n_3623;
	wire n_3624;
	wire n_3625;
	wire n_3626;
	wire n_3627;
	wire n_3628;
	wire n_3629;
	wire n_3630;
	wire n_3631;
	wire n_3632;
	wire n_3633;
	wire n_3634;
	wire n_3635;
	wire n_3636;
	wire n_3637;
	wire n_3638;
	wire n_3639;
	wire n_3640;
	wire n_3641;
	wire n_3642;
	wire n_3643;
	wire n_3644;
	wire n_3645;
	wire n_3646;
	wire n_3647;
	wire n_3648;
	wire n_3649;
	wire n_3650;
	wire n_3651;
	wire n_3652;
	wire n_3653;
	wire n_3654;
	wire n_3655;
	wire n_3656;
	wire n_3657;
	wire n_3658;
	wire n_3659;
	wire n_3660;
	wire n_3661;
	wire n_3662;
	wire n_3663;
	wire n_3664;
	wire n_3665;
	wire n_3666;
	wire n_3667;
	wire n_3668;
	wire n_3669;
	wire n_3670;
	wire n_3671;
	wire n_3672;
	wire n_3673;
	wire n_3674;
	wire n_3675;
	wire n_3676;
	wire n_3677;
	wire n_3678;
	wire n_3679;
	wire n_3680;
	wire n_3681;
	wire n_3682;
	wire n_3683;
	wire n_3684;
	wire n_3685;
	wire n_3686;
	wire n_3687;
	wire n_3688;
	wire n_3689;
	wire n_3690;
	wire n_3691;
	wire n_3692;
	wire n_3693;
	wire n_3694;
	wire n_3695;
	wire n_3696;
	wire n_3697;
	wire n_3698;
	wire n_3699;
	wire n_3700;
	wire n_3701;
	wire n_3702;
	wire n_3703;
	wire n_3704;
	wire n_3705;
	wire n_3706;
	wire n_3707;
	wire n_3708;
	wire n_3709;
	wire n_3710;
	wire n_3711;
	wire n_3712;
	wire n_3713;
	wire n_3714;
	wire n_3715;
	wire n_3716;
	wire n_3717;
	wire n_3718;
	wire n_3719;
	wire n_3720;
	wire n_3721;
	wire n_3722;
	wire n_3723;
	wire n_3724;
	wire n_3725;
	wire n_3726;
	wire n_3727;
	wire n_3728;
	wire n_3729;
	wire n_3730;
	wire n_3731;
	wire n_3732;
	wire n_3733;
	wire n_3734;
	wire n_3735;
	wire n_3736;
	wire n_3737;
	wire n_3738;
	wire n_3739;
	wire n_3740;
	wire n_3741;
	wire n_3742;
	wire n_3743;
	wire n_3744;
	wire n_3745;
	wire n_3746;
	wire n_3747;
	wire n_3748;
	wire n_3749;
	wire n_3750;
	wire n_3751;
	wire n_3752;
	wire n_3753;
	wire n_3754;
	wire n_3755;
	wire n_3756;
	wire n_3757;
	wire n_3758;
	wire n_3759;
	wire n_3760;
	wire n_3761;
	wire n_3762;
	wire n_3763;
	wire n_3764;
	wire n_3765;
	wire n_3766;
	wire n_3767;
	wire n_3768;
	wire n_3769;
	wire n_3770;
	wire n_3771;
	wire n_3772;
	wire n_3773;
	wire n_3774;
	wire n_3775;
	wire n_3776;
	wire n_3777;
	wire n_3778;
	wire n_3779;
	wire n_3780;
	wire n_3781;
	wire n_3782;
	wire n_3783;
	wire n_3784;
	wire n_3785;
	wire n_3786;
	wire n_3787;
	wire n_3788;
	wire n_3789;
	wire n_3790;
	wire n_3791;
	wire n_3792;
	wire n_3793;
	wire n_3794;
	wire n_3795;
	wire n_3796;
	wire n_3797;
	wire n_3798;
	wire n_3799;
	wire n_3800;
	wire n_3801;
	wire n_3802;
	wire n_3803;
	wire n_3804;
	wire n_3805;
	wire n_3806;
	wire n_3807;
	wire n_3808;
	wire n_3809;
	wire n_3810;
	wire n_3811;
	wire n_3812;
	wire n_3813;
	wire n_3814;
	wire n_3815;
	wire n_3816;
	wire n_3817;
	wire n_3818;
	wire n_3819;
	wire n_3820;
	wire n_3821;
	wire n_3822;
	wire n_3823;
	wire n_3824;
	wire n_3825;
	wire n_3826;
	wire n_3827;
	wire n_3828;
	wire n_3829;
	wire n_3830;
	wire n_3831;
	wire n_3832;
	wire n_3833;
	wire n_3834;
	wire n_3835;
	wire n_3836;
	wire n_3837;
	wire n_3838;
	wire n_3839;
	wire n_3840;
	wire n_3841;
	wire n_3842;
	wire n_3843;
	wire n_3844;
	wire n_3845;
	wire n_3846;
	wire n_3847;
	wire n_3848;
	wire n_3849;
	wire n_3850;
	wire n_3851;
	wire n_3852;
	wire n_3853;
	wire n_3854;
	wire n_3855;
	wire n_3856;
	wire n_3857;
	wire n_3858;
	wire n_3859;
	wire n_3860;
	wire n_3861;
	wire n_3862;
	wire n_3863;
	wire n_3864;
	wire n_3865;
	wire n_3866;
	wire n_3867;
	wire n_3868;
	wire n_3869;
	wire n_3870;
	wire n_3871;
	wire n_3872;
	wire n_3873;
	wire n_3874;
	wire n_3875;
	wire n_3876;
	wire n_3877;
	wire n_3878;
	wire n_3879;
	wire n_3880;
	wire n_3881;
	wire n_3882;
	wire n_3883;
	wire n_3884;
	wire n_3885;
	wire n_3886;
	wire n_3887;
	wire n_3888;
	wire n_3889;
	wire n_3890;
	wire n_3891;
	wire n_3892;
	wire n_3893;
	wire n_3894;
	wire n_3895;
	wire n_3896;
	wire n_3897;
	wire n_3898;
	wire n_3899;
	wire n_3900;
	wire n_3901;
	wire n_3902;
	wire n_3903;
	wire n_3904;
	wire n_3905;
	wire n_3906;
	wire n_3907;
	wire n_3908;
	wire n_3909;
	wire n_3910;
	wire n_3911;
	wire n_3912;
	wire n_3913;
	wire n_3914;
	wire n_3915;
	wire n_3916;
	wire n_3917;
	wire n_3918;
	wire n_3919;
	wire n_3920;
	wire n_3921;
	wire n_3922;
	wire n_3923;
	wire n_3924;
	wire n_3925;
	wire n_3926;
	wire n_3927;
	wire n_3928;
	wire n_3929;
	wire n_3930;
	wire n_3931;
	wire n_3932;
	wire n_3933;
	wire n_3934;
	wire n_3935;
	wire n_3936;
	wire n_3937;
	wire n_3938;
	wire n_3939;
	wire n_3940;
	wire n_3941;
	wire n_3942;
	wire n_3943;
	wire n_3944;
	wire n_3945;
	wire n_3946;
	wire n_3947;
	wire n_3948;
	wire n_3949;
	wire n_3950;
	wire n_3951;
	wire n_3952;
	wire n_3953;
	wire n_3954;
	wire n_3955;
	wire n_3956;
	wire n_3957;
	wire n_3958;
	wire n_3959;
	wire n_3960;
	wire n_3961;
	wire n_3962;
	wire n_3963;
	wire n_3964;
	wire n_3965;
	wire n_3966;
	wire n_3967;
	wire n_3968;
	wire n_3969;
	wire n_3970;
	wire n_3971;
	wire n_3972;
	wire n_3973;
	wire n_3974;
	wire n_3975;
	wire n_3976;
	wire n_3977;
	wire n_3978;
	wire n_3979;
	wire n_3980;
	wire n_3981;
	wire n_3982;
	wire n_3983;
	wire n_3984;
	wire n_3985;
	wire n_3986;
	wire n_3987;
	wire n_3988;
	wire n_3989;
	wire n_3990;
	wire n_3991;
	wire n_3992;
	wire n_3993;
	wire n_3994;
	wire n_3995;
	wire n_3996;
	wire n_3997;
	wire n_3998;
	wire n_3999;
	wire n_4000;
	wire n_4001;
	wire n_4002;
	wire n_4003;
	wire n_4004;
	wire n_4005;
	wire n_4006;
	wire n_4007;
	wire n_4008;
	wire n_4009;
	wire n_4010;
	wire n_4011;
	wire n_4012;
	wire n_4013;
	wire n_4014;
	wire n_4015;
	wire n_4016;
	wire n_4017;
	wire n_4018;
	wire n_4019;
	wire n_4020;
	wire n_4021;
	wire n_4022;
	wire n_4023;
	wire n_4024;
	wire n_4025;
	wire n_4026;
	wire n_4027;
	wire n_4028;
	wire n_4029;
	wire n_4030;
	wire n_4031;
	wire n_4032;
	wire n_4033;
	wire n_4034;
	wire n_4035;
	wire n_4036;
	wire n_4037;
	wire n_4038;
	wire n_4039;
	wire n_4040;
	wire n_4041;
	wire n_4042;
	wire n_4043;
	wire n_4044;
	wire n_4045;
	wire n_4046;
	wire n_4047;
	wire n_4048;
	wire n_4049;
	wire n_4050;
	wire n_4051;
	wire n_4052;
	wire n_4053;
	wire n_4054;
	wire n_4055;
	wire n_4056;
	wire n_4057;
	wire n_4058;
	wire n_4059;
	wire n_4060;
	wire n_4061;
	wire n_4062;
	wire n_4063;
	wire n_4064;
	wire n_4065;
	wire n_4066;
	wire n_4067;
	wire n_4068;
	wire n_4069;
	wire n_4070;
	wire n_4071;
	wire n_4072;
	wire n_4073;
	wire n_4074;
	wire n_4075;
	wire n_4076;
	wire n_4077;
	wire n_4078;
	wire n_4079;
	wire n_4080;
	wire n_4081;
	wire n_4082;
	wire n_4083;
	wire n_4084;
	wire n_4085;
	wire n_4086;
	wire n_4087;
	wire n_4088;
	wire n_4089;
	wire n_4090;
	wire n_4091;
	wire n_4092;
	wire n_4093;
	wire n_4094;
	wire n_4095;
	wire n_4096;
	wire n_4097;
	wire n_4098;
	wire n_4099;
	wire n_4100;
	wire n_4101;
	wire n_4102;
	wire n_4103;
	wire n_4104;
	wire n_4105;
	wire n_4106;
	wire n_4107;
	wire n_4108;
	wire n_4109;
	wire n_4110;
	wire n_4111;
	wire n_4112;
	wire n_4113;
	wire n_4114;
	wire n_4115;
	wire n_4116;
	wire n_4117;
	wire n_4118;
	wire n_4119;
	wire n_4120;
	wire n_4121;
	wire n_4122;
	wire n_4123;
	wire n_4124;
	wire n_4125;
	wire n_4126;
	wire n_4127;
	wire n_4128;
	wire n_4129;
	wire n_4130;
	wire n_4131;
	wire n_4132;
	wire n_4133;
	wire n_4134;
	wire n_4135;
	wire n_4136;
	wire n_4137;
	wire n_4138;
	wire n_4139;
	wire n_4140;
	wire n_4141;
	wire n_4142;
	wire n_4143;
	wire n_4144;
	wire n_4145;
	wire n_4146;
	wire n_4147;
	wire n_4148;
	wire n_4149;
	wire n_4150;
	wire n_4151;
	wire n_4152;
	wire n_4153;
	wire n_4154;
	wire n_4155;
	wire n_4156;
	wire n_4157;
	wire n_4158;
	wire n_4159;
	wire n_4160;
	wire n_4161;
	wire n_4162;
	wire n_4163;
	wire n_4164;
	wire n_4165;
	wire n_4166;
	wire n_4167;
	wire n_4168;
	wire n_4169;
	wire n_4170;
	wire n_4171;
	wire n_4172;
	wire n_4173;
	wire n_4174;
	wire n_4175;
	wire n_4176;
	wire n_4177;
	wire n_4178;
	wire n_4179;
	wire n_4180;
	wire n_4181;
	wire n_4182;
	wire n_4183;
	wire n_4184;
	wire n_4185;
	wire n_4186;
	wire n_4187;
	wire n_4188;
	wire n_4189;
	wire n_4190;
	wire n_4191;
	wire n_4192;
	wire n_4193;
	wire n_4194;
	wire n_4195;
	wire n_4196;
	wire n_4197;
	wire n_4198;
	wire n_4199;
	wire n_4200;
	wire n_4201;
	wire n_4202;
	wire n_4203;
	wire n_4204;
	wire n_4205;
	wire n_4206;
	wire n_4207;
	wire n_4208;
	wire n_4209;
	wire n_4210;
	wire n_4211;
	wire n_4212;
	wire n_4213;
	wire n_4214;
	wire n_4215;
	wire n_4216;
	wire n_4217;
	wire n_4218;
	wire n_4219;
	wire n_4220;
	wire n_4221;
	wire n_4222;
	wire n_4223;
	wire n_4224;
	wire n_4225;
	wire n_4226;
	wire n_4227;
	wire n_4228;
	wire n_4229;
	wire n_4230;
	wire n_4231;
	wire n_4232;
	wire n_4233;
	wire n_4234;
	wire n_4235;
	wire n_4236;
	wire n_4237;
	wire n_4238;
	wire n_4239;
	wire n_4240;
	wire n_4241;
	wire n_4242;
	wire n_4243;
	wire n_4244;
	wire n_4245;
	wire n_4246;
	wire n_4247;
	wire n_4248;
	wire n_4249;
	wire n_4250;
	wire n_4251;
	wire n_4252;
	wire n_4253;
	wire n_4254;
	wire n_4255;
	wire n_4256;
	wire n_4257;
	wire n_4258;
	wire n_4259;
	wire n_4260;
	wire n_4261;
	wire n_4262;
	wire n_4263;
	wire n_4264;
	wire n_4265;
	wire n_4266;
	wire n_4267;
	wire n_4268;
	wire n_4269;
	wire n_4270;
	wire n_4271;
	wire n_4272;
	wire n_4273;
	wire n_4274;
	wire n_4275;
	wire n_4276;
	wire n_4277;
	wire n_4278;
	wire n_4279;
	wire n_4280;
	wire n_4281;
	wire n_4282;
	wire n_4283;
	wire n_4284;
	wire n_4285;
	wire n_4286;
	wire n_4287;
	wire n_4288;
	wire n_4289;
	wire n_4290;
	wire n_4291;
	wire n_4292;
	wire n_4293;
	wire n_4294;
	wire n_4295;
	wire n_4296;
	wire n_4297;
	wire n_4298;
	wire n_4299;
	wire n_4300;
	wire n_4301;
	wire n_4302;
	wire n_4303;
	wire n_4304;
	wire n_4305;
	wire n_4306;
	wire n_4307;
	wire n_4308;
	wire n_4309;
	wire n_4310;
	wire n_4311;
	wire n_4312;
	wire n_4313;
	wire n_4314;
	wire n_4315;
	wire n_4316;
	wire n_4317;
	wire n_4318;
	wire n_4319;
	wire n_4320;
	wire n_4321;
	wire n_4322;
	wire n_4323;
	wire n_4324;
	wire n_4325;
	wire n_4326;
	wire n_4327;
	wire n_4328;
	wire n_4329;
	wire n_4330;
	wire n_4331;
	wire n_4332;
	wire n_4333;
	wire n_4334;
	wire n_4335;
	wire n_4336;
	wire n_4337;
	wire n_4338;
	wire n_4339;
	wire n_4340;
	wire n_4341;
	wire n_4342;
	wire n_4343;
	wire n_4344;
	wire n_4345;
	wire n_4346;
	wire n_4347;
	wire n_4348;
	wire n_4349;
	wire n_4350;
	wire n_4351;
	wire n_4352;
	wire n_4353;
	wire n_4354;
	wire n_4355;
	wire n_4356;
	wire n_4357;
	wire n_4358;
	wire n_4359;
	wire n_4360;
	wire n_4361;
	wire n_4362;
	wire n_4363;
	wire n_4364;
	wire n_4365;
	wire n_4366;
	wire n_4367;
	wire n_4368;
	wire n_4369;
	wire n_4370;
	wire n_4371;
	wire n_4372;
	wire n_4373;
	wire n_4374;
	wire n_4375;
	wire n_4376;
	wire n_4377;
	wire n_4378;
	wire n_4379;
	wire n_4380;
	wire n_4381;
	wire n_4382;
	wire n_4383;
	wire n_4384;
	wire n_4385;
	wire n_4386;
	wire n_4387;
	wire n_4388;
	wire n_4389;
	wire n_4390;
	wire n_4391;
	wire n_4392;
	wire n_4393;
	wire n_4394;
	wire n_4395;
	wire n_4396;
	wire n_4397;
	wire n_4398;
	wire n_4399;
	wire n_4400;
	wire n_4401;
	wire n_4402;
	wire n_4403;
	wire n_4404;
	wire n_4405;
	wire n_4406;
	wire n_4407;
	wire n_4408;
	wire n_4409;
	wire n_4410;
	wire n_4411;
	wire n_4412;
	wire n_4413;
	wire n_4414;
	wire n_4415;
	wire n_4416;
	wire n_4417;
	wire n_4418;
	wire n_4419;
	wire n_4420;
	wire n_4421;
	wire n_4422;
	wire n_4423;
	wire n_4424;
	wire n_4425;
	wire n_4426;
	wire n_4427;
	wire n_4428;
	wire n_4429;
	wire n_4430;
	wire n_4431;
	wire n_4432;
	wire n_4433;
	wire n_4434;
	wire n_4435;
	wire n_4436;
	wire n_4437;
	wire n_4438;
	wire n_4439;
	wire n_4440;
	wire n_4441;
	wire n_4442;
	wire n_4443;
	wire n_4444;
	wire n_4445;
	wire n_4446;
	wire n_4447;
	wire n_4448;
	wire n_4449;
	wire n_4450;
	wire n_4451;
	wire n_4452;
	wire n_4453;
	wire n_4454;
	wire n_4455;
	wire n_4456;
	wire n_4457;
	wire n_4458;
	wire n_4459;
	wire n_4460;
	wire n_4461;
	wire n_4462;
	wire n_4463;
	wire n_4464;
	wire n_4465;
	wire n_4466;
	wire n_4467;
	wire n_4468;
	wire n_4469;
	wire n_4470;
	wire n_4471;
	wire n_4472;
	wire n_4473;
	wire n_4474;
	wire n_4475;
	wire n_4476;
	wire n_4477;
	wire n_4478;
	wire n_4479;
	wire n_4480;
	wire n_4481;
	wire n_4482;
	wire n_4483;
	wire n_4484;
	wire n_4485;
	wire n_4486;
	wire n_4487;
	wire n_4488;
	wire n_4489;
	wire n_4490;
	wire n_4491;
	wire n_4492;
	wire n_4493;
	wire n_4494;
	wire n_4495;
	wire n_4496;
	wire n_4497;
	wire n_4498;
	wire n_4499;
	wire n_4500;
	wire n_4501;
	wire n_4502;
	wire n_4503;
	wire n_4504;
	wire n_4505;
	wire n_4506;
	wire n_4507;
	wire n_4508;
	wire n_4509;
	wire n_4510;
	wire n_4511;
	wire n_4512;
	wire n_4513;
	wire n_4514;
	wire n_4515;
	wire n_4516;
	wire n_4517;
	wire n_4518;
	wire n_4519;
	wire n_4520;
	wire n_4521;
	wire n_4522;
	wire n_4523;
	wire n_4524;
	wire n_4525;
	wire n_4526;
	wire n_4527;
	wire n_4528;
	wire n_4529;
	wire n_4530;
	wire n_4531;
	wire n_4532;
	wire n_4533;
	wire n_4534;
	wire n_4535;
	wire n_4536;
	wire n_4537;
	wire n_4538;
	wire n_4539;
	wire n_4540;
	wire n_4541;
	wire n_4542;
	wire n_4543;
	wire n_4544;
	wire n_4545;
	wire n_4546;
	wire n_4547;
	wire n_4548;
	wire n_4549;
	wire n_4550;
	wire n_4551;
	wire n_4552;
	wire n_4553;
	wire n_4554;
	wire n_4555;
	wire n_4556;
	wire n_4557;
	wire n_4558;
	wire n_4559;
	wire n_4560;
	wire n_4561;
	wire n_4562;
	wire n_4563;
	wire n_4564;
	wire n_4565;
	wire n_4566;
	wire n_4567;
	wire n_4568;
	wire n_4569;
	wire n_4570;
	wire n_4571;
	wire n_4572;
	wire n_4573;
	wire n_4574;
	wire n_4575;
	wire n_4576;
	wire n_4577;
	wire n_4578;
	wire n_4579;
	wire n_4580;
	wire n_4581;
	wire n_4582;
	wire n_4583;
	wire n_4584;
	wire n_4585;
	wire n_4586;
	wire n_4587;
	wire n_4588;
	wire n_4589;
	wire n_4590;
	wire n_4591;
	wire n_4592;
	wire n_4593;
	wire n_4594;
	wire n_4595;
	wire n_4596;
	wire n_4597;
	wire n_4598;
	wire n_4599;
	wire n_4600;
	wire n_4601;
	wire n_4602;
	wire n_4603;
	wire n_4604;
	wire n_4605;
	wire n_4606;
	wire n_4607;
	wire n_4608;
	wire n_4609;
	wire n_4610;
	wire n_4611;
	wire n_4612;
	wire n_4613;
	wire n_4614;
	wire n_4615;
	wire n_4616;
	wire n_4617;
	wire n_4618;
	wire n_4619;
	wire n_4620;
	wire n_4621;
	wire n_4622;
	wire n_4623;
	wire n_4624;
	wire n_4625;
	wire n_4626;
	wire n_4627;
	wire n_4628;
	wire n_4629;
	wire n_4630;
	wire n_4631;
	wire n_4632;
	wire n_4633;
	wire n_4634;
	wire n_4635;
	wire n_4636;
	wire n_4637;
	wire n_4638;
	wire n_4639;
	wire n_4640;
	wire n_4641;
	wire n_4642;
	wire n_4643;
	wire n_4644;
	wire n_4645;
	wire n_4646;
	wire n_4647;
	wire n_4648;
	wire n_4649;
	wire n_4650;
	wire n_4651;
	wire n_4652;
	wire n_4653;
	wire n_4654;
	wire n_4655;
	wire n_4656;
	wire n_4657;
	wire n_4658;
	wire n_4659;
	wire n_4660;
	wire n_4661;
	wire n_4662;
	wire n_4663;
	wire n_4664;
	wire n_4665;
	wire n_4666;
	wire n_4667;
	wire n_4668;
	wire n_4669;
	wire n_4670;
	wire n_4671;
	wire n_4672;
	wire n_4673;
	wire n_4674;
	wire n_4675;
	wire n_4676;
	wire n_4677;
	wire n_4678;
	wire n_4679;
	wire n_4680;
	wire n_4681;
	wire n_4682;
	wire n_4683;
	wire n_4684;
	wire n_4685;
	wire n_4686;
	wire n_4687;
	wire n_4688;
	wire n_4689;
	wire n_4690;
	wire n_4691;
	wire n_4692;
	wire n_4693;
	wire n_4694;
	wire n_4695;
	wire n_4696;
	wire n_4697;
	wire n_4698;
	wire n_4699;
	wire n_4700;
	wire n_4701;
	wire n_4702;
	wire n_4703;
	wire n_4704;
	wire n_4705;
	wire n_4706;
	wire n_4707;
	wire n_4708;
	wire n_4709;
	wire n_4710;
	wire n_4711;
	wire n_4712;
	wire n_4713;
	wire n_4714;
	wire n_4715;
	wire n_4716;
	wire n_4717;
	wire n_4718;
	wire n_4719;
	wire n_4720;
	wire n_4721;
	wire n_4722;
	wire n_4723;
	wire n_4724;
	wire n_4725;
	wire n_4726;
	wire n_4727;
	wire n_4728;
	wire n_4729;
	wire n_4730;
	wire n_4731;
	wire n_4732;
	wire n_4733;
	wire n_4734;
	wire n_4735;
	wire n_4736;
	wire n_4737;
	wire n_4738;
	wire n_4739;
	wire n_4740;
	wire n_4741;
	wire n_4742;
	wire n_4743;
	wire n_4744;
	wire n_4745;
	wire n_4746;
	wire n_4747;
	wire n_4748;
	wire n_4749;
	wire n_4750;
	wire n_4751;
	wire n_4752;
	wire n_4753;
	wire n_4754;
	wire n_4755;
	wire n_4756;
	wire n_4757;
	wire n_4758;
	wire n_4759;
	wire n_4760;
	wire n_4761;
	wire n_4762;
	wire n_4763;
	wire n_4764;
	wire n_4765;
	wire n_4766;
	wire n_4767;
	wire n_4768;
	wire n_4769;
	wire n_4770;
	wire n_4771;
	wire n_4772;
	wire n_4773;
	wire n_4774;
	wire n_4775;
	wire n_4776;
	wire n_4777;
	wire n_4778;
	wire n_4779;
	wire n_4780;
	wire n_4781;
	wire n_4782;
	wire n_4783;
	wire n_4784;
	wire n_4785;
	wire n_4786;
	wire n_4787;
	wire n_4788;
	wire n_4789;
	wire n_4790;
	wire n_4791;
	wire n_4792;
	wire n_4793;
	wire n_4794;
	wire n_4795;
	wire n_4796;
	wire n_4797;
	wire n_4798;
	wire n_4799;
	wire n_4800;
	wire n_4801;
	wire n_4802;
	wire n_4803;
	wire n_4804;
	wire n_4805;
	wire n_4806;
	wire n_4807;
	wire n_4808;
	wire n_4809;
	wire n_4810;
	wire n_4811;
	wire n_4812;
	wire n_4813;
	wire n_4814;
	wire n_4815;
	wire n_4816;
	wire n_4817;
	wire n_4818;
	wire n_4819;
	wire n_4820;
	wire n_4821;
	wire n_4822;
	wire n_4823;
	wire n_4824;
	wire n_4825;
	wire n_4826;
	wire n_4827;
	wire n_4828;
	wire n_4829;
	wire n_4830;
	wire n_4831;
	wire n_4832;
	wire n_4833;
	wire n_4834;
	wire n_4835;
	wire n_4836;
	wire n_4837;
	wire n_4838;
	wire n_4839;
	wire n_4840;
	wire n_4841;
	wire n_4842;
	wire n_4843;
	wire n_4844;
	wire n_4845;
	wire n_4846;
	wire n_4847;
	wire n_4848;
	wire n_4849;
	wire n_4850;
	wire n_4851;
	wire n_4852;
	wire n_4853;
	wire n_4854;
	wire n_4855;
	wire n_4856;
	wire n_4857;
	wire n_4858;
	wire n_4859;
	wire n_4860;
	wire n_4861;
	wire n_4862;
	wire n_4863;
	wire n_4864;
	wire n_4865;
	wire n_4866;
	wire n_4867;
	wire n_4868;
	wire n_4869;
	wire n_4870;
	wire n_4871;
	wire n_4872;
	wire n_4873;
	wire n_4874;
	wire n_4875;
	wire n_4876;
	wire n_4877;
	wire n_4878;
	wire n_4879;
	wire n_4880;
	wire n_4881;
	wire n_4882;
	wire n_4883;
	wire n_4884;
	wire n_4885;
	wire n_4886;
	wire n_4887;
	wire n_4888;
	wire n_4889;
	wire n_4890;
	wire n_4891;
	wire n_4892;
	wire n_4893;
	wire n_4894;
	wire n_4895;
	wire n_4896;
	wire n_4897;
	wire n_4898;
	wire n_4899;
	wire n_4900;
	wire n_4901;
	wire n_4902;
	wire n_4903;
	wire n_4904;
	wire n_4905;
	wire n_4906;
	wire n_4907;
	wire n_4908;
	wire n_4909;
	wire n_4910;
	wire n_4911;
	wire n_4912;
	wire n_4913;
	wire n_4914;
	wire n_4915;
	wire n_4916;
	wire n_4917;
	wire n_4918;
	wire n_4919;
	wire n_4920;
	wire n_4921;
	wire n_4922;
	wire n_4923;
	wire n_4924;
	wire n_4925;
	wire n_4926;
	wire n_4927;
	wire n_4928;
	wire n_4929;
	wire n_4930;
	wire n_4931;
	wire n_4932;
	wire n_4933;
	wire n_4934;
	wire n_4935;
	wire n_4936;
	wire n_4937;
	wire n_4938;
	wire n_4939;
	wire n_4940;
	wire n_4941;
	wire n_4942;
	wire n_4943;
	wire n_4944;
	wire n_4945;
	wire n_4946;
	wire n_4947;
	wire n_4948;
	wire n_4949;
	wire n_4950;
	wire n_4951;
	wire n_4952;
	wire n_4953;
	wire n_4954;
	wire n_4955;
	wire n_4956;
	wire n_4957;
	wire n_4958;
	wire n_4959;
	wire n_4960;
	wire n_4961;
	wire n_4962;
	wire n_4963;
	wire n_4964;
	wire n_4965;
	wire n_4966;
	wire n_4967;
	wire n_4968;
	wire n_4969;
	wire n_4970;
	wire n_4971;
	wire n_4972;
	wire n_4973;
	wire n_4974;
	wire n_4975;
	wire n_4976;
	wire n_4977;
	wire n_4978;
	wire n_4979;
	wire n_4980;
	wire n_4981;
	wire n_4982;
	wire n_4983;
	wire n_4984;
	wire n_4985;
	wire n_4986;
	wire n_4987;
	wire n_4988;
	wire n_4989;
	wire n_4990;
	wire n_4991;
	wire n_4992;
	wire n_4993;
	wire n_4994;
	wire n_4995;
	wire n_4996;
	wire n_4997;
	wire n_4998;
	wire n_4999;
	wire n_5000;
	wire n_5001;
	wire n_5002;
	wire n_5003;
	wire n_5004;
	wire n_5005;
	wire n_5006;
	wire n_5007;
	wire n_5008;
	wire n_5009;
	wire n_5010;
	wire n_5011;
	wire n_5012;
	wire n_5013;
	wire n_5014;
	wire n_5015;
	wire n_5016;
	wire n_5017;
	wire n_5018;
	wire n_5019;
	wire n_5020;
	wire n_5021;
	wire n_5022;
	wire n_5023;
	wire n_5024;
	wire n_5025;
	wire n_5026;
	wire n_5027;
	wire n_5028;
	wire n_5029;
	wire n_5030;
	wire n_5031;
	wire n_5032;
	wire n_5033;
	wire n_5034;
	wire n_5035;
	wire n_5036;
	wire n_5037;
	wire n_5038;
	wire n_5039;
	wire n_5040;
	wire n_5041;
	wire n_5042;
	wire n_5043;
	wire n_5044;
	wire n_5045;
	wire n_5046;
	wire n_5047;
	wire n_5048;
	wire n_5049;
	wire n_5050;
	wire n_5051;
	wire n_5052;
	wire n_5053;
	wire n_5054;
	wire n_5055;
	wire n_5056;
	wire n_5057;
	wire n_5058;
	wire n_5059;
	wire n_5060;
	wire n_5061;
	wire n_5062;
	wire n_5063;
	wire n_5064;
	wire n_5065;
	wire n_5066;
	wire n_5067;
	wire n_5068;
	wire n_5069;
	wire n_5070;
	wire n_5071;
	wire n_5072;
	wire n_5073;
	wire n_5074;
	wire n_5075;
	wire n_5076;
	wire n_5077;
	wire n_5078;
	wire n_5079;
	wire n_5080;
	wire n_5081;
	wire n_5082;
	wire n_5083;
	wire n_5084;
	wire n_5085;
	wire n_5086;
	wire n_5087;
	wire n_5088;
	wire n_5089;
	wire n_5090;
	wire n_5091;
	wire n_5092;
	wire n_5093;
	wire n_5094;
	wire n_5095;
	wire n_5096;
	wire n_5097;
	wire n_5098;
	wire n_5099;
	wire n_5100;
	wire n_5101;
	wire n_5102;
	wire n_5103;
	wire n_5104;
	wire n_5105;
	wire n_5106;
	wire n_5107;
	wire n_5108;
	wire n_5109;
	wire n_5110;
	wire n_5111;
	wire n_5112;
	wire n_5113;
	wire n_5114;
	wire n_5115;
	wire n_5116;
	wire n_5117;
	wire n_5118;
	wire n_5119;
	wire n_5120;
	wire n_5121;
	wire n_5122;
	wire n_5123;
	wire n_5124;
	wire n_5125;
	wire n_5126;
	wire n_5127;
	wire n_5128;
	wire n_5129;
	wire n_5130;
	wire n_5131;
	wire n_5132;
	wire n_5133;
	wire n_5134;
	wire n_5135;
	wire n_5136;
	wire n_5137;
	wire n_5138;
	wire n_5139;
	wire n_5140;
	wire n_5141;
	wire n_5142;
	wire n_5143;
	wire n_5144;
	wire n_5145;
	wire n_5146;
	wire n_5147;
	wire n_5148;
	wire n_5149;
	wire n_5150;
	wire n_5151;
	wire n_5152;
	wire n_5153;
	wire n_5154;
	wire n_5155;
	wire n_5156;
	wire n_5157;
	wire n_5158;
	wire n_5159;
	wire n_5160;
	wire n_5161;
	wire n_5162;
	wire n_5163;
	wire n_5164;
	wire n_5165;
	wire n_5166;
	wire n_5167;
	wire n_5168;
	wire n_5169;
	wire n_5170;
	wire n_5171;
	wire n_5172;
	wire n_5173;
	wire n_5174;
	wire n_5175;
	wire n_5176;
	wire n_5177;
	wire n_5178;
	wire n_5179;
	wire n_5180;
	wire n_5181;
	wire n_5182;
	wire n_5183;
	wire n_5184;
	wire n_5185;
	wire n_5186;
	wire n_5187;
	wire n_5188;
	wire n_5189;
	wire n_5190;
	wire n_5191;
	wire n_5192;
	wire n_5193;
	wire n_5194;
	wire n_5195;
	wire n_5196;
	wire n_5197;
	wire n_5198;
	wire n_5199;
	wire n_5200;
	wire n_5201;
	wire n_5202;
	wire n_5203;
	wire n_5204;
	wire n_5205;
	wire n_5206;
	wire n_5207;
	wire n_5208;
	wire n_5209;
	wire n_5210;
	wire n_5211;
	wire n_5212;
	wire n_5213;
	wire n_5214;
	wire n_5215;
	wire n_5216;
	wire n_5217;
	wire n_5218;
	wire n_5219;
	wire n_5220;
	wire n_5221;
	wire n_5222;
	wire n_5223;
	wire n_5224;
	wire n_5225;
	wire n_5226;
	wire n_5227;
	wire n_5228;
	wire n_5229;
	wire n_5230;
	wire n_5231;
	wire n_5232;
	wire n_5233;
	wire n_5234;
	wire n_5235;
	wire n_5236;
	wire n_5237;
	wire n_5238;
	wire n_5239;
	wire n_5240;
	wire n_5241;
	wire n_5242;
	wire n_5243;
	wire n_5244;
	wire n_5245;
	wire n_5246;
	wire n_5247;
	wire n_5248;
	wire n_5249;
	wire n_5250;
	wire n_5251;
	wire n_5252;
	wire n_5253;
	wire n_5254;
	wire n_5255;
	wire n_5256;
	wire n_5257;
	wire n_5258;
	wire n_5259;
	wire n_5260;
	wire n_5261;
	wire n_5262;
	wire n_5263;
	wire n_5264;
	wire n_5265;
	wire n_5266;
	wire n_5267;
	wire n_5268;
	wire n_5269;
	wire n_5270;
	wire n_5271;
	wire n_5272;
	wire n_5273;
	wire n_5274;
	wire n_5275;
	wire n_5276;
	wire n_5277;
	wire n_5278;
	wire n_5279;
	wire n_5280;
	wire n_5281;
	wire n_5282;
	wire n_5283;
	wire n_5284;
	wire n_5285;
	wire n_5286;
	wire n_5287;
	wire n_5288;
	wire n_5289;
	wire n_5290;
	wire n_5291;
	wire n_5292;
	wire n_5293;
	wire n_5294;
	wire n_5295;
	wire n_5296;
	wire n_5297;
	wire n_5298;
	wire n_5299;
	wire n_5300;
	wire n_5301;
	wire n_5302;
	wire n_5303;
	wire n_5304;
	wire n_5305;
	wire n_5306;
	wire n_5307;
	wire n_5308;
	wire n_5309;
	wire n_5310;
	wire n_5311;
	wire n_5312;
	wire n_5313;
	wire n_5314;
	wire n_5315;
	wire n_5316;
	wire n_5317;
	wire n_5318;
	wire n_5319;
	wire n_5320;
	wire n_5321;
	wire n_5322;
	wire n_5323;
	wire n_5324;
	wire n_5325;
	wire n_5326;
	wire n_5327;
	wire n_5328;
	wire n_5329;
	wire n_5330;
	wire n_5331;
	wire n_5332;
	wire n_5333;
	wire n_5334;
	wire n_5335;
	wire n_5336;
	wire n_5337;
	wire n_5338;
	wire n_5339;
	wire n_5340;
	wire n_5341;
	wire n_5342;
	wire n_5343;
	wire n_5344;
	wire n_5345;
	wire n_5346;
	wire n_5347;
	wire n_5348;
	wire n_5349;
	wire n_5350;
	wire n_5351;
	wire n_5352;
	wire n_5353;
	wire n_5354;
	wire n_5355;
	wire n_5356;
	wire n_5357;
	wire n_5358;
	wire n_5359;
	wire n_5360;
	wire n_5361;
	wire n_5362;
	wire n_5363;
	wire n_5364;
	wire n_5365;
	wire n_5366;
	wire n_5367;
	wire n_5368;
	wire n_5369;
	wire n_5370;
	wire n_5371;
	wire n_5372;
	wire n_5373;
	wire n_5374;
	wire n_5375;
	wire n_5376;
	wire n_5377;
	wire n_5378;
	wire n_5379;
	wire n_5380;
	wire n_5381;
	wire n_5382;
	wire n_5383;
	wire n_5384;
	wire n_5385;
	wire n_5386;
	wire n_5387;
	wire n_5388;
	wire n_5389;
	wire n_5390;
	wire n_5391;
	wire n_5392;
	wire n_5393;
	wire n_5394;
	wire n_5395;
	wire n_5396;
	wire n_5397;
	wire n_5398;
	wire n_5399;
	wire n_5400;
	wire n_5401;
	wire n_5402;
	wire n_5403;
	wire n_5404;
	wire n_5405;
	wire n_5406;
	wire n_5407;
	wire n_5408;
	wire n_5409;
	wire n_5410;
	wire n_5411;
	wire n_5412;
	wire n_5413;
	wire n_5414;
	wire n_5415;
	wire n_5416;
	wire n_5417;
	wire n_5418;
	wire n_5419;
	wire n_5420;
	wire n_5421;
	wire n_5422;
	wire n_5423;
	wire n_5424;
	wire n_5425;
	wire n_5426;
	wire n_5427;
	wire n_5428;
	wire n_5429;
	wire n_5430;
	wire n_5431;
	wire n_5432;
	wire n_5433;
	wire n_5434;
	wire n_5435;
	wire n_5436;
	wire n_5437;
	wire n_5438;
	wire n_5439;
	wire n_5440;
	wire n_5441;
	wire n_5442;
	wire n_5443;
	wire n_5444;
	wire n_5445;
	wire n_5446;
	wire n_5447;
	wire n_5448;
	wire n_5449;
	wire n_5450;
	wire n_5451;
	wire n_5452;
	wire n_5453;
	wire n_5454;
	wire n_5455;
	wire n_5456;
	wire n_5457;
	wire n_5458;
	wire n_5459;
	wire n_5460;
	wire n_5461;
	wire n_5462;
	wire n_5463;
	wire n_5464;
	wire n_5465;
	wire n_5466;
	wire n_5467;
	wire n_5468;
	wire n_5469;
	wire n_5470;
	wire n_5471;
	wire n_5472;
	wire n_5473;
	wire n_5474;
	wire n_5475;
	wire n_5476;
	wire n_5477;
	wire n_5478;
	wire n_5479;
	wire n_5480;
	wire n_5481;
	wire n_5482;
	wire n_5483;
	wire n_5484;
	wire n_5485;
	wire n_5486;
	wire n_5487;
	wire n_5488;
	wire n_5489;
	wire n_5490;
	wire n_5491;
	wire n_5492;
	wire n_5493;
	wire n_5494;
	wire n_5495;
	wire n_5496;
	wire n_5497;
	wire n_5498;
	wire n_5499;
	wire n_5500;
	wire n_5501;
	wire n_5502;
	wire n_5503;
	wire n_5504;
	wire n_5505;
	wire n_5506;
	wire n_5507;
	wire n_5508;
	wire n_5509;
	wire n_5510;
	wire n_5511;
	wire n_5512;
	wire n_5513;
	wire n_5514;
	wire n_5515;
	wire n_5516;
	wire n_5517;
	wire n_5518;
	wire n_5519;
	wire n_5520;
	wire n_5521;
	wire n_5522;
	wire n_5523;
	wire n_5524;
	wire n_5525;
	wire n_5526;
	wire n_5527;
	wire n_5528;
	wire n_5529;
	wire n_5530;
	wire n_5531;
	wire n_5532;
	wire n_5533;
	wire n_5534;
	wire n_5535;
	wire n_5536;
	wire n_5537;
	wire n_5538;
	wire n_5539;
	wire n_5540;
	wire n_5541;
	wire n_5542;
	wire n_5543;
	wire n_5544;
	wire n_5545;
	wire n_5546;
	wire n_5547;
	wire n_5548;
	wire n_5549;
	wire n_5550;
	wire n_5551;
	wire n_5552;
	wire n_5553;
	wire n_5554;
	wire n_5555;
	wire n_5556;
	wire n_5557;
	wire n_5558;
	wire n_5559;
	wire n_5560;
	wire n_5561;
	wire n_5562;
	wire n_5563;
	wire n_5564;
	wire n_5565;
	wire n_5566;
	wire n_5567;
	wire n_5568;
	wire n_5569;
	wire n_5570;
	wire n_5571;
	wire n_5572;
	wire n_5573;
	wire n_5574;
	wire n_5575;
	wire n_5576;
	wire n_5577;
	wire n_5578;
	wire n_5579;
	wire n_5580;
	wire n_5581;
	wire n_5582;
	wire n_5583;
	wire n_5584;
	wire n_5585;
	wire n_5586;
	wire n_5587;
	wire n_5588;
	wire n_5589;
	wire n_5590;
	wire n_5591;
	wire n_5592;
	wire n_5593;
	wire n_5594;
	wire n_5595;
	wire n_5596;
	wire n_5597;
	wire n_5598;
	wire n_5599;
	wire n_5600;
	wire n_5601;
	wire n_5602;
	wire n_5603;
	wire n_5604;
	wire n_5605;
	wire n_5606;
	wire n_5607;
	wire n_5608;
	wire n_5609;
	wire n_5610;
	wire n_5611;
	wire n_5612;
	wire n_5613;
	wire n_5614;
	wire n_5615;
	wire n_5616;
	wire n_5617;
	wire n_5618;
	wire n_5619;
	wire n_5620;
	wire n_5621;
	wire n_5622;
	wire n_5623;
	wire n_5624;
	wire n_5625;
	wire n_5626;
	wire n_5627;
	wire n_5628;
	wire n_5629;
	wire n_5630;
	wire n_5631;
	wire n_5632;
	wire n_5633;
	wire n_5634;
	wire n_5635;
	wire n_5636;
	wire n_5637;
	wire n_5638;
	wire n_5639;
	wire n_5640;
	wire n_5641;
	wire n_5642;
	wire n_5643;
	wire n_5644;
	wire n_5645;
	wire n_5646;
	wire n_5647;
	wire n_5648;
	wire n_5649;
	wire n_5650;
	wire n_5651;
	wire n_5652;
	wire n_5653;
	wire n_5654;
	wire n_5655;
	wire n_5656;
	wire n_5657;
	wire n_5658;
	wire n_5659;
	wire n_5660;
	wire n_5661;
	wire n_5662;
	wire n_5663;
	wire n_5664;
	wire n_5665;
	wire n_5666;
	wire n_5667;
	wire n_5668;
	wire n_5669;
	wire n_5670;
	wire n_5671;
	wire n_5672;
	wire n_5673;
	wire n_5674;
	wire n_5675;
	wire n_5676;
	wire n_5677;
	wire n_5678;
	wire n_5679;
	wire n_5680;
	wire n_5681;
	wire n_5682;
	wire n_5683;
	wire n_5684;
	wire n_5685;
	wire n_5686;
	wire n_5687;
	wire n_5688;
	wire n_5689;
	wire n_5690;
	wire n_5691;
	wire n_5692;
	wire n_5693;
	wire n_5694;
	wire n_5695;
	wire n_5696;
	wire n_5697;
	wire n_5698;
	wire n_5699;
	wire n_5700;
	wire n_5701;
	wire n_5702;
	wire n_5703;
	wire n_5704;
	wire n_5705;
	wire n_5706;
	wire n_5707;
	wire n_5708;
	wire n_5709;
	wire n_5710;
	wire n_5711;
	wire n_5712;
	wire n_5713;
	wire n_5714;
	wire n_5715;
	wire n_5716;
	wire n_5717;
	wire n_5718;
	wire n_5719;
	wire n_5720;
	wire n_5721;
	wire n_5722;
	wire n_5723;
	wire n_5724;
	wire n_5725;
	wire n_5726;
	wire n_5727;
	wire n_5728;
	wire n_5729;
	wire n_5730;
	wire n_5731;
	wire n_5732;
	wire n_5733;
	wire n_5734;
	wire n_5735;
	wire n_5736;
	wire n_5737;
	wire n_5738;
	wire n_5739;
	wire n_5740;
	wire n_5741;
	wire n_5742;
	wire n_5743;
	wire n_5744;
	wire n_5745;
	wire n_5746;
	wire n_5747;
	wire n_5748;
	wire n_5749;
	wire n_5750;
	wire n_5751;
	wire n_5752;
	wire n_5753;
	wire n_5754;
	wire n_5755;
	wire n_5756;
	wire n_5757;
	wire n_5758;
	wire n_5759;
	wire n_5760;
	wire n_5761;
	wire n_5762;
	wire n_5763;
	wire n_5764;
	wire n_5765;
	wire n_5766;
	wire n_5767;
	wire n_5768;
	wire n_5769;
	wire n_5770;
	wire n_5771;
	wire n_5772;
	wire n_5773;
	wire n_5774;
	wire n_5775;
	wire n_5776;
	wire n_5777;
	wire n_5778;
	wire n_5779;
	wire n_5780;
	wire n_5781;
	wire n_5782;
	wire n_5783;
	wire n_5784;
	wire n_5785;
	wire n_5786;
	wire n_5787;
	wire n_5788;
	wire n_5789;
	wire n_5790;
	wire n_5791;
	wire n_5792;
	wire n_5793;
	wire n_5794;
	wire n_5795;
	wire n_5796;
	wire n_5797;
	wire n_5798;
	wire n_5799;
	wire n_5800;
	wire n_5801;
	wire n_5802;
	wire n_5803;
	wire n_5804;
	wire n_5805;
	wire n_5806;
	wire n_5807;
	wire n_5808;
	wire n_5809;
	wire n_5810;
	wire n_5811;
	wire n_5812;
	wire n_5813;
	wire n_5814;
	wire n_5815;
	wire n_5816;
	wire n_5817;
	wire n_5818;
	wire n_5819;
	wire n_5820;
	wire n_5821;
	wire n_5822;
	wire n_5823;
	wire n_5824;
	wire n_5825;
	wire n_5826;
	wire n_5827;
	wire n_5828;
	wire n_5829;
	wire n_5830;
	wire n_5831;
	wire n_5832;
	wire n_5833;
	wire n_5834;
	wire n_5835;
	wire n_5836;
	wire n_5837;
	wire n_5838;
	wire n_5839;
	wire n_5840;
	wire n_5841;
	wire n_5842;
	wire n_5843;
	wire n_5844;
	wire n_5845;
	wire n_5846;
	wire n_5847;
	wire n_5848;
	wire n_5849;
	wire n_5850;
	wire n_5851;
	wire n_5852;
	wire n_5853;
	wire n_5854;
	wire n_5855;
	wire n_5856;
	wire n_5857;
	wire n_5858;
	wire n_5859;
	wire n_5860;
	wire n_5861;
	wire n_5862;
	wire n_5863;
	wire n_5864;
	wire n_5865;
	wire n_5866;
	wire n_5867;
	wire n_5868;
	wire n_5869;
	wire n_5870;
	wire n_5871;
	wire n_5872;
	wire n_5873;
	wire n_5874;
	wire n_5875;
	wire n_5876;
	wire n_5877;
	wire n_5878;
	wire n_5879;
	wire n_5880;
	wire n_5881;
	wire n_5882;
	wire n_5883;
	wire n_5884;
	wire n_5885;
	wire n_5886;
	wire n_5887;
	wire n_5888;
	wire n_5889;
	wire n_5890;
	wire n_5891;
	wire n_5892;
	wire n_5893;
	wire n_5894;
	wire n_5895;
	wire n_5896;
	wire n_5897;
	wire n_5898;
	wire n_5899;
	wire n_5900;
	wire n_5901;
	wire n_5902;
	wire n_5903;
	wire n_5904;
	wire n_5905;
	wire n_5906;
	wire n_5907;
	wire n_5908;
	wire n_5909;
	wire n_5910;
	wire n_5911;
	wire n_5912;
	wire n_5913;
	wire n_5914;
	wire n_5915;
	wire n_5916;
	wire n_5917;
	wire n_5918;
	wire n_5919;
	wire n_5920;
	wire n_5921;
	wire n_5922;
	wire n_5923;
	wire n_5924;
	wire n_5925;
	wire n_5926;
	wire n_5927;
	wire n_5928;
	wire n_5929;
	wire n_5930;
	wire n_5931;
	wire n_5932;
	wire n_5933;
	wire n_5934;
	wire n_5935;
	wire n_5936;
	wire n_5937;
	wire n_5938;
	wire n_5939;
	wire n_5940;
	wire n_5941;
	wire n_5942;
	wire n_5943;
	wire n_5944;
	wire n_5945;
	wire n_5946;
	wire n_5947;
	wire n_5948;
	wire n_5949;
	wire n_5950;
	wire n_5951;
	wire n_5952;
	wire n_5953;
	wire n_5954;
	wire n_5955;
	wire n_5956;
	wire n_5957;
	wire n_5958;
	wire n_5959;
	wire n_5960;
	wire n_5961;
	wire n_5962;
	wire n_5963;
	wire n_5964;
	wire n_5965;
	wire n_5966;
	wire n_5967;
	wire n_5968;
	wire n_5969;
	wire n_5970;
	wire n_5971;
	wire n_5972;
	wire n_5973;
	wire n_5974;
	wire n_5975;
	wire n_5976;
	wire n_5977;
	wire n_5978;
	wire n_5979;
	wire n_5980;
	wire n_5981;
	wire n_5982;
	wire n_5983;
	wire n_5984;
	wire n_5985;
	wire n_5986;
	wire n_5987;
	wire n_5988;
	wire n_5989;
	wire n_5990;
	wire n_5991;
	wire n_5992;
	wire n_5993;
	wire n_5994;
	wire n_5995;
	wire n_5996;
	wire n_5997;
	wire n_5998;
	wire n_5999;
	wire n_6000;
	wire n_6001;
	wire n_6002;
	wire n_6003;
	wire n_6004;
	wire n_6005;
	wire n_6006;
	wire n_6007;
	wire n_6008;
	wire n_6009;
	wire n_6010;
	wire n_6011;
	wire n_6012;
	wire n_6013;
	wire n_6014;
	wire n_6015;
	wire n_6016;
	wire n_6017;
	wire n_6018;
	wire n_6019;
	wire n_6020;
	wire n_6021;
	wire n_6022;
	wire n_6023;
	wire n_6024;
	wire n_6025;
	wire n_6026;
	wire n_6027;
	wire n_6028;
	wire n_6029;
	wire n_6030;
	wire n_6031;
	wire n_6032;
	wire n_6033;
	wire n_6034;
	wire n_6035;
	wire n_6036;
	wire n_6037;
	wire n_6038;
	wire n_6039;
	wire n_6040;
	wire n_6041;
	wire n_6042;
	wire n_6043;
	wire n_6044;
	wire n_6045;
	wire n_6046;
	wire n_6047;
	wire n_6048;
	wire n_6049;
	wire n_6050;
	wire n_6051;
	wire n_6052;
	wire n_6053;
	wire n_6054;
	wire n_6055;
	wire n_6056;
	wire n_6057;
	wire n_6058;
	wire n_6059;
	wire n_6060;
	wire n_6061;
	wire n_6062;
	wire n_6063;
	wire n_6064;
	wire n_6065;
	wire n_6066;
	wire n_6067;
	wire n_6068;
	wire n_6069;
	wire n_6070;
	wire n_6071;
	wire n_6072;
	wire n_6073;
	wire n_6074;
	wire n_6075;
	wire n_6076;
	wire n_6077;
	wire n_6078;
	wire n_6079;
	wire n_6080;
	wire n_6081;
	wire n_6082;
	wire n_6083;
	wire n_6084;
	wire n_6085;
	wire n_6086;
	wire n_6087;
	wire n_6088;
	wire n_6089;
	wire n_6090;
	wire n_6091;
	wire n_6092;
	wire n_6093;
	wire n_6094;
	wire n_6095;
	wire n_6096;
	wire n_6097;
	wire n_6098;
	wire n_6099;
	wire n_6100;
	wire n_6101;
	wire n_6102;
	wire n_6103;
	wire n_6104;
	wire n_6105;
	wire n_6106;
	wire n_6107;
	wire n_6108;
	wire n_6109;
	wire n_6110;
	wire n_6111;
	wire n_6112;
	wire n_6113;
	wire n_6114;
	wire n_6115;
	wire n_6116;
	wire n_6117;
	wire n_6118;
	wire n_6119;
	wire n_6120;
	wire n_6121;
	wire n_6122;
	wire n_6123;
	wire n_6124;
	wire n_6125;
	wire n_6126;
	wire n_6127;
	wire n_6128;
	wire n_6129;
	wire n_6130;
	wire n_6131;
	wire n_6132;
	wire n_6133;
	wire n_6134;
	wire n_6135;
	wire n_6136;
	wire n_6137;
	wire n_6138;
	wire n_6139;
	wire n_6140;
	wire n_6141;
	wire n_6142;
	wire n_6143;
	wire n_6144;
	wire n_6145;
	wire n_6146;
	wire n_6147;
	wire n_6148;
	wire n_6149;
	wire n_6150;
	wire n_6151;
	wire n_6152;
	wire n_6153;
	wire n_6154;
	wire n_6155;
	wire n_6156;
	wire n_6157;
	wire n_6158;
	wire n_6159;
	wire n_6160;
	wire n_6161;
	wire n_6162;
	wire n_6163;
	wire n_6164;
	wire n_6165;
	wire n_6166;
	wire n_6167;
	wire n_6168;
	wire n_6169;
	wire n_6170;
	wire n_6171;
	wire n_6172;
	wire n_6173;
	wire n_6174;
	wire n_6175;
	wire n_6176;
	wire n_6177;
	wire n_6178;
	wire n_6179;
	wire n_6180;
	wire n_6181;
	wire n_6182;
	wire n_6183;
	wire n_6184;
	wire n_6185;
	wire n_6186;
	wire n_6187;
	wire n_6188;
	wire n_6189;
	wire n_6190;
	wire n_6191;
	wire n_6192;
	wire n_6193;
	wire n_6194;
	wire n_6195;
	wire n_6196;
	wire n_6197;
	wire n_6198;
	wire n_6199;
	wire n_6200;
	wire n_6201;
	wire n_6202;
	wire n_6203;
	wire n_6204;
	wire n_6205;
	wire n_6206;
	wire n_6207;
	wire n_6208;
	wire n_6209;
	wire n_6210;
	wire n_6211;
	wire n_6212;
	wire n_6213;
	wire n_6214;
	wire n_6215;
	wire n_6216;
	wire n_6217;
	wire n_6218;
	wire n_6219;
	wire n_6220;
	wire n_6221;
	wire n_6222;
	wire n_6223;
	wire n_6224;
	wire n_6225;
	wire n_6226;
	wire n_6227;
	wire n_6228;
	wire n_6229;
	wire n_6230;
	wire n_6231;
	wire n_6232;
	wire n_6233;
	wire n_6234;
	wire n_6235;
	wire n_6236;
	wire n_6237;
	wire n_6238;
	wire n_6239;
	wire n_6240;
	wire n_6241;
	wire n_6242;
	wire n_6243;
	wire n_6244;
	wire n_6245;
	wire n_6246;
	wire n_6247;
	wire n_6248;
	wire n_6249;
	wire n_6250;
	wire n_6251;
	wire n_6252;
	wire n_6253;
	wire n_6254;
	wire n_6255;
	wire n_6256;
	wire n_6257;
	wire n_6258;
	wire n_6259;
	wire n_6260;
	wire n_6261;
	wire n_6262;
	wire n_6263;
	wire n_6264;
	wire n_6265;
	wire n_6266;
	wire n_6267;
	wire n_6268;
	wire n_6269;
	wire n_6270;
	wire n_6271;
	wire n_6272;
	wire n_6273;
	wire n_6274;
	wire n_6275;
	wire n_6276;
	wire n_6277;
	wire n_6278;
	wire n_6279;
	wire n_6280;
	wire n_6281;
	wire n_6282;
	wire n_6283;
	wire n_6284;
	wire n_6285;
	wire n_6286;
	wire n_6287;
	wire n_6288;
	wire n_6289;
	wire n_6290;
	wire n_6291;
	wire n_6292;
	wire n_6293;
	wire n_6294;
	wire n_6295;
	wire n_6296;
	wire n_6297;
	wire n_6298;
	wire n_6299;
	wire n_6300;
	wire n_6301;
	wire n_6302;
	wire n_6303;
	wire n_6304;
	wire n_6305;
	wire n_6306;
	wire n_6307;
	wire n_6308;
	wire n_6309;
	wire n_6310;
	wire n_6311;
	wire n_6312;
	wire n_6313;
	wire n_6314;
	wire n_6315;
	wire n_6316;
	wire n_6317;
	wire n_6318;
	wire n_6319;
	wire n_6320;
	wire n_6321;
	wire n_6322;
	wire n_6323;
	wire n_6324;
	wire n_6325;
	wire n_6326;
	wire n_6327;
	wire n_6328;
	wire n_6329;
	wire n_6330;
	wire n_6331;
	wire n_6332;
	wire n_6333;
	wire n_6334;
	wire n_6335;
	wire n_6336;
	wire n_6337;
	wire n_6338;
	wire n_6339;
	wire n_6340;
	wire n_6341;
	wire n_6342;
	wire n_6343;
	wire n_6344;
	wire n_6345;
	wire n_6346;
	wire n_6347;
	wire n_6348;
	wire n_6349;
	wire n_6350;
	wire n_6351;
	wire n_6352;
	wire n_6353;
	wire n_6354;
	wire n_6355;
	wire n_6356;
	wire n_6357;
	wire n_6358;
	wire n_6359;
	wire n_6360;
	wire n_6361;
	wire n_6362;
	wire n_6363;
	wire n_6364;
	wire n_6365;
	wire n_6366;
	wire n_6367;
	wire n_6368;
	wire n_6369;
	wire n_6370;
	wire n_6371;
	wire n_6372;
	wire n_6373;
	wire n_6374;
	wire n_6375;
	wire n_6376;
	wire n_6377;
	wire n_6378;
	wire n_6379;
	wire n_6380;
	wire n_6381;
	wire n_6382;
	wire n_6383;
	wire n_6384;
	wire n_6385;
	wire n_6386;
	wire n_6387;
	wire n_6388;
	wire n_6389;
	wire n_6390;
	wire n_6391;
	wire n_6392;
	wire n_6393;
	wire n_6394;
	wire n_6395;
	wire n_6396;
	wire n_6397;
	wire n_6398;
	wire n_6399;
	wire n_6400;
	wire n_6401;
	wire n_6402;
	wire n_6403;
	wire n_6404;
	wire n_6405;
	wire n_6406;
	wire n_6407;
	wire n_6408;
	wire n_6409;
	wire n_6410;
	wire n_6411;
	wire n_6412;
	wire n_6413;
	wire n_6414;
	wire n_6415;
	wire n_6416;
	wire n_6417;
	wire n_6418;
	wire n_6419;
	wire n_6420;
	wire n_6421;
	wire n_6422;
	wire n_6423;
	wire n_6424;
	wire n_6425;
	wire n_6426;
	wire n_6427;
	wire n_6428;
	wire n_6429;
	wire n_6430;
	wire n_6431;
	wire n_6432;
	wire n_6433;
	wire n_6434;
	wire n_6435;
	wire n_6436;
	wire n_6437;
	wire n_6438;
	wire n_6439;
	wire n_6440;
	wire n_6441;
	wire n_6442;
	wire n_6443;
	wire n_6444;
	wire n_6445;
	wire n_6446;
	wire n_6447;
	wire n_6448;
	wire n_6449;
	wire n_6450;
	wire n_6451;
	wire n_6452;
	wire n_6453;
	wire n_6454;
	wire n_6455;
	wire n_6456;
	wire n_6457;
	wire n_6458;
	wire n_6459;
	wire n_6460;
	wire n_6461;
	wire n_6462;
	wire n_6463;
	wire n_6464;
	wire n_6465;
	wire n_6466;
	wire n_6467;
	wire n_6468;
	wire n_6469;
	wire n_6470;
	wire n_6471;
	wire n_6472;
	wire n_6473;
	wire n_6474;
	wire n_6475;
	wire n_6476;
	wire n_6477;
	wire n_6478;
	wire n_6479;
	wire n_6480;
	wire n_6481;
	wire n_6482;
	wire n_6483;
	wire n_6484;
	wire n_6485;
	wire n_6486;
	wire n_6487;
	wire n_6488;
	wire n_6489;
	wire n_6490;
	wire n_6491;
	wire n_6492;
	wire n_6493;
	wire n_6494;
	wire n_6495;
	wire n_6496;
	wire n_6497;
	wire n_6498;
	wire n_6499;
	wire n_6500;
	wire n_6501;
	wire n_6502;
	wire n_6503;
	wire n_6504;
	wire n_6505;
	wire n_6506;
	wire n_6507;
	wire n_6508;
	wire n_6509;
	wire n_6510;
	wire n_6511;
	wire n_6512;
	wire n_6513;
	wire n_6514;
	wire n_6515;
	wire n_6516;
	wire n_6517;
	wire n_6518;
	wire n_6519;
	wire n_6520;
	wire n_6521;
	wire n_6522;
	wire n_6523;
	wire n_6524;
	wire n_6525;
	wire n_6526;
	wire n_6527;
	wire n_6528;
	wire n_6529;
	wire n_6530;
	wire n_6531;
	wire n_6532;
	wire n_6533;
	wire n_6534;
	wire n_6535;
	wire n_6536;
	wire n_6537;
	wire n_6538;
	wire n_6539;
	wire n_6540;
	wire n_6541;
	wire n_6542;
	wire n_6543;
	wire n_6544;
	wire n_6545;
	wire n_6546;
	wire n_6547;
	wire n_6548;
	wire n_6549;
	wire n_6550;
	wire n_6551;
	wire n_6552;
	wire n_6553;
	wire n_6554;
	wire n_6555;
	wire n_6556;
	wire n_6557;
	wire n_6558;
	wire n_6559;
	wire n_6560;
	wire n_6561;
	wire n_6562;
	wire n_6563;
	wire n_6564;
	wire n_6565;
	wire n_6566;
	wire n_6567;
	wire n_6568;
	wire n_6569;
	wire n_6570;
	wire n_6571;
	wire n_6572;
	wire n_6573;
	wire n_6574;
	wire n_6575;
	wire n_6576;
	wire n_6577;
	wire n_6578;
	wire n_6579;
	wire n_6580;
	wire n_6581;
	wire n_6582;
	wire n_6583;
	wire n_6584;
	wire n_6585;
	wire n_6586;
	wire n_6587;
	wire n_6588;
	wire n_6589;
	wire n_6590;
	wire n_6591;
	wire n_6592;
	wire n_6593;
	wire n_6594;
	wire n_6595;
	wire n_6596;
	wire n_6597;
	wire n_6598;
	wire n_6599;
	wire n_6600;
	wire n_6601;
	wire n_6602;
	wire n_6603;
	wire n_6604;
	wire n_6605;
	wire n_6606;
	wire n_6607;
	wire n_6608;
	wire n_6609;
	wire n_6610;
	wire n_6611;
	wire n_6612;
	wire n_6613;
	wire n_6614;
	wire n_6615;
	wire n_6616;
	wire n_6617;
	wire n_6618;
	wire n_6619;
	wire n_6620;
	wire n_6621;
	wire n_6622;
	wire n_6623;
	wire n_6624;
	wire n_6625;
	wire n_6626;
	wire n_6627;
	wire n_6628;
	wire n_6629;
	wire n_6630;
	wire n_6631;
	wire n_6632;
	wire n_6633;
	wire n_6634;
	wire n_6635;
	wire n_6636;
	wire n_6637;
	wire n_6638;
	wire n_6639;
	wire n_6640;
	wire n_6641;
	wire n_6642;
	wire n_6643;
	wire n_6644;
	wire n_6645;
	wire n_6646;
	wire n_6647;
	wire n_6648;
	wire n_6649;
	wire n_6650;
	wire n_6651;
	wire n_6652;
	wire n_6653;
	wire n_6654;
	wire n_6655;
	wire n_6656;
	wire n_6657;
	wire n_6658;
	wire n_6659;
	wire n_6660;
	wire n_6661;
	wire n_6662;
	wire n_6663;
	wire n_6664;
	wire n_6665;
	wire n_6666;
	wire n_6667;
	wire n_6668;
	wire n_6669;
	wire n_6670;
	wire n_6671;
	wire n_6672;
	wire n_6673;
	wire n_6674;
	wire n_6675;
	wire n_6676;
	wire n_6677;
	wire n_6678;
	wire n_6679;
	wire n_6680;
	wire n_6681;
	wire n_6682;
	wire n_6683;
	wire n_6684;
	wire n_6685;
	wire n_6686;
	wire n_6687;
	wire n_6688;
	wire n_6689;
	wire n_6690;
	wire n_6691;
	wire n_6692;
	wire n_6693;
	wire n_6694;
	wire n_6695;
	wire n_6696;
	wire n_6697;
	wire n_6698;
	wire n_6699;
	wire n_6700;
	wire n_6701;
	wire n_6702;
	wire n_6703;
	wire n_6704;
	wire n_6705;
	wire n_6706;
	wire n_6707;
	wire n_6708;
	wire n_6709;
	wire n_6710;
	wire n_6711;
	wire n_6712;
	wire n_6713;
	wire n_6714;
	wire n_6715;
	wire n_6716;
	wire n_6717;
	wire n_6718;
	wire n_6719;
	wire n_6720;
	wire n_6721;
	wire n_6722;
	wire n_6723;
	wire n_6724;
	wire n_6725;
	wire n_6726;
	wire n_6727;
	wire n_6728;
	wire n_6729;
	wire n_6730;
	wire n_6731;
	wire n_6732;
	wire n_6733;
	wire n_6734;
	wire n_6735;
	wire n_6736;
	wire n_6737;
	wire n_6738;
	wire n_6739;
	wire n_6740;
	wire n_6741;
	wire n_6742;
	wire n_6743;
	wire n_6744;
	wire n_6745;
	wire n_6746;
	wire n_6747;
	wire n_6748;
	wire n_6749;
	wire n_6750;
	wire n_6751;
	wire n_6752;
	wire n_6753;
	wire n_6754;
	wire n_6755;
	wire n_6756;
	wire n_6757;
	wire n_6758;
	wire n_6759;
	wire n_6760;
	wire n_6761;
	wire n_6762;
	wire n_6763;
	wire n_6764;
	wire n_6765;
	wire n_6766;
	wire n_6767;
	wire n_6768;
	wire n_6769;
	wire n_6770;
	wire n_6771;
	wire n_6772;
	wire n_6773;
	wire n_6774;
	wire n_6775;
	wire n_6776;
	wire n_6777;
	wire n_6778;
	wire n_6779;
	wire n_6780;
	wire n_6781;
	wire n_6782;
	wire n_6783;
	wire n_6784;
	wire n_6785;
	wire n_6786;
	wire n_6787;
	wire n_6788;
	wire n_6789;
	wire n_6790;
	wire n_6791;
	wire n_6792;
	wire n_6793;
	wire n_6794;
	wire n_6795;
	wire n_6796;
	wire n_6797;
	wire n_6798;
	wire n_6799;
	wire n_6800;
	wire n_6801;
	wire n_6802;
	wire n_6803;
	wire n_6804;
	wire n_6805;
	wire n_6806;
	wire n_6807;
	wire n_6808;
	wire n_6809;
	wire n_6810;
	wire n_6811;
	wire n_6812;
	wire n_6813;
	wire n_6814;
	wire n_6815;
	wire n_6816;
	wire n_6817;
	wire n_6818;
	wire n_6819;
	wire n_6820;
	wire n_6821;
	wire n_6822;
	wire n_6823;
	wire n_6824;
	wire n_6825;
	wire n_6826;
	wire n_6827;
	wire n_6828;
	wire n_6829;
	wire n_6830;
	wire n_6831;
	wire n_6832;
	wire n_6833;
	wire n_6834;
	wire n_6835;
	wire n_6836;
	wire n_6837;
	wire n_6838;
	wire n_6839;
	wire n_6840;
	wire n_6841;
	wire n_6842;
	wire n_6843;
	wire n_6844;
	wire n_6845;
	wire n_6846;
	wire n_6847;
	wire n_6848;
	wire n_6849;
	wire n_6850;
	wire n_6851;
	wire n_6852;
	wire n_6853;
	wire n_6854;
	wire n_6855;
	wire n_6856;
	wire n_6857;
	wire n_6858;
	wire n_6859;
	wire n_6860;
	wire n_6861;
	wire n_6862;
	wire n_6863;
	wire n_6864;
	wire n_6865;
	wire n_6866;
	wire n_6867;
	wire n_6868;
	wire n_6869;
	wire n_6870;
	wire n_6871;
	wire n_6872;
	wire n_6873;
	wire n_6874;
	wire n_6875;
	wire n_6876;
	wire n_6877;
	wire n_6878;
	wire n_6879;
	wire n_6880;
	wire n_6881;
	wire n_6882;
	wire n_6883;
	wire n_6884;
	wire n_6885;
	wire n_6886;
	wire n_6887;
	wire n_6888;
	wire n_6889;
	wire n_6890;
	wire n_6891;
	wire n_6892;
	wire n_6893;
	wire n_6894;
	wire n_6895;
	wire n_6896;
	wire n_6897;
	wire n_6898;
	wire n_6899;
	wire n_6900;
	wire n_6901;
	wire n_6902;
	wire n_6903;
	wire n_6904;
	wire n_6905;
	wire n_6906;
	wire n_6907;
	wire n_6908;
	wire n_6909;
	wire n_6910;
	wire n_6911;
	wire n_6912;
	wire n_6913;
	wire n_6914;
	wire n_6915;
	wire n_6916;
	wire n_6917;
	wire n_6918;
	wire n_6919;
	wire n_6920;
	wire n_6921;
	wire n_6922;
	wire n_6923;
	wire n_6924;
	wire n_6925;
	wire n_6926;
	wire n_6927;
	wire n_6928;
	wire n_6929;
	wire n_6930;
	wire n_6931;
	wire n_6932;
	wire n_6933;
	wire n_6934;
	wire n_6935;
	wire n_6936;
	wire n_6937;
	wire n_6938;
	wire n_6939;
	wire n_6940;
	wire n_6941;
	wire n_6942;
	wire n_6943;
	wire n_6944;
	wire n_6945;
	wire n_6946;
	wire n_6947;
	wire n_6948;
	wire n_6949;
	wire n_6950;
	wire n_6951;
	wire n_6952;
	wire n_6953;
	wire n_6954;
	wire n_6955;
	wire n_6956;
	wire n_6957;
	wire n_6958;
	wire n_6959;
	wire n_6960;
	wire n_6961;
	wire n_6962;
	wire n_6963;
	wire n_6964;
	wire n_6965;
	wire n_6966;
	wire n_6967;
	wire n_6968;
	wire n_6969;
	wire n_6970;
	wire n_6971;
	wire n_6972;
	wire n_6973;
	wire n_6974;
	wire n_6975;
	wire n_6976;
	wire n_6977;
	wire n_6978;
	wire n_6979;
	wire n_6980;
	wire n_6981;
	wire n_6982;
	wire n_6983;
	wire n_6984;
	wire n_6985;
	wire n_6986;
	wire n_6987;
	wire n_6988;
	wire n_6989;
	wire n_6990;
	wire n_6991;
	wire n_6992;
	wire n_6993;
	wire n_6994;
	wire n_6995;
	wire n_6996;
	wire n_6997;
	wire n_6998;
	wire n_6999;
	wire n_7000;
	wire n_7001;
	wire n_7002;
	wire n_7003;
	wire n_7004;
	wire n_7005;
	wire n_7006;
	wire n_7007;
	wire n_7008;
	wire n_7009;
	wire n_7010;
	wire n_7011;
	wire n_7012;
	wire n_7013;
	wire n_7014;
	wire n_7015;
	wire n_7016;
	wire n_7017;
	wire n_7018;
	wire n_7019;
	wire n_7020;
	wire n_7021;
	wire n_7022;
	wire n_7023;
	wire n_7024;
	wire n_7025;
	wire n_7026;
	wire n_7027;
	wire n_7028;
	wire n_7029;
	wire n_7030;
	wire n_7031;
	wire n_7032;
	wire n_7033;
	wire n_7034;
	wire n_7035;
	wire n_7036;
	wire n_7037;
	wire n_7038;
	wire n_7039;
	wire n_7040;
	wire n_7041;
	wire n_7042;
	wire n_7043;
	wire n_7044;
	wire n_7045;
	wire n_7046;
	wire n_7047;
	wire n_7048;
	wire n_7049;
	wire n_7050;
	wire n_7051;
	wire n_7052;
	wire n_7053;
	wire n_7054;
	wire n_7055;
	wire n_7056;
	wire n_7057;
	wire n_7058;
	wire n_7059;
	wire n_7060;
	wire n_7061;
	wire n_7062;
	wire n_7063;
	wire n_7064;
	wire n_7065;
	wire n_7066;
	wire n_7067;
	wire n_7068;
	wire n_7069;
	wire n_7070;
	wire n_7071;
	wire n_7072;
	wire n_7073;
	wire n_7074;
	wire n_7075;
	wire n_7076;
	wire n_7077;
	wire n_7078;
	wire n_7079;
	wire n_7080;
	wire n_7081;
	wire n_7082;
	wire n_7083;
	wire n_7084;
	wire n_7085;
	wire n_7086;
	wire n_7087;
	wire n_7088;
	wire n_7089;
	wire n_7090;
	wire n_7091;
	wire n_7092;
	wire n_7093;
	wire n_7094;
	wire n_7095;
	wire n_7096;
	wire n_7097;
	wire n_7098;
	wire n_7099;
	wire n_7100;
	wire n_7101;
	wire n_7102;
	wire n_7103;
	wire n_7104;
	wire n_7105;
	wire n_7106;
	wire n_7107;
	wire n_7108;
	wire n_7109;
	wire n_7110;
	wire n_7111;
	wire n_7112;
	wire n_7113;
	wire n_7114;
	wire n_7115;
	wire n_7116;
	wire n_7117;
	wire n_7118;
	wire n_7119;
	wire n_7120;
	wire n_7121;
	wire n_7122;
	wire n_7123;
	wire n_7124;
	wire n_7125;
	wire n_7126;
	wire n_7127;
	wire n_7128;
	wire n_7129;
	wire n_7130;
	wire n_7131;
	wire n_7132;
	wire n_7133;
	wire n_7134;
	wire n_7135;
	wire n_7136;
	wire n_7137;
	wire n_7138;
	wire n_7139;
	wire n_7140;
	wire n_7141;
	wire n_7142;
	wire n_7143;
	wire n_7144;
	wire n_7145;
	wire n_7146;
	wire n_7147;
	wire n_7148;
	wire n_7149;
	wire n_7150;
	wire n_7151;
	wire n_7152;
	wire n_7153;
	wire n_7154;
	wire n_7155;
	wire n_7156;
	wire n_7157;
	wire n_7158;
	wire n_7159;
	wire n_7160;
	wire n_7161;
	wire n_7162;
	wire n_7163;
	wire n_7164;
	wire n_7165;
	wire n_7166;
	wire n_7167;
	wire n_7168;
	wire n_7169;
	wire n_7170;
	wire n_7171;
	wire n_7172;
	wire n_7173;
	wire n_7174;
	wire n_7175;
	wire n_7176;
	wire n_7177;
	wire n_7178;
	wire n_7179;
	wire n_7180;
	wire n_7181;
	wire n_7182;
	wire n_7183;
	wire n_7184;
	wire n_7185;
	wire n_7186;
	wire n_7187;
	wire n_7188;
	wire n_7189;
	wire n_7190;
	wire n_7191;
	wire n_7192;
	wire n_7193;
	wire n_7194;
	wire n_7195;
	wire n_7196;
	wire n_7197;
	wire n_7198;
	wire n_7199;
	wire n_7200;
	wire n_7201;
	wire n_7202;
	wire n_7203;
	wire n_7204;
	wire n_7205;
	wire n_7206;
	wire n_7207;
	wire n_7208;
	wire n_7209;
	wire n_7210;
	wire n_7211;
	wire n_7212;
	wire n_7213;
	wire n_7214;
	wire n_7215;
	wire n_7216;
	wire n_7217;
	wire n_7218;
	wire n_7219;
	wire n_7220;
	wire n_7221;
	wire n_7222;
	wire n_7223;
	wire n_7224;
	wire n_7225;
	wire n_7226;
	wire n_7227;
	wire n_7228;
	wire n_7229;
	wire n_7230;
	wire n_7231;
	wire n_7232;
	wire n_7233;
	wire n_7234;
	wire n_7235;
	wire n_7236;
	wire n_7237;
	wire n_7238;
	wire n_7239;
	wire n_7240;
	wire n_7241;
	wire n_7242;
	wire n_7243;
	wire n_7244;
	wire n_7245;
	wire n_7246;
	wire n_7247;
	wire n_7248;
	wire n_7249;
	wire n_7250;
	wire n_7251;
	wire n_7252;
	wire n_7253;
	wire n_7254;
	wire n_7255;
	wire n_7256;
	wire n_7257;
	wire n_7258;
	wire n_7259;
	wire n_7260;
	wire n_7261;
	wire n_7262;
	wire n_7263;
	wire n_7264;
	wire n_7265;
	wire n_7266;
	wire n_7267;
	wire n_7268;
	wire n_7269;
	wire n_7270;
	wire n_7271;
	wire n_7272;
	wire n_7273;
	wire n_7274;
	wire n_7275;
	wire n_7276;
	wire n_7277;
	wire n_7278;
	wire n_7279;
	wire n_7280;
	wire n_7281;
	wire n_7282;
	wire n_7283;
	wire n_7284;
	wire n_7285;
	wire n_7286;
	wire n_7287;
	wire n_7288;
	wire n_7289;
	wire n_7290;
	wire n_7291;
	wire n_7292;
	wire n_7293;
	wire n_7294;
	wire n_7295;
	wire n_7296;
	wire n_7297;
	wire n_7298;
	wire n_7299;
	wire n_7300;
	wire n_7301;
	wire n_7302;
	wire n_7303;
	wire n_7304;
	wire n_7305;
	wire n_7306;
	wire n_7307;
	wire n_7308;
	wire n_7309;
	wire n_7310;
	wire n_7311;
	wire n_7312;
	wire n_7313;
	wire n_7314;
	wire n_7315;
	wire n_7316;
	wire n_7317;
	wire n_7318;
	wire n_7319;
	wire n_7320;
	wire n_7321;
	wire n_7322;
	wire n_7323;
	wire n_7324;
	wire n_7325;
	wire n_7326;
	wire n_7327;
	wire n_7328;
	wire n_7329;
	wire n_7330;
	wire n_7331;
	wire n_7332;
	wire n_7333;
	wire n_7334;
	wire n_7335;
	wire n_7336;
	wire n_7337;
	wire n_7338;
	wire n_7339;
	wire n_7340;
	wire n_7341;
	wire n_7342;
	wire n_7343;
	wire n_7344;
	wire n_7345;
	wire n_7346;
	wire n_7347;
	wire n_7348;
	wire n_7349;
	wire n_7350;
	wire n_7351;
	wire n_7352;
	wire n_7353;
	wire n_7354;
	wire n_7355;
	wire n_7356;
	wire n_7357;
	wire n_7358;
	wire n_7359;
	wire n_7360;
	wire n_7361;
	wire n_7362;
	wire n_7363;
	wire n_7364;
	wire n_7365;
	wire n_7366;
	wire n_7367;
	wire n_7368;
	wire n_7369;
	wire n_7370;
	wire n_7371;
	wire n_7372;
	wire n_7373;
	wire n_7374;
	wire n_7375;
	wire n_7376;
	wire n_7377;
	wire n_7378;
	wire n_7379;
	wire n_7380;
	wire n_7381;
	wire n_7382;
	wire n_7383;
	wire n_7384;
	wire n_7385;
	wire n_7386;
	wire n_7387;
	wire n_7388;
	wire n_7389;
	wire n_7390;
	wire n_7391;
	wire n_7392;
	wire n_7393;
	wire n_7394;
	wire n_7395;
	wire n_7396;
	wire n_7397;
	wire n_7398;
	wire n_7399;
	wire n_7400;
	wire n_7401;
	wire n_7402;
	wire n_7403;
	wire n_7404;
	wire n_7405;
	wire n_7406;
	wire n_7407;
	wire n_7408;
	wire n_7409;
	wire n_7410;
	wire n_7411;
	wire n_7412;
	wire n_7413;
	wire n_7414;
	wire n_7415;
	wire n_7416;
	wire n_7417;
	wire n_7418;
	wire n_7419;
	wire n_7420;
	wire n_7421;
	wire n_7422;
	wire n_7423;
	wire n_7424;
	wire n_7425;
	wire n_7426;
	wire n_7427;
	wire n_7428;
	wire n_7429;
	wire n_7430;
	wire n_7431;
	wire n_7432;
	wire n_7433;
	wire n_7434;
	wire n_7435;
	wire n_7436;
	wire n_7437;
	wire n_7438;
	wire n_7439;
	wire n_7440;
	wire n_7441;
	wire n_7442;
	wire n_7443;
	wire n_7444;
	wire n_7445;
	wire n_7446;
	wire n_7447;
	wire n_7448;
	wire n_7449;
	wire n_7450;
	wire n_7451;
	wire n_7452;
	wire n_7453;
	wire n_7454;
	wire n_7455;
	wire n_7456;
	wire n_7457;
	wire n_7458;
	wire n_7459;
	wire n_7460;
	wire n_7461;
	wire n_7462;
	wire n_7463;
	wire n_7464;
	wire n_7465;
	wire n_7466;
	wire n_7467;
	wire n_7468;
	wire n_7469;
	wire n_7470;
	wire n_7471;
	wire n_7472;
	wire n_7473;
	wire n_7474;
	wire n_7475;
	wire n_7476;
	wire n_7477;
	wire n_7478;
	wire n_7479;
	wire n_7480;
	wire n_7481;
	wire n_7482;
	wire n_7483;
	wire n_7484;
	wire n_7485;
	wire n_7486;
	wire n_7487;
	wire n_7488;
	wire n_7489;
	wire n_7490;
	wire n_7491;
	wire n_7492;
	wire n_7493;
	wire n_7494;
	wire n_7495;
	wire n_7496;
	wire n_7497;
	wire n_7498;
	wire n_7499;
	wire n_7500;
	wire n_7501;
	wire n_7502;
	wire n_7503;
	wire n_7504;
	wire n_7505;
	wire n_7506;
	wire n_7507;
	wire n_7508;
	wire n_7509;
	wire n_7510;
	wire n_7511;
	wire n_7512;
	wire n_7513;
	wire n_7514;
	wire n_7515;
	wire n_7516;
	wire n_7517;
	wire n_7518;
	wire n_7519;
	wire n_7520;
	wire n_7521;
	wire n_7522;
	wire n_7523;
	wire n_7524;
	wire n_7525;
	wire n_7526;
	wire n_7527;
	wire n_7528;
	wire n_7529;
	wire n_7530;
	wire n_7531;
	wire n_7532;
	wire n_7533;
	wire n_7534;
	wire n_7535;
	wire n_7536;
	wire n_7537;
	wire n_7538;
	wire n_7539;
	wire n_7540;
	wire n_7541;
	wire n_7542;
	wire n_7543;
	wire n_7544;
	wire n_7545;
	wire n_7546;
	wire n_7547;
	wire n_7548;
	wire n_7549;
	wire n_7550;
	wire n_7551;
	wire n_7552;
	wire n_7553;
	wire n_7554;
	wire n_7555;
	wire n_7556;
	wire n_7557;
	wire n_7558;
	wire n_7559;
	wire n_7560;
	wire n_7561;
	wire n_7562;
	wire n_7563;
	wire n_7564;
	wire n_7565;
	wire n_7566;
	wire n_7567;
	wire n_7568;
	wire n_7569;
	wire n_7570;
	wire n_7571;
	wire n_7572;
	wire n_7573;
	wire n_7574;
	wire n_7575;
	wire n_7576;
	wire n_7577;
	wire n_7578;
	wire n_7579;
	wire n_7580;
	wire n_7581;
	wire n_7582;
	wire n_7583;
	wire n_7584;
	wire n_7585;
	wire n_7586;
	wire n_7587;
	wire n_7588;
	wire n_7589;
	wire n_7590;
	wire n_7591;
	wire n_7592;
	wire n_7593;
	wire n_7594;
	wire n_7595;
	wire n_7596;
	wire n_7597;
	wire n_7598;
	wire n_7599;
	wire n_7600;
	wire n_7601;
	wire n_7602;
	wire n_7603;
	wire n_7604;
	wire n_7605;
	wire n_7606;
	wire n_7607;
	wire n_7608;
	wire n_7609;
	wire n_7610;
	wire n_7611;
	wire n_7612;
	wire n_7613;
	wire n_7614;
	wire n_7615;
	wire n_7616;
	wire n_7617;
	wire n_7618;
	wire n_7619;
	wire n_7620;
	wire n_7621;
	wire n_7622;
	wire n_7623;
	wire n_7624;
	wire n_7625;
	wire n_7626;
	wire n_7627;
	wire n_7628;
	wire n_7629;
	wire n_7630;
	wire n_7631;
	wire n_7632;
	wire n_7633;
	wire n_7634;
	wire n_7635;
	wire n_7636;
	wire n_7637;
	wire n_7638;
	wire n_7639;
	wire n_7640;
	wire n_7641;
	wire n_7642;
	wire n_7643;
	wire n_7644;
	wire n_7645;
	wire n_7646;
	wire n_7647;
	wire n_7648;
	wire n_7649;
	wire n_7650;
	wire n_7651;
	wire n_7652;
	wire n_7653;
	wire n_7654;
	wire n_7655;
	wire n_7656;
	wire n_7657;
	wire n_7658;
	wire n_7659;
	wire n_7660;
	wire n_7661;
	wire n_7662;
	wire n_7663;
	wire n_7664;
	wire n_7665;
	wire n_7666;
	wire n_7667;
	wire n_7668;
	wire n_7669;
	wire n_7670;
	wire n_7671;
	wire n_7672;
	wire n_7673;
	wire n_7674;
	wire n_7675;
	wire n_7676;
	wire n_7677;
	wire n_7678;
	wire n_7679;
	wire n_7680;
	wire n_7681;
	wire n_7682;
	wire n_7683;
	wire n_7684;
	wire n_7685;
	wire n_7686;
	wire n_7687;
	wire n_7688;
	wire n_7689;
	wire n_7690;
	wire n_7691;
	wire n_7692;
	wire n_7693;
	wire n_7694;
	wire n_7695;
	wire n_7696;
	wire n_7697;
	wire n_7698;
	wire n_7699;
	wire n_7700;
	wire n_7701;
	wire n_7702;
	wire n_7703;
	wire n_7704;
	wire n_7705;
	wire n_7706;
	wire n_7707;
	wire n_7708;
	wire n_7709;
	wire n_7710;
	wire n_7711;
	wire n_7712;
	wire n_7713;
	wire n_7714;
	wire n_7715;
	wire n_7716;
	wire n_7717;
	wire n_7718;
	wire n_7719;
	wire n_7720;
	wire n_7721;
	wire n_7722;
	wire n_7723;
	wire n_7724;
	wire n_7725;
	wire n_7726;
	wire n_7727;
	wire n_7728;
	wire n_7729;
	wire n_7730;
	wire n_7731;
	wire n_7732;
	wire n_7733;
	wire n_7734;
	wire n_7735;
	wire n_7736;
	wire n_7737;
	wire n_7738;
	wire n_7739;
	wire n_7740;
	wire n_7741;
	wire n_7742;
	wire n_7743;
	wire n_7744;
	wire n_7745;
	wire n_7746;
	wire n_7747;
	wire n_7748;
	wire n_7749;
	wire n_7750;
	wire n_7751;
	wire n_7752;
	wire n_7753;
	wire n_7754;
	wire n_7755;
	wire n_7756;
	wire n_7757;
	wire n_7758;
	wire n_7759;
	wire n_7760;
	wire n_7761;
	wire n_7762;
	wire n_7763;
	wire n_7764;
	wire n_7765;
	wire n_7766;
	wire n_7767;
	wire n_7768;
	wire n_7769;
	wire n_7770;
	wire n_7771;
	wire n_7772;
	wire n_7773;
	wire n_7774;
	wire n_7775;
	wire n_7776;
	wire n_7777;
	wire n_7778;
	wire n_7779;
	wire n_7780;
	wire n_7781;
	wire n_7782;
	wire n_7783;
	wire n_7784;
	wire n_7785;
	wire n_7786;
	wire n_7787;
	wire n_7788;
	wire n_7789;
	wire n_7790;
	wire n_7791;
	wire n_7792;
	wire n_7793;
	wire n_7794;
	wire n_7795;
	wire n_7796;
	wire n_7797;
	wire n_7798;
	wire n_7799;
	wire n_7800;
	wire n_7801;
	wire n_7802;
	wire n_7803;
	wire n_7804;
	wire n_7805;
	wire n_7806;
	wire n_7807;
	wire n_7808;
	wire n_7809;
	wire n_7810;
	wire n_7811;
	wire n_7812;
	wire n_7813;
	wire n_7814;
	wire n_7815;
	wire n_7816;
	wire n_7817;
	wire n_7818;
	wire n_7819;
	wire n_7820;
	wire n_7821;
	wire n_7822;
	wire n_7823;
	wire n_7824;
	wire n_7825;
	wire n_7826;
	wire n_7827;
	wire n_7828;
	wire n_7829;
	wire n_7830;
	wire n_7831;
	wire n_7832;
	wire n_7833;
	wire n_7834;
	wire n_7835;
	wire n_7836;
	wire n_7837;
	wire n_7838;
	wire n_7839;
	wire n_7840;
	wire n_7841;
	wire n_7842;
	wire n_7843;
	wire n_7844;
	wire n_7845;
	wire n_7846;
	wire n_7847;
	wire n_7848;
	wire n_7849;
	wire n_7850;
	wire n_7851;
	wire n_7852;
	wire n_7853;
	wire n_7854;
	wire n_7855;
	wire n_7856;
	wire n_7857;
	wire n_7858;
	wire n_7859;
	wire n_7860;
	wire n_7861;
	wire n_7862;
	wire n_7863;
	wire n_7864;
	wire n_7865;
	wire n_7866;
	wire n_7867;
	wire n_7868;
	wire n_7869;
	wire n_7870;
	wire n_7871;
	wire n_7872;
	wire n_7873;
	wire n_7874;
	wire n_7875;
	wire n_7876;
	wire n_7877;
	wire n_7878;
	wire n_7879;
	wire n_7880;
	wire n_7881;
	wire n_7882;
	wire n_7883;
	wire n_7884;
	wire n_7885;
	wire n_7886;
	wire n_7887;
	wire n_7888;
	wire n_7889;
	wire n_7890;
	wire n_7891;
	wire n_7892;
	wire n_7893;
	wire n_7894;
	wire n_7895;
	wire n_7896;
	wire n_7897;
	wire n_7898;
	wire n_7899;
	wire n_7900;
	wire n_7901;
	wire n_7902;
	wire n_7903;
	wire n_7904;
	wire n_7905;
	wire n_7906;
	wire n_7907;
	wire n_7908;
	wire n_7909;
	wire n_7910;
	wire n_7911;
	wire n_7912;
	wire n_7913;
	wire n_7914;
	wire n_7915;
	wire n_7916;
	wire n_7917;
	wire n_7918;
	wire n_7919;
	wire n_7920;
	wire n_7921;
	wire n_7922;
	wire n_7923;
	wire n_7924;
	wire n_7925;
	wire n_7926;
	wire n_7927;
	wire n_7928;
	wire n_7929;
	wire n_7930;
	wire n_7931;
	wire n_7932;
	wire n_7933;
	wire n_7934;
	wire n_7935;
	wire n_7936;
	wire n_7937;
	wire n_7938;
	wire n_7939;
	wire n_7940;
	wire n_7941;
	wire n_7942;
	wire n_7943;
	wire n_7944;
	wire n_7945;
	wire n_7946;
	wire n_7947;
	wire n_7948;
	wire n_7949;
	wire n_7950;
	wire n_7951;
	wire n_7952;
	wire n_7953;
	wire n_7954;
	wire n_7955;
	wire n_7956;
	wire n_7957;
	wire n_7958;
	wire n_7959;
	wire n_7960;
	wire n_7961;
	wire n_7962;
	wire n_7963;
	wire n_7964;
	wire n_7965;
	wire n_7966;
	wire n_7967;
	wire n_7968;
	wire n_7969;
	wire n_7970;
	wire n_7971;
	wire n_7972;
	wire n_7973;
	wire n_7974;
	wire n_7975;
	wire n_7976;
	wire n_7977;
	wire n_7978;
	wire n_7979;
	wire n_7980;
	wire n_7981;
	wire n_7982;
	wire n_7983;
	wire n_7984;
	wire n_7985;
	wire n_7986;
	wire n_7987;
	wire n_7988;
	wire n_7989;
	wire n_7990;
	wire n_7991;
	wire n_7992;
	wire n_7993;
	wire n_7994;
	wire n_7995;
	wire n_7996;
	wire n_7997;
	wire n_7998;
	wire n_7999;
	wire n_8000;
	wire n_8001;
	wire n_8002;
	wire n_8003;
	wire n_8004;
	wire n_8005;
	wire n_8006;
	wire n_8007;
	wire n_8008;
	wire n_8009;
	wire n_8010;
	wire n_8011;
	wire n_8012;
	wire n_8013;
	wire n_8014;
	wire n_8015;
	wire n_8016;
	wire n_8017;
	wire n_8018;
	wire n_8019;
	wire n_8020;
	wire n_8021;
	wire n_8022;
	wire n_8023;
	wire n_8024;
	wire n_8025;
	wire n_8026;
	wire n_8027;
	wire n_8028;
	wire n_8029;
	wire n_8030;
	wire n_8031;
	wire n_8032;
	wire n_8033;
	wire n_8034;
	wire n_8035;
	wire n_8036;
	wire n_8037;
	wire n_8038;
	wire n_8039;
	wire n_8040;
	wire n_8041;
	wire n_8042;
	wire n_8043;
	wire n_8044;
	wire n_8045;
	wire n_8046;
	wire n_8047;
	wire n_8048;
	wire n_8049;
	wire n_8050;
	wire n_8051;
	wire n_8052;
	wire n_8053;
	wire n_8054;
	wire n_8055;
	wire n_8056;
	wire n_8057;
	wire n_8058;
	wire n_8059;
	wire n_8060;
	wire n_8061;
	wire n_8062;
	wire n_8063;
	wire n_8064;
	wire n_8065;
	wire n_8066;
	wire n_8067;
	wire n_8068;
	wire n_8069;
	wire n_8070;
	wire n_8071;
	wire n_8072;
	wire n_8073;
	wire n_8074;
	wire n_8075;
	wire n_8076;
	wire n_8077;
	wire n_8078;
	wire n_8079;
	wire n_8080;
	wire n_8081;
	wire n_8082;
	wire n_8083;
	wire n_8084;
	wire n_8085;
	wire n_8086;
	wire n_8087;
	wire n_8088;
	wire n_8089;
	wire n_8090;
	wire n_8091;
	wire n_8092;
	wire n_8093;
	wire n_8094;
	wire n_8095;
	wire n_8096;
	wire n_8097;
	wire n_8098;
	wire n_8099;
	wire n_8100;
	wire n_8101;
	wire n_8102;
	wire n_8103;
	wire n_8104;
	wire n_8105;
	wire n_8106;
	wire n_8107;
	wire n_8108;
	wire n_8109;
	wire n_8110;
	wire n_8111;
	wire n_8112;
	wire n_8113;
	wire n_8114;
	wire n_8115;
	wire n_8116;
	wire n_8117;
	wire n_8118;
	wire n_8119;
	wire n_8120;
	wire n_8121;
	wire n_8122;
	wire n_8123;
	wire n_8124;
	wire n_8125;
	wire n_8126;
	wire n_8127;
	wire n_8128;
	wire n_8129;
	wire n_8130;
	wire n_8131;
	wire n_8132;
	wire n_8133;
	wire n_8134;
	wire n_8135;
	wire n_8136;
	wire n_8137;
	wire n_8138;
	wire n_8139;
	wire n_8140;
	wire n_8141;
	wire n_8142;
	wire n_8143;
	wire n_8144;
	wire n_8145;
	wire n_8146;
	wire n_8147;
	wire n_8148;
	wire n_8149;
	wire n_8150;
	wire n_8151;
	wire n_8152;
	wire n_8153;
	wire n_8154;
	wire n_8155;
	wire n_8156;
	wire n_8157;
	wire n_8158;
	wire n_8159;
	wire n_8160;
	wire n_8161;
	wire n_8162;
	wire n_8163;
	wire n_8164;
	wire n_8165;
	wire n_8166;
	wire n_8167;
	wire n_8168;
	wire n_8169;
	wire n_8170;
	wire n_8171;
	wire n_8172;
	wire n_8173;
	wire n_8174;
	wire n_8175;
	wire n_8176;
	wire n_8177;
	wire n_8178;
	wire n_8179;
	wire n_8180;
	wire n_8181;
	wire n_8182;
	wire n_8183;
	wire n_8184;
	wire n_8185;
	wire n_8186;
	wire n_8187;
	wire n_8188;
	wire n_8189;
	wire n_8190;
	wire n_8191;
	wire n_8192;
	wire n_8193;
	wire n_8194;
	wire n_8195;
	wire n_8196;
	wire n_8197;
	wire n_8198;
	wire n_8199;
	wire n_8200;
	wire n_8201;
	wire n_8202;
	wire n_8203;
	wire n_8204;
	wire n_8205;
	wire n_8206;
	wire n_8207;
	wire n_8208;
	wire n_8209;
	wire n_8210;
	wire n_8211;
	wire n_8212;
	wire n_8213;
	wire n_8214;
	wire n_8215;
	wire n_8216;
	wire n_8217;
	wire n_8218;
	wire n_8219;
	wire n_8220;
	wire n_8221;
	wire n_8222;
	wire n_8223;
	wire n_8224;
	wire n_8225;
	wire n_8226;
	wire n_8227;
	wire n_8228;
	wire n_8229;
	wire n_8230;
	wire n_8231;
	wire n_8232;
	wire n_8233;
	wire n_8234;
	wire n_8235;
	wire n_8236;
	wire n_8237;
	wire n_8238;
	wire n_8239;
	wire n_8240;
	wire n_8241;
	wire n_8242;
	wire n_8243;
	wire n_8244;
	wire n_8245;
	wire n_8246;
	wire n_8247;
	wire n_8248;
	wire n_8249;
	wire n_8250;
	wire n_8251;
	wire n_8252;
	wire n_8253;
	wire n_8254;
	wire n_8255;
	wire n_8256;
	wire n_8257;
	wire n_8258;
	wire n_8259;
	wire n_8260;
	wire n_8261;
	wire n_8262;
	wire n_8263;
	wire n_8264;
	wire n_8265;
	wire n_8266;
	wire n_8267;
	wire n_8268;
	wire n_8269;
	wire n_8270;
	wire n_8271;
	wire n_8272;
	wire n_8273;
	wire n_8274;
	wire n_8275;
	wire n_8276;
	wire n_8277;
	wire n_8278;
	wire n_8279;
	wire n_8280;
	wire n_8281;
	wire n_8282;
	wire n_8283;
	wire n_8284;
	wire n_8285;
	wire n_8286;
	wire n_8287;
	wire n_8288;
	wire n_8289;
	wire n_8290;
	wire n_8291;
	wire n_8292;
	wire n_8293;
	wire n_8294;
	wire n_8295;
	wire n_8296;
	wire n_8297;
	wire n_8298;
	wire n_8299;
	wire n_8300;
	wire n_8301;
	wire n_8302;
	wire n_8303;
	wire n_8304;
	wire n_8305;
	wire n_8306;
	wire n_8307;
	wire n_8308;
	wire n_8309;
	wire n_8310;
	wire n_8311;
	wire n_8312;
	wire n_8313;
	wire n_8314;
	wire n_8315;
	wire n_8316;
	wire n_8317;
	wire n_8318;
	wire n_8319;
	wire n_8320;
	wire n_8321;
	wire n_8322;
	wire n_8323;
	wire n_8324;
	wire n_8325;
	wire n_8326;
	wire n_8327;
	wire n_8328;
	wire n_8329;
	wire n_8330;
	wire n_8331;
	wire n_8332;
	wire n_8333;
	wire n_8334;
	wire n_8335;
	wire n_8336;
	wire n_8337;
	wire n_8338;
	wire n_8339;
	wire n_8340;
	wire n_8341;
	wire n_8342;
	wire n_8343;
	wire n_8344;
	wire n_8345;
	wire n_8346;
	wire n_8347;
	wire n_8348;
	wire n_8349;
	wire n_8350;
	wire n_8351;
	wire n_8352;
	wire n_8353;
	wire n_8354;
	wire n_8355;
	wire n_8356;
	wire n_8357;
	wire n_8358;
	wire n_8359;
	wire n_8360;
	wire n_8361;
	wire n_8362;
	wire n_8363;
	wire n_8364;
	wire n_8365;
	wire n_8366;
	wire n_8367;
	wire n_8368;
	wire n_8369;
	wire n_8370;
	wire n_8371;
	wire n_8372;
	wire n_8373;
	wire n_8374;
	wire n_8375;
	wire n_8376;
	wire n_8377;
	wire n_8378;
	wire n_8379;
	wire n_8380;
	wire n_8381;
	wire n_8382;
	wire n_8383;
	wire n_8384;
	wire n_8385;
	wire n_8386;
	wire n_8387;
	wire n_8388;
	wire n_8389;
	wire n_8390;
	wire n_8391;
	wire n_8392;
	wire n_8393;
	wire n_8394;
	wire n_8395;
	wire n_8396;
	wire n_8397;
	wire n_8398;
	wire n_8399;
	wire n_8400;
	wire n_8401;
	wire n_8402;
	output o_1;
	assign n_706 = (x_298 & ~x_718) ;
	assign n_702 = (~x_718 & x_804) ;
	assign n_707 = (~x_101 & ~n_706) ;
	assign n_705 = (x_651 & x_718) ;
	assign n_703 = (x_101 & ~n_702) ;
	assign n_701 = (x_603 & x_718) ;
	assign n_718 = (x_367 & ~x_718) ;
	assign n_714 = (~x_718 & x_781) ;
	assign n_708 = (~n_705 & n_707) ;
	assign n_704 = (~n_701 & n_703) ;
	assign n_719 = (~x_101 & ~n_718) ;
	assign n_717 = (x_172 & x_718) ;
	assign n_715 = (x_101 & ~n_714) ;
	assign n_713 = (x_682 & x_718) ;
	assign n_709 = (~n_704 & ~n_708) ;
	assign n_720 = (~n_717 & n_719) ;
	assign n_716 = (~n_713 & n_715) ;
	assign n_710 = (x_576 & n_709) ;
	assign n_731 = (x_450 & ~x_718) ;
	assign n_727 = (x_702 & ~x_718) ;
	assign n_721 = (~n_716 & ~n_720) ;
	assign n_712 = (x_493 & n_710) ;
	assign n_732 = (~x_101 & ~n_731) ;
	assign n_730 = (x_250 & x_718) ;
	assign n_728 = (x_101 & ~n_727) ;
	assign n_726 = (x_150 & x_718) ;
	assign n_722 = (~n_712 & ~n_721) ;
	assign n_711 = (~x_493 & ~n_710) ;
	assign n_733 = (~n_730 & n_732) ;
	assign n_729 = (~n_726 & n_728) ;
	assign n_723 = (~n_711 & ~n_722) ;
	assign n_744 = (x_377 & ~x_718) ;
	assign n_740 = (x_106 & ~x_718) ;
	assign n_734 = (~n_729 & ~n_733) ;
	assign n_725 = (x_320 & n_723) ;
	assign n_745 = (~x_101 & ~n_744) ;
	assign n_743 = (x_329 & x_718) ;
	assign n_741 = (x_101 & ~n_740) ;
	assign n_739 = (x_718 & x_818) ;
	assign n_735 = (~n_725 & ~n_734) ;
	assign n_724 = (~x_320 & ~n_723) ;
	assign n_746 = (~n_743 & n_745) ;
	assign n_742 = (~n_739 & n_741) ;
	assign n_736 = (~n_724 & ~n_735) ;
	assign n_757 = (x_310 & ~x_718) ;
	assign n_753 = (x_197 & ~x_718) ;
	assign n_747 = (~n_742 & ~n_746) ;
	assign n_738 = (x_391 & n_736) ;
	assign n_758 = (~x_101 & ~n_757) ;
	assign n_756 = (x_499 & x_718) ;
	assign n_754 = (x_101 & ~n_753) ;
	assign n_752 = (x_718 & x_749) ;
	assign n_748 = (~n_738 & ~n_747) ;
	assign n_737 = (~x_391 & ~n_736) ;
	assign n_759 = (~n_756 & n_758) ;
	assign n_755 = (~n_752 & n_754) ;
	assign n_749 = (~n_737 & ~n_748) ;
	assign n_770 = (x_503 & ~x_718) ;
	assign n_766 = (x_635 & ~x_718) ;
	assign n_760 = (~n_755 & ~n_759) ;
	assign n_751 = (x_436 & n_749) ;
	assign n_771 = (~x_101 & ~n_770) ;
	assign n_769 = (x_428 & x_718) ;
	assign n_767 = (x_101 & ~n_766) ;
	assign n_765 = (x_718 & x_817) ;
	assign n_761 = (~n_751 & ~n_760) ;
	assign n_750 = (~x_436 & ~n_749) ;
	assign n_772 = (~n_769 & n_771) ;
	assign n_768 = (~n_765 & n_767) ;
	assign n_762 = (~n_750 & ~n_761) ;
	assign n_783 = (x_590 & ~x_718) ;
	assign n_779 = (x_549 & ~x_718) ;
	assign n_773 = (~n_768 & ~n_772) ;
	assign n_764 = (x_359 & n_762) ;
	assign n_784 = (~x_101 & ~n_783) ;
	assign n_782 = (x_381 & x_718) ;
	assign n_780 = (x_101 & ~n_779) ;
	assign n_778 = (x_718 & x_766) ;
	assign n_774 = (~n_764 & ~n_773) ;
	assign n_763 = (~x_359 & ~n_762) ;
	assign n_9 = (~x_255 & ~x_578) ;
	assign n_13 = (x_255 & x_578) ;
	assign n_147 = (x_77 & ~x_255) ;
	assign n_146 = (x_99 & ~x_578) ;
	assign n_138 = (~x_527 & x_706) ;
	assign n_137 = (x_277 & x_527) ;
	assign n_785 = (~n_782 & n_784) ;
	assign n_781 = (~n_778 & n_780) ;
	assign n_775 = (~n_763 & ~n_774) ;
	assign n_151 = (x_595 & n_9) ;
	assign n_150 = (x_290 & n_13) ;
	assign n_148 = (~n_146 & ~n_147) ;
	assign n_142 = (~x_527 & x_641) ;
	assign n_141 = (x_340 & x_527) ;
	assign n_139 = (~n_137 & ~n_138) ;
	assign n_796 = (x_246 & ~x_718) ;
	assign n_792 = (x_267 & ~x_718) ;
	assign n_786 = (~n_781 & ~n_785) ;
	assign n_777 = (x_447 & n_775) ;
	assign n_152 = (~n_150 & ~n_151) ;
	assign n_149 = (~n_9 & ~n_148) ;
	assign n_143 = (~n_141 & ~n_142) ;
	assign n_140 = (x_726 & ~n_139) ;
	assign n_797 = (~x_101 & ~n_796) ;
	assign n_795 = (x_459 & x_718) ;
	assign n_793 = (x_101 & ~n_792) ;
	assign n_791 = (x_684 & x_718) ;
	assign n_787 = (~n_777 & ~n_786) ;
	assign n_776 = (~x_447 & ~n_775) ;
	assign n_153 = (~n_149 & n_152) ;
	assign n_145 = (n_140 & ~n_143) ;
	assign n_127 = (x_183 & ~x_578) ;
	assign n_126 = (~x_255 & x_741) ;
	assign n_798 = (~n_795 & n_797) ;
	assign n_794 = (~n_791 & n_793) ;
	assign n_788 = (~n_776 & ~n_787) ;
	assign n_154 = (~n_145 & n_153) ;
	assign n_144 = (~n_140 & n_143) ;
	assign n_135 = (x_162 & ~x_527) ;
	assign n_134 = (x_392 & x_527) ;
	assign n_131 = (x_512 & n_9) ;
	assign n_130 = (x_213 & n_13) ;
	assign n_128 = (~n_126 & ~n_127) ;
	assign n_809 = (x_165 & ~x_718) ;
	assign n_805 = (x_348 & ~x_718) ;
	assign n_799 = (~n_794 & ~n_798) ;
	assign n_790 = (x_529 & n_788) ;
	assign n_155 = (~n_144 & ~n_154) ;
	assign n_136 = (~n_134 & ~n_135) ;
	assign n_132 = (~n_130 & ~n_131) ;
	assign n_129 = (~n_9 & ~n_128) ;
	assign n_119 = (~x_578 & x_646) ;
	assign n_118 = (~x_255 & x_805) ;
	assign n_810 = (~x_101 & ~n_809) ;
	assign n_808 = (x_364 & x_718) ;
	assign n_806 = (x_101 & ~n_805) ;
	assign n_804 = (x_126 & x_718) ;
	assign n_800 = (~n_790 & ~n_799) ;
	assign n_789 = (~x_529 & ~n_788) ;
	assign n_156 = (~n_136 & n_155) ;
	assign n_133 = (~n_129 & n_132) ;
	assign n_123 = (x_440 & n_9) ;
	assign n_122 = (x_608 & n_13) ;
	assign n_120 = (~n_118 & ~n_119) ;
	assign n_811 = (~n_808 & n_810) ;
	assign n_807 = (~n_804 & n_806) ;
	assign n_801 = (~n_789 & ~n_800) ;
	assign n_158 = (n_136 & ~n_155) ;
	assign n_157 = (n_133 & ~n_156) ;
	assign n_124 = (~n_122 & ~n_123) ;
	assign n_121 = (~n_9 & ~n_120) ;
	assign n_822 = (x_657 & ~x_718) ;
	assign n_818 = (x_482 & ~x_718) ;
	assign n_812 = (~n_807 & ~n_811) ;
	assign n_803 = (x_307 & n_801) ;
	assign n_168 = (x_564 & ~x_578) ;
	assign n_167 = (~x_255 & x_776) ;
	assign n_163 = (x_524 & ~x_527) ;
	assign n_162 = (x_446 & x_527) ;
	assign n_159 = (~n_157 & ~n_158) ;
	assign n_125 = (~n_121 & n_124) ;
	assign n_823 = (~x_101 & ~n_822) ;
	assign n_821 = (x_291 & x_718) ;
	assign n_819 = (x_101 & ~n_818) ;
	assign n_817 = (x_218 & x_718) ;
	assign n_813 = (~n_803 & ~n_812) ;
	assign n_802 = (~x_307 & ~n_801) ;
	assign n_172 = (x_374 & n_9) ;
	assign n_171 = (x_688 & n_13) ;
	assign n_169 = (~n_167 & ~n_168) ;
	assign n_164 = (~n_162 & ~n_163) ;
	assign n_161 = (~n_125 & n_159) ;
	assign n_824 = (~n_821 & n_823) ;
	assign n_820 = (~n_817 & n_819) ;
	assign n_814 = (~n_802 & ~n_813) ;
	assign n_173 = (~n_171 & ~n_172) ;
	assign n_170 = (~n_9 & ~n_169) ;
	assign n_165 = (~n_161 & n_164) ;
	assign n_160 = (n_125 & ~n_159) ;
	assign n_109 = (x_252 & ~x_578) ;
	assign n_108 = (~x_255 & x_694) ;
	assign n_835 = (x_412 & ~x_718) ;
	assign n_831 = (x_128 & ~x_718) ;
	assign n_825 = (~n_820 & ~n_824) ;
	assign n_816 = (x_220 & n_814) ;
	assign n_178 = (~x_527 & x_591) ;
	assign n_177 = (x_511 & x_527) ;
	assign n_174 = (~n_170 & n_173) ;
	assign n_166 = (~n_160 & ~n_165) ;
	assign n_113 = (x_445 & n_9) ;
	assign n_112 = (x_143 & n_13) ;
	assign n_110 = (~n_108 & ~n_109) ;
	assign n_836 = (~x_101 & ~n_835) ;
	assign n_834 = (x_544 & x_718) ;
	assign n_832 = (x_101 & ~n_831) ;
	assign n_830 = (x_718 & x_816) ;
	assign n_826 = (~n_816 & ~n_825) ;
	assign n_815 = (~x_220 & ~n_814) ;
	assign n_179 = (~n_177 & ~n_178) ;
	assign n_176 = (n_166 & ~n_174) ;
	assign n_114 = (~n_112 & ~n_113) ;
	assign n_111 = (~n_9 & ~n_110) ;
	assign n_106 = (~x_527 & x_658) ;
	assign n_105 = (x_125 & x_527) ;
	assign n_837 = (~n_834 & n_836) ;
	assign n_833 = (~n_830 & n_832) ;
	assign n_827 = (~n_815 & ~n_826) ;
	assign n_180 = (~n_176 & n_179) ;
	assign n_175 = (~n_166 & n_174) ;
	assign n_115 = (~n_111 & n_114) ;
	assign n_107 = (~n_105 & ~n_106) ;
	assign n_98 = (x_114 & ~x_255) ;
	assign n_97 = (x_334 & ~x_578) ;
	assign n_848 = (x_400 & ~x_718) ;
	assign n_844 = (~x_718 & x_808) ;
	assign n_838 = (~n_833 & ~n_837) ;
	assign n_829 = (x_247 & n_827) ;
	assign n_181 = (~n_175 & ~n_180) ;
	assign n_117 = (n_107 & n_115) ;
	assign n_102 = (x_375 & n_9) ;
	assign n_101 = (x_813 & n_13) ;
	assign n_99 = (~n_97 & ~n_98) ;
	assign n_849 = (~x_101 & ~n_848) ;
	assign n_847 = (x_620 & x_718) ;
	assign n_845 = (x_101 & ~n_844) ;
	assign n_843 = (x_146 & x_718) ;
	assign n_839 = (~n_829 & ~n_838) ;
	assign n_828 = (~x_247 & ~n_827) ;
	assign n_182 = (~n_117 & n_181) ;
	assign n_116 = (~n_107 & ~n_115) ;
	assign n_103 = (~n_101 & ~n_102) ;
	assign n_100 = (~n_9 & ~n_99) ;
	assign n_850 = (~n_847 & n_849) ;
	assign n_846 = (~n_843 & n_845) ;
	assign n_840 = (~n_828 & ~n_839) ;
	assign n_192 = (x_203 & ~x_255) ;
	assign n_191 = (x_496 & ~x_578) ;
	assign n_187 = (~x_527 & x_725) ;
	assign n_186 = (x_199 & x_527) ;
	assign n_183 = (~n_116 & ~n_182) ;
	assign n_104 = (~n_100 & n_103) ;
	assign n_861 = (x_474 & ~x_718) ;
	assign n_857 = (~x_718 & x_760) ;
	assign n_851 = (~n_846 & ~n_850) ;
	assign n_842 = (x_166 & n_840) ;
	assign n_196 = (x_309 & n_9) ;
	assign n_195 = (x_752 & n_13) ;
	assign n_193 = (~n_191 & ~n_192) ;
	assign n_188 = (~n_186 & ~n_187) ;
	assign n_185 = (n_104 & n_183) ;
	assign n_862 = (~x_101 & ~n_861) ;
	assign n_860 = (x_211 & x_718) ;
	assign n_858 = (x_101 & ~n_857) ;
	assign n_856 = (x_685 & x_718) ;
	assign n_852 = (~n_842 & ~n_851) ;
	assign n_841 = (~x_166 & ~n_840) ;
	assign n_197 = (~n_195 & ~n_196) ;
	assign n_194 = (~n_9 & ~n_193) ;
	assign n_189 = (~n_185 & ~n_188) ;
	assign n_184 = (~n_104 & ~n_183) ;
	assign n_863 = (~n_860 & n_862) ;
	assign n_859 = (~n_856 & n_858) ;
	assign n_853 = (~n_841 & ~n_852) ;
	assign n_207 = (x_424 & ~x_578) ;
	assign n_206 = (~x_255 & x_625) ;
	assign n_202 = (~x_527 & x_785) ;
	assign n_201 = (x_527 & x_654) ;
	assign n_198 = (~n_194 & n_197) ;
	assign n_190 = (~n_184 & ~n_189) ;
	assign n_874 = (x_555 & ~x_718) ;
	assign n_870 = (x_73 & ~x_718) ;
	assign n_864 = (~n_859 & ~n_863) ;
	assign n_855 = (x_659 & n_853) ;
	assign n_211 = (x_506 & n_9) ;
	assign n_210 = (x_820 & n_13) ;
	assign n_208 = (~n_206 & ~n_207) ;
	assign n_203 = (~n_201 & ~n_202) ;
	assign n_200 = (n_190 & n_198) ;
	assign n_875 = (~x_101 & ~n_874) ;
	assign n_873 = (x_120 & x_718) ;
	assign n_871 = (x_101 & ~n_870) ;
	assign n_869 = (x_601 & x_718) ;
	assign n_865 = (~n_855 & ~n_864) ;
	assign n_854 = (~x_659 & ~n_853) ;
	assign n_212 = (~n_210 & ~n_211) ;
	assign n_209 = (~n_9 & ~n_208) ;
	assign n_204 = (~n_200 & ~n_203) ;
	assign n_199 = (~n_190 & ~n_198) ;
	assign n_88 = (x_385 & ~x_578) ;
	assign n_87 = (~x_255 & x_548) ;
	assign n_876 = (~n_873 & n_875) ;
	assign n_872 = (~n_869 & n_871) ;
	assign n_866 = (~n_854 & ~n_865) ;
	assign n_217 = (x_83 & ~x_527) ;
	assign n_216 = (x_527 & x_586) ;
	assign n_213 = (~n_209 & n_212) ;
	assign n_205 = (~n_199 & ~n_204) ;
	assign n_92 = (x_593 & n_9) ;
	assign n_91 = (x_762 & n_13) ;
	assign n_89 = (~n_87 & ~n_88) ;
	assign n_888 = (x_281 & ~x_718) ;
	assign n_884 = (~x_718 & x_755) ;
	assign n_877 = (~n_872 & ~n_876) ;
	assign n_868 = (x_738 & n_866) ;
	assign n_218 = (~n_216 & ~n_217) ;
	assign n_215 = (n_205 & n_213) ;
	assign n_93 = (~n_91 & ~n_92) ;
	assign n_90 = (~n_9 & ~n_89) ;
	assign n_85 = (~x_527 & x_764) ;
	assign n_84 = (x_518 & x_527) ;
	assign n_889 = (~x_101 & ~n_888) ;
	assign n_887 = (x_689 & x_718) ;
	assign n_885 = (x_101 & ~n_884) ;
	assign n_883 = (x_219 & x_718) ;
	assign n_878 = (~n_868 & ~n_877) ;
	assign n_867 = (~x_738 & ~n_866) ;
	assign n_219 = (~n_215 & ~n_218) ;
	assign n_214 = (~n_205 & ~n_213) ;
	assign n_94 = (~n_90 & n_93) ;
	assign n_86 = (~n_84 & ~n_85) ;
	assign n_77 = (x_111 & ~x_255) ;
	assign n_76 = (x_559 & ~x_578) ;
	assign n_890 = (~n_887 & n_889) ;
	assign n_886 = (~n_883 & n_885) ;
	assign n_879 = (~n_867 & ~n_878) ;
	assign n_220 = (~n_214 & ~n_219) ;
	assign n_96 = (n_86 & n_94) ;
	assign n_81 = (x_346 & n_9) ;
	assign n_80 = (x_79 & n_13) ;
	assign n_78 = (~n_76 & ~n_77) ;
	assign n_1141 = (x_193 & ~x_718) ;
	assign n_1137 = (x_675 & ~x_718) ;
	assign n_891 = (~n_886 & ~n_890) ;
	assign n_881 = (x_806 & n_879) ;
	assign n_221 = (~n_96 & ~n_220) ;
	assign n_95 = (~n_86 & ~n_94) ;
	assign n_82 = (~n_80 & ~n_81) ;
	assign n_79 = (~n_9 & ~n_78) ;
	assign n_1142 = (~x_101 & ~n_1141) ;
	assign n_1140 = (x_718 & x_768) ;
	assign n_1138 = (x_101 & ~n_1137) ;
	assign n_1136 = (x_300 & x_718) ;
	assign n_1131 = (~n_881 & ~n_891) ;
	assign n_880 = (~x_806 & ~n_879) ;
	assign n_231 = (x_276 & ~x_578) ;
	assign n_230 = (~x_255 & x_693) ;
	assign n_226 = (~x_527 & x_696) ;
	assign n_225 = (x_455 & x_527) ;
	assign n_222 = (~n_95 & ~n_221) ;
	assign n_83 = (~n_79 & n_82) ;
	assign n_1143 = (~n_1140 & n_1142) ;
	assign n_1139 = (~n_1136 & n_1138) ;
	assign n_1132 = (~n_880 & ~n_1131) ;
	assign n_235 = (x_413 & n_9) ;
	assign n_234 = (x_748 & n_13) ;
	assign n_232 = (~n_230 & ~n_231) ;
	assign n_227 = (~n_225 & ~n_226) ;
	assign n_224 = (n_83 & n_222) ;
	assign n_1788 = (x_618 & ~x_718) ;
	assign n_1784 = (x_145 & ~x_718) ;
	assign n_1144 = (~n_1139 & ~n_1143) ;
	assign n_1134 = (x_775 & n_1132) ;
	assign n_236 = (~n_234 & ~n_235) ;
	assign n_233 = (~n_9 & ~n_232) ;
	assign n_228 = (~n_224 & ~n_227) ;
	assign n_223 = (~n_83 & ~n_222) ;
	assign n_1789 = (~x_101 & ~n_1788) ;
	assign n_1787 = (x_718 & x_811) ;
	assign n_1785 = (x_101 & ~n_1784) ;
	assign n_1783 = (x_536 & x_718) ;
	assign n_1778 = (~n_1134 & ~n_1144) ;
	assign n_1133 = (~x_775 & ~n_1132) ;
	assign n_246 = (x_189 & ~x_578) ;
	assign n_245 = (~x_255 & x_774) ;
	assign n_241 = (~x_527 & x_629) ;
	assign n_240 = (x_396 & x_527) ;
	assign n_237 = (~n_233 & n_236) ;
	assign n_229 = (~n_223 & ~n_228) ;
	assign n_1790 = (~n_1787 & n_1789) ;
	assign n_1786 = (~n_1783 & n_1785) ;
	assign n_1779 = (~n_1133 & ~n_1778) ;
	assign n_250 = (x_489 & n_9) ;
	assign n_249 = (x_667 & n_13) ;
	assign n_247 = (~n_245 & ~n_246) ;
	assign n_242 = (~n_240 & ~n_241) ;
	assign n_239 = (n_229 & n_237) ;
	assign n_1920 = (x_708 & ~x_718) ;
	assign n_1916 = (x_231 & ~x_718) ;
	assign n_1791 = (~n_1786 & ~n_1790) ;
	assign n_1781 = (x_699 & n_1779) ;
	assign n_251 = (~n_249 & ~n_250) ;
	assign n_248 = (~n_9 & ~n_247) ;
	assign n_243 = (~n_239 & ~n_242) ;
	assign n_238 = (~n_229 & ~n_237) ;
	assign n_1921 = (~x_101 & ~n_1920) ;
	assign n_1919 = (x_718 & x_744) ;
	assign n_1917 = (x_101 & ~n_1916) ;
	assign n_1915 = (x_456 & x_718) ;
	assign n_1911 = (~n_1781 & ~n_1791) ;
	assign n_1780 = (~x_699 & ~n_1779) ;
	assign n_261 = (~x_578 & x_621) ;
	assign n_260 = (~x_255 & x_807) ;
	assign n_256 = (~x_527 & x_565) ;
	assign n_255 = (x_343 & x_527) ;
	assign n_252 = (~n_248 & n_251) ;
	assign n_244 = (~n_238 & ~n_243) ;
	assign n_1922 = (~n_1919 & n_1921) ;
	assign n_1918 = (~n_1915 & n_1917) ;
	assign n_1912 = (~n_1780 & ~n_1911) ;
	assign n_46 = (x_101 & ~x_697) ;
	assign n_7619 = (x_140 & n_94) ;
	assign n_7618 = (~x_140 & ~n_94) ;
	assign n_265 = (x_342 & n_9) ;
	assign n_264 = (x_152 & n_13) ;
	assign n_262 = (~n_260 & ~n_261) ;
	assign n_257 = (~n_255 & ~n_256) ;
	assign n_254 = (n_244 & n_252) ;
	assign n_1933 = (x_121 & ~x_718) ;
	assign n_1929 = (x_606 & ~x_718) ;
	assign n_1923 = (~n_1918 & ~n_1922) ;
	assign n_1914 = (x_112 & n_1912) ;
	assign n_62 = (i_1 & ~i_2) ;
	assign n_47 = (x_718 & n_46) ;
	assign n_44 = (~x_101 & ~x_718) ;
	assign n_7620 = (~n_7618 & ~n_7619) ;
	assign n_266 = (~n_264 & ~n_265) ;
	assign n_263 = (~n_9 & ~n_262) ;
	assign n_258 = (~n_254 & ~n_257) ;
	assign n_253 = (~n_244 & ~n_252) ;
	assign n_1934 = (~x_101 & ~n_1933) ;
	assign n_1932 = (x_69 & x_718) ;
	assign n_1930 = (x_101 & ~n_1929) ;
	assign n_1928 = (x_356 & x_718) ;
	assign n_1924 = (~n_1914 & ~n_1923) ;
	assign n_1913 = (~x_112 & ~n_1912) ;
	assign n_1 = (~x_168 & ~x_664) ;
	assign n_63 = (~i_3 & n_62) ;
	assign n_48 = (x_777 & ~n_47) ;
	assign n_45 = (x_697 & n_44) ;
	assign n_4 = (~i_1 & ~i_2) ;
	assign n_2 = (~i_1 & i_2) ;
	assign n_7622 = (n_220 & n_7620) ;
	assign n_527 = (~x_332 & x_664) ;
	assign n_276 = (~x_578 & x_710) ;
	assign n_275 = (~x_255 & x_740) ;
	assign n_271 = (x_205 & ~x_527) ;
	assign n_270 = (x_462 & x_527) ;
	assign n_267 = (~n_263 & n_266) ;
	assign n_259 = (~n_253 & ~n_258) ;
	assign n_1935 = (~n_1932 & n_1934) ;
	assign n_1931 = (~n_1928 & n_1930) ;
	assign n_1925 = (~n_1913 & ~n_1924) ;
	assign n_64 = (n_63 & n_1) ;
	assign n_59 = (x_168 & ~x_664) ;
	assign n_49 = (~n_45 & n_48) ;
	assign n_43 = (x_638 & x_777) ;
	assign n_5 = (i_3 & n_4) ;
	assign n_3 = (~i_3 & n_2) ;
	assign n_7623 = (n_527 & ~n_7622) ;
	assign n_7621 = (~n_220 & ~n_7620) ;
	assign n_280 = (x_261 & n_9) ;
	assign n_279 = (x_236 & n_13) ;
	assign n_277 = (~n_275 & ~n_276) ;
	assign n_272 = (~n_270 & ~n_271) ;
	assign n_269 = (n_259 & n_267) ;
	assign n_1946 = (~x_718 & x_798) ;
	assign n_1942 = (x_522 & ~x_718) ;
	assign n_1936 = (~n_1931 & ~n_1935) ;
	assign n_1927 = (x_201 & n_1925) ;
	assign n_65 = (~n_59 & ~n_64) ;
	assign n_50 = (n_43 & ~n_49) ;
	assign n_6 = (~n_3 & ~n_5) ;
	assign n_7624 = (~n_7621 & n_7623) ;
	assign n_14 = (x_332 & ~n_13) ;
	assign n_12 = (~x_168 & x_664) ;
	assign n_10 = (x_332 & ~n_9) ;
	assign n_8 = (x_168 & x_664) ;
	assign n_281 = (~n_279 & ~n_280) ;
	assign n_278 = (~n_9 & ~n_277) ;
	assign n_273 = (~n_269 & ~n_272) ;
	assign n_268 = (~n_259 & ~n_267) ;
	assign n_1947 = (~x_101 & ~n_1946) ;
	assign n_1945 = (x_157 & x_718) ;
	assign n_1943 = (x_101 & ~n_1942) ;
	assign n_1941 = (x_433 & x_718) ;
	assign n_1937 = (~n_1927 & ~n_1936) ;
	assign n_1926 = (~x_201 & ~n_1925) ;
	assign n_7643 = (i_65 & n_59) ;
	assign n_66 = (i_5 & ~n_65) ;
	assign n_60 = (i_5 & ~n_59) ;
	assign n_53 = (i_5 & n_50) ;
	assign n_51 = (i_5 & ~n_50) ;
	assign n_5833 = (~i_45 & ~n_6) ;
	assign n_947 = (i_5 & n_1) ;
	assign n_7626 = (n_86 & ~n_7624) ;
	assign n_29 = (i_5 & ~n_1) ;
	assign n_629 = (~x_697 & ~x_777) ;
	assign n_15 = (n_12 & n_14) ;
	assign n_11 = (n_8 & n_10) ;
	assign n_282 = (~n_278 & n_281) ;
	assign n_274 = (~n_268 & ~n_273) ;
	assign n_1948 = (~n_1945 & n_1947) ;
	assign n_1944 = (~n_1941 & n_1943) ;
	assign n_1938 = (~n_1926 & ~n_1937) ;
	assign n_7644 = (n_66 & n_7643) ;
	assign n_7642 = (x_517 & n_60) ;
	assign n_7637 = (x_416 & n_53) ;
	assign n_7636 = (x_516 & n_51) ;
	assign n_7630 = (n_947 & ~n_5833) ;
	assign n_7629 = (n_6 & n_86) ;
	assign n_7627 = (n_29 & ~n_7626) ;
	assign n_7625 = (~n_86 & n_7624) ;
	assign n_936 = (n_629 & n_3) ;
	assign n_7 = (n_1 & ~n_6) ;
	assign n_16 = (~n_11 & ~n_15) ;
	assign n_284 = (n_274 & n_282) ;
	assign n_283 = (~n_274 & ~n_282) ;
	assign n_1960 = (x_93 & ~x_718) ;
	assign n_1956 = (x_577 & ~x_718) ;
	assign n_1949 = (~n_1944 & ~n_1948) ;
	assign n_1940 = (x_627 & n_1938) ;
	assign n_7645 = (~n_7642 & ~n_7644) ;
	assign n_7638 = (~n_7636 & ~n_7637) ;
	assign n_7631 = (~n_7629 & n_7630) ;
	assign n_7628 = (~n_7625 & n_7627) ;
	assign n_7612 = (~x_519 & ~n_936) ;
	assign n_7604 = (i_20 & n_7) ;
	assign n_7603 = (x_341 & ~n_16) ;
	assign n_17 = (~n_7 & n_16) ;
	assign n_7560 = (~n_283 & ~n_284) ;
	assign n_1961 = (~x_101 & ~n_1960) ;
	assign n_1959 = (x_98 & x_718) ;
	assign n_1957 = (x_101 & ~n_1956) ;
	assign n_1955 = (x_380 & x_718) ;
	assign n_1950 = (~n_1940 & ~n_1949) ;
	assign n_1939 = (~x_627 & ~n_1938) ;
	assign n_7647 = (~x_517 & n_7645) ;
	assign n_7646 = (x_517 & ~n_7645) ;
	assign n_7640 = (~x_516 & n_7638) ;
	assign n_7639 = (x_516 & ~n_7638) ;
	assign n_7632 = (~n_7628 & ~n_7631) ;
	assign n_7613 = (i_5 & ~n_7612) ;
	assign n_7611 = (~i_56 & n_936) ;
	assign n_7605 = (~n_7603 & ~n_7604) ;
	assign n_20 = (i_5 & ~n_17) ;
	assign n_18 = (i_5 & n_17) ;
	assign n_944 = (n_1 & n_3) ;
	assign n_286 = (x_130 & ~x_527) ;
	assign n_285 = (x_525 & x_527) ;
	assign n_7562 = (~x_669 & ~n_7560) ;
	assign n_1962 = (~n_1959 & n_1961) ;
	assign n_1958 = (~n_1955 & n_1957) ;
	assign n_1951 = (~n_1939 & ~n_1950) ;
	assign n_7648 = (~n_7646 & ~n_7647) ;
	assign n_7641 = (~n_7639 & ~n_7640) ;
	assign n_7634 = (~x_518 & n_7632) ;
	assign n_7633 = (x_518 & ~n_7632) ;
	assign n_7614 = (~n_7611 & n_7613) ;
	assign n_7606 = (n_20 & ~n_7605) ;
	assign n_7602 = (x_520 & n_18) ;
	assign n_948 = (n_3 & n_947) ;
	assign n_945 = (i_5 & ~n_944) ;
	assign n_544 = (x_697 & ~x_777) ;
	assign n_287 = (~n_285 & ~n_286) ;
	assign n_7563 = (~x_332 & ~n_7562) ;
	assign n_7561 = (x_669 & n_7560) ;
	assign n_2664 = (~x_718 & x_720) ;
	assign n_2660 = (x_492 & ~x_718) ;
	assign n_1963 = (~n_1958 & ~n_1962) ;
	assign n_1953 = (x_683 & n_1951) ;
	assign n_7649 = (~n_7641 & ~n_7648) ;
	assign n_7635 = (~n_7633 & ~n_7634) ;
	assign n_7616 = (~x_519 & ~n_7614) ;
	assign n_7615 = (x_519 & n_7614) ;
	assign n_7607 = (~n_7602 & ~n_7606) ;
	assign n_7597 = (i_11 & n_948) ;
	assign n_7596 = (x_521 & n_945) ;
	assign n_7590 = (~x_522 & ~n_544) ;
	assign n_7570 = (n_6 & n_287) ;
	assign n_7564 = (~n_7561 & n_7563) ;
	assign n_2665 = (~x_101 & ~n_2664) ;
	assign n_2663 = (x_718 & x_730) ;
	assign n_2661 = (x_101 & ~n_2660) ;
	assign n_2659 = (x_454 & x_718) ;
	assign n_2654 = (~n_1953 & ~n_1963) ;
	assign n_1952 = (~x_683 & ~n_1951) ;
	assign n_7650 = (~n_7635 & n_7649) ;
	assign n_7617 = (~n_7615 & ~n_7616) ;
	assign n_7609 = (~x_520 & n_7607) ;
	assign n_7608 = (x_520 & ~n_7607) ;
	assign n_7598 = (~n_7596 & ~n_7597) ;
	assign n_7591 = (i_5 & ~n_7590) ;
	assign n_7589 = (~i_62 & n_544) ;
	assign n_7583 = (~x_523 & ~n_936) ;
	assign n_7571 = (n_1 & ~n_7570) ;
	assign n_903 = (~i_61 & ~n_6) ;
	assign n_7566 = (n_287 & ~n_7564) ;
	assign n_2666 = (~n_2663 & n_2665) ;
	assign n_2662 = (~n_2659 & n_2661) ;
	assign n_2655 = (~n_1952 & ~n_2654) ;
	assign n_7651 = (~n_7617 & n_7650) ;
	assign n_7610 = (~n_7608 & ~n_7609) ;
	assign n_7600 = (~x_521 & n_7598) ;
	assign n_7599 = (x_521 & ~n_7598) ;
	assign n_7592 = (~n_7589 & n_7591) ;
	assign n_7584 = (i_5 & ~n_7583) ;
	assign n_7582 = (~i_23 & n_936) ;
	assign n_7572 = (~n_903 & n_7571) ;
	assign n_7569 = (n_59 & ~n_287) ;
	assign n_7567 = (x_664 & ~n_7566) ;
	assign n_7565 = (~n_287 & n_7564) ;
	assign n_7523 = (~x_691 & n_799) ;
	assign n_7522 = (x_691 & ~n_799) ;
	assign n_2808 = (~x_718 & x_790) ;
	assign n_2804 = (x_317 & ~x_718) ;
	assign n_2667 = (~n_2662 & ~n_2666) ;
	assign n_2657 = (x_600 & n_2655) ;
	assign n_7652 = (~n_7610 & n_7651) ;
	assign n_7601 = (~n_7599 & ~n_7600) ;
	assign n_7594 = (~x_522 & ~n_7592) ;
	assign n_7593 = (x_522 & n_7592) ;
	assign n_7585 = (~n_7582 & n_7584) ;
	assign n_7573 = (~n_7569 & ~n_7572) ;
	assign n_7568 = (~n_7565 & n_7567) ;
	assign n_697 = (~x_638 & x_777) ;
	assign n_7524 = (~n_7522 & ~n_7523) ;
	assign n_7521 = (~n_789 & ~n_790) ;
	assign n_2809 = (~x_101 & ~n_2808) ;
	assign n_2807 = (x_649 & x_718) ;
	assign n_2805 = (x_101 & ~n_2804) ;
	assign n_2803 = (x_369 & x_718) ;
	assign n_2799 = (~n_2657 & ~n_2667) ;
	assign n_2656 = (~x_600 & ~n_2655) ;
	assign n_7653 = (~n_7601 & n_7652) ;
	assign n_7595 = (~n_7593 & ~n_7594) ;
	assign n_7587 = (~x_523 & ~n_7585) ;
	assign n_7586 = (x_523 & n_7585) ;
	assign n_7574 = (~n_7568 & n_7573) ;
	assign n_7554 = (~x_526 & ~n_697) ;
	assign n_7533 = (i_8 & ~n_6) ;
	assign n_698 = (i_5 & ~n_697) ;
	assign n_669 = (n_629 & ~n_6) ;
	assign n_7526 = (n_7521 & ~n_7524) ;
	assign n_2810 = (~n_2807 & n_2809) ;
	assign n_2806 = (~n_2803 & n_2805) ;
	assign n_2800 = (~n_2656 & ~n_2799) ;
	assign n_7654 = (~n_7595 & n_7653) ;
	assign n_7588 = (~n_7586 & ~n_7587) ;
	assign n_7580 = (~x_524 & n_164) ;
	assign n_7579 = (x_524 & ~n_164) ;
	assign n_7575 = (i_5 & ~n_7574) ;
	assign n_7555 = (i_5 & ~n_7554) ;
	assign n_7553 = (~x_447 & n_697) ;
	assign n_7534 = (n_629 & ~n_7533) ;
	assign n_7532 = (x_529 & n_6) ;
	assign n_699 = (~n_669 & n_698) ;
	assign n_7529 = (x_529 & ~n_697) ;
	assign n_7527 = (n_697 & ~n_7526) ;
	assign n_7525 = (~n_7521 & n_7524) ;
	assign n_32 = (n_12 & ~n_14) ;
	assign n_30 = (x_332 & n_9) ;
	assign n_2821 = (~x_718 & x_791) ;
	assign n_2817 = (x_393 & ~x_718) ;
	assign n_2811 = (~n_2806 & ~n_2810) ;
	assign n_2802 = (x_216 & n_2800) ;
	assign n_7655 = (~n_7588 & n_7654) ;
	assign n_7581 = (~n_7579 & ~n_7580) ;
	assign n_7577 = (~x_525 & ~n_7575) ;
	assign n_7576 = (x_525 & n_7575) ;
	assign n_7556 = (~n_7553 & n_7555) ;
	assign n_4363 = (i_5 & ~n_7) ;
	assign n_7543 = (i_64 & n_59) ;
	assign n_7535 = (~n_7532 & n_7534) ;
	assign n_902 = (i_5 & ~n_699) ;
	assign n_7530 = (~n_629 & ~n_7529) ;
	assign n_7528 = (~n_7525 & n_7527) ;
	assign n_33 = (x_332 & n_32) ;
	assign n_31 = (n_8 & n_30) ;
	assign n_2822 = (~x_101 & ~n_2821) ;
	assign n_2820 = (x_568 & x_718) ;
	assign n_2818 = (x_101 & ~n_2817) ;
	assign n_2816 = (x_301 & x_718) ;
	assign n_2812 = (~n_2802 & ~n_2811) ;
	assign n_2801 = (~x_216 & ~n_2800) ;
	assign n_7656 = (~n_7581 & n_7655) ;
	assign n_7578 = (~n_7576 & ~n_7577) ;
	assign n_7558 = (~x_526 & ~n_7556) ;
	assign n_7557 = (x_526 & n_7556) ;
	assign n_7549 = (~n_527 & n_4363) ;
	assign n_7544 = (n_66 & n_7543) ;
	assign n_7542 = (x_528 & n_60) ;
	assign n_7536 = (n_902 & ~n_7535) ;
	assign n_7531 = (~n_7528 & n_7530) ;
	assign n_34 = (~n_31 & ~n_33) ;
	assign n_2834 = (~x_718 & x_719) ;
	assign n_2830 = (x_434 & ~x_718) ;
	assign n_2823 = (~n_2820 & n_2822) ;
	assign n_2819 = (~n_2816 & n_2818) ;
	assign n_2813 = (~n_2801 & ~n_2812) ;
	assign n_7657 = (~n_7578 & n_7656) ;
	assign n_7559 = (~n_7557 & ~n_7558) ;
	assign n_7551 = (~x_527 & n_7549) ;
	assign n_7550 = (x_527 & ~n_7549) ;
	assign n_7545 = (~n_7542 & ~n_7544) ;
	assign n_7537 = (~n_7531 & n_7536) ;
	assign n_7520 = (x_529 & n_699) ;
	assign n_7514 = (~x_530 & ~n_544) ;
	assign n_35 = (n_29 & ~n_34) ;
	assign n_3575 = (i_56 & ~n_6) ;
	assign n_7496 = (i_56 & n_1) ;
	assign n_2835 = (~x_101 & ~n_2834) ;
	assign n_2833 = (x_251 & x_718) ;
	assign n_2831 = (x_101 & ~n_2830) ;
	assign n_2829 = (x_514 & x_718) ;
	assign n_2824 = (~n_2819 & ~n_2823) ;
	assign n_2815 = (x_299 & n_2813) ;
	assign n_7658 = (~n_7559 & n_7657) ;
	assign n_7552 = (~n_7550 & ~n_7551) ;
	assign n_7547 = (~x_528 & n_7545) ;
	assign n_7546 = (x_528 & ~n_7545) ;
	assign n_7538 = (~n_7520 & ~n_7537) ;
	assign n_7515 = (i_5 & ~n_7514) ;
	assign n_7513 = (~i_15 & n_544) ;
	assign n_36 = (i_5 & ~n_35) ;
	assign n_7500 = (x_97 & ~n_16) ;
	assign n_7499 = (n_1 & n_3575) ;
	assign n_7497 = (~n_17 & ~n_7496) ;
	assign n_2836 = (~n_2833 & n_2835) ;
	assign n_2832 = (~n_2829 & n_2831) ;
	assign n_2825 = (~n_2815 & ~n_2824) ;
	assign n_2814 = (~x_299 & ~n_2813) ;
	assign n_7659 = (~n_7552 & n_7658) ;
	assign n_7548 = (~n_7546 & ~n_7547) ;
	assign n_7540 = (~x_529 & n_7538) ;
	assign n_7539 = (x_529 & ~n_7538) ;
	assign n_7516 = (~n_7513 & n_7515) ;
	assign n_7508 = (x_350 & n_35) ;
	assign n_7507 = (x_531 & n_36) ;
	assign n_7501 = (~n_7499 & ~n_7500) ;
	assign n_7498 = (x_532 & ~n_7497) ;
	assign n_2837 = (~n_2832 & ~n_2836) ;
	assign n_2826 = (~n_2814 & ~n_2825) ;
	assign n_7660 = (~n_7548 & n_7659) ;
	assign n_7541 = (~n_7539 & ~n_7540) ;
	assign n_7518 = (~x_530 & ~n_7516) ;
	assign n_7517 = (x_530 & n_7516) ;
	assign n_7509 = (~n_7507 & ~n_7508) ;
	assign n_7502 = (~n_7498 & n_7501) ;
	assign n_7446 = (~x_262 & n_2837) ;
	assign n_7445 = (x_262 & ~n_2837) ;
	assign n_2828 = (x_538 & n_2826) ;
	assign n_2827 = (~x_538 & ~n_2826) ;
	assign n_7661 = (~n_7541 & n_7660) ;
	assign n_7519 = (~n_7517 & ~n_7518) ;
	assign n_7511 = (~x_531 & n_7509) ;
	assign n_7510 = (x_531 & ~n_7509) ;
	assign n_7503 = (i_5 & ~n_7502) ;
	assign n_7491 = (i_28 & n_948) ;
	assign n_7490 = (x_533 & n_945) ;
	assign n_7447 = (~n_7445 & ~n_7446) ;
	assign n_7444 = (~n_2827 & ~n_2828) ;
	assign n_7662 = (~n_7519 & n_7661) ;
	assign n_7512 = (~n_7510 & ~n_7511) ;
	assign n_7505 = (~x_532 & ~n_7503) ;
	assign n_7504 = (x_532 & n_7503) ;
	assign n_7492 = (~n_7490 & ~n_7491) ;
	assign n_7485 = (x_432 & n_53) ;
	assign n_7484 = (x_534 & n_51) ;
	assign n_7478 = (i_24 & n_59) ;
	assign n_7455 = (~x_538 & n_6) ;
	assign n_6350 = (~i_13 & ~n_6) ;
	assign n_7449 = (n_7444 & ~n_7447) ;
	assign n_7663 = (~n_7512 & n_7662) ;
	assign n_7506 = (~n_7504 & ~n_7505) ;
	assign n_7494 = (~x_533 & n_7492) ;
	assign n_7493 = (x_533 & ~n_7492) ;
	assign n_7486 = (~n_7484 & ~n_7485) ;
	assign n_7479 = (n_66 & n_7478) ;
	assign n_7477 = (x_535 & n_60) ;
	assign n_7471 = (~x_536 & ~n_544) ;
	assign n_7456 = (~n_6350 & ~n_7455) ;
	assign n_7452 = (x_538 & ~n_697) ;
	assign n_7450 = (n_697 & ~n_7449) ;
	assign n_7448 = (~n_7444 & n_7447) ;
	assign n_7664 = (~n_7506 & n_7663) ;
	assign n_7495 = (~n_7493 & ~n_7494) ;
	assign n_7488 = (~x_534 & n_7486) ;
	assign n_7487 = (x_534 & ~n_7486) ;
	assign n_7480 = (~n_7477 & ~n_7479) ;
	assign n_7472 = (i_5 & ~n_7471) ;
	assign n_7470 = (~i_65 & n_544) ;
	assign n_7457 = (n_629 & ~n_7456) ;
	assign n_7453 = (~n_629 & ~n_7452) ;
	assign n_7451 = (~n_7448 & n_7450) ;
	assign n_7665 = (~n_7495 & n_7664) ;
	assign n_7489 = (~n_7487 & ~n_7488) ;
	assign n_7482 = (~x_535 & n_7480) ;
	assign n_7481 = (x_535 & ~n_7480) ;
	assign n_7473 = (~n_7470 & n_7472) ;
	assign n_7465 = (i_63 & n_948) ;
	assign n_7464 = (x_537 & n_945) ;
	assign n_7458 = (n_902 & ~n_7457) ;
	assign n_7454 = (~n_7451 & n_7453) ;
	assign n_7666 = (~n_7489 & n_7665) ;
	assign n_7483 = (~n_7481 & ~n_7482) ;
	assign n_7475 = (~x_536 & ~n_7473) ;
	assign n_7474 = (x_536 & n_7473) ;
	assign n_7466 = (~n_7464 & ~n_7465) ;
	assign n_7459 = (~n_7454 & n_7458) ;
	assign n_7443 = (x_538 & n_699) ;
	assign n_7437 = (~x_539 & ~n_697) ;
	assign n_291 = (x_71 & ~x_255) ;
	assign n_290 = (x_116 & ~x_578) ;
	assign n_7667 = (~n_7483 & n_7666) ;
	assign n_7476 = (~n_7474 & ~n_7475) ;
	assign n_7468 = (~x_537 & n_7466) ;
	assign n_7467 = (x_537 & ~n_7466) ;
	assign n_7460 = (~n_7443 & ~n_7459) ;
	assign n_7438 = (i_5 & ~n_7437) ;
	assign n_7436 = (~x_302 & n_697) ;
	assign n_1577 = (i_56 & n_59) ;
	assign n_630 = (n_63 & n_629) ;
	assign n_662 = (x_638 & n_49) ;
	assign n_295 = (x_554 & n_9) ;
	assign n_294 = (x_599 & n_13) ;
	assign n_292 = (~n_290 & ~n_291) ;
	assign n_7668 = (~n_7476 & n_7667) ;
	assign n_7469 = (~n_7467 & ~n_7468) ;
	assign n_7462 = (~x_538 & n_7460) ;
	assign n_7461 = (x_538 & ~n_7460) ;
	assign n_7439 = (~n_7436 & n_7438) ;
	assign n_1578 = (n_66 & n_1577) ;
	assign n_1576 = (x_540 & n_60) ;
	assign n_7427 = (~x_541 & ~n_630) ;
	assign n_7419 = (~i_27 & n_669) ;
	assign n_664 = (n_629 & n_6) ;
	assign n_663 = (~n_629 & ~n_662) ;
	assign n_296 = (~n_294 & ~n_295) ;
	assign n_293 = (~n_9 & ~n_292) ;
	assign n_288 = (~n_284 & ~n_287) ;
	assign n_7669 = (~n_7469 & n_7668) ;
	assign n_7463 = (~n_7461 & ~n_7462) ;
	assign n_7441 = (~x_539 & ~n_7439) ;
	assign n_7440 = (x_539 & n_7439) ;
	assign n_1579 = (~n_1576 & ~n_1578) ;
	assign n_7428 = (i_5 & ~n_7427) ;
	assign n_7426 = (~i_54 & n_630) ;
	assign n_7420 = (i_5 & ~n_7419) ;
	assign n_7418 = (~x_135 & n_662) ;
	assign n_665 = (~n_663 & ~n_664) ;
	assign n_306 = (x_167 & ~x_255) ;
	assign n_305 = (~x_578 & x_796) ;
	assign n_301 = (~x_527 & x_662) ;
	assign n_300 = (x_398 & x_527) ;
	assign n_297 = (~n_293 & n_296) ;
	assign n_289 = (~n_283 & ~n_288) ;
	assign n_7670 = (~n_7463 & n_7669) ;
	assign n_7442 = (~n_7440 & ~n_7441) ;
	assign n_7434 = (~x_540 & n_1579) ;
	assign n_7433 = (x_540 & ~n_1579) ;
	assign n_7429 = (~n_7426 & n_7428) ;
	assign n_7421 = (~n_7418 & n_7420) ;
	assign n_7417 = (~x_542 & ~n_665) ;
	assign n_7411 = (~x_543 & ~n_544) ;
	assign n_310 = (x_642 & n_9) ;
	assign n_309 = (x_517 & n_13) ;
	assign n_307 = (~n_305 & ~n_306) ;
	assign n_302 = (~n_300 & ~n_301) ;
	assign n_299 = (n_289 & n_297) ;
	assign n_7671 = (~n_7442 & n_7670) ;
	assign n_7435 = (~n_7433 & ~n_7434) ;
	assign n_7431 = (~x_541 & ~n_7429) ;
	assign n_7430 = (x_541 & n_7429) ;
	assign n_7422 = (~n_7417 & n_7421) ;
	assign n_7412 = (i_5 & ~n_7411) ;
	assign n_7410 = (~i_23 & n_544) ;
	assign n_7404 = (~x_544 & ~n_630) ;
	assign n_420 = (x_192 & ~x_527) ;
	assign n_419 = (x_84 & x_527) ;
	assign n_311 = (~n_309 & ~n_310) ;
	assign n_308 = (~n_9 & ~n_307) ;
	assign n_303 = (~n_299 & ~n_302) ;
	assign n_298 = (~n_289 & ~n_297) ;
	assign n_7672 = (~n_7435 & n_7671) ;
	assign n_7432 = (~n_7430 & ~n_7431) ;
	assign n_7424 = (~x_542 & ~n_7422) ;
	assign n_7423 = (x_542 & n_7422) ;
	assign n_7413 = (~n_7410 & n_7412) ;
	assign n_7405 = (i_5 & ~n_7404) ;
	assign n_7403 = (~i_16 & n_630) ;
	assign n_421 = (~n_419 & ~n_420) ;
	assign n_321 = (~x_255 & x_672) ;
	assign n_320 = (~x_578 & x_770) ;
	assign n_316 = (~x_527 & x_731) ;
	assign n_315 = (x_345 & x_527) ;
	assign n_312 = (~n_308 & n_311) ;
	assign n_304 = (~n_298 & ~n_303) ;
	assign n_7673 = (~n_7432 & n_7672) ;
	assign n_7425 = (~n_7423 & ~n_7424) ;
	assign n_7415 = (~x_543 & ~n_7413) ;
	assign n_7414 = (x_543 & n_7413) ;
	assign n_7406 = (~n_7403 & n_7405) ;
	assign n_7398 = (n_35 & ~n_421) ;
	assign n_7397 = (x_545 & n_36) ;
	assign n_325 = (x_195 & n_9) ;
	assign n_324 = (x_297 & n_13) ;
	assign n_322 = (~n_320 & ~n_321) ;
	assign n_317 = (~n_315 & ~n_316) ;
	assign n_314 = (n_304 & n_312) ;
	assign n_7674 = (~n_7425 & n_7673) ;
	assign n_7416 = (~n_7414 & ~n_7415) ;
	assign n_7408 = (~x_544 & ~n_7406) ;
	assign n_7407 = (x_544 & n_7406) ;
	assign n_7399 = (~n_7397 & ~n_7398) ;
	assign n_7392 = (~n_272 & n_35) ;
	assign n_7391 = (x_546 & n_36) ;
	assign n_1009 = (i_5 & n_527) ;
	assign n_1007 = (i_5 & ~n_527) ;
	assign n_7362 = (i_28 & ~n_6) ;
	assign n_326 = (~n_324 & ~n_325) ;
	assign n_323 = (~n_9 & ~n_322) ;
	assign n_318 = (~n_314 & ~n_317) ;
	assign n_313 = (~n_304 & ~n_312) ;
	assign n_7675 = (~n_7416 & n_7674) ;
	assign n_7409 = (~n_7407 & ~n_7408) ;
	assign n_7401 = (~x_545 & n_7399) ;
	assign n_7400 = (x_545 & ~n_7399) ;
	assign n_7393 = (~n_7391 & ~n_7392) ;
	assign n_7386 = (~n_242 & n_1009) ;
	assign n_7385 = (x_547 & n_1007) ;
	assign n_7379 = (i_45 & n_59) ;
	assign n_7363 = (n_629 & ~n_7362) ;
	assign n_7361 = (x_550 & n_6) ;
	assign n_336 = (x_86 & ~x_578) ;
	assign n_335 = (~x_255 & x_589) ;
	assign n_331 = (~x_527 & x_787) ;
	assign n_330 = (x_282 & x_527) ;
	assign n_327 = (~n_323 & n_326) ;
	assign n_319 = (~n_313 & ~n_318) ;
	assign n_7676 = (~n_7409 & n_7675) ;
	assign n_7402 = (~n_7400 & ~n_7401) ;
	assign n_7395 = (~x_546 & n_7393) ;
	assign n_7394 = (x_546 & ~n_7393) ;
	assign n_7387 = (~n_7385 & ~n_7386) ;
	assign n_7380 = (n_66 & n_7379) ;
	assign n_7378 = (x_548 & n_60) ;
	assign n_7372 = (~x_549 & ~n_544) ;
	assign n_7364 = (~n_7361 & n_7363) ;
	assign n_340 = (x_104 & n_9) ;
	assign n_339 = (x_373 & n_13) ;
	assign n_337 = (~n_335 & ~n_336) ;
	assign n_332 = (~n_330 & ~n_331) ;
	assign n_329 = (n_319 & n_327) ;
	assign n_7677 = (~n_7402 & n_7676) ;
	assign n_7396 = (~n_7394 & ~n_7395) ;
	assign n_7389 = (~x_547 & n_7387) ;
	assign n_7388 = (x_547 & ~n_7387) ;
	assign n_7381 = (~n_7378 & ~n_7380) ;
	assign n_7373 = (i_5 & ~n_7372) ;
	assign n_7371 = (~i_59 & n_544) ;
	assign n_7365 = (i_5 & ~n_7364) ;
	assign n_7360 = (~x_717 & n_662) ;
	assign n_341 = (~n_339 & ~n_340) ;
	assign n_338 = (~n_9 & ~n_337) ;
	assign n_333 = (~n_329 & ~n_332) ;
	assign n_328 = (~n_319 & ~n_327) ;
	assign n_7678 = (~n_7396 & n_7677) ;
	assign n_7390 = (~n_7388 & ~n_7389) ;
	assign n_7383 = (~x_548 & n_7381) ;
	assign n_7382 = (x_548 & ~n_7381) ;
	assign n_7374 = (~n_7371 & n_7373) ;
	assign n_7366 = (~n_7360 & n_7365) ;
	assign n_7359 = (~x_550 & n_663) ;
	assign n_7353 = (i_42 & n_64) ;
	assign n_978 = (i_5 & ~n_64) ;
	assign n_351 = (x_229 & ~x_255) ;
	assign n_350 = (~x_578 & x_742) ;
	assign n_346 = (x_92 & ~x_527) ;
	assign n_345 = (x_212 & x_527) ;
	assign n_342 = (~n_338 & n_341) ;
	assign n_334 = (~n_328 & ~n_333) ;
	assign n_7679 = (~n_7390 & n_7678) ;
	assign n_7384 = (~n_7382 & ~n_7383) ;
	assign n_7376 = (~x_549 & ~n_7374) ;
	assign n_7375 = (x_549 & n_7374) ;
	assign n_7367 = (~n_7359 & n_7366) ;
	assign n_7354 = (n_66 & n_7353) ;
	assign n_7352 = (x_551 & n_978) ;
	assign n_355 = (x_705 & n_9) ;
	assign n_354 = (x_443 & n_13) ;
	assign n_352 = (~n_350 & ~n_351) ;
	assign n_347 = (~n_345 & ~n_346) ;
	assign n_344 = (n_334 & n_342) ;
	assign n_7680 = (~n_7384 & n_7679) ;
	assign n_7377 = (~n_7375 & ~n_7376) ;
	assign n_7369 = (~x_550 & ~n_7367) ;
	assign n_7368 = (x_550 & n_7367) ;
	assign n_7355 = (~n_7352 & ~n_7354) ;
	assign n_7347 = (~n_143 & n_35) ;
	assign n_7346 = (x_552 & n_36) ;
	assign n_356 = (~n_354 & ~n_355) ;
	assign n_353 = (~n_9 & ~n_352) ;
	assign n_348 = (~n_344 & ~n_347) ;
	assign n_343 = (~n_334 & ~n_342) ;
	assign n_7681 = (~n_7377 & n_7680) ;
	assign n_7370 = (~n_7368 & ~n_7369) ;
	assign n_7357 = (~x_551 & n_7355) ;
	assign n_7356 = (x_551 & ~n_7355) ;
	assign n_7348 = (~n_7346 & ~n_7347) ;
	assign n_406 = (~x_527 & x_553) ;
	assign n_405 = (x_527 & x_784) ;
	assign n_7337 = (i_60 & n_64) ;
	assign n_366 = (x_176 & ~x_255) ;
	assign n_365 = (~x_578 & x_786) ;
	assign n_361 = (x_160 & ~x_527) ;
	assign n_360 = (x_138 & x_527) ;
	assign n_357 = (~n_353 & n_356) ;
	assign n_349 = (~n_343 & ~n_348) ;
	assign n_7682 = (~n_7370 & n_7681) ;
	assign n_7358 = (~n_7356 & ~n_7357) ;
	assign n_7350 = (~x_552 & n_7348) ;
	assign n_7349 = (x_552 & ~n_7348) ;
	assign n_407 = (~n_405 & ~n_406) ;
	assign n_7338 = (n_66 & n_7337) ;
	assign n_7336 = (x_554 & n_978) ;
	assign n_7330 = (~x_555 & ~n_630) ;
	assign n_370 = (x_653 & n_9) ;
	assign n_369 = (x_399 & n_13) ;
	assign n_367 = (~n_365 & ~n_366) ;
	assign n_362 = (~n_360 & ~n_361) ;
	assign n_359 = (n_349 & n_357) ;
	assign n_7683 = (~n_7358 & n_7682) ;
	assign n_7351 = (~n_7349 & ~n_7350) ;
	assign n_7344 = (~x_553 & n_407) ;
	assign n_7343 = (x_553 & ~n_407) ;
	assign n_7339 = (~n_7336 & ~n_7338) ;
	assign n_7331 = (i_5 & ~n_7330) ;
	assign n_7329 = (~i_26 & n_630) ;
	assign n_435 = (x_122 & ~x_527) ;
	assign n_434 = (x_155 & x_527) ;
	assign n_371 = (~n_369 & ~n_370) ;
	assign n_368 = (~n_9 & ~n_367) ;
	assign n_363 = (~n_359 & ~n_362) ;
	assign n_358 = (~n_349 & ~n_357) ;
	assign n_7684 = (~n_7351 & n_7683) ;
	assign n_7345 = (~n_7343 & ~n_7344) ;
	assign n_7341 = (~x_554 & n_7339) ;
	assign n_7340 = (x_554 & ~n_7339) ;
	assign n_7332 = (~n_7329 & n_7331) ;
	assign n_7324 = (~n_227 & n_35) ;
	assign n_7323 = (x_556 & n_36) ;
	assign n_436 = (~n_434 & ~n_435) ;
	assign n_381 = (~x_255 & x_256) ;
	assign n_380 = (~x_578 & x_716) ;
	assign n_372 = (~n_368 & n_371) ;
	assign n_364 = (~n_358 & ~n_363) ;
	assign n_375 = (x_228 & ~x_527) ;
	assign n_374 = (x_76 & x_527) ;
	assign n_7685 = (~n_7345 & n_7684) ;
	assign n_7342 = (~n_7340 & ~n_7341) ;
	assign n_7334 = (~x_555 & ~n_7332) ;
	assign n_7333 = (x_555 & n_7332) ;
	assign n_7325 = (~n_7323 & ~n_7324) ;
	assign n_7318 = (n_1009 & ~n_436) ;
	assign n_7317 = (x_557 & n_1007) ;
	assign n_7311 = (~x_558 & ~n_697) ;
	assign n_385 = (x_734 & n_9) ;
	assign n_384 = (x_430 & n_13) ;
	assign n_382 = (~n_380 & ~n_381) ;
	assign n_377 = (n_364 & n_372) ;
	assign n_376 = (~n_374 & ~n_375) ;
	assign n_7686 = (~n_7342 & n_7685) ;
	assign n_7335 = (~n_7333 & ~n_7334) ;
	assign n_7327 = (~x_556 & n_7325) ;
	assign n_7326 = (x_556 & ~n_7325) ;
	assign n_7319 = (~n_7317 & ~n_7318) ;
	assign n_7312 = (i_5 & ~n_7311) ;
	assign n_7310 = (~x_806 & n_697) ;
	assign n_7304 = (i_16 & n_64) ;
	assign n_386 = (~n_384 & ~n_385) ;
	assign n_383 = (~n_9 & ~n_382) ;
	assign n_378 = (~n_376 & ~n_377) ;
	assign n_373 = (~n_364 & ~n_372) ;
	assign n_7687 = (~n_7335 & n_7686) ;
	assign n_7328 = (~n_7326 & ~n_7327) ;
	assign n_7321 = (~x_557 & n_7319) ;
	assign n_7320 = (x_557 & ~n_7319) ;
	assign n_7313 = (~n_7310 & n_7312) ;
	assign n_7305 = (n_66 & n_7304) ;
	assign n_7303 = (x_559 & n_978) ;
	assign n_7297 = (~x_560 & ~n_936) ;
	assign n_396 = (~x_255 & x_336) ;
	assign n_395 = (~x_578 & x_632) ;
	assign n_391 = (x_293 & ~x_527) ;
	assign n_390 = (x_527 & x_724) ;
	assign n_387 = (~n_383 & n_386) ;
	assign n_379 = (~n_373 & ~n_378) ;
	assign n_7688 = (~n_7328 & n_7687) ;
	assign n_7322 = (~n_7320 & ~n_7321) ;
	assign n_7315 = (~x_558 & ~n_7313) ;
	assign n_7314 = (x_558 & n_7313) ;
	assign n_7306 = (~n_7303 & ~n_7305) ;
	assign n_7298 = (i_5 & ~n_7297) ;
	assign n_7296 = (~i_47 & n_936) ;
	assign n_7290 = (i_23 & n_59) ;
	assign n_400 = (x_95 & n_9) ;
	assign n_399 = (x_353 & n_13) ;
	assign n_397 = (~n_395 & ~n_396) ;
	assign n_392 = (~n_390 & ~n_391) ;
	assign n_389 = (n_379 & n_387) ;
	assign n_7689 = (~n_7322 & n_7688) ;
	assign n_7316 = (~n_7314 & ~n_7315) ;
	assign n_7308 = (~x_559 & n_7306) ;
	assign n_7307 = (x_559 & ~n_7306) ;
	assign n_7299 = (~n_7296 & n_7298) ;
	assign n_7291 = (n_66 & n_7290) ;
	assign n_7289 = (x_561 & n_60) ;
	assign n_7283 = (~x_562 & ~n_936) ;
	assign n_401 = (~n_399 & ~n_400) ;
	assign n_398 = (~n_9 & ~n_397) ;
	assign n_393 = (~n_389 & ~n_392) ;
	assign n_388 = (~n_379 & ~n_387) ;
	assign n_7690 = (~n_7316 & n_7689) ;
	assign n_7309 = (~n_7307 & ~n_7308) ;
	assign n_7301 = (~x_560 & ~n_7299) ;
	assign n_7300 = (x_560 & n_7299) ;
	assign n_7292 = (~n_7289 & ~n_7291) ;
	assign n_7284 = (i_5 & ~n_7283) ;
	assign n_7282 = (~i_31 & n_936) ;
	assign n_7276 = (i_28 & n_64) ;
	assign n_411 = (x_185 & ~x_578) ;
	assign n_410 = (~x_255 & x_490) ;
	assign n_402 = (~n_398 & n_401) ;
	assign n_394 = (~n_388 & ~n_393) ;
	assign n_7691 = (~n_7309 & n_7690) ;
	assign n_7302 = (~n_7300 & ~n_7301) ;
	assign n_7294 = (~x_561 & n_7292) ;
	assign n_7293 = (x_561 & ~n_7292) ;
	assign n_7285 = (~n_7282 & n_7284) ;
	assign n_7277 = (n_66 & n_7276) ;
	assign n_7275 = (x_563 & n_978) ;
	assign n_7269 = (i_68 & n_64) ;
	assign n_415 = (x_780 & n_9) ;
	assign n_414 = (x_453 & n_13) ;
	assign n_412 = (~n_410 & ~n_411) ;
	assign n_404 = (n_394 & n_402) ;
	assign n_7692 = (~n_7302 & n_7691) ;
	assign n_7295 = (~n_7293 & ~n_7294) ;
	assign n_7287 = (~x_562 & ~n_7285) ;
	assign n_7286 = (x_562 & n_7285) ;
	assign n_7278 = (~n_7275 & ~n_7277) ;
	assign n_7270 = (n_66 & n_7269) ;
	assign n_7268 = (x_564 & n_978) ;
	assign n_416 = (~n_414 & ~n_415) ;
	assign n_413 = (~n_9 & ~n_412) ;
	assign n_408 = (~n_404 & ~n_407) ;
	assign n_403 = (~n_394 & ~n_402) ;
	assign n_7693 = (~n_7295 & n_7692) ;
	assign n_7288 = (~n_7286 & ~n_7287) ;
	assign n_7280 = (~x_563 & n_7278) ;
	assign n_7279 = (x_563 & ~n_7278) ;
	assign n_7271 = (~n_7268 & ~n_7270) ;
	assign n_426 = (x_269 & ~x_578) ;
	assign n_425 = (~x_255 & x_417) ;
	assign n_417 = (~n_413 & n_416) ;
	assign n_409 = (~n_403 & ~n_408) ;
	assign n_7694 = (~n_7288 & n_7693) ;
	assign n_7281 = (~n_7279 & ~n_7280) ;
	assign n_7273 = (~x_564 & n_7271) ;
	assign n_7272 = (x_564 & ~n_7271) ;
	assign n_7260 = (x_613 & n_53) ;
	assign n_7259 = (x_566 & n_51) ;
	assign n_7253 = (~x_567 & ~n_697) ;
	assign n_430 = (x_701 & n_9) ;
	assign n_429 = (x_535 & n_13) ;
	assign n_427 = (~n_425 & ~n_426) ;
	assign n_422 = (n_409 & n_417) ;
	assign n_7695 = (~n_7281 & n_7694) ;
	assign n_7274 = (~n_7272 & ~n_7273) ;
	assign n_7266 = (~x_565 & n_257) ;
	assign n_7265 = (x_565 & ~n_257) ;
	assign n_7261 = (~n_7259 & ~n_7260) ;
	assign n_7254 = (i_5 & ~n_7253) ;
	assign n_7252 = (~x_323 & n_697) ;
	assign n_7246 = (~x_568 & ~n_630) ;
	assign n_431 = (~n_429 & ~n_430) ;
	assign n_428 = (~n_9 & ~n_427) ;
	assign n_423 = (~n_421 & ~n_422) ;
	assign n_418 = (~n_409 & ~n_417) ;
	assign n_7696 = (~n_7274 & n_7695) ;
	assign n_7267 = (~n_7265 & ~n_7266) ;
	assign n_7263 = (~x_566 & n_7261) ;
	assign n_7262 = (x_566 & ~n_7261) ;
	assign n_7255 = (~n_7252 & n_7254) ;
	assign n_7247 = (i_5 & ~n_7246) ;
	assign n_7245 = (~i_21 & n_630) ;
	assign n_441 = (~x_255 & x_390) ;
	assign n_440 = (x_563 & ~x_578) ;
	assign n_432 = (~n_428 & n_431) ;
	assign n_424 = (~n_418 & ~n_423) ;
	assign n_7697 = (~n_7267 & n_7696) ;
	assign n_7264 = (~n_7262 & ~n_7263) ;
	assign n_7257 = (~x_567 & ~n_7255) ;
	assign n_7256 = (x_567 & n_7255) ;
	assign n_7248 = (~n_7245 & n_7247) ;
	assign n_7240 = (~n_164 & n_1009) ;
	assign n_7239 = (x_569 & n_1007) ;
	assign n_7233 = (~x_570 & ~n_630) ;
	assign n_7225 = (~i_6 & n_669) ;
	assign n_445 = (x_105 & n_9) ;
	assign n_444 = (x_296 & n_13) ;
	assign n_442 = (~n_440 & ~n_441) ;
	assign n_437 = (n_424 & n_432) ;
	assign n_7698 = (~n_7264 & n_7697) ;
	assign n_7258 = (~n_7256 & ~n_7257) ;
	assign n_7250 = (~x_568 & ~n_7248) ;
	assign n_7249 = (x_568 & n_7248) ;
	assign n_7241 = (~n_7239 & ~n_7240) ;
	assign n_7234 = (i_5 & ~n_7233) ;
	assign n_7232 = (~i_42 & n_630) ;
	assign n_7226 = (i_5 & ~n_7225) ;
	assign n_7224 = (~x_558 & n_662) ;
	assign n_7180 = (~x_576 & ~n_709) ;
	assign n_446 = (~n_444 & ~n_445) ;
	assign n_443 = (~n_9 & ~n_442) ;
	assign n_438 = (~n_436 & ~n_437) ;
	assign n_433 = (~n_424 & ~n_432) ;
	assign n_7699 = (~n_7258 & n_7698) ;
	assign n_7251 = (~n_7249 & ~n_7250) ;
	assign n_7243 = (~x_569 & n_7241) ;
	assign n_7242 = (x_569 & ~n_7241) ;
	assign n_7235 = (~n_7232 & n_7234) ;
	assign n_7227 = (~n_7224 & n_7226) ;
	assign n_7223 = (~x_571 & ~n_665) ;
	assign n_7181 = (~n_710 & ~n_7180) ;
	assign n_456 = (~x_255 & x_470) ;
	assign n_455 = (x_479 & ~x_578) ;
	assign n_451 = (~x_527 & x_814) ;
	assign n_450 = (x_510 & x_527) ;
	assign n_447 = (~n_443 & n_446) ;
	assign n_439 = (~n_433 & ~n_438) ;
	assign n_7700 = (~n_7251 & n_7699) ;
	assign n_7244 = (~n_7242 & ~n_7243) ;
	assign n_7237 = (~x_570 & ~n_7235) ;
	assign n_7236 = (x_570 & n_7235) ;
	assign n_7228 = (~n_7223 & n_7227) ;
	assign n_7218 = (x_717 & n_53) ;
	assign n_7217 = (x_572 & n_51) ;
	assign n_4905 = (i_49 & ~n_6) ;
	assign n_7183 = (x_423 & n_7181) ;
	assign n_1558 = (x_168 & x_255) ;
	assign n_1538 = (x_332 & x_664) ;
	assign n_460 = (x_200 & n_9) ;
	assign n_459 = (x_215 & n_13) ;
	assign n_457 = (~n_455 & ~n_456) ;
	assign n_452 = (~n_450 & ~n_451) ;
	assign n_449 = (n_439 & n_447) ;
	assign n_7701 = (~n_7244 & n_7700) ;
	assign n_7238 = (~n_7236 & ~n_7237) ;
	assign n_7230 = (~x_571 & ~n_7228) ;
	assign n_7229 = (x_571 & n_7228) ;
	assign n_7219 = (~n_7217 & ~n_7218) ;
	assign n_7212 = (x_631 & n_35) ;
	assign n_7211 = (x_573 & n_36) ;
	assign n_7205 = (~x_574 & ~n_936) ;
	assign n_7190 = (n_629 & ~n_4905) ;
	assign n_7189 = (x_576 & n_6) ;
	assign n_7186 = (x_576 & ~n_697) ;
	assign n_7184 = (n_697 & ~n_7183) ;
	assign n_7182 = (~x_423 & ~n_7181) ;
	assign n_1559 = (n_1538 & ~n_1558) ;
	assign n_461 = (~n_459 & ~n_460) ;
	assign n_458 = (~n_9 & ~n_457) ;
	assign n_453 = (~n_449 & ~n_452) ;
	assign n_448 = (~n_439 & ~n_447) ;
	assign n_7702 = (~n_7238 & n_7701) ;
	assign n_7231 = (~n_7229 & ~n_7230) ;
	assign n_7221 = (~x_572 & n_7219) ;
	assign n_7220 = (x_572 & ~n_7219) ;
	assign n_7213 = (~n_7211 & ~n_7212) ;
	assign n_7206 = (i_5 & ~n_7205) ;
	assign n_7204 = (~i_61 & n_936) ;
	assign n_7191 = (~n_7189 & n_7190) ;
	assign n_7187 = (~n_629 & ~n_7186) ;
	assign n_7185 = (~n_7182 & n_7184) ;
	assign n_1560 = (x_578 & ~n_1559) ;
	assign n_1557 = (~x_168 & n_10) ;
	assign n_462 = (~n_458 & n_461) ;
	assign n_454 = (~n_448 & ~n_453) ;
	assign n_7703 = (~n_7231 & n_7702) ;
	assign n_7222 = (~n_7220 & ~n_7221) ;
	assign n_7215 = (~x_573 & n_7213) ;
	assign n_7214 = (x_573 & ~n_7213) ;
	assign n_7207 = (~n_7204 & n_7206) ;
	assign n_7199 = (i_36 & n_948) ;
	assign n_7198 = (x_575 & n_945) ;
	assign n_7192 = (n_902 & ~n_7191) ;
	assign n_7188 = (~n_7185 & n_7187) ;
	assign n_1563 = (~x_578 & ~n_3) ;
	assign n_1542 = (n_1 & ~n_5) ;
	assign n_1561 = (~n_1557 & ~n_1560) ;
	assign n_464 = (n_454 & n_462) ;
	assign n_463 = (~n_454 & ~n_462) ;
	assign n_7704 = (~n_7222 & n_7703) ;
	assign n_7216 = (~n_7214 & ~n_7215) ;
	assign n_7209 = (~x_574 & ~n_7207) ;
	assign n_7208 = (x_574 & n_7207) ;
	assign n_7200 = (~n_7198 & ~n_7199) ;
	assign n_7193 = (~n_7188 & n_7192) ;
	assign n_7179 = (x_576 & n_699) ;
	assign n_7173 = (~x_577 & ~n_544) ;
	assign n_1564 = (n_1542 & ~n_1563) ;
	assign n_1562 = (~n_1 & ~n_1561) ;
	assign n_7134 = (~n_463 & ~n_464) ;
	assign n_7705 = (~n_7216 & n_7704) ;
	assign n_7210 = (~n_7208 & ~n_7209) ;
	assign n_7202 = (~x_575 & n_7200) ;
	assign n_7201 = (x_575 & ~n_7200) ;
	assign n_7194 = (~n_7179 & ~n_7193) ;
	assign n_7174 = (i_5 & ~n_7173) ;
	assign n_7172 = (~i_39 & n_544) ;
	assign n_1565 = (~n_1562 & ~n_1564) ;
	assign n_466 = (~x_527 & x_763) ;
	assign n_465 = (x_527 & x_582) ;
	assign n_7136 = (~x_520 & ~n_7134) ;
	assign n_7706 = (~n_7210 & n_7705) ;
	assign n_7203 = (~n_7201 & ~n_7202) ;
	assign n_7196 = (~x_576 & n_7194) ;
	assign n_7195 = (x_576 & ~n_7194) ;
	assign n_7175 = (~n_7172 & n_7174) ;
	assign n_1567 = (x_578 & n_18) ;
	assign n_1566 = (n_20 & ~n_1565) ;
	assign n_467 = (~n_465 & ~n_466) ;
	assign n_7137 = (n_527 & ~n_7136) ;
	assign n_7135 = (x_520 & n_7134) ;
	assign n_7707 = (~n_7203 & n_7706) ;
	assign n_7197 = (~n_7195 & ~n_7196) ;
	assign n_7177 = (~x_577 & ~n_7175) ;
	assign n_7176 = (x_577 & n_7175) ;
	assign n_1568 = (~n_1566 & ~n_1567) ;
	assign n_7164 = (x_458 & n_53) ;
	assign n_7163 = (x_579 & n_51) ;
	assign n_3935 = (i_5 & n_936) ;
	assign n_3933 = (i_5 & ~n_936) ;
	assign n_7143 = (n_6 & n_467) ;
	assign n_3966 = (~i_14 & ~n_6) ;
	assign n_7138 = (~n_7135 & n_7137) ;
	assign n_7093 = (~n_214 & ~n_215) ;
	assign n_7708 = (~n_7197 & n_7707) ;
	assign n_7178 = (~n_7176 & ~n_7177) ;
	assign n_7170 = (~x_578 & n_1568) ;
	assign n_7169 = (x_578 & ~n_1568) ;
	assign n_7165 = (~n_7163 & ~n_7164) ;
	assign n_7158 = (i_40 & n_3935) ;
	assign n_7157 = (x_580 & n_3933) ;
	assign n_7144 = (~n_3966 & ~n_7143) ;
	assign n_7140 = (n_467 & n_7138) ;
	assign n_7095 = (~x_670 & ~n_7093) ;
	assign n_7709 = (~n_7178 & n_7708) ;
	assign n_7171 = (~n_7169 & ~n_7170) ;
	assign n_7167 = (~x_579 & n_7165) ;
	assign n_7166 = (x_579 & ~n_7165) ;
	assign n_7159 = (~n_7157 & ~n_7158) ;
	assign n_7152 = (x_429 & n_35) ;
	assign n_7151 = (x_581 & n_36) ;
	assign n_7145 = (n_1 & ~n_7144) ;
	assign n_7141 = (~n_1 & ~n_7140) ;
	assign n_7139 = (~n_467 & ~n_7138) ;
	assign n_7127 = (x_202 & ~n_16) ;
	assign n_7126 = (i_40 & n_7) ;
	assign n_7096 = (~x_332 & ~n_7095) ;
	assign n_7094 = (x_670 & n_7093) ;
	assign n_7710 = (~n_7171 & n_7709) ;
	assign n_7168 = (~n_7166 & ~n_7167) ;
	assign n_7161 = (~x_580 & n_7159) ;
	assign n_7160 = (x_580 & ~n_7159) ;
	assign n_7153 = (~n_7151 & ~n_7152) ;
	assign n_7146 = (i_5 & ~n_7145) ;
	assign n_7142 = (~n_7139 & n_7141) ;
	assign n_7128 = (~n_7126 & ~n_7127) ;
	assign n_4639 = (~i_53 & ~n_6) ;
	assign n_7097 = (~n_7094 & n_7096) ;
	assign n_7711 = (~n_7168 & n_7710) ;
	assign n_7162 = (~n_7160 & ~n_7161) ;
	assign n_7155 = (~x_581 & n_7153) ;
	assign n_7154 = (x_581 & ~n_7153) ;
	assign n_7147 = (~n_7142 & n_7146) ;
	assign n_7129 = (n_20 & ~n_7128) ;
	assign n_7125 = (x_583 & n_18) ;
	assign n_7104 = (n_1 & ~n_4639) ;
	assign n_7103 = (n_6 & n_218) ;
	assign n_7099 = (n_218 & ~n_7097) ;
	assign n_7712 = (~n_7162 & n_7711) ;
	assign n_7156 = (~n_7154 & ~n_7155) ;
	assign n_7149 = (~x_582 & ~n_7147) ;
	assign n_7148 = (x_582 & n_7147) ;
	assign n_7130 = (~n_7125 & ~n_7129) ;
	assign n_7120 = (i_61 & n_948) ;
	assign n_7119 = (x_584 & n_945) ;
	assign n_7113 = (~x_585 & ~n_936) ;
	assign n_7105 = (~n_7103 & n_7104) ;
	assign n_7102 = (n_59 & ~n_218) ;
	assign n_7100 = (x_664 & ~n_7099) ;
	assign n_7098 = (~n_218 & n_7097) ;
	assign n_7713 = (~n_7156 & n_7712) ;
	assign n_7150 = (~n_7148 & ~n_7149) ;
	assign n_7132 = (~x_583 & n_7130) ;
	assign n_7131 = (x_583 & ~n_7130) ;
	assign n_7121 = (~n_7119 & ~n_7120) ;
	assign n_7114 = (i_5 & ~n_7113) ;
	assign n_7112 = (~i_36 & n_936) ;
	assign n_7106 = (~n_7102 & ~n_7105) ;
	assign n_7101 = (~n_7098 & n_7100) ;
	assign n_7714 = (~n_7150 & n_7713) ;
	assign n_7133 = (~n_7131 & ~n_7132) ;
	assign n_7123 = (~x_584 & n_7121) ;
	assign n_7122 = (x_584 & ~n_7121) ;
	assign n_7115 = (~n_7112 & n_7114) ;
	assign n_7107 = (~n_7101 & n_7106) ;
	assign n_7715 = (~n_7133 & n_7714) ;
	assign n_7124 = (~n_7122 & ~n_7123) ;
	assign n_7117 = (~x_585 & ~n_7115) ;
	assign n_7116 = (x_585 & n_7115) ;
	assign n_7108 = (i_5 & ~n_7107) ;
	assign n_7088 = (x_370 & n_53) ;
	assign n_7087 = (x_587 & n_51) ;
	assign n_7081 = (~x_588 & ~n_936) ;
	assign n_7716 = (~n_7124 & n_7715) ;
	assign n_7118 = (~n_7116 & ~n_7117) ;
	assign n_7110 = (~x_586 & ~n_7108) ;
	assign n_7109 = (x_586 & n_7108) ;
	assign n_7089 = (~n_7087 & ~n_7088) ;
	assign n_7082 = (i_5 & ~n_7081) ;
	assign n_7080 = (~i_9 & n_936) ;
	assign n_7074 = (i_36 & n_59) ;
	assign n_7717 = (~n_7118 & n_7716) ;
	assign n_7111 = (~n_7109 & ~n_7110) ;
	assign n_7091 = (~x_587 & n_7089) ;
	assign n_7090 = (x_587 & ~n_7089) ;
	assign n_7083 = (~n_7080 & n_7082) ;
	assign n_7075 = (n_66 & n_7074) ;
	assign n_7073 = (x_589 & n_60) ;
	assign n_7067 = (~x_590 & ~n_630) ;
	assign n_7718 = (~n_7111 & n_7717) ;
	assign n_7092 = (~n_7090 & ~n_7091) ;
	assign n_7085 = (~x_588 & ~n_7083) ;
	assign n_7084 = (x_588 & n_7083) ;
	assign n_7076 = (~n_7073 & ~n_7075) ;
	assign n_7068 = (i_5 & ~n_7067) ;
	assign n_7066 = (~i_59 & n_630) ;
	assign n_7719 = (~n_7092 & n_7718) ;
	assign n_7086 = (~n_7084 & ~n_7085) ;
	assign n_7078 = (~x_589 & n_7076) ;
	assign n_7077 = (x_589 & ~n_7076) ;
	assign n_7069 = (~n_7066 & n_7068) ;
	assign n_7720 = (~n_7086 & n_7719) ;
	assign n_7079 = (~n_7077 & ~n_7078) ;
	assign n_7071 = (~x_590 & ~n_7069) ;
	assign n_7070 = (x_590 & n_7069) ;
	assign n_7058 = (x_352 & n_35) ;
	assign n_7057 = (x_592 & n_36) ;
	assign n_7051 = (i_45 & n_64) ;
	assign n_7721 = (~n_7079 & n_7720) ;
	assign n_7072 = (~n_7070 & ~n_7071) ;
	assign n_7064 = (~x_591 & n_179) ;
	assign n_7063 = (x_591 & ~n_179) ;
	assign n_7059 = (~n_7057 & ~n_7058) ;
	assign n_7052 = (n_66 & n_7051) ;
	assign n_7050 = (x_593 & n_978) ;
	assign n_7722 = (~n_7072 & n_7721) ;
	assign n_7065 = (~n_7063 & ~n_7064) ;
	assign n_7061 = (~x_592 & n_7059) ;
	assign n_7060 = (x_592 & ~n_7059) ;
	assign n_7053 = (~n_7050 & ~n_7052) ;
	assign n_7045 = (i_16 & n_948) ;
	assign n_7044 = (x_594 & n_945) ;
	assign n_7038 = (i_11 & n_64) ;
	assign n_7723 = (~n_7065 & n_7722) ;
	assign n_7062 = (~n_7060 & ~n_7061) ;
	assign n_7055 = (~x_593 & n_7053) ;
	assign n_7054 = (x_593 & ~n_7053) ;
	assign n_7046 = (~n_7044 & ~n_7045) ;
	assign n_7039 = (n_66 & n_7038) ;
	assign n_7037 = (x_595 & n_978) ;
	assign n_7724 = (~n_7062 & n_7723) ;
	assign n_7056 = (~n_7054 & ~n_7055) ;
	assign n_7048 = (~x_594 & n_7046) ;
	assign n_7047 = (x_594 & ~n_7046) ;
	assign n_7040 = (~n_7037 & ~n_7039) ;
	assign n_7032 = (i_47 & n_948) ;
	assign n_7031 = (x_596 & n_945) ;
	assign n_7025 = (~x_597 & ~n_544) ;
	assign n_7725 = (~n_7056 & n_7724) ;
	assign n_7049 = (~n_7047 & ~n_7048) ;
	assign n_7042 = (~x_595 & n_7040) ;
	assign n_7041 = (x_595 & ~n_7040) ;
	assign n_7033 = (~n_7031 & ~n_7032) ;
	assign n_7026 = (i_5 & ~n_7025) ;
	assign n_7024 = (~i_28 & n_544) ;
	assign n_7018 = (i_38 & n_59) ;
	assign n_7726 = (~n_7049 & n_7725) ;
	assign n_7043 = (~n_7041 & ~n_7042) ;
	assign n_7035 = (~x_596 & n_7033) ;
	assign n_7034 = (x_596 & ~n_7033) ;
	assign n_7027 = (~n_7024 & n_7026) ;
	assign n_7019 = (n_66 & n_7018) ;
	assign n_7017 = (x_598 & n_60) ;
	assign n_7011 = (~x_69 & ~n_630) ;
	assign n_7727 = (~n_7043 & n_7726) ;
	assign n_7036 = (~n_7034 & ~n_7035) ;
	assign n_7029 = (~x_597 & ~n_7027) ;
	assign n_7028 = (x_597 & n_7027) ;
	assign n_7020 = (~n_7017 & ~n_7019) ;
	assign n_7012 = (i_5 & ~n_7011) ;
	assign n_7010 = (~i_25 & n_630) ;
	assign n_7004 = (~x_70 & ~n_697) ;
	assign n_6951 = (~n_377 & ~n_373) ;
	assign n_7728 = (~n_7036 & n_7727) ;
	assign n_7030 = (~n_7028 & ~n_7029) ;
	assign n_7022 = (~x_598 & n_7020) ;
	assign n_7021 = (x_598 & ~n_7020) ;
	assign n_7013 = (~n_7010 & n_7012) ;
	assign n_7005 = (i_5 & ~n_7004) ;
	assign n_7003 = (~x_576 & n_697) ;
	assign n_6997 = (i_60 & n_59) ;
	assign n_6953 = (~x_823 & ~n_6951) ;
	assign n_7729 = (~n_7030 & n_7728) ;
	assign n_7023 = (~n_7021 & ~n_7022) ;
	assign n_7015 = (~x_69 & ~n_7013) ;
	assign n_7014 = (x_69 & n_7013) ;
	assign n_7006 = (~n_7003 & n_7005) ;
	assign n_6998 = (n_66 & n_6997) ;
	assign n_6996 = (x_71 & n_60) ;
	assign n_6954 = (~x_332 & ~n_6953) ;
	assign n_6952 = (x_823 & n_6951) ;
	assign n_7730 = (~n_7023 & n_7729) ;
	assign n_7016 = (~n_7014 & ~n_7015) ;
	assign n_7008 = (~x_70 & ~n_7006) ;
	assign n_7007 = (x_70 & n_7006) ;
	assign n_6999 = (~n_6996 & ~n_6998) ;
	assign n_6991 = (x_504 & n_53) ;
	assign n_6990 = (x_72 & n_51) ;
	assign n_6984 = (~x_73 & ~n_544) ;
	assign n_1605 = (~n_3 & n_1542) ;
	assign n_6955 = (~n_6952 & n_6954) ;
	assign n_7731 = (~n_7016 & n_7730) ;
	assign n_7009 = (~n_7007 & ~n_7008) ;
	assign n_7001 = (~x_71 & n_6999) ;
	assign n_7000 = (x_71 & ~n_6999) ;
	assign n_6992 = (~n_6990 & ~n_6991) ;
	assign n_6985 = (i_5 & ~n_6984) ;
	assign n_6983 = (~i_26 & n_544) ;
	assign n_6970 = (i_44 & n_7) ;
	assign n_6969 = (x_401 & ~n_16) ;
	assign n_1606 = (~n_59 & ~n_1605) ;
	assign n_6957 = (n_376 & ~n_6955) ;
	assign n_7732 = (~n_7009 & n_7731) ;
	assign n_7002 = (~n_7000 & ~n_7001) ;
	assign n_6994 = (~x_72 & n_6992) ;
	assign n_6993 = (x_72 & ~n_6992) ;
	assign n_6986 = (~n_6983 & n_6985) ;
	assign n_6978 = (i_8 & n_948) ;
	assign n_6977 = (x_74 & n_945) ;
	assign n_6971 = (~n_6969 & ~n_6970) ;
	assign n_6961 = (~n_376 & ~n_1606) ;
	assign n_6960 = (i_39 & n_7) ;
	assign n_6958 = (x_664 & ~n_6957) ;
	assign n_6956 = (~n_376 & n_6955) ;
	assign n_7733 = (~n_7002 & n_7732) ;
	assign n_6995 = (~n_6993 & ~n_6994) ;
	assign n_6988 = (~x_73 & ~n_6986) ;
	assign n_6987 = (x_73 & n_6986) ;
	assign n_6979 = (~n_6977 & ~n_6978) ;
	assign n_6972 = (n_20 & ~n_6971) ;
	assign n_6968 = (x_75 & n_18) ;
	assign n_6962 = (~n_6960 & ~n_6961) ;
	assign n_6959 = (~n_6956 & n_6958) ;
	assign n_7734 = (~n_6995 & n_7733) ;
	assign n_6989 = (~n_6987 & ~n_6988) ;
	assign n_6981 = (~x_74 & n_6979) ;
	assign n_6980 = (x_74 & ~n_6979) ;
	assign n_6973 = (~n_6968 & ~n_6972) ;
	assign n_6963 = (~n_6959 & n_6962) ;
	assign n_6945 = (i_11 & n_59) ;
	assign n_6921 = (x_80 & ~n_14) ;
	assign n_7735 = (~n_6989 & n_7734) ;
	assign n_6982 = (~n_6980 & ~n_6981) ;
	assign n_6975 = (~x_75 & n_6973) ;
	assign n_6974 = (x_75 & ~n_6973) ;
	assign n_6964 = (i_5 & ~n_6963) ;
	assign n_6946 = (n_66 & n_6945) ;
	assign n_6944 = (x_77 & n_60) ;
	assign n_6938 = (~x_78 & ~n_936) ;
	assign n_6922 = (n_12 & ~n_6921) ;
	assign n_6920 = (x_779 & n_14) ;
	assign n_6917 = (x_779 & n_11) ;
	assign n_7736 = (~n_6982 & n_7735) ;
	assign n_6976 = (~n_6974 & ~n_6975) ;
	assign n_6966 = (~x_76 & ~n_6964) ;
	assign n_6965 = (x_76 & n_6964) ;
	assign n_6947 = (~n_6944 & ~n_6946) ;
	assign n_6939 = (i_5 & ~n_6938) ;
	assign n_6937 = (~i_4 & n_936) ;
	assign n_6931 = (i_16 & n_59) ;
	assign n_6923 = (~n_6920 & n_6922) ;
	assign n_6918 = (x_168 & ~n_6917) ;
	assign n_6916 = (x_80 & ~n_11) ;
	assign n_6913 = (~x_80 & n_6) ;
	assign n_4406 = (~i_65 & ~n_6) ;
	assign n_6881 = (~n_422 & ~n_418) ;
	assign n_7737 = (~n_6976 & n_7736) ;
	assign n_6967 = (~n_6965 & ~n_6966) ;
	assign n_6949 = (~x_77 & n_6947) ;
	assign n_6948 = (x_77 & ~n_6947) ;
	assign n_6940 = (~n_6937 & n_6939) ;
	assign n_6932 = (n_66 & n_6931) ;
	assign n_6930 = (x_79 & n_60) ;
	assign n_6924 = (i_5 & ~n_6923) ;
	assign n_6919 = (~n_6916 & n_6918) ;
	assign n_6914 = (~n_4406 & ~n_6913) ;
	assign n_6883 = (~x_141 & ~n_6881) ;
	assign n_7738 = (~n_6967 & n_7737) ;
	assign n_6950 = (~n_6948 & ~n_6949) ;
	assign n_6942 = (~x_78 & ~n_6940) ;
	assign n_6941 = (x_78 & n_6940) ;
	assign n_6933 = (~n_6930 & ~n_6932) ;
	assign n_6925 = (~n_6919 & n_6924) ;
	assign n_6915 = (n_1 & ~n_6914) ;
	assign n_6884 = (n_527 & ~n_6883) ;
	assign n_6882 = (x_141 & n_6881) ;
	assign n_7739 = (~n_6950 & n_7738) ;
	assign n_6943 = (~n_6941 & ~n_6942) ;
	assign n_6935 = (~x_79 & n_6933) ;
	assign n_6934 = (x_79 & ~n_6933) ;
	assign n_6926 = (~n_6915 & n_6925) ;
	assign n_6908 = (i_18 & n_948) ;
	assign n_6907 = (x_81 & n_945) ;
	assign n_6890 = (n_6 & n_421) ;
	assign n_4732 = (~i_35 & ~n_6) ;
	assign n_6885 = (~n_6882 & n_6884) ;
	assign n_7740 = (~n_6943 & n_7739) ;
	assign n_6936 = (~n_6934 & ~n_6935) ;
	assign n_6928 = (~x_80 & ~n_6926) ;
	assign n_6927 = (x_80 & n_6926) ;
	assign n_6909 = (~n_6907 & ~n_6908) ;
	assign n_6902 = (x_485 & n_35) ;
	assign n_6901 = (x_82 & n_36) ;
	assign n_6891 = (~n_4732 & ~n_6890) ;
	assign n_6887 = (n_421 & n_6885) ;
	assign n_7741 = (~n_6936 & n_7740) ;
	assign n_6929 = (~n_6927 & ~n_6928) ;
	assign n_6911 = (~x_81 & n_6909) ;
	assign n_6910 = (x_81 & ~n_6909) ;
	assign n_6903 = (~n_6901 & ~n_6902) ;
	assign n_6892 = (n_1 & ~n_6891) ;
	assign n_6888 = (~n_1 & ~n_6887) ;
	assign n_6886 = (~n_421 & ~n_6885) ;
	assign n_7742 = (~n_6929 & n_7741) ;
	assign n_6912 = (~n_6910 & ~n_6911) ;
	assign n_6905 = (~x_82 & n_6903) ;
	assign n_6904 = (x_82 & ~n_6903) ;
	assign n_6893 = (i_5 & ~n_6892) ;
	assign n_6889 = (~n_6886 & n_6888) ;
	assign n_7743 = (~n_6912 & n_7742) ;
	assign n_6906 = (~n_6904 & ~n_6905) ;
	assign n_6899 = (~x_83 & n_218) ;
	assign n_6898 = (x_83 & ~n_218) ;
	assign n_6894 = (~n_6889 & n_6893) ;
	assign n_6876 = (i_37 & n_948) ;
	assign n_6875 = (x_85 & n_945) ;
	assign n_6869 = (i_25 & n_64) ;
	assign n_7744 = (~n_6906 & n_7743) ;
	assign n_6900 = (~n_6898 & ~n_6899) ;
	assign n_6896 = (~x_84 & ~n_6894) ;
	assign n_6895 = (x_84 & n_6894) ;
	assign n_6877 = (~n_6875 & ~n_6876) ;
	assign n_6870 = (n_66 & n_6869) ;
	assign n_6868 = (x_86 & n_978) ;
	assign n_7745 = (~n_6900 & n_7744) ;
	assign n_6897 = (~n_6895 & ~n_6896) ;
	assign n_6879 = (~x_85 & n_6877) ;
	assign n_6878 = (x_85 & ~n_6877) ;
	assign n_6871 = (~n_6868 & ~n_6870) ;
	assign n_6863 = (x_758 & n_53) ;
	assign n_6862 = (x_87 & n_51) ;
	assign n_7746 = (~n_6897 & n_7745) ;
	assign n_6880 = (~n_6878 & ~n_6879) ;
	assign n_6873 = (~x_86 & n_6871) ;
	assign n_6872 = (x_86 & ~n_6871) ;
	assign n_6864 = (~n_6862 & ~n_6863) ;
	assign n_6857 = (i_9 & n_948) ;
	assign n_6856 = (x_88 & n_945) ;
	assign n_7747 = (~n_6880 & n_7746) ;
	assign n_6874 = (~n_6872 & ~n_6873) ;
	assign n_6866 = (~x_87 & n_6864) ;
	assign n_6865 = (x_87 & ~n_6864) ;
	assign n_6858 = (~n_6856 & ~n_6857) ;
	assign n_6851 = (~n_86 & n_35) ;
	assign n_6850 = (x_89 & n_36) ;
	assign n_7748 = (~n_6874 & n_7747) ;
	assign n_6867 = (~n_6865 & ~n_6866) ;
	assign n_6860 = (~x_88 & n_6858) ;
	assign n_6859 = (x_88 & ~n_6858) ;
	assign n_6852 = (~n_6850 & ~n_6851) ;
	assign n_6845 = (~n_332 & n_1009) ;
	assign n_6844 = (x_90 & n_1007) ;
	assign n_6838 = (~x_91 & ~n_697) ;
	assign n_7749 = (~n_6867 & n_7748) ;
	assign n_6861 = (~n_6859 & ~n_6860) ;
	assign n_6854 = (~x_89 & n_6852) ;
	assign n_6853 = (x_89 & ~n_6852) ;
	assign n_6846 = (~n_6844 & ~n_6845) ;
	assign n_6839 = (i_5 & ~n_6838) ;
	assign n_6837 = (~x_600 & n_697) ;
	assign n_7750 = (~n_6861 & n_7749) ;
	assign n_6855 = (~n_6853 & ~n_6854) ;
	assign n_6848 = (~x_90 & n_6846) ;
	assign n_6847 = (x_90 & ~n_6846) ;
	assign n_6840 = (~n_6837 & n_6839) ;
	assign n_6828 = (~x_93 & ~n_630) ;
	assign n_7751 = (~n_6855 & n_7750) ;
	assign n_6849 = (~n_6847 & ~n_6848) ;
	assign n_6842 = (~x_91 & ~n_6840) ;
	assign n_6841 = (x_91 & n_6840) ;
	assign n_6829 = (i_5 & ~n_6828) ;
	assign n_6827 = (~i_39 & n_630) ;
	assign n_7752 = (~n_6849 & n_7751) ;
	assign n_6843 = (~n_6841 & ~n_6842) ;
	assign n_6835 = (~x_92 & n_347) ;
	assign n_6834 = (x_92 & ~n_347) ;
	assign n_6830 = (~n_6827 & n_6829) ;
	assign n_6822 = (x_709 & n_53) ;
	assign n_6821 = (x_94 & n_51) ;
	assign n_6815 = (i_17 & n_64) ;
	assign n_6807 = (~i_19 & n_669) ;
	assign n_7753 = (~n_6843 & n_7752) ;
	assign n_6836 = (~n_6834 & ~n_6835) ;
	assign n_6832 = (~x_93 & ~n_6830) ;
	assign n_6831 = (x_93 & n_6830) ;
	assign n_6823 = (~n_6821 & ~n_6822) ;
	assign n_6816 = (n_66 & n_6815) ;
	assign n_6814 = (x_95 & n_978) ;
	assign n_6808 = (i_5 & ~n_6807) ;
	assign n_6806 = (~x_407 & n_662) ;
	assign n_7754 = (~n_6836 & n_7753) ;
	assign n_6833 = (~n_6831 & ~n_6832) ;
	assign n_6825 = (~x_94 & n_6823) ;
	assign n_6824 = (x_94 & ~n_6823) ;
	assign n_6817 = (~n_6814 & ~n_6816) ;
	assign n_6809 = (~n_6806 & n_6808) ;
	assign n_6805 = (~x_96 & ~n_665) ;
	assign n_7755 = (~n_6833 & n_7754) ;
	assign n_6826 = (~n_6824 & ~n_6825) ;
	assign n_6819 = (~x_95 & n_6817) ;
	assign n_6818 = (x_95 & ~n_6817) ;
	assign n_6810 = (~n_6805 & n_6809) ;
	assign n_6800 = (~n_139 & n_1009) ;
	assign n_6799 = (x_97 & n_1007) ;
	assign n_6793 = (~x_98 & ~n_630) ;
	assign n_6770 = (~x_697 & ~n_44) ;
	assign n_1653 = (~x_718 & n_662) ;
	assign n_7756 = (~n_6826 & n_7755) ;
	assign n_6820 = (~n_6818 & ~n_6819) ;
	assign n_6812 = (~x_96 & ~n_6810) ;
	assign n_6811 = (x_96 & n_6810) ;
	assign n_6801 = (~n_6799 & ~n_6800) ;
	assign n_6794 = (i_5 & ~n_6793) ;
	assign n_6792 = (~i_41 & n_630) ;
	assign n_6786 = (i_29 & n_64) ;
	assign n_6771 = (n_662 & n_6770) ;
	assign n_6769 = (x_101 & ~n_1653) ;
	assign n_7757 = (~n_6820 & n_7756) ;
	assign n_6813 = (~n_6811 & ~n_6812) ;
	assign n_6803 = (~x_97 & n_6801) ;
	assign n_6802 = (x_97 & ~n_6801) ;
	assign n_6795 = (~n_6792 & n_6794) ;
	assign n_6787 = (n_66 & n_6786) ;
	assign n_6785 = (x_99 & n_978) ;
	assign n_6772 = (~n_6769 & ~n_6771) ;
	assign n_6767 = (~x_101 & ~n_3) ;
	assign n_1650 = (n_629 & ~n_5) ;
	assign n_7758 = (~n_6813 & n_7757) ;
	assign n_6804 = (~n_6802 & ~n_6803) ;
	assign n_6797 = (~x_98 & ~n_6795) ;
	assign n_6796 = (x_98 & n_6795) ;
	assign n_6788 = (~n_6785 & ~n_6787) ;
	assign n_6780 = (x_436 & n_53) ;
	assign n_6779 = (x_100 & n_51) ;
	assign n_6773 = (~n_629 & ~n_6772) ;
	assign n_6768 = (n_1650 & ~n_6767) ;
	assign n_7759 = (~n_6804 & n_7758) ;
	assign n_6798 = (~n_6796 & ~n_6797) ;
	assign n_6790 = (~x_99 & n_6788) ;
	assign n_6789 = (x_99 & ~n_6788) ;
	assign n_6781 = (~n_6779 & ~n_6780) ;
	assign n_6774 = (~n_6768 & ~n_6773) ;
	assign n_7760 = (~n_6798 & n_7759) ;
	assign n_6791 = (~n_6789 & ~n_6790) ;
	assign n_6783 = (~x_100 & n_6781) ;
	assign n_6782 = (x_100 & ~n_6781) ;
	assign n_6775 = (i_5 & ~n_6774) ;
	assign n_6762 = (~n_392 & n_1009) ;
	assign n_6761 = (x_102 & n_1007) ;
	assign n_7761 = (~n_6791 & n_7760) ;
	assign n_6784 = (~n_6782 & ~n_6783) ;
	assign n_6777 = (~x_101 & ~n_6775) ;
	assign n_6776 = (x_101 & n_6775) ;
	assign n_6763 = (~n_6761 & ~n_6762) ;
	assign n_6756 = (x_622 & n_53) ;
	assign n_6755 = (x_103 & n_51) ;
	assign n_6749 = (i_36 & n_64) ;
	assign n_7762 = (~n_6784 & n_7761) ;
	assign n_6778 = (~n_6776 & ~n_6777) ;
	assign n_6765 = (~x_102 & n_6763) ;
	assign n_6764 = (x_102 & ~n_6763) ;
	assign n_6757 = (~n_6755 & ~n_6756) ;
	assign n_6750 = (n_66 & n_6749) ;
	assign n_6748 = (x_104 & n_978) ;
	assign n_6742 = (i_63 & n_64) ;
	assign n_7763 = (~n_6778 & n_7762) ;
	assign n_6766 = (~n_6764 & ~n_6765) ;
	assign n_6759 = (~x_103 & n_6757) ;
	assign n_6758 = (x_103 & ~n_6757) ;
	assign n_6751 = (~n_6748 & ~n_6750) ;
	assign n_6743 = (n_66 & n_6742) ;
	assign n_6741 = (x_105 & n_978) ;
	assign n_6735 = (~x_106 & ~n_544) ;
	assign n_6727 = (~i_66 & n_669) ;
	assign n_6725 = (~x_270 & ~n_544) ;
	assign n_7764 = (~n_6766 & n_7763) ;
	assign n_6760 = (~n_6758 & ~n_6759) ;
	assign n_6753 = (~x_104 & n_6751) ;
	assign n_6752 = (x_104 & ~n_6751) ;
	assign n_6744 = (~n_6741 & ~n_6743) ;
	assign n_6736 = (i_5 & ~n_6735) ;
	assign n_6734 = (~i_30 & n_544) ;
	assign n_6728 = (i_5 & ~n_6727) ;
	assign n_6726 = (n_662 & n_6725) ;
	assign n_6678 = (~x_498 & n_1923) ;
	assign n_6677 = (x_498 & ~n_1923) ;
	assign n_7765 = (~n_6760 & n_7764) ;
	assign n_6754 = (~n_6752 & ~n_6753) ;
	assign n_6746 = (~x_105 & n_6744) ;
	assign n_6745 = (x_105 & ~n_6744) ;
	assign n_6737 = (~n_6734 & n_6736) ;
	assign n_6729 = (~n_6726 & n_6728) ;
	assign n_6724 = (~x_107 & ~n_665) ;
	assign n_6679 = (~n_6677 & ~n_6678) ;
	assign n_6676 = (~n_1913 & ~n_1914) ;
	assign n_7766 = (~n_6754 & n_7765) ;
	assign n_6747 = (~n_6745 & ~n_6746) ;
	assign n_6739 = (~x_106 & ~n_6737) ;
	assign n_6738 = (x_106 & n_6737) ;
	assign n_6730 = (~n_6724 & n_6729) ;
	assign n_6719 = (x_659 & n_53) ;
	assign n_6718 = (x_108 & n_51) ;
	assign n_6712 = (~x_109 & ~n_936) ;
	assign n_6688 = (i_10 & ~n_6) ;
	assign n_6681 = (n_6676 & ~n_6679) ;
	assign n_7767 = (~n_6747 & n_7766) ;
	assign n_6740 = (~n_6738 & ~n_6739) ;
	assign n_6732 = (~x_107 & ~n_6730) ;
	assign n_6731 = (x_107 & n_6730) ;
	assign n_6720 = (~n_6718 & ~n_6719) ;
	assign n_6713 = (i_5 & ~n_6712) ;
	assign n_6711 = (~i_49 & n_936) ;
	assign n_6705 = (~x_110 & ~n_697) ;
	assign n_6689 = (n_629 & ~n_6688) ;
	assign n_6687 = (x_112 & n_6) ;
	assign n_6684 = (x_112 & ~n_697) ;
	assign n_6682 = (n_697 & ~n_6681) ;
	assign n_6680 = (~n_6676 & n_6679) ;
	assign n_7768 = (~n_6740 & n_7767) ;
	assign n_6733 = (~n_6731 & ~n_6732) ;
	assign n_6722 = (~x_108 & n_6720) ;
	assign n_6721 = (x_108 & ~n_6720) ;
	assign n_6714 = (~n_6711 & n_6713) ;
	assign n_6706 = (i_5 & ~n_6705) ;
	assign n_6704 = (~x_538 & n_697) ;
	assign n_6698 = (i_32 & n_59) ;
	assign n_6690 = (~n_6687 & n_6689) ;
	assign n_6685 = (~n_629 & ~n_6684) ;
	assign n_6683 = (~n_6680 & n_6682) ;
	assign n_7769 = (~n_6733 & n_7768) ;
	assign n_6723 = (~n_6721 & ~n_6722) ;
	assign n_6716 = (~x_109 & ~n_6714) ;
	assign n_6715 = (x_109 & n_6714) ;
	assign n_6707 = (~n_6704 & n_6706) ;
	assign n_6699 = (n_66 & n_6698) ;
	assign n_6697 = (x_111 & n_60) ;
	assign n_6691 = (~n_6690 & n_902) ;
	assign n_6686 = (~n_6683 & n_6685) ;
	assign n_7770 = (~n_6723 & n_7769) ;
	assign n_6717 = (~n_6715 & ~n_6716) ;
	assign n_6709 = (~x_110 & ~n_6707) ;
	assign n_6708 = (x_110 & n_6707) ;
	assign n_6700 = (~n_6697 & ~n_6699) ;
	assign n_6692 = (~n_6686 & n_6691) ;
	assign n_6675 = (x_112 & n_699) ;
	assign n_471 = (x_331 & ~x_578) ;
	assign n_470 = (~x_255 & x_360) ;
	assign n_7771 = (~n_6717 & n_7770) ;
	assign n_6710 = (~n_6708 & ~n_6709) ;
	assign n_6702 = (~x_111 & n_6700) ;
	assign n_6701 = (x_111 & ~n_6700) ;
	assign n_6693 = (~n_6675 & ~n_6692) ;
	assign n_6670 = (~n_287 & n_1009) ;
	assign n_6669 = (x_113 & n_1007) ;
	assign n_6663 = (i_59 & n_59) ;
	assign n_475 = (x_637 & n_9) ;
	assign n_474 = (x_598 & n_13) ;
	assign n_472 = (~n_470 & ~n_471) ;
	assign n_7772 = (~n_6710 & n_7771) ;
	assign n_6703 = (~n_6701 & ~n_6702) ;
	assign n_6695 = (~x_112 & n_6693) ;
	assign n_6694 = (x_112 & ~n_6693) ;
	assign n_6671 = (~n_6669 & ~n_6670) ;
	assign n_6664 = (n_66 & n_6663) ;
	assign n_6662 = (x_114 & n_60) ;
	assign n_6656 = (i_12 & n_59) ;
	assign n_476 = (~n_474 & ~n_475) ;
	assign n_473 = (~n_9 & ~n_472) ;
	assign n_468 = (~n_464 & ~n_467) ;
	assign n_7773 = (~n_6703 & n_7772) ;
	assign n_6696 = (~n_6694 & ~n_6695) ;
	assign n_6673 = (~x_113 & n_6671) ;
	assign n_6672 = (x_113 & ~n_6671) ;
	assign n_6665 = (~n_6662 & ~n_6664) ;
	assign n_6657 = (n_66 & n_6656) ;
	assign n_6655 = (x_115 & n_60) ;
	assign n_6649 = (i_37 & n_64) ;
	assign n_486 = (~x_255 & x_285) ;
	assign n_485 = (x_406 & ~x_578) ;
	assign n_481 = (~x_527 & x_695) ;
	assign n_480 = (x_527 & x_645) ;
	assign n_477 = (~n_473 & n_476) ;
	assign n_469 = (~n_463 & ~n_468) ;
	assign n_7774 = (~n_6696 & n_7773) ;
	assign n_6674 = (~n_6672 & ~n_6673) ;
	assign n_6667 = (~x_114 & n_6665) ;
	assign n_6666 = (x_114 & ~n_6665) ;
	assign n_6658 = (~n_6655 & ~n_6657) ;
	assign n_6650 = (n_66 & n_6649) ;
	assign n_6648 = (x_116 & n_978) ;
	assign n_6642 = (~x_117 & ~n_697) ;
	assign n_490 = (x_551 & n_9) ;
	assign n_489 = (x_686 & n_13) ;
	assign n_487 = (~n_485 & ~n_486) ;
	assign n_482 = (~n_480 & ~n_481) ;
	assign n_479 = (n_469 & n_477) ;
	assign n_7775 = (~n_6674 & n_7774) ;
	assign n_6668 = (~n_6666 & ~n_6667) ;
	assign n_6660 = (~x_115 & n_6658) ;
	assign n_6659 = (x_115 & ~n_6658) ;
	assign n_6651 = (~n_6648 & ~n_6650) ;
	assign n_6643 = (i_5 & ~n_6642) ;
	assign n_6641 = (~x_627 & n_697) ;
	assign n_6635 = (~x_118 & ~n_936) ;
	assign n_491 = (~n_489 & ~n_490) ;
	assign n_488 = (~n_9 & ~n_487) ;
	assign n_483 = (~n_479 & ~n_482) ;
	assign n_478 = (~n_469 & ~n_477) ;
	assign n_7776 = (~n_6668 & n_7775) ;
	assign n_6661 = (~n_6659 & ~n_6660) ;
	assign n_6653 = (~x_116 & n_6651) ;
	assign n_6652 = (x_116 & ~n_6651) ;
	assign n_6644 = (~n_6641 & n_6643) ;
	assign n_6636 = (i_5 & ~n_6635) ;
	assign n_6634 = (~i_38 & n_936) ;
	assign n_501 = (x_421 & ~x_578) ;
	assign n_500 = (~x_255 & x_528) ;
	assign n_496 = (~x_527 & x_628) ;
	assign n_495 = (x_204 & x_527) ;
	assign n_492 = (~n_488 & n_491) ;
	assign n_484 = (~n_478 & ~n_483) ;
	assign n_7777 = (~n_6661 & n_7776) ;
	assign n_6654 = (~n_6652 & ~n_6653) ;
	assign n_6646 = (~x_117 & ~n_6644) ;
	assign n_6645 = (x_117 & n_6644) ;
	assign n_6637 = (~n_6634 & n_6636) ;
	assign n_6629 = (i_25 & n_948) ;
	assign n_6628 = (x_119 & n_945) ;
	assign n_6622 = (~x_120 & ~n_630) ;
	assign n_6582 = (x_759 & n_181) ;
	assign n_6581 = (~x_759 & ~n_181) ;
	assign n_505 = (x_263 & n_9) ;
	assign n_504 = (x_151 & n_13) ;
	assign n_502 = (~n_500 & ~n_501) ;
	assign n_497 = (~n_495 & ~n_496) ;
	assign n_494 = (n_484 & n_492) ;
	assign n_7778 = (~n_6654 & n_7777) ;
	assign n_6647 = (~n_6645 & ~n_6646) ;
	assign n_6639 = (~x_118 & ~n_6637) ;
	assign n_6638 = (x_118 & n_6637) ;
	assign n_6630 = (~n_6628 & ~n_6629) ;
	assign n_6623 = (i_5 & ~n_6622) ;
	assign n_6621 = (~i_40 & n_630) ;
	assign n_6615 = (~x_121 & ~n_630) ;
	assign n_6583 = (~n_6581 & ~n_6582) ;
	assign n_506 = (~n_504 & ~n_505) ;
	assign n_503 = (~n_9 & ~n_502) ;
	assign n_498 = (~n_494 & ~n_497) ;
	assign n_493 = (~n_484 & ~n_492) ;
	assign n_7779 = (~n_6647 & n_7778) ;
	assign n_6640 = (~n_6638 & ~n_6639) ;
	assign n_6632 = (~x_119 & n_6630) ;
	assign n_6631 = (x_119 & ~n_6630) ;
	assign n_6624 = (~n_6621 & n_6623) ;
	assign n_6616 = (i_5 & ~n_6615) ;
	assign n_6614 = (~i_36 & n_630) ;
	assign n_6585 = (n_115 & ~n_527) ;
	assign n_6584 = (n_527 & ~n_6583) ;
	assign n_507 = (~n_503 & n_506) ;
	assign n_499 = (~n_493 & ~n_498) ;
	assign n_7780 = (~n_6640 & n_7779) ;
	assign n_6633 = (~n_6631 & ~n_6632) ;
	assign n_6626 = (~x_120 & ~n_6624) ;
	assign n_6625 = (x_120 & n_6624) ;
	assign n_6617 = (~n_6614 & n_6616) ;
	assign n_6586 = (~n_6584 & ~n_6585) ;
	assign n_6580 = (~n_116 & ~n_117) ;
	assign n_508 = (~n_499 & ~n_507) ;
	assign n_512 = (n_499 & n_507) ;
	assign n_7781 = (~n_6633 & n_7780) ;
	assign n_6627 = (~n_6625 & ~n_6626) ;
	assign n_6619 = (~x_121 & ~n_6617) ;
	assign n_6618 = (x_121 & n_6617) ;
	assign n_6606 = (x_401 & n_35) ;
	assign n_6605 = (x_123 & n_36) ;
	assign n_6599 = (~x_124 & ~n_936) ;
	assign n_4147 = (~i_31 & ~n_6) ;
	assign n_6588 = (~n_6580 & ~n_6586) ;
	assign n_6543 = (~n_512 & ~n_508) ;
	assign n_7782 = (~n_6627 & n_7781) ;
	assign n_6620 = (~n_6618 & ~n_6619) ;
	assign n_6612 = (~x_122 & n_436) ;
	assign n_6611 = (x_122 & ~n_436) ;
	assign n_6607 = (~n_6605 & ~n_6606) ;
	assign n_6600 = (i_5 & ~n_6599) ;
	assign n_6598 = (~i_13 & n_936) ;
	assign n_6592 = (n_947 & ~n_4147) ;
	assign n_6591 = (n_6 & n_107) ;
	assign n_6589 = (n_29 & ~n_6588) ;
	assign n_6587 = (n_6580 & n_6586) ;
	assign n_510 = (x_173 & ~x_527) ;
	assign n_509 = (x_129 & x_527) ;
	assign n_6545 = (~x_460 & ~n_6543) ;
	assign n_7783 = (~n_6620 & n_7782) ;
	assign n_6613 = (~n_6611 & ~n_6612) ;
	assign n_6609 = (~x_123 & n_6607) ;
	assign n_6608 = (x_123 & ~n_6607) ;
	assign n_6601 = (~n_6598 & n_6600) ;
	assign n_6593 = (~n_6591 & n_6592) ;
	assign n_6590 = (~n_6587 & n_6589) ;
	assign n_6574 = (~x_126 & ~n_544) ;
	assign n_511 = (~n_509 & ~n_510) ;
	assign n_6546 = (n_527 & ~n_6545) ;
	assign n_6544 = (x_460 & n_6543) ;
	assign n_7784 = (~n_6613 & n_7783) ;
	assign n_6610 = (~n_6608 & ~n_6609) ;
	assign n_6603 = (~x_124 & ~n_6601) ;
	assign n_6602 = (x_124 & n_6601) ;
	assign n_6594 = (~n_6590 & ~n_6593) ;
	assign n_6575 = (i_5 & ~n_6574) ;
	assign n_6573 = (~i_22 & n_544) ;
	assign n_4440 = (~i_64 & ~n_6) ;
	assign n_6552 = (n_6 & n_511) ;
	assign n_6547 = (~n_6544 & n_6546) ;
	assign n_7785 = (~n_6610 & n_7784) ;
	assign n_6604 = (~n_6602 & ~n_6603) ;
	assign n_6596 = (~x_125 & n_6594) ;
	assign n_6595 = (x_125 & ~n_6594) ;
	assign n_6576 = (~n_6573 & n_6575) ;
	assign n_6568 = (i_53 & n_948) ;
	assign n_6567 = (x_127 & n_945) ;
	assign n_6561 = (~x_128 & ~n_544) ;
	assign n_6553 = (~n_6552 & ~n_4440) ;
	assign n_6549 = (n_511 & n_6547) ;
	assign n_7786 = (~n_6604 & n_7785) ;
	assign n_6597 = (~n_6595 & ~n_6596) ;
	assign n_6578 = (~x_126 & ~n_6576) ;
	assign n_6577 = (x_126 & n_6576) ;
	assign n_6569 = (~n_6567 & ~n_6568) ;
	assign n_6562 = (i_5 & ~n_6561) ;
	assign n_6560 = (~i_32 & n_544) ;
	assign n_6554 = (n_1 & ~n_6553) ;
	assign n_6550 = (~n_1 & ~n_6549) ;
	assign n_6548 = (~n_511 & ~n_6547) ;
	assign n_7787 = (~n_6597 & n_7786) ;
	assign n_6579 = (~n_6577 & ~n_6578) ;
	assign n_6571 = (~x_127 & n_6569) ;
	assign n_6570 = (x_127 & ~n_6569) ;
	assign n_6563 = (~n_6560 & n_6562) ;
	assign n_6555 = (i_5 & ~n_6554) ;
	assign n_6551 = (~n_6548 & n_6550) ;
	assign n_7788 = (~n_6579 & n_7787) ;
	assign n_6572 = (~n_6570 & ~n_6571) ;
	assign n_6565 = (~x_128 & ~n_6563) ;
	assign n_6564 = (x_128 & n_6563) ;
	assign n_6556 = (~n_6551 & n_6555) ;
	assign n_6527 = (i_27 & n_7) ;
	assign n_6526 = (x_569 & ~n_16) ;
	assign n_7789 = (~n_6572 & n_7788) ;
	assign n_6566 = (~n_6564 & ~n_6565) ;
	assign n_6558 = (~x_129 & ~n_6556) ;
	assign n_6557 = (x_129 & n_6556) ;
	assign n_6535 = (x_97 & n_35) ;
	assign n_6534 = (x_131 & n_36) ;
	assign n_6528 = (~n_6526 & ~n_6527) ;
	assign n_7790 = (~n_6566 & n_7789) ;
	assign n_6559 = (~n_6557 & ~n_6558) ;
	assign n_6541 = (~x_130 & n_287) ;
	assign n_6540 = (x_130 & ~n_287) ;
	assign n_6536 = (~n_6534 & ~n_6535) ;
	assign n_6529 = (n_20 & ~n_6528) ;
	assign n_6525 = (x_132 & n_18) ;
	assign n_6519 = (~x_133 & ~n_544) ;
	assign n_6472 = (~n_358 & ~n_359) ;
	assign n_7791 = (~n_6559 & n_7790) ;
	assign n_6542 = (~n_6540 & ~n_6541) ;
	assign n_6538 = (~x_131 & n_6536) ;
	assign n_6537 = (x_131 & ~n_6536) ;
	assign n_6530 = (~n_6525 & ~n_6529) ;
	assign n_6520 = (i_5 & ~n_6519) ;
	assign n_6518 = (~i_12 & n_544) ;
	assign n_6474 = (~x_782 & ~n_6472) ;
	assign n_7792 = (~n_6542 & n_7791) ;
	assign n_6539 = (~n_6537 & ~n_6538) ;
	assign n_6532 = (~x_132 & n_6530) ;
	assign n_6531 = (x_132 & ~n_6530) ;
	assign n_6521 = (~n_6518 & n_6520) ;
	assign n_6513 = (~n_203 & n_35) ;
	assign n_6512 = (x_134 & n_36) ;
	assign n_6506 = (x_391 & n_697) ;
	assign n_2348 = (i_5 & ~n_629) ;
	assign n_6475 = (n_527 & ~n_6474) ;
	assign n_6473 = (x_782 & n_6472) ;
	assign n_7793 = (~n_6539 & n_7792) ;
	assign n_6533 = (~n_6531 & ~n_6532) ;
	assign n_6523 = (~x_133 & ~n_6521) ;
	assign n_6522 = (x_133 & n_6521) ;
	assign n_6514 = (~n_6512 & ~n_6513) ;
	assign n_6507 = (n_2348 & n_6506) ;
	assign n_6505 = (x_135 & n_698) ;
	assign n_6492 = (~i_22 & n_669) ;
	assign n_6490 = (~x_363 & ~n_544) ;
	assign n_2393 = (~i_62 & ~n_6) ;
	assign n_6481 = (n_6 & n_362) ;
	assign n_6476 = (~n_6473 & n_6475) ;
	assign n_7794 = (~n_6533 & n_7793) ;
	assign n_6524 = (~n_6522 & ~n_6523) ;
	assign n_6516 = (~x_134 & n_6514) ;
	assign n_6515 = (x_134 & ~n_6514) ;
	assign n_6508 = (~n_6505 & ~n_6507) ;
	assign n_6500 = (x_102 & n_35) ;
	assign n_6499 = (x_136 & n_36) ;
	assign n_6493 = (i_5 & ~n_6492) ;
	assign n_6491 = (n_662 & n_6490) ;
	assign n_6482 = (~n_6481 & ~n_2393) ;
	assign n_6478 = (n_362 & n_6476) ;
	assign n_7795 = (~n_6524 & n_7794) ;
	assign n_6517 = (~n_6515 & ~n_6516) ;
	assign n_6510 = (~x_135 & n_6508) ;
	assign n_6509 = (x_135 & ~n_6508) ;
	assign n_6501 = (~n_6499 & ~n_6500) ;
	assign n_6494 = (~n_6491 & n_6493) ;
	assign n_6489 = (~x_137 & ~n_665) ;
	assign n_6483 = (n_1 & ~n_6482) ;
	assign n_6479 = (~n_1 & ~n_6478) ;
	assign n_6477 = (~n_362 & ~n_6476) ;
	assign n_6458 = (i_57 & n_1) ;
	assign n_6457 = (~x_140 & n_6) ;
	assign n_7796 = (~n_6517 & n_7795) ;
	assign n_6511 = (~n_6509 & ~n_6510) ;
	assign n_6503 = (~x_136 & n_6501) ;
	assign n_6502 = (x_136 & ~n_6501) ;
	assign n_6495 = (~n_6489 & n_6494) ;
	assign n_6484 = (i_5 & ~n_6483) ;
	assign n_6480 = (~n_6477 & n_6479) ;
	assign n_6459 = (~n_6457 & n_6458) ;
	assign n_6456 = (x_463 & ~n_16) ;
	assign n_6447 = (i_21 & n_1) ;
	assign n_6446 = (~x_141 & n_6) ;
	assign n_7797 = (~n_6511 & n_7796) ;
	assign n_6504 = (~n_6502 & ~n_6503) ;
	assign n_6497 = (~x_137 & ~n_6495) ;
	assign n_6496 = (x_137 & n_6495) ;
	assign n_6485 = (~n_6480 & n_6484) ;
	assign n_6467 = (i_58 & n_948) ;
	assign n_6466 = (x_139 & n_945) ;
	assign n_6460 = (~n_6456 & ~n_6459) ;
	assign n_6455 = (x_140 & n_17) ;
	assign n_6448 = (~n_6446 & n_6447) ;
	assign n_6445 = (x_644 & ~n_16) ;
	assign n_7798 = (~n_6504 & n_7797) ;
	assign n_6498 = (~n_6496 & ~n_6497) ;
	assign n_6487 = (~x_138 & ~n_6485) ;
	assign n_6486 = (x_138 & n_6485) ;
	assign n_6468 = (~n_6466 & ~n_6467) ;
	assign n_6461 = (~n_6455 & n_6460) ;
	assign n_6449 = (~n_6445 & ~n_6448) ;
	assign n_6444 = (x_141 & n_17) ;
	assign n_7799 = (~n_6498 & n_7798) ;
	assign n_6488 = (~n_6486 & ~n_6487) ;
	assign n_6470 = (~x_139 & n_6468) ;
	assign n_6469 = (x_139 & ~n_6468) ;
	assign n_6462 = (i_5 & ~n_6461) ;
	assign n_6450 = (~n_6444 & n_6449) ;
	assign n_7800 = (~n_6488 & n_7799) ;
	assign n_6471 = (~n_6469 & ~n_6470) ;
	assign n_6464 = (~x_140 & ~n_6462) ;
	assign n_6463 = (x_140 & n_6462) ;
	assign n_6451 = (i_5 & ~n_6450) ;
	assign n_6439 = (x_447 & n_53) ;
	assign n_6438 = (x_142 & n_51) ;
	assign n_6432 = (i_7 & n_59) ;
	assign n_7801 = (~n_6471 & n_7800) ;
	assign n_6465 = (~n_6463 & ~n_6464) ;
	assign n_6453 = (~x_141 & ~n_6451) ;
	assign n_6452 = (x_141 & n_6451) ;
	assign n_6440 = (~n_6438 & ~n_6439) ;
	assign n_6433 = (n_66 & n_6432) ;
	assign n_6431 = (x_143 & n_60) ;
	assign n_6425 = (~x_144 & ~n_936) ;
	assign n_7802 = (~n_6465 & n_7801) ;
	assign n_6454 = (~n_6452 & ~n_6453) ;
	assign n_6442 = (~x_142 & n_6440) ;
	assign n_6441 = (x_142 & ~n_6440) ;
	assign n_6434 = (~n_6431 & ~n_6433) ;
	assign n_6426 = (i_5 & ~n_6425) ;
	assign n_6424 = (~i_42 & n_936) ;
	assign n_6418 = (~x_145 & ~n_544) ;
	assign n_7803 = (~n_6454 & n_7802) ;
	assign n_6443 = (~n_6441 & ~n_6442) ;
	assign n_6436 = (~x_143 & n_6434) ;
	assign n_6435 = (x_143 & ~n_6434) ;
	assign n_6427 = (~n_6424 & n_6426) ;
	assign n_6419 = (i_5 & ~n_6418) ;
	assign n_6417 = (~i_33 & n_544) ;
	assign n_6411 = (~x_146 & ~n_544) ;
	assign n_7804 = (~n_6443 & n_7803) ;
	assign n_6437 = (~n_6435 & ~n_6436) ;
	assign n_6429 = (~x_144 & ~n_6427) ;
	assign n_6428 = (x_144 & n_6427) ;
	assign n_6420 = (~n_6417 & n_6419) ;
	assign n_6412 = (i_5 & ~n_6411) ;
	assign n_6410 = (~i_19 & n_544) ;
	assign n_7805 = (~n_6437 & n_7804) ;
	assign n_6430 = (~n_6428 & ~n_6429) ;
	assign n_6422 = (~x_145 & ~n_6420) ;
	assign n_6421 = (x_145 & n_6420) ;
	assign n_6413 = (~n_6410 & n_6412) ;
	assign n_6405 = (x_600 & n_53) ;
	assign n_6404 = (x_147 & n_51) ;
	assign n_7806 = (~n_6430 & n_7805) ;
	assign n_6423 = (~n_6421 & ~n_6422) ;
	assign n_6415 = (~x_146 & ~n_6413) ;
	assign n_6414 = (x_146 & n_6413) ;
	assign n_6406 = (~n_6404 & ~n_6405) ;
	assign n_6399 = (n_35 & ~n_407) ;
	assign n_6398 = (x_148 & n_36) ;
	assign n_6392 = (~x_149 & ~n_544) ;
	assign n_7807 = (~n_6423 & n_7806) ;
	assign n_6416 = (~n_6414 & ~n_6415) ;
	assign n_6408 = (~x_147 & n_6406) ;
	assign n_6407 = (x_147 & ~n_6406) ;
	assign n_6400 = (~n_6398 & ~n_6399) ;
	assign n_6393 = (i_5 & ~n_6392) ;
	assign n_6391 = (~i_38 & n_544) ;
	assign n_6385 = (~x_150 & ~n_544) ;
	assign n_6340 = (~n_433 & ~n_437) ;
	assign n_7808 = (~n_6416 & n_7807) ;
	assign n_6409 = (~n_6407 & ~n_6408) ;
	assign n_6402 = (~x_148 & n_6400) ;
	assign n_6401 = (x_148 & ~n_6400) ;
	assign n_6394 = (~n_6391 & n_6393) ;
	assign n_6386 = (i_5 & ~n_6385) ;
	assign n_6384 = (~i_52 & n_544) ;
	assign n_6378 = (i_34 & n_59) ;
	assign n_6342 = (~x_227 & ~n_6340) ;
	assign n_7809 = (~n_6409 & n_7808) ;
	assign n_6403 = (~n_6401 & ~n_6402) ;
	assign n_6396 = (~x_149 & ~n_6394) ;
	assign n_6395 = (x_149 & n_6394) ;
	assign n_6387 = (~n_6384 & n_6386) ;
	assign n_6379 = (n_66 & n_6378) ;
	assign n_6377 = (x_151 & n_60) ;
	assign n_6371 = (i_40 & n_59) ;
	assign n_6343 = (n_527 & ~n_6342) ;
	assign n_6341 = (x_227 & n_6340) ;
	assign n_7810 = (~n_6403 & n_7809) ;
	assign n_6397 = (~n_6395 & ~n_6396) ;
	assign n_6389 = (~x_150 & ~n_6387) ;
	assign n_6388 = (x_150 & n_6387) ;
	assign n_6380 = (~n_6377 & ~n_6379) ;
	assign n_6372 = (n_66 & n_6371) ;
	assign n_6370 = (x_152 & n_60) ;
	assign n_6349 = (n_6 & n_436) ;
	assign n_6344 = (~n_6341 & n_6343) ;
	assign n_7811 = (~n_6397 & n_7810) ;
	assign n_6390 = (~n_6388 & ~n_6389) ;
	assign n_6382 = (~x_151 & n_6380) ;
	assign n_6381 = (x_151 & ~n_6380) ;
	assign n_6373 = (~n_6370 & ~n_6372) ;
	assign n_6365 = (i_41 & n_948) ;
	assign n_6364 = (x_153 & n_945) ;
	assign n_6351 = (~n_6349 & ~n_6350) ;
	assign n_6346 = (n_436 & n_6344) ;
	assign n_7812 = (~n_6390 & n_7811) ;
	assign n_6383 = (~n_6381 & ~n_6382) ;
	assign n_6375 = (~x_152 & n_6373) ;
	assign n_6374 = (x_152 & ~n_6373) ;
	assign n_6366 = (~n_6364 & ~n_6365) ;
	assign n_6359 = (x_408 & n_35) ;
	assign n_6358 = (x_154 & n_36) ;
	assign n_6352 = (n_1 & ~n_6351) ;
	assign n_6347 = (~n_1 & ~n_6346) ;
	assign n_6345 = (~n_436 & ~n_6344) ;
	assign n_7813 = (~n_6383 & n_7812) ;
	assign n_6376 = (~n_6374 & ~n_6375) ;
	assign n_6368 = (~x_153 & n_6366) ;
	assign n_6367 = (x_153 & ~n_6366) ;
	assign n_6360 = (~n_6358 & ~n_6359) ;
	assign n_6353 = (i_5 & ~n_6352) ;
	assign n_6348 = (~n_6345 & n_6347) ;
	assign n_7814 = (~n_6376 & n_7813) ;
	assign n_6369 = (~n_6367 & ~n_6368) ;
	assign n_6362 = (~x_154 & n_6360) ;
	assign n_6361 = (x_154 & ~n_6360) ;
	assign n_6354 = (~n_6348 & n_6353) ;
	assign n_6335 = (i_68 & n_948) ;
	assign n_6334 = (x_156 & n_945) ;
	assign n_6328 = (~x_157 & ~n_630) ;
	assign n_7815 = (~n_6369 & n_7814) ;
	assign n_6363 = (~n_6361 & ~n_6362) ;
	assign n_6356 = (~x_155 & ~n_6354) ;
	assign n_6355 = (x_155 & n_6354) ;
	assign n_6336 = (~n_6334 & ~n_6335) ;
	assign n_6329 = (i_5 & ~n_6328) ;
	assign n_6327 = (~i_48 & n_630) ;
	assign n_7816 = (~n_6363 & n_7815) ;
	assign n_6357 = (~n_6355 & ~n_6356) ;
	assign n_6338 = (~x_156 & n_6336) ;
	assign n_6337 = (x_156 & ~n_6336) ;
	assign n_6330 = (~n_6327 & n_6329) ;
	assign n_6322 = (i_51 & n_948) ;
	assign n_6321 = (x_158 & n_945) ;
	assign n_7817 = (~n_6357 & n_7816) ;
	assign n_6339 = (~n_6337 & ~n_6338) ;
	assign n_6332 = (~x_157 & ~n_6330) ;
	assign n_6331 = (x_157 & n_6330) ;
	assign n_6323 = (~n_6321 & ~n_6322) ;
	assign n_6316 = (x_275 & n_53) ;
	assign n_6315 = (x_159 & n_51) ;
	assign n_7818 = (~n_6339 & n_7817) ;
	assign n_6333 = (~n_6331 & ~n_6332) ;
	assign n_6325 = (~x_158 & n_6323) ;
	assign n_6324 = (x_158 & ~n_6323) ;
	assign n_6317 = (~n_6315 & ~n_6316) ;
	assign n_6306 = (~x_161 & ~n_936) ;
	assign n_6267 = (~x_96 & n_851) ;
	assign n_6266 = (x_96 & ~n_851) ;
	assign n_7819 = (~n_6333 & n_7818) ;
	assign n_6326 = (~n_6324 & ~n_6325) ;
	assign n_6319 = (~x_159 & n_6317) ;
	assign n_6318 = (x_159 & ~n_6317) ;
	assign n_6307 = (i_5 & ~n_6306) ;
	assign n_6305 = (~i_57 & n_936) ;
	assign n_6268 = (~n_6266 & ~n_6267) ;
	assign n_6265 = (~n_841 & ~n_842) ;
	assign n_7820 = (~n_6326 & n_7819) ;
	assign n_6320 = (~n_6318 & ~n_6319) ;
	assign n_6313 = (~x_160 & n_362) ;
	assign n_6312 = (x_160 & ~n_362) ;
	assign n_6308 = (~n_6305 & n_6307) ;
	assign n_6277 = (i_18 & ~n_6) ;
	assign n_6270 = (n_6265 & ~n_6268) ;
	assign n_7821 = (~n_6320 & n_7820) ;
	assign n_6314 = (~n_6312 & ~n_6313) ;
	assign n_6310 = (~x_161 & ~n_6308) ;
	assign n_6309 = (x_161 & n_6308) ;
	assign n_6297 = (~n_332 & n_35) ;
	assign n_6296 = (x_163 & n_36) ;
	assign n_1582 = (i_49 & n_59) ;
	assign n_6278 = (n_629 & ~n_6277) ;
	assign n_6276 = (x_166 & n_6) ;
	assign n_6273 = (x_166 & ~n_697) ;
	assign n_6271 = (n_697 & ~n_6270) ;
	assign n_6269 = (~n_6265 & n_6268) ;
	assign n_7822 = (~n_6314 & n_7821) ;
	assign n_6311 = (~n_6309 & ~n_6310) ;
	assign n_6303 = (~x_162 & n_136) ;
	assign n_6302 = (x_162 & ~n_136) ;
	assign n_6298 = (~n_6296 & ~n_6297) ;
	assign n_1583 = (n_66 & n_1582) ;
	assign n_1581 = (x_164 & n_60) ;
	assign n_6287 = (~x_165 & ~n_630) ;
	assign n_6279 = (~n_6276 & n_6278) ;
	assign n_6274 = (~n_629 & ~n_6273) ;
	assign n_6272 = (~n_6269 & n_6271) ;
	assign n_7823 = (~n_6311 & n_7822) ;
	assign n_6304 = (~n_6302 & ~n_6303) ;
	assign n_6300 = (~x_163 & n_6298) ;
	assign n_6299 = (x_163 & ~n_6298) ;
	assign n_1584 = (~n_1581 & ~n_1583) ;
	assign n_6288 = (i_5 & ~n_6287) ;
	assign n_6286 = (~i_53 & n_630) ;
	assign n_6280 = (n_902 & ~n_6279) ;
	assign n_6275 = (~n_6272 & n_6274) ;
	assign n_7824 = (~n_6304 & n_7823) ;
	assign n_6301 = (~n_6299 & ~n_6300) ;
	assign n_6294 = (~x_164 & n_1584) ;
	assign n_6293 = (x_164 & ~n_1584) ;
	assign n_6289 = (~n_6286 & n_6288) ;
	assign n_6281 = (~n_6275 & n_6280) ;
	assign n_6264 = (x_166 & n_699) ;
	assign n_6258 = (i_33 & n_59) ;
	assign n_1818 = (~n_63 & ~n_3) ;
	assign n_7825 = (~n_6301 & n_7824) ;
	assign n_6295 = (~n_6293 & ~n_6294) ;
	assign n_6291 = (~x_165 & ~n_6289) ;
	assign n_6290 = (x_165 & n_6289) ;
	assign n_6282 = (~n_6264 & ~n_6281) ;
	assign n_6259 = (n_66 & n_6258) ;
	assign n_6257 = (x_167 & n_60) ;
	assign n_6251 = (n_1542 & ~n_1818) ;
	assign n_6250 = (n_8 & ~n_30) ;
	assign n_6243 = (i_37 & n_7) ;
	assign n_6242 = (x_792 & ~n_16) ;
	assign n_7826 = (~n_6295 & n_7825) ;
	assign n_6292 = (~n_6290 & ~n_6291) ;
	assign n_6284 = (~x_166 & n_6282) ;
	assign n_6283 = (x_166 & ~n_6282) ;
	assign n_6260 = (~n_6257 & ~n_6259) ;
	assign n_6252 = (~n_6250 & ~n_6251) ;
	assign n_6244 = (~n_6242 & ~n_6243) ;
	assign n_7827 = (~n_6292 & n_7826) ;
	assign n_6285 = (~n_6283 & ~n_6284) ;
	assign n_6262 = (~x_167 & n_6260) ;
	assign n_6261 = (x_167 & ~n_6260) ;
	assign n_6253 = (i_5 & ~n_6252) ;
	assign n_6245 = (n_20 & ~n_6244) ;
	assign n_6241 = (x_169 & n_18) ;
	assign n_7828 = (~n_6285 & n_7827) ;
	assign n_6263 = (~n_6261 & ~n_6262) ;
	assign n_6255 = (~x_168 & ~n_6253) ;
	assign n_6254 = (x_168 & n_6253) ;
	assign n_6246 = (~n_6241 & ~n_6245) ;
	assign n_6236 = (i_46 & n_948) ;
	assign n_6235 = (x_170 & n_945) ;
	assign n_6229 = (~x_171 & ~n_936) ;
	assign n_7829 = (~n_6263 & n_7828) ;
	assign n_6256 = (~n_6254 & ~n_6255) ;
	assign n_6248 = (~x_169 & n_6246) ;
	assign n_6247 = (x_169 & ~n_6246) ;
	assign n_6237 = (~n_6235 & ~n_6236) ;
	assign n_6230 = (i_5 & ~n_6229) ;
	assign n_6228 = (~i_39 & n_936) ;
	assign n_6222 = (~x_172 & ~n_630) ;
	assign n_7830 = (~n_6256 & n_7829) ;
	assign n_6249 = (~n_6247 & ~n_6248) ;
	assign n_6239 = (~x_170 & n_6237) ;
	assign n_6238 = (x_170 & ~n_6237) ;
	assign n_6231 = (~n_6228 & n_6230) ;
	assign n_6223 = (i_5 & ~n_6222) ;
	assign n_6221 = (~i_29 & n_630) ;
	assign n_7831 = (~n_6249 & n_7830) ;
	assign n_6240 = (~n_6238 & ~n_6239) ;
	assign n_6233 = (~x_171 & ~n_6231) ;
	assign n_6232 = (x_171 & n_6231) ;
	assign n_6224 = (~n_6221 & n_6223) ;
	assign n_7832 = (~n_6240 & n_7831) ;
	assign n_6234 = (~n_6232 & ~n_6233) ;
	assign n_6226 = (~x_172 & ~n_6224) ;
	assign n_6225 = (x_172 & n_6224) ;
	assign n_6213 = (x_178 & n_53) ;
	assign n_6212 = (x_174 & n_51) ;
	assign n_6206 = (~x_175 & ~n_936) ;
	assign n_7833 = (~n_6234 & n_7832) ;
	assign n_6227 = (~n_6225 & ~n_6226) ;
	assign n_6219 = (~x_173 & n_511) ;
	assign n_6218 = (x_173 & ~n_511) ;
	assign n_6214 = (~n_6212 & ~n_6213) ;
	assign n_6207 = (i_5 & ~n_6206) ;
	assign n_6205 = (~i_19 & n_936) ;
	assign n_6199 = (i_39 & n_59) ;
	assign n_7834 = (~n_6227 & n_7833) ;
	assign n_6220 = (~n_6218 & ~n_6219) ;
	assign n_6216 = (~x_174 & n_6214) ;
	assign n_6215 = (x_174 & ~n_6214) ;
	assign n_6208 = (~n_6205 & n_6207) ;
	assign n_6200 = (n_66 & n_6199) ;
	assign n_6198 = (x_176 & n_60) ;
	assign n_6192 = (~x_177 & ~n_936) ;
	assign n_7835 = (~n_6220 & n_7834) ;
	assign n_6217 = (~n_6215 & ~n_6216) ;
	assign n_6210 = (~x_175 & ~n_6208) ;
	assign n_6209 = (x_175 & n_6208) ;
	assign n_6201 = (~n_6198 & ~n_6200) ;
	assign n_6193 = (i_5 & ~n_6192) ;
	assign n_6191 = (~i_33 & n_936) ;
	assign n_6185 = (~x_178 & ~n_697) ;
	assign n_6170 = (~x_180 & n_6) ;
	assign n_5727 = (~i_51 & ~n_6) ;
	assign n_6166 = (~x_337 & ~n_544) ;
	assign n_7836 = (~n_6217 & n_7835) ;
	assign n_6211 = (~n_6209 & ~n_6210) ;
	assign n_6203 = (~x_176 & n_6201) ;
	assign n_6202 = (x_176 & ~n_6201) ;
	assign n_6194 = (~n_6191 & n_6193) ;
	assign n_6186 = (i_5 & ~n_6185) ;
	assign n_6184 = (~x_683 & n_697) ;
	assign n_6171 = (~n_5727 & ~n_6170) ;
	assign n_6167 = (n_662 & ~n_6166) ;
	assign n_7837 = (~n_6211 & n_7836) ;
	assign n_6204 = (~n_6202 & ~n_6203) ;
	assign n_6196 = (~x_177 & ~n_6194) ;
	assign n_6195 = (x_177 & n_6194) ;
	assign n_6187 = (~n_6184 & n_6186) ;
	assign n_6179 = (x_376 & n_53) ;
	assign n_6178 = (x_179 & n_51) ;
	assign n_6172 = (n_629 & ~n_6171) ;
	assign n_6168 = (~n_629 & ~n_6167) ;
	assign n_6165 = (x_180 & ~n_662) ;
	assign n_7838 = (~n_6204 & n_7837) ;
	assign n_6197 = (~n_6195 & ~n_6196) ;
	assign n_6189 = (~x_178 & ~n_6187) ;
	assign n_6188 = (x_178 & n_6187) ;
	assign n_6180 = (~n_6178 & ~n_6179) ;
	assign n_6173 = (i_5 & ~n_6172) ;
	assign n_6169 = (~n_6165 & n_6168) ;
	assign n_7839 = (~n_6197 & n_7838) ;
	assign n_6190 = (~n_6188 & ~n_6189) ;
	assign n_6182 = (~x_179 & n_6180) ;
	assign n_6181 = (x_179 & ~n_6180) ;
	assign n_6174 = (~n_6169 & n_6173) ;
	assign n_6160 = (~n_143 & n_1009) ;
	assign n_6159 = (x_181 & n_1007) ;
	assign n_6153 = (~x_182 & ~n_630) ;
	assign n_7840 = (~n_6190 & n_7839) ;
	assign n_6183 = (~n_6181 & ~n_6182) ;
	assign n_6176 = (~x_180 & ~n_6174) ;
	assign n_6175 = (x_180 & n_6174) ;
	assign n_6161 = (~n_6159 & ~n_6160) ;
	assign n_6154 = (i_5 & ~n_6153) ;
	assign n_6152 = (~i_14 & n_630) ;
	assign n_6146 = (i_52 & n_64) ;
	assign n_7841 = (~n_6183 & n_7840) ;
	assign n_6177 = (~n_6175 & ~n_6176) ;
	assign n_6163 = (~x_181 & n_6161) ;
	assign n_6162 = (x_181 & ~n_6161) ;
	assign n_6155 = (~n_6152 & n_6154) ;
	assign n_6147 = (n_66 & n_6146) ;
	assign n_6145 = (x_183 & n_978) ;
	assign n_6139 = (~x_184 & ~n_936) ;
	assign n_7842 = (~n_6177 & n_7841) ;
	assign n_6164 = (~n_6162 & ~n_6163) ;
	assign n_6157 = (~x_182 & ~n_6155) ;
	assign n_6156 = (x_182 & n_6155) ;
	assign n_6148 = (~n_6145 & ~n_6147) ;
	assign n_6140 = (i_5 & ~n_6139) ;
	assign n_6138 = (~i_30 & n_936) ;
	assign n_6132 = (i_21 & n_64) ;
	assign n_7843 = (~n_6164 & n_7842) ;
	assign n_6158 = (~n_6156 & ~n_6157) ;
	assign n_6150 = (~x_183 & n_6148) ;
	assign n_6149 = (x_183 & ~n_6148) ;
	assign n_6141 = (~n_6138 & n_6140) ;
	assign n_6133 = (n_66 & n_6132) ;
	assign n_6131 = (x_185 & n_978) ;
	assign n_6125 = (~x_186 & ~n_697) ;
	assign n_7844 = (~n_6158 & n_7843) ;
	assign n_6151 = (~n_6149 & ~n_6150) ;
	assign n_6143 = (~x_184 & ~n_6141) ;
	assign n_6142 = (x_184 & n_6141) ;
	assign n_6134 = (~n_6131 & ~n_6133) ;
	assign n_6126 = (i_5 & ~n_6125) ;
	assign n_6124 = (~x_432 & n_697) ;
	assign n_7845 = (~n_6151 & n_7844) ;
	assign n_6144 = (~n_6142 & ~n_6143) ;
	assign n_6136 = (~x_185 & n_6134) ;
	assign n_6135 = (x_185 & ~n_6134) ;
	assign n_6127 = (~n_6124 & n_6126) ;
	assign n_6119 = (i_64 & n_948) ;
	assign n_6118 = (x_187 & n_945) ;
	assign n_7846 = (~n_6144 & n_7845) ;
	assign n_6137 = (~n_6135 & ~n_6136) ;
	assign n_6129 = (~x_186 & ~n_6127) ;
	assign n_6128 = (x_186 & n_6127) ;
	assign n_6120 = (~n_6118 & ~n_6119) ;
	assign n_6113 = (~n_407 & n_1009) ;
	assign n_6112 = (x_188 & n_1007) ;
	assign n_6106 = (i_51 & n_64) ;
	assign n_7847 = (~n_6137 & n_7846) ;
	assign n_6130 = (~n_6128 & ~n_6129) ;
	assign n_6122 = (~x_187 & n_6120) ;
	assign n_6121 = (x_187 & ~n_6120) ;
	assign n_6114 = (~n_6112 & ~n_6113) ;
	assign n_6107 = (n_66 & n_6106) ;
	assign n_6105 = (x_189 & n_978) ;
	assign n_6099 = (~x_190 & ~n_697) ;
	assign n_7848 = (~n_6130 & n_7847) ;
	assign n_6123 = (~n_6121 & ~n_6122) ;
	assign n_6116 = (~x_188 & n_6114) ;
	assign n_6115 = (x_188 & ~n_6114) ;
	assign n_6108 = (~n_6105 & ~n_6107) ;
	assign n_6100 = (i_5 & ~n_6099) ;
	assign n_6098 = (~x_699 & n_697) ;
	assign n_6092 = (~x_191 & ~n_936) ;
	assign n_7849 = (~n_6123 & n_7848) ;
	assign n_6117 = (~n_6115 & ~n_6116) ;
	assign n_6110 = (~x_189 & n_6108) ;
	assign n_6109 = (x_189 & ~n_6108) ;
	assign n_6101 = (~n_6098 & n_6100) ;
	assign n_6093 = (i_5 & ~n_6092) ;
	assign n_6091 = (~i_24 & n_936) ;
	assign n_7850 = (~n_6117 & n_7849) ;
	assign n_6111 = (~n_6109 & ~n_6110) ;
	assign n_6103 = (~x_190 & ~n_6101) ;
	assign n_6102 = (x_190 & n_6101) ;
	assign n_6094 = (~n_6091 & n_6093) ;
	assign n_6082 = (~x_193 & ~n_630) ;
	assign n_6026 = (~n_184 & ~n_185) ;
	assign n_7851 = (~n_6111 & n_7850) ;
	assign n_6104 = (~n_6102 & ~n_6103) ;
	assign n_6096 = (~x_191 & ~n_6094) ;
	assign n_6095 = (x_191 & n_6094) ;
	assign n_6083 = (i_5 & ~n_6082) ;
	assign n_6081 = (~i_60 & n_630) ;
	assign n_6028 = (~x_75 & ~n_6026) ;
	assign n_7852 = (~n_6104 & n_7851) ;
	assign n_6097 = (~n_6095 & ~n_6096) ;
	assign n_6089 = (~x_192 & n_421) ;
	assign n_6088 = (x_192 & ~n_421) ;
	assign n_6084 = (~n_6081 & n_6083) ;
	assign n_6076 = (x_683 & n_53) ;
	assign n_6075 = (x_194 & n_51) ;
	assign n_6069 = (i_10 & n_64) ;
	assign n_6029 = (~x_332 & ~n_6028) ;
	assign n_6027 = (x_75 & n_6026) ;
	assign n_7853 = (~n_6097 & n_7852) ;
	assign n_6090 = (~n_6088 & ~n_6089) ;
	assign n_6086 = (~x_193 & ~n_6084) ;
	assign n_6085 = (x_193 & n_6084) ;
	assign n_6077 = (~n_6075 & ~n_6076) ;
	assign n_6070 = (n_66 & n_6069) ;
	assign n_6068 = (x_195 & n_978) ;
	assign n_6062 = (~x_196 & ~n_936) ;
	assign n_3363 = (~i_59 & ~n_6) ;
	assign n_6030 = (~n_6027 & n_6029) ;
	assign n_6000 = (~x_427 & n_1936) ;
	assign n_5999 = (x_427 & ~n_1936) ;
	assign n_7854 = (~n_6090 & n_7853) ;
	assign n_6087 = (~n_6085 & ~n_6086) ;
	assign n_6079 = (~x_194 & n_6077) ;
	assign n_6078 = (x_194 & ~n_6077) ;
	assign n_6071 = (~n_6068 & ~n_6070) ;
	assign n_6063 = (i_5 & ~n_6062) ;
	assign n_6061 = (~i_15 & n_936) ;
	assign n_6055 = (~x_197 & ~n_544) ;
	assign n_6047 = (i_38 & n_669) ;
	assign n_6046 = (x_186 & n_662) ;
	assign n_6037 = (n_1 & ~n_3363) ;
	assign n_6036 = (n_6 & n_188) ;
	assign n_6032 = (n_188 & ~n_6030) ;
	assign n_6001 = (~n_5999 & ~n_6000) ;
	assign n_5998 = (~n_1926 & ~n_1927) ;
	assign n_7855 = (~n_6087 & n_7854) ;
	assign n_6080 = (~n_6078 & ~n_6079) ;
	assign n_6073 = (~x_195 & n_6071) ;
	assign n_6072 = (x_195 & ~n_6071) ;
	assign n_6064 = (~n_6061 & n_6063) ;
	assign n_6056 = (i_5 & ~n_6055) ;
	assign n_6054 = (~i_58 & n_544) ;
	assign n_6048 = (~n_6046 & ~n_6047) ;
	assign n_6045 = (x_198 & ~n_665) ;
	assign n_6038 = (~n_6036 & n_6037) ;
	assign n_6035 = (n_59 & ~n_188) ;
	assign n_6033 = (x_664 & ~n_6032) ;
	assign n_6031 = (~n_188 & n_6030) ;
	assign n_6010 = (i_36 & ~n_6) ;
	assign n_6003 = (n_5998 & ~n_6001) ;
	assign n_7856 = (~n_6080 & n_7855) ;
	assign n_6074 = (~n_6072 & ~n_6073) ;
	assign n_6066 = (~x_196 & ~n_6064) ;
	assign n_6065 = (x_196 & n_6064) ;
	assign n_6057 = (~n_6054 & n_6056) ;
	assign n_6049 = (~n_6045 & n_6048) ;
	assign n_6039 = (~n_6035 & ~n_6038) ;
	assign n_6034 = (~n_6031 & n_6033) ;
	assign n_6011 = (n_629 & ~n_6010) ;
	assign n_6009 = (x_201 & n_6) ;
	assign n_6006 = (x_201 & ~n_697) ;
	assign n_6004 = (n_697 & ~n_6003) ;
	assign n_6002 = (~n_5998 & n_6001) ;
	assign n_5967 = (~n_493 & ~n_494) ;
	assign n_7857 = (~n_6074 & n_7856) ;
	assign n_6067 = (~n_6065 & ~n_6066) ;
	assign n_6059 = (~x_197 & ~n_6057) ;
	assign n_6058 = (x_197 & n_6057) ;
	assign n_6050 = (i_5 & ~n_6049) ;
	assign n_6040 = (~n_6034 & n_6039) ;
	assign n_6020 = (i_14 & n_64) ;
	assign n_6012 = (~n_6009 & n_6011) ;
	assign n_6007 = (~n_629 & ~n_6006) ;
	assign n_6005 = (~n_6002 & n_6004) ;
	assign n_5969 = (~x_366 & ~n_5967) ;
	assign n_7858 = (~n_6067 & n_7857) ;
	assign n_6060 = (~n_6058 & ~n_6059) ;
	assign n_6052 = (~x_198 & ~n_6050) ;
	assign n_6051 = (x_198 & n_6050) ;
	assign n_6041 = (i_5 & ~n_6040) ;
	assign n_6021 = (n_66 & n_6020) ;
	assign n_6019 = (x_200 & n_978) ;
	assign n_6013 = (n_902 & ~n_6012) ;
	assign n_6008 = (~n_6005 & n_6007) ;
	assign n_5970 = (n_527 & ~n_5969) ;
	assign n_5968 = (x_366 & n_5967) ;
	assign n_7859 = (~n_6060 & n_7858) ;
	assign n_6053 = (~n_6051 & ~n_6052) ;
	assign n_6043 = (~x_199 & ~n_6041) ;
	assign n_6042 = (x_199 & n_6041) ;
	assign n_6022 = (~n_6019 & ~n_6021) ;
	assign n_6014 = (~n_6008 & n_6013) ;
	assign n_5997 = (x_201 & n_699) ;
	assign n_2901 = (~i_42 & ~n_6) ;
	assign n_5976 = (n_6 & n_497) ;
	assign n_5971 = (~n_5968 & n_5970) ;
	assign n_7860 = (~n_6053 & n_7859) ;
	assign n_6044 = (~n_6042 & ~n_6043) ;
	assign n_6024 = (~x_200 & n_6022) ;
	assign n_6023 = (x_200 & ~n_6022) ;
	assign n_6015 = (~n_5997 & ~n_6014) ;
	assign n_5992 = (~n_272 & n_1009) ;
	assign n_5991 = (x_202 & n_1007) ;
	assign n_5985 = (i_8 & n_59) ;
	assign n_5977 = (~n_5976 & ~n_2901) ;
	assign n_5973 = (n_497 & n_5971) ;
	assign n_7861 = (~n_6044 & n_7860) ;
	assign n_6025 = (~n_6023 & ~n_6024) ;
	assign n_6017 = (~x_201 & n_6015) ;
	assign n_6016 = (x_201 & ~n_6015) ;
	assign n_5993 = (~n_5991 & ~n_5992) ;
	assign n_5986 = (n_66 & n_5985) ;
	assign n_5984 = (x_203 & n_60) ;
	assign n_5978 = (n_1 & ~n_5977) ;
	assign n_5974 = (~n_1 & ~n_5973) ;
	assign n_5972 = (~n_497 & ~n_5971) ;
	assign n_7862 = (~n_6025 & n_7861) ;
	assign n_6018 = (~n_6016 & ~n_6017) ;
	assign n_5995 = (~x_202 & n_5993) ;
	assign n_5994 = (x_202 & ~n_5993) ;
	assign n_5987 = (~n_5984 & ~n_5986) ;
	assign n_5979 = (i_5 & ~n_5978) ;
	assign n_5975 = (~n_5972 & n_5974) ;
	assign n_7863 = (~n_6018 & n_7862) ;
	assign n_5996 = (~n_5994 & ~n_5995) ;
	assign n_5989 = (~x_203 & n_5987) ;
	assign n_5988 = (x_203 & ~n_5987) ;
	assign n_5980 = (~n_5975 & n_5979) ;
	assign n_5958 = (i_67 & n_59) ;
	assign n_5950 = (~i_7 & n_669) ;
	assign n_5948 = (~x_610 & ~n_544) ;
	assign n_5905 = (~n_343 & ~n_344) ;
	assign n_7864 = (~n_5996 & n_7863) ;
	assign n_5990 = (~n_5988 & ~n_5989) ;
	assign n_5982 = (~x_204 & ~n_5980) ;
	assign n_5981 = (x_204 & n_5980) ;
	assign n_5959 = (n_66 & n_5958) ;
	assign n_5957 = (x_206 & n_60) ;
	assign n_5951 = (i_5 & ~n_5950) ;
	assign n_5949 = (n_662 & n_5948) ;
	assign n_5907 = (~x_803 & ~n_5905) ;
	assign n_7865 = (~n_5990 & n_7864) ;
	assign n_5983 = (~n_5981 & ~n_5982) ;
	assign n_5965 = (~x_205 & n_272) ;
	assign n_5964 = (x_205 & ~n_272) ;
	assign n_5960 = (~n_5957 & ~n_5959) ;
	assign n_5952 = (~n_5949 & n_5951) ;
	assign n_5947 = (~x_207 & ~n_665) ;
	assign n_5908 = (~x_332 & ~n_5907) ;
	assign n_5906 = (x_803 & n_5905) ;
	assign n_7866 = (~n_5983 & n_7865) ;
	assign n_5966 = (~n_5964 & ~n_5965) ;
	assign n_5962 = (~x_206 & n_5960) ;
	assign n_5961 = (x_206 & ~n_5960) ;
	assign n_5953 = (~n_5947 & n_5952) ;
	assign n_5942 = (i_48 & n_948) ;
	assign n_5941 = (x_208 & n_945) ;
	assign n_5909 = (~n_5906 & n_5908) ;
	assign n_7867 = (~n_5966 & n_7866) ;
	assign n_5963 = (~n_5961 & ~n_5962) ;
	assign n_5955 = (~x_207 & ~n_5953) ;
	assign n_5954 = (x_207 & n_5953) ;
	assign n_5943 = (~n_5941 & ~n_5942) ;
	assign n_5936 = (~n_107 & n_35) ;
	assign n_5935 = (x_209 & n_36) ;
	assign n_5911 = (n_347 & ~n_5909) ;
	assign n_7868 = (~n_5963 & n_7867) ;
	assign n_5956 = (~n_5954 & ~n_5955) ;
	assign n_5945 = (~x_208 & n_5943) ;
	assign n_5944 = (x_208 & ~n_5943) ;
	assign n_5937 = (~n_5935 & ~n_5936) ;
	assign n_5930 = (x_627 & n_53) ;
	assign n_5929 = (x_210 & n_51) ;
	assign n_5923 = (~x_211 & ~n_630) ;
	assign n_5915 = (~n_347 & ~n_1606) ;
	assign n_5914 = (i_36 & n_7) ;
	assign n_5912 = (x_664 & ~n_5911) ;
	assign n_5910 = (~n_347 & n_5909) ;
	assign n_5866 = (~x_481 & n_2811) ;
	assign n_5865 = (x_481 & ~n_2811) ;
	assign n_7869 = (~n_5956 & n_7868) ;
	assign n_5946 = (~n_5944 & ~n_5945) ;
	assign n_5939 = (~x_209 & n_5937) ;
	assign n_5938 = (x_209 & ~n_5937) ;
	assign n_5931 = (~n_5929 & ~n_5930) ;
	assign n_5924 = (i_5 & ~n_5923) ;
	assign n_5922 = (~i_51 & n_630) ;
	assign n_5916 = (~n_5914 & ~n_5915) ;
	assign n_5913 = (~n_5910 & n_5912) ;
	assign n_5867 = (~n_5865 & ~n_5866) ;
	assign n_5864 = (~n_2802 & ~n_2801) ;
	assign n_7870 = (~n_5946 & n_7869) ;
	assign n_5940 = (~n_5938 & ~n_5939) ;
	assign n_5933 = (~x_210 & n_5931) ;
	assign n_5932 = (x_210 & ~n_5931) ;
	assign n_5925 = (~n_5922 & n_5924) ;
	assign n_5917 = (~n_5913 & n_5916) ;
	assign n_5899 = (i_52 & n_59) ;
	assign n_5875 = (~x_216 & n_6) ;
	assign n_1065 = (~i_17 & ~n_6) ;
	assign n_5869 = (n_5864 & ~n_5867) ;
	assign n_7871 = (~n_5940 & n_7870) ;
	assign n_5934 = (~n_5932 & ~n_5933) ;
	assign n_5927 = (~x_211 & ~n_5925) ;
	assign n_5926 = (x_211 & n_5925) ;
	assign n_5918 = (i_5 & ~n_5917) ;
	assign n_5900 = (n_66 & n_5899) ;
	assign n_5898 = (x_213 & n_60) ;
	assign n_5892 = (i_54 & n_64) ;
	assign n_5876 = (~n_1065 & ~n_5875) ;
	assign n_5872 = (x_216 & ~n_697) ;
	assign n_5870 = (n_697 & ~n_5869) ;
	assign n_5868 = (~n_5864 & n_5867) ;
	assign n_7872 = (~n_5934 & n_7871) ;
	assign n_5928 = (~n_5926 & ~n_5927) ;
	assign n_5920 = (~x_212 & ~n_5918) ;
	assign n_5919 = (x_212 & n_5918) ;
	assign n_5901 = (~n_5898 & ~n_5900) ;
	assign n_5893 = (n_66 & n_5892) ;
	assign n_5891 = (x_214 & n_978) ;
	assign n_5885 = (i_20 & n_59) ;
	assign n_5877 = (n_629 & ~n_5876) ;
	assign n_5873 = (~n_629 & ~n_5872) ;
	assign n_5871 = (~n_5868 & n_5870) ;
	assign n_5824 = (~x_810 & n_825) ;
	assign n_5823 = (x_810 & ~n_825) ;
	assign n_7873 = (~n_5928 & n_7872) ;
	assign n_5921 = (~n_5919 & ~n_5920) ;
	assign n_5903 = (~x_213 & n_5901) ;
	assign n_5902 = (x_213 & ~n_5901) ;
	assign n_5894 = (~n_5891 & ~n_5893) ;
	assign n_5886 = (n_66 & n_5885) ;
	assign n_5884 = (x_215 & n_60) ;
	assign n_5878 = (n_902 & ~n_5877) ;
	assign n_5874 = (~n_5871 & n_5873) ;
	assign n_5825 = (~n_5823 & ~n_5824) ;
	assign n_5822 = (~n_815 & ~n_816) ;
	assign n_7874 = (~n_5921 & n_7873) ;
	assign n_5904 = (~n_5902 & ~n_5903) ;
	assign n_5896 = (~x_214 & n_5894) ;
	assign n_5895 = (x_214 & ~n_5894) ;
	assign n_5887 = (~n_5884 & ~n_5886) ;
	assign n_5879 = (~n_5874 & n_5878) ;
	assign n_5863 = (x_216 & n_699) ;
	assign n_5834 = (~x_220 & n_6) ;
	assign n_5827 = (n_5822 & ~n_5825) ;
	assign n_7875 = (~n_5904 & n_7874) ;
	assign n_5897 = (~n_5895 & ~n_5896) ;
	assign n_5889 = (~x_215 & n_5887) ;
	assign n_5888 = (x_215 & ~n_5887) ;
	assign n_5880 = (~n_5863 & ~n_5879) ;
	assign n_5858 = (i_15 & n_948) ;
	assign n_5857 = (x_217 & n_945) ;
	assign n_5851 = (~x_218 & ~n_544) ;
	assign n_5835 = (~n_5833 & ~n_5834) ;
	assign n_5830 = (x_220 & ~n_697) ;
	assign n_5828 = (n_697 & ~n_5827) ;
	assign n_5826 = (~n_5822 & n_5825) ;
	assign n_7876 = (~n_5897 & n_7875) ;
	assign n_5890 = (~n_5888 & ~n_5889) ;
	assign n_5882 = (~x_216 & n_5880) ;
	assign n_5881 = (x_216 & ~n_5880) ;
	assign n_5859 = (~n_5857 & ~n_5858) ;
	assign n_5852 = (i_5 & ~n_5851) ;
	assign n_5850 = (~i_57 & n_544) ;
	assign n_5844 = (~x_219 & ~n_544) ;
	assign n_5836 = (n_629 & ~n_5835) ;
	assign n_5831 = (~n_629 & ~n_5830) ;
	assign n_5829 = (~n_5826 & n_5828) ;
	assign n_7877 = (~n_5890 & n_7876) ;
	assign n_5883 = (~n_5881 & ~n_5882) ;
	assign n_5861 = (~x_217 & n_5859) ;
	assign n_5860 = (x_217 & ~n_5859) ;
	assign n_5853 = (~n_5850 & n_5852) ;
	assign n_5845 = (i_5 & ~n_5844) ;
	assign n_5843 = (~i_6 & n_544) ;
	assign n_5837 = (n_902 & ~n_5836) ;
	assign n_5832 = (~n_5829 & n_5831) ;
	assign n_7878 = (~n_5883 & n_7877) ;
	assign n_5862 = (~n_5860 & ~n_5861) ;
	assign n_5855 = (~x_218 & ~n_5853) ;
	assign n_5854 = (x_218 & n_5853) ;
	assign n_5846 = (~n_5843 & n_5845) ;
	assign n_5838 = (~n_5832 & n_5837) ;
	assign n_5821 = (x_220 & n_699) ;
	assign n_7879 = (~n_5862 & n_7878) ;
	assign n_5856 = (~n_5854 & ~n_5855) ;
	assign n_5848 = (~x_219 & ~n_5846) ;
	assign n_5847 = (x_219 & n_5846) ;
	assign n_5839 = (~n_5821 & ~n_5838) ;
	assign n_5816 = (i_21 & n_948) ;
	assign n_5815 = (x_221 & n_945) ;
	assign n_5802 = (i_52 & n_7) ;
	assign n_5801 = (x_264 & ~n_16) ;
	assign n_7880 = (~n_5856 & n_7879) ;
	assign n_5849 = (~n_5847 & ~n_5848) ;
	assign n_5841 = (~x_220 & n_5839) ;
	assign n_5840 = (x_220 & ~n_5839) ;
	assign n_5817 = (~n_5815 & ~n_5816) ;
	assign n_5810 = (x_202 & n_35) ;
	assign n_5809 = (x_222 & n_36) ;
	assign n_5803 = (~n_5801 & ~n_5802) ;
	assign n_7881 = (~n_5849 & n_7880) ;
	assign n_5842 = (~n_5840 & ~n_5841) ;
	assign n_5819 = (~x_221 & n_5817) ;
	assign n_5818 = (x_221 & ~n_5817) ;
	assign n_5811 = (~n_5809 & ~n_5810) ;
	assign n_5804 = (n_20 & ~n_5803) ;
	assign n_5800 = (x_223 & n_18) ;
	assign n_5794 = (~x_224 & ~n_544) ;
	assign n_7882 = (~n_5842 & n_7881) ;
	assign n_5820 = (~n_5818 & ~n_5819) ;
	assign n_5813 = (~x_222 & n_5811) ;
	assign n_5812 = (x_222 & ~n_5811) ;
	assign n_5805 = (~n_5800 & ~n_5804) ;
	assign n_5795 = (i_5 & ~n_5794) ;
	assign n_5793 = (~i_64 & n_544) ;
	assign n_5787 = (~x_225 & ~n_697) ;
	assign n_5772 = (i_24 & n_1) ;
	assign n_5771 = (~x_227 & n_6) ;
	assign n_7883 = (~n_5820 & n_7882) ;
	assign n_5814 = (~n_5812 & ~n_5813) ;
	assign n_5807 = (~x_223 & n_5805) ;
	assign n_5806 = (x_223 & ~n_5805) ;
	assign n_5796 = (~n_5793 & n_5795) ;
	assign n_5788 = (i_5 & ~n_5787) ;
	assign n_5786 = (~x_436 & n_697) ;
	assign n_5773 = (~n_5771 & n_5772) ;
	assign n_5770 = (x_557 & ~n_16) ;
	assign n_5706 = (x_622 & ~x_640) ;
	assign n_5705 = (~x_765 & x_773) ;
	assign n_5703 = (x_765 & ~x_773) ;
	assign n_5702 = (x_605 & ~x_613) ;
	assign n_5699 = (x_186 & ~x_196) ;
	assign n_5698 = (~x_519 & x_576) ;
	assign n_5696 = (x_519 & ~x_576) ;
	assign n_5695 = (~x_622 & x_640) ;
	assign n_5691 = (x_715 & ~x_758) ;
	assign n_5690 = (~x_523 & x_539) ;
	assign n_5688 = (x_363 & ~x_451) ;
	assign n_5687 = (x_248 & ~x_307) ;
	assign n_5684 = (~x_480 & x_526) ;
	assign n_5683 = (~x_78 & x_91) ;
	assign n_5681 = (x_78 & ~x_91) ;
	assign n_5680 = (~x_715 & x_758) ;
	assign n_5675 = (~x_171 & x_178) ;
	assign n_5674 = (~x_112 & x_469) ;
	assign n_5672 = (x_617 & ~x_633) ;
	assign n_5671 = (x_70 & ~x_109) ;
	assign n_5668 = (x_529 & ~x_588) ;
	assign n_5667 = (~x_278 & x_299) ;
	assign n_5665 = (~x_387 & x_699) ;
	assign n_5664 = (x_166 & ~x_175) ;
	assign n_5660 = (~x_491 & x_806) ;
	assign n_5659 = (~x_286 & x_627) ;
	assign n_5657 = (~x_110 & x_124) ;
	assign n_5656 = (~x_135 & x_184) ;
	assign n_5653 = (x_302 & ~x_794) ;
	assign n_5652 = (~x_289 & x_330) ;
	assign n_5650 = (x_323 & ~x_727) ;
	assign n_5649 = (~x_585 & x_709) ;
	assign n_5643 = (x_118 & ~x_432) ;
	assign n_5642 = (x_112 & ~x_469) ;
	assign n_5640 = (x_476 & ~x_600) ;
	assign n_5639 = (x_258 & ~x_659) ;
	assign n_5636 = (x_480 & ~x_526) ;
	assign n_5635 = (x_225 & ~x_268) ;
	assign n_5633 = (x_161 & ~x_220) ;
	assign n_5632 = (~x_370 & x_778) ;
	assign n_5628 = (~x_397 & x_407) ;
	assign n_5627 = (x_397 & ~x_407) ;
	assign n_5625 = (x_339 & ~x_683) ;
	assign n_5624 = (x_289 & ~x_330) ;
	assign n_5621 = (~x_376 & x_711) ;
	assign n_5620 = (~x_339 & x_683) ;
	assign n_5618 = (~x_391 & x_442) ;
	assign n_5617 = (~x_312 & x_359) ;
	assign n_5612 = (x_585 & ~x_709) ;
	assign n_5611 = (x_416 & ~x_431) ;
	assign n_5609 = (x_191 & ~x_538) ;
	assign n_5608 = (x_704 & ~x_717) ;
	assign n_5605 = (~x_216 & x_560) ;
	assign n_5604 = (~x_248 & x_307) ;
	assign n_5602 = (x_324 & ~x_337) ;
	assign n_5601 = (~x_605 & x_613) ;
	assign n_5597 = (~x_558 & x_574) ;
	assign n_5596 = (x_387 & ~x_699) ;
	assign n_5594 = (~x_580 & x_738) ;
	assign n_5593 = (~x_379 & x_436) ;
	assign n_5590 = (~x_704 & x_717) ;
	assign n_5589 = (~x_225 & x_268) ;
	assign n_5587 = (~x_323 & x_727) ;
	assign n_5586 = (x_117 & ~x_666) ;
	assign n_7884 = (~n_5814 & n_7883) ;
	assign n_5808 = (~n_5806 & ~n_5807) ;
	assign n_5798 = (~x_224 & ~n_5796) ;
	assign n_5797 = (x_224 & n_5796) ;
	assign n_5789 = (~n_5786 & n_5788) ;
	assign n_5781 = (i_30 & n_948) ;
	assign n_5780 = (x_226 & n_945) ;
	assign n_5774 = (~n_5770 & ~n_5773) ;
	assign n_5769 = (x_227 & n_17) ;
	assign n_5707 = (~n_5705 & ~n_5706) ;
	assign n_5704 = (~n_5702 & ~n_5703) ;
	assign n_5700 = (~n_5698 & ~n_5699) ;
	assign n_5697 = (~n_5695 & ~n_5696) ;
	assign n_5692 = (~n_5690 & ~n_5691) ;
	assign n_5689 = (~n_5687 & ~n_5688) ;
	assign n_5685 = (~n_5683 & ~n_5684) ;
	assign n_5682 = (~n_5680 & ~n_5681) ;
	assign n_5676 = (~n_5674 & ~n_5675) ;
	assign n_5673 = (~n_5671 & ~n_5672) ;
	assign n_5669 = (~n_5667 & ~n_5668) ;
	assign n_5666 = (~n_5664 & ~n_5665) ;
	assign n_5661 = (~n_5659 & ~n_5660) ;
	assign n_5658 = (~n_5656 & ~n_5657) ;
	assign n_5654 = (~n_5652 & ~n_5653) ;
	assign n_5651 = (~n_5649 & ~n_5650) ;
	assign n_5644 = (~n_5642 & ~n_5643) ;
	assign n_5641 = (~n_5639 & ~n_5640) ;
	assign n_5637 = (~n_5635 & ~n_5636) ;
	assign n_5634 = (~n_5632 & ~n_5633) ;
	assign n_5629 = (~n_5627 & ~n_5628) ;
	assign n_5626 = (~n_5624 & ~n_5625) ;
	assign n_5622 = (~n_5620 & ~n_5621) ;
	assign n_5619 = (~n_5617 & ~n_5618) ;
	assign n_5613 = (~n_5611 & ~n_5612) ;
	assign n_5610 = (~n_5608 & ~n_5609) ;
	assign n_5606 = (~n_5604 & ~n_5605) ;
	assign n_5603 = (~n_5601 & ~n_5602) ;
	assign n_5598 = (~n_5596 & ~n_5597) ;
	assign n_5595 = (~n_5593 & ~n_5594) ;
	assign n_5591 = (~n_5589 & ~n_5590) ;
	assign n_5588 = (~n_5586 & ~n_5587) ;
	assign n_5580 = (x_247 & ~x_643) ;
	assign n_5579 = (x_491 & ~x_806) ;
	assign n_5577 = (x_320 & ~x_371) ;
	assign n_5576 = (x_201 & ~x_361) ;
	assign n_5573 = (x_458 & ~x_623) ;
	assign n_5572 = (x_379 & ~x_436) ;
	assign n_5570 = (~x_504 & x_795) ;
	assign n_5569 = (~x_191 & x_538) ;
	assign n_5565 = (~x_144 & x_270) ;
	assign n_5564 = (~x_161 & x_220) ;
	assign n_5561 = (~x_529 & x_588) ;
	assign n_5560 = (~x_117 & x_666) ;
	assign n_5558 = (x_420 & ~x_775) ;
	assign n_5557 = (~x_630 & x_677) ;
	assign n_5538 = (~x_476 & x_600) ;
	assign n_5537 = (~x_201 & x_361) ;
	assign n_5535 = (~x_617 & x_633) ;
	assign n_5534 = (x_110 & ~x_124) ;
	assign n_5531 = (~x_420 & x_775) ;
	assign n_5530 = (~x_166 & x_175) ;
	assign n_5528 = (~x_793 & x_802) ;
	assign n_5527 = (x_630 & ~x_677) ;
	assign n_5523 = (~x_70 & x_109) ;
	assign n_5522 = (x_370 & ~x_778) ;
	assign n_5520 = (x_278 & ~x_299) ;
	assign n_5519 = (~x_186 & x_196) ;
	assign n_5516 = (~x_320 & x_371) ;
	assign n_5515 = (x_286 & ~x_627) ;
	assign n_5513 = (~x_562 & x_610) ;
	assign n_5512 = (x_171 & ~x_178) ;
	assign n_5507 = (x_562 & ~x_610) ;
	assign n_5506 = (x_177 & ~x_190) ;
	assign n_5504 = (x_523 & ~x_539) ;
	assign n_5503 = (x_558 & ~x_574) ;
	assign n_5500 = (~x_230 & x_567) ;
	assign n_5499 = (~x_302 & x_794) ;
	assign n_5497 = (~x_416 & x_431) ;
	assign n_5496 = (~x_177 & x_190) ;
	assign n_5492 = (~x_447 & x_502) ;
	assign n_5491 = (x_391 & ~x_442) ;
	assign n_5489 = (x_376 & ~x_711) ;
	assign n_5488 = (x_216 & ~x_560) ;
	assign n_5485 = (~x_258 & x_659) ;
	assign n_5484 = (x_144 & ~x_270) ;
	assign n_5482 = (~x_363 & x_451) ;
	assign n_5481 = (~x_324 & x_337) ;
	assign n_7885 = (~n_5808 & n_7884) ;
	assign n_5799 = (~n_5797 & ~n_5798) ;
	assign n_5791 = (~x_225 & ~n_5789) ;
	assign n_5790 = (x_225 & n_5789) ;
	assign n_5782 = (~n_5780 & ~n_5781) ;
	assign n_5775 = (~n_5769 & n_5774) ;
	assign n_5708 = (n_5704 & n_5707) ;
	assign n_5701 = (n_5697 & n_5700) ;
	assign n_5693 = (n_5689 & n_5692) ;
	assign n_5686 = (n_5682 & n_5685) ;
	assign n_5677 = (n_5673 & n_5676) ;
	assign n_5670 = (n_5666 & n_5669) ;
	assign n_5662 = (n_5658 & n_5661) ;
	assign n_5655 = (n_5651 & n_5654) ;
	assign n_5645 = (n_5641 & n_5644) ;
	assign n_5638 = (n_5634 & n_5637) ;
	assign n_5630 = (n_5626 & n_5629) ;
	assign n_5623 = (n_5619 & n_5622) ;
	assign n_5614 = (n_5610 & n_5613) ;
	assign n_5607 = (n_5603 & n_5606) ;
	assign n_5599 = (n_5595 & n_5598) ;
	assign n_5592 = (n_5588 & n_5591) ;
	assign n_5581 = (~n_5579 & ~n_5580) ;
	assign n_5578 = (~n_5576 & ~n_5577) ;
	assign n_5574 = (~n_5572 & ~n_5573) ;
	assign n_5571 = (~n_5569 & ~n_5570) ;
	assign n_5566 = (~n_5564 & ~n_5565) ;
	assign n_5562 = (~n_5560 & ~n_5561) ;
	assign n_5559 = (~n_5557 & ~n_5558) ;
	assign n_5553 = (x_477 & x_486) ;
	assign n_5552 = (~x_477 & ~x_486) ;
	assign n_5550 = (x_259 & x_275) ;
	assign n_5549 = (~x_259 & ~x_275) ;
	assign n_5546 = (x_354 & x_465) ;
	assign n_5545 = (~x_354 & ~x_465) ;
	assign n_5539 = (~n_5537 & ~n_5538) ;
	assign n_5536 = (~n_5534 & ~n_5535) ;
	assign n_5532 = (~n_5530 & ~n_5531) ;
	assign n_5529 = (~n_5527 & ~n_5528) ;
	assign n_5524 = (~n_5522 & ~n_5523) ;
	assign n_5521 = (~n_5519 & ~n_5520) ;
	assign n_5517 = (~n_5515 & ~n_5516) ;
	assign n_5514 = (~n_5512 & ~n_5513) ;
	assign n_5508 = (~n_5506 & ~n_5507) ;
	assign n_5505 = (~n_5503 & ~n_5504) ;
	assign n_5501 = (~n_5499 & ~n_5500) ;
	assign n_5498 = (~n_5496 & ~n_5497) ;
	assign n_5493 = (~n_5491 & ~n_5492) ;
	assign n_5490 = (~n_5488 & ~n_5489) ;
	assign n_5486 = (~n_5484 & ~n_5485) ;
	assign n_5483 = (~n_5481 & ~n_5482) ;
	assign n_5476 = (x_793 & ~x_802) ;
	assign n_5475 = (x_441 & ~x_493) ;
	assign n_5473 = (~x_458 & x_623) ;
	assign n_5472 = (~x_441 & x_493) ;
	assign n_5468 = (x_504 & ~x_795) ;
	assign n_5467 = (x_580 & ~x_738) ;
	assign n_5465 = (~x_118 & x_432) ;
	assign n_5464 = (x_312 & ~x_359) ;
	assign n_5461 = (x_230 & ~x_567) ;
	assign n_5460 = (x_135 & ~x_184) ;
	assign n_5458 = (~x_247 & x_643) ;
	assign n_5457 = (x_447 & ~x_502) ;
	assign n_7886 = (~n_5799 & n_7885) ;
	assign n_5792 = (~n_5790 & ~n_5791) ;
	assign n_5784 = (~x_226 & n_5782) ;
	assign n_5783 = (x_226 & ~n_5782) ;
	assign n_5776 = (i_5 & ~n_5775) ;
	assign n_5760 = (i_62 & n_59) ;
	assign n_5736 = (x_232 & ~n_14) ;
	assign n_5709 = (n_5701 & n_5708) ;
	assign n_5694 = (n_5686 & n_5693) ;
	assign n_5678 = (n_5670 & n_5677) ;
	assign n_5663 = (n_5655 & n_5662) ;
	assign n_5646 = (n_5638 & n_5645) ;
	assign n_5631 = (n_5623 & n_5630) ;
	assign n_5615 = (n_5607 & n_5614) ;
	assign n_5600 = (n_5592 & n_5599) ;
	assign n_5582 = (n_5578 & n_5581) ;
	assign n_5575 = (n_5571 & n_5574) ;
	assign n_5567 = (n_43 & n_5566) ;
	assign n_5563 = (n_5559 & n_5562) ;
	assign n_5554 = (~n_5552 & ~n_5553) ;
	assign n_5551 = (~n_5549 & ~n_5550) ;
	assign n_5547 = (~n_5545 & ~n_5546) ;
	assign n_5540 = (n_5536 & n_5539) ;
	assign n_5533 = (n_5529 & n_5532) ;
	assign n_5525 = (n_5521 & n_5524) ;
	assign n_5518 = (n_5514 & n_5517) ;
	assign n_5509 = (n_5505 & n_5508) ;
	assign n_5502 = (n_5498 & n_5501) ;
	assign n_5494 = (n_5490 & n_5493) ;
	assign n_5487 = (n_5483 & n_5486) ;
	assign n_5477 = (~n_5475 & ~n_5476) ;
	assign n_5474 = (~n_5472 & ~n_5473) ;
	assign n_5469 = (~n_5467 & ~n_5468) ;
	assign n_5466 = (~n_5464 & ~n_5465) ;
	assign n_5462 = (~n_5460 & ~n_5461) ;
	assign n_5459 = (~n_5457 & ~n_5458) ;
	assign n_7887 = (~n_5792 & n_7886) ;
	assign n_5785 = (~n_5783 & ~n_5784) ;
	assign n_5778 = (~x_227 & ~n_5776) ;
	assign n_5777 = (x_227 & n_5776) ;
	assign n_5761 = (n_66 & n_5760) ;
	assign n_5759 = (x_229 & n_60) ;
	assign n_5753 = (~x_230 & ~n_936) ;
	assign n_5737 = (n_12 & ~n_5736) ;
	assign n_5735 = (x_631 & n_14) ;
	assign n_5732 = (x_631 & n_11) ;
	assign n_5710 = (n_5694 & n_5709) ;
	assign n_5679 = (n_5663 & n_5678) ;
	assign n_5647 = (n_5631 & n_5646) ;
	assign n_5616 = (n_5600 & n_5615) ;
	assign n_5583 = (n_5575 & n_5582) ;
	assign n_5568 = (n_5563 & n_5567) ;
	assign n_5555 = (~n_5551 & ~n_5554) ;
	assign n_5548 = (n_45 & ~n_5547) ;
	assign n_5541 = (n_5533 & n_5540) ;
	assign n_5526 = (n_5518 & n_5525) ;
	assign n_5510 = (n_5502 & n_5509) ;
	assign n_5495 = (n_5487 & n_5494) ;
	assign n_5478 = (n_5474 & n_5477) ;
	assign n_1820 = (n_43 & n_45) ;
	assign n_5470 = (n_5466 & n_5469) ;
	assign n_5463 = (n_5459 & n_5462) ;
	assign n_7888 = (~n_5785 & n_7887) ;
	assign n_5779 = (~n_5777 & ~n_5778) ;
	assign n_5767 = (~x_228 & n_376) ;
	assign n_5766 = (x_228 & ~n_376) ;
	assign n_5762 = (~n_5759 & ~n_5761) ;
	assign n_5754 = (i_5 & ~n_5753) ;
	assign n_5752 = (~i_64 & n_936) ;
	assign n_5746 = (~x_231 & ~n_544) ;
	assign n_5738 = (~n_5735 & n_5737) ;
	assign n_5733 = (x_168 & ~n_5732) ;
	assign n_5731 = (x_232 & ~n_11) ;
	assign n_5728 = (~x_232 & n_6) ;
	assign n_5711 = (n_5679 & n_5710) ;
	assign n_5648 = (n_5616 & n_5647) ;
	assign n_5584 = (n_5568 & n_5583) ;
	assign n_5556 = (n_5548 & n_5555) ;
	assign n_5542 = (n_5526 & n_5541) ;
	assign n_5511 = (n_5495 & n_5510) ;
	assign n_5479 = (n_1820 & n_5478) ;
	assign n_5471 = (n_5463 & n_5470) ;
	assign n_7889 = (~n_5779 & n_7888) ;
	assign n_5768 = (~n_5766 & ~n_5767) ;
	assign n_5764 = (~x_229 & n_5762) ;
	assign n_5763 = (x_229 & ~n_5762) ;
	assign n_5755 = (~n_5752 & n_5754) ;
	assign n_5747 = (i_5 & ~n_5746) ;
	assign n_5745 = (~i_10 & n_544) ;
	assign n_5739 = (i_5 & ~n_5738) ;
	assign n_5734 = (~n_5731 & n_5733) ;
	assign n_5729 = (~n_5727 & ~n_5728) ;
	assign n_5712 = (n_5648 & n_5711) ;
	assign n_5585 = (n_5556 & n_5584) ;
	assign n_5543 = (n_5511 & n_5542) ;
	assign n_5480 = (n_5471 & n_5479) ;
	assign n_7890 = (~n_5768 & n_7889) ;
	assign n_5765 = (~n_5763 & ~n_5764) ;
	assign n_5757 = (~x_230 & ~n_5755) ;
	assign n_5756 = (x_230 & n_5755) ;
	assign n_5748 = (~n_5745 & n_5747) ;
	assign n_5740 = (~n_5734 & n_5739) ;
	assign n_5730 = (n_1 & ~n_5729) ;
	assign n_5721 = (~x_233 & ~n_544) ;
	assign n_5713 = (n_5585 & n_5712) ;
	assign n_5544 = (n_5480 & n_5543) ;
	assign n_7891 = (~n_5765 & n_7890) ;
	assign n_5758 = (~n_5756 & ~n_5757) ;
	assign n_5750 = (~x_231 & ~n_5748) ;
	assign n_5749 = (x_231 & n_5748) ;
	assign n_5741 = (~n_5730 & n_5740) ;
	assign n_5722 = (i_5 & ~n_5721) ;
	assign n_5720 = (~i_20 & n_544) ;
	assign n_5714 = (n_5544 & n_5713) ;
	assign n_5456 = (x_234 & ~n_1820) ;
	assign n_7892 = (~n_5758 & n_7891) ;
	assign n_5751 = (~n_5749 & ~n_5750) ;
	assign n_5743 = (~x_232 & ~n_5741) ;
	assign n_5742 = (x_232 & n_5741) ;
	assign n_5723 = (~n_5720 & n_5722) ;
	assign n_5715 = (~n_5456 & ~n_5714) ;
	assign n_7893 = (~n_5751 & n_7892) ;
	assign n_5744 = (~n_5742 & ~n_5743) ;
	assign n_5725 = (~x_233 & ~n_5723) ;
	assign n_5724 = (x_233 & n_5723) ;
	assign n_5716 = (i_5 & ~n_5715) ;
	assign n_5451 = (i_60 & n_948) ;
	assign n_5450 = (x_235 & n_945) ;
	assign n_5444 = (i_6 & n_59) ;
	assign n_7894 = (~n_5744 & n_7893) ;
	assign n_5726 = (~n_5724 & ~n_5725) ;
	assign n_5718 = (~x_234 & ~n_5716) ;
	assign n_5717 = (x_234 & n_5716) ;
	assign n_5452 = (~n_5450 & ~n_5451) ;
	assign n_5445 = (n_66 & n_5444) ;
	assign n_5443 = (x_236 & n_60) ;
	assign n_7895 = (~n_5726 & n_7894) ;
	assign n_5719 = (~n_5717 & ~n_5718) ;
	assign n_5454 = (~x_235 & n_5452) ;
	assign n_5453 = (x_235 & ~n_5452) ;
	assign n_5446 = (~n_5443 & ~n_5445) ;
	assign n_5438 = (x_113 & n_35) ;
	assign n_5437 = (x_237 & n_36) ;
	assign n_7896 = (~n_5719 & n_7895) ;
	assign n_5455 = (~n_5453 & ~n_5454) ;
	assign n_5448 = (~x_236 & n_5446) ;
	assign n_5447 = (x_236 & ~n_5446) ;
	assign n_5439 = (~n_5437 & ~n_5438) ;
	assign n_5432 = (n_35 & ~n_511) ;
	assign n_5431 = (x_238 & n_36) ;
	assign n_1570 = (i_49 & n_64) ;
	assign n_7897 = (~n_5455 & n_7896) ;
	assign n_5449 = (~n_5447 & ~n_5448) ;
	assign n_5441 = (~x_237 & n_5439) ;
	assign n_5440 = (x_237 & ~n_5439) ;
	assign n_5433 = (~n_5431 & ~n_5432) ;
	assign n_1571 = (n_66 & n_1570) ;
	assign n_1569 = (x_239 & n_978) ;
	assign n_7898 = (~n_5449 & n_7897) ;
	assign n_5442 = (~n_5440 & ~n_5441) ;
	assign n_5435 = (~x_238 & n_5433) ;
	assign n_5434 = (x_238 & ~n_5433) ;
	assign n_1572 = (~n_1569 & ~n_1571) ;
	assign n_74 = (x_240 & ~x_527) ;
	assign n_73 = (x_527 & x_819) ;
	assign n_7899 = (~n_5442 & n_7898) ;
	assign n_5436 = (~n_5434 & ~n_5435) ;
	assign n_5429 = (~x_239 & n_1572) ;
	assign n_5428 = (x_239 & ~n_1572) ;
	assign n_75 = (~n_73 & ~n_74) ;
	assign n_5420 = (i_27 & n_948) ;
	assign n_5419 = (x_241 & n_945) ;
	assign n_5369 = (~x_722 & n_838) ;
	assign n_5368 = (x_722 & ~n_838) ;
	assign n_7900 = (~n_5436 & n_7899) ;
	assign n_5430 = (~n_5428 & ~n_5429) ;
	assign n_5426 = (~x_240 & n_75) ;
	assign n_5425 = (x_240 & ~n_75) ;
	assign n_5421 = (~n_5419 & ~n_5420) ;
	assign n_5414 = (x_363 & n_53) ;
	assign n_5413 = (x_242 & n_51) ;
	assign n_5370 = (~n_5368 & ~n_5369) ;
	assign n_5367 = (~n_828 & ~n_829) ;
	assign n_7901 = (~n_5430 & n_7900) ;
	assign n_5427 = (~n_5425 & ~n_5426) ;
	assign n_5423 = (~x_241 & n_5421) ;
	assign n_5422 = (x_241 & ~n_5421) ;
	assign n_5415 = (~n_5413 & ~n_5414) ;
	assign n_5408 = (i_19 & n_948) ;
	assign n_5407 = (x_243 & n_945) ;
	assign n_5379 = (i_32 & ~n_6) ;
	assign n_5372 = (n_5367 & ~n_5370) ;
	assign n_7902 = (~n_5427 & n_7901) ;
	assign n_5424 = (~n_5422 & ~n_5423) ;
	assign n_5417 = (~x_242 & n_5415) ;
	assign n_5416 = (x_242 & ~n_5415) ;
	assign n_5409 = (~n_5407 & ~n_5408) ;
	assign n_5402 = (x_135 & n_53) ;
	assign n_5401 = (x_244 & n_51) ;
	assign n_5380 = (n_629 & ~n_5379) ;
	assign n_5378 = (x_247 & n_6) ;
	assign n_5375 = (x_247 & ~n_697) ;
	assign n_5373 = (n_697 & ~n_5372) ;
	assign n_5371 = (~n_5367 & n_5370) ;
	assign n_7903 = (~n_5424 & n_7902) ;
	assign n_5418 = (~n_5416 & ~n_5417) ;
	assign n_5411 = (~x_243 & n_5409) ;
	assign n_5410 = (x_243 & ~n_5409) ;
	assign n_5403 = (~n_5401 & ~n_5402) ;
	assign n_5396 = (n_35 & ~n_75) ;
	assign n_5395 = (x_245 & n_36) ;
	assign n_5389 = (~x_246 & ~n_630) ;
	assign n_5381 = (~n_5378 & n_5380) ;
	assign n_5376 = (~n_629 & ~n_5375) ;
	assign n_5374 = (~n_5371 & n_5373) ;
	assign n_7904 = (~n_5418 & n_7903) ;
	assign n_5412 = (~n_5410 & ~n_5411) ;
	assign n_5405 = (~x_244 & n_5403) ;
	assign n_5404 = (x_244 & ~n_5403) ;
	assign n_5397 = (~n_5395 & ~n_5396) ;
	assign n_5390 = (i_5 & ~n_5389) ;
	assign n_5388 = (~i_8 & n_630) ;
	assign n_5382 = (n_902 & ~n_5381) ;
	assign n_5377 = (~n_5374 & n_5376) ;
	assign n_7905 = (~n_5412 & n_7904) ;
	assign n_5406 = (~n_5404 & ~n_5405) ;
	assign n_5399 = (~x_245 & n_5397) ;
	assign n_5398 = (x_245 & ~n_5397) ;
	assign n_5391 = (~n_5388 & n_5390) ;
	assign n_5383 = (~n_5377 & n_5382) ;
	assign n_5366 = (x_247 & n_699) ;
	assign n_5360 = (~x_248 & ~n_936) ;
	assign n_5352 = (~i_37 & n_669) ;
	assign n_7906 = (~n_5406 & n_7905) ;
	assign n_5400 = (~n_5398 & ~n_5399) ;
	assign n_5393 = (~x_246 & ~n_5391) ;
	assign n_5392 = (x_246 & n_5391) ;
	assign n_5384 = (~n_5366 & ~n_5383) ;
	assign n_5361 = (i_5 & ~n_5360) ;
	assign n_5359 = (~i_22 & n_936) ;
	assign n_5353 = (i_5 & ~n_5352) ;
	assign n_5351 = (~x_275 & n_662) ;
	assign n_7907 = (~n_5400 & n_7906) ;
	assign n_5394 = (~n_5392 & ~n_5393) ;
	assign n_5386 = (~x_247 & n_5384) ;
	assign n_5385 = (x_247 & ~n_5384) ;
	assign n_5362 = (~n_5359 & n_5361) ;
	assign n_5354 = (~n_5351 & n_5353) ;
	assign n_5350 = (~x_249 & ~n_665) ;
	assign n_5344 = (~x_250 & ~n_630) ;
	assign n_7908 = (~n_5394 & n_7907) ;
	assign n_5387 = (~n_5385 & ~n_5386) ;
	assign n_5364 = (~x_248 & ~n_5362) ;
	assign n_5363 = (x_248 & n_5362) ;
	assign n_5355 = (~n_5350 & n_5354) ;
	assign n_5345 = (i_5 & ~n_5344) ;
	assign n_5343 = (~i_52 & n_630) ;
	assign n_5337 = (~x_251 & ~n_630) ;
	assign n_1539 = (~x_168 & n_1538) ;
	assign n_1543 = (~n_59 & ~n_527) ;
	assign n_7909 = (~n_5387 & n_7908) ;
	assign n_5365 = (~n_5363 & ~n_5364) ;
	assign n_5357 = (~x_249 & ~n_5355) ;
	assign n_5356 = (x_249 & n_5355) ;
	assign n_5346 = (~n_5343 & n_5345) ;
	assign n_5338 = (i_5 & ~n_5337) ;
	assign n_5336 = (~i_24 & n_630) ;
	assign n_5330 = (i_7 & n_64) ;
	assign n_1546 = (x_578 & n_1539) ;
	assign n_1544 = (~n_1542 & n_1543) ;
	assign n_1222 = (x_308 & ~x_527) ;
	assign n_1221 = (x_527 & x_767) ;
	assign n_7910 = (~n_5365 & n_7909) ;
	assign n_5358 = (~n_5356 & ~n_5357) ;
	assign n_5348 = (~x_250 & ~n_5346) ;
	assign n_5347 = (x_250 & n_5346) ;
	assign n_5339 = (~n_5336 & n_5338) ;
	assign n_5331 = (n_66 & n_5330) ;
	assign n_5329 = (x_252 & n_978) ;
	assign n_1547 = (~n_944 & ~n_1546) ;
	assign n_1545 = (x_255 & ~n_1544) ;
	assign n_1540 = (~n_11 & ~n_1539) ;
	assign n_1223 = (~n_1221 & ~n_1222) ;
	assign n_5153 = (~x_463 & x_801) ;
	assign n_5152 = (~x_313 & x_779) ;
	assign n_5147 = (~x_389 & x_626) ;
	assign n_5146 = (~x_273 & x_419) ;
	assign n_5144 = (~x_272 & x_736) ;
	assign n_5143 = (~x_139 & x_485) ;
	assign n_5140 = (x_463 & ~x_801) ;
	assign n_5139 = (x_74 & ~x_429) ;
	assign n_5137 = (x_254 & ~x_537) ;
	assign n_5136 = (~x_575 & x_737) ;
	assign n_5123 = (~x_97 & x_294) ;
	assign n_5122 = (x_575 & ~x_737) ;
	assign n_5120 = (x_139 & ~x_485) ;
	assign n_5119 = (~x_113 & x_584) ;
	assign n_5116 = (~x_328 & x_673) ;
	assign n_5115 = (x_170 & ~x_631) ;
	assign n_5113 = (x_328 & ~x_673) ;
	assign n_5112 = (~x_170 & x_631) ;
	assign n_5108 = (~x_418 & x_713) ;
	assign n_5107 = (~x_127 & x_352) ;
	assign n_5105 = (~x_217 & x_408) ;
	assign n_5104 = (x_217 & ~x_408) ;
	assign n_5101 = (~x_264 & x_607) ;
	assign n_5100 = (x_273 & ~x_419) ;
	assign n_5098 = (x_188 & ~x_471) ;
	assign n_5097 = (~x_181 & x_521) ;
	assign n_5092 = (x_113 & ~x_584) ;
	assign n_5091 = (x_264 & ~x_607) ;
	assign n_5089 = (x_418 & ~x_713) ;
	assign n_5088 = (~x_283 & x_557) ;
	assign n_5085 = (~x_322 & x_712) ;
	assign n_5084 = (x_487 & ~x_656) ;
	assign n_5082 = (~x_341 & x_614) ;
	assign n_5081 = (x_341 & ~x_614) ;
	assign n_5077 = (x_389 & ~x_626) ;
	assign n_5076 = (~x_487 & x_656) ;
	assign n_5074 = (~x_188 & x_471) ;
	assign n_5073 = (x_283 & ~x_557) ;
	assign n_5070 = (x_81 & ~x_547) ;
	assign n_5069 = (x_127 & ~x_352) ;
	assign n_5067 = (~x_81 & x_547) ;
	assign n_5066 = (~x_235 & x_792) ;
	assign n_7911 = (~n_5358 & n_7910) ;
	assign n_5349 = (~n_5347 & ~n_5348) ;
	assign n_5341 = (~x_251 & ~n_5339) ;
	assign n_5340 = (x_251 & n_5339) ;
	assign n_5332 = (~n_5329 & ~n_5331) ;
	assign n_5324 = (x_289 & n_53) ;
	assign n_5323 = (x_253 & n_51) ;
	assign n_1548 = (~n_1545 & n_1547) ;
	assign n_1541 = (~x_255 & ~n_1540) ;
	assign n_5273 = (x_743 & n_188) ;
	assign n_5272 = (~x_596 & ~n_407) ;
	assign n_5270 = (~x_509 & ~n_511) ;
	assign n_5269 = (~x_85 & ~n_302) ;
	assign n_5266 = (~x_771 & ~n_317) ;
	assign n_5265 = (~x_533 & ~n_452) ;
	assign n_5263 = (~x_208 & ~n_362) ;
	assign n_5262 = (~x_439 & ~n_497) ;
	assign n_5258 = (~x_243 & ~n_242) ;
	assign n_5257 = (x_304 & n_436) ;
	assign n_5255 = (x_680 & n_392) ;
	assign n_5254 = (~x_660 & ~n_107) ;
	assign n_5251 = (x_357 & n_482) ;
	assign n_5250 = (x_596 & n_407) ;
	assign n_5248 = (x_88 & n_203) ;
	assign n_5247 = (~x_153 & ~n_376) ;
	assign n_5242 = (x_797 & n_86) ;
	assign n_5241 = (x_661 & n_272) ;
	assign n_5239 = (~x_747 & ~n_287) ;
	assign n_5238 = (~x_461 & ~n_75) ;
	assign n_5235 = (x_509 & n_511) ;
	assign n_5234 = (x_660 & n_107) ;
	assign n_5232 = (x_594 & n_227) ;
	assign n_5231 = (x_692 & n_332) ;
	assign n_5218 = (~x_772 & ~n_218) ;
	assign n_5217 = (~x_357 & ~n_482) ;
	assign n_5215 = (x_158 & n_257) ;
	assign n_5214 = (x_772 & n_218) ;
	assign n_5211 = (x_461 & n_75) ;
	assign n_5210 = (~x_158 & ~n_257) ;
	assign n_5208 = (x_156 & n_179) ;
	assign n_5207 = (~x_88 & ~n_203) ;
	assign n_5203 = (~x_797 & ~n_86) ;
	assign n_5202 = (x_85 & n_302) ;
	assign n_5200 = (x_365 & n_1223) ;
	assign n_5199 = (x_435 & n_139) ;
	assign n_5196 = (~x_692 & ~n_332) ;
	assign n_5195 = (~x_594 & ~n_227) ;
	assign n_5193 = (x_771 & n_317) ;
	assign n_5192 = (~x_119 & ~n_347) ;
	assign n_5187 = (~x_221 & ~n_421) ;
	assign n_5186 = (~x_661 & ~n_272) ;
	assign n_5184 = (~x_304 & ~n_436) ;
	assign n_5183 = (~x_505 & ~n_143) ;
	assign n_5180 = (x_153 & n_376) ;
	assign n_5179 = (~x_743 & ~n_188) ;
	assign n_5177 = (~x_449 & ~n_467) ;
	assign n_5176 = (~x_365 & ~n_1223) ;
	assign n_5172 = (~x_241 & ~n_164) ;
	assign n_5171 = (~x_435 & ~n_139) ;
	assign n_5169 = (x_241 & n_164) ;
	assign n_5168 = (x_321 & n_136) ;
	assign n_5165 = (x_505 & n_143) ;
	assign n_5164 = (x_221 & n_421) ;
	assign n_5162 = (~x_321 & ~n_136) ;
	assign n_5161 = (x_243 & n_242) ;
	assign n_5154 = (~n_5152 & ~n_5153) ;
	assign n_5151 = (x_202 & ~x_665) ;
	assign n_5148 = (~n_5146 & ~n_5147) ;
	assign n_5145 = (~n_5143 & ~n_5144) ;
	assign n_5141 = (~n_5139 & ~n_5140) ;
	assign n_5138 = (~n_5136 & ~n_5137) ;
	assign n_5124 = (~n_5122 & ~n_5123) ;
	assign n_5121 = (~n_5119 & ~n_5120) ;
	assign n_5117 = (~n_5115 & ~n_5116) ;
	assign n_5114 = (~n_5112 & ~n_5113) ;
	assign n_5109 = (~n_5107 & ~n_5108) ;
	assign n_5106 = (~n_5104 & ~n_5105) ;
	assign n_5102 = (~n_5100 & ~n_5101) ;
	assign n_5099 = (~n_5097 & ~n_5098) ;
	assign n_5093 = (~n_5091 & ~n_5092) ;
	assign n_5090 = (~n_5088 & ~n_5089) ;
	assign n_5086 = (~n_5084 & ~n_5085) ;
	assign n_5083 = (~n_5081 & ~n_5082) ;
	assign n_5078 = (~n_5076 & ~n_5077) ;
	assign n_5075 = (~n_5073 & ~n_5074) ;
	assign n_5071 = (~n_5069 & ~n_5070) ;
	assign n_5068 = (~n_5066 & ~n_5067) ;
	assign n_5060 = (x_181 & ~x_521) ;
	assign n_5059 = (~x_102 & x_394) ;
	assign n_5057 = (x_272 & ~x_736) ;
	assign n_5056 = (~x_202 & x_665) ;
	assign n_5053 = (x_97 & ~x_294) ;
	assign n_5052 = (~x_254 & x_537) ;
	assign n_5050 = (x_187 & ~x_350) ;
	assign n_5049 = (x_401 & ~x_757) ;
	assign n_5045 = (x_313 & ~x_779) ;
	assign n_5044 = (~x_90 & x_513) ;
	assign n_5042 = (x_355 & ~x_644) ;
	assign n_5041 = (~x_355 & x_644) ;
	assign n_5038 = (x_102 & ~x_394) ;
	assign n_5037 = (~x_401 & x_757) ;
	assign n_5035 = (~x_74 & x_429) ;
	assign n_5034 = (~x_187 & x_350) ;
	assign n_7912 = (~n_5349 & n_7911) ;
	assign n_5342 = (~n_5340 & ~n_5341) ;
	assign n_5334 = (~x_252 & n_5332) ;
	assign n_5333 = (x_252 & ~n_5332) ;
	assign n_5325 = (~n_5323 & ~n_5324) ;
	assign n_5318 = (n_1009 & ~n_452) ;
	assign n_5317 = (x_254 & n_1007) ;
	assign n_1549 = (~n_1541 & n_1548) ;
	assign n_5274 = (~n_5272 & ~n_5273) ;
	assign n_5271 = (~n_5269 & ~n_5270) ;
	assign n_5267 = (~n_5265 & ~n_5266) ;
	assign n_5264 = (~n_5262 & ~n_5263) ;
	assign n_5259 = (~n_5257 & ~n_5258) ;
	assign n_5256 = (~n_5254 & ~n_5255) ;
	assign n_5252 = (~n_5250 & ~n_5251) ;
	assign n_5249 = (~n_5247 & ~n_5248) ;
	assign n_5243 = (~n_5241 & ~n_5242) ;
	assign n_5240 = (~n_5238 & ~n_5239) ;
	assign n_5236 = (~n_5234 & ~n_5235) ;
	assign n_5233 = (~n_5231 & ~n_5232) ;
	assign n_5228 = (x_533 & n_452) ;
	assign n_5227 = (x_119 & n_347) ;
	assign n_5225 = (x_449 & n_467) ;
	assign n_5224 = (x_208 & n_362) ;
	assign n_5219 = (~n_5217 & ~n_5218) ;
	assign n_5216 = (~n_5214 & ~n_5215) ;
	assign n_5212 = (~n_5210 & ~n_5211) ;
	assign n_5209 = (~n_5207 & ~n_5208) ;
	assign n_5204 = (~n_5202 & ~n_5203) ;
	assign n_5201 = (~n_5199 & ~n_5200) ;
	assign n_5197 = (~n_5195 & ~n_5196) ;
	assign n_5194 = (~n_5192 & ~n_5193) ;
	assign n_5188 = (~n_5186 & ~n_5187) ;
	assign n_5185 = (~n_5183 & ~n_5184) ;
	assign n_5181 = (~n_5179 & ~n_5180) ;
	assign n_5178 = (~n_5176 & ~n_5177) ;
	assign n_5173 = (~n_5171 & ~n_5172) ;
	assign n_5170 = (~n_5168 & ~n_5169) ;
	assign n_5166 = (~n_5164 & ~n_5165) ;
	assign n_5163 = (~n_5161 & ~n_5162) ;
	assign n_5155 = (~n_5151 & n_5154) ;
	assign n_5149 = (n_5145 & n_5148) ;
	assign n_5142 = (n_5138 & n_5141) ;
	assign n_5133 = (~x_156 & ~n_179) ;
	assign n_5132 = (x_747 & n_287) ;
	assign n_5130 = (~x_680 & ~n_392) ;
	assign n_5129 = (x_439 & n_497) ;
	assign n_5125 = (n_5121 & n_5124) ;
	assign n_5118 = (n_5114 & n_5117) ;
	assign n_5110 = (n_5106 & n_5109) ;
	assign n_5103 = (n_5099 & n_5102) ;
	assign n_5094 = (n_5090 & n_5093) ;
	assign n_5087 = (n_5083 & n_5086) ;
	assign n_5079 = (n_5075 & n_5078) ;
	assign n_5072 = (n_5068 & n_5071) ;
	assign n_5061 = (~n_5059 & ~n_5060) ;
	assign n_5058 = (~n_5056 & ~n_5057) ;
	assign n_5054 = (~n_5052 & ~n_5053) ;
	assign n_5051 = (~n_5049 & ~n_5050) ;
	assign n_5046 = (~n_5044 & ~n_5045) ;
	assign n_5043 = (~n_5041 & ~n_5042) ;
	assign n_5039 = (~n_5037 & ~n_5038) ;
	assign n_5036 = (~n_5034 & ~n_5035) ;
	assign n_5030 = (x_90 & ~x_513) ;
	assign n_5029 = (x_235 & ~x_792) ;
	assign n_5027 = (x_322 & ~x_712) ;
	assign n_7913 = (~n_5342 & n_7912) ;
	assign n_5335 = (~n_5333 & ~n_5334) ;
	assign n_5327 = (~x_253 & n_5325) ;
	assign n_5326 = (x_253 & ~n_5325) ;
	assign n_5319 = (~n_5317 & ~n_5318) ;
	assign n_1550 = (n_20 & ~n_1549) ;
	assign n_1537 = (x_255 & n_18) ;
	assign n_5308 = (i_4 & n_59) ;
	assign n_5275 = (n_5271 & n_5274) ;
	assign n_5268 = (n_5264 & n_5267) ;
	assign n_5260 = (n_5256 & n_5259) ;
	assign n_5253 = (n_5249 & n_5252) ;
	assign n_5244 = (n_5240 & n_5243) ;
	assign n_5237 = (n_5233 & n_5236) ;
	assign n_5229 = (~n_5227 & ~n_5228) ;
	assign n_5226 = (~n_5224 & ~n_5225) ;
	assign n_5220 = (n_5216 & n_5219) ;
	assign n_5213 = (n_5209 & n_5212) ;
	assign n_5205 = (n_5201 & n_5204) ;
	assign n_5198 = (n_5194 & n_5197) ;
	assign n_5189 = (n_5185 & n_5188) ;
	assign n_5182 = (n_5178 & n_5181) ;
	assign n_5174 = (n_5170 & n_5173) ;
	assign n_5167 = (n_5163 & n_5166) ;
	assign n_5156 = (n_31 & n_5155) ;
	assign n_5150 = (n_5142 & n_5149) ;
	assign n_5134 = (~n_5132 & ~n_5133) ;
	assign n_5131 = (~n_5129 & ~n_5130) ;
	assign n_5126 = (n_5118 & n_5125) ;
	assign n_5111 = (n_5103 & n_5110) ;
	assign n_5095 = (n_5087 & n_5094) ;
	assign n_5080 = (n_5072 & n_5079) ;
	assign n_5062 = (n_5058 & n_5061) ;
	assign n_5055 = (n_5051 & n_5054) ;
	assign n_5047 = (n_5043 & n_5046) ;
	assign n_5040 = (n_5036 & n_5039) ;
	assign n_5031 = (~n_5029 & ~n_5030) ;
	assign n_5028 = (i_5 & ~n_5027) ;
	assign n_5025 = (x_226 & x_569) ;
	assign n_5024 = (~x_226 & ~x_569) ;
	assign n_7914 = (~n_5335 & n_7913) ;
	assign n_5328 = (~n_5326 & ~n_5327) ;
	assign n_5321 = (~x_254 & n_5319) ;
	assign n_5320 = (x_254 & ~n_5319) ;
	assign n_1551 = (~n_1537 & ~n_1550) ;
	assign n_5309 = (n_66 & n_5308) ;
	assign n_5307 = (x_256 & n_60) ;
	assign n_5276 = (n_5268 & n_5275) ;
	assign n_5261 = (n_5253 & n_5260) ;
	assign n_5245 = (n_5237 & n_5244) ;
	assign n_5230 = (n_5226 & n_5229) ;
	assign n_5221 = (n_5213 & n_5220) ;
	assign n_5206 = (n_5198 & n_5205) ;
	assign n_5190 = (n_5182 & n_5189) ;
	assign n_5175 = (n_5167 & n_5174) ;
	assign n_5157 = (n_5150 & n_5156) ;
	assign n_5135 = (n_5131 & n_5134) ;
	assign n_5127 = (n_5111 & n_5126) ;
	assign n_5096 = (n_5080 & n_5095) ;
	assign n_5063 = (n_5055 & n_5062) ;
	assign n_5048 = (n_5040 & n_5047) ;
	assign n_5032 = (n_5028 & n_5031) ;
	assign n_5026 = (~n_5024 & ~n_5025) ;
	assign n_7915 = (~n_5328 & n_7914) ;
	assign n_5322 = (~n_5320 & ~n_5321) ;
	assign n_5315 = (~x_255 & n_1551) ;
	assign n_5314 = (x_255 & ~n_1551) ;
	assign n_5310 = (~n_5307 & ~n_5309) ;
	assign n_5302 = (n_35 & ~n_452) ;
	assign n_5301 = (x_257 & n_36) ;
	assign n_5295 = (~x_258 & ~n_936) ;
	assign n_5277 = (n_5261 & n_5276) ;
	assign n_5246 = (n_5230 & n_5245) ;
	assign n_5222 = (n_5206 & n_5221) ;
	assign n_5191 = (n_5175 & n_5190) ;
	assign n_5158 = (n_5135 & n_5157) ;
	assign n_5128 = (n_5096 & n_5127) ;
	assign n_5064 = (n_5048 & n_5063) ;
	assign n_5033 = (~n_5026 & n_5032) ;
	assign n_7916 = (~n_5322 & n_7915) ;
	assign n_5316 = (~n_5314 & ~n_5315) ;
	assign n_5312 = (~x_256 & n_5310) ;
	assign n_5311 = (x_256 & ~n_5310) ;
	assign n_5303 = (~n_5301 & ~n_5302) ;
	assign n_5296 = (i_5 & ~n_5295) ;
	assign n_5294 = (~i_51 & n_936) ;
	assign n_5288 = (~x_259 & ~n_936) ;
	assign n_5278 = (n_5246 & n_5277) ;
	assign n_5223 = (n_5191 & n_5222) ;
	assign n_5159 = (n_5128 & n_5158) ;
	assign n_5065 = (n_5033 & n_5064) ;
	assign n_7917 = (~n_5316 & n_7916) ;
	assign n_5313 = (~n_5311 & ~n_5312) ;
	assign n_5305 = (~x_257 & n_5303) ;
	assign n_5304 = (x_257 & ~n_5303) ;
	assign n_5297 = (~n_5294 & n_5296) ;
	assign n_5289 = (i_5 & ~n_5288) ;
	assign n_5287 = (~i_60 & n_936) ;
	assign n_5281 = (i_5 & x_260) ;
	assign n_5279 = (n_5223 & n_5278) ;
	assign n_5160 = (n_5065 & n_5159) ;
	assign n_7918 = (~n_5313 & n_7917) ;
	assign n_5306 = (~n_5304 & ~n_5305) ;
	assign n_5299 = (~x_258 & ~n_5297) ;
	assign n_5298 = (x_258 & n_5297) ;
	assign n_5290 = (~n_5287 & n_5289) ;
	assign n_5282 = (~n_31 & n_5281) ;
	assign n_5280 = (n_5160 & n_5279) ;
	assign n_5018 = (i_61 & n_64) ;
	assign n_5010 = (~i_24 & n_669) ;
	assign n_5008 = (~x_110 & ~n_544) ;
	assign n_7919 = (~n_5306 & n_7918) ;
	assign n_5300 = (~n_5298 & ~n_5299) ;
	assign n_5292 = (~x_259 & ~n_5290) ;
	assign n_5291 = (x_259 & n_5290) ;
	assign n_5283 = (~n_5280 & ~n_5282) ;
	assign n_5019 = (n_66 & n_5018) ;
	assign n_5017 = (x_261 & n_978) ;
	assign n_5011 = (i_5 & ~n_5010) ;
	assign n_5009 = (n_662 & n_5008) ;
	assign n_7920 = (~n_5300 & n_7919) ;
	assign n_5293 = (~n_5291 & ~n_5292) ;
	assign n_5285 = (~x_260 & n_5283) ;
	assign n_5284 = (x_260 & ~n_5283) ;
	assign n_5020 = (~n_5017 & ~n_5019) ;
	assign n_5012 = (~n_5009 & n_5011) ;
	assign n_5007 = (~x_262 & ~n_665) ;
	assign n_5001 = (i_64 & n_64) ;
	assign n_7921 = (~n_5293 & n_7920) ;
	assign n_5286 = (~n_5284 & ~n_5285) ;
	assign n_5022 = (~x_261 & n_5020) ;
	assign n_5021 = (x_261 & ~n_5020) ;
	assign n_5013 = (~n_5007 & n_5012) ;
	assign n_5002 = (n_66 & n_5001) ;
	assign n_5000 = (x_263 & n_978) ;
	assign n_7922 = (~n_5286 & n_7921) ;
	assign n_5023 = (~n_5021 & ~n_5022) ;
	assign n_5015 = (~x_262 & ~n_5013) ;
	assign n_5014 = (x_262 & n_5013) ;
	assign n_5003 = (~n_5000 & ~n_5002) ;
	assign n_4995 = (~n_136 & n_1009) ;
	assign n_4994 = (x_264 & n_1007) ;
	assign n_4988 = (~x_265 & ~n_630) ;
	assign n_7923 = (~n_5023 & n_7922) ;
	assign n_5016 = (~n_5014 & ~n_5015) ;
	assign n_5005 = (~x_263 & n_5003) ;
	assign n_5004 = (x_263 & ~n_5003) ;
	assign n_4996 = (~n_4994 & ~n_4995) ;
	assign n_4989 = (i_5 & ~n_4988) ;
	assign n_4987 = (~i_15 & n_630) ;
	assign n_7924 = (~n_5016 & n_7923) ;
	assign n_5006 = (~n_5004 & ~n_5005) ;
	assign n_4998 = (~x_264 & n_4996) ;
	assign n_4997 = (x_264 & ~n_4996) ;
	assign n_4990 = (~n_4987 & n_4989) ;
	assign n_4982 = (x_337 & n_53) ;
	assign n_4981 = (x_266 & n_51) ;
	assign n_4975 = (~x_267 & ~n_544) ;
	assign n_7925 = (~n_5006 & n_7924) ;
	assign n_4999 = (~n_4997 & ~n_4998) ;
	assign n_4992 = (~x_265 & ~n_4990) ;
	assign n_4991 = (x_265 & n_4990) ;
	assign n_4983 = (~n_4981 & ~n_4982) ;
	assign n_4976 = (i_5 & ~n_4975) ;
	assign n_4974 = (~i_8 & n_544) ;
	assign n_4968 = (~x_268 & ~n_936) ;
	assign n_7926 = (~n_4999 & n_7925) ;
	assign n_4993 = (~n_4991 & ~n_4992) ;
	assign n_4985 = (~x_266 & n_4983) ;
	assign n_4984 = (x_266 & ~n_4983) ;
	assign n_4977 = (~n_4974 & n_4976) ;
	assign n_4969 = (i_5 & ~n_4968) ;
	assign n_4967 = (~i_58 & n_936) ;
	assign n_4961 = (i_24 & n_64) ;
	assign n_7927 = (~n_4993 & n_7926) ;
	assign n_4986 = (~n_4984 & ~n_4985) ;
	assign n_4979 = (~x_267 & ~n_4977) ;
	assign n_4978 = (x_267 & n_4977) ;
	assign n_4970 = (~n_4967 & n_4969) ;
	assign n_4962 = (n_66 & n_4961) ;
	assign n_4960 = (x_269 & n_978) ;
	assign n_4954 = (~x_270 & ~n_697) ;
	assign n_7928 = (~n_4986 & n_7927) ;
	assign n_4980 = (~n_4978 & ~n_4979) ;
	assign n_4972 = (~x_268 & ~n_4970) ;
	assign n_4971 = (x_268 & n_4970) ;
	assign n_4963 = (~n_4960 & ~n_4962) ;
	assign n_4955 = (i_5 & ~n_4954) ;
	assign n_4953 = (~x_504 & n_697) ;
	assign n_7929 = (~n_4980 & n_7928) ;
	assign n_4973 = (~n_4971 & ~n_4972) ;
	assign n_4965 = (~x_269 & n_4963) ;
	assign n_4964 = (x_269 & ~n_4963) ;
	assign n_4956 = (~n_4953 & n_4955) ;
	assign n_4948 = (x_389 & n_35) ;
	assign n_4947 = (x_271 & n_36) ;
	assign n_7930 = (~n_4973 & n_7929) ;
	assign n_4966 = (~n_4964 & ~n_4965) ;
	assign n_4958 = (~x_270 & ~n_4956) ;
	assign n_4957 = (x_270 & n_4956) ;
	assign n_4949 = (~n_4947 & ~n_4948) ;
	assign n_4942 = (~n_227 & n_1009) ;
	assign n_4941 = (x_272 & n_1007) ;
	assign n_4900 = (x_532 & ~x_726) ;
	assign n_4899 = (~x_532 & x_726) ;
	assign n_7931 = (~n_4966 & n_7930) ;
	assign n_4959 = (~n_4957 & ~n_4958) ;
	assign n_4951 = (~x_271 & n_4949) ;
	assign n_4950 = (x_271 & ~n_4949) ;
	assign n_4943 = (~n_4941 & ~n_4942) ;
	assign n_4936 = (i_42 & n_948) ;
	assign n_4935 = (x_273 & n_945) ;
	assign n_4929 = (~x_274 & ~n_544) ;
	assign n_4901 = (~n_4899 & ~n_4900) ;
	assign n_2847 = (x_634 & ~x_718) ;
	assign n_2843 = (x_358 & ~x_718) ;
	assign n_7932 = (~n_4959 & n_7931) ;
	assign n_4952 = (~n_4950 & ~n_4951) ;
	assign n_4945 = (~x_272 & n_4943) ;
	assign n_4944 = (x_272 & ~n_4943) ;
	assign n_4937 = (~n_4935 & ~n_4936) ;
	assign n_4930 = (i_5 & ~n_4929) ;
	assign n_4928 = (~i_54 & n_544) ;
	assign n_4922 = (~x_275 & ~n_697) ;
	assign n_4902 = (n_527 & ~n_4901) ;
	assign n_2848 = (~x_101 & ~n_2847) ;
	assign n_2846 = (x_333 & x_718) ;
	assign n_2844 = (x_101 & ~n_2843) ;
	assign n_2842 = (x_597 & x_718) ;
	assign n_2838 = (~n_2828 & ~n_2837) ;
	assign n_7933 = (~n_4952 & n_7932) ;
	assign n_4946 = (~n_4944 & ~n_4945) ;
	assign n_4939 = (~x_273 & n_4937) ;
	assign n_4938 = (x_273 & ~n_4937) ;
	assign n_4931 = (~n_4928 & n_4930) ;
	assign n_4923 = (i_5 & ~n_4922) ;
	assign n_4921 = (~x_775 & n_697) ;
	assign n_4915 = (i_19 & n_64) ;
	assign n_4907 = (n_139 & n_4902) ;
	assign n_4906 = (n_1 & n_4905) ;
	assign n_4903 = (~n_139 & ~n_4902) ;
	assign n_4855 = (~n_328 & ~n_329) ;
	assign n_2849 = (~n_2846 & n_2848) ;
	assign n_2845 = (~n_2842 & n_2844) ;
	assign n_2839 = (~n_2827 & ~n_2838) ;
	assign n_7934 = (~n_4946 & n_7933) ;
	assign n_4940 = (~n_4938 & ~n_4939) ;
	assign n_4933 = (~x_274 & ~n_4931) ;
	assign n_4932 = (x_274 & n_4931) ;
	assign n_4924 = (~n_4921 & n_4923) ;
	assign n_4916 = (n_66 & n_4915) ;
	assign n_4914 = (x_276 & n_978) ;
	assign n_4908 = (~n_4906 & ~n_4907) ;
	assign n_4904 = (~n_7 & n_4903) ;
	assign n_4857 = (~x_735 & ~n_4855) ;
	assign n_2860 = (x_182 & ~x_718) ;
	assign n_2856 = (x_448 & ~x_718) ;
	assign n_2850 = (~n_2845 & ~n_2849) ;
	assign n_2841 = (x_458 & n_2839) ;
	assign n_7935 = (~n_4940 & n_7934) ;
	assign n_4934 = (~n_4932 & ~n_4933) ;
	assign n_4926 = (~x_275 & ~n_4924) ;
	assign n_4925 = (x_275 & n_4924) ;
	assign n_4917 = (~n_4914 & ~n_4916) ;
	assign n_4909 = (~n_4904 & n_4908) ;
	assign n_4893 = (~x_278 & ~n_936) ;
	assign n_4858 = (~x_332 & ~n_4857) ;
	assign n_4856 = (x_735 & n_4855) ;
	assign n_2861 = (~x_101 & ~n_2860) ;
	assign n_2859 = (x_497 & x_718) ;
	assign n_2857 = (x_101 & ~n_2856) ;
	assign n_2855 = (x_233 & x_718) ;
	assign n_2851 = (~n_2841 & ~n_2850) ;
	assign n_2840 = (~x_458 & ~n_2839) ;
	assign n_7936 = (~n_4934 & n_7935) ;
	assign n_4927 = (~n_4925 & ~n_4926) ;
	assign n_4919 = (~x_276 & n_4917) ;
	assign n_4918 = (x_276 & ~n_4917) ;
	assign n_4910 = (i_5 & ~n_4909) ;
	assign n_4894 = (i_5 & ~n_4893) ;
	assign n_4892 = (~i_21 & n_936) ;
	assign n_4886 = (~x_279 & ~n_630) ;
	assign n_4859 = (~n_4856 & n_4858) ;
	assign n_2862 = (~n_2859 & n_2861) ;
	assign n_2858 = (~n_2855 & n_2857) ;
	assign n_2852 = (~n_2840 & ~n_2851) ;
	assign n_7937 = (~n_4927 & n_7936) ;
	assign n_4920 = (~n_4918 & ~n_4919) ;
	assign n_4912 = (~x_277 & ~n_4910) ;
	assign n_4911 = (x_277 & n_4910) ;
	assign n_4895 = (~n_4892 & n_4894) ;
	assign n_4887 = (i_5 & ~n_4886) ;
	assign n_4885 = (~i_23 & n_630) ;
	assign n_4861 = (n_332 & ~n_4859) ;
	assign n_2873 = (x_265 & ~x_718) ;
	assign n_2869 = (x_530 & ~x_718) ;
	assign n_2863 = (~n_2858 & ~n_2862) ;
	assign n_2854 = (x_376 & n_2852) ;
	assign n_7938 = (~n_4920 & n_7937) ;
	assign n_4913 = (~n_4911 & ~n_4912) ;
	assign n_4897 = (~x_278 & ~n_4895) ;
	assign n_4896 = (x_278 & n_4895) ;
	assign n_4888 = (~n_4885 & n_4887) ;
	assign n_4880 = (x_493 & n_53) ;
	assign n_4879 = (x_280 & n_51) ;
	assign n_4873 = (~x_281 & ~n_630) ;
	assign n_4865 = (~n_332 & ~n_1606) ;
	assign n_4864 = (i_10 & n_7) ;
	assign n_4862 = (x_664 & ~n_4861) ;
	assign n_4860 = (~n_332 & n_4859) ;
	assign n_2874 = (~x_101 & ~n_2873) ;
	assign n_2872 = (x_425 & x_718) ;
	assign n_2870 = (x_101 & ~n_2869) ;
	assign n_2868 = (x_149 & x_718) ;
	assign n_2864 = (~n_2854 & ~n_2863) ;
	assign n_2853 = (~x_376 & ~n_2852) ;
	assign n_7939 = (~n_4913 & n_7938) ;
	assign n_4898 = (~n_4896 & ~n_4897) ;
	assign n_4890 = (~x_279 & ~n_4888) ;
	assign n_4889 = (x_279 & n_4888) ;
	assign n_4881 = (~n_4879 & ~n_4880) ;
	assign n_4874 = (i_5 & ~n_4873) ;
	assign n_4872 = (~i_61 & n_630) ;
	assign n_4866 = (~n_4864 & ~n_4865) ;
	assign n_4863 = (~n_4860 & n_4862) ;
	assign n_2875 = (~n_2872 & n_2874) ;
	assign n_2871 = (~n_2868 & n_2870) ;
	assign n_2865 = (~n_2853 & ~n_2864) ;
	assign n_7940 = (~n_4898 & n_7939) ;
	assign n_4891 = (~n_4889 & ~n_4890) ;
	assign n_4883 = (~x_280 & n_4881) ;
	assign n_4882 = (x_280 & ~n_4881) ;
	assign n_4875 = (~n_4872 & n_4874) ;
	assign n_4867 = (~n_4863 & n_4866) ;
	assign n_2887 = (x_570 & ~x_718) ;
	assign n_2883 = (x_306 & ~x_718) ;
	assign n_2876 = (~n_2871 & ~n_2875) ;
	assign n_2867 = (x_432 & n_2865) ;
	assign n_7941 = (~n_4891 & n_7940) ;
	assign n_4884 = (~n_4882 & ~n_4883) ;
	assign n_4877 = (~x_281 & ~n_4875) ;
	assign n_4876 = (x_281 & n_4875) ;
	assign n_4868 = (i_5 & ~n_4867) ;
	assign n_4850 = (i_13 & n_948) ;
	assign n_4849 = (x_283 & n_945) ;
	assign n_4820 = (i_68 & ~n_6) ;
	assign n_2888 = (~x_101 & ~n_2887) ;
	assign n_2886 = (x_384 & x_718) ;
	assign n_2884 = (x_101 & ~n_2883) ;
	assign n_2882 = (x_668 & x_718) ;
	assign n_2877 = (~n_2867 & ~n_2876) ;
	assign n_2866 = (~x_432 & ~n_2865) ;
	assign n_7942 = (~n_4884 & n_7941) ;
	assign n_4878 = (~n_4876 & ~n_4877) ;
	assign n_4870 = (~x_282 & ~n_4868) ;
	assign n_4869 = (x_282 & n_4868) ;
	assign n_4851 = (~n_4849 & ~n_4850) ;
	assign n_4844 = (x_738 & n_53) ;
	assign n_4843 = (x_284 & n_51) ;
	assign n_4837 = (i_42 & n_59) ;
	assign n_4821 = (n_629 & ~n_4820) ;
	assign n_4819 = (x_287 & n_6) ;
	assign n_2889 = (~n_2886 & n_2888) ;
	assign n_2885 = (~n_2882 & n_2884) ;
	assign n_2878 = (~n_2866 & ~n_2877) ;
	assign n_7943 = (~n_4878 & n_7942) ;
	assign n_4871 = (~n_4869 & ~n_4870) ;
	assign n_4853 = (~x_283 & n_4851) ;
	assign n_4852 = (x_283 & ~n_4851) ;
	assign n_4845 = (~n_4843 & ~n_4844) ;
	assign n_4838 = (n_66 & n_4837) ;
	assign n_4836 = (x_285 & n_60) ;
	assign n_4830 = (~x_286 & ~n_936) ;
	assign n_4822 = (~n_4819 & n_4821) ;
	assign n_4020 = (x_483 & ~x_718) ;
	assign n_4016 = (x_224 & ~x_718) ;
	assign n_2890 = (~n_2885 & ~n_2889) ;
	assign n_2880 = (x_504 & n_2878) ;
	assign n_7944 = (~n_4871 & n_7943) ;
	assign n_4854 = (~n_4852 & ~n_4853) ;
	assign n_4847 = (~x_284 & n_4845) ;
	assign n_4846 = (x_284 & ~n_4845) ;
	assign n_4839 = (~n_4836 & ~n_4838) ;
	assign n_4831 = (i_5 & ~n_4830) ;
	assign n_4829 = (~i_48 & n_936) ;
	assign n_4823 = (i_5 & ~n_4822) ;
	assign n_4818 = (~x_225 & n_662) ;
	assign n_4021 = (~x_101 & ~n_4020) ;
	assign n_4019 = (x_466 & x_718) ;
	assign n_4017 = (x_101 & ~n_4016) ;
	assign n_4015 = (x_718 & x_751) ;
	assign n_4011 = (~n_2880 & ~n_2890) ;
	assign n_2879 = (~x_504 & ~n_2878) ;
	assign n_7945 = (~n_4854 & n_7944) ;
	assign n_4848 = (~n_4846 & ~n_4847) ;
	assign n_4841 = (~x_285 & n_4839) ;
	assign n_4840 = (x_285 & ~n_4839) ;
	assign n_4832 = (~n_4829 & n_4831) ;
	assign n_4824 = (~n_4818 & n_4823) ;
	assign n_4817 = (~x_287 & n_663) ;
	assign n_4022 = (~n_4019 & n_4021) ;
	assign n_4018 = (~n_4015 & n_4017) ;
	assign n_4012 = (~n_2879 & ~n_4011) ;
	assign n_7946 = (~n_4848 & n_7945) ;
	assign n_4842 = (~n_4840 & ~n_4841) ;
	assign n_4834 = (~x_286 & ~n_4832) ;
	assign n_4833 = (x_286 & n_4832) ;
	assign n_4825 = (~n_4817 & n_4824) ;
	assign n_4812 = (x_299 & n_53) ;
	assign n_4811 = (x_288 & n_51) ;
	assign n_4805 = (~x_289 & ~n_697) ;
	assign n_4034 = (x_541 & ~x_718) ;
	assign n_4030 = (x_274 & ~x_718) ;
	assign n_4023 = (~n_4018 & ~n_4022) ;
	assign n_4014 = (x_323 & n_4012) ;
	assign n_7947 = (~n_4842 & n_7946) ;
	assign n_4835 = (~n_4833 & ~n_4834) ;
	assign n_4827 = (~x_287 & ~n_4825) ;
	assign n_4826 = (x_287 & n_4825) ;
	assign n_4813 = (~n_4811 & ~n_4812) ;
	assign n_4806 = (i_5 & ~n_4805) ;
	assign n_4804 = (~x_529 & n_697) ;
	assign n_4798 = (i_29 & n_59) ;
	assign n_4035 = (~x_101 & ~n_4034) ;
	assign n_4033 = (x_414 & x_718) ;
	assign n_4031 = (x_101 & ~n_4030) ;
	assign n_4029 = (x_700 & x_718) ;
	assign n_4024 = (~n_4014 & ~n_4023) ;
	assign n_4013 = (~x_323 & ~n_4012) ;
	assign n_7948 = (~n_4835 & n_7947) ;
	assign n_4828 = (~n_4826 & ~n_4827) ;
	assign n_4815 = (~x_288 & n_4813) ;
	assign n_4814 = (x_288 & ~n_4813) ;
	assign n_4807 = (~n_4804 & n_4806) ;
	assign n_4799 = (n_66 & n_4798) ;
	assign n_4797 = (x_290 & n_60) ;
	assign n_4791 = (~x_291 & ~n_630) ;
	assign n_4036 = (~n_4033 & n_4035) ;
	assign n_4032 = (~n_4029 & n_4031) ;
	assign n_4025 = (~n_4013 & ~n_4024) ;
	assign n_7949 = (~n_4828 & n_7948) ;
	assign n_4816 = (~n_4814 & ~n_4815) ;
	assign n_4809 = (~x_289 & ~n_4807) ;
	assign n_4808 = (x_289 & n_4807) ;
	assign n_4800 = (~n_4797 & ~n_4799) ;
	assign n_4792 = (i_5 & ~n_4791) ;
	assign n_4790 = (~i_57 & n_630) ;
	assign n_4784 = (i_23 & n_64) ;
	assign n_4037 = (~n_4032 & ~n_4036) ;
	assign n_4027 = (x_370 & n_4025) ;
	assign n_7950 = (~n_4816 & n_7949) ;
	assign n_4810 = (~n_4808 & ~n_4809) ;
	assign n_4802 = (~x_290 & n_4800) ;
	assign n_4801 = (x_290 & ~n_4800) ;
	assign n_4793 = (~n_4790 & n_4792) ;
	assign n_4785 = (n_66 & n_4784) ;
	assign n_4783 = (x_292 & n_978) ;
	assign n_4763 = (i_38 & n_1) ;
	assign n_4684 = (~n_4027 & ~n_4037) ;
	assign n_4026 = (~x_370 & ~n_4025) ;
	assign n_4680 = (x_279 & ~x_718) ;
	assign n_4676 = (x_543 & ~x_718) ;
	assign n_7951 = (~n_4810 & n_7950) ;
	assign n_4803 = (~n_4801 & ~n_4802) ;
	assign n_4795 = (~x_291 & ~n_4793) ;
	assign n_4794 = (x_291 & n_4793) ;
	assign n_4786 = (~n_4783 & ~n_4785) ;
	assign n_4767 = (x_408 & ~n_16) ;
	assign n_4766 = (i_38 & n_7) ;
	assign n_4764 = (~n_17 & ~n_4763) ;
	assign n_4723 = (~x_349 & n_2824) ;
	assign n_4722 = (x_349 & ~n_2824) ;
	assign n_4685 = (~n_4026 & ~n_4684) ;
	assign n_4681 = (~x_101 & ~n_4680) ;
	assign n_4679 = (x_411 & x_718) ;
	assign n_4677 = (x_101 & ~n_4676) ;
	assign n_4675 = (x_133 & x_718) ;
	assign n_7952 = (~n_4803 & n_7951) ;
	assign n_4796 = (~n_4794 & ~n_4795) ;
	assign n_4788 = (~x_292 & n_4786) ;
	assign n_4787 = (x_292 & ~n_4786) ;
	assign n_4775 = (i_49 & n_948) ;
	assign n_4774 = (x_294 & n_945) ;
	assign n_4768 = (~n_4766 & ~n_4767) ;
	assign n_4765 = (x_295 & ~n_4764) ;
	assign n_4724 = (~n_4722 & ~n_4723) ;
	assign n_4721 = (~n_2814 & ~n_2815) ;
	assign n_4687 = (~x_728 & n_4685) ;
	assign n_4686 = (x_728 & ~n_4685) ;
	assign n_4682 = (~n_4679 & n_4681) ;
	assign n_4678 = (~n_4675 & n_4677) ;
	assign n_7953 = (~n_4796 & n_7952) ;
	assign n_4789 = (~n_4787 & ~n_4788) ;
	assign n_4781 = (~x_293 & n_392) ;
	assign n_4780 = (x_293 & ~n_392) ;
	assign n_4776 = (~n_4774 & ~n_4775) ;
	assign n_4769 = (~n_4765 & n_4768) ;
	assign n_4757 = (i_28 & n_59) ;
	assign n_4733 = (~x_299 & n_6) ;
	assign n_4726 = (n_4721 & ~n_4724) ;
	assign n_4688 = (~n_4686 & ~n_4687) ;
	assign n_4683 = (~n_4678 & ~n_4682) ;
	assign n_7954 = (~n_4789 & n_7953) ;
	assign n_4782 = (~n_4780 & ~n_4781) ;
	assign n_4778 = (~x_294 & n_4776) ;
	assign n_4777 = (x_294 & ~n_4776) ;
	assign n_4770 = (i_5 & ~n_4769) ;
	assign n_4758 = (n_66 & n_4757) ;
	assign n_4756 = (x_296 & n_60) ;
	assign n_4750 = (i_50 & n_59) ;
	assign n_4734 = (~n_4732 & ~n_4733) ;
	assign n_4729 = (x_299 & ~n_697) ;
	assign n_4727 = (n_697 & ~n_4726) ;
	assign n_4725 = (~n_4721 & n_4724) ;
	assign n_4690 = (~n_4683 & n_4688) ;
	assign n_7955 = (~n_4782 & n_7954) ;
	assign n_4779 = (~n_4777 & ~n_4778) ;
	assign n_4772 = (~x_295 & ~n_4770) ;
	assign n_4771 = (x_295 & n_4770) ;
	assign n_4759 = (~n_4756 & ~n_4758) ;
	assign n_4751 = (n_66 & n_4750) ;
	assign n_4749 = (x_297 & n_60) ;
	assign n_4743 = (~x_298 & ~n_630) ;
	assign n_4735 = (n_629 & ~n_4734) ;
	assign n_4730 = (~n_629 & ~n_4729) ;
	assign n_4728 = (~n_4725 & n_4727) ;
	assign n_4691 = (n_697 & ~n_4690) ;
	assign n_4689 = (n_4683 & ~n_4688) ;
	assign n_7956 = (~n_4779 & n_7955) ;
	assign n_4773 = (~n_4771 & ~n_4772) ;
	assign n_4761 = (~x_296 & n_4759) ;
	assign n_4760 = (x_296 & ~n_4759) ;
	assign n_4752 = (~n_4749 & ~n_4751) ;
	assign n_4744 = (i_5 & ~n_4743) ;
	assign n_4742 = (~i_49 & n_630) ;
	assign n_4736 = (n_902 & ~n_4735) ;
	assign n_4731 = (~n_4728 & n_4730) ;
	assign n_4697 = (~x_302 & n_6) ;
	assign n_1237 = (~i_23 & ~n_6) ;
	assign n_4692 = (~n_4689 & n_4691) ;
	assign n_7957 = (~n_4773 & n_7956) ;
	assign n_4762 = (~n_4760 & ~n_4761) ;
	assign n_4754 = (~x_297 & n_4752) ;
	assign n_4753 = (x_297 & ~n_4752) ;
	assign n_4745 = (~n_4742 & n_4744) ;
	assign n_4737 = (~n_4731 & n_4736) ;
	assign n_4720 = (x_299 & n_699) ;
	assign n_4714 = (~x_300 & ~n_544) ;
	assign n_4698 = (~n_1237 & ~n_4697) ;
	assign n_4694 = (~x_302 & n_4692) ;
	assign n_7958 = (~n_4762 & n_7957) ;
	assign n_4755 = (~n_4753 & ~n_4754) ;
	assign n_4747 = (~x_298 & ~n_4745) ;
	assign n_4746 = (x_298 & n_4745) ;
	assign n_4738 = (~n_4720 & ~n_4737) ;
	assign n_4715 = (i_5 & ~n_4714) ;
	assign n_4713 = (~i_37 & n_544) ;
	assign n_4707 = (~x_301 & ~n_544) ;
	assign n_4699 = (n_629 & ~n_4698) ;
	assign n_4695 = (~n_629 & ~n_4694) ;
	assign n_4693 = (x_302 & ~n_4692) ;
	assign n_7959 = (~n_4755 & n_7958) ;
	assign n_4748 = (~n_4746 & ~n_4747) ;
	assign n_4740 = (~x_299 & n_4738) ;
	assign n_4739 = (x_299 & ~n_4738) ;
	assign n_4716 = (~n_4713 & n_4715) ;
	assign n_4708 = (i_5 & ~n_4707) ;
	assign n_4706 = (~i_21 & n_544) ;
	assign n_4700 = (n_902 & ~n_4699) ;
	assign n_4696 = (~n_4693 & n_4695) ;
	assign n_4630 = (~x_137 & n_812) ;
	assign n_4629 = (x_137 & ~n_812) ;
	assign n_7960 = (~n_4748 & n_7959) ;
	assign n_4741 = (~n_4739 & ~n_4740) ;
	assign n_4718 = (~x_300 & ~n_4716) ;
	assign n_4717 = (x_300 & n_4716) ;
	assign n_4709 = (~n_4706 & n_4708) ;
	assign n_4701 = (~n_4696 & n_4700) ;
	assign n_4674 = (x_302 & n_699) ;
	assign n_4631 = (~n_4629 & ~n_4630) ;
	assign n_4628 = (~n_802 & ~n_803) ;
	assign n_7961 = (~n_4741 & n_7960) ;
	assign n_4719 = (~n_4717 & ~n_4718) ;
	assign n_4711 = (~x_301 & ~n_4709) ;
	assign n_4710 = (x_301 & n_4709) ;
	assign n_4702 = (~n_4674 & ~n_4701) ;
	assign n_4669 = (n_35 & ~n_482) ;
	assign n_4668 = (x_303 & n_36) ;
	assign n_4640 = (~x_307 & n_6) ;
	assign n_4633 = (n_4628 & ~n_4631) ;
	assign n_7962 = (~n_4719 & n_7961) ;
	assign n_4712 = (~n_4710 & ~n_4711) ;
	assign n_4704 = (~x_302 & n_4702) ;
	assign n_4703 = (x_302 & ~n_4702) ;
	assign n_4670 = (~n_4668 & ~n_4669) ;
	assign n_4663 = (i_24 & n_948) ;
	assign n_4662 = (x_304 & n_945) ;
	assign n_4641 = (~n_4639 & ~n_4640) ;
	assign n_4636 = (x_307 & ~n_697) ;
	assign n_4634 = (n_697 & ~n_4633) ;
	assign n_4632 = (~n_4628 & n_4631) ;
	assign n_7963 = (~n_4712 & n_7962) ;
	assign n_4705 = (~n_4703 & ~n_4704) ;
	assign n_4672 = (~x_303 & n_4670) ;
	assign n_4671 = (x_303 & ~n_4670) ;
	assign n_4664 = (~n_4662 & ~n_4663) ;
	assign n_4657 = (x_567 & n_53) ;
	assign n_4656 = (x_305 & n_51) ;
	assign n_4650 = (~x_306 & ~n_544) ;
	assign n_4642 = (n_629 & ~n_4641) ;
	assign n_4637 = (~n_629 & ~n_4636) ;
	assign n_4635 = (~n_4632 & n_4634) ;
	assign n_7964 = (~n_4705 & n_7963) ;
	assign n_4673 = (~n_4671 & ~n_4672) ;
	assign n_4666 = (~x_304 & n_4664) ;
	assign n_4665 = (x_304 & ~n_4664) ;
	assign n_4658 = (~n_4656 & ~n_4657) ;
	assign n_4651 = (i_5 & ~n_4650) ;
	assign n_4649 = (~i_42 & n_544) ;
	assign n_4643 = (n_902 & ~n_4642) ;
	assign n_4638 = (~n_4635 & n_4637) ;
	assign n_7965 = (~n_4673 & n_7964) ;
	assign n_4667 = (~n_4665 & ~n_4666) ;
	assign n_4660 = (~x_305 & n_4658) ;
	assign n_4659 = (x_305 & ~n_4658) ;
	assign n_4652 = (~n_4649 & n_4651) ;
	assign n_4644 = (~n_4638 & n_4643) ;
	assign n_4627 = (x_307 & n_699) ;
	assign n_7966 = (~n_4667 & n_7965) ;
	assign n_4661 = (~n_4659 & ~n_4660) ;
	assign n_4654 = (~x_306 & ~n_4652) ;
	assign n_4653 = (x_306 & n_4652) ;
	assign n_4645 = (~n_4627 & ~n_4644) ;
	assign n_4618 = (i_8 & n_64) ;
	assign n_4578 = (~x_355 & ~x_357) ;
	assign n_4577 = (~x_322 & x_332) ;
	assign n_4575 = (~x_435 & ~x_439) ;
	assign n_4574 = (~x_365 & ~x_394) ;
	assign n_4571 = (~x_273 & ~x_283) ;
	assign n_4570 = (~x_241 & ~x_243) ;
	assign n_4568 = (~x_313 & ~x_321) ;
	assign n_4567 = (~x_294 & ~x_304) ;
	assign n_4563 = (~x_575 & ~x_584) ;
	assign n_4562 = (~x_533 & ~x_537) ;
	assign n_4560 = (~x_607 & ~x_614) ;
	assign n_4559 = (~x_594 & ~x_596) ;
	assign n_4556 = (~x_471 & ~x_487) ;
	assign n_4555 = (~x_449 & ~x_461) ;
	assign n_4553 = (~x_513 & ~x_521) ;
	assign n_4552 = (~x_505 & ~x_509) ;
	assign n_7967 = (~n_4661 & n_7966) ;
	assign n_4655 = (~n_4653 & ~n_4654) ;
	assign n_4647 = (~x_307 & n_4645) ;
	assign n_4646 = (x_307 & ~n_4645) ;
	assign n_4619 = (n_66 & n_4618) ;
	assign n_4617 = (x_309 & n_978) ;
	assign n_4611 = (~x_310 & ~n_630) ;
	assign n_4579 = (n_4577 & n_4578) ;
	assign n_4576 = (n_4574 & n_4575) ;
	assign n_4572 = (n_4570 & n_4571) ;
	assign n_4569 = (n_4567 & n_4568) ;
	assign n_4564 = (n_4562 & n_4563) ;
	assign n_4561 = (n_4559 & n_4560) ;
	assign n_4557 = (n_4555 & n_4556) ;
	assign n_4554 = (n_4552 & n_4553) ;
	assign n_4548 = (~x_747 & ~x_757) ;
	assign n_4547 = (~x_736 & ~x_743) ;
	assign n_4545 = (~x_797 & ~x_801) ;
	assign n_4544 = (~x_771 & ~x_772) ;
	assign n_4541 = (~x_661 & ~x_665) ;
	assign n_4540 = (~x_626 & ~x_660) ;
	assign n_4538 = (~x_692 & ~x_713) ;
	assign n_4537 = (~x_673 & ~x_680) ;
	assign n_4532 = (~x_187 & ~x_208) ;
	assign n_4531 = (~x_158 & ~x_170) ;
	assign n_4529 = (~x_226 & ~x_235) ;
	assign n_4528 = (~x_217 & ~x_221) ;
	assign n_4525 = (~x_88 & ~x_119) ;
	assign n_4524 = (~x_81 & ~x_85) ;
	assign n_4522 = (~x_153 & ~x_156) ;
	assign n_4521 = (~x_127 & ~x_139) ;
	assign n_7968 = (~n_4655 & n_7967) ;
	assign n_4648 = (~n_4646 & ~n_4647) ;
	assign n_4625 = (~x_308 & n_1223) ;
	assign n_4624 = (x_308 & ~n_1223) ;
	assign n_4620 = (~n_4617 & ~n_4619) ;
	assign n_4612 = (i_5 & ~n_4611) ;
	assign n_4610 = (~i_58 & n_630) ;
	assign n_4580 = (n_4576 & n_4579) ;
	assign n_4573 = (n_4569 & n_4572) ;
	assign n_4565 = (n_4561 & n_4564) ;
	assign n_4558 = (n_4554 & n_4557) ;
	assign n_4549 = (n_4547 & n_4548) ;
	assign n_4546 = (n_4544 & n_4545) ;
	assign n_4542 = (n_4540 & n_4541) ;
	assign n_4539 = (n_4537 & n_4538) ;
	assign n_4533 = (n_4531 & n_4532) ;
	assign n_4530 = (n_4528 & n_4529) ;
	assign n_4526 = (n_4524 & n_4525) ;
	assign n_4523 = (n_4521 & n_4522) ;
	assign n_4518 = (i_5 & ~x_74) ;
	assign n_7969 = (~n_4648 & n_7968) ;
	assign n_4626 = (~n_4624 & ~n_4625) ;
	assign n_4622 = (~x_309 & n_4620) ;
	assign n_4621 = (x_309 & ~n_4620) ;
	assign n_4613 = (~n_4610 & n_4612) ;
	assign n_4605 = (x_547 & n_35) ;
	assign n_4604 = (x_311 & n_36) ;
	assign n_4598 = (~x_312 & ~n_936) ;
	assign n_4581 = (n_4573 & n_4580) ;
	assign n_4566 = (n_4558 & n_4565) ;
	assign n_4550 = (n_4546 & n_4549) ;
	assign n_4543 = (n_4539 & n_4542) ;
	assign n_4534 = (n_4530 & n_4533) ;
	assign n_4527 = (n_4523 & n_4526) ;
	assign n_4519 = (n_8 & n_4518) ;
	assign n_7970 = (~n_4626 & n_7969) ;
	assign n_4623 = (~n_4621 & ~n_4622) ;
	assign n_4615 = (~x_310 & ~n_4613) ;
	assign n_4614 = (x_310 & n_4613) ;
	assign n_4606 = (~n_4604 & ~n_4605) ;
	assign n_4599 = (i_5 & ~n_4598) ;
	assign n_4597 = (~i_7 & n_936) ;
	assign n_4582 = (n_4566 & n_4581) ;
	assign n_4551 = (n_4543 & n_4550) ;
	assign n_4535 = (n_4527 & n_4534) ;
	assign n_4520 = (n_9 & n_4519) ;
	assign n_7971 = (~n_4623 & n_7970) ;
	assign n_4616 = (~n_4614 & ~n_4615) ;
	assign n_4608 = (~x_311 & n_4606) ;
	assign n_4607 = (x_311 & ~n_4606) ;
	assign n_4600 = (~n_4597 & n_4599) ;
	assign n_4592 = (i_33 & n_948) ;
	assign n_4591 = (x_313 & n_945) ;
	assign n_4585 = (x_314 & n_29) ;
	assign n_4583 = (n_4551 & n_4582) ;
	assign n_4536 = (n_4520 & n_4535) ;
	assign n_7972 = (~n_4616 & n_7971) ;
	assign n_4609 = (~n_4607 & ~n_4608) ;
	assign n_4602 = (~x_312 & ~n_4600) ;
	assign n_4601 = (x_312 & n_4600) ;
	assign n_4593 = (~n_4591 & ~n_4592) ;
	assign n_4586 = (~n_31 & n_4585) ;
	assign n_4584 = (n_4536 & n_4583) ;
	assign n_4505 = (i_19 & n_7) ;
	assign n_4504 = (x_547 & ~n_16) ;
	assign n_4465 = (~x_464 & n_734) ;
	assign n_4464 = (x_464 & ~n_734) ;
	assign n_7973 = (~n_4609 & n_7972) ;
	assign n_4603 = (~n_4601 & ~n_4602) ;
	assign n_4595 = (~x_313 & n_4593) ;
	assign n_4594 = (x_313 & ~n_4593) ;
	assign n_4587 = (~n_4584 & ~n_4586) ;
	assign n_4513 = (x_272 & n_35) ;
	assign n_4512 = (x_315 & n_36) ;
	assign n_4506 = (~n_4504 & ~n_4505) ;
	assign n_4466 = (~n_4464 & ~n_4465) ;
	assign n_4463 = (~n_724 & ~n_725) ;
	assign n_7974 = (~n_4603 & n_7973) ;
	assign n_4596 = (~n_4594 & ~n_4595) ;
	assign n_4589 = (~x_314 & n_4587) ;
	assign n_4588 = (x_314 & ~n_4587) ;
	assign n_4514 = (~n_4512 & ~n_4513) ;
	assign n_4507 = (n_20 & ~n_4506) ;
	assign n_4503 = (x_316 & n_18) ;
	assign n_4497 = (~x_317 & ~n_544) ;
	assign n_4475 = (i_55 & ~n_6) ;
	assign n_4468 = (n_4463 & ~n_4466) ;
	assign n_7975 = (~n_4596 & n_7974) ;
	assign n_4590 = (~n_4588 & ~n_4589) ;
	assign n_4516 = (~x_315 & n_4514) ;
	assign n_4515 = (x_315 & ~n_4514) ;
	assign n_4508 = (~n_4503 & ~n_4507) ;
	assign n_4498 = (i_5 & ~n_4497) ;
	assign n_4496 = (~i_17 & n_544) ;
	assign n_4476 = (n_629 & ~n_4475) ;
	assign n_4474 = (x_320 & n_6) ;
	assign n_4471 = (x_320 & ~n_697) ;
	assign n_4469 = (n_697 & ~n_4468) ;
	assign n_4467 = (~n_4463 & n_4466) ;
	assign n_4431 = (~x_703 & n_4023) ;
	assign n_4430 = (x_703 & ~n_4023) ;
	assign n_7976 = (~n_4590 & n_7975) ;
	assign n_4517 = (~n_4515 & ~n_4516) ;
	assign n_4510 = (~x_316 & n_4508) ;
	assign n_4509 = (x_316 & ~n_4508) ;
	assign n_4499 = (~n_4496 & n_4498) ;
	assign n_4491 = (x_70 & n_53) ;
	assign n_4490 = (x_318 & n_51) ;
	assign n_4477 = (~n_4474 & n_4476) ;
	assign n_4472 = (~n_629 & ~n_4471) ;
	assign n_4470 = (~n_4467 & n_4469) ;
	assign n_4432 = (~n_4430 & ~n_4431) ;
	assign n_4429 = (~n_4013 & ~n_4014) ;
	assign n_7977 = (~n_4517 & n_7976) ;
	assign n_4511 = (~n_4509 & ~n_4510) ;
	assign n_4501 = (~x_317 & ~n_4499) ;
	assign n_4500 = (x_317 & n_4499) ;
	assign n_4492 = (~n_4490 & ~n_4491) ;
	assign n_4485 = (~n_242 & n_35) ;
	assign n_4484 = (x_319 & n_36) ;
	assign n_4478 = (n_902 & ~n_4477) ;
	assign n_4473 = (~n_4470 & n_4472) ;
	assign n_4441 = (~x_323 & n_6) ;
	assign n_4434 = (n_4429 & ~n_4432) ;
	assign n_7978 = (~n_4511 & n_7977) ;
	assign n_4502 = (~n_4500 & ~n_4501) ;
	assign n_4494 = (~x_318 & n_4492) ;
	assign n_4493 = (x_318 & ~n_4492) ;
	assign n_4486 = (~n_4484 & ~n_4485) ;
	assign n_4479 = (~n_4473 & n_4478) ;
	assign n_4462 = (x_320 & n_699) ;
	assign n_4442 = (~n_4440 & ~n_4441) ;
	assign n_4437 = (x_323 & ~n_697) ;
	assign n_4435 = (n_697 & ~n_4434) ;
	assign n_4433 = (~n_4429 & n_4432) ;
	assign n_7979 = (~n_4502 & n_7978) ;
	assign n_4495 = (~n_4493 & ~n_4494) ;
	assign n_4488 = (~x_319 & n_4486) ;
	assign n_4487 = (x_319 & ~n_4486) ;
	assign n_4480 = (~n_4462 & ~n_4479) ;
	assign n_4457 = (i_52 & n_948) ;
	assign n_4456 = (x_321 & n_945) ;
	assign n_4443 = (n_629 & ~n_4442) ;
	assign n_4438 = (~n_629 & ~n_4437) ;
	assign n_4436 = (~n_4433 & n_4435) ;
	assign n_7980 = (~n_4495 & n_7979) ;
	assign n_4489 = (~n_4487 & ~n_4488) ;
	assign n_4482 = (~x_320 & n_4480) ;
	assign n_4481 = (x_320 & ~n_4480) ;
	assign n_4458 = (~n_4456 & ~n_4457) ;
	assign n_4451 = (i_39 & n_948) ;
	assign n_4450 = (x_322 & n_945) ;
	assign n_4444 = (n_902 & ~n_4443) ;
	assign n_4439 = (~n_4436 & n_4438) ;
	assign n_7981 = (~n_4489 & n_7980) ;
	assign n_4483 = (~n_4481 & ~n_4482) ;
	assign n_4460 = (~x_321 & n_4458) ;
	assign n_4459 = (x_321 & ~n_4458) ;
	assign n_4452 = (~n_4450 & ~n_4451) ;
	assign n_4445 = (~n_4439 & n_4444) ;
	assign n_4428 = (x_323 & n_699) ;
	assign n_4422 = (~x_324 & ~n_936) ;
	assign n_4407 = (~x_326 & n_6) ;
	assign n_4402 = (~x_190 & ~n_544) ;
	assign n_7982 = (~n_4483 & n_7981) ;
	assign n_4461 = (~n_4459 & ~n_4460) ;
	assign n_4454 = (~x_322 & n_4452) ;
	assign n_4453 = (x_322 & ~n_4452) ;
	assign n_4446 = (~n_4428 & ~n_4445) ;
	assign n_4423 = (i_5 & ~n_4422) ;
	assign n_4421 = (~i_46 & n_936) ;
	assign n_4408 = (~n_4406 & ~n_4407) ;
	assign n_4403 = (n_662 & ~n_4402) ;
	assign n_7983 = (~n_4461 & n_7982) ;
	assign n_4455 = (~n_4453 & ~n_4454) ;
	assign n_4448 = (~x_323 & n_4446) ;
	assign n_4447 = (x_323 & ~n_4446) ;
	assign n_4424 = (~n_4421 & n_4423) ;
	assign n_4416 = (x_779 & n_35) ;
	assign n_4415 = (x_325 & n_36) ;
	assign n_4409 = (n_629 & ~n_4408) ;
	assign n_4404 = (~n_629 & ~n_4403) ;
	assign n_4401 = (x_326 & ~n_662) ;
	assign n_7984 = (~n_4455 & n_7983) ;
	assign n_4449 = (~n_4447 & ~n_4448) ;
	assign n_4426 = (~x_324 & ~n_4424) ;
	assign n_4425 = (x_324 & n_4424) ;
	assign n_4417 = (~n_4415 & ~n_4416) ;
	assign n_4410 = (i_5 & ~n_4409) ;
	assign n_4405 = (~n_4401 & n_4404) ;
	assign n_7985 = (~n_4449 & n_7984) ;
	assign n_4427 = (~n_4425 & ~n_4426) ;
	assign n_4419 = (~x_325 & n_4417) ;
	assign n_4418 = (x_325 & ~n_4417) ;
	assign n_4411 = (~n_4405 & n_4410) ;
	assign n_4396 = (x_633 & n_53) ;
	assign n_4395 = (x_327 & n_51) ;
	assign n_7986 = (~n_4427 & n_7985) ;
	assign n_4420 = (~n_4418 & ~n_4419) ;
	assign n_4413 = (~x_326 & ~n_4411) ;
	assign n_4412 = (x_326 & n_4411) ;
	assign n_4397 = (~n_4395 & ~n_4396) ;
	assign n_4390 = (~n_107 & n_1009) ;
	assign n_4389 = (x_328 & n_1007) ;
	assign n_4383 = (~x_329 & ~n_630) ;
	assign n_7987 = (~n_4420 & n_7986) ;
	assign n_4414 = (~n_4412 & ~n_4413) ;
	assign n_4399 = (~x_327 & n_4397) ;
	assign n_4398 = (x_327 & ~n_4397) ;
	assign n_4391 = (~n_4389 & ~n_4390) ;
	assign n_4384 = (i_5 & ~n_4383) ;
	assign n_4382 = (~i_27 & n_630) ;
	assign n_4376 = (~x_330 & ~n_936) ;
	assign n_7988 = (~n_4414 & n_7987) ;
	assign n_4400 = (~n_4398 & ~n_4399) ;
	assign n_4393 = (~x_328 & n_4391) ;
	assign n_4392 = (x_328 & ~n_4391) ;
	assign n_4385 = (~n_4382 & n_4384) ;
	assign n_4377 = (i_5 & ~n_4376) ;
	assign n_4375 = (~i_8 & n_936) ;
	assign n_4369 = (i_38 & n_64) ;
	assign n_7989 = (~n_4400 & n_7988) ;
	assign n_4394 = (~n_4392 & ~n_4393) ;
	assign n_4387 = (~x_329 & ~n_4385) ;
	assign n_4386 = (x_329 & n_4385) ;
	assign n_4378 = (~n_4375 & n_4377) ;
	assign n_4370 = (n_66 & n_4369) ;
	assign n_4368 = (x_331 & n_978) ;
	assign n_4361 = (x_332 & ~x_664) ;
	assign n_7990 = (~n_4394 & n_7989) ;
	assign n_4388 = (~n_4386 & ~n_4387) ;
	assign n_4380 = (~x_330 & ~n_4378) ;
	assign n_4379 = (x_330 & n_4378) ;
	assign n_4371 = (~n_4368 & ~n_4370) ;
	assign n_4362 = (~n_527 & ~n_4361) ;
	assign n_4355 = (~x_333 & ~n_630) ;
	assign n_7991 = (~n_4388 & n_7990) ;
	assign n_4381 = (~n_4379 & ~n_4380) ;
	assign n_4373 = (~x_331 & n_4371) ;
	assign n_4372 = (x_331 & ~n_4371) ;
	assign n_4364 = (~n_4362 & n_4363) ;
	assign n_4356 = (i_5 & ~n_4355) ;
	assign n_4354 = (~i_28 & n_630) ;
	assign n_4348 = (i_44 & n_64) ;
	assign n_7992 = (~n_4381 & n_7991) ;
	assign n_4374 = (~n_4372 & ~n_4373) ;
	assign n_4366 = (~x_332 & ~n_4364) ;
	assign n_4365 = (x_332 & n_4364) ;
	assign n_4357 = (~n_4354 & n_4356) ;
	assign n_4349 = (n_66 & n_4348) ;
	assign n_4347 = (x_334 & n_978) ;
	assign n_7993 = (~n_4374 & n_7992) ;
	assign n_4367 = (~n_4365 & ~n_4366) ;
	assign n_4359 = (~x_333 & ~n_4357) ;
	assign n_4358 = (x_333 & n_4357) ;
	assign n_4350 = (~n_4347 & ~n_4349) ;
	assign n_4342 = (~n_139 & n_35) ;
	assign n_4341 = (x_335 & n_36) ;
	assign n_4335 = (i_17 & n_59) ;
	assign n_4299 = (~x_612 & n_153) ;
	assign n_4298 = (x_612 & ~n_153) ;
	assign n_7994 = (~n_4367 & n_7993) ;
	assign n_4360 = (~n_4358 & ~n_4359) ;
	assign n_4352 = (~x_334 & n_4350) ;
	assign n_4351 = (x_334 & ~n_4350) ;
	assign n_4343 = (~n_4341 & ~n_4342) ;
	assign n_4336 = (n_66 & n_4335) ;
	assign n_4334 = (x_336 & n_60) ;
	assign n_4328 = (~x_337 & ~n_697) ;
	assign n_1234 = (~n_1 & ~n_527) ;
	assign n_4300 = (~n_4298 & ~n_4299) ;
	assign n_4297 = (~n_144 & ~n_145) ;
	assign n_4267 = (~n_253 & ~n_254) ;
	assign n_7995 = (~n_4360 & n_7994) ;
	assign n_4353 = (~n_4351 & ~n_4352) ;
	assign n_4345 = (~x_335 & n_4343) ;
	assign n_4344 = (x_335 & ~n_4343) ;
	assign n_4337 = (~n_4334 & ~n_4336) ;
	assign n_4329 = (i_5 & ~n_4328) ;
	assign n_4327 = (~x_659 & n_697) ;
	assign n_4306 = (~n_1605 & ~n_1234) ;
	assign n_4302 = (n_4297 & n_4300) ;
	assign n_4269 = (~x_232 & ~n_4267) ;
	assign n_7996 = (~n_4353 & n_7995) ;
	assign n_4346 = (~n_4344 & ~n_4345) ;
	assign n_4339 = (~x_336 & n_4337) ;
	assign n_4338 = (x_336 & ~n_4337) ;
	assign n_4330 = (~n_4327 & n_4329) ;
	assign n_4322 = (x_419 & n_35) ;
	assign n_4321 = (x_338 & n_36) ;
	assign n_4315 = (~x_339 & ~n_936) ;
	assign n_4307 = (~n_143 & ~n_4306) ;
	assign n_4305 = (i_11 & n_7) ;
	assign n_4303 = (n_527 & ~n_4302) ;
	assign n_4301 = (~n_4297 & ~n_4300) ;
	assign n_4270 = (~x_332 & ~n_4269) ;
	assign n_4268 = (x_232 & n_4267) ;
	assign n_4244 = (~n_313 & ~n_314) ;
	assign n_7997 = (~n_4346 & n_7996) ;
	assign n_4340 = (~n_4338 & ~n_4339) ;
	assign n_4332 = (~x_337 & ~n_4330) ;
	assign n_4331 = (x_337 & n_4330) ;
	assign n_4323 = (~n_4321 & ~n_4322) ;
	assign n_4316 = (i_5 & ~n_4315) ;
	assign n_4314 = (~i_41 & n_936) ;
	assign n_4308 = (~n_4305 & ~n_4307) ;
	assign n_4304 = (~n_4301 & n_4303) ;
	assign n_4271 = (~n_4268 & n_4270) ;
	assign n_4246 = (~x_80 & ~n_4244) ;
	assign n_7998 = (~n_4340 & n_7997) ;
	assign n_4333 = (~n_4331 & ~n_4332) ;
	assign n_4325 = (~x_338 & n_4323) ;
	assign n_4324 = (x_338 & ~n_4323) ;
	assign n_4317 = (~n_4314 & n_4316) ;
	assign n_4309 = (~n_4304 & n_4308) ;
	assign n_4273 = (n_257 & ~n_4271) ;
	assign n_4247 = (~x_332 & ~n_4246) ;
	assign n_4245 = (x_80 & n_4244) ;
	assign n_7999 = (~n_4333 & n_7998) ;
	assign n_4326 = (~n_4324 & ~n_4325) ;
	assign n_4319 = (~x_339 & ~n_4317) ;
	assign n_4318 = (x_339 & n_4317) ;
	assign n_4310 = (i_5 & ~n_4309) ;
	assign n_4292 = (n_1009 & ~n_467) ;
	assign n_4291 = (x_341 & n_1007) ;
	assign n_4285 = (i_26 & n_64) ;
	assign n_4277 = (~n_257 & ~n_1606) ;
	assign n_4276 = (i_46 & n_7) ;
	assign n_4274 = (x_664 & ~n_4273) ;
	assign n_4272 = (~n_257 & n_4271) ;
	assign n_4248 = (~n_4245 & n_4247) ;
	assign n_8000 = (~n_4326 & n_7999) ;
	assign n_4320 = (~n_4318 & ~n_4319) ;
	assign n_4312 = (~x_340 & ~n_4310) ;
	assign n_4311 = (x_340 & n_4310) ;
	assign n_4293 = (~n_4291 & ~n_4292) ;
	assign n_4286 = (n_66 & n_4285) ;
	assign n_4284 = (x_342 & n_978) ;
	assign n_4278 = (~n_4276 & ~n_4277) ;
	assign n_4275 = (~n_4272 & n_4274) ;
	assign n_4250 = (n_317 & ~n_4248) ;
	assign n_8001 = (~n_4320 & n_8000) ;
	assign n_4313 = (~n_4311 & ~n_4312) ;
	assign n_4295 = (~x_341 & n_4293) ;
	assign n_4294 = (x_341 & ~n_4293) ;
	assign n_4287 = (~n_4284 & ~n_4286) ;
	assign n_4279 = (~n_4275 & n_4278) ;
	assign n_4254 = (~n_317 & ~n_1606) ;
	assign n_4253 = (i_33 & n_7) ;
	assign n_4251 = (x_664 & ~n_4250) ;
	assign n_4249 = (~n_317 & n_4248) ;
	assign n_8002 = (~n_4313 & n_8001) ;
	assign n_4296 = (~n_4294 & ~n_4295) ;
	assign n_4289 = (~x_342 & n_4287) ;
	assign n_4288 = (x_342 & ~n_4287) ;
	assign n_4280 = (i_5 & ~n_4279) ;
	assign n_4262 = (x_539 & n_53) ;
	assign n_4261 = (x_344 & n_51) ;
	assign n_4255 = (~n_4253 & ~n_4254) ;
	assign n_4252 = (~n_4249 & n_4251) ;
	assign n_8003 = (~n_4296 & n_8002) ;
	assign n_4290 = (~n_4288 & ~n_4289) ;
	assign n_4282 = (~x_343 & ~n_4280) ;
	assign n_4281 = (x_343 & n_4280) ;
	assign n_4263 = (~n_4261 & ~n_4262) ;
	assign n_4256 = (~n_4252 & n_4255) ;
	assign n_4238 = (i_32 & n_64) ;
	assign n_8004 = (~n_4290 & n_8003) ;
	assign n_4283 = (~n_4281 & ~n_4282) ;
	assign n_4265 = (~x_344 & n_4263) ;
	assign n_4264 = (x_344 & ~n_4263) ;
	assign n_4257 = (i_5 & ~n_4256) ;
	assign n_4239 = (n_66 & n_4238) ;
	assign n_4237 = (x_346 & n_978) ;
	assign n_8005 = (~n_4283 & n_8004) ;
	assign n_4266 = (~n_4264 & ~n_4265) ;
	assign n_4259 = (~x_345 & ~n_4257) ;
	assign n_4258 = (x_345 & n_4257) ;
	assign n_4240 = (~n_4237 & ~n_4239) ;
	assign n_4232 = (x_391 & n_53) ;
	assign n_4231 = (x_347 & n_51) ;
	assign n_4225 = (~x_348 & ~n_544) ;
	assign n_4217 = (i_21 & n_669) ;
	assign n_4216 = (x_793 & n_662) ;
	assign n_8006 = (~n_4266 & n_8005) ;
	assign n_4260 = (~n_4258 & ~n_4259) ;
	assign n_4242 = (~x_346 & n_4240) ;
	assign n_4241 = (x_346 & ~n_4240) ;
	assign n_4233 = (~n_4231 & ~n_4232) ;
	assign n_4226 = (i_5 & ~n_4225) ;
	assign n_4224 = (~i_53 & n_544) ;
	assign n_4218 = (~n_4216 & ~n_4217) ;
	assign n_4215 = (x_349 & ~n_665) ;
	assign n_8007 = (~n_4260 & n_8006) ;
	assign n_4243 = (~n_4241 & ~n_4242) ;
	assign n_4235 = (~x_347 & n_4233) ;
	assign n_4234 = (x_347 & ~n_4233) ;
	assign n_4227 = (~n_4224 & n_4226) ;
	assign n_4219 = (~n_4215 & n_4218) ;
	assign n_8008 = (~n_4243 & n_8007) ;
	assign n_4236 = (~n_4234 & ~n_4235) ;
	assign n_4229 = (~x_348 & ~n_4227) ;
	assign n_4228 = (x_348 & n_4227) ;
	assign n_4220 = (i_5 & ~n_4219) ;
	assign n_4210 = (n_1009 & ~n_511) ;
	assign n_4209 = (x_350 & n_1007) ;
	assign n_8009 = (~n_4236 & n_8008) ;
	assign n_4230 = (~n_4228 & ~n_4229) ;
	assign n_4222 = (~x_349 & ~n_4220) ;
	assign n_4221 = (x_349 & n_4220) ;
	assign n_4211 = (~n_4209 & ~n_4210) ;
	assign n_4204 = (x_610 & n_53) ;
	assign n_4203 = (x_351 & n_51) ;
	assign n_8010 = (~n_4230 & n_8009) ;
	assign n_4223 = (~n_4221 & ~n_4222) ;
	assign n_4213 = (~x_350 & n_4211) ;
	assign n_4212 = (x_350 & ~n_4211) ;
	assign n_4205 = (~n_4203 & ~n_4204) ;
	assign n_4198 = (~n_218 & n_1009) ;
	assign n_4197 = (x_352 & n_1007) ;
	assign n_4191 = (i_47 & n_59) ;
	assign n_8011 = (~n_4223 & n_8010) ;
	assign n_4214 = (~n_4212 & ~n_4213) ;
	assign n_4207 = (~x_351 & n_4205) ;
	assign n_4206 = (x_351 & ~n_4205) ;
	assign n_4199 = (~n_4197 & ~n_4198) ;
	assign n_4192 = (n_66 & n_4191) ;
	assign n_4190 = (x_353 & n_60) ;
	assign n_4184 = (~x_354 & ~n_936) ;
	assign n_4138 = (~x_207 & n_773) ;
	assign n_4137 = (x_207 & ~n_773) ;
	assign n_8012 = (~n_4214 & n_8011) ;
	assign n_4208 = (~n_4206 & ~n_4207) ;
	assign n_4201 = (~x_352 & n_4199) ;
	assign n_4200 = (x_352 & ~n_4199) ;
	assign n_4193 = (~n_4190 & ~n_4192) ;
	assign n_4185 = (i_5 & ~n_4184) ;
	assign n_4183 = (~i_45 & n_936) ;
	assign n_4139 = (~n_4137 & ~n_4138) ;
	assign n_4136 = (~n_763 & ~n_764) ;
	assign n_8013 = (~n_4208 & n_8012) ;
	assign n_4202 = (~n_4200 & ~n_4201) ;
	assign n_4195 = (~x_353 & n_4193) ;
	assign n_4194 = (x_353 & ~n_4193) ;
	assign n_4186 = (~n_4183 & n_4185) ;
	assign n_4178 = (i_35 & n_948) ;
	assign n_4177 = (x_355 & n_945) ;
	assign n_4171 = (~x_356 & ~n_544) ;
	assign n_4148 = (~x_359 & n_6) ;
	assign n_4141 = (n_4136 & ~n_4139) ;
	assign n_8014 = (~n_4202 & n_8013) ;
	assign n_4196 = (~n_4194 & ~n_4195) ;
	assign n_4188 = (~x_354 & ~n_4186) ;
	assign n_4187 = (x_354 & n_4186) ;
	assign n_4179 = (~n_4177 & ~n_4178) ;
	assign n_4172 = (i_5 & ~n_4171) ;
	assign n_4170 = (~i_25 & n_544) ;
	assign n_4149 = (~n_4147 & ~n_4148) ;
	assign n_4144 = (x_359 & ~n_697) ;
	assign n_4142 = (n_697 & ~n_4141) ;
	assign n_4140 = (~n_4136 & n_4139) ;
	assign n_8015 = (~n_4196 & n_8014) ;
	assign n_4189 = (~n_4187 & ~n_4188) ;
	assign n_4181 = (~x_355 & n_4179) ;
	assign n_4180 = (x_355 & ~n_4179) ;
	assign n_4173 = (~n_4170 & n_4172) ;
	assign n_4165 = (i_38 & n_948) ;
	assign n_4164 = (x_357 & n_945) ;
	assign n_4158 = (~x_358 & ~n_544) ;
	assign n_4150 = (n_629 & ~n_4149) ;
	assign n_4145 = (~n_629 & ~n_4144) ;
	assign n_4143 = (~n_4140 & n_4142) ;
	assign n_8016 = (~n_4189 & n_8015) ;
	assign n_4182 = (~n_4180 & ~n_4181) ;
	assign n_4175 = (~x_356 & ~n_4173) ;
	assign n_4174 = (x_356 & n_4173) ;
	assign n_4166 = (~n_4164 & ~n_4165) ;
	assign n_4159 = (i_5 & ~n_4158) ;
	assign n_4157 = (~i_63 & n_544) ;
	assign n_4151 = (n_902 & ~n_4150) ;
	assign n_4146 = (~n_4143 & n_4145) ;
	assign n_8017 = (~n_4182 & n_8016) ;
	assign n_4176 = (~n_4174 & ~n_4175) ;
	assign n_4168 = (~x_357 & n_4166) ;
	assign n_4167 = (x_357 & ~n_4166) ;
	assign n_4160 = (~n_4157 & n_4159) ;
	assign n_4152 = (~n_4146 & n_4151) ;
	assign n_4135 = (x_359 & n_699) ;
	assign n_4129 = (i_15 & n_59) ;
	assign n_8018 = (~n_4176 & n_8017) ;
	assign n_4169 = (~n_4167 & ~n_4168) ;
	assign n_4162 = (~x_358 & ~n_4160) ;
	assign n_4161 = (x_358 & n_4160) ;
	assign n_4153 = (~n_4135 & ~n_4152) ;
	assign n_4130 = (n_66 & n_4129) ;
	assign n_4128 = (x_360 & n_60) ;
	assign n_4122 = (~x_361 & ~n_936) ;
	assign n_8019 = (~n_4169 & n_8018) ;
	assign n_4163 = (~n_4161 & ~n_4162) ;
	assign n_4155 = (~x_359 & n_4153) ;
	assign n_4154 = (x_359 & ~n_4153) ;
	assign n_4131 = (~n_4128 & ~n_4130) ;
	assign n_4123 = (i_5 & ~n_4122) ;
	assign n_4121 = (~i_25 & n_936) ;
	assign n_8020 = (~n_4163 & n_8019) ;
	assign n_4156 = (~n_4154 & ~n_4155) ;
	assign n_4133 = (~x_360 & n_4131) ;
	assign n_4132 = (x_360 & ~n_4131) ;
	assign n_4124 = (~n_4121 & n_4123) ;
	assign n_4116 = (x_302 & n_53) ;
	assign n_4115 = (x_362 & n_51) ;
	assign n_4109 = (~x_363 & ~n_697) ;
	assign n_4086 = (x_366 & ~n_14) ;
	assign n_8021 = (~n_4156 & n_8020) ;
	assign n_4134 = (~n_4132 & ~n_4133) ;
	assign n_4126 = (~x_361 & ~n_4124) ;
	assign n_4125 = (x_361 & n_4124) ;
	assign n_4117 = (~n_4115 & ~n_4116) ;
	assign n_4110 = (i_5 & ~n_4109) ;
	assign n_4108 = (~x_307 & n_697) ;
	assign n_4102 = (~x_364 & ~n_630) ;
	assign n_4087 = (n_12 & ~n_4086) ;
	assign n_4085 = (x_419 & n_14) ;
	assign n_4082 = (x_419 & n_11) ;
	assign n_8022 = (~n_4134 & n_8021) ;
	assign n_4127 = (~n_4125 & ~n_4126) ;
	assign n_4119 = (~x_362 & n_4117) ;
	assign n_4118 = (x_362 & ~n_4117) ;
	assign n_4111 = (~n_4108 & n_4110) ;
	assign n_4103 = (i_5 & ~n_4102) ;
	assign n_4101 = (~i_22 & n_630) ;
	assign n_4088 = (~n_4085 & n_4087) ;
	assign n_4083 = (x_168 & ~n_4082) ;
	assign n_4081 = (x_366 & ~n_11) ;
	assign n_4078 = (x_366 & n_6) ;
	assign n_4039 = (~x_648 & n_4037) ;
	assign n_4038 = (x_648 & ~n_4037) ;
	assign n_8023 = (~n_4127 & n_8022) ;
	assign n_4120 = (~n_4118 & ~n_4119) ;
	assign n_4113 = (~x_363 & ~n_4111) ;
	assign n_4112 = (x_363 & n_4111) ;
	assign n_4104 = (~n_4101 & n_4103) ;
	assign n_4096 = (i_12 & n_948) ;
	assign n_4095 = (x_365 & n_945) ;
	assign n_4089 = (i_5 & ~n_4088) ;
	assign n_4084 = (~n_4081 & n_4083) ;
	assign n_4079 = (n_1 & ~n_4078) ;
	assign n_4077 = (i_66 & ~n_6) ;
	assign n_4040 = (~n_4038 & ~n_4039) ;
	assign n_4028 = (~n_4026 & ~n_4027) ;
	assign n_8024 = (~n_4120 & n_8023) ;
	assign n_4114 = (~n_4112 & ~n_4113) ;
	assign n_4106 = (~x_364 & ~n_4104) ;
	assign n_4105 = (x_364 & n_4104) ;
	assign n_4097 = (~n_4095 & ~n_4096) ;
	assign n_4090 = (~n_4084 & n_4089) ;
	assign n_4080 = (~n_4077 & n_4079) ;
	assign n_4071 = (~x_367 & ~n_630) ;
	assign n_4048 = (~x_370 & n_6) ;
	assign n_535 = (~i_54 & ~n_6) ;
	assign n_4042 = (n_4028 & ~n_4040) ;
	assign n_8025 = (~n_4114 & n_8024) ;
	assign n_4107 = (~n_4105 & ~n_4106) ;
	assign n_4099 = (~x_365 & n_4097) ;
	assign n_4098 = (x_365 & ~n_4097) ;
	assign n_4091 = (~n_4080 & n_4090) ;
	assign n_4072 = (i_5 & ~n_4071) ;
	assign n_4070 = (~i_11 & n_630) ;
	assign n_4049 = (~n_535 & ~n_4048) ;
	assign n_4045 = (x_370 & ~n_697) ;
	assign n_4043 = (n_697 & ~n_4042) ;
	assign n_4041 = (~n_4028 & n_4040) ;
	assign n_8026 = (~n_4107 & n_8025) ;
	assign n_4100 = (~n_4098 & ~n_4099) ;
	assign n_4093 = (~x_366 & ~n_4091) ;
	assign n_4092 = (x_366 & n_4091) ;
	assign n_4073 = (~n_4070 & n_4072) ;
	assign n_4065 = (x_699 & n_53) ;
	assign n_4064 = (x_368 & n_51) ;
	assign n_4058 = (~x_369 & ~n_544) ;
	assign n_4050 = (n_629 & ~n_4049) ;
	assign n_4046 = (~n_629 & ~n_4045) ;
	assign n_4044 = (~n_4041 & n_4043) ;
	assign n_8027 = (~n_4100 & n_8026) ;
	assign n_4094 = (~n_4092 & ~n_4093) ;
	assign n_4075 = (~x_367 & ~n_4073) ;
	assign n_4074 = (x_367 & n_4073) ;
	assign n_4066 = (~n_4064 & ~n_4065) ;
	assign n_4059 = (i_5 & ~n_4058) ;
	assign n_4057 = (~i_47 & n_544) ;
	assign n_4051 = (n_902 & ~n_4050) ;
	assign n_4047 = (~n_4044 & n_4046) ;
	assign n_8028 = (~n_4094 & n_8027) ;
	assign n_4076 = (~n_4074 & ~n_4075) ;
	assign n_4068 = (~x_368 & n_4066) ;
	assign n_4067 = (x_368 & ~n_4066) ;
	assign n_4060 = (~n_4057 & n_4059) ;
	assign n_4052 = (~n_4047 & n_4051) ;
	assign n_4010 = (x_370 & n_699) ;
	assign n_4004 = (~x_371 & ~n_936) ;
	assign n_3957 = (~x_636 & n_2863) ;
	assign n_3956 = (x_636 & ~n_2863) ;
	assign n_8029 = (~n_4076 & n_8028) ;
	assign n_4069 = (~n_4067 & ~n_4068) ;
	assign n_4062 = (~x_369 & ~n_4060) ;
	assign n_4061 = (x_369 & n_4060) ;
	assign n_4053 = (~n_4010 & ~n_4052) ;
	assign n_4005 = (i_5 & ~n_4004) ;
	assign n_4003 = (~i_52 & n_936) ;
	assign n_3958 = (~n_3956 & ~n_3957) ;
	assign n_3955 = (~n_2853 & ~n_2854) ;
	assign n_8030 = (~n_4069 & n_8029) ;
	assign n_4063 = (~n_4061 & ~n_4062) ;
	assign n_4055 = (~x_370 & n_4053) ;
	assign n_4054 = (x_370 & ~n_4053) ;
	assign n_4006 = (~n_4003 & n_4005) ;
	assign n_3998 = (~n_218 & n_35) ;
	assign n_3997 = (x_372 & n_36) ;
	assign n_3991 = (i_25 & n_59) ;
	assign n_3967 = (~x_376 & n_6) ;
	assign n_3960 = (n_3955 & ~n_3958) ;
	assign n_8031 = (~n_4063 & n_8030) ;
	assign n_4056 = (~n_4054 & ~n_4055) ;
	assign n_4008 = (~x_371 & ~n_4006) ;
	assign n_4007 = (x_371 & n_4006) ;
	assign n_3999 = (~n_3997 & ~n_3998) ;
	assign n_3992 = (n_66 & n_3991) ;
	assign n_3990 = (x_373 & n_60) ;
	assign n_3984 = (i_58 & n_64) ;
	assign n_3968 = (~n_3966 & ~n_3967) ;
	assign n_3963 = (x_376 & ~n_697) ;
	assign n_3961 = (n_697 & ~n_3960) ;
	assign n_3959 = (~n_3955 & n_3958) ;
	assign n_8032 = (~n_4056 & n_8031) ;
	assign n_4009 = (~n_4007 & ~n_4008) ;
	assign n_4001 = (~x_372 & n_3999) ;
	assign n_4000 = (x_372 & ~n_3999) ;
	assign n_3993 = (~n_3990 & ~n_3992) ;
	assign n_3985 = (n_66 & n_3984) ;
	assign n_3983 = (x_374 & n_978) ;
	assign n_3977 = (i_59 & n_64) ;
	assign n_3969 = (n_629 & ~n_3968) ;
	assign n_3964 = (~n_629 & ~n_3963) ;
	assign n_3962 = (~n_3959 & n_3961) ;
	assign n_8033 = (~n_4009 & n_8032) ;
	assign n_4002 = (~n_4000 & ~n_4001) ;
	assign n_3995 = (~x_373 & n_3993) ;
	assign n_3994 = (x_373 & ~n_3993) ;
	assign n_3986 = (~n_3983 & ~n_3985) ;
	assign n_3978 = (n_66 & n_3977) ;
	assign n_3976 = (x_375 & n_978) ;
	assign n_3970 = (n_902 & ~n_3969) ;
	assign n_3965 = (~n_3962 & n_3964) ;
	assign n_8034 = (~n_4002 & n_8033) ;
	assign n_3996 = (~n_3994 & ~n_3995) ;
	assign n_3988 = (~x_374 & n_3986) ;
	assign n_3987 = (x_374 & ~n_3986) ;
	assign n_3979 = (~n_3976 & ~n_3978) ;
	assign n_3971 = (~n_3965 & n_3970) ;
	assign n_3954 = (x_376 & n_699) ;
	assign n_3948 = (~x_377 & ~n_630) ;
	assign n_8035 = (~n_3996 & n_8034) ;
	assign n_3989 = (~n_3987 & ~n_3988) ;
	assign n_3981 = (~x_375 & n_3979) ;
	assign n_3980 = (x_375 & ~n_3979) ;
	assign n_3972 = (~n_3954 & ~n_3971) ;
	assign n_3949 = (i_5 & ~n_3948) ;
	assign n_3947 = (~i_30 & n_630) ;
	assign n_8036 = (~n_3989 & n_8035) ;
	assign n_3982 = (~n_3980 & ~n_3981) ;
	assign n_3974 = (~x_376 & n_3972) ;
	assign n_3973 = (x_376 & ~n_3972) ;
	assign n_3950 = (~n_3947 & n_3949) ;
	assign n_3942 = (x_264 & n_35) ;
	assign n_3941 = (x_378 & n_36) ;
	assign n_8037 = (~n_3982 & n_8036) ;
	assign n_3975 = (~n_3973 & ~n_3974) ;
	assign n_3952 = (~x_377 & ~n_3950) ;
	assign n_3951 = (x_377 & n_3950) ;
	assign n_3943 = (~n_3941 & ~n_3942) ;
	assign n_3936 = (i_68 & n_3935) ;
	assign n_3934 = (x_379 & n_3933) ;
	assign n_3927 = (~x_380 & ~n_544) ;
	assign n_8038 = (~n_3975 & n_8037) ;
	assign n_3953 = (~n_3951 & ~n_3952) ;
	assign n_3945 = (~x_378 & n_3943) ;
	assign n_3944 = (x_378 & ~n_3943) ;
	assign n_3937 = (~n_3934 & ~n_3936) ;
	assign n_3928 = (i_5 & ~n_3927) ;
	assign n_3926 = (~i_41 & n_544) ;
	assign n_3920 = (~x_381 & ~n_630) ;
	assign n_3912 = (~i_48 & n_669) ;
	assign n_3910 = (~x_117 & ~n_544) ;
	assign n_8039 = (~n_3953 & n_8038) ;
	assign n_3946 = (~n_3944 & ~n_3945) ;
	assign n_3939 = (~x_379 & n_3937) ;
	assign n_3938 = (x_379 & ~n_3937) ;
	assign n_3929 = (~n_3926 & n_3928) ;
	assign n_3921 = (i_5 & ~n_3920) ;
	assign n_3919 = (~i_44 & n_630) ;
	assign n_3913 = (i_5 & ~n_3912) ;
	assign n_3911 = (n_662 & n_3910) ;
	assign n_3902 = (~i_29 & n_669) ;
	assign n_3900 = (~x_758 & ~n_544) ;
	assign n_8040 = (~n_3946 & n_8039) ;
	assign n_3940 = (~n_3938 & ~n_3939) ;
	assign n_3931 = (~x_380 & ~n_3929) ;
	assign n_3930 = (x_380 & n_3929) ;
	assign n_3922 = (~n_3919 & n_3921) ;
	assign n_3914 = (~n_3911 & n_3913) ;
	assign n_3909 = (~x_382 & ~n_665) ;
	assign n_3903 = (i_5 & ~n_3902) ;
	assign n_3901 = (n_662 & n_3900) ;
	assign n_8041 = (~n_3940 & n_8040) ;
	assign n_3932 = (~n_3930 & ~n_3931) ;
	assign n_3924 = (~x_381 & ~n_3922) ;
	assign n_3923 = (x_381 & n_3922) ;
	assign n_3915 = (~n_3909 & n_3914) ;
	assign n_3904 = (~n_3901 & n_3903) ;
	assign n_3899 = (~x_383 & ~n_665) ;
	assign n_3893 = (~x_384 & ~n_630) ;
	assign n_8042 = (~n_3932 & n_8041) ;
	assign n_3925 = (~n_3923 & ~n_3924) ;
	assign n_3917 = (~x_382 & ~n_3915) ;
	assign n_3916 = (x_382 & n_3915) ;
	assign n_3905 = (~n_3899 & n_3904) ;
	assign n_3894 = (i_5 & ~n_3893) ;
	assign n_3892 = (~i_66 & n_630) ;
	assign n_3886 = (i_57 & n_64) ;
	assign n_3813 = (x_223 & n_133) ;
	assign n_3812 = (~x_223 & ~n_133) ;
	assign n_8043 = (~n_3925 & n_8042) ;
	assign n_3918 = (~n_3916 & ~n_3917) ;
	assign n_3907 = (~x_383 & ~n_3905) ;
	assign n_3906 = (x_383 & n_3905) ;
	assign n_3895 = (~n_3892 & n_3894) ;
	assign n_3887 = (n_66 & n_3886) ;
	assign n_3885 = (x_385 & n_978) ;
	assign n_3834 = (~x_542 & n_747) ;
	assign n_3833 = (x_542 & ~n_747) ;
	assign n_3814 = (~n_3812 & ~n_3813) ;
	assign n_8044 = (~n_3918 & n_8043) ;
	assign n_3908 = (~n_3906 & ~n_3907) ;
	assign n_3897 = (~x_384 & ~n_3895) ;
	assign n_3896 = (x_384 & n_3895) ;
	assign n_3888 = (~n_3885 & ~n_3887) ;
	assign n_3880 = (x_254 & n_35) ;
	assign n_3879 = (x_386 & n_36) ;
	assign n_3873 = (~x_387 & ~n_936) ;
	assign n_3835 = (~n_3833 & ~n_3834) ;
	assign n_3832 = (~n_737 & ~n_738) ;
	assign n_3816 = (n_155 & ~n_3814) ;
	assign n_8045 = (~n_3908 & n_8044) ;
	assign n_3898 = (~n_3896 & ~n_3897) ;
	assign n_3890 = (~x_385 & n_3888) ;
	assign n_3889 = (x_385 & ~n_3888) ;
	assign n_3881 = (~n_3879 & ~n_3880) ;
	assign n_3874 = (i_5 & ~n_3873) ;
	assign n_3872 = (~i_65 & n_936) ;
	assign n_3844 = (i_30 & ~n_6) ;
	assign n_3837 = (n_3832 & ~n_3835) ;
	assign n_3817 = (~x_332 & ~n_3816) ;
	assign n_3815 = (~n_155 & n_3814) ;
	assign n_8046 = (~n_3898 & n_8045) ;
	assign n_3891 = (~n_3889 & ~n_3890) ;
	assign n_3883 = (~x_386 & n_3881) ;
	assign n_3882 = (x_386 & ~n_3881) ;
	assign n_3875 = (~n_3872 & n_3874) ;
	assign n_3867 = (~n_347 & n_35) ;
	assign n_3866 = (x_388 & n_36) ;
	assign n_3845 = (n_629 & ~n_3844) ;
	assign n_3843 = (x_391 & n_6) ;
	assign n_3840 = (x_391 & ~n_697) ;
	assign n_3838 = (n_697 & ~n_3837) ;
	assign n_3836 = (~n_3832 & n_3835) ;
	assign n_3818 = (~n_3815 & n_3817) ;
	assign n_8047 = (~n_3891 & n_8046) ;
	assign n_3884 = (~n_3882 & ~n_3883) ;
	assign n_3877 = (~x_387 & ~n_3875) ;
	assign n_3876 = (x_387 & n_3875) ;
	assign n_3868 = (~n_3866 & ~n_3867) ;
	assign n_3861 = (n_1009 & ~n_75) ;
	assign n_3860 = (x_389 & n_1007) ;
	assign n_3854 = (i_63 & n_59) ;
	assign n_3846 = (~n_3843 & n_3845) ;
	assign n_3841 = (~n_629 & ~n_3840) ;
	assign n_3839 = (~n_3836 & n_3838) ;
	assign n_3820 = (n_136 & ~n_3818) ;
	assign n_3775 = (~n_238 & ~n_239) ;
	assign n_8048 = (~n_3884 & n_8047) ;
	assign n_3878 = (~n_3876 & ~n_3877) ;
	assign n_3870 = (~x_388 & n_3868) ;
	assign n_3869 = (x_388 & ~n_3868) ;
	assign n_3862 = (~n_3860 & ~n_3861) ;
	assign n_3855 = (n_66 & n_3854) ;
	assign n_3853 = (x_390 & n_60) ;
	assign n_3847 = (n_902 & ~n_3846) ;
	assign n_3842 = (~n_3839 & n_3841) ;
	assign n_3824 = (~n_136 & ~n_1606) ;
	assign n_3823 = (i_55 & n_7) ;
	assign n_3821 = (x_664 & ~n_3820) ;
	assign n_3819 = (~n_136 & n_3818) ;
	assign n_3777 = (~x_316 & ~n_3775) ;
	assign n_8049 = (~n_3878 & n_8048) ;
	assign n_3871 = (~n_3869 & ~n_3870) ;
	assign n_3864 = (~x_389 & n_3862) ;
	assign n_3863 = (x_389 & ~n_3862) ;
	assign n_3856 = (~n_3853 & ~n_3855) ;
	assign n_3848 = (~n_3842 & n_3847) ;
	assign n_3831 = (x_391 & n_699) ;
	assign n_3825 = (~n_3823 & ~n_3824) ;
	assign n_3822 = (~n_3819 & n_3821) ;
	assign n_3778 = (~x_332 & ~n_3777) ;
	assign n_3776 = (x_316 & n_3775) ;
	assign n_3749 = (~n_298 & ~n_299) ;
	assign n_8050 = (~n_3871 & n_8049) ;
	assign n_3865 = (~n_3863 & ~n_3864) ;
	assign n_3858 = (~x_390 & n_3856) ;
	assign n_3857 = (x_390 & ~n_3856) ;
	assign n_3849 = (~n_3831 & ~n_3848) ;
	assign n_3826 = (~n_3822 & n_3825) ;
	assign n_3806 = (~x_393 & ~n_544) ;
	assign n_3779 = (~n_3776 & n_3778) ;
	assign n_3751 = (~x_169 & ~n_3749) ;
	assign n_8051 = (~n_3865 & n_8050) ;
	assign n_3859 = (~n_3857 & ~n_3858) ;
	assign n_3851 = (~x_391 & n_3849) ;
	assign n_3850 = (x_391 & ~n_3849) ;
	assign n_3827 = (i_5 & ~n_3826) ;
	assign n_3807 = (i_5 & ~n_3806) ;
	assign n_3805 = (~i_35 & n_544) ;
	assign n_3781 = (n_242 & ~n_3779) ;
	assign n_3752 = (~x_332 & ~n_3751) ;
	assign n_3750 = (x_169 & n_3749) ;
	assign n_8052 = (~n_3859 & n_8051) ;
	assign n_3852 = (~n_3850 & ~n_3851) ;
	assign n_3829 = (~x_392 & ~n_3827) ;
	assign n_3828 = (x_392 & n_3827) ;
	assign n_3808 = (~n_3805 & n_3807) ;
	assign n_3800 = (i_4 & n_948) ;
	assign n_3799 = (x_394 & n_945) ;
	assign n_3793 = (i_12 & n_64) ;
	assign n_3785 = (~n_242 & ~n_1606) ;
	assign n_3784 = (i_18 & n_7) ;
	assign n_3782 = (x_664 & ~n_3781) ;
	assign n_3780 = (~n_242 & n_3779) ;
	assign n_3759 = (n_6 & n_302) ;
	assign n_3753 = (~n_3750 & n_3752) ;
	assign n_8053 = (~n_3852 & n_8052) ;
	assign n_3830 = (~n_3828 & ~n_3829) ;
	assign n_3810 = (~x_393 & ~n_3808) ;
	assign n_3809 = (x_393 & n_3808) ;
	assign n_3801 = (~n_3799 & ~n_3800) ;
	assign n_3794 = (n_66 & n_3793) ;
	assign n_3792 = (x_395 & n_978) ;
	assign n_3786 = (~n_3784 & ~n_3785) ;
	assign n_3783 = (~n_3780 & n_3782) ;
	assign n_3760 = (n_1 & ~n_3759) ;
	assign n_1155 = (~i_60 & ~n_6) ;
	assign n_3755 = (n_302 & ~n_3753) ;
	assign n_8054 = (~n_3830 & n_8053) ;
	assign n_3811 = (~n_3809 & ~n_3810) ;
	assign n_3803 = (~x_394 & n_3801) ;
	assign n_3802 = (x_394 & ~n_3801) ;
	assign n_3795 = (~n_3792 & ~n_3794) ;
	assign n_3787 = (~n_3783 & n_3786) ;
	assign n_3769 = (~x_397 & ~n_936) ;
	assign n_3761 = (~n_1155 & n_3760) ;
	assign n_3758 = (n_59 & ~n_302) ;
	assign n_3756 = (x_664 & ~n_3755) ;
	assign n_3754 = (~n_302 & n_3753) ;
	assign n_8055 = (~n_3811 & n_8054) ;
	assign n_3804 = (~n_3802 & ~n_3803) ;
	assign n_3797 = (~x_395 & n_3795) ;
	assign n_3796 = (x_395 & ~n_3795) ;
	assign n_3788 = (i_5 & ~n_3787) ;
	assign n_3770 = (i_5 & ~n_3769) ;
	assign n_3768 = (~i_18 & n_936) ;
	assign n_3762 = (~n_3758 & ~n_3761) ;
	assign n_3757 = (~n_3754 & n_3756) ;
	assign n_8056 = (~n_3804 & n_8055) ;
	assign n_3798 = (~n_3796 & ~n_3797) ;
	assign n_3790 = (~x_396 & ~n_3788) ;
	assign n_3789 = (x_396 & n_3788) ;
	assign n_3771 = (~n_3768 & n_3770) ;
	assign n_3763 = (~n_3757 & n_3762) ;
	assign n_3743 = (i_41 & n_59) ;
	assign n_8057 = (~n_3798 & n_8056) ;
	assign n_3791 = (~n_3789 & ~n_3790) ;
	assign n_3773 = (~x_397 & ~n_3771) ;
	assign n_3772 = (x_397 & n_3771) ;
	assign n_3764 = (i_5 & ~n_3763) ;
	assign n_3744 = (n_66 & n_3743) ;
	assign n_3742 = (x_399 & n_60) ;
	assign n_3736 = (~x_400 & ~n_630) ;
	assign n_8058 = (~n_3791 & n_8057) ;
	assign n_3774 = (~n_3772 & ~n_3773) ;
	assign n_3766 = (~x_398 & ~n_3764) ;
	assign n_3765 = (x_398 & n_3764) ;
	assign n_3745 = (~n_3742 & ~n_3744) ;
	assign n_3737 = (i_5 & ~n_3736) ;
	assign n_3735 = (~i_18 & n_630) ;
	assign n_3722 = (~i_41 & n_669) ;
	assign n_3720 = (~x_178 & ~n_544) ;
	assign n_8059 = (~n_3774 & n_8058) ;
	assign n_3767 = (~n_3765 & ~n_3766) ;
	assign n_3747 = (~x_399 & n_3745) ;
	assign n_3746 = (x_399 & ~n_3745) ;
	assign n_3738 = (~n_3735 & n_3737) ;
	assign n_3730 = (~n_188 & n_1009) ;
	assign n_3729 = (x_401 & n_1007) ;
	assign n_3723 = (i_5 & ~n_3722) ;
	assign n_3721 = (n_662 & n_3720) ;
	assign n_8060 = (~n_3767 & n_8059) ;
	assign n_3748 = (~n_3746 & ~n_3747) ;
	assign n_3740 = (~x_400 & ~n_3738) ;
	assign n_3739 = (x_400 & n_3738) ;
	assign n_3731 = (~n_3729 & ~n_3730) ;
	assign n_3724 = (~n_3721 & n_3723) ;
	assign n_3719 = (~x_402 & ~n_665) ;
	assign n_8061 = (~n_3748 & n_8060) ;
	assign n_3741 = (~n_3739 & ~n_3740) ;
	assign n_3733 = (~x_401 & n_3731) ;
	assign n_3732 = (x_401 & ~n_3731) ;
	assign n_3725 = (~n_3719 & n_3724) ;
	assign n_3714 = (x_117 & n_53) ;
	assign n_3713 = (x_403 & n_51) ;
	assign n_8062 = (~n_3741 & n_8061) ;
	assign n_3734 = (~n_3732 & ~n_3733) ;
	assign n_3727 = (~x_402 & ~n_3725) ;
	assign n_3726 = (x_402 & n_3725) ;
	assign n_3715 = (~n_3713 & ~n_3714) ;
	assign n_3708 = (x_558 & n_53) ;
	assign n_3707 = (x_404 & n_51) ;
	assign n_8063 = (~n_3734 & n_8062) ;
	assign n_3728 = (~n_3726 & ~n_3727) ;
	assign n_3717 = (~x_403 & n_3715) ;
	assign n_3716 = (x_403 & ~n_3715) ;
	assign n_3709 = (~n_3707 & ~n_3708) ;
	assign n_3702 = (x_644 & n_35) ;
	assign n_3701 = (x_405 & n_36) ;
	assign n_3695 = (i_66 & n_64) ;
	assign n_8064 = (~n_3728 & n_8063) ;
	assign n_3718 = (~n_3716 & ~n_3717) ;
	assign n_3711 = (~x_404 & n_3709) ;
	assign n_3710 = (x_404 & ~n_3709) ;
	assign n_3703 = (~n_3701 & ~n_3702) ;
	assign n_3696 = (n_66 & n_3695) ;
	assign n_3694 = (x_406 & n_978) ;
	assign n_3688 = (~x_407 & ~n_697) ;
	assign n_8065 = (~n_3718 & n_8064) ;
	assign n_3712 = (~n_3710 & ~n_3711) ;
	assign n_3705 = (~x_405 & n_3703) ;
	assign n_3704 = (x_405 & ~n_3703) ;
	assign n_3697 = (~n_3694 & ~n_3696) ;
	assign n_3689 = (i_5 & ~n_3688) ;
	assign n_3687 = (~x_166 & n_697) ;
	assign n_8066 = (~n_3712 & n_8065) ;
	assign n_3706 = (~n_3704 & ~n_3705) ;
	assign n_3699 = (~x_406 & n_3697) ;
	assign n_3698 = (x_406 & ~n_3697) ;
	assign n_3690 = (~n_3687 & n_3689) ;
	assign n_3682 = (n_1009 & ~n_482) ;
	assign n_3681 = (x_408 & n_1007) ;
	assign n_3668 = (~i_43 & n_669) ;
	assign n_3666 = (~x_91 & ~n_544) ;
	assign n_8067 = (~n_3706 & n_8066) ;
	assign n_3700 = (~n_3698 & ~n_3699) ;
	assign n_3692 = (~x_407 & ~n_3690) ;
	assign n_3691 = (x_407 & n_3690) ;
	assign n_3683 = (~n_3681 & ~n_3682) ;
	assign n_3676 = (x_806 & n_53) ;
	assign n_3675 = (x_409 & n_51) ;
	assign n_3669 = (i_5 & ~n_3668) ;
	assign n_3667 = (n_662 & n_3666) ;
	assign n_8068 = (~n_3700 & n_8067) ;
	assign n_3693 = (~n_3691 & ~n_3692) ;
	assign n_3685 = (~x_408 & n_3683) ;
	assign n_3684 = (x_408 & ~n_3683) ;
	assign n_3677 = (~n_3675 & ~n_3676) ;
	assign n_3670 = (~n_3667 & n_3669) ;
	assign n_3665 = (~x_410 & ~n_665) ;
	assign n_3659 = (~x_411 & ~n_630) ;
	assign n_8069 = (~n_3693 & n_8068) ;
	assign n_3686 = (~n_3684 & ~n_3685) ;
	assign n_3679 = (~x_409 & n_3677) ;
	assign n_3678 = (x_409 & ~n_3677) ;
	assign n_3671 = (~n_3665 & n_3670) ;
	assign n_3660 = (i_5 & ~n_3659) ;
	assign n_3658 = (~i_12 & n_630) ;
	assign n_3652 = (~x_412 & ~n_630) ;
	assign n_8070 = (~n_3686 & n_8069) ;
	assign n_3680 = (~n_3678 & ~n_3679) ;
	assign n_3673 = (~x_410 & ~n_3671) ;
	assign n_3672 = (x_410 & n_3671) ;
	assign n_3661 = (~n_3658 & n_3660) ;
	assign n_3653 = (i_5 & ~n_3652) ;
	assign n_3651 = (~i_32 & n_630) ;
	assign n_3645 = (i_18 & n_64) ;
	assign n_8071 = (~n_3680 & n_8070) ;
	assign n_3674 = (~n_3672 & ~n_3673) ;
	assign n_3663 = (~x_411 & ~n_3661) ;
	assign n_3662 = (x_411 & n_3661) ;
	assign n_3654 = (~n_3651 & n_3653) ;
	assign n_3646 = (n_66 & n_3645) ;
	assign n_3644 = (x_413 & n_978) ;
	assign n_3638 = (~x_414 & ~n_630) ;
	assign n_8072 = (~n_3674 & n_8071) ;
	assign n_3664 = (~n_3662 & ~n_3663) ;
	assign n_3656 = (~x_412 & ~n_3654) ;
	assign n_3655 = (x_412 & n_3654) ;
	assign n_3647 = (~n_3644 & ~n_3646) ;
	assign n_3639 = (i_5 & ~n_3638) ;
	assign n_3637 = (~i_67 & n_630) ;
	assign n_8073 = (~n_3664 & n_8072) ;
	assign n_3657 = (~n_3655 & ~n_3656) ;
	assign n_3649 = (~x_413 & n_3647) ;
	assign n_3648 = (x_413 & ~n_3647) ;
	assign n_3640 = (~n_3637 & n_3639) ;
	assign n_3632 = (~n_287 & n_35) ;
	assign n_3631 = (x_415 & n_36) ;
	assign n_3625 = (~x_416 & ~n_697) ;
	assign n_8074 = (~n_3657 & n_8073) ;
	assign n_3650 = (~n_3648 & ~n_3649) ;
	assign n_3642 = (~x_414 & ~n_3640) ;
	assign n_3641 = (x_414 & n_3640) ;
	assign n_3633 = (~n_3631 & ~n_3632) ;
	assign n_3626 = (i_5 & ~n_3625) ;
	assign n_3624 = (~x_247 & n_697) ;
	assign n_3618 = (i_13 & n_59) ;
	assign n_8075 = (~n_3650 & n_8074) ;
	assign n_3643 = (~n_3641 & ~n_3642) ;
	assign n_3635 = (~x_415 & n_3633) ;
	assign n_3634 = (x_415 & ~n_3633) ;
	assign n_3627 = (~n_3624 & n_3626) ;
	assign n_3619 = (n_66 & n_3618) ;
	assign n_3617 = (x_417 & n_60) ;
	assign n_8076 = (~n_3643 & n_8075) ;
	assign n_3636 = (~n_3634 & ~n_3635) ;
	assign n_3629 = (~x_416 & ~n_3627) ;
	assign n_3628 = (x_416 & n_3627) ;
	assign n_3620 = (~n_3617 & ~n_3619) ;
	assign n_3612 = (n_1009 & ~n_1223) ;
	assign n_3611 = (x_418 & n_1007) ;
	assign n_8077 = (~n_3636 & n_8076) ;
	assign n_3630 = (~n_3628 & ~n_3629) ;
	assign n_3622 = (~x_417 & n_3620) ;
	assign n_3621 = (x_417 & ~n_3620) ;
	assign n_3613 = (~n_3611 & ~n_3612) ;
	assign n_3606 = (n_1009 & ~n_497) ;
	assign n_3605 = (x_419 & n_1007) ;
	assign n_3599 = (~x_420 & ~n_936) ;
	assign n_3576 = (x_423 & n_6) ;
	assign n_8078 = (~n_3630 & n_8077) ;
	assign n_3623 = (~n_3621 & ~n_3622) ;
	assign n_3615 = (~x_418 & n_3613) ;
	assign n_3614 = (x_418 & ~n_3613) ;
	assign n_3607 = (~n_3605 & ~n_3606) ;
	assign n_3600 = (i_5 & ~n_3599) ;
	assign n_3598 = (~i_37 & n_936) ;
	assign n_3592 = (i_34 & n_64) ;
	assign n_3577 = (n_629 & ~n_3576) ;
	assign n_8079 = (~n_3623 & n_8078) ;
	assign n_3616 = (~n_3614 & ~n_3615) ;
	assign n_3609 = (~x_419 & n_3607) ;
	assign n_3608 = (x_419 & ~n_3607) ;
	assign n_3601 = (~n_3598 & n_3600) ;
	assign n_3593 = (n_66 & n_3592) ;
	assign n_3591 = (x_421 & n_978) ;
	assign n_3578 = (~n_3575 & n_3577) ;
	assign n_8080 = (~n_3616 & n_8079) ;
	assign n_3610 = (~n_3608 & ~n_3609) ;
	assign n_3603 = (~x_420 & ~n_3601) ;
	assign n_3602 = (x_420 & n_3601) ;
	assign n_3594 = (~n_3591 & ~n_3593) ;
	assign n_3586 = (x_793 & n_53) ;
	assign n_3585 = (x_422 & n_51) ;
	assign n_3579 = (i_5 & ~n_3578) ;
	assign n_3574 = (~x_70 & n_662) ;
	assign n_8081 = (~n_3610 & n_8080) ;
	assign n_3604 = (~n_3602 & ~n_3603) ;
	assign n_3596 = (~x_421 & n_3594) ;
	assign n_3595 = (x_421 & ~n_3594) ;
	assign n_3587 = (~n_3585 & ~n_3586) ;
	assign n_3580 = (~n_3574 & n_3579) ;
	assign n_3573 = (~x_423 & n_663) ;
	assign n_3567 = (i_22 & n_64) ;
	assign n_8082 = (~n_3604 & n_8081) ;
	assign n_3597 = (~n_3595 & ~n_3596) ;
	assign n_3589 = (~x_422 & n_3587) ;
	assign n_3588 = (x_422 & ~n_3587) ;
	assign n_3581 = (~n_3573 & n_3580) ;
	assign n_3568 = (n_66 & n_3567) ;
	assign n_3566 = (x_424 & n_978) ;
	assign n_3560 = (~x_425 & ~n_630) ;
	assign n_8083 = (~n_3597 & n_8082) ;
	assign n_3590 = (~n_3588 & ~n_3589) ;
	assign n_3583 = (~x_423 & ~n_3581) ;
	assign n_3582 = (x_423 & n_3581) ;
	assign n_3569 = (~n_3566 & ~n_3568) ;
	assign n_3561 = (i_5 & ~n_3560) ;
	assign n_3559 = (~i_38 & n_630) ;
	assign n_3546 = (~i_25 & n_669) ;
	assign n_3544 = (~x_709 & ~n_544) ;
	assign n_8084 = (~n_3590 & n_8083) ;
	assign n_3584 = (~n_3582 & ~n_3583) ;
	assign n_3571 = (~x_424 & n_3569) ;
	assign n_3570 = (x_424 & ~n_3569) ;
	assign n_3562 = (~n_3559 & n_3561) ;
	assign n_3554 = (x_656 & n_35) ;
	assign n_3553 = (x_426 & n_36) ;
	assign n_3547 = (i_5 & ~n_3546) ;
	assign n_3545 = (n_662 & n_3544) ;
	assign n_3498 = (~x_198 & n_2876) ;
	assign n_3497 = (x_198 & ~n_2876) ;
	assign n_8085 = (~n_3584 & n_8084) ;
	assign n_3572 = (~n_3570 & ~n_3571) ;
	assign n_3564 = (~x_425 & ~n_3562) ;
	assign n_3563 = (x_425 & n_3562) ;
	assign n_3555 = (~n_3553 & ~n_3554) ;
	assign n_3548 = (~n_3545 & n_3547) ;
	assign n_3543 = (~x_427 & ~n_665) ;
	assign n_3537 = (~x_428 & ~n_630) ;
	assign n_3499 = (~n_3497 & ~n_3498) ;
	assign n_3496 = (~n_2866 & ~n_2867) ;
	assign n_8086 = (~n_3572 & n_8085) ;
	assign n_3565 = (~n_3563 & ~n_3564) ;
	assign n_3557 = (~x_426 & n_3555) ;
	assign n_3556 = (x_426 & ~n_3555) ;
	assign n_3549 = (~n_3543 & n_3548) ;
	assign n_3538 = (i_5 & ~n_3537) ;
	assign n_3536 = (~i_7 & n_630) ;
	assign n_3507 = (~x_432 & n_6) ;
	assign n_2266 = (~i_15 & ~n_6) ;
	assign n_3501 = (n_3496 & ~n_3499) ;
	assign n_8087 = (~n_3565 & n_8086) ;
	assign n_3558 = (~n_3556 & ~n_3557) ;
	assign n_3551 = (~x_427 & ~n_3549) ;
	assign n_3550 = (x_427 & n_3549) ;
	assign n_3539 = (~n_3536 & n_3538) ;
	assign n_3531 = (~n_203 & n_1009) ;
	assign n_3530 = (x_429 & n_1007) ;
	assign n_3524 = (i_43 & n_59) ;
	assign n_3508 = (~n_2266 & ~n_3507) ;
	assign n_3504 = (x_432 & ~n_697) ;
	assign n_3502 = (n_697 & ~n_3501) ;
	assign n_3500 = (~n_3496 & n_3499) ;
	assign n_8088 = (~n_3558 & n_8087) ;
	assign n_3552 = (~n_3550 & ~n_3551) ;
	assign n_3541 = (~x_428 & ~n_3539) ;
	assign n_3540 = (x_428 & n_3539) ;
	assign n_3532 = (~n_3530 & ~n_3531) ;
	assign n_3525 = (n_66 & n_3524) ;
	assign n_3523 = (x_430 & n_60) ;
	assign n_3517 = (~x_431 & ~n_936) ;
	assign n_3509 = (n_629 & ~n_3508) ;
	assign n_3505 = (~n_629 & ~n_3504) ;
	assign n_3503 = (~n_3500 & n_3502) ;
	assign n_3457 = (~x_287 & n_760) ;
	assign n_3456 = (x_287 & ~n_760) ;
	assign n_8089 = (~n_3552 & n_8088) ;
	assign n_3542 = (~n_3540 & ~n_3541) ;
	assign n_3534 = (~x_429 & n_3532) ;
	assign n_3533 = (x_429 & ~n_3532) ;
	assign n_3526 = (~n_3523 & ~n_3525) ;
	assign n_3518 = (i_5 & ~n_3517) ;
	assign n_3516 = (~i_32 & n_936) ;
	assign n_3510 = (n_902 & ~n_3509) ;
	assign n_3506 = (~n_3503 & n_3505) ;
	assign n_3458 = (~n_3456 & ~n_3457) ;
	assign n_3455 = (~n_750 & ~n_751) ;
	assign n_8090 = (~n_3542 & n_8089) ;
	assign n_3535 = (~n_3533 & ~n_3534) ;
	assign n_3528 = (~x_430 & n_3526) ;
	assign n_3527 = (x_430 & ~n_3526) ;
	assign n_3519 = (~n_3516 & n_3518) ;
	assign n_3511 = (~n_3506 & n_3510) ;
	assign n_3495 = (x_432 & n_699) ;
	assign n_3489 = (~x_433 & ~n_544) ;
	assign n_3466 = (~x_436 & n_6) ;
	assign n_2735 = (~i_58 & ~n_6) ;
	assign n_3460 = (n_3455 & ~n_3458) ;
	assign n_8091 = (~n_3535 & n_8090) ;
	assign n_3529 = (~n_3527 & ~n_3528) ;
	assign n_3521 = (~x_431 & ~n_3519) ;
	assign n_3520 = (x_431 & n_3519) ;
	assign n_3512 = (~n_3495 & ~n_3511) ;
	assign n_3490 = (i_5 & ~n_3489) ;
	assign n_3488 = (~i_48 & n_544) ;
	assign n_3482 = (~x_434 & ~n_544) ;
	assign n_3467 = (~n_2735 & ~n_3466) ;
	assign n_3463 = (x_436 & ~n_697) ;
	assign n_3461 = (n_697 & ~n_3460) ;
	assign n_3459 = (~n_3455 & n_3458) ;
	assign n_8092 = (~n_3529 & n_8091) ;
	assign n_3522 = (~n_3520 & ~n_3521) ;
	assign n_3514 = (~x_432 & n_3512) ;
	assign n_3513 = (x_432 & ~n_3512) ;
	assign n_3491 = (~n_3488 & n_3490) ;
	assign n_3483 = (i_5 & ~n_3482) ;
	assign n_3481 = (~i_13 & n_544) ;
	assign n_3468 = (n_629 & ~n_3467) ;
	assign n_3464 = (~n_629 & ~n_3463) ;
	assign n_3462 = (~n_3459 & n_3461) ;
	assign n_8093 = (~n_3522 & n_8092) ;
	assign n_3515 = (~n_3513 & ~n_3514) ;
	assign n_3493 = (~x_433 & ~n_3491) ;
	assign n_3492 = (x_433 & n_3491) ;
	assign n_3484 = (~n_3481 & n_3483) ;
	assign n_3476 = (i_56 & n_948) ;
	assign n_3475 = (x_435 & n_945) ;
	assign n_3469 = (n_902 & ~n_3468) ;
	assign n_3465 = (~n_3462 & n_3464) ;
	assign n_3437 = (i_12 & n_1) ;
	assign n_8094 = (~n_3515 & n_8093) ;
	assign n_3494 = (~n_3492 & ~n_3493) ;
	assign n_3486 = (~x_434 & ~n_3484) ;
	assign n_3485 = (x_434 & n_3484) ;
	assign n_3477 = (~n_3475 & ~n_3476) ;
	assign n_3470 = (~n_3465 & n_3469) ;
	assign n_3454 = (x_436 & n_699) ;
	assign n_3441 = (x_418 & ~n_16) ;
	assign n_3440 = (i_12 & n_7) ;
	assign n_3438 = (~n_17 & ~n_3437) ;
	assign n_8095 = (~n_3494 & n_8094) ;
	assign n_3487 = (~n_3485 & ~n_3486) ;
	assign n_3479 = (~x_435 & n_3477) ;
	assign n_3478 = (x_435 & ~n_3477) ;
	assign n_3471 = (~n_3454 & ~n_3470) ;
	assign n_3449 = (x_201 & n_53) ;
	assign n_3448 = (x_437 & n_51) ;
	assign n_3442 = (~n_3440 & ~n_3441) ;
	assign n_3439 = (x_438 & ~n_3438) ;
	assign n_8096 = (~n_3487 & n_8095) ;
	assign n_3480 = (~n_3478 & ~n_3479) ;
	assign n_3473 = (~x_436 & n_3471) ;
	assign n_3472 = (x_436 & ~n_3471) ;
	assign n_3450 = (~n_3448 & ~n_3449) ;
	assign n_3443 = (~n_3439 & n_3442) ;
	assign n_8097 = (~n_3480 & n_8096) ;
	assign n_3474 = (~n_3472 & ~n_3473) ;
	assign n_3452 = (~x_437 & n_3450) ;
	assign n_3451 = (x_437 & ~n_3450) ;
	assign n_3444 = (i_5 & ~n_3443) ;
	assign n_3432 = (i_66 & n_948) ;
	assign n_3431 = (x_439 & n_945) ;
	assign n_3425 = (i_30 & n_64) ;
	assign n_3373 = (~n_160 & ~n_161) ;
	assign n_8098 = (~n_3474 & n_8097) ;
	assign n_3453 = (~n_3451 & ~n_3452) ;
	assign n_3446 = (~x_438 & ~n_3444) ;
	assign n_3445 = (x_438 & n_3444) ;
	assign n_3433 = (~n_3431 & ~n_3432) ;
	assign n_3426 = (n_66 & n_3425) ;
	assign n_3424 = (x_440 & n_978) ;
	assign n_3418 = (~x_441 & ~n_936) ;
	assign n_3375 = (x_132 & n_3373) ;
	assign n_8099 = (~n_3453 & n_8098) ;
	assign n_3447 = (~n_3445 & ~n_3446) ;
	assign n_3435 = (~x_439 & n_3433) ;
	assign n_3434 = (x_439 & ~n_3433) ;
	assign n_3427 = (~n_3424 & ~n_3426) ;
	assign n_3419 = (i_5 & ~n_3418) ;
	assign n_3417 = (~i_29 & n_936) ;
	assign n_3411 = (~x_442 & ~n_936) ;
	assign n_3376 = (~x_332 & ~n_3375) ;
	assign n_3374 = (~x_132 & ~n_3373) ;
	assign n_3354 = (~x_609 & n_786) ;
	assign n_3353 = (x_609 & ~n_786) ;
	assign n_8100 = (~n_3447 & n_8099) ;
	assign n_3436 = (~n_3434 & ~n_3435) ;
	assign n_3429 = (~x_440 & n_3427) ;
	assign n_3428 = (x_440 & ~n_3427) ;
	assign n_3420 = (~n_3417 & n_3419) ;
	assign n_3412 = (i_5 & ~n_3411) ;
	assign n_3410 = (~i_27 & n_936) ;
	assign n_3404 = (i_48 & n_59) ;
	assign n_3377 = (~n_3374 & n_3376) ;
	assign n_3355 = (~n_3353 & ~n_3354) ;
	assign n_3352 = (~n_776 & ~n_777) ;
	assign n_8101 = (~n_3436 & n_8100) ;
	assign n_3430 = (~n_3428 & ~n_3429) ;
	assign n_3422 = (~x_441 & ~n_3420) ;
	assign n_3421 = (x_441 & n_3420) ;
	assign n_3413 = (~n_3410 & n_3412) ;
	assign n_3405 = (n_66 & n_3404) ;
	assign n_3403 = (x_443 & n_60) ;
	assign n_3379 = (n_164 & ~n_3377) ;
	assign n_3364 = (~x_447 & n_6) ;
	assign n_3357 = (n_3352 & ~n_3355) ;
	assign n_8102 = (~n_3430 & n_8101) ;
	assign n_3423 = (~n_3421 & ~n_3422) ;
	assign n_3415 = (~x_442 & ~n_3413) ;
	assign n_3414 = (x_442 & n_3413) ;
	assign n_3406 = (~n_3403 & ~n_3405) ;
	assign n_3398 = (x_677 & n_53) ;
	assign n_3397 = (x_444 & n_51) ;
	assign n_3391 = (i_31 & n_64) ;
	assign n_3383 = (~n_164 & ~n_1606) ;
	assign n_3382 = (i_30 & n_7) ;
	assign n_3380 = (x_664 & ~n_3379) ;
	assign n_3378 = (~n_164 & n_3377) ;
	assign n_3365 = (~n_3363 & ~n_3364) ;
	assign n_3360 = (x_447 & ~n_697) ;
	assign n_3358 = (n_697 & ~n_3357) ;
	assign n_3356 = (~n_3352 & n_3355) ;
	assign n_8103 = (~n_3423 & n_8102) ;
	assign n_3416 = (~n_3414 & ~n_3415) ;
	assign n_3408 = (~x_443 & n_3406) ;
	assign n_3407 = (x_443 & ~n_3406) ;
	assign n_3399 = (~n_3397 & ~n_3398) ;
	assign n_3392 = (n_66 & n_3391) ;
	assign n_3390 = (x_445 & n_978) ;
	assign n_3384 = (~n_3382 & ~n_3383) ;
	assign n_3381 = (~n_3378 & n_3380) ;
	assign n_3366 = (n_629 & ~n_3365) ;
	assign n_3361 = (~n_629 & ~n_3360) ;
	assign n_3359 = (~n_3356 & n_3358) ;
	assign n_8104 = (~n_3416 & n_8103) ;
	assign n_3409 = (~n_3407 & ~n_3408) ;
	assign n_3401 = (~x_444 & n_3399) ;
	assign n_3400 = (x_444 & ~n_3399) ;
	assign n_3393 = (~n_3390 & ~n_3392) ;
	assign n_3385 = (~n_3381 & n_3384) ;
	assign n_3367 = (n_902 & ~n_3366) ;
	assign n_3362 = (~n_3359 & n_3361) ;
	assign n_8105 = (~n_3409 & n_8104) ;
	assign n_3402 = (~n_3400 & ~n_3401) ;
	assign n_3395 = (~x_445 & n_3393) ;
	assign n_3394 = (x_445 & ~n_3393) ;
	assign n_3386 = (i_5 & ~n_3385) ;
	assign n_3368 = (~n_3362 & n_3367) ;
	assign n_3351 = (x_447 & n_699) ;
	assign n_3345 = (~x_448 & ~n_544) ;
	assign n_8106 = (~n_3402 & n_8105) ;
	assign n_3396 = (~n_3394 & ~n_3395) ;
	assign n_3388 = (~x_446 & ~n_3386) ;
	assign n_3387 = (x_446 & n_3386) ;
	assign n_3369 = (~n_3351 & ~n_3368) ;
	assign n_3346 = (i_5 & ~n_3345) ;
	assign n_3344 = (~i_14 & n_544) ;
	assign n_3287 = (~n_223 & ~n_224) ;
	assign n_8107 = (~n_3396 & n_8106) ;
	assign n_3389 = (~n_3387 & ~n_3388) ;
	assign n_3371 = (~x_447 & n_3369) ;
	assign n_3370 = (x_447 & ~n_3369) ;
	assign n_3347 = (~n_3344 & n_3346) ;
	assign n_3339 = (i_20 & n_948) ;
	assign n_3338 = (x_449 & n_945) ;
	assign n_3332 = (~x_450 & ~n_630) ;
	assign n_3289 = (~x_515 & ~n_3287) ;
	assign n_8108 = (~n_3389 & n_8107) ;
	assign n_3372 = (~n_3370 & ~n_3371) ;
	assign n_3349 = (~x_448 & ~n_3347) ;
	assign n_3348 = (x_448 & n_3347) ;
	assign n_3340 = (~n_3338 & ~n_3339) ;
	assign n_3333 = (i_5 & ~n_3332) ;
	assign n_3331 = (~i_55 & n_630) ;
	assign n_3325 = (~x_451 & ~n_936) ;
	assign n_3290 = (~x_332 & ~n_3289) ;
	assign n_3288 = (x_515 & n_3287) ;
	assign n_8109 = (~n_3372 & n_8108) ;
	assign n_3350 = (~n_3348 & ~n_3349) ;
	assign n_3342 = (~x_449 & n_3340) ;
	assign n_3341 = (x_449 & ~n_3340) ;
	assign n_3334 = (~n_3331 & n_3333) ;
	assign n_3326 = (i_5 & ~n_3325) ;
	assign n_3324 = (~i_53 & n_936) ;
	assign n_3291 = (~n_3288 & n_3290) ;
	assign n_8110 = (~n_3350 & n_8109) ;
	assign n_3343 = (~n_3341 & ~n_3342) ;
	assign n_3336 = (~x_450 & ~n_3334) ;
	assign n_3335 = (x_450 & n_3334) ;
	assign n_3327 = (~n_3324 & n_3326) ;
	assign n_3319 = (x_307 & n_53) ;
	assign n_3318 = (x_452 & n_51) ;
	assign n_3312 = (i_21 & n_59) ;
	assign n_3293 = (n_227 & ~n_3291) ;
	assign n_3256 = (~x_550 & n_2850) ;
	assign n_3255 = (x_550 & ~n_2850) ;
	assign n_8111 = (~n_3343 & n_8110) ;
	assign n_3337 = (~n_3335 & ~n_3336) ;
	assign n_3329 = (~x_451 & ~n_3327) ;
	assign n_3328 = (x_451 & n_3327) ;
	assign n_3320 = (~n_3318 & ~n_3319) ;
	assign n_3313 = (n_66 & n_3312) ;
	assign n_3311 = (x_453 & n_60) ;
	assign n_3305 = (~x_454 & ~n_544) ;
	assign n_3297 = (~n_227 & ~n_1606) ;
	assign n_3296 = (i_32 & n_7) ;
	assign n_3294 = (x_664 & ~n_3293) ;
	assign n_3292 = (~n_227 & n_3291) ;
	assign n_3257 = (~n_3255 & ~n_3256) ;
	assign n_3254 = (~n_2840 & ~n_2841) ;
	assign n_8112 = (~n_3337 & n_8111) ;
	assign n_3330 = (~n_3328 & ~n_3329) ;
	assign n_3322 = (~x_452 & n_3320) ;
	assign n_3321 = (x_452 & ~n_3320) ;
	assign n_3314 = (~n_3311 & ~n_3313) ;
	assign n_3306 = (i_5 & ~n_3305) ;
	assign n_3304 = (~i_43 & n_544) ;
	assign n_3298 = (~n_3296 & ~n_3297) ;
	assign n_3295 = (~n_3292 & n_3294) ;
	assign n_3265 = (~x_458 & n_6) ;
	assign n_2753 = (~i_63 & ~n_6) ;
	assign n_3259 = (n_3254 & ~n_3257) ;
	assign n_8113 = (~n_3330 & n_8112) ;
	assign n_3323 = (~n_3321 & ~n_3322) ;
	assign n_3316 = (~x_453 & n_3314) ;
	assign n_3315 = (x_453 & ~n_3314) ;
	assign n_3307 = (~n_3304 & n_3306) ;
	assign n_3299 = (~n_3295 & n_3298) ;
	assign n_3281 = (~x_456 & ~n_544) ;
	assign n_3266 = (~n_2753 & ~n_3265) ;
	assign n_3262 = (x_458 & ~n_697) ;
	assign n_3260 = (n_697 & ~n_3259) ;
	assign n_3258 = (~n_3254 & n_3257) ;
	assign n_3214 = (~n_268 & ~n_269) ;
	assign n_8114 = (~n_3323 & n_8113) ;
	assign n_3317 = (~n_3315 & ~n_3316) ;
	assign n_3309 = (~x_454 & ~n_3307) ;
	assign n_3308 = (x_454 & n_3307) ;
	assign n_3300 = (i_5 & ~n_3299) ;
	assign n_3282 = (i_5 & ~n_3281) ;
	assign n_3280 = (~i_50 & n_544) ;
	assign n_3267 = (n_629 & ~n_3266) ;
	assign n_3263 = (~n_629 & ~n_3262) ;
	assign n_3261 = (~n_3258 & n_3260) ;
	assign n_3216 = (~x_583 & ~n_3214) ;
	assign n_8115 = (~n_3317 & n_8114) ;
	assign n_3310 = (~n_3308 & ~n_3309) ;
	assign n_3302 = (~x_455 & ~n_3300) ;
	assign n_3301 = (x_455 & n_3300) ;
	assign n_3283 = (~n_3280 & n_3282) ;
	assign n_3275 = (~n_317 & n_35) ;
	assign n_3274 = (x_457 & n_36) ;
	assign n_3268 = (n_902 & ~n_3267) ;
	assign n_3264 = (~n_3261 & n_3263) ;
	assign n_3217 = (~x_332 & ~n_3216) ;
	assign n_3215 = (x_583 & n_3214) ;
	assign n_8116 = (~n_3310 & n_8115) ;
	assign n_3303 = (~n_3301 & ~n_3302) ;
	assign n_3285 = (~x_456 & ~n_3283) ;
	assign n_3284 = (x_456 & n_3283) ;
	assign n_3276 = (~n_3274 & ~n_3275) ;
	assign n_3269 = (~n_3264 & n_3268) ;
	assign n_3253 = (x_458 & n_699) ;
	assign n_3247 = (~x_459 & ~n_630) ;
	assign n_3239 = (i_34 & n_7) ;
	assign n_3238 = (x_350 & ~n_16) ;
	assign n_3218 = (~n_3215 & n_3217) ;
	assign n_8117 = (~n_3303 & n_8116) ;
	assign n_3286 = (~n_3284 & ~n_3285) ;
	assign n_3278 = (~x_457 & n_3276) ;
	assign n_3277 = (x_457 & ~n_3276) ;
	assign n_3270 = (~n_3253 & ~n_3269) ;
	assign n_3248 = (i_5 & ~n_3247) ;
	assign n_3246 = (~i_9 & n_630) ;
	assign n_3240 = (~n_3238 & ~n_3239) ;
	assign n_3220 = (n_272 & ~n_3218) ;
	assign n_8118 = (~n_3286 & n_8117) ;
	assign n_3279 = (~n_3277 & ~n_3278) ;
	assign n_3272 = (~x_458 & n_3270) ;
	assign n_3271 = (x_458 & ~n_3270) ;
	assign n_3249 = (~n_3246 & n_3248) ;
	assign n_3241 = (n_20 & ~n_3240) ;
	assign n_3237 = (x_460 & n_18) ;
	assign n_3224 = (~n_272 & ~n_1606) ;
	assign n_3223 = (i_26 & n_7) ;
	assign n_3221 = (x_664 & ~n_3220) ;
	assign n_3219 = (~n_272 & n_3218) ;
	assign n_8119 = (~n_3279 & n_8118) ;
	assign n_3273 = (~n_3271 & ~n_3272) ;
	assign n_3251 = (~x_459 & ~n_3249) ;
	assign n_3250 = (x_459 & n_3249) ;
	assign n_3242 = (~n_3237 & ~n_3241) ;
	assign n_3232 = (i_67 & n_948) ;
	assign n_3231 = (x_461 & n_945) ;
	assign n_3225 = (~n_3223 & ~n_3224) ;
	assign n_3222 = (~n_3219 & n_3221) ;
	assign n_8120 = (~n_3273 & n_8119) ;
	assign n_3252 = (~n_3250 & ~n_3251) ;
	assign n_3244 = (~x_460 & n_3242) ;
	assign n_3243 = (x_460 & ~n_3242) ;
	assign n_3233 = (~n_3231 & ~n_3232) ;
	assign n_3226 = (~n_3222 & n_3225) ;
	assign n_3201 = (~i_52 & n_669) ;
	assign n_3199 = (~x_677 & ~n_544) ;
	assign n_8121 = (~n_3252 & n_8120) ;
	assign n_3245 = (~n_3243 & ~n_3244) ;
	assign n_3235 = (~x_461 & n_3233) ;
	assign n_3234 = (x_461 & ~n_3233) ;
	assign n_3227 = (i_5 & ~n_3226) ;
	assign n_3209 = (~n_86 & n_1009) ;
	assign n_3208 = (x_463 & n_1007) ;
	assign n_3202 = (i_5 & ~n_3201) ;
	assign n_3200 = (n_662 & n_3199) ;
	assign n_8122 = (~n_3245 & n_8121) ;
	assign n_3236 = (~n_3234 & ~n_3235) ;
	assign n_3229 = (~x_462 & ~n_3227) ;
	assign n_3228 = (x_462 & n_3227) ;
	assign n_3210 = (~n_3208 & ~n_3209) ;
	assign n_3203 = (~n_3200 & n_3202) ;
	assign n_3198 = (~x_464 & ~n_665) ;
	assign n_3192 = (~x_465 & ~n_697) ;
	assign n_8123 = (~n_3236 & n_8122) ;
	assign n_3230 = (~n_3228 & ~n_3229) ;
	assign n_3212 = (~x_463 & n_3210) ;
	assign n_3211 = (x_463 & ~n_3210) ;
	assign n_3204 = (~n_3198 & n_3203) ;
	assign n_3193 = (i_5 & ~n_3192) ;
	assign n_3191 = (~x_220 & n_697) ;
	assign n_3185 = (~x_466 & ~n_630) ;
	assign n_8124 = (~n_3230 & n_8123) ;
	assign n_3213 = (~n_3211 & ~n_3212) ;
	assign n_3206 = (~x_464 & ~n_3204) ;
	assign n_3205 = (x_464 & n_3204) ;
	assign n_3194 = (~n_3191 & n_3193) ;
	assign n_3186 = (i_5 & ~n_3185) ;
	assign n_3184 = (~i_34 & n_630) ;
	assign n_8125 = (~n_3213 & n_8124) ;
	assign n_3207 = (~n_3205 & ~n_3206) ;
	assign n_3196 = (~x_465 & ~n_3194) ;
	assign n_3195 = (x_465 & n_3194) ;
	assign n_3187 = (~n_3184 & n_3186) ;
	assign n_3179 = (x_188 & n_35) ;
	assign n_3178 = (x_467 & n_36) ;
	assign n_8126 = (~n_3207 & n_8125) ;
	assign n_3197 = (~n_3195 & ~n_3196) ;
	assign n_3189 = (~x_466 & ~n_3187) ;
	assign n_3188 = (x_466 & n_3187) ;
	assign n_3180 = (~n_3178 & ~n_3179) ;
	assign n_3173 = (n_35 & ~n_1223) ;
	assign n_3172 = (x_468 & n_36) ;
	assign n_3166 = (~x_469 & ~n_936) ;
	assign n_8127 = (~n_3197 & n_8126) ;
	assign n_3190 = (~n_3188 & ~n_3189) ;
	assign n_3182 = (~x_467 & n_3180) ;
	assign n_3181 = (x_467 & ~n_3180) ;
	assign n_3174 = (~n_3172 & ~n_3173) ;
	assign n_3167 = (i_5 & ~n_3166) ;
	assign n_3165 = (~i_50 & n_936) ;
	assign n_3159 = (i_14 & n_59) ;
	assign n_8128 = (~n_3190 & n_8127) ;
	assign n_3183 = (~n_3181 & ~n_3182) ;
	assign n_3176 = (~x_468 & n_3174) ;
	assign n_3175 = (x_468 & ~n_3174) ;
	assign n_3168 = (~n_3165 & n_3167) ;
	assign n_3160 = (n_66 & n_3159) ;
	assign n_3158 = (x_470 & n_60) ;
	assign n_8129 = (~n_3183 & n_8128) ;
	assign n_3177 = (~n_3175 & ~n_3176) ;
	assign n_3170 = (~x_469 & ~n_3168) ;
	assign n_3169 = (x_469 & n_3168) ;
	assign n_3161 = (~n_3158 & ~n_3160) ;
	assign n_3153 = (i_17 & n_948) ;
	assign n_3152 = (x_471 & n_945) ;
	assign n_3146 = (i_67 & n_64) ;
	assign n_8130 = (~n_3177 & n_8129) ;
	assign n_3171 = (~n_3169 & ~n_3170) ;
	assign n_3163 = (~x_470 & n_3161) ;
	assign n_3162 = (x_470 & ~n_3161) ;
	assign n_3154 = (~n_3152 & ~n_3153) ;
	assign n_3147 = (n_66 & n_3146) ;
	assign n_3145 = (x_472 & n_978) ;
	assign n_8131 = (~n_3171 & n_8130) ;
	assign n_3164 = (~n_3162 & ~n_3163) ;
	assign n_3156 = (~x_471 & n_3154) ;
	assign n_3155 = (x_471 & ~n_3154) ;
	assign n_3148 = (~n_3145 & ~n_3147) ;
	assign n_3140 = (x_407 & n_53) ;
	assign n_3139 = (x_473 & n_51) ;
	assign n_3133 = (~x_474 & ~n_630) ;
	assign n_8132 = (~n_3164 & n_8131) ;
	assign n_3157 = (~n_3155 & ~n_3156) ;
	assign n_3150 = (~x_472 & n_3148) ;
	assign n_3149 = (x_472 & ~n_3148) ;
	assign n_3141 = (~n_3139 & ~n_3140) ;
	assign n_3134 = (i_5 & ~n_3133) ;
	assign n_3132 = (~i_46 & n_630) ;
	assign n_8133 = (~n_3157 & n_8132) ;
	assign n_3151 = (~n_3149 & ~n_3150) ;
	assign n_3143 = (~x_473 & n_3141) ;
	assign n_3142 = (x_473 & ~n_3141) ;
	assign n_3135 = (~n_3132 & n_3134) ;
	assign n_3127 = (x_328 & n_35) ;
	assign n_3126 = (x_475 & n_36) ;
	assign n_3120 = (~x_476 & ~n_936) ;
	assign n_8134 = (~n_3151 & n_8133) ;
	assign n_3144 = (~n_3142 & ~n_3143) ;
	assign n_3137 = (~x_474 & ~n_3135) ;
	assign n_3136 = (x_474 & n_3135) ;
	assign n_3128 = (~n_3126 & ~n_3127) ;
	assign n_3121 = (i_5 & ~n_3120) ;
	assign n_3119 = (~i_43 & n_936) ;
	assign n_3113 = (~x_477 & ~n_697) ;
	assign n_8135 = (~n_3144 & n_8134) ;
	assign n_3138 = (~n_3136 & ~n_3137) ;
	assign n_3130 = (~x_475 & n_3128) ;
	assign n_3129 = (x_475 & ~n_3128) ;
	assign n_3122 = (~n_3119 & n_3121) ;
	assign n_3114 = (i_5 & ~n_3113) ;
	assign n_3112 = (~x_738 & n_697) ;
	assign n_3106 = (i_54 & n_59) ;
	assign n_3082 = (i_47 & ~n_6) ;
	assign n_8136 = (~n_3138 & n_8135) ;
	assign n_3131 = (~n_3129 & ~n_3130) ;
	assign n_3124 = (~x_476 & ~n_3122) ;
	assign n_3123 = (x_476 & n_3122) ;
	assign n_3115 = (~n_3112 & n_3114) ;
	assign n_3107 = (n_66 & n_3106) ;
	assign n_3105 = (x_478 & n_60) ;
	assign n_3099 = (i_20 & n_64) ;
	assign n_3083 = (n_629 & ~n_3082) ;
	assign n_3081 = (x_481 & n_6) ;
	assign n_8137 = (~n_3131 & n_8136) ;
	assign n_3125 = (~n_3123 & ~n_3124) ;
	assign n_3117 = (~x_477 & ~n_3115) ;
	assign n_3116 = (x_477 & n_3115) ;
	assign n_3108 = (~n_3105 & ~n_3107) ;
	assign n_3100 = (n_66 & n_3099) ;
	assign n_3098 = (x_479 & n_978) ;
	assign n_3092 = (~x_480 & ~n_936) ;
	assign n_3084 = (~n_3081 & n_3083) ;
	assign n_8138 = (~n_3125 & n_8137) ;
	assign n_3118 = (~n_3116 & ~n_3117) ;
	assign n_3110 = (~x_478 & n_3108) ;
	assign n_3109 = (x_478 & ~n_3108) ;
	assign n_3101 = (~n_3098 & ~n_3100) ;
	assign n_3093 = (i_5 & ~n_3092) ;
	assign n_3091 = (~i_59 & n_936) ;
	assign n_3085 = (i_5 & ~n_3084) ;
	assign n_3080 = (~x_773 & n_662) ;
	assign n_8139 = (~n_3118 & n_8138) ;
	assign n_3111 = (~n_3109 & ~n_3110) ;
	assign n_3103 = (~x_479 & n_3101) ;
	assign n_3102 = (x_479 & ~n_3101) ;
	assign n_3094 = (~n_3091 & n_3093) ;
	assign n_3086 = (~n_3080 & n_3085) ;
	assign n_3079 = (~x_481 & n_663) ;
	assign n_3073 = (~x_482 & ~n_544) ;
	assign n_8140 = (~n_3111 & n_8139) ;
	assign n_3104 = (~n_3102 & ~n_3103) ;
	assign n_3096 = (~x_480 & ~n_3094) ;
	assign n_3095 = (x_480 & n_3094) ;
	assign n_3087 = (~n_3079 & n_3086) ;
	assign n_3074 = (i_5 & ~n_3073) ;
	assign n_3072 = (~i_45 & n_544) ;
	assign n_3066 = (~x_483 & ~n_630) ;
	assign n_8141 = (~n_3104 & n_8140) ;
	assign n_3097 = (~n_3095 & ~n_3096) ;
	assign n_3089 = (~x_481 & ~n_3087) ;
	assign n_3088 = (x_481 & n_3087) ;
	assign n_3075 = (~n_3072 & n_3074) ;
	assign n_3067 = (i_5 & ~n_3066) ;
	assign n_3065 = (~i_64 & n_630) ;
	assign n_8142 = (~n_3097 & n_8141) ;
	assign n_3090 = (~n_3088 & ~n_3089) ;
	assign n_3077 = (~x_482 & ~n_3075) ;
	assign n_3076 = (x_482 & n_3075) ;
	assign n_3068 = (~n_3065 & n_3067) ;
	assign n_3060 = (~n_164 & n_35) ;
	assign n_3059 = (x_484 & n_36) ;
	assign n_8143 = (~n_3090 & n_8142) ;
	assign n_3078 = (~n_3076 & ~n_3077) ;
	assign n_3070 = (~x_483 & ~n_3068) ;
	assign n_3069 = (x_483 & n_3068) ;
	assign n_3061 = (~n_3059 & ~n_3060) ;
	assign n_3054 = (~n_179 & n_1009) ;
	assign n_3053 = (x_485 & n_1007) ;
	assign n_3047 = (~x_486 & ~n_936) ;
	assign n_8144 = (~n_3078 & n_8143) ;
	assign n_3071 = (~n_3069 & ~n_3070) ;
	assign n_3063 = (~x_484 & n_3061) ;
	assign n_3062 = (x_484 & ~n_3061) ;
	assign n_3055 = (~n_3053 & ~n_3054) ;
	assign n_3048 = (i_5 & ~n_3047) ;
	assign n_3046 = (~i_26 & n_936) ;
	assign n_8145 = (~n_3071 & n_8144) ;
	assign n_3064 = (~n_3062 & ~n_3063) ;
	assign n_3057 = (~x_485 & n_3055) ;
	assign n_3056 = (x_485 & ~n_3055) ;
	assign n_3049 = (~n_3046 & n_3048) ;
	assign n_3041 = (i_62 & n_948) ;
	assign n_3040 = (x_487 & n_945) ;
	assign n_2987 = (~x_383 & n_721) ;
	assign n_2986 = (x_383 & ~n_721) ;
	assign n_8146 = (~n_3064 & n_8145) ;
	assign n_3058 = (~n_3056 & ~n_3057) ;
	assign n_3051 = (~x_486 & ~n_3049) ;
	assign n_3050 = (x_486 & n_3049) ;
	assign n_3042 = (~n_3040 & ~n_3041) ;
	assign n_3035 = (x_418 & n_35) ;
	assign n_3034 = (x_488 & n_36) ;
	assign n_3028 = (i_46 & n_64) ;
	assign n_2988 = (~n_2986 & ~n_2987) ;
	assign n_2985 = (~n_711 & ~n_712) ;
	assign n_8147 = (~n_3058 & n_8146) ;
	assign n_3052 = (~n_3050 & ~n_3051) ;
	assign n_3044 = (~x_487 & n_3042) ;
	assign n_3043 = (x_487 & ~n_3042) ;
	assign n_3036 = (~n_3034 & ~n_3035) ;
	assign n_3029 = (n_66 & n_3028) ;
	assign n_3027 = (x_489 & n_978) ;
	assign n_3021 = (i_35 & n_59) ;
	assign n_2997 = (i_11 & ~n_6) ;
	assign n_2990 = (n_2985 & ~n_2988) ;
	assign n_8148 = (~n_3052 & n_8147) ;
	assign n_3045 = (~n_3043 & ~n_3044) ;
	assign n_3038 = (~x_488 & n_3036) ;
	assign n_3037 = (x_488 & ~n_3036) ;
	assign n_3030 = (~n_3027 & ~n_3029) ;
	assign n_3022 = (n_66 & n_3021) ;
	assign n_3020 = (x_490 & n_60) ;
	assign n_3014 = (~x_491 & ~n_936) ;
	assign n_2998 = (n_629 & ~n_2997) ;
	assign n_2996 = (x_493 & n_6) ;
	assign n_2993 = (x_493 & ~n_697) ;
	assign n_2991 = (n_697 & ~n_2990) ;
	assign n_2989 = (~n_2985 & n_2988) ;
	assign n_8149 = (~n_3045 & n_8148) ;
	assign n_3039 = (~n_3037 & ~n_3038) ;
	assign n_3032 = (~x_489 & n_3030) ;
	assign n_3031 = (x_489 & ~n_3030) ;
	assign n_3023 = (~n_3020 & ~n_3022) ;
	assign n_3015 = (i_5 & ~n_3014) ;
	assign n_3013 = (~i_6 & n_936) ;
	assign n_3007 = (~x_492 & ~n_544) ;
	assign n_2999 = (~n_2996 & n_2998) ;
	assign n_2994 = (~n_629 & ~n_2993) ;
	assign n_2992 = (~n_2989 & n_2991) ;
	assign n_8150 = (~n_3039 & n_8149) ;
	assign n_3033 = (~n_3031 & ~n_3032) ;
	assign n_3025 = (~x_490 & n_3023) ;
	assign n_3024 = (x_490 & ~n_3023) ;
	assign n_3016 = (~n_3013 & n_3015) ;
	assign n_3008 = (i_5 & ~n_3007) ;
	assign n_3006 = (~i_4 & n_544) ;
	assign n_3000 = (n_902 & ~n_2999) ;
	assign n_2995 = (~n_2992 & n_2994) ;
	assign n_8151 = (~n_3033 & n_8150) ;
	assign n_3026 = (~n_3024 & ~n_3025) ;
	assign n_3018 = (~x_491 & ~n_3016) ;
	assign n_3017 = (x_491 & n_3016) ;
	assign n_3009 = (~n_3006 & n_3008) ;
	assign n_3001 = (~n_2995 & n_3000) ;
	assign n_2984 = (x_493 & n_699) ;
	assign n_8152 = (~n_3026 & n_8151) ;
	assign n_3019 = (~n_3017 & ~n_3018) ;
	assign n_3011 = (~x_492 & ~n_3009) ;
	assign n_3010 = (x_492 & n_3009) ;
	assign n_3002 = (~n_2984 & ~n_3001) ;
	assign n_2979 = (x_270 & n_53) ;
	assign n_2978 = (x_494 & n_51) ;
	assign n_8153 = (~n_3019 & n_8152) ;
	assign n_3012 = (~n_3010 & ~n_3011) ;
	assign n_3004 = (~x_493 & n_3002) ;
	assign n_3003 = (x_493 & ~n_3002) ;
	assign n_2980 = (~n_2978 & ~n_2979) ;
	assign n_2973 = (x_576 & n_53) ;
	assign n_2972 = (x_495 & n_51) ;
	assign n_2966 = (i_9 & n_64) ;
	assign n_2950 = (~x_498 & ~n_662) ;
	assign n_2948 = (~x_622 & ~n_544) ;
	assign n_2945 = (~i_50 & ~n_6) ;
	assign n_8154 = (~n_3012 & n_8153) ;
	assign n_3005 = (~n_3003 & ~n_3004) ;
	assign n_2982 = (~x_494 & n_2980) ;
	assign n_2981 = (x_494 & ~n_2980) ;
	assign n_2974 = (~n_2972 & ~n_2973) ;
	assign n_2967 = (n_66 & n_2966) ;
	assign n_2965 = (x_496 & n_978) ;
	assign n_2959 = (~x_497 & ~n_630) ;
	assign n_2951 = (~n_629 & ~n_2950) ;
	assign n_2949 = (n_662 & n_2948) ;
	assign n_2946 = (n_629 & ~n_2945) ;
	assign n_2944 = (~x_498 & n_6) ;
	assign n_8155 = (~n_3005 & n_8154) ;
	assign n_2983 = (~n_2981 & ~n_2982) ;
	assign n_2976 = (~x_495 & n_2974) ;
	assign n_2975 = (x_495 & ~n_2974) ;
	assign n_2968 = (~n_2965 & ~n_2967) ;
	assign n_2960 = (i_5 & ~n_2959) ;
	assign n_2958 = (~i_20 & n_630) ;
	assign n_2952 = (~n_2949 & n_2951) ;
	assign n_2947 = (~n_2944 & n_2946) ;
	assign n_8156 = (~n_2983 & n_8155) ;
	assign n_2977 = (~n_2975 & ~n_2976) ;
	assign n_2970 = (~x_496 & n_2968) ;
	assign n_2969 = (x_496 & ~n_2968) ;
	assign n_2961 = (~n_2958 & n_2960) ;
	assign n_2953 = (~n_2947 & ~n_2952) ;
	assign n_2938 = (~x_499 & ~n_630) ;
	assign n_2892 = (~x_107 & n_2890) ;
	assign n_2891 = (x_107 & ~n_2890) ;
	assign n_8157 = (~n_2977 & n_8156) ;
	assign n_2971 = (~n_2969 & ~n_2970) ;
	assign n_2963 = (~x_497 & ~n_2961) ;
	assign n_2962 = (x_497 & n_2961) ;
	assign n_2954 = (i_5 & ~n_2953) ;
	assign n_2939 = (i_5 & ~n_2938) ;
	assign n_2937 = (~i_68 & n_630) ;
	assign n_2893 = (~n_2891 & ~n_2892) ;
	assign n_2881 = (~n_2879 & ~n_2880) ;
	assign n_8158 = (~n_2971 & n_8157) ;
	assign n_2964 = (~n_2962 & ~n_2963) ;
	assign n_2956 = (~x_498 & ~n_2954) ;
	assign n_2955 = (x_498 & n_2954) ;
	assign n_2940 = (~n_2937 & n_2939) ;
	assign n_2932 = (x_341 & n_35) ;
	assign n_2931 = (x_500 & n_36) ;
	assign n_2902 = (~x_504 & n_6) ;
	assign n_2895 = (n_2881 & ~n_2893) ;
	assign n_8159 = (~n_2964 & n_8158) ;
	assign n_2957 = (~n_2955 & ~n_2956) ;
	assign n_2942 = (~x_499 & ~n_2940) ;
	assign n_2941 = (x_499 & n_2940) ;
	assign n_2933 = (~n_2931 & ~n_2932) ;
	assign n_2926 = (x_190 & n_53) ;
	assign n_2925 = (x_501 & n_51) ;
	assign n_2919 = (~x_502 & ~n_936) ;
	assign n_2903 = (~n_2901 & ~n_2902) ;
	assign n_2898 = (x_504 & ~n_697) ;
	assign n_2896 = (n_697 & ~n_2895) ;
	assign n_2894 = (~n_2881 & n_2893) ;
	assign n_8160 = (~n_2957 & n_8159) ;
	assign n_2943 = (~n_2941 & ~n_2942) ;
	assign n_2935 = (~x_500 & n_2933) ;
	assign n_2934 = (x_500 & ~n_2933) ;
	assign n_2927 = (~n_2925 & ~n_2926) ;
	assign n_2920 = (i_5 & ~n_2919) ;
	assign n_2918 = (~i_44 & n_936) ;
	assign n_2912 = (~x_503 & ~n_630) ;
	assign n_2904 = (n_629 & ~n_2903) ;
	assign n_2899 = (~n_629 & ~n_2898) ;
	assign n_2897 = (~n_2894 & n_2896) ;
	assign n_8161 = (~n_2943 & n_8160) ;
	assign n_2936 = (~n_2934 & ~n_2935) ;
	assign n_2929 = (~x_501 & n_2927) ;
	assign n_2928 = (x_501 & ~n_2927) ;
	assign n_2921 = (~n_2918 & n_2920) ;
	assign n_2913 = (i_5 & ~n_2912) ;
	assign n_2911 = (~i_31 & n_630) ;
	assign n_2905 = (n_902 & ~n_2904) ;
	assign n_2900 = (~n_2897 & n_2899) ;
	assign n_8162 = (~n_2936 & n_8161) ;
	assign n_2930 = (~n_2928 & ~n_2929) ;
	assign n_2923 = (~x_502 & ~n_2921) ;
	assign n_2922 = (x_502 & n_2921) ;
	assign n_2914 = (~n_2911 & n_2913) ;
	assign n_2906 = (~n_2900 & n_2905) ;
	assign n_2798 = (x_504 & n_699) ;
	assign n_2744 = (~n_448 & ~n_449) ;
	assign n_2724 = (~n_175 & ~n_176) ;
	assign n_8163 = (~n_2930 & n_8162) ;
	assign n_2924 = (~n_2922 & ~n_2923) ;
	assign n_2916 = (~x_503 & ~n_2914) ;
	assign n_2915 = (x_503 & n_2914) ;
	assign n_2907 = (~n_2798 & ~n_2906) ;
	assign n_2793 = (i_29 & n_948) ;
	assign n_2792 = (x_505 & n_945) ;
	assign n_2786 = (i_53 & n_64) ;
	assign n_2771 = (i_67 & n_1) ;
	assign n_2770 = (~x_508 & n_6) ;
	assign n_2746 = (~x_604 & ~n_2744) ;
	assign n_2726 = (~x_678 & ~n_2724) ;
	assign n_8164 = (~n_2924 & n_8163) ;
	assign n_2917 = (~n_2915 & ~n_2916) ;
	assign n_2909 = (~x_504 & n_2907) ;
	assign n_2908 = (x_504 & ~n_2907) ;
	assign n_2794 = (~n_2792 & ~n_2793) ;
	assign n_2787 = (n_66 & n_2786) ;
	assign n_2785 = (x_506 & n_978) ;
	assign n_2772 = (~n_2770 & n_2771) ;
	assign n_2769 = (x_389 & ~n_16) ;
	assign n_2747 = (n_527 & ~n_2746) ;
	assign n_2745 = (x_604 & n_2744) ;
	assign n_2727 = (~x_332 & ~n_2726) ;
	assign n_2725 = (x_678 & n_2724) ;
	assign n_8165 = (~n_2917 & n_8164) ;
	assign n_2910 = (~n_2908 & ~n_2909) ;
	assign n_2796 = (~x_505 & n_2794) ;
	assign n_2795 = (x_505 & ~n_2794) ;
	assign n_2788 = (~n_2785 & ~n_2787) ;
	assign n_2780 = (x_166 & n_53) ;
	assign n_2779 = (x_507 & n_51) ;
	assign n_2773 = (~n_2769 & ~n_2772) ;
	assign n_2768 = (x_508 & n_17) ;
	assign n_2754 = (n_6 & n_452) ;
	assign n_2748 = (~n_2745 & n_2747) ;
	assign n_2728 = (~n_2725 & n_2727) ;
	assign n_8166 = (~n_2910 & n_8165) ;
	assign n_2797 = (~n_2795 & ~n_2796) ;
	assign n_2790 = (~x_506 & n_2788) ;
	assign n_2789 = (x_506 & ~n_2788) ;
	assign n_2781 = (~n_2779 & ~n_2780) ;
	assign n_2774 = (~n_2768 & n_2773) ;
	assign n_2755 = (~n_2753 & ~n_2754) ;
	assign n_2750 = (n_452 & n_2748) ;
	assign n_2736 = (n_1 & ~n_2735) ;
	assign n_2734 = (n_6 & n_179) ;
	assign n_2730 = (n_179 & ~n_2728) ;
	assign n_8167 = (~n_2797 & n_8166) ;
	assign n_2791 = (~n_2789 & ~n_2790) ;
	assign n_2783 = (~x_507 & n_2781) ;
	assign n_2782 = (x_507 & ~n_2781) ;
	assign n_2775 = (i_5 & ~n_2774) ;
	assign n_2763 = (i_34 & n_948) ;
	assign n_2762 = (x_509 & n_945) ;
	assign n_2756 = (n_1 & ~n_2755) ;
	assign n_2751 = (~n_1 & ~n_2750) ;
	assign n_2749 = (~n_452 & ~n_2748) ;
	assign n_2737 = (~n_2734 & n_2736) ;
	assign n_2733 = (n_59 & ~n_179) ;
	assign n_2731 = (x_664 & ~n_2730) ;
	assign n_2729 = (~n_179 & n_2728) ;
	assign n_8168 = (~n_2791 & n_8167) ;
	assign n_2784 = (~n_2782 & ~n_2783) ;
	assign n_2777 = (~x_508 & ~n_2775) ;
	assign n_2776 = (x_508 & n_2775) ;
	assign n_2764 = (~n_2762 & ~n_2763) ;
	assign n_2757 = (i_5 & ~n_2756) ;
	assign n_2752 = (~n_2749 & n_2751) ;
	assign n_2738 = (~n_2733 & ~n_2737) ;
	assign n_2732 = (~n_2729 & n_2731) ;
	assign n_8169 = (~n_2784 & n_8168) ;
	assign n_2778 = (~n_2776 & ~n_2777) ;
	assign n_2766 = (~x_509 & n_2764) ;
	assign n_2765 = (x_509 & ~n_2764) ;
	assign n_2758 = (~n_2752 & n_2757) ;
	assign n_2739 = (~n_2732 & n_2738) ;
	assign n_2718 = (i_55 & n_64) ;
	assign n_2669 = (~x_410 & n_2667) ;
	assign n_2668 = (x_410 & ~n_2667) ;
	assign n_8170 = (~n_2778 & n_8169) ;
	assign n_2767 = (~n_2765 & ~n_2766) ;
	assign n_2760 = (~x_510 & ~n_2758) ;
	assign n_2759 = (x_510 & n_2758) ;
	assign n_2740 = (i_5 & ~n_2739) ;
	assign n_2719 = (n_66 & n_2718) ;
	assign n_2717 = (x_512 & n_978) ;
	assign n_2670 = (~n_2668 & ~n_2669) ;
	assign n_2658 = (~n_2656 & ~n_2657) ;
	assign n_8171 = (~n_2767 & n_8170) ;
	assign n_2761 = (~n_2759 & ~n_2760) ;
	assign n_2742 = (~x_511 & ~n_2740) ;
	assign n_2741 = (x_511 & n_2740) ;
	assign n_2720 = (~n_2717 & ~n_2719) ;
	assign n_2712 = (i_10 & n_948) ;
	assign n_2711 = (x_513 & n_945) ;
	assign n_2705 = (~x_514 & ~n_544) ;
	assign n_2697 = (i_16 & n_7) ;
	assign n_2696 = (x_272 & ~n_16) ;
	assign n_2679 = (i_4 & ~n_6) ;
	assign n_2672 = (n_2658 & ~n_2670) ;
	assign n_8172 = (~n_2761 & n_8171) ;
	assign n_2743 = (~n_2741 & ~n_2742) ;
	assign n_2722 = (~x_512 & n_2720) ;
	assign n_2721 = (x_512 & ~n_2720) ;
	assign n_2713 = (~n_2711 & ~n_2712) ;
	assign n_2706 = (i_5 & ~n_2705) ;
	assign n_2704 = (~i_24 & n_544) ;
	assign n_2698 = (~n_2696 & ~n_2697) ;
	assign n_2680 = (n_629 & ~n_2679) ;
	assign n_2678 = (x_600 & n_6) ;
	assign n_2675 = (x_600 & ~n_697) ;
	assign n_2673 = (n_697 & ~n_2672) ;
	assign n_2671 = (~n_2658 & n_2670) ;
	assign n_8173 = (~n_2743 & n_8172) ;
	assign n_2723 = (~n_2721 & ~n_2722) ;
	assign n_2715 = (~x_513 & n_2713) ;
	assign n_2714 = (x_513 & ~n_2713) ;
	assign n_2707 = (~n_2704 & n_2706) ;
	assign n_2699 = (n_20 & ~n_2698) ;
	assign n_2695 = (x_515 & n_18) ;
	assign n_2689 = (i_37 & n_59) ;
	assign n_2681 = (~n_2678 & n_2680) ;
	assign n_2676 = (~n_629 & ~n_2675) ;
	assign n_2674 = (~n_2671 & n_2673) ;
	assign n_8174 = (~n_2723 & n_8173) ;
	assign n_2716 = (~n_2714 & ~n_2715) ;
	assign n_2709 = (~x_514 & ~n_2707) ;
	assign n_2708 = (x_514 & n_2707) ;
	assign n_2700 = (~n_2695 & ~n_2699) ;
	assign n_2690 = (n_66 & n_2689) ;
	assign n_2688 = (x_599 & n_60) ;
	assign n_2682 = (n_902 & ~n_2681) ;
	assign n_2677 = (~n_2674 & n_2676) ;
	assign n_8175 = (~n_2716 & n_8174) ;
	assign n_2710 = (~n_2708 & ~n_2709) ;
	assign n_2702 = (~x_515 & n_2700) ;
	assign n_2701 = (x_515 & ~n_2700) ;
	assign n_2691 = (~n_2688 & ~n_2690) ;
	assign n_2683 = (~n_2677 & n_2682) ;
	assign n_2653 = (x_600 & n_699) ;
	assign n_2647 = (~x_601 & ~n_544) ;
	assign n_8176 = (~n_2710 & n_8175) ;
	assign n_2703 = (~n_2701 & ~n_2702) ;
	assign n_2693 = (~x_599 & n_2691) ;
	assign n_2692 = (x_599 & ~n_2691) ;
	assign n_2684 = (~n_2653 & ~n_2683) ;
	assign n_2648 = (i_5 & ~n_2647) ;
	assign n_2646 = (~i_40 & n_544) ;
	assign n_8177 = (~n_2703 & n_8176) ;
	assign n_2694 = (~n_2692 & ~n_2693) ;
	assign n_2686 = (~x_600 & n_2684) ;
	assign n_2685 = (x_600 & ~n_2684) ;
	assign n_2649 = (~n_2646 & n_2648) ;
	assign n_2641 = (x_323 & n_53) ;
	assign n_2640 = (x_602 & n_51) ;
	assign n_2634 = (~x_603 & ~n_544) ;
	assign n_2626 = (i_28 & n_7) ;
	assign n_2625 = (x_254 & ~n_16) ;
	assign n_8178 = (~n_2694 & n_8177) ;
	assign n_2687 = (~n_2685 & ~n_2686) ;
	assign n_2651 = (~x_601 & ~n_2649) ;
	assign n_2650 = (x_601 & n_2649) ;
	assign n_2642 = (~n_2640 & ~n_2641) ;
	assign n_2635 = (i_5 & ~n_2634) ;
	assign n_2633 = (~i_56 & n_544) ;
	assign n_2627 = (~n_2625 & ~n_2626) ;
	assign n_8179 = (~n_2687 & n_8178) ;
	assign n_2652 = (~n_2650 & ~n_2651) ;
	assign n_2644 = (~x_602 & n_2642) ;
	assign n_2643 = (x_602 & ~n_2642) ;
	assign n_2636 = (~n_2633 & n_2635) ;
	assign n_2628 = (n_20 & ~n_2627) ;
	assign n_2624 = (x_604 & n_18) ;
	assign n_2618 = (~x_605 & ~n_936) ;
	assign n_8180 = (~n_2652 & n_8179) ;
	assign n_2645 = (~n_2643 & ~n_2644) ;
	assign n_2638 = (~x_603 & ~n_2636) ;
	assign n_2637 = (x_603 & n_2636) ;
	assign n_2629 = (~n_2624 & ~n_2628) ;
	assign n_2619 = (i_5 & ~n_2618) ;
	assign n_2617 = (~i_54 & n_936) ;
	assign n_2611 = (~x_606 & ~n_544) ;
	assign n_2588 = (i_44 & ~n_6) ;
	assign n_8181 = (~n_2645 & n_8180) ;
	assign n_2639 = (~n_2637 & ~n_2638) ;
	assign n_2631 = (~x_604 & n_2629) ;
	assign n_2630 = (x_604 & ~n_2629) ;
	assign n_2620 = (~n_2617 & n_2619) ;
	assign n_2612 = (i_5 & ~n_2611) ;
	assign n_2610 = (~i_36 & n_544) ;
	assign n_2589 = (n_629 & ~n_2588) ;
	assign n_2587 = (x_609 & n_6) ;
	assign n_8182 = (~n_2639 & n_8181) ;
	assign n_2632 = (~n_2630 & ~n_2631) ;
	assign n_2622 = (~x_605 & ~n_2620) ;
	assign n_2621 = (x_605 & n_2620) ;
	assign n_2613 = (~n_2610 & n_2612) ;
	assign n_2605 = (i_55 & n_948) ;
	assign n_2604 = (x_607 & n_945) ;
	assign n_2598 = (i_27 & n_59) ;
	assign n_2590 = (~n_2587 & n_2589) ;
	assign n_8183 = (~n_2632 & n_8182) ;
	assign n_2623 = (~n_2621 & ~n_2622) ;
	assign n_2615 = (~x_606 & ~n_2613) ;
	assign n_2614 = (x_606 & n_2613) ;
	assign n_2606 = (~n_2604 & ~n_2605) ;
	assign n_2599 = (n_66 & n_2598) ;
	assign n_2597 = (x_608 & n_60) ;
	assign n_2591 = (i_5 & ~n_2590) ;
	assign n_2586 = (~x_526 & n_662) ;
	assign n_8184 = (~n_2623 & n_8183) ;
	assign n_2616 = (~n_2614 & ~n_2615) ;
	assign n_2608 = (~x_607 & n_2606) ;
	assign n_2607 = (x_607 & ~n_2606) ;
	assign n_2600 = (~n_2597 & ~n_2599) ;
	assign n_2592 = (~n_2586 & n_2591) ;
	assign n_2585 = (~x_609 & n_663) ;
	assign n_2579 = (~x_610 & ~n_697) ;
	assign n_623 = (~i_47 & ~i_48) ;
	assign n_622 = (~i_45 & ~i_46) ;
	assign n_620 = (~i_51 & ~i_52) ;
	assign n_619 = (~i_49 & ~i_50) ;
	assign n_616 = (~i_39 & ~i_40) ;
	assign n_615 = (~i_37 & ~i_38) ;
	assign n_613 = (~i_43 & ~i_44) ;
	assign n_612 = (~i_41 & ~i_42) ;
	assign n_608 = (~i_63 & ~i_64) ;
	assign n_607 = (~i_61 & ~i_62) ;
	assign n_605 = (~i_67 & ~i_68) ;
	assign n_604 = (~i_65 & ~i_66) ;
	assign n_601 = (~i_55 & ~i_56) ;
	assign n_600 = (~i_53 & ~i_54) ;
	assign n_598 = (~i_59 & ~i_60) ;
	assign n_597 = (~i_57 & ~i_58) ;
	assign n_592 = (~i_15 & ~i_16) ;
	assign n_591 = (~i_13 & ~i_14) ;
	assign n_589 = (~i_19 & ~i_20) ;
	assign n_588 = (~i_17 & ~i_18) ;
	assign n_585 = (~i_7 & ~i_8) ;
	assign n_584 = (~i_4 & ~i_6) ;
	assign n_582 = (~i_11 & ~i_12) ;
	assign n_581 = (~i_9 & ~i_10) ;
	assign n_577 = (~i_31 & ~i_32) ;
	assign n_576 = (~i_29 & ~i_30) ;
	assign n_574 = (~i_35 & ~i_36) ;
	assign n_573 = (~i_33 & ~i_34) ;
	assign n_570 = (~i_23 & ~i_24) ;
	assign n_569 = (~i_21 & ~i_22) ;
	assign n_567 = (~i_27 & ~i_28) ;
	assign n_566 = (~i_25 & ~i_26) ;
	assign n_2529 = (~x_431 & ~x_441) ;
	assign n_2528 = (~x_397 & ~x_420) ;
	assign n_2526 = (~x_469 & ~x_476) ;
	assign n_2525 = (~x_442 & ~x_451) ;
	assign n_2522 = (~x_339 & ~x_354) ;
	assign n_2521 = (~x_324 & ~x_330) ;
	assign n_2519 = (~x_379 & ~x_387) ;
	assign n_2518 = (~x_361 & ~x_371) ;
	assign n_2514 = (~x_585 & ~x_588) ;
	assign n_2513 = (~x_574 & ~x_580) ;
	assign n_2511 = (~x_623 & ~x_630) ;
	assign n_2510 = (~x_605 & ~x_617) ;
	assign n_2507 = (~x_491 & ~x_502) ;
	assign n_2506 = (~x_480 & ~x_486) ;
	assign n_2504 = (~x_560 & ~x_562) ;
	assign n_2503 = (~x_519 & ~x_523) ;
	assign n_8185 = (~n_2616 & n_8184) ;
	assign n_2609 = (~n_2607 & ~n_2608) ;
	assign n_2602 = (~x_608 & n_2600) ;
	assign n_2601 = (x_608 & ~n_2600) ;
	assign n_2593 = (~n_2585 & n_2592) ;
	assign n_2580 = (i_5 & ~n_2579) ;
	assign n_2578 = (~x_359 & n_697) ;
	assign n_2565 = (i_29 & n_7) ;
	assign n_2564 = (x_181 & ~n_16) ;
	assign n_624 = (n_622 & n_623) ;
	assign n_621 = (n_619 & n_620) ;
	assign n_617 = (n_615 & n_616) ;
	assign n_614 = (n_612 & n_613) ;
	assign n_609 = (n_607 & n_608) ;
	assign n_606 = (n_604 & n_605) ;
	assign n_602 = (n_600 & n_601) ;
	assign n_599 = (n_597 & n_598) ;
	assign n_593 = (n_591 & n_592) ;
	assign n_590 = (n_588 & n_589) ;
	assign n_586 = (n_584 & n_585) ;
	assign n_583 = (n_581 & n_582) ;
	assign n_578 = (n_576 & n_577) ;
	assign n_575 = (n_573 & n_574) ;
	assign n_571 = (n_569 & n_570) ;
	assign n_568 = (n_566 & n_567) ;
	assign n_2530 = (n_2528 & n_2529) ;
	assign n_2527 = (n_2525 & n_2526) ;
	assign n_2523 = (n_2521 & n_2522) ;
	assign n_2520 = (n_2518 & n_2519) ;
	assign n_2515 = (n_2513 & n_2514) ;
	assign n_2512 = (n_2510 & n_2511) ;
	assign n_2508 = (n_2506 & n_2507) ;
	assign n_2505 = (n_2503 & n_2504) ;
	assign n_2499 = (~x_666 & ~x_704) ;
	assign n_2498 = (~x_640 & ~x_643) ;
	assign n_2496 = (~x_727 & ~x_765) ;
	assign n_2495 = (~x_711 & ~x_715) ;
	assign n_2487 = (~x_118 & ~x_124) ;
	assign n_2486 = (~x_78 & ~x_109) ;
	assign n_2482 = (~x_258 & ~x_259) ;
	assign n_2481 = (~x_230 & ~x_248) ;
	assign n_2479 = (~x_286 & ~x_312) ;
	assign n_2478 = (~x_268 & ~x_278) ;
	assign n_2475 = (~x_171 & ~x_175) ;
	assign n_2474 = (~x_144 & ~x_161) ;
	assign n_2472 = (~x_191 & ~x_196) ;
	assign n_2471 = (~x_177 & ~x_184) ;
	assign n_8186 = (~n_2609 & n_8185) ;
	assign n_2603 = (~n_2601 & ~n_2602) ;
	assign n_2595 = (~x_609 & ~n_2593) ;
	assign n_2594 = (x_609 & n_2593) ;
	assign n_2581 = (~n_2578 & n_2580) ;
	assign n_2573 = (x_477 & n_53) ;
	assign n_2572 = (x_611 & n_51) ;
	assign n_2566 = (~n_2564 & ~n_2565) ;
	assign n_625 = (n_621 & n_624) ;
	assign n_618 = (n_614 & n_617) ;
	assign n_610 = (n_606 & n_609) ;
	assign n_603 = (n_599 & n_602) ;
	assign n_594 = (n_590 & n_593) ;
	assign n_587 = (n_583 & n_586) ;
	assign n_579 = (n_575 & n_578) ;
	assign n_572 = (n_568 & n_571) ;
	assign n_2531 = (n_2527 & n_2530) ;
	assign n_2524 = (n_2520 & n_2523) ;
	assign n_2516 = (n_2512 & n_2515) ;
	assign n_2509 = (n_2505 & n_2508) ;
	assign n_2500 = (n_2498 & n_2499) ;
	assign n_2497 = (n_2495 & n_2496) ;
	assign n_2493 = (~x_795 & ~x_802) ;
	assign n_2492 = (~x_778 & ~x_794) ;
	assign n_2488 = (n_2486 & n_2487) ;
	assign n_2483 = (n_2481 & n_2482) ;
	assign n_2480 = (n_2478 & n_2479) ;
	assign n_2476 = (n_2474 & n_2475) ;
	assign n_2473 = (n_2471 & n_2472) ;
	assign n_8187 = (~n_2603 & n_8186) ;
	assign n_2596 = (~n_2594 & ~n_2595) ;
	assign n_2583 = (~x_610 & ~n_2581) ;
	assign n_2582 = (x_610 & n_2581) ;
	assign n_2574 = (~n_2572 & ~n_2573) ;
	assign n_2567 = (n_20 & ~n_2566) ;
	assign n_2563 = (x_612 & n_18) ;
	assign n_2557 = (~x_613 & ~n_697) ;
	assign n_626 = (n_618 & n_625) ;
	assign n_611 = (n_603 & n_610) ;
	assign n_595 = (n_587 & n_594) ;
	assign n_580 = (n_572 & n_579) ;
	assign n_2532 = (n_2524 & n_2531) ;
	assign n_2517 = (n_2509 & n_2516) ;
	assign n_2501 = (n_2497 & n_2500) ;
	assign n_2494 = (n_2492 & n_2493) ;
	assign n_2489 = (~n_544 & n_2488) ;
	assign n_2484 = (n_2480 & n_2483) ;
	assign n_2477 = (n_2473 & n_2476) ;
	assign n_8188 = (~n_2596 & n_8187) ;
	assign n_2584 = (~n_2582 & ~n_2583) ;
	assign n_2576 = (~x_611 & n_2574) ;
	assign n_2575 = (x_611 & ~n_2574) ;
	assign n_2568 = (~n_2563 & ~n_2567) ;
	assign n_2558 = (i_5 & ~n_2557) ;
	assign n_2556 = (~x_370 & n_697) ;
	assign n_2543 = (~x_615 & ~n_64) ;
	assign n_627 = (n_611 & n_626) ;
	assign n_596 = (n_580 & n_595) ;
	assign n_2533 = (n_2517 & n_2532) ;
	assign n_2502 = (n_2494 & n_2501) ;
	assign n_2490 = (n_1820 & n_2489) ;
	assign n_2485 = (n_2477 & n_2484) ;
	assign n_8189 = (~n_2584 & n_8188) ;
	assign n_2577 = (~n_2575 & ~n_2576) ;
	assign n_2570 = (~x_612 & n_2568) ;
	assign n_2569 = (x_612 & ~n_2568) ;
	assign n_2559 = (~n_2556 & n_2558) ;
	assign n_2551 = (i_14 & n_948) ;
	assign n_2550 = (x_614 & n_945) ;
	assign n_2544 = (n_66 & ~n_2543) ;
	assign n_628 = (n_596 & n_627) ;
	assign n_2541 = (x_615 & ~n_59) ;
	assign n_2534 = (n_2502 & n_2533) ;
	assign n_2491 = (n_2485 & n_2490) ;
	assign n_8190 = (~n_2577 & n_8189) ;
	assign n_2571 = (~n_2569 & ~n_2570) ;
	assign n_2561 = (~x_613 & ~n_2559) ;
	assign n_2560 = (x_613 & n_2559) ;
	assign n_2552 = (~n_2550 & ~n_2551) ;
	assign n_2545 = (n_628 & n_2544) ;
	assign n_2542 = (n_978 & n_2541) ;
	assign n_2535 = (n_2491 & n_2534) ;
	assign n_2470 = (x_616 & ~n_1820) ;
	assign n_8191 = (~n_2571 & n_8190) ;
	assign n_2562 = (~n_2560 & ~n_2561) ;
	assign n_2554 = (~x_614 & n_2552) ;
	assign n_2553 = (x_614 & ~n_2552) ;
	assign n_2546 = (~n_2542 & ~n_2545) ;
	assign n_2536 = (~n_2470 & ~n_2535) ;
	assign n_2464 = (~x_617 & ~n_936) ;
	assign n_8192 = (~n_2562 & n_8191) ;
	assign n_2555 = (~n_2553 & ~n_2554) ;
	assign n_2548 = (~x_615 & n_2546) ;
	assign n_2547 = (x_615 & ~n_2546) ;
	assign n_2537 = (n_2348 & ~n_2536) ;
	assign n_2465 = (i_5 & ~n_2464) ;
	assign n_2463 = (~i_14 & n_936) ;
	assign n_2457 = (~x_618 & ~n_630) ;
	assign n_8193 = (~n_2555 & n_8192) ;
	assign n_2549 = (~n_2547 & ~n_2548) ;
	assign n_2539 = (~x_616 & ~n_2537) ;
	assign n_2538 = (x_616 & n_2537) ;
	assign n_2466 = (~n_2463 & n_2465) ;
	assign n_2458 = (i_5 & ~n_2457) ;
	assign n_2456 = (~i_33 & n_630) ;
	assign n_8194 = (~n_2549 & n_8193) ;
	assign n_2540 = (~n_2538 & ~n_2539) ;
	assign n_2468 = (~x_617 & ~n_2466) ;
	assign n_2467 = (x_617 & n_2466) ;
	assign n_2459 = (~n_2456 & n_2458) ;
	assign n_2451 = (~n_362 & n_35) ;
	assign n_2450 = (x_619 & n_36) ;
	assign n_2444 = (~x_620 & ~n_630) ;
	assign n_8195 = (~n_2540 & n_8194) ;
	assign n_2469 = (~n_2467 & ~n_2468) ;
	assign n_2461 = (~x_618 & ~n_2459) ;
	assign n_2460 = (x_618 & n_2459) ;
	assign n_2452 = (~n_2450 & ~n_2451) ;
	assign n_2445 = (i_5 & ~n_2444) ;
	assign n_2443 = (~i_19 & n_630) ;
	assign n_2437 = (i_40 & n_64) ;
	assign n_8196 = (~n_2469 & n_8195) ;
	assign n_2462 = (~n_2460 & ~n_2461) ;
	assign n_2454 = (~x_619 & n_2452) ;
	assign n_2453 = (x_619 & ~n_2452) ;
	assign n_2446 = (~n_2443 & n_2445) ;
	assign n_2438 = (n_66 & n_2437) ;
	assign n_2436 = (x_621 & n_978) ;
	assign n_2430 = (~x_622 & ~n_697) ;
	assign n_2384 = (~x_382 & n_1949) ;
	assign n_2383 = (x_382 & ~n_1949) ;
	assign n_8197 = (~n_2462 & n_8196) ;
	assign n_2455 = (~n_2453 & ~n_2454) ;
	assign n_2448 = (~x_620 & ~n_2446) ;
	assign n_2447 = (x_620 & n_2446) ;
	assign n_2439 = (~n_2436 & ~n_2438) ;
	assign n_2431 = (i_5 & ~n_2430) ;
	assign n_2429 = (~x_112 & n_697) ;
	assign n_2423 = (~x_623 & ~n_936) ;
	assign n_2385 = (~n_2383 & ~n_2384) ;
	assign n_2382 = (~n_1939 & ~n_1940) ;
	assign n_8198 = (~n_2455 & n_8197) ;
	assign n_2449 = (~n_2447 & ~n_2448) ;
	assign n_2441 = (~x_621 & n_2439) ;
	assign n_2440 = (x_621 & ~n_2439) ;
	assign n_2432 = (~n_2429 & n_2431) ;
	assign n_2424 = (i_5 & ~n_2423) ;
	assign n_2422 = (~i_28 & n_936) ;
	assign n_2394 = (~x_627 & n_6) ;
	assign n_2387 = (n_2382 & ~n_2385) ;
	assign n_8199 = (~n_2449 & n_8198) ;
	assign n_2442 = (~n_2440 & ~n_2441) ;
	assign n_2434 = (~x_622 & ~n_2432) ;
	assign n_2433 = (x_622 & n_2432) ;
	assign n_2425 = (~n_2422 & n_2424) ;
	assign n_2417 = (x_359 & n_53) ;
	assign n_2416 = (x_624 & n_51) ;
	assign n_2410 = (i_53 & n_59) ;
	assign n_2395 = (~n_2393 & ~n_2394) ;
	assign n_2390 = (x_627 & ~n_697) ;
	assign n_2388 = (n_697 & ~n_2387) ;
	assign n_2386 = (~n_2382 & n_2385) ;
	assign n_8200 = (~n_2442 & n_8199) ;
	assign n_2435 = (~n_2433 & ~n_2434) ;
	assign n_2427 = (~x_623 & ~n_2425) ;
	assign n_2426 = (x_623 & n_2425) ;
	assign n_2418 = (~n_2416 & ~n_2417) ;
	assign n_2411 = (n_66 & n_2410) ;
	assign n_2409 = (x_625 & n_60) ;
	assign n_2396 = (n_629 & ~n_2395) ;
	assign n_2391 = (~n_629 & ~n_2390) ;
	assign n_2389 = (~n_2386 & n_2388) ;
	assign n_8201 = (~n_2435 & n_8200) ;
	assign n_2428 = (~n_2426 & ~n_2427) ;
	assign n_2420 = (~x_624 & n_2418) ;
	assign n_2419 = (x_624 & ~n_2418) ;
	assign n_2412 = (~n_2409 & ~n_2411) ;
	assign n_2404 = (i_54 & n_948) ;
	assign n_2403 = (x_626 & n_945) ;
	assign n_2397 = (n_902 & ~n_2396) ;
	assign n_2392 = (~n_2389 & n_2391) ;
	assign n_8202 = (~n_2428 & n_8201) ;
	assign n_2421 = (~n_2419 & ~n_2420) ;
	assign n_2414 = (~x_625 & n_2412) ;
	assign n_2413 = (x_625 & ~n_2412) ;
	assign n_2405 = (~n_2403 & ~n_2404) ;
	assign n_2398 = (~n_2392 & n_2397) ;
	assign n_2381 = (x_627 & n_699) ;
	assign n_8203 = (~n_2421 & n_8202) ;
	assign n_2415 = (~n_2413 & ~n_2414) ;
	assign n_2407 = (~x_626 & n_2405) ;
	assign n_2406 = (x_626 & ~n_2405) ;
	assign n_2399 = (~n_2381 & ~n_2398) ;
	assign n_8204 = (~n_2415 & n_8203) ;
	assign n_2408 = (~n_2406 & ~n_2407) ;
	assign n_2401 = (~x_627 & n_2399) ;
	assign n_2400 = (x_627 & ~n_2399) ;
	assign n_2369 = (~x_630 & ~n_936) ;
	assign n_8205 = (~n_2408 & n_8204) ;
	assign n_2402 = (~n_2400 & ~n_2401) ;
	assign n_2379 = (~x_628 & n_497) ;
	assign n_2378 = (x_628 & ~n_497) ;
	assign n_2370 = (i_5 & ~n_2369) ;
	assign n_2368 = (~i_55 & n_936) ;
	assign n_8206 = (~n_2402 & n_8205) ;
	assign n_2380 = (~n_2378 & ~n_2379) ;
	assign n_2376 = (~x_629 & n_242) ;
	assign n_2375 = (x_629 & ~n_242) ;
	assign n_2371 = (~n_2368 & n_2370) ;
	assign n_2363 = (~n_257 & n_1009) ;
	assign n_2362 = (x_631 & n_1007) ;
	assign n_2356 = (i_47 & n_64) ;
	assign n_8207 = (~n_2380 & n_8206) ;
	assign n_2377 = (~n_2375 & ~n_2376) ;
	assign n_2373 = (~x_630 & ~n_2371) ;
	assign n_2372 = (x_630 & n_2371) ;
	assign n_2364 = (~n_2362 & ~n_2363) ;
	assign n_2357 = (n_66 & n_2356) ;
	assign n_2355 = (x_632 & n_978) ;
	assign n_2349 = (x_376 & n_697) ;
	assign n_8208 = (~n_2377 & n_8207) ;
	assign n_2374 = (~n_2372 & ~n_2373) ;
	assign n_2366 = (~x_631 & n_2364) ;
	assign n_2365 = (x_631 & ~n_2364) ;
	assign n_2358 = (~n_2355 & ~n_2357) ;
	assign n_2350 = (n_2348 & n_2349) ;
	assign n_2347 = (x_633 & n_698) ;
	assign n_2341 = (~x_634 & ~n_630) ;
	assign n_8209 = (~n_2374 & n_8208) ;
	assign n_2367 = (~n_2365 & ~n_2366) ;
	assign n_2360 = (~x_632 & n_2358) ;
	assign n_2359 = (x_632 & ~n_2358) ;
	assign n_2351 = (~n_2347 & ~n_2350) ;
	assign n_2342 = (i_5 & ~n_2341) ;
	assign n_2340 = (~i_63 & n_630) ;
	assign n_2334 = (~x_635 & ~n_544) ;
	assign n_2326 = (~i_20 & n_669) ;
	assign n_8210 = (~n_2367 & n_8209) ;
	assign n_2361 = (~n_2359 & ~n_2360) ;
	assign n_2353 = (~x_633 & n_2351) ;
	assign n_2352 = (x_633 & ~n_2351) ;
	assign n_2343 = (~n_2340 & n_2342) ;
	assign n_2335 = (i_5 & ~n_2334) ;
	assign n_2333 = (~i_31 & n_544) ;
	assign n_2327 = (i_5 & ~n_2326) ;
	assign n_2325 = (~x_633 & n_662) ;
	assign n_8211 = (~n_2361 & n_8210) ;
	assign n_2354 = (~n_2352 & ~n_2353) ;
	assign n_2345 = (~x_634 & ~n_2343) ;
	assign n_2344 = (x_634 & n_2343) ;
	assign n_2336 = (~n_2333 & n_2335) ;
	assign n_2328 = (~n_2325 & n_2327) ;
	assign n_2324 = (~x_636 & ~n_665) ;
	assign n_2318 = (i_15 & n_64) ;
	assign n_1118 = (~x_777 & ~n_669) ;
	assign n_8212 = (~n_2354 & n_8211) ;
	assign n_2346 = (~n_2344 & ~n_2345) ;
	assign n_2338 = (~x_635 & ~n_2336) ;
	assign n_2337 = (x_635 & n_2336) ;
	assign n_2329 = (~n_2324 & n_2328) ;
	assign n_2319 = (n_66 & n_2318) ;
	assign n_2317 = (x_637 & n_978) ;
	assign n_2311 = (x_638 & n_1118) ;
	assign n_8213 = (~n_2346 & n_8212) ;
	assign n_2339 = (~n_2337 & ~n_2338) ;
	assign n_2331 = (~x_636 & ~n_2329) ;
	assign n_2330 = (x_636 & n_2329) ;
	assign n_2320 = (~n_2317 & ~n_2319) ;
	assign n_2312 = (~n_697 & ~n_2311) ;
	assign n_8214 = (~n_2339 & n_8213) ;
	assign n_2332 = (~n_2330 & ~n_2331) ;
	assign n_2322 = (~x_637 & n_2320) ;
	assign n_2321 = (x_637 & ~n_2320) ;
	assign n_2313 = (i_5 & ~n_2312) ;
	assign n_2306 = (~n_376 & n_35) ;
	assign n_2305 = (x_639 & n_36) ;
	assign n_2299 = (~x_640 & ~n_936) ;
	assign n_2257 = (~n_478 & ~n_479) ;
	assign n_8215 = (~n_2332 & n_8214) ;
	assign n_2323 = (~n_2321 & ~n_2322) ;
	assign n_2315 = (~x_638 & ~n_2313) ;
	assign n_2314 = (x_638 & n_2313) ;
	assign n_2307 = (~n_2305 & ~n_2306) ;
	assign n_2300 = (i_5 & ~n_2299) ;
	assign n_2298 = (~i_10 & n_936) ;
	assign n_2259 = (~x_295 & ~n_2257) ;
	assign n_8216 = (~n_2323 & n_8215) ;
	assign n_2316 = (~n_2314 & ~n_2315) ;
	assign n_2309 = (~x_639 & n_2307) ;
	assign n_2308 = (x_639 & ~n_2307) ;
	assign n_2301 = (~n_2298 & n_2300) ;
	assign n_2289 = (i_33 & n_64) ;
	assign n_2260 = (n_527 & ~n_2259) ;
	assign n_2258 = (x_295 & n_2257) ;
	assign n_8217 = (~n_2316 & n_8216) ;
	assign n_2310 = (~n_2308 & ~n_2309) ;
	assign n_2303 = (~x_640 & ~n_2301) ;
	assign n_2302 = (x_640 & n_2301) ;
	assign n_2290 = (n_66 & n_2289) ;
	assign n_2288 = (x_642 & n_978) ;
	assign n_2282 = (~x_643 & ~n_936) ;
	assign n_2267 = (n_6 & n_482) ;
	assign n_2261 = (~n_2258 & n_2260) ;
	assign n_8218 = (~n_2310 & n_8217) ;
	assign n_2304 = (~n_2302 & ~n_2303) ;
	assign n_2296 = (~x_641 & n_143) ;
	assign n_2295 = (x_641 & ~n_143) ;
	assign n_2291 = (~n_2288 & ~n_2290) ;
	assign n_2283 = (i_5 & ~n_2282) ;
	assign n_2281 = (~i_16 & n_936) ;
	assign n_2268 = (~n_2266 & ~n_2267) ;
	assign n_2263 = (n_482 & n_2261) ;
	assign n_8219 = (~n_2304 & n_8218) ;
	assign n_2297 = (~n_2295 & ~n_2296) ;
	assign n_2293 = (~x_642 & n_2291) ;
	assign n_2292 = (x_642 & ~n_2291) ;
	assign n_2284 = (~n_2281 & n_2283) ;
	assign n_2276 = (~n_421 & n_1009) ;
	assign n_2275 = (x_644 & n_1007) ;
	assign n_2269 = (n_1 & ~n_2268) ;
	assign n_2264 = (~n_1 & ~n_2263) ;
	assign n_2262 = (~n_482 & ~n_2261) ;
	assign n_8220 = (~n_2297 & n_8219) ;
	assign n_2294 = (~n_2292 & ~n_2293) ;
	assign n_2286 = (~x_643 & ~n_2284) ;
	assign n_2285 = (x_643 & n_2284) ;
	assign n_2277 = (~n_2275 & ~n_2276) ;
	assign n_2270 = (i_5 & ~n_2269) ;
	assign n_2265 = (~n_2262 & n_2264) ;
	assign n_2251 = (i_27 & n_64) ;
	assign n_8221 = (~n_2294 & n_8220) ;
	assign n_2287 = (~n_2285 & ~n_2286) ;
	assign n_2279 = (~x_644 & n_2277) ;
	assign n_2278 = (x_644 & ~n_2277) ;
	assign n_2271 = (~n_2265 & n_2270) ;
	assign n_2252 = (n_66 & n_2251) ;
	assign n_2250 = (x_646 & n_978) ;
	assign n_2237 = (~i_67 & n_669) ;
	assign n_2235 = (~x_613 & ~n_544) ;
	assign n_8222 = (~n_2287 & n_8221) ;
	assign n_2280 = (~n_2278 & ~n_2279) ;
	assign n_2273 = (~x_645 & ~n_2271) ;
	assign n_2272 = (x_645 & n_2271) ;
	assign n_2253 = (~n_2250 & ~n_2252) ;
	assign n_2245 = (x_773 & n_53) ;
	assign n_2244 = (x_647 & n_51) ;
	assign n_2238 = (i_5 & ~n_2237) ;
	assign n_2236 = (n_662 & n_2235) ;
	assign n_2184 = (~n_199 & ~n_200) ;
	assign n_8223 = (~n_2280 & n_8222) ;
	assign n_2274 = (~n_2272 & ~n_2273) ;
	assign n_2255 = (~x_646 & n_2253) ;
	assign n_2254 = (x_646 & ~n_2253) ;
	assign n_2246 = (~n_2244 & ~n_2245) ;
	assign n_2239 = (~n_2236 & n_2238) ;
	assign n_2234 = (~x_648 & ~n_665) ;
	assign n_2228 = (~x_649 & ~n_630) ;
	assign n_2186 = (~x_756 & ~n_2184) ;
	assign n_8224 = (~n_2274 & n_8223) ;
	assign n_2256 = (~n_2254 & ~n_2255) ;
	assign n_2248 = (~x_647 & n_2246) ;
	assign n_2247 = (x_647 & ~n_2246) ;
	assign n_2240 = (~n_2234 & n_2239) ;
	assign n_2229 = (i_5 & ~n_2228) ;
	assign n_2227 = (~i_47 & n_630) ;
	assign n_2187 = (~x_332 & ~n_2186) ;
	assign n_2185 = (x_756 & n_2184) ;
	assign n_8225 = (~n_2256 & n_8224) ;
	assign n_2249 = (~n_2247 & ~n_2248) ;
	assign n_2242 = (~x_648 & ~n_2240) ;
	assign n_2241 = (x_648 & n_2240) ;
	assign n_2230 = (~n_2227 & n_2229) ;
	assign n_2222 = (n_35 & ~n_467) ;
	assign n_2221 = (x_650 & n_36) ;
	assign n_2215 = (~x_651 & ~n_630) ;
	assign n_2188 = (~n_2185 & n_2187) ;
	assign n_8226 = (~n_2249 & n_8225) ;
	assign n_2243 = (~n_2241 & ~n_2242) ;
	assign n_2232 = (~x_649 & ~n_2230) ;
	assign n_2231 = (x_649 & n_2230) ;
	assign n_2223 = (~n_2221 & ~n_2222) ;
	assign n_2216 = (i_5 & ~n_2215) ;
	assign n_2214 = (~i_56 & n_630) ;
	assign n_2190 = (n_203 & ~n_2188) ;
	assign n_8227 = (~n_2243 & n_8226) ;
	assign n_2233 = (~n_2231 & ~n_2232) ;
	assign n_2225 = (~x_650 & n_2223) ;
	assign n_2224 = (x_650 & ~n_2223) ;
	assign n_2217 = (~n_2214 & n_2216) ;
	assign n_2209 = (n_35 & ~n_436) ;
	assign n_2208 = (x_652 & n_36) ;
	assign n_2202 = (i_39 & n_64) ;
	assign n_2194 = (~n_203 & ~n_1606) ;
	assign n_2193 = (i_8 & n_7) ;
	assign n_2191 = (x_664 & ~n_2190) ;
	assign n_2189 = (~n_203 & n_2188) ;
	assign n_8228 = (~n_2233 & n_8227) ;
	assign n_2226 = (~n_2224 & ~n_2225) ;
	assign n_2219 = (~x_651 & ~n_2217) ;
	assign n_2218 = (x_651 & n_2217) ;
	assign n_2210 = (~n_2208 & ~n_2209) ;
	assign n_2203 = (n_66 & n_2202) ;
	assign n_2201 = (x_653 & n_978) ;
	assign n_2195 = (~n_2193 & ~n_2194) ;
	assign n_2192 = (~n_2189 & n_2191) ;
	assign n_2177 = (~i_40 & n_669) ;
	assign n_2175 = (~x_477 & ~n_544) ;
	assign n_2139 = (~x_180 & n_864) ;
	assign n_2138 = (x_180 & ~n_864) ;
	assign n_8229 = (~n_2226 & n_8228) ;
	assign n_2220 = (~n_2218 & ~n_2219) ;
	assign n_2212 = (~x_652 & n_2210) ;
	assign n_2211 = (x_652 & ~n_2210) ;
	assign n_2204 = (~n_2201 & ~n_2203) ;
	assign n_2196 = (~n_2192 & n_2195) ;
	assign n_2178 = (i_5 & ~n_2177) ;
	assign n_2176 = (n_662 & n_2175) ;
	assign n_2140 = (~n_2138 & ~n_2139) ;
	assign n_2137 = (~n_854 & ~n_855) ;
	assign n_8230 = (~n_2220 & n_8229) ;
	assign n_2213 = (~n_2211 & ~n_2212) ;
	assign n_2206 = (~x_653 & n_2204) ;
	assign n_2205 = (x_653 & ~n_2204) ;
	assign n_2197 = (i_5 & ~n_2196) ;
	assign n_2179 = (~n_2176 & n_2178) ;
	assign n_2174 = (~x_655 & ~n_665) ;
	assign n_2149 = (i_46 & ~n_6) ;
	assign n_2142 = (n_2137 & ~n_2140) ;
	assign n_8231 = (~n_2213 & n_8230) ;
	assign n_2207 = (~n_2205 & ~n_2206) ;
	assign n_2199 = (~x_654 & ~n_2197) ;
	assign n_2198 = (x_654 & n_2197) ;
	assign n_2180 = (~n_2174 & n_2179) ;
	assign n_2169 = (~n_362 & n_1009) ;
	assign n_2168 = (x_656 & n_1007) ;
	assign n_2162 = (~x_657 & ~n_630) ;
	assign n_2150 = (n_629 & ~n_2149) ;
	assign n_2148 = (x_659 & n_6) ;
	assign n_2145 = (x_659 & ~n_697) ;
	assign n_2143 = (n_697 & ~n_2142) ;
	assign n_2141 = (~n_2137 & n_2140) ;
	assign n_8232 = (~n_2207 & n_8231) ;
	assign n_2200 = (~n_2198 & ~n_2199) ;
	assign n_2182 = (~x_655 & ~n_2180) ;
	assign n_2181 = (x_655 & n_2180) ;
	assign n_2170 = (~n_2168 & ~n_2169) ;
	assign n_2163 = (i_5 & ~n_2162) ;
	assign n_2161 = (~i_45 & n_630) ;
	assign n_2151 = (~n_2148 & n_2150) ;
	assign n_2146 = (~n_629 & ~n_2145) ;
	assign n_2144 = (~n_2141 & n_2143) ;
	assign n_8233 = (~n_2200 & n_8232) ;
	assign n_2183 = (~n_2181 & ~n_2182) ;
	assign n_2172 = (~x_656 & n_2170) ;
	assign n_2171 = (x_656 & ~n_2170) ;
	assign n_2164 = (~n_2161 & n_2163) ;
	assign n_2152 = (n_902 & ~n_2151) ;
	assign n_2147 = (~n_2144 & n_2146) ;
	assign n_8234 = (~n_2183 & n_8233) ;
	assign n_2173 = (~n_2171 & ~n_2172) ;
	assign n_2166 = (~x_657 & ~n_2164) ;
	assign n_2165 = (x_657 & n_2164) ;
	assign n_2153 = (~n_2147 & n_2152) ;
	assign n_2136 = (x_659 & n_699) ;
	assign n_8235 = (~n_2173 & n_8234) ;
	assign n_2167 = (~n_2165 & ~n_2166) ;
	assign n_2159 = (~x_658 & n_107) ;
	assign n_2158 = (x_658 & ~n_107) ;
	assign n_2154 = (~n_2136 & ~n_2153) ;
	assign n_2131 = (i_7 & n_948) ;
	assign n_2130 = (x_660 & n_945) ;
	assign n_8236 = (~n_2167 & n_8235) ;
	assign n_2160 = (~n_2158 & ~n_2159) ;
	assign n_2156 = (~x_659 & n_2154) ;
	assign n_2155 = (x_659 & ~n_2154) ;
	assign n_2132 = (~n_2130 & ~n_2131) ;
	assign n_2125 = (i_40 & n_948) ;
	assign n_2124 = (x_661 & n_945) ;
	assign n_8237 = (~n_2160 & n_8236) ;
	assign n_2157 = (~n_2155 & ~n_2156) ;
	assign n_2134 = (~x_660 & n_2132) ;
	assign n_2133 = (x_660 & ~n_2132) ;
	assign n_2126 = (~n_2124 & ~n_2125) ;
	assign n_8238 = (~n_2157 & n_8237) ;
	assign n_2135 = (~n_2133 & ~n_2134) ;
	assign n_2128 = (~x_661 & n_2126) ;
	assign n_2127 = (x_661 & ~n_2126) ;
	assign n_2116 = (x_712 & n_35) ;
	assign n_2115 = (x_663 & n_36) ;
	assign n_8239 = (~n_2135 & n_8238) ;
	assign n_2129 = (~n_2127 & ~n_2128) ;
	assign n_2122 = (~x_662 & n_302) ;
	assign n_2121 = (x_662 & ~n_302) ;
	assign n_2117 = (~n_2115 & ~n_2116) ;
	assign n_8240 = (~n_2129 & n_8239) ;
	assign n_2123 = (~n_2121 & ~n_2122) ;
	assign n_2119 = (~x_663 & n_2117) ;
	assign n_2118 = (x_663 & ~n_2117) ;
	assign n_2111 = (~n_20 & ~n_1009) ;
	assign n_2106 = (i_26 & n_948) ;
	assign n_2105 = (x_665 & n_945) ;
	assign n_2099 = (~x_666 & ~n_936) ;
	assign n_8241 = (~n_2123 & n_8240) ;
	assign n_2120 = (~n_2118 & ~n_2119) ;
	assign n_2113 = (~x_664 & n_2111) ;
	assign n_2112 = (x_664 & ~n_2111) ;
	assign n_2107 = (~n_2105 & ~n_2106) ;
	assign n_2100 = (i_5 & ~n_2099) ;
	assign n_2098 = (~i_62 & n_936) ;
	assign n_2092 = (i_51 & n_59) ;
	assign n_8242 = (~n_2120 & n_8241) ;
	assign n_2114 = (~n_2112 & ~n_2113) ;
	assign n_2109 = (~x_665 & n_2107) ;
	assign n_2108 = (x_665 & ~n_2107) ;
	assign n_2101 = (~n_2098 & n_2100) ;
	assign n_2093 = (n_66 & n_2092) ;
	assign n_2091 = (x_667 & n_60) ;
	assign n_2085 = (~x_668 & ~n_544) ;
	assign n_2077 = (i_6 & n_7) ;
	assign n_2076 = (x_113 & ~n_16) ;
	assign n_8243 = (~n_2114 & n_8242) ;
	assign n_2110 = (~n_2108 & ~n_2109) ;
	assign n_2103 = (~x_666 & ~n_2101) ;
	assign n_2102 = (x_666 & n_2101) ;
	assign n_2094 = (~n_2091 & ~n_2093) ;
	assign n_2086 = (i_5 & ~n_2085) ;
	assign n_2084 = (~i_66 & n_544) ;
	assign n_2078 = (~n_2076 & ~n_2077) ;
	assign n_2068 = (i_22 & n_7) ;
	assign n_2067 = (x_352 & ~n_16) ;
	assign n_8244 = (~n_2110 & n_8243) ;
	assign n_2104 = (~n_2102 & ~n_2103) ;
	assign n_2096 = (~x_667 & n_2094) ;
	assign n_2095 = (x_667 & ~n_2094) ;
	assign n_2087 = (~n_2084 & n_2086) ;
	assign n_2079 = (n_20 & ~n_2078) ;
	assign n_2075 = (x_669 & n_18) ;
	assign n_2069 = (~n_2067 & ~n_2068) ;
	assign n_2059 = (i_47 & n_7) ;
	assign n_2058 = (x_188 & ~n_16) ;
	assign n_8245 = (~n_2104 & n_8244) ;
	assign n_2097 = (~n_2095 & ~n_2096) ;
	assign n_2089 = (~x_668 & ~n_2087) ;
	assign n_2088 = (x_668 & n_2087) ;
	assign n_2080 = (~n_2075 & ~n_2079) ;
	assign n_2070 = (n_20 & ~n_2069) ;
	assign n_2066 = (x_670 & n_18) ;
	assign n_2060 = (~n_2058 & ~n_2059) ;
	assign n_8246 = (~n_2097 & n_8245) ;
	assign n_2090 = (~n_2088 & ~n_2089) ;
	assign n_2082 = (~x_669 & n_2080) ;
	assign n_2081 = (x_669 & ~n_2080) ;
	assign n_2071 = (~n_2066 & ~n_2070) ;
	assign n_2061 = (n_20 & ~n_2060) ;
	assign n_2057 = (x_671 & n_18) ;
	assign n_2051 = (i_10 & n_59) ;
	assign n_8247 = (~n_2090 & n_8246) ;
	assign n_2083 = (~n_2081 & ~n_2082) ;
	assign n_2073 = (~x_670 & n_2071) ;
	assign n_2072 = (x_670 & ~n_2071) ;
	assign n_2062 = (~n_2057 & ~n_2061) ;
	assign n_2052 = (n_66 & n_2051) ;
	assign n_2050 = (x_672 & n_60) ;
	assign n_8248 = (~n_2083 & n_8247) ;
	assign n_2074 = (~n_2072 & ~n_2073) ;
	assign n_2064 = (~x_671 & n_2062) ;
	assign n_2063 = (x_671 & ~n_2062) ;
	assign n_2053 = (~n_2050 & ~n_2052) ;
	assign n_2045 = (i_31 & n_948) ;
	assign n_2044 = (x_673 & n_945) ;
	assign n_8249 = (~n_2074 & n_8248) ;
	assign n_2065 = (~n_2063 & ~n_2064) ;
	assign n_2055 = (~x_672 & n_2053) ;
	assign n_2054 = (x_672 & ~n_2053) ;
	assign n_2046 = (~n_2044 & ~n_2045) ;
	assign n_2039 = (x_112 & n_53) ;
	assign n_2038 = (x_674 & n_51) ;
	assign n_2032 = (~x_675 & ~n_544) ;
	assign n_8250 = (~n_2065 & n_8249) ;
	assign n_2056 = (~n_2054 & ~n_2055) ;
	assign n_2048 = (~x_673 & n_2046) ;
	assign n_2047 = (x_673 & ~n_2046) ;
	assign n_2040 = (~n_2038 & ~n_2039) ;
	assign n_2033 = (i_5 & ~n_2032) ;
	assign n_2031 = (~i_60 & n_544) ;
	assign n_8251 = (~n_2056 & n_8250) ;
	assign n_2049 = (~n_2047 & ~n_2048) ;
	assign n_2042 = (~x_674 & n_2040) ;
	assign n_2041 = (x_674 & ~n_2040) ;
	assign n_2034 = (~n_2031 & n_2033) ;
	assign n_2026 = (x_792 & n_35) ;
	assign n_2025 = (x_676 & n_36) ;
	assign n_2019 = (~x_677 & ~n_697) ;
	assign n_2011 = (i_68 & n_7) ;
	assign n_2010 = (x_485 & ~n_16) ;
	assign n_8252 = (~n_2049 & n_8251) ;
	assign n_2043 = (~n_2041 & ~n_2042) ;
	assign n_2036 = (~x_675 & ~n_2034) ;
	assign n_2035 = (x_675 & n_2034) ;
	assign n_2027 = (~n_2025 & ~n_2026) ;
	assign n_2020 = (i_5 & ~n_2019) ;
	assign n_2018 = (~x_320 & n_697) ;
	assign n_2012 = (~n_2010 & ~n_2011) ;
	assign n_1965 = (~x_402 & n_1963) ;
	assign n_1964 = (x_402 & ~n_1963) ;
	assign n_8253 = (~n_2043 & n_8252) ;
	assign n_2037 = (~n_2035 & ~n_2036) ;
	assign n_2029 = (~x_676 & n_2027) ;
	assign n_2028 = (x_676 & ~n_2027) ;
	assign n_2021 = (~n_2018 & n_2020) ;
	assign n_2013 = (n_20 & ~n_2012) ;
	assign n_2009 = (x_678 & n_18) ;
	assign n_1966 = (~n_1964 & ~n_1965) ;
	assign n_1954 = (~n_1952 & ~n_1953) ;
	assign n_8254 = (~n_2037 & n_8253) ;
	assign n_2030 = (~n_2028 & ~n_2029) ;
	assign n_2023 = (~x_677 & ~n_2021) ;
	assign n_2022 = (x_677 & n_2021) ;
	assign n_2014 = (~n_2009 & ~n_2013) ;
	assign n_2004 = (x_186 & n_53) ;
	assign n_2003 = (x_679 & n_51) ;
	assign n_1975 = (i_39 & ~n_6) ;
	assign n_1968 = (n_1954 & ~n_1966) ;
	assign n_8255 = (~n_2030 & n_8254) ;
	assign n_2024 = (~n_2022 & ~n_2023) ;
	assign n_2016 = (~x_678 & n_2014) ;
	assign n_2015 = (x_678 & ~n_2014) ;
	assign n_2005 = (~n_2003 & ~n_2004) ;
	assign n_1998 = (i_43 & n_948) ;
	assign n_1997 = (x_680 & n_945) ;
	assign n_1976 = (n_629 & ~n_1975) ;
	assign n_1974 = (x_683 & n_6) ;
	assign n_1971 = (x_683 & ~n_697) ;
	assign n_1969 = (n_697 & ~n_1968) ;
	assign n_1967 = (~n_1954 & n_1966) ;
	assign n_8256 = (~n_2024 & n_8255) ;
	assign n_2017 = (~n_2015 & ~n_2016) ;
	assign n_2007 = (~x_679 & n_2005) ;
	assign n_2006 = (x_679 & ~n_2005) ;
	assign n_1999 = (~n_1997 & ~n_1998) ;
	assign n_1992 = (x_216 & n_53) ;
	assign n_1991 = (x_681 & n_51) ;
	assign n_1985 = (~x_682 & ~n_544) ;
	assign n_1977 = (~n_1974 & n_1976) ;
	assign n_1972 = (~n_629 & ~n_1971) ;
	assign n_1970 = (~n_1967 & n_1969) ;
	assign n_8257 = (~n_2017 & n_8256) ;
	assign n_2008 = (~n_2006 & ~n_2007) ;
	assign n_2001 = (~x_680 & n_1999) ;
	assign n_2000 = (x_680 & ~n_1999) ;
	assign n_1993 = (~n_1991 & ~n_1992) ;
	assign n_1986 = (i_5 & ~n_1985) ;
	assign n_1984 = (~i_29 & n_544) ;
	assign n_1978 = (n_902 & ~n_1977) ;
	assign n_1973 = (~n_1970 & n_1972) ;
	assign n_8258 = (~n_2008 & n_8257) ;
	assign n_2002 = (~n_2000 & ~n_2001) ;
	assign n_1995 = (~x_681 & n_1993) ;
	assign n_1994 = (x_681 & ~n_1993) ;
	assign n_1987 = (~n_1984 & n_1986) ;
	assign n_1979 = (~n_1973 & n_1978) ;
	assign n_1910 = (x_683 & n_699) ;
	assign n_1904 = (~x_684 & ~n_544) ;
	assign n_8259 = (~n_2002 & n_8258) ;
	assign n_1996 = (~n_1994 & ~n_1995) ;
	assign n_1989 = (~x_682 & ~n_1987) ;
	assign n_1988 = (x_682 & n_1987) ;
	assign n_1980 = (~n_1910 & ~n_1979) ;
	assign n_1905 = (i_5 & ~n_1904) ;
	assign n_1903 = (~i_9 & n_544) ;
	assign n_1897 = (~x_685 & ~n_544) ;
	assign n_8260 = (~n_1996 & n_8259) ;
	assign n_1990 = (~n_1988 & ~n_1989) ;
	assign n_1982 = (~x_683 & n_1980) ;
	assign n_1981 = (x_683 & ~n_1980) ;
	assign n_1906 = (~n_1903 & n_1905) ;
	assign n_1898 = (i_5 & ~n_1897) ;
	assign n_1896 = (~i_51 & n_544) ;
	assign n_1890 = (i_66 & n_59) ;
	assign n_8261 = (~n_1990 & n_8260) ;
	assign n_1983 = (~n_1981 & ~n_1982) ;
	assign n_1908 = (~x_684 & ~n_1906) ;
	assign n_1907 = (x_684 & n_1906) ;
	assign n_1899 = (~n_1896 & n_1898) ;
	assign n_1891 = (n_66 & n_1890) ;
	assign n_1889 = (x_686 & n_60) ;
	assign n_8262 = (~n_1983 & n_8261) ;
	assign n_1909 = (~n_1907 & ~n_1908) ;
	assign n_1901 = (~x_685 & ~n_1899) ;
	assign n_1900 = (x_685 & n_1899) ;
	assign n_1892 = (~n_1889 & ~n_1891) ;
	assign n_1884 = (~n_188 & n_35) ;
	assign n_1883 = (x_687 & n_36) ;
	assign n_1877 = (i_68 & n_59) ;
	assign n_8263 = (~n_1909 & n_8262) ;
	assign n_1902 = (~n_1900 & ~n_1901) ;
	assign n_1894 = (~x_686 & n_1892) ;
	assign n_1893 = (x_686 & ~n_1892) ;
	assign n_1885 = (~n_1883 & ~n_1884) ;
	assign n_1878 = (n_66 & n_1877) ;
	assign n_1876 = (x_688 & n_60) ;
	assign n_1870 = (~x_689 & ~n_630) ;
	assign n_1308 = (~i_9 & ~n_6) ;
	assign n_8264 = (~n_1902 & n_8263) ;
	assign n_1895 = (~n_1893 & ~n_1894) ;
	assign n_1887 = (~x_687 & n_1885) ;
	assign n_1886 = (x_687 & ~n_1885) ;
	assign n_1879 = (~n_1876 & ~n_1878) ;
	assign n_1871 = (i_5 & ~n_1870) ;
	assign n_1869 = (~i_6 & n_630) ;
	assign n_1856 = (n_629 & n_1308) ;
	assign n_8265 = (~n_1895 & n_8264) ;
	assign n_1888 = (~n_1886 & ~n_1887) ;
	assign n_1881 = (~x_688 & n_1879) ;
	assign n_1880 = (x_688 & ~n_1879) ;
	assign n_1872 = (~n_1869 & n_1871) ;
	assign n_1864 = (x_91 & n_53) ;
	assign n_1863 = (x_690 & n_51) ;
	assign n_1857 = (i_5 & ~n_1856) ;
	assign n_1855 = (~x_289 & n_662) ;
	assign n_8266 = (~n_1888 & n_8265) ;
	assign n_1882 = (~n_1880 & ~n_1881) ;
	assign n_1874 = (~x_689 & ~n_1872) ;
	assign n_1873 = (x_689 & n_1872) ;
	assign n_1865 = (~n_1863 & ~n_1864) ;
	assign n_1858 = (~n_1855 & n_1857) ;
	assign n_1854 = (~x_691 & ~n_665) ;
	assign n_8267 = (~n_1882 & n_8266) ;
	assign n_1875 = (~n_1873 & ~n_1874) ;
	assign n_1867 = (~x_690 & n_1865) ;
	assign n_1866 = (x_690 & ~n_1865) ;
	assign n_1859 = (~n_1854 & n_1858) ;
	assign n_1849 = (i_50 & n_948) ;
	assign n_1848 = (x_692 & n_945) ;
	assign n_1842 = (i_18 & n_59) ;
	assign n_8268 = (~n_1875 & n_8267) ;
	assign n_1868 = (~n_1866 & ~n_1867) ;
	assign n_1861 = (~x_691 & ~n_1859) ;
	assign n_1860 = (x_691 & n_1859) ;
	assign n_1850 = (~n_1848 & ~n_1849) ;
	assign n_1843 = (n_66 & n_1842) ;
	assign n_1841 = (x_693 & n_60) ;
	assign n_1835 = (i_31 & n_59) ;
	assign n_1793 = (~x_326 & n_1791) ;
	assign n_1792 = (x_326 & ~n_1791) ;
	assign n_8269 = (~n_1868 & n_8268) ;
	assign n_1862 = (~n_1860 & ~n_1861) ;
	assign n_1852 = (~x_692 & n_1850) ;
	assign n_1851 = (x_692 & ~n_1850) ;
	assign n_1844 = (~n_1841 & ~n_1843) ;
	assign n_1836 = (n_66 & n_1835) ;
	assign n_1834 = (x_694 & n_60) ;
	assign n_1794 = (~n_1792 & ~n_1793) ;
	assign n_1782 = (~n_1780 & ~n_1781) ;
	assign n_8270 = (~n_1862 & n_8269) ;
	assign n_1853 = (~n_1851 & ~n_1852) ;
	assign n_1846 = (~x_693 & n_1844) ;
	assign n_1845 = (x_693 & ~n_1844) ;
	assign n_1837 = (~n_1834 & ~n_1836) ;
	assign n_1821 = (x_697 & x_777) ;
	assign n_1803 = (i_33 & ~n_6) ;
	assign n_1796 = (n_1782 & ~n_1794) ;
	assign n_8271 = (~n_1853 & n_8270) ;
	assign n_1847 = (~n_1845 & ~n_1846) ;
	assign n_1839 = (~x_694 & n_1837) ;
	assign n_1838 = (x_694 & ~n_1837) ;
	assign n_1822 = (~n_1820 & n_1821) ;
	assign n_1819 = (n_1650 & ~n_1818) ;
	assign n_1804 = (n_629 & ~n_1803) ;
	assign n_1802 = (x_699 & n_6) ;
	assign n_1799 = (x_699 & ~n_697) ;
	assign n_1797 = (n_697 & ~n_1796) ;
	assign n_1795 = (~n_1782 & n_1794) ;
	assign n_8272 = (~n_1847 & n_8271) ;
	assign n_1840 = (~n_1838 & ~n_1839) ;
	assign n_1832 = (~x_695 & n_482) ;
	assign n_1831 = (x_695 & ~n_482) ;
	assign n_1823 = (~n_1819 & ~n_1822) ;
	assign n_1805 = (~n_1802 & n_1804) ;
	assign n_1800 = (~n_629 & ~n_1799) ;
	assign n_1798 = (~n_1795 & n_1797) ;
	assign n_8273 = (~n_1840 & n_8272) ;
	assign n_1833 = (~n_1831 & ~n_1832) ;
	assign n_1829 = (~x_696 & n_227) ;
	assign n_1828 = (x_696 & ~n_227) ;
	assign n_1824 = (i_5 & ~n_1823) ;
	assign n_1813 = (x_529 & n_53) ;
	assign n_1812 = (x_698 & n_51) ;
	assign n_1806 = (n_902 & ~n_1805) ;
	assign n_1801 = (~n_1798 & n_1800) ;
	assign n_8274 = (~n_1833 & n_8273) ;
	assign n_1830 = (~n_1828 & ~n_1829) ;
	assign n_1826 = (~x_697 & ~n_1824) ;
	assign n_1825 = (x_697 & n_1824) ;
	assign n_1814 = (~n_1812 & ~n_1813) ;
	assign n_1807 = (~n_1801 & n_1806) ;
	assign n_1777 = (x_699 & n_699) ;
	assign n_1771 = (~x_700 & ~n_544) ;
	assign n_8275 = (~n_1830 & n_8274) ;
	assign n_1827 = (~n_1825 & ~n_1826) ;
	assign n_1816 = (~x_698 & n_1814) ;
	assign n_1815 = (x_698 & ~n_1814) ;
	assign n_1808 = (~n_1777 & ~n_1807) ;
	assign n_1772 = (i_5 & ~n_1771) ;
	assign n_1770 = (~i_67 & n_544) ;
	assign n_1764 = (i_13 & n_64) ;
	assign n_8276 = (~n_1827 & n_8275) ;
	assign n_1817 = (~n_1815 & ~n_1816) ;
	assign n_1810 = (~x_699 & n_1808) ;
	assign n_1809 = (x_699 & ~n_1808) ;
	assign n_1773 = (~n_1770 & n_1772) ;
	assign n_1765 = (n_66 & n_1764) ;
	assign n_1763 = (x_701 & n_978) ;
	assign n_1757 = (~x_702 & ~n_544) ;
	assign n_1749 = (~i_34 & n_669) ;
	assign n_8277 = (~n_1817 & n_8276) ;
	assign n_1811 = (~n_1809 & ~n_1810) ;
	assign n_1775 = (~x_700 & ~n_1773) ;
	assign n_1774 = (x_700 & n_1773) ;
	assign n_1766 = (~n_1763 & ~n_1765) ;
	assign n_1758 = (i_5 & ~n_1757) ;
	assign n_1756 = (~i_55 & n_544) ;
	assign n_1750 = (i_5 & ~n_1749) ;
	assign n_1748 = (~x_567 & n_662) ;
	assign n_8278 = (~n_1811 & n_8277) ;
	assign n_1776 = (~n_1774 & ~n_1775) ;
	assign n_1768 = (~x_701 & n_1766) ;
	assign n_1767 = (x_701 & ~n_1766) ;
	assign n_1759 = (~n_1756 & n_1758) ;
	assign n_1751 = (~n_1748 & n_1750) ;
	assign n_1747 = (~x_703 & ~n_665) ;
	assign n_1741 = (~x_704 & ~n_936) ;
	assign n_8279 = (~n_1776 & n_8278) ;
	assign n_1769 = (~n_1767 & ~n_1768) ;
	assign n_1761 = (~x_702 & ~n_1759) ;
	assign n_1760 = (x_702 & n_1759) ;
	assign n_1752 = (~n_1747 & n_1751) ;
	assign n_1742 = (i_5 & ~n_1741) ;
	assign n_1740 = (~i_63 & n_936) ;
	assign n_1734 = (i_62 & n_64) ;
	assign n_8280 = (~n_1769 & n_8279) ;
	assign n_1762 = (~n_1760 & ~n_1761) ;
	assign n_1754 = (~x_703 & ~n_1752) ;
	assign n_1753 = (x_703 & n_1752) ;
	assign n_1743 = (~n_1740 & n_1742) ;
	assign n_1735 = (n_66 & n_1734) ;
	assign n_1733 = (x_705 & n_978) ;
	assign n_8281 = (~n_1762 & n_8280) ;
	assign n_1755 = (~n_1753 & ~n_1754) ;
	assign n_1745 = (~x_704 & ~n_1743) ;
	assign n_1744 = (x_704 & n_1743) ;
	assign n_1736 = (~n_1733 & ~n_1735) ;
	assign n_8282 = (~n_1755 & n_8281) ;
	assign n_1746 = (~n_1744 & ~n_1745) ;
	assign n_1738 = (~x_705 & n_1736) ;
	assign n_1737 = (x_705 & ~n_1736) ;
	assign n_1725 = (x_526 & n_53) ;
	assign n_1724 = (x_707 & n_51) ;
	assign n_1718 = (~x_708 & ~n_630) ;
	assign n_8283 = (~n_1746 & n_8282) ;
	assign n_1739 = (~n_1737 & ~n_1738) ;
	assign n_1731 = (~x_706 & n_139) ;
	assign n_1730 = (x_706 & ~n_139) ;
	assign n_1726 = (~n_1724 & ~n_1725) ;
	assign n_1719 = (i_5 & ~n_1718) ;
	assign n_1717 = (~i_10 & n_630) ;
	assign n_1711 = (~x_709 & ~n_697) ;
	assign n_8284 = (~n_1739 & n_8283) ;
	assign n_1732 = (~n_1730 & ~n_1731) ;
	assign n_1728 = (~x_707 & n_1726) ;
	assign n_1727 = (x_707 & ~n_1726) ;
	assign n_1720 = (~n_1717 & n_1719) ;
	assign n_1712 = (i_5 & ~n_1711) ;
	assign n_1710 = (~x_201 & n_697) ;
	assign n_1704 = (i_6 & n_64) ;
	assign n_8285 = (~n_1732 & n_8284) ;
	assign n_1729 = (~n_1727 & ~n_1728) ;
	assign n_1722 = (~x_708 & ~n_1720) ;
	assign n_1721 = (x_708 & n_1720) ;
	assign n_1713 = (~n_1710 & n_1712) ;
	assign n_1705 = (n_66 & n_1704) ;
	assign n_1703 = (x_710 & n_978) ;
	assign n_1697 = (~x_711 & ~n_936) ;
	assign n_8286 = (~n_1729 & n_8285) ;
	assign n_1723 = (~n_1721 & ~n_1722) ;
	assign n_1715 = (~x_709 & ~n_1713) ;
	assign n_1714 = (x_709 & n_1713) ;
	assign n_1706 = (~n_1703 & ~n_1705) ;
	assign n_1698 = (i_5 & ~n_1697) ;
	assign n_1696 = (~i_20 & n_936) ;
	assign n_8287 = (~n_1723 & n_8286) ;
	assign n_1716 = (~n_1714 & ~n_1715) ;
	assign n_1708 = (~x_710 & n_1706) ;
	assign n_1707 = (x_710 & ~n_1706) ;
	assign n_1699 = (~n_1696 & n_1698) ;
	assign n_1691 = (~n_376 & n_1009) ;
	assign n_1690 = (x_712 & n_1007) ;
	assign n_8288 = (~n_1716 & n_8287) ;
	assign n_1709 = (~n_1707 & ~n_1708) ;
	assign n_1701 = (~x_711 & ~n_1699) ;
	assign n_1700 = (x_711 & n_1699) ;
	assign n_1692 = (~n_1690 & ~n_1691) ;
	assign n_1685 = (i_23 & n_948) ;
	assign n_1684 = (x_713 & n_945) ;
	assign n_1553 = (i_56 & n_64) ;
	assign n_8289 = (~n_1709 & n_8288) ;
	assign n_1702 = (~n_1700 & ~n_1701) ;
	assign n_1694 = (~x_712 & n_1692) ;
	assign n_1693 = (x_712 & ~n_1692) ;
	assign n_1686 = (~n_1684 & ~n_1685) ;
	assign n_1554 = (n_66 & n_1553) ;
	assign n_1552 = (x_714 & n_978) ;
	assign n_1675 = (~x_715 & ~n_936) ;
	assign n_8290 = (~n_1702 & n_8289) ;
	assign n_1695 = (~n_1693 & ~n_1694) ;
	assign n_1688 = (~x_713 & n_1686) ;
	assign n_1687 = (x_713 & ~n_1686) ;
	assign n_1555 = (~n_1552 & ~n_1554) ;
	assign n_1676 = (i_5 & ~n_1675) ;
	assign n_1674 = (~i_11 & n_936) ;
	assign n_1668 = (i_43 & n_64) ;
	assign n_8291 = (~n_1695 & n_8290) ;
	assign n_1689 = (~n_1687 & ~n_1688) ;
	assign n_1682 = (~x_714 & n_1555) ;
	assign n_1681 = (x_714 & ~n_1555) ;
	assign n_1677 = (~n_1674 & n_1676) ;
	assign n_1669 = (n_66 & n_1668) ;
	assign n_1667 = (x_716 & n_978) ;
	assign n_1661 = (~x_717 & ~n_697) ;
	assign n_1651 = (~n_663 & ~n_1650) ;
	assign n_8292 = (~n_1689 & n_8291) ;
	assign n_1683 = (~n_1681 & ~n_1682) ;
	assign n_1679 = (~x_715 & ~n_1677) ;
	assign n_1678 = (x_715 & n_1677) ;
	assign n_1670 = (~n_1667 & ~n_1669) ;
	assign n_1662 = (i_5 & ~n_1661) ;
	assign n_1660 = (~x_458 & n_697) ;
	assign n_1654 = (~n_936 & ~n_1653) ;
	assign n_1652 = (x_718 & ~n_1651) ;
	assign n_1595 = (~n_388 & ~n_389) ;
	assign n_8293 = (~n_1683 & n_8292) ;
	assign n_1680 = (~n_1678 & ~n_1679) ;
	assign n_1672 = (~x_716 & n_1670) ;
	assign n_1671 = (x_716 & ~n_1670) ;
	assign n_1663 = (~n_1660 & n_1662) ;
	assign n_1655 = (~n_1652 & n_1654) ;
	assign n_1644 = (~x_719 & ~n_630) ;
	assign n_1597 = (~x_754 & ~n_1595) ;
	assign n_8294 = (~n_1680 & n_8293) ;
	assign n_1673 = (~n_1671 & ~n_1672) ;
	assign n_1665 = (~x_717 & ~n_1663) ;
	assign n_1664 = (x_717 & n_1663) ;
	assign n_1656 = (i_5 & ~n_1655) ;
	assign n_1645 = (i_5 & ~n_1644) ;
	assign n_1643 = (~i_13 & n_630) ;
	assign n_1637 = (~x_720 & ~n_630) ;
	assign n_1598 = (~x_332 & ~n_1597) ;
	assign n_1596 = (x_754 & n_1595) ;
	assign n_8295 = (~n_1673 & n_8294) ;
	assign n_1666 = (~n_1664 & ~n_1665) ;
	assign n_1658 = (~x_718 & ~n_1656) ;
	assign n_1657 = (x_718 & n_1656) ;
	assign n_1646 = (~n_1643 & n_1645) ;
	assign n_1638 = (i_5 & ~n_1637) ;
	assign n_1636 = (~i_4 & n_630) ;
	assign n_1623 = (~i_16 & n_669) ;
	assign n_1621 = (~x_416 & ~n_544) ;
	assign n_1599 = (~n_1596 & n_1598) ;
	assign n_8296 = (~n_1666 & n_8295) ;
	assign n_1659 = (~n_1657 & ~n_1658) ;
	assign n_1648 = (~x_719 & ~n_1646) ;
	assign n_1647 = (x_719 & n_1646) ;
	assign n_1639 = (~n_1636 & n_1638) ;
	assign n_1631 = (~n_257 & n_35) ;
	assign n_1630 = (x_721 & n_36) ;
	assign n_1624 = (i_5 & ~n_1623) ;
	assign n_1622 = (n_662 & n_1621) ;
	assign n_1601 = (n_392 & ~n_1599) ;
	assign n_8297 = (~n_1659 & n_8296) ;
	assign n_1649 = (~n_1647 & ~n_1648) ;
	assign n_1641 = (~x_720 & ~n_1639) ;
	assign n_1640 = (x_720 & n_1639) ;
	assign n_1632 = (~n_1630 & ~n_1631) ;
	assign n_1625 = (~n_1622 & n_1624) ;
	assign n_1620 = (~x_722 & ~n_665) ;
	assign n_1607 = (~n_1606 & ~n_392) ;
	assign n_1604 = (i_4 & n_7) ;
	assign n_1602 = (x_664 & ~n_1601) ;
	assign n_1600 = (~n_392 & n_1599) ;
	assign n_8298 = (~n_1649 & n_8297) ;
	assign n_1642 = (~n_1640 & ~n_1641) ;
	assign n_1634 = (~x_721 & n_1632) ;
	assign n_1633 = (x_721 & ~n_1632) ;
	assign n_1626 = (~n_1620 & n_1625) ;
	assign n_1615 = (x_90 & n_35) ;
	assign n_1614 = (x_723 & n_36) ;
	assign n_1608 = (~n_1604 & ~n_1607) ;
	assign n_1603 = (~n_1600 & n_1602) ;
	assign n_8299 = (~n_1642 & n_8298) ;
	assign n_1635 = (~n_1633 & ~n_1634) ;
	assign n_1628 = (~x_722 & ~n_1626) ;
	assign n_1627 = (x_722 & n_1626) ;
	assign n_1616 = (~n_1614 & ~n_1615) ;
	assign n_1609 = (~n_1603 & n_1608) ;
	assign n_1585 = (~n_1584 & n_1551) ;
	assign n_1573 = (~n_1572 & n_1551) ;
	assign n_8300 = (~n_1635 & n_8299) ;
	assign n_1629 = (~n_1627 & ~n_1628) ;
	assign n_1618 = (~x_723 & n_1616) ;
	assign n_1617 = (x_723 & ~n_1616) ;
	assign n_1610 = (i_5 & ~n_1609) ;
	assign n_1586 = (~n_1568 & ~n_1585) ;
	assign n_1580 = (~n_1551 & ~n_1579) ;
	assign n_1574 = (n_1568 & ~n_1573) ;
	assign n_1556 = (~n_1551 & ~n_1555) ;
	assign n_8301 = (~n_1629 & n_8300) ;
	assign n_1619 = (~n_1617 & ~n_1618) ;
	assign n_1612 = (~x_724 & ~n_1610) ;
	assign n_1611 = (x_724 & n_1610) ;
	assign n_1587 = (~n_1580 & n_1586) ;
	assign n_1575 = (~n_1556 & n_1574) ;
	assign n_1531 = (~x_727 & ~n_936) ;
	assign n_1523 = (~i_12 & n_669) ;
	assign n_1521 = (~x_539 & ~n_544) ;
	assign n_8302 = (~n_1619 & n_8301) ;
	assign n_1613 = (~n_1611 & ~n_1612) ;
	assign n_1593 = (~x_725 & n_188) ;
	assign n_1592 = (x_725 & ~n_188) ;
	assign n_1588 = (~n_1575 & ~n_1587) ;
	assign n_1532 = (i_5 & ~n_1531) ;
	assign n_1530 = (~i_34 & n_936) ;
	assign n_1524 = (i_5 & ~n_1523) ;
	assign n_1522 = (n_662 & n_1521) ;
	assign n_8303 = (~n_1613 & n_8302) ;
	assign n_1594 = (~n_1592 & ~n_1593) ;
	assign n_1590 = (~x_726 & ~n_1588) ;
	assign n_1589 = (x_726 & n_1588) ;
	assign n_1533 = (~n_1530 & n_1532) ;
	assign n_1525 = (~n_1522 & n_1524) ;
	assign n_1520 = (~x_728 & ~n_665) ;
	assign n_8304 = (~n_1594 & n_8303) ;
	assign n_1591 = (~n_1589 & ~n_1590) ;
	assign n_1535 = (~x_727 & ~n_1533) ;
	assign n_1534 = (x_727 & n_1533) ;
	assign n_1526 = (~n_1520 & n_1525) ;
	assign n_1515 = (~n_179 & n_35) ;
	assign n_1514 = (x_729 & n_36) ;
	assign n_1508 = (~x_730 & ~n_630) ;
	assign n_8305 = (~n_1591 & n_8304) ;
	assign n_1536 = (~n_1534 & ~n_1535) ;
	assign n_1528 = (~x_728 & ~n_1526) ;
	assign n_1527 = (x_728 & n_1526) ;
	assign n_1516 = (~n_1514 & ~n_1515) ;
	assign n_1509 = (i_5 & ~n_1508) ;
	assign n_1507 = (~i_43 & n_630) ;
	assign n_8306 = (~n_1536 & n_8305) ;
	assign n_1529 = (~n_1527 & ~n_1528) ;
	assign n_1518 = (~x_729 & n_1516) ;
	assign n_1517 = (x_729 & ~n_1516) ;
	assign n_1510 = (~n_1507 & n_1509) ;
	assign n_8307 = (~n_1529 & n_8306) ;
	assign n_1519 = (~n_1517 & ~n_1518) ;
	assign n_1512 = (~x_730 & ~n_1510) ;
	assign n_1511 = (x_730 & n_1510) ;
	assign n_1499 = (n_35 & ~n_392) ;
	assign n_1498 = (x_732 & n_36) ;
	assign n_1477 = (i_50 & n_1) ;
	assign n_1476 = (~x_735 & n_6) ;
	assign n_1443 = (~x_655 & n_877) ;
	assign n_1442 = (x_655 & ~n_877) ;
	assign n_8308 = (~n_1519 & n_8307) ;
	assign n_1513 = (~n_1511 & ~n_1512) ;
	assign n_1505 = (~x_731 & n_317) ;
	assign n_1504 = (x_731 & ~n_317) ;
	assign n_1500 = (~n_1498 & ~n_1499) ;
	assign n_1493 = (x_737 & n_35) ;
	assign n_1492 = (x_733 & n_36) ;
	assign n_1486 = (i_4 & n_64) ;
	assign n_1478 = (~n_1476 & n_1477) ;
	assign n_1475 = (x_90 & ~n_16) ;
	assign n_1444 = (~n_1442 & ~n_1443) ;
	assign n_1441 = (~n_867 & ~n_868) ;
	assign n_8309 = (~n_1513 & n_8308) ;
	assign n_1506 = (~n_1504 & ~n_1505) ;
	assign n_1502 = (~x_732 & n_1500) ;
	assign n_1501 = (x_732 & ~n_1500) ;
	assign n_1494 = (~n_1492 & ~n_1493) ;
	assign n_1487 = (n_66 & n_1486) ;
	assign n_1485 = (x_734 & n_978) ;
	assign n_1479 = (~n_1475 & ~n_1478) ;
	assign n_1474 = (x_735 & n_17) ;
	assign n_1453 = (i_26 & ~n_6) ;
	assign n_1446 = (n_1441 & ~n_1444) ;
	assign n_8310 = (~n_1506 & n_8309) ;
	assign n_1503 = (~n_1501 & ~n_1502) ;
	assign n_1496 = (~x_733 & n_1494) ;
	assign n_1495 = (x_733 & ~n_1494) ;
	assign n_1488 = (~n_1485 & ~n_1487) ;
	assign n_1480 = (~n_1474 & n_1479) ;
	assign n_1454 = (n_629 & ~n_1453) ;
	assign n_1452 = (x_738 & n_6) ;
	assign n_1449 = (x_738 & ~n_697) ;
	assign n_1447 = (n_697 & ~n_1446) ;
	assign n_1445 = (~n_1441 & n_1444) ;
	assign n_8311 = (~n_1503 & n_8310) ;
	assign n_1497 = (~n_1495 & ~n_1496) ;
	assign n_1490 = (~x_734 & n_1488) ;
	assign n_1489 = (x_734 & ~n_1488) ;
	assign n_1481 = (i_5 & ~n_1480) ;
	assign n_1469 = (i_32 & n_948) ;
	assign n_1468 = (x_736 & n_945) ;
	assign n_1455 = (~n_1452 & n_1454) ;
	assign n_1450 = (~n_629 & ~n_1449) ;
	assign n_1448 = (~n_1445 & n_1447) ;
	assign n_8312 = (~n_1497 & n_8311) ;
	assign n_1491 = (~n_1489 & ~n_1490) ;
	assign n_1483 = (~x_735 & ~n_1481) ;
	assign n_1482 = (x_735 & n_1481) ;
	assign n_1470 = (~n_1468 & ~n_1469) ;
	assign n_1463 = (~n_347 & n_1009) ;
	assign n_1462 = (x_737 & n_1007) ;
	assign n_1456 = (n_902 & ~n_1455) ;
	assign n_1451 = (~n_1448 & n_1450) ;
	assign n_8313 = (~n_1491 & n_8312) ;
	assign n_1484 = (~n_1482 & ~n_1483) ;
	assign n_1472 = (~x_736 & n_1470) ;
	assign n_1471 = (x_736 & ~n_1470) ;
	assign n_1464 = (~n_1462 & ~n_1463) ;
	assign n_1457 = (~n_1451 & n_1456) ;
	assign n_1440 = (x_738 & n_699) ;
	assign n_8314 = (~n_1484 & n_8313) ;
	assign n_1473 = (~n_1471 & ~n_1472) ;
	assign n_1466 = (~x_737 & n_1464) ;
	assign n_1465 = (x_737 & ~n_1464) ;
	assign n_1458 = (~n_1440 & ~n_1457) ;
	assign n_1435 = (x_220 & n_53) ;
	assign n_1434 = (x_739 & n_51) ;
	assign n_1428 = (i_61 & n_59) ;
	assign n_8315 = (~n_1473 & n_8314) ;
	assign n_1467 = (~n_1465 & ~n_1466) ;
	assign n_1460 = (~x_738 & n_1458) ;
	assign n_1459 = (x_738 & ~n_1458) ;
	assign n_1436 = (~n_1434 & ~n_1435) ;
	assign n_1429 = (n_66 & n_1428) ;
	assign n_1427 = (x_740 & n_60) ;
	assign n_1421 = (i_55 & n_59) ;
	assign n_8316 = (~n_1467 & n_8315) ;
	assign n_1461 = (~n_1459 & ~n_1460) ;
	assign n_1438 = (~x_739 & n_1436) ;
	assign n_1437 = (x_739 & ~n_1436) ;
	assign n_1430 = (~n_1427 & ~n_1429) ;
	assign n_1422 = (n_66 & n_1421) ;
	assign n_1420 = (x_741 & n_60) ;
	assign n_1414 = (i_48 & n_64) ;
	assign n_8317 = (~n_1461 & n_8316) ;
	assign n_1439 = (~n_1437 & ~n_1438) ;
	assign n_1432 = (~x_740 & n_1430) ;
	assign n_1431 = (x_740 & ~n_1430) ;
	assign n_1423 = (~n_1420 & ~n_1422) ;
	assign n_1415 = (n_66 & n_1414) ;
	assign n_1413 = (x_742 & n_978) ;
	assign n_8318 = (~n_1439 & n_8317) ;
	assign n_1433 = (~n_1431 & ~n_1432) ;
	assign n_1425 = (~x_741 & n_1423) ;
	assign n_1424 = (x_741 & ~n_1423) ;
	assign n_1416 = (~n_1413 & ~n_1415) ;
	assign n_1408 = (i_44 & n_948) ;
	assign n_1407 = (x_743 & n_945) ;
	assign n_1401 = (~x_744 & ~n_630) ;
	assign n_8319 = (~n_1433 & n_8318) ;
	assign n_1426 = (~n_1424 & ~n_1425) ;
	assign n_1418 = (~x_742 & n_1416) ;
	assign n_1417 = (x_742 & ~n_1416) ;
	assign n_1409 = (~n_1407 & ~n_1408) ;
	assign n_1402 = (i_5 & ~n_1401) ;
	assign n_1400 = (~i_50 & n_630) ;
	assign n_8320 = (~n_1426 & n_8319) ;
	assign n_1419 = (~n_1417 & ~n_1418) ;
	assign n_1411 = (~x_743 & n_1409) ;
	assign n_1410 = (x_743 & ~n_1409) ;
	assign n_1403 = (~n_1400 & n_1402) ;
	assign n_1395 = (x_247 & n_53) ;
	assign n_1394 = (x_745 & n_51) ;
	assign n_8321 = (~n_1419 & n_8320) ;
	assign n_1412 = (~n_1410 & ~n_1411) ;
	assign n_1405 = (~x_744 & ~n_1403) ;
	assign n_1404 = (x_744 & n_1403) ;
	assign n_1396 = (~n_1394 & ~n_1395) ;
	assign n_1389 = (x_181 & n_35) ;
	assign n_1388 = (x_746 & n_36) ;
	assign n_8322 = (~n_1412 & n_8321) ;
	assign n_1406 = (~n_1404 & ~n_1405) ;
	assign n_1398 = (~x_745 & n_1396) ;
	assign n_1397 = (x_745 & ~n_1396) ;
	assign n_1390 = (~n_1388 & ~n_1389) ;
	assign n_1383 = (i_6 & n_948) ;
	assign n_1382 = (x_747 & n_945) ;
	assign n_1376 = (i_19 & n_59) ;
	assign n_8323 = (~n_1406 & n_8322) ;
	assign n_1399 = (~n_1397 & ~n_1398) ;
	assign n_1392 = (~x_746 & n_1390) ;
	assign n_1391 = (x_746 & ~n_1390) ;
	assign n_1384 = (~n_1382 & ~n_1383) ;
	assign n_1377 = (n_66 & n_1376) ;
	assign n_1375 = (x_748 & n_60) ;
	assign n_1369 = (~x_749 & ~n_544) ;
	assign n_8324 = (~n_1399 & n_8323) ;
	assign n_1393 = (~n_1391 & ~n_1392) ;
	assign n_1386 = (~x_747 & n_1384) ;
	assign n_1385 = (x_747 & ~n_1384) ;
	assign n_1378 = (~n_1375 & ~n_1377) ;
	assign n_1370 = (i_5 & ~n_1369) ;
	assign n_1368 = (~i_68 & n_544) ;
	assign n_8325 = (~n_1393 & n_8324) ;
	assign n_1387 = (~n_1385 & ~n_1386) ;
	assign n_1380 = (~x_748 & n_1378) ;
	assign n_1379 = (x_748 & ~n_1378) ;
	assign n_1371 = (~n_1368 & n_1370) ;
	assign n_1363 = (x_225 & n_53) ;
	assign n_1362 = (x_750 & n_51) ;
	assign n_1356 = (~x_751 & ~n_544) ;
	assign n_8326 = (~n_1387 & n_8325) ;
	assign n_1381 = (~n_1379 & ~n_1380) ;
	assign n_1373 = (~x_749 & ~n_1371) ;
	assign n_1372 = (x_749 & n_1371) ;
	assign n_1364 = (~n_1362 & ~n_1363) ;
	assign n_1357 = (i_5 & ~n_1356) ;
	assign n_1355 = (~i_34 & n_544) ;
	assign n_1349 = (i_9 & n_59) ;
	assign n_8327 = (~n_1381 & n_8326) ;
	assign n_1374 = (~n_1372 & ~n_1373) ;
	assign n_1366 = (~x_750 & n_1364) ;
	assign n_1365 = (x_750 & ~n_1364) ;
	assign n_1358 = (~n_1355 & n_1357) ;
	assign n_1350 = (n_66 & n_1349) ;
	assign n_1348 = (x_752 & n_60) ;
	assign n_1335 = (x_102 & ~n_16) ;
	assign n_1334 = (i_43 & n_7) ;
	assign n_1317 = (x_756 & ~n_14) ;
	assign n_8328 = (~n_1374 & n_8327) ;
	assign n_1367 = (~n_1365 & ~n_1366) ;
	assign n_1360 = (~x_751 & ~n_1358) ;
	assign n_1359 = (x_751 & n_1358) ;
	assign n_1351 = (~n_1348 & ~n_1350) ;
	assign n_1343 = (n_35 & ~n_497) ;
	assign n_1342 = (x_753 & n_36) ;
	assign n_1336 = (~n_1334 & ~n_1335) ;
	assign n_1318 = (n_12 & ~n_1317) ;
	assign n_1316 = (x_429 & n_14) ;
	assign n_1313 = (x_429 & n_11) ;
	assign n_8329 = (~n_1367 & n_8328) ;
	assign n_1361 = (~n_1359 & ~n_1360) ;
	assign n_1353 = (~x_752 & n_1351) ;
	assign n_1352 = (x_752 & ~n_1351) ;
	assign n_1344 = (~n_1342 & ~n_1343) ;
	assign n_1337 = (n_20 & ~n_1336) ;
	assign n_1333 = (x_754 & n_18) ;
	assign n_1327 = (~x_755 & ~n_544) ;
	assign n_1319 = (~n_1316 & n_1318) ;
	assign n_1314 = (x_168 & ~n_1313) ;
	assign n_1312 = (x_756 & ~n_11) ;
	assign n_1309 = (~x_756 & n_6) ;
	assign n_8330 = (~n_1361 & n_8329) ;
	assign n_1354 = (~n_1352 & ~n_1353) ;
	assign n_1346 = (~x_753 & n_1344) ;
	assign n_1345 = (x_753 & ~n_1344) ;
	assign n_1338 = (~n_1333 & ~n_1337) ;
	assign n_1328 = (i_5 & ~n_1327) ;
	assign n_1326 = (~i_61 & n_544) ;
	assign n_1320 = (i_5 & ~n_1319) ;
	assign n_1315 = (~n_1312 & n_1314) ;
	assign n_1310 = (~n_1308 & ~n_1309) ;
	assign n_8331 = (~n_1354 & n_8330) ;
	assign n_1347 = (~n_1345 & ~n_1346) ;
	assign n_1340 = (~x_754 & n_1338) ;
	assign n_1339 = (x_754 & ~n_1338) ;
	assign n_1329 = (~n_1326 & n_1328) ;
	assign n_1321 = (~n_1315 & n_1320) ;
	assign n_1311 = (n_1 & ~n_1310) ;
	assign n_8332 = (~n_1347 & n_8331) ;
	assign n_1341 = (~n_1339 & ~n_1340) ;
	assign n_1331 = (~x_755 & ~n_1329) ;
	assign n_1330 = (x_755 & n_1329) ;
	assign n_1322 = (~n_1311 & n_1321) ;
	assign n_1303 = (i_59 & n_948) ;
	assign n_1302 = (x_757 & n_945) ;
	assign n_1296 = (~x_758 & ~n_697) ;
	assign n_1288 = (i_7 & n_7) ;
	assign n_1287 = (x_328 & ~n_16) ;
	assign n_516 = (x_472 & ~x_578) ;
	assign n_515 = (~x_255 & x_478) ;
	assign n_8333 = (~n_1341 & n_8332) ;
	assign n_1332 = (~n_1330 & ~n_1331) ;
	assign n_1324 = (~x_756 & ~n_1322) ;
	assign n_1323 = (x_756 & n_1322) ;
	assign n_1304 = (~n_1302 & ~n_1303) ;
	assign n_1297 = (i_5 & ~n_1296) ;
	assign n_1295 = (~x_493 & n_697) ;
	assign n_1289 = (~n_1287 & ~n_1288) ;
	assign n_1214 = (x_395 & ~x_578) ;
	assign n_1213 = (~x_255 & x_561) ;
	assign n_520 = (x_214 & n_9) ;
	assign n_519 = (x_206 & n_13) ;
	assign n_517 = (~n_515 & ~n_516) ;
	assign n_8334 = (~n_1332 & n_8333) ;
	assign n_1325 = (~n_1323 & ~n_1324) ;
	assign n_1306 = (~x_757 & n_1304) ;
	assign n_1305 = (x_757 & ~n_1304) ;
	assign n_1298 = (~n_1295 & n_1297) ;
	assign n_1290 = (n_20 & ~n_1289) ;
	assign n_1286 = (x_759 & n_18) ;
	assign n_1280 = (~x_760 & ~n_544) ;
	assign n_1218 = (x_292 & n_9) ;
	assign n_1217 = (x_115 & n_13) ;
	assign n_1215 = (~n_1213 & ~n_1214) ;
	assign n_521 = (~n_519 & ~n_520) ;
	assign n_518 = (~n_9 & ~n_517) ;
	assign n_513 = (~n_511 & ~n_512) ;
	assign n_8335 = (~n_1325 & n_8334) ;
	assign n_1307 = (~n_1305 & ~n_1306) ;
	assign n_1300 = (~x_758 & ~n_1298) ;
	assign n_1299 = (x_758 & n_1298) ;
	assign n_1291 = (~n_1286 & ~n_1290) ;
	assign n_1281 = (i_5 & ~n_1280) ;
	assign n_1279 = (~i_46 & n_544) ;
	assign n_1225 = (~x_438 & n_1223) ;
	assign n_1224 = (x_438 & ~n_1223) ;
	assign n_1219 = (~n_1217 & ~n_1218) ;
	assign n_1216 = (~n_9 & ~n_1215) ;
	assign n_522 = (~n_518 & n_521) ;
	assign n_514 = (~n_508 & ~n_513) ;
	assign n_8336 = (~n_1307 & n_8335) ;
	assign n_1301 = (~n_1299 & ~n_1300) ;
	assign n_1293 = (~x_759 & n_1291) ;
	assign n_1292 = (x_759 & ~n_1291) ;
	assign n_1282 = (~n_1279 & n_1281) ;
	assign n_1274 = (x_465 & n_53) ;
	assign n_1273 = (x_761 & n_51) ;
	assign n_1267 = (i_57 & n_59) ;
	assign n_1226 = (~n_1224 & ~n_1225) ;
	assign n_1220 = (~n_1216 & n_1219) ;
	assign n_524 = (n_514 & n_522) ;
	assign n_8337 = (~n_1301 & n_8336) ;
	assign n_1294 = (~n_1292 & ~n_1293) ;
	assign n_1284 = (~x_760 & ~n_1282) ;
	assign n_1283 = (x_760 & n_1282) ;
	assign n_1275 = (~n_1273 & ~n_1274) ;
	assign n_1268 = (n_66 & n_1267) ;
	assign n_1266 = (x_762 & n_60) ;
	assign n_1228 = (~n_1220 & ~n_1226) ;
	assign n_1227 = (n_1220 & n_1226) ;
	assign n_1211 = (~n_75 & ~n_524) ;
	assign n_523 = (~n_514 & ~n_522) ;
	assign n_8338 = (~n_1294 & n_8337) ;
	assign n_1285 = (~n_1283 & ~n_1284) ;
	assign n_1277 = (~x_761 & n_1275) ;
	assign n_1276 = (x_761 & ~n_1275) ;
	assign n_1269 = (~n_1266 & ~n_1268) ;
	assign n_1229 = (~n_1227 & ~n_1228) ;
	assign n_1212 = (~n_523 & ~n_1211) ;
	assign n_8339 = (~n_1285 & n_8338) ;
	assign n_1278 = (~n_1276 & ~n_1277) ;
	assign n_1271 = (~x_762 & n_1269) ;
	assign n_1270 = (x_762 & ~n_1269) ;
	assign n_1254 = (~x_765 & ~n_936) ;
	assign n_1238 = (n_1 & ~n_1237) ;
	assign n_1236 = (n_6 & n_1223) ;
	assign n_1231 = (n_1212 & n_1229) ;
	assign n_8340 = (~n_1278 & n_8339) ;
	assign n_1272 = (~n_1270 & ~n_1271) ;
	assign n_1264 = (~x_763 & n_467) ;
	assign n_1263 = (x_763 & ~n_467) ;
	assign n_1255 = (i_5 & ~n_1254) ;
	assign n_1253 = (~i_17 & n_936) ;
	assign n_1247 = (~x_766 & ~n_544) ;
	assign n_1239 = (~n_1236 & n_1238) ;
	assign n_1235 = (~n_1223 & n_1234) ;
	assign n_1232 = (n_527 & ~n_1231) ;
	assign n_1230 = (~n_1212 & ~n_1229) ;
	assign n_8341 = (~n_1272 & n_8340) ;
	assign n_1265 = (~n_1263 & ~n_1264) ;
	assign n_1261 = (~x_764 & n_86) ;
	assign n_1260 = (x_764 & ~n_86) ;
	assign n_1256 = (~n_1253 & n_1255) ;
	assign n_1248 = (i_5 & ~n_1247) ;
	assign n_1246 = (~i_44 & n_544) ;
	assign n_1240 = (~n_1235 & ~n_1239) ;
	assign n_1233 = (~n_1230 & n_1232) ;
	assign n_8342 = (~n_1265 & n_8341) ;
	assign n_1262 = (~n_1260 & ~n_1261) ;
	assign n_1258 = (~x_765 & ~n_1256) ;
	assign n_1257 = (x_765 & n_1256) ;
	assign n_1249 = (~n_1246 & n_1248) ;
	assign n_1241 = (~n_1233 & n_1240) ;
	assign n_1205 = (~x_768 & ~n_630) ;
	assign n_8343 = (~n_1262 & n_8342) ;
	assign n_1259 = (~n_1257 & ~n_1258) ;
	assign n_1251 = (~x_766 & ~n_1249) ;
	assign n_1250 = (x_766 & n_1249) ;
	assign n_1242 = (i_5 & ~n_1241) ;
	assign n_1206 = (i_5 & ~n_1205) ;
	assign n_1204 = (~i_37 & n_630) ;
	assign n_8344 = (~n_1259 & n_8343) ;
	assign n_1252 = (~n_1250 & ~n_1251) ;
	assign n_1244 = (~x_767 & ~n_1242) ;
	assign n_1243 = (x_767 & n_1242) ;
	assign n_1207 = (~n_1204 & n_1206) ;
	assign n_1199 = (x_775 & n_53) ;
	assign n_1198 = (x_769 & n_51) ;
	assign n_1192 = (i_50 & n_64) ;
	assign n_1146 = (~x_249 & n_1144) ;
	assign n_1145 = (x_249 & ~n_1144) ;
	assign n_8345 = (~n_1252 & n_8344) ;
	assign n_1245 = (~n_1243 & ~n_1244) ;
	assign n_1209 = (~x_768 & ~n_1207) ;
	assign n_1208 = (x_768 & n_1207) ;
	assign n_1200 = (~n_1198 & ~n_1199) ;
	assign n_1193 = (n_66 & n_1192) ;
	assign n_1191 = (x_770 & n_978) ;
	assign n_1147 = (~n_1145 & ~n_1146) ;
	assign n_1135 = (~n_1133 & ~n_1134) ;
	assign n_8346 = (~n_1245 & n_8345) ;
	assign n_1210 = (~n_1208 & ~n_1209) ;
	assign n_1202 = (~x_769 & n_1200) ;
	assign n_1201 = (x_769 & ~n_1200) ;
	assign n_1194 = (~n_1191 & ~n_1193) ;
	assign n_1186 = (i_65 & n_948) ;
	assign n_1185 = (x_771 & n_945) ;
	assign n_1156 = (~x_775 & n_6) ;
	assign n_1149 = (n_1135 & ~n_1147) ;
	assign n_8347 = (~n_1210 & n_8346) ;
	assign n_1203 = (~n_1201 & ~n_1202) ;
	assign n_1196 = (~x_770 & n_1194) ;
	assign n_1195 = (x_770 & ~n_1194) ;
	assign n_1187 = (~n_1185 & ~n_1186) ;
	assign n_1180 = (i_22 & n_948) ;
	assign n_1179 = (x_772 & n_945) ;
	assign n_1173 = (~x_773 & ~n_697) ;
	assign n_1157 = (~n_1155 & ~n_1156) ;
	assign n_1152 = (x_775 & ~n_697) ;
	assign n_1150 = (n_697 & ~n_1149) ;
	assign n_1148 = (~n_1135 & n_1147) ;
	assign n_8348 = (~n_1203 & n_8347) ;
	assign n_1197 = (~n_1195 & ~n_1196) ;
	assign n_1189 = (~x_771 & n_1187) ;
	assign n_1188 = (x_771 & ~n_1187) ;
	assign n_1181 = (~n_1179 & ~n_1180) ;
	assign n_1174 = (i_5 & ~n_1173) ;
	assign n_1172 = (~x_216 & n_697) ;
	assign n_1166 = (i_46 & n_59) ;
	assign n_1158 = (n_629 & ~n_1157) ;
	assign n_1153 = (~n_629 & ~n_1152) ;
	assign n_1151 = (~n_1148 & n_1150) ;
	assign n_8349 = (~n_1197 & n_8348) ;
	assign n_1190 = (~n_1188 & ~n_1189) ;
	assign n_1183 = (~x_772 & n_1181) ;
	assign n_1182 = (x_772 & ~n_1181) ;
	assign n_1175 = (~n_1172 & n_1174) ;
	assign n_1167 = (n_66 & n_1166) ;
	assign n_1165 = (x_774 & n_60) ;
	assign n_1159 = (n_902 & ~n_1158) ;
	assign n_1154 = (~n_1151 & n_1153) ;
	assign n_8350 = (~n_1190 & n_8349) ;
	assign n_1184 = (~n_1182 & ~n_1183) ;
	assign n_1177 = (~x_773 & ~n_1175) ;
	assign n_1176 = (x_773 & n_1175) ;
	assign n_1168 = (~n_1165 & ~n_1167) ;
	assign n_1160 = (~n_1154 & n_1159) ;
	assign n_1130 = (x_775 & n_699) ;
	assign n_1124 = (i_58 & n_59) ;
	assign n_8351 = (~n_1184 & n_8350) ;
	assign n_1178 = (~n_1176 & ~n_1177) ;
	assign n_1170 = (~x_774 & n_1168) ;
	assign n_1169 = (x_774 & ~n_1168) ;
	assign n_1161 = (~n_1130 & ~n_1160) ;
	assign n_1125 = (n_66 & n_1124) ;
	assign n_1123 = (x_776 & n_60) ;
	assign n_8352 = (~n_1178 & n_8351) ;
	assign n_1171 = (~n_1169 & ~n_1170) ;
	assign n_1163 = (~x_775 & n_1161) ;
	assign n_1162 = (x_775 & ~n_1161) ;
	assign n_1126 = (~n_1123 & ~n_1125) ;
	assign n_1112 = (~x_778 & ~n_936) ;
	assign n_1054 = (~n_403 & ~n_404) ;
	assign n_8353 = (~n_1171 & n_8352) ;
	assign n_1164 = (~n_1162 & ~n_1163) ;
	assign n_1128 = (~x_776 & n_1126) ;
	assign n_1127 = (x_776 & ~n_1126) ;
	assign n_1119 = (n_51 & ~n_1118) ;
	assign n_1113 = (i_5 & ~n_1112) ;
	assign n_1111 = (~i_67 & n_936) ;
	assign n_1056 = (~x_671 & ~n_1054) ;
	assign n_8354 = (~n_1164 & n_8353) ;
	assign n_1129 = (~n_1127 & ~n_1128) ;
	assign n_1121 = (~x_777 & ~n_1119) ;
	assign n_1120 = (x_777 & n_1119) ;
	assign n_1114 = (~n_1111 & n_1113) ;
	assign n_1106 = (~n_317 & n_1009) ;
	assign n_1105 = (x_779 & n_1007) ;
	assign n_1099 = (i_35 & n_64) ;
	assign n_1083 = (i_48 & n_1) ;
	assign n_1082 = (~x_782 & n_6) ;
	assign n_1057 = (~x_332 & ~n_1056) ;
	assign n_1055 = (x_671 & n_1054) ;
	assign n_8355 = (~n_1129 & n_8354) ;
	assign n_1122 = (~n_1120 & ~n_1121) ;
	assign n_1116 = (~x_778 & ~n_1114) ;
	assign n_1115 = (x_778 & n_1114) ;
	assign n_1107 = (~n_1105 & ~n_1106) ;
	assign n_1100 = (n_66 & n_1099) ;
	assign n_1098 = (x_780 & n_978) ;
	assign n_1092 = (~x_781 & ~n_544) ;
	assign n_1084 = (~n_1082 & n_1083) ;
	assign n_1081 = (x_656 & ~n_16) ;
	assign n_1058 = (~n_1055 & n_1057) ;
	assign n_8356 = (~n_1122 & n_8355) ;
	assign n_1117 = (~n_1115 & ~n_1116) ;
	assign n_1109 = (~x_779 & n_1107) ;
	assign n_1108 = (x_779 & ~n_1107) ;
	assign n_1101 = (~n_1098 & ~n_1100) ;
	assign n_1093 = (i_5 & ~n_1092) ;
	assign n_1091 = (~i_11 & n_544) ;
	assign n_1085 = (~n_1081 & ~n_1084) ;
	assign n_1080 = (x_782 & n_17) ;
	assign n_1066 = (n_1 & ~n_1065) ;
	assign n_1064 = (n_6 & n_407) ;
	assign n_1060 = (n_407 & ~n_1058) ;
	assign n_8357 = (~n_1117 & n_8356) ;
	assign n_1110 = (~n_1108 & ~n_1109) ;
	assign n_1103 = (~x_780 & n_1101) ;
	assign n_1102 = (x_780 & ~n_1101) ;
	assign n_1094 = (~n_1091 & n_1093) ;
	assign n_1086 = (~n_1080 & n_1085) ;
	assign n_1067 = (~n_1064 & n_1066) ;
	assign n_1063 = (n_59 & ~n_407) ;
	assign n_1061 = (x_664 & ~n_1060) ;
	assign n_1059 = (~n_407 & n_1058) ;
	assign n_8358 = (~n_1110 & n_8357) ;
	assign n_1104 = (~n_1102 & ~n_1103) ;
	assign n_1096 = (~x_781 & ~n_1094) ;
	assign n_1095 = (x_781 & n_1094) ;
	assign n_1087 = (i_5 & ~n_1086) ;
	assign n_1075 = (x_110 & n_53) ;
	assign n_1074 = (x_783 & n_51) ;
	assign n_1068 = (~n_1063 & ~n_1067) ;
	assign n_1062 = (~n_1059 & n_1061) ;
	assign n_8359 = (~n_1104 & n_8358) ;
	assign n_1097 = (~n_1095 & ~n_1096) ;
	assign n_1089 = (~x_782 & ~n_1087) ;
	assign n_1088 = (x_782 & n_1087) ;
	assign n_1076 = (~n_1074 & ~n_1075) ;
	assign n_1069 = (~n_1062 & n_1068) ;
	assign n_8360 = (~n_1097 & n_8359) ;
	assign n_1090 = (~n_1088 & ~n_1089) ;
	assign n_1078 = (~x_783 & n_1076) ;
	assign n_1077 = (x_783 & ~n_1076) ;
	assign n_1070 = (i_5 & ~n_1069) ;
	assign n_1045 = (i_41 & n_64) ;
	assign n_8361 = (~n_1090 & n_8360) ;
	assign n_1079 = (~n_1077 & ~n_1078) ;
	assign n_1072 = (~x_784 & ~n_1070) ;
	assign n_1071 = (x_784 & n_1070) ;
	assign n_1046 = (n_66 & n_1045) ;
	assign n_1044 = (x_786 & n_978) ;
	assign n_8362 = (~n_1079 & n_8361) ;
	assign n_1073 = (~n_1071 & ~n_1072) ;
	assign n_1052 = (~x_785 & n_203) ;
	assign n_1051 = (x_785 & ~n_203) ;
	assign n_1047 = (~n_1044 & ~n_1046) ;
	assign n_8363 = (~n_1073 & n_8362) ;
	assign n_1053 = (~n_1051 & ~n_1052) ;
	assign n_1049 = (~x_786 & n_1047) ;
	assign n_1048 = (x_786 & ~n_1047) ;
	assign n_1036 = (~n_136 & n_35) ;
	assign n_1035 = (x_788 & n_36) ;
	assign n_8364 = (~n_1053 & n_8363) ;
	assign n_1050 = (~n_1048 & ~n_1049) ;
	assign n_1042 = (~x_787 & n_332) ;
	assign n_1041 = (x_787 & ~n_332) ;
	assign n_1037 = (~n_1035 & ~n_1036) ;
	assign n_1030 = (x_320 & n_53) ;
	assign n_1029 = (x_789 & n_51) ;
	assign n_1023 = (~x_790 & ~n_630) ;
	assign n_8365 = (~n_1050 & n_8364) ;
	assign n_1043 = (~n_1041 & ~n_1042) ;
	assign n_1039 = (~x_788 & n_1037) ;
	assign n_1038 = (x_788 & ~n_1037) ;
	assign n_1031 = (~n_1029 & ~n_1030) ;
	assign n_1024 = (i_5 & ~n_1023) ;
	assign n_1022 = (~i_17 & n_630) ;
	assign n_1016 = (~x_791 & ~n_630) ;
	assign n_8366 = (~n_1043 & n_8365) ;
	assign n_1040 = (~n_1038 & ~n_1039) ;
	assign n_1033 = (~x_789 & n_1031) ;
	assign n_1032 = (x_789 & ~n_1031) ;
	assign n_1025 = (~n_1022 & n_1024) ;
	assign n_1017 = (i_5 & ~n_1016) ;
	assign n_1015 = (~i_35 & n_630) ;
	assign n_8367 = (~n_1040 & n_8366) ;
	assign n_1034 = (~n_1032 & ~n_1033) ;
	assign n_1027 = (~x_790 & ~n_1025) ;
	assign n_1026 = (x_790 & n_1025) ;
	assign n_1018 = (~n_1015 & n_1017) ;
	assign n_1010 = (~n_302 & n_1009) ;
	assign n_1008 = (x_792 & n_1007) ;
	assign n_1001 = (~x_793 & ~n_697) ;
	assign n_8368 = (~n_1034 & n_8367) ;
	assign n_1028 = (~n_1026 & ~n_1027) ;
	assign n_1020 = (~x_791 & ~n_1018) ;
	assign n_1019 = (x_791 & n_1018) ;
	assign n_1011 = (~n_1008 & ~n_1010) ;
	assign n_1002 = (i_5 & ~n_1001) ;
	assign n_1000 = (~x_299 & n_697) ;
	assign n_994 = (~x_794 & ~n_936) ;
	assign n_8369 = (~n_1028 & n_8368) ;
	assign n_1021 = (~n_1019 & ~n_1020) ;
	assign n_1013 = (~x_792 & n_1011) ;
	assign n_1012 = (x_792 & ~n_1011) ;
	assign n_1003 = (~n_1000 & n_1002) ;
	assign n_995 = (i_5 & ~n_994) ;
	assign n_993 = (~i_12 & n_936) ;
	assign n_987 = (~x_795 & ~n_936) ;
	assign n_8370 = (~n_1021 & n_8369) ;
	assign n_1014 = (~n_1012 & ~n_1013) ;
	assign n_1005 = (~x_793 & ~n_1003) ;
	assign n_1004 = (x_793 & n_1003) ;
	assign n_996 = (~n_993 & n_995) ;
	assign n_988 = (i_5 & ~n_987) ;
	assign n_986 = (~i_66 & n_936) ;
	assign n_980 = (i_65 & n_64) ;
	assign n_8371 = (~n_1014 & n_8370) ;
	assign n_1006 = (~n_1004 & ~n_1005) ;
	assign n_998 = (~x_794 & ~n_996) ;
	assign n_997 = (x_794 & n_996) ;
	assign n_989 = (~n_986 & n_988) ;
	assign n_981 = (n_66 & n_980) ;
	assign n_979 = (x_796 & n_978) ;
	assign n_8372 = (~n_1006 & n_8371) ;
	assign n_999 = (~n_997 & ~n_998) ;
	assign n_991 = (~x_795 & ~n_989) ;
	assign n_990 = (x_795 & n_989) ;
	assign n_982 = (~n_979 & ~n_981) ;
	assign n_973 = (i_57 & n_948) ;
	assign n_972 = (x_797 & n_945) ;
	assign n_966 = (~x_798 & ~n_630) ;
	assign n_8373 = (~n_999 & n_8372) ;
	assign n_992 = (~n_990 & ~n_991) ;
	assign n_984 = (~x_796 & n_982) ;
	assign n_983 = (x_796 & ~n_982) ;
	assign n_974 = (~n_972 & ~n_973) ;
	assign n_967 = (i_5 & ~n_966) ;
	assign n_965 = (~i_62 & n_630) ;
	assign n_8374 = (~n_992 & n_8373) ;
	assign n_985 = (~n_983 & ~n_984) ;
	assign n_976 = (~x_797 & n_974) ;
	assign n_975 = (x_797 & ~n_974) ;
	assign n_968 = (~n_965 & n_967) ;
	assign n_960 = (~x_799 & ~n_629) ;
	assign n_8375 = (~n_985 & n_8374) ;
	assign n_977 = (~n_975 & ~n_976) ;
	assign n_970 = (~x_798 & ~n_968) ;
	assign n_969 = (x_798 & n_968) ;
	assign n_961 = (i_5 & ~n_960) ;
	assign n_955 = (x_557 & n_35) ;
	assign n_954 = (x_800 & n_36) ;
	assign n_893 = (~x_571 & n_891) ;
	assign n_892 = (x_571 & ~n_891) ;
	assign n_8376 = (~n_977 & n_8375) ;
	assign n_971 = (~n_969 & ~n_970) ;
	assign n_963 = (~x_799 & ~n_961) ;
	assign n_962 = (x_799 & n_961) ;
	assign n_956 = (~n_954 & ~n_955) ;
	assign n_949 = (i_45 & n_948) ;
	assign n_946 = (x_801 & n_945) ;
	assign n_938 = (~x_802 & ~n_936) ;
	assign n_929 = (i_25 & n_7) ;
	assign n_928 = (x_737 & ~n_16) ;
	assign n_894 = (~n_892 & ~n_893) ;
	assign n_882 = (~n_880 & ~n_881) ;
	assign n_8377 = (~n_971 & n_8376) ;
	assign n_964 = (~n_962 & ~n_963) ;
	assign n_958 = (~x_800 & n_956) ;
	assign n_957 = (x_800 & ~n_956) ;
	assign n_950 = (~n_946 & ~n_949) ;
	assign n_939 = (i_5 & ~n_938) ;
	assign n_937 = (~i_35 & n_936) ;
	assign n_930 = (~n_928 & ~n_929) ;
	assign n_904 = (~x_806 & n_6) ;
	assign n_896 = (n_882 & ~n_894) ;
	assign n_8378 = (~n_964 & n_8377) ;
	assign n_959 = (~n_957 & ~n_958) ;
	assign n_952 = (~x_801 & n_950) ;
	assign n_951 = (x_801 & ~n_950) ;
	assign n_940 = (~n_937 & n_939) ;
	assign n_931 = (n_20 & ~n_930) ;
	assign n_927 = (x_803 & n_18) ;
	assign n_921 = (~x_804 & ~n_544) ;
	assign n_905 = (~n_903 & ~n_904) ;
	assign n_899 = (x_806 & ~n_697) ;
	assign n_897 = (n_697 & ~n_896) ;
	assign n_895 = (~n_882 & n_894) ;
	assign n_8379 = (~n_959 & n_8378) ;
	assign n_953 = (~n_951 & ~n_952) ;
	assign n_942 = (~x_802 & ~n_940) ;
	assign n_941 = (x_802 & n_940) ;
	assign n_932 = (~n_927 & ~n_931) ;
	assign n_922 = (i_5 & ~n_921) ;
	assign n_920 = (~i_49 & n_544) ;
	assign n_914 = (i_30 & n_59) ;
	assign n_906 = (n_629 & ~n_905) ;
	assign n_900 = (~n_629 & ~n_899) ;
	assign n_898 = (~n_895 & n_897) ;
	assign n_8380 = (~n_953 & n_8379) ;
	assign n_943 = (~n_941 & ~n_942) ;
	assign n_934 = (~x_803 & n_932) ;
	assign n_933 = (x_803 & ~n_932) ;
	assign n_923 = (~n_920 & n_922) ;
	assign n_915 = (n_66 & n_914) ;
	assign n_913 = (x_805 & n_60) ;
	assign n_907 = (n_902 & ~n_906) ;
	assign n_901 = (~n_898 & n_900) ;
	assign n_8381 = (~n_943 & n_8380) ;
	assign n_935 = (~n_933 & ~n_934) ;
	assign n_925 = (~x_804 & ~n_923) ;
	assign n_924 = (x_804 & n_923) ;
	assign n_916 = (~n_913 & ~n_915) ;
	assign n_908 = (~n_901 & n_907) ;
	assign n_700 = (x_806 & n_699) ;
	assign n_691 = (i_26 & n_59) ;
	assign n_8382 = (~n_935 & n_8381) ;
	assign n_926 = (~n_924 & ~n_925) ;
	assign n_918 = (~x_805 & n_916) ;
	assign n_917 = (x_805 & ~n_916) ;
	assign n_909 = (~n_700 & ~n_908) ;
	assign n_692 = (n_66 & n_691) ;
	assign n_690 = (x_807 & n_60) ;
	assign n_684 = (~x_808 & ~n_544) ;
	assign n_8383 = (~n_926 & n_8382) ;
	assign n_919 = (~n_917 & ~n_918) ;
	assign n_911 = (~x_806 & n_909) ;
	assign n_910 = (x_806 & ~n_909) ;
	assign n_693 = (~n_690 & ~n_692) ;
	assign n_685 = (i_5 & ~n_684) ;
	assign n_683 = (~i_18 & n_544) ;
	assign n_670 = (~i_57 & n_669) ;
	assign n_667 = (~x_465 & ~n_544) ;
	assign n_8384 = (~n_919 & n_8383) ;
	assign n_912 = (~n_910 & ~n_911) ;
	assign n_695 = (~x_807 & n_693) ;
	assign n_694 = (x_807 & ~n_693) ;
	assign n_686 = (~n_683 & n_685) ;
	assign n_678 = (~n_302 & n_35) ;
	assign n_677 = (x_809 & n_36) ;
	assign n_671 = (i_5 & ~n_670) ;
	assign n_668 = (n_662 & n_667) ;
	assign n_8385 = (~n_912 & n_8384) ;
	assign n_696 = (~n_694 & ~n_695) ;
	assign n_688 = (~x_808 & ~n_686) ;
	assign n_687 = (x_808 & n_686) ;
	assign n_679 = (~n_677 & ~n_678) ;
	assign n_672 = (~n_668 & n_671) ;
	assign n_666 = (~x_810 & ~n_665) ;
	assign n_656 = (~x_811 & ~n_630) ;
	assign n_8386 = (~n_696 & n_8385) ;
	assign n_689 = (~n_687 & ~n_688) ;
	assign n_681 = (~x_809 & n_679) ;
	assign n_680 = (x_809 & ~n_679) ;
	assign n_673 = (~n_666 & n_672) ;
	assign n_657 = (i_5 & ~n_656) ;
	assign n_655 = (~i_65 & n_630) ;
	assign n_8387 = (~n_689 & n_8386) ;
	assign n_682 = (~n_680 & ~n_681) ;
	assign n_675 = (~x_810 & ~n_673) ;
	assign n_674 = (x_810 & n_673) ;
	assign n_658 = (~n_655 & n_657) ;
	assign n_650 = (x_569 & n_35) ;
	assign n_649 = (x_812 & n_36) ;
	assign n_643 = (i_44 & n_59) ;
	assign n_8388 = (~n_682 & n_8387) ;
	assign n_676 = (~n_674 & ~n_675) ;
	assign n_660 = (~x_811 & ~n_658) ;
	assign n_659 = (x_811 & n_658) ;
	assign n_651 = (~n_649 & ~n_650) ;
	assign n_644 = (n_66 & n_643) ;
	assign n_642 = (x_813 & n_60) ;
	assign n_525 = (~n_523 & ~n_524) ;
	assign n_8389 = (~n_676 & n_8388) ;
	assign n_661 = (~n_659 & ~n_660) ;
	assign n_653 = (~x_812 & n_651) ;
	assign n_652 = (x_812 & ~n_651) ;
	assign n_645 = (~n_642 & ~n_644) ;
	assign n_633 = (~x_815 & ~n_630) ;
	assign n_631 = (~n_630 & ~n_544) ;
	assign n_528 = (~x_508 & ~n_525) ;
	assign n_8390 = (~n_661 & n_8389) ;
	assign n_654 = (~n_652 & ~n_653) ;
	assign n_647 = (~x_813 & n_645) ;
	assign n_646 = (x_813 & ~n_645) ;
	assign n_634 = (i_5 & ~n_633) ;
	assign n_632 = (~n_628 & ~n_631) ;
	assign n_560 = (~x_816 & ~n_544) ;
	assign n_529 = (n_527 & ~n_528) ;
	assign n_526 = (x_508 & n_525) ;
	assign n_8391 = (~n_654 & n_8390) ;
	assign n_648 = (~n_646 & ~n_647) ;
	assign n_640 = (~x_814 & n_452) ;
	assign n_639 = (x_814 & ~n_452) ;
	assign n_635 = (~n_632 & n_634) ;
	assign n_561 = (i_5 & ~n_560) ;
	assign n_559 = (~i_16 & n_544) ;
	assign n_553 = (~x_817 & ~n_544) ;
	assign n_536 = (n_6 & n_75) ;
	assign n_530 = (~n_526 & n_529) ;
	assign n_8392 = (~n_648 & n_8391) ;
	assign n_641 = (~n_639 & ~n_640) ;
	assign n_637 = (~x_815 & ~n_635) ;
	assign n_636 = (x_815 & n_635) ;
	assign n_562 = (~n_559 & n_561) ;
	assign n_554 = (i_5 & ~n_553) ;
	assign n_552 = (~i_7 & n_544) ;
	assign n_546 = (~x_818 & ~n_544) ;
	assign n_537 = (~n_535 & ~n_536) ;
	assign n_532 = (n_75 & n_530) ;
	assign n_8393 = (~n_641 & n_8392) ;
	assign n_638 = (~n_636 & ~n_637) ;
	assign n_564 = (~x_816 & ~n_562) ;
	assign n_563 = (x_816 & n_562) ;
	assign n_555 = (~n_552 & n_554) ;
	assign n_547 = (i_5 & ~n_546) ;
	assign n_545 = (~i_27 & n_544) ;
	assign n_538 = (n_1 & ~n_537) ;
	assign n_533 = (~n_1 & ~n_532) ;
	assign n_531 = (~n_75 & ~n_530) ;
	assign n_8394 = (~n_638 & n_8393) ;
	assign n_565 = (~n_563 & ~n_564) ;
	assign n_557 = (~x_817 & ~n_555) ;
	assign n_556 = (x_817 & n_555) ;
	assign n_548 = (~n_545 & n_547) ;
	assign n_539 = (i_5 & ~n_538) ;
	assign n_534 = (~n_531 & n_533) ;
	assign n_67 = (i_22 & n_59) ;
	assign n_8395 = (~n_565 & n_8394) ;
	assign n_558 = (~n_556 & ~n_557) ;
	assign n_550 = (~x_818 & ~n_548) ;
	assign n_549 = (x_818 & n_548) ;
	assign n_540 = (~n_534 & n_539) ;
	assign n_68 = (n_66 & n_67) ;
	assign n_61 = (x_820 & n_60) ;
	assign n_8396 = (~n_558 & n_8395) ;
	assign n_551 = (~n_549 & ~n_550) ;
	assign n_542 = (~x_819 & ~n_540) ;
	assign n_541 = (x_819 & n_540) ;
	assign n_69 = (~n_61 & ~n_68) ;
	assign n_54 = (x_538 & n_53) ;
	assign n_52 = (x_821 & n_51) ;
	assign n_22 = (i_41 & n_7) ;
	assign n_21 = (x_712 & ~n_16) ;
	assign n_8397 = (~n_551 & n_8396) ;
	assign n_543 = (~n_541 & ~n_542) ;
	assign n_71 = (~x_820 & n_69) ;
	assign n_70 = (x_820 & ~n_69) ;
	assign n_55 = (~n_52 & ~n_54) ;
	assign n_38 = (x_463 & n_35) ;
	assign n_37 = (x_822 & n_36) ;
	assign n_23 = (~n_21 & ~n_22) ;
	assign n_8398 = (~n_543 & n_8397) ;
	assign n_72 = (~n_70 & ~n_71) ;
	assign n_57 = (~x_821 & n_55) ;
	assign n_56 = (x_821 & ~n_55) ;
	assign n_39 = (~n_37 & ~n_38) ;
	assign n_24 = (n_20 & ~n_23) ;
	assign n_19 = (x_823 & n_18) ;
	assign n_8399 = (~n_72 & n_8398) ;
	assign n_58 = (~n_56 & ~n_57) ;
	assign n_41 = (~x_822 & n_39) ;
	assign n_40 = (x_822 & ~n_39) ;
	assign n_25 = (~n_19 & ~n_24) ;
	assign n_8400 = (~n_58 & n_8399) ;
	assign n_42 = (~n_40 & ~n_41) ;
	assign n_27 = (~x_823 & n_25) ;
	assign n_26 = (x_823 & ~n_25) ;
	assign n_8401 = (~n_42 & n_8400) ;
	assign n_28 = (~n_26 & ~n_27) ;
	assign n_8402 = (~n_28 & n_8401) ;
	assign o_1 = ~n_8402 ;
endmodule
