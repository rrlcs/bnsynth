// skolem function for order file variables
// Generated using findDep.cpp 
module small-bug1-fixpoint-5 (v_1, v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_12, v_13, v_14, v_15, v_16, v_17, v_18, v_19, v_20, v_21, v_22, v_23, v_24, v_25, v_26, v_27, v_28, v_29, v_30, v_31, o_1);
input v_1;
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_13;
input v_14;
input v_15;
input v_16;
input v_17;
input v_18;
input v_19;
input v_20;
input v_21;
input v_22;
input v_23;
input v_24;
input v_25;
input v_26;
input v_27;
input v_28;
input v_29;
input v_30;
input v_31;
output o_1;
wire v_32;
wire v_33;
wire v_34;
wire v_35;
wire v_36;
wire v_37;
wire v_38;
wire v_39;
wire v_40;
wire v_41;
wire v_42;
wire v_43;
wire v_44;
wire v_45;
wire v_46;
wire v_47;
wire v_48;
wire v_49;
wire v_50;
wire v_51;
wire v_52;
wire v_53;
wire v_54;
wire v_55;
wire v_56;
wire v_57;
wire v_58;
wire v_59;
wire v_60;
wire v_61;
wire v_62;
wire v_63;
wire v_64;
wire v_65;
wire v_66;
wire v_67;
wire v_68;
wire v_69;
wire v_70;
wire v_71;
wire v_72;
wire v_73;
wire v_74;
wire v_75;
wire v_76;
wire v_77;
wire v_78;
wire v_79;
wire v_80;
wire v_81;
wire v_82;
wire v_83;
wire v_84;
wire v_85;
wire v_86;
wire v_87;
wire v_88;
wire v_89;
wire v_90;
wire v_91;
wire x_1;
assign v_32 = ~v_1 & v_9;
assign v_33 = ~v_8 & v_32;
assign v_36 = ~v_2 & v_7;
assign v_37 = ~v_11 & v_36;
assign v_40 = ~v_3 & v_10;
assign v_41 = ~v_13 & v_40;
assign v_44 = ~v_4 & v_12;
assign v_45 = ~v_15 & v_44;
assign v_48 = ~v_5 & v_14;
assign v_49 = ~v_17 & v_48;
assign v_52 = v_87 & v_88 & v_89;
assign v_53 = ~v_18 & v_25;
assign v_54 = ~v_24 & v_53;
assign v_57 = ~v_19 & v_23;
assign v_58 = ~v_27 & v_57;
assign v_61 = ~v_20 & v_26;
assign v_62 = ~v_29 & v_61;
assign v_65 = ~v_21 & v_28;
assign v_66 = ~v_31 & v_65;
assign v_69 = v_90 & v_91;
assign v_72 = ~v_70 & ~v_71;
assign v_75 = ~v_73 & ~v_74;
assign v_78 = ~v_76 & ~v_77;
assign v_81 = ~v_79 & ~v_80;
assign v_84 = ~v_82 & ~v_83;
assign v_86 = v_69 & v_85;
assign v_87 = ~v_1 & ~v_2 & ~v_3 & ~v_4 & ~v_5;
assign v_88 = ~v_6 & ~v_35 & ~v_39 & ~v_43 & ~v_47;
assign v_89 = ~v_51;
assign v_90 = ~v_18 & ~v_19 & ~v_20 & ~v_21 & ~v_22;
assign v_91 = ~v_56 & ~v_60 & ~v_64 & ~v_68;
assign v_34 = v_8 | v_33;
assign v_38 = v_11 | v_37;
assign v_42 = v_13 | v_41;
assign v_46 = v_15 | v_45;
assign v_50 = v_17 | v_49;
assign v_55 = v_24 | v_54;
assign v_59 = v_27 | v_58;
assign v_63 = v_29 | v_62;
assign v_67 = v_31 | v_66;
assign v_85 = v_72 | v_75 | v_78 | v_81 | v_84;
assign v_35 = v_34 ^ v_7;
assign v_39 = v_38 ^ v_10;
assign v_43 = v_42 ^ v_12;
assign v_47 = v_46 ^ v_14;
assign v_51 = v_50 ^ v_16;
assign v_56 = v_55 ^ v_23;
assign v_60 = v_59 ^ v_26;
assign v_64 = v_63 ^ v_28;
assign v_68 = v_67 ^ v_30;
assign v_70 = v_18 ^ v_6;
assign v_71 = v_25 ^ v_16;
assign v_73 = v_19 ^ v_6;
assign v_74 = v_23 ^ v_16;
assign v_76 = v_20 ^ v_6;
assign v_77 = v_26 ^ v_16;
assign v_79 = v_21 ^ v_6;
assign v_80 = v_28 ^ v_16;
assign v_82 = v_22 ^ v_6;
assign v_83 = v_30 ^ v_16;
assign x_1 = v_86 | ~v_52;
assign o_1 = x_1;
endmodule
