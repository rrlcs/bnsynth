// skolem function for order file variables
// Generated using findDep.cpp 
module rankfunc56_signed_64 (v_1, v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_12, v_13, v_14, v_15, v_16, v_17, v_18, v_19, v_20, v_21, v_22, v_23, v_24, v_25, v_26, v_27, v_28, v_29, v_30, v_31, v_32, v_33, v_34, v_35, v_36, v_37, v_38, v_39, v_40, v_41, v_42, v_43, v_44, v_45, v_46, v_47, v_48, v_49, v_50, v_51, v_52, v_53, v_54, v_55, v_56, v_57, v_58, v_59, v_60, v_61, v_62, v_63, v_64, v_65, v_66, v_67, v_68, v_69, v_70, v_71, v_72, v_73, v_74, v_75, v_76, v_77, v_78, v_79, v_80, v_81, v_82, v_83, v_84, v_85, v_86, v_87, v_88, v_89, v_90, v_91, v_92, v_93, v_94, v_95, v_96, v_97, v_98, v_99, v_100, v_101, v_102, v_103, v_104, v_105, v_106, v_107, v_108, v_109, v_110, v_111, v_112, v_113, v_114, v_115, v_116, v_117, v_118, v_119, v_120, v_121, v_122, v_123, v_124, v_125, v_126, v_127, v_128, v_129, v_130, v_131, v_132, v_133, v_134, v_135, v_136, v_137, v_138, v_139, v_140, v_141, v_142, v_143, v_144, v_145, v_146, v_147, v_148, v_149, v_150, v_151, v_152, v_153, v_154, v_155, v_156, v_157, v_158, v_159, v_160, v_161, v_162, v_163, v_164, v_165, v_166, v_167, v_168, v_169, v_170, v_171, v_172, v_173, v_174, v_175, v_176, v_177, v_178, v_179, v_180, v_181, v_182, v_183, v_184, v_185, v_186, v_187, v_188, v_189, v_190, v_191, v_192, v_193, v_194, v_195, v_196, v_197, v_198, v_199, v_200, v_201, v_202, v_203, v_204, v_205, v_206, v_207, v_208, v_209, v_210, v_211, v_212, v_213, v_214, v_215, v_216, v_217, v_218, v_219, v_220, v_221, v_222, v_223, v_224, v_225, v_226, v_227, v_228, v_229, v_230, v_231, v_232, v_233, v_234, v_235, v_236, v_237, v_238, v_239, v_240, v_241, v_242, v_243, v_244, v_245, v_246, v_247, v_248, v_249, v_250, v_251, v_252, v_253, v_254, v_255, v_256, v_257, v_258, v_259, v_260, v_261, v_262, v_263, v_264, v_265, v_266, v_267, v_268, v_269, v_270, v_271, v_272, v_273, v_274, v_275, v_276, v_277, v_278, v_279, v_280, v_281, v_282, v_283, v_284, v_285, v_286, v_287, v_288, v_289, v_290, v_291, v_292, v_293, v_294, v_295, v_296, v_297, v_298, v_299, v_300, v_301, v_302, v_303, v_304, v_305, v_306, v_307, v_308, v_309, v_310, v_311, v_312, v_313, v_314, v_315, v_316, v_317, v_318, v_319, v_320, v_449, v_451, v_452, v_453, v_454, v_455, v_456, v_457, v_458, v_459, v_460, v_461, v_462, v_463, v_464, v_465, v_466, v_467, v_468, v_469, v_470, v_471, v_472, v_473, v_474, v_475, v_476, v_477, v_478, v_479, v_480, v_481, v_482, v_483, v_484, v_485, v_486, v_487, v_488, v_489, v_490, v_491, v_492, v_493, v_494, v_495, v_496, v_497, v_498, v_499, v_500, v_501, v_502, v_503, v_504, v_505, v_506, v_507, v_508, v_509, v_510, v_511, v_512, v_513, v_514, v_517, v_780, v_781, v_782, v_783, v_784, v_785, v_786, v_787, v_788, v_789, v_790, v_791, v_792, v_793, v_794, v_795, v_796, v_797, v_798, v_799, v_800, v_801, v_802, v_803, v_804, v_805, v_806, v_807, v_808, v_809, v_810, v_811, v_812, v_813, v_814, v_815, v_816, v_817, v_818, v_819, v_820, v_821, v_822, v_823, v_824, v_825, v_826, v_827, v_828, v_829, v_830, v_831, v_832, v_833, v_834, v_835, v_836, v_837, v_838, v_839, v_840, v_841, v_842, v_843, v_844, v_845, v_846, v_847, v_848, v_849, v_850, v_851, v_852, v_853, v_854, v_855, v_856, v_857, v_858, v_859, v_860, v_861, v_862, v_863, v_864, v_865, v_866, v_867, v_868, v_869, v_870, v_871, v_872, v_873, v_874, v_875, v_876, v_877, v_878, v_879, v_880, v_881, v_882, v_883, v_884, v_885, v_886, v_887, v_888, v_889, v_890, v_891, v_892, v_893, v_894, v_895, v_896, v_897, v_898, v_899, v_900, v_901, v_902, v_903, v_904, v_905, v_906, v_907, v_1162, v_1164, v_1165, v_1166, v_1167, v_1168, v_1169, v_1170, v_1171, v_1172, v_1173, v_1174, v_1175, v_1176, v_1177, v_1178, v_1179, v_1180, v_1181, v_1182, v_1183, v_1184, v_1185, v_1186, v_1187, v_1188, v_1189, v_1190, v_1191, v_1192, v_1193, v_1194, v_1195, v_1196, v_1197, v_1198, v_1199, v_1200, v_1201, v_1202, v_1203, v_1204, v_1205, v_1206, v_1207, v_1208, v_1209, v_1210, v_1211, v_1212, v_1213, v_1214, v_1215, v_1216, v_1217, v_1218, v_1219, v_1220, v_1221, v_1222, v_1223, v_1224, v_1225, v_1226, v_1227, v_1228, v_1229, v_1230, v_1231, v_1232, v_1233, v_1234, v_1235, v_1236, v_1237, v_1238, v_1239, v_1240, v_1241, v_1242, v_1243, v_1244, v_1245, v_1246, v_1247, v_1248, v_1249, v_1250, v_1251, v_1252, v_1253, v_1254, v_1255, v_1256, v_1257, v_1258, v_1259, v_1260, v_1261, v_1262, v_1263, v_1264, v_1265, v_1266, v_1267, v_1268, v_1269, v_1270, v_1271, v_1272, v_1273, v_1274, v_1275, v_1276, v_1277, v_1278, v_1279, v_1280, v_1281, v_1282, v_1283, v_1284, v_1285, v_1286, v_1287, v_1288, v_1289, v_1290, v_1291, v_1546, o_1);
input v_1;
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_13;
input v_14;
input v_15;
input v_16;
input v_17;
input v_18;
input v_19;
input v_20;
input v_21;
input v_22;
input v_23;
input v_24;
input v_25;
input v_26;
input v_27;
input v_28;
input v_29;
input v_30;
input v_31;
input v_32;
input v_33;
input v_34;
input v_35;
input v_36;
input v_37;
input v_38;
input v_39;
input v_40;
input v_41;
input v_42;
input v_43;
input v_44;
input v_45;
input v_46;
input v_47;
input v_48;
input v_49;
input v_50;
input v_51;
input v_52;
input v_53;
input v_54;
input v_55;
input v_56;
input v_57;
input v_58;
input v_59;
input v_60;
input v_61;
input v_62;
input v_63;
input v_64;
input v_65;
input v_66;
input v_67;
input v_68;
input v_69;
input v_70;
input v_71;
input v_72;
input v_73;
input v_74;
input v_75;
input v_76;
input v_77;
input v_78;
input v_79;
input v_80;
input v_81;
input v_82;
input v_83;
input v_84;
input v_85;
input v_86;
input v_87;
input v_88;
input v_89;
input v_90;
input v_91;
input v_92;
input v_93;
input v_94;
input v_95;
input v_96;
input v_97;
input v_98;
input v_99;
input v_100;
input v_101;
input v_102;
input v_103;
input v_104;
input v_105;
input v_106;
input v_107;
input v_108;
input v_109;
input v_110;
input v_111;
input v_112;
input v_113;
input v_114;
input v_115;
input v_116;
input v_117;
input v_118;
input v_119;
input v_120;
input v_121;
input v_122;
input v_123;
input v_124;
input v_125;
input v_126;
input v_127;
input v_128;
input v_129;
input v_130;
input v_131;
input v_132;
input v_133;
input v_134;
input v_135;
input v_136;
input v_137;
input v_138;
input v_139;
input v_140;
input v_141;
input v_142;
input v_143;
input v_144;
input v_145;
input v_146;
input v_147;
input v_148;
input v_149;
input v_150;
input v_151;
input v_152;
input v_153;
input v_154;
input v_155;
input v_156;
input v_157;
input v_158;
input v_159;
input v_160;
input v_161;
input v_162;
input v_163;
input v_164;
input v_165;
input v_166;
input v_167;
input v_168;
input v_169;
input v_170;
input v_171;
input v_172;
input v_173;
input v_174;
input v_175;
input v_176;
input v_177;
input v_178;
input v_179;
input v_180;
input v_181;
input v_182;
input v_183;
input v_184;
input v_185;
input v_186;
input v_187;
input v_188;
input v_189;
input v_190;
input v_191;
input v_192;
input v_193;
input v_194;
input v_195;
input v_196;
input v_197;
input v_198;
input v_199;
input v_200;
input v_201;
input v_202;
input v_203;
input v_204;
input v_205;
input v_206;
input v_207;
input v_208;
input v_209;
input v_210;
input v_211;
input v_212;
input v_213;
input v_214;
input v_215;
input v_216;
input v_217;
input v_218;
input v_219;
input v_220;
input v_221;
input v_222;
input v_223;
input v_224;
input v_225;
input v_226;
input v_227;
input v_228;
input v_229;
input v_230;
input v_231;
input v_232;
input v_233;
input v_234;
input v_235;
input v_236;
input v_237;
input v_238;
input v_239;
input v_240;
input v_241;
input v_242;
input v_243;
input v_244;
input v_245;
input v_246;
input v_247;
input v_248;
input v_249;
input v_250;
input v_251;
input v_252;
input v_253;
input v_254;
input v_255;
input v_256;
input v_257;
input v_258;
input v_259;
input v_260;
input v_261;
input v_262;
input v_263;
input v_264;
input v_265;
input v_266;
input v_267;
input v_268;
input v_269;
input v_270;
input v_271;
input v_272;
input v_273;
input v_274;
input v_275;
input v_276;
input v_277;
input v_278;
input v_279;
input v_280;
input v_281;
input v_282;
input v_283;
input v_284;
input v_285;
input v_286;
input v_287;
input v_288;
input v_289;
input v_290;
input v_291;
input v_292;
input v_293;
input v_294;
input v_295;
input v_296;
input v_297;
input v_298;
input v_299;
input v_300;
input v_301;
input v_302;
input v_303;
input v_304;
input v_305;
input v_306;
input v_307;
input v_308;
input v_309;
input v_310;
input v_311;
input v_312;
input v_313;
input v_314;
input v_315;
input v_316;
input v_317;
input v_318;
input v_319;
input v_320;
input v_449;
input v_451;
input v_452;
input v_453;
input v_454;
input v_455;
input v_456;
input v_457;
input v_458;
input v_459;
input v_460;
input v_461;
input v_462;
input v_463;
input v_464;
input v_465;
input v_466;
input v_467;
input v_468;
input v_469;
input v_470;
input v_471;
input v_472;
input v_473;
input v_474;
input v_475;
input v_476;
input v_477;
input v_478;
input v_479;
input v_480;
input v_481;
input v_482;
input v_483;
input v_484;
input v_485;
input v_486;
input v_487;
input v_488;
input v_489;
input v_490;
input v_491;
input v_492;
input v_493;
input v_494;
input v_495;
input v_496;
input v_497;
input v_498;
input v_499;
input v_500;
input v_501;
input v_502;
input v_503;
input v_504;
input v_505;
input v_506;
input v_507;
input v_508;
input v_509;
input v_510;
input v_511;
input v_512;
input v_513;
input v_514;
input v_517;
input v_780;
input v_781;
input v_782;
input v_783;
input v_784;
input v_785;
input v_786;
input v_787;
input v_788;
input v_789;
input v_790;
input v_791;
input v_792;
input v_793;
input v_794;
input v_795;
input v_796;
input v_797;
input v_798;
input v_799;
input v_800;
input v_801;
input v_802;
input v_803;
input v_804;
input v_805;
input v_806;
input v_807;
input v_808;
input v_809;
input v_810;
input v_811;
input v_812;
input v_813;
input v_814;
input v_815;
input v_816;
input v_817;
input v_818;
input v_819;
input v_820;
input v_821;
input v_822;
input v_823;
input v_824;
input v_825;
input v_826;
input v_827;
input v_828;
input v_829;
input v_830;
input v_831;
input v_832;
input v_833;
input v_834;
input v_835;
input v_836;
input v_837;
input v_838;
input v_839;
input v_840;
input v_841;
input v_842;
input v_843;
input v_844;
input v_845;
input v_846;
input v_847;
input v_848;
input v_849;
input v_850;
input v_851;
input v_852;
input v_853;
input v_854;
input v_855;
input v_856;
input v_857;
input v_858;
input v_859;
input v_860;
input v_861;
input v_862;
input v_863;
input v_864;
input v_865;
input v_866;
input v_867;
input v_868;
input v_869;
input v_870;
input v_871;
input v_872;
input v_873;
input v_874;
input v_875;
input v_876;
input v_877;
input v_878;
input v_879;
input v_880;
input v_881;
input v_882;
input v_883;
input v_884;
input v_885;
input v_886;
input v_887;
input v_888;
input v_889;
input v_890;
input v_891;
input v_892;
input v_893;
input v_894;
input v_895;
input v_896;
input v_897;
input v_898;
input v_899;
input v_900;
input v_901;
input v_902;
input v_903;
input v_904;
input v_905;
input v_906;
input v_907;
input v_1162;
input v_1164;
input v_1165;
input v_1166;
input v_1167;
input v_1168;
input v_1169;
input v_1170;
input v_1171;
input v_1172;
input v_1173;
input v_1174;
input v_1175;
input v_1176;
input v_1177;
input v_1178;
input v_1179;
input v_1180;
input v_1181;
input v_1182;
input v_1183;
input v_1184;
input v_1185;
input v_1186;
input v_1187;
input v_1188;
input v_1189;
input v_1190;
input v_1191;
input v_1192;
input v_1193;
input v_1194;
input v_1195;
input v_1196;
input v_1197;
input v_1198;
input v_1199;
input v_1200;
input v_1201;
input v_1202;
input v_1203;
input v_1204;
input v_1205;
input v_1206;
input v_1207;
input v_1208;
input v_1209;
input v_1210;
input v_1211;
input v_1212;
input v_1213;
input v_1214;
input v_1215;
input v_1216;
input v_1217;
input v_1218;
input v_1219;
input v_1220;
input v_1221;
input v_1222;
input v_1223;
input v_1224;
input v_1225;
input v_1226;
input v_1227;
input v_1228;
input v_1229;
input v_1230;
input v_1231;
input v_1232;
input v_1233;
input v_1234;
input v_1235;
input v_1236;
input v_1237;
input v_1238;
input v_1239;
input v_1240;
input v_1241;
input v_1242;
input v_1243;
input v_1244;
input v_1245;
input v_1246;
input v_1247;
input v_1248;
input v_1249;
input v_1250;
input v_1251;
input v_1252;
input v_1253;
input v_1254;
input v_1255;
input v_1256;
input v_1257;
input v_1258;
input v_1259;
input v_1260;
input v_1261;
input v_1262;
input v_1263;
input v_1264;
input v_1265;
input v_1266;
input v_1267;
input v_1268;
input v_1269;
input v_1270;
input v_1271;
input v_1272;
input v_1273;
input v_1274;
input v_1275;
input v_1276;
input v_1277;
input v_1278;
input v_1279;
input v_1280;
input v_1281;
input v_1282;
input v_1283;
input v_1284;
input v_1285;
input v_1286;
input v_1287;
input v_1288;
input v_1289;
input v_1290;
input v_1291;
input v_1546;
output o_1;
wire v_321;
wire v_322;
wire v_323;
wire v_324;
wire v_325;
wire v_326;
wire v_327;
wire v_328;
wire v_329;
wire v_330;
wire v_331;
wire v_332;
wire v_333;
wire v_334;
wire v_335;
wire v_336;
wire v_337;
wire v_338;
wire v_339;
wire v_340;
wire v_341;
wire v_342;
wire v_343;
wire v_344;
wire v_345;
wire v_346;
wire v_347;
wire v_348;
wire v_349;
wire v_350;
wire v_351;
wire v_352;
wire v_353;
wire v_354;
wire v_355;
wire v_356;
wire v_357;
wire v_358;
wire v_359;
wire v_360;
wire v_361;
wire v_362;
wire v_363;
wire v_364;
wire v_365;
wire v_366;
wire v_367;
wire v_368;
wire v_369;
wire v_370;
wire v_371;
wire v_372;
wire v_373;
wire v_374;
wire v_375;
wire v_376;
wire v_377;
wire v_378;
wire v_379;
wire v_380;
wire v_381;
wire v_382;
wire v_383;
wire v_384;
wire v_385;
wire v_386;
wire v_387;
wire v_388;
wire v_389;
wire v_390;
wire v_391;
wire v_392;
wire v_393;
wire v_394;
wire v_395;
wire v_396;
wire v_397;
wire v_398;
wire v_399;
wire v_400;
wire v_401;
wire v_402;
wire v_403;
wire v_404;
wire v_405;
wire v_406;
wire v_407;
wire v_408;
wire v_409;
wire v_410;
wire v_411;
wire v_412;
wire v_413;
wire v_414;
wire v_415;
wire v_416;
wire v_417;
wire v_418;
wire v_419;
wire v_420;
wire v_421;
wire v_422;
wire v_423;
wire v_424;
wire v_425;
wire v_426;
wire v_427;
wire v_428;
wire v_429;
wire v_430;
wire v_431;
wire v_432;
wire v_433;
wire v_434;
wire v_435;
wire v_436;
wire v_437;
wire v_438;
wire v_439;
wire v_440;
wire v_441;
wire v_442;
wire v_443;
wire v_444;
wire v_445;
wire v_446;
wire v_447;
wire v_448;
wire v_450;
wire v_515;
wire v_516;
wire v_518;
wire v_519;
wire v_520;
wire v_521;
wire v_522;
wire v_523;
wire v_524;
wire v_525;
wire v_526;
wire v_527;
wire v_528;
wire v_529;
wire v_530;
wire v_531;
wire v_532;
wire v_533;
wire v_534;
wire v_535;
wire v_536;
wire v_537;
wire v_538;
wire v_539;
wire v_540;
wire v_541;
wire v_542;
wire v_543;
wire v_544;
wire v_545;
wire v_546;
wire v_547;
wire v_548;
wire v_549;
wire v_550;
wire v_551;
wire v_552;
wire v_553;
wire v_554;
wire v_555;
wire v_556;
wire v_557;
wire v_558;
wire v_559;
wire v_560;
wire v_561;
wire v_562;
wire v_563;
wire v_564;
wire v_565;
wire v_566;
wire v_567;
wire v_568;
wire v_569;
wire v_570;
wire v_571;
wire v_572;
wire v_573;
wire v_574;
wire v_575;
wire v_576;
wire v_577;
wire v_578;
wire v_579;
wire v_580;
wire v_581;
wire v_582;
wire v_583;
wire v_584;
wire v_585;
wire v_586;
wire v_587;
wire v_588;
wire v_589;
wire v_590;
wire v_591;
wire v_592;
wire v_593;
wire v_594;
wire v_595;
wire v_596;
wire v_597;
wire v_598;
wire v_599;
wire v_600;
wire v_601;
wire v_602;
wire v_603;
wire v_604;
wire v_605;
wire v_606;
wire v_607;
wire v_608;
wire v_609;
wire v_610;
wire v_611;
wire v_612;
wire v_613;
wire v_614;
wire v_615;
wire v_616;
wire v_617;
wire v_618;
wire v_619;
wire v_620;
wire v_621;
wire v_622;
wire v_623;
wire v_624;
wire v_625;
wire v_626;
wire v_627;
wire v_628;
wire v_629;
wire v_630;
wire v_631;
wire v_632;
wire v_633;
wire v_634;
wire v_635;
wire v_636;
wire v_637;
wire v_638;
wire v_639;
wire v_640;
wire v_641;
wire v_642;
wire v_643;
wire v_644;
wire v_645;
wire v_646;
wire v_647;
wire v_648;
wire v_649;
wire v_650;
wire v_651;
wire v_652;
wire v_653;
wire v_654;
wire v_655;
wire v_656;
wire v_657;
wire v_658;
wire v_659;
wire v_660;
wire v_661;
wire v_662;
wire v_663;
wire v_664;
wire v_665;
wire v_666;
wire v_667;
wire v_668;
wire v_669;
wire v_670;
wire v_671;
wire v_672;
wire v_673;
wire v_674;
wire v_675;
wire v_676;
wire v_677;
wire v_678;
wire v_679;
wire v_680;
wire v_681;
wire v_682;
wire v_683;
wire v_684;
wire v_685;
wire v_686;
wire v_687;
wire v_688;
wire v_689;
wire v_690;
wire v_691;
wire v_692;
wire v_693;
wire v_694;
wire v_695;
wire v_696;
wire v_697;
wire v_698;
wire v_699;
wire v_700;
wire v_701;
wire v_702;
wire v_703;
wire v_704;
wire v_705;
wire v_706;
wire v_707;
wire v_708;
wire v_709;
wire v_710;
wire v_711;
wire v_712;
wire v_713;
wire v_714;
wire v_715;
wire v_716;
wire v_717;
wire v_718;
wire v_719;
wire v_720;
wire v_721;
wire v_722;
wire v_723;
wire v_724;
wire v_725;
wire v_726;
wire v_727;
wire v_728;
wire v_729;
wire v_730;
wire v_731;
wire v_732;
wire v_733;
wire v_734;
wire v_735;
wire v_736;
wire v_737;
wire v_738;
wire v_739;
wire v_740;
wire v_741;
wire v_742;
wire v_743;
wire v_744;
wire v_745;
wire v_746;
wire v_747;
wire v_748;
wire v_749;
wire v_750;
wire v_751;
wire v_752;
wire v_753;
wire v_754;
wire v_755;
wire v_756;
wire v_757;
wire v_758;
wire v_759;
wire v_760;
wire v_761;
wire v_762;
wire v_763;
wire v_764;
wire v_765;
wire v_766;
wire v_767;
wire v_768;
wire v_769;
wire v_770;
wire v_771;
wire v_772;
wire v_773;
wire v_774;
wire v_775;
wire v_776;
wire v_777;
wire v_778;
wire v_779;
wire v_908;
wire v_909;
wire v_910;
wire v_911;
wire v_912;
wire v_913;
wire v_914;
wire v_915;
wire v_916;
wire v_917;
wire v_918;
wire v_919;
wire v_920;
wire v_921;
wire v_922;
wire v_923;
wire v_924;
wire v_925;
wire v_926;
wire v_927;
wire v_928;
wire v_929;
wire v_930;
wire v_931;
wire v_932;
wire v_933;
wire v_934;
wire v_935;
wire v_936;
wire v_937;
wire v_938;
wire v_939;
wire v_940;
wire v_941;
wire v_942;
wire v_943;
wire v_944;
wire v_945;
wire v_946;
wire v_947;
wire v_948;
wire v_949;
wire v_950;
wire v_951;
wire v_952;
wire v_953;
wire v_954;
wire v_955;
wire v_956;
wire v_957;
wire v_958;
wire v_959;
wire v_960;
wire v_961;
wire v_962;
wire v_963;
wire v_964;
wire v_965;
wire v_966;
wire v_967;
wire v_968;
wire v_969;
wire v_970;
wire v_971;
wire v_972;
wire v_973;
wire v_974;
wire v_975;
wire v_976;
wire v_977;
wire v_978;
wire v_979;
wire v_980;
wire v_981;
wire v_982;
wire v_983;
wire v_984;
wire v_985;
wire v_986;
wire v_987;
wire v_988;
wire v_989;
wire v_990;
wire v_991;
wire v_992;
wire v_993;
wire v_994;
wire v_995;
wire v_996;
wire v_997;
wire v_998;
wire v_999;
wire v_1000;
wire v_1001;
wire v_1002;
wire v_1003;
wire v_1004;
wire v_1005;
wire v_1006;
wire v_1007;
wire v_1008;
wire v_1009;
wire v_1010;
wire v_1011;
wire v_1012;
wire v_1013;
wire v_1014;
wire v_1015;
wire v_1016;
wire v_1017;
wire v_1018;
wire v_1019;
wire v_1020;
wire v_1021;
wire v_1022;
wire v_1023;
wire v_1024;
wire v_1025;
wire v_1026;
wire v_1027;
wire v_1028;
wire v_1029;
wire v_1030;
wire v_1031;
wire v_1032;
wire v_1033;
wire v_1034;
wire v_1035;
wire v_1036;
wire v_1037;
wire v_1038;
wire v_1039;
wire v_1040;
wire v_1041;
wire v_1042;
wire v_1043;
wire v_1044;
wire v_1045;
wire v_1046;
wire v_1047;
wire v_1048;
wire v_1049;
wire v_1050;
wire v_1051;
wire v_1052;
wire v_1053;
wire v_1054;
wire v_1055;
wire v_1056;
wire v_1057;
wire v_1058;
wire v_1059;
wire v_1060;
wire v_1061;
wire v_1062;
wire v_1063;
wire v_1064;
wire v_1065;
wire v_1066;
wire v_1067;
wire v_1068;
wire v_1069;
wire v_1070;
wire v_1071;
wire v_1072;
wire v_1073;
wire v_1074;
wire v_1075;
wire v_1076;
wire v_1077;
wire v_1078;
wire v_1079;
wire v_1080;
wire v_1081;
wire v_1082;
wire v_1083;
wire v_1084;
wire v_1085;
wire v_1086;
wire v_1087;
wire v_1088;
wire v_1089;
wire v_1090;
wire v_1091;
wire v_1092;
wire v_1093;
wire v_1094;
wire v_1095;
wire v_1096;
wire v_1097;
wire v_1098;
wire v_1099;
wire v_1100;
wire v_1101;
wire v_1102;
wire v_1103;
wire v_1104;
wire v_1105;
wire v_1106;
wire v_1107;
wire v_1108;
wire v_1109;
wire v_1110;
wire v_1111;
wire v_1112;
wire v_1113;
wire v_1114;
wire v_1115;
wire v_1116;
wire v_1117;
wire v_1118;
wire v_1119;
wire v_1120;
wire v_1121;
wire v_1122;
wire v_1123;
wire v_1124;
wire v_1125;
wire v_1126;
wire v_1127;
wire v_1128;
wire v_1129;
wire v_1130;
wire v_1131;
wire v_1132;
wire v_1133;
wire v_1134;
wire v_1135;
wire v_1136;
wire v_1137;
wire v_1138;
wire v_1139;
wire v_1140;
wire v_1141;
wire v_1142;
wire v_1143;
wire v_1144;
wire v_1145;
wire v_1146;
wire v_1147;
wire v_1148;
wire v_1149;
wire v_1150;
wire v_1151;
wire v_1152;
wire v_1153;
wire v_1154;
wire v_1155;
wire v_1156;
wire v_1157;
wire v_1158;
wire v_1159;
wire v_1160;
wire v_1161;
wire v_1163;
wire v_1292;
wire v_1293;
wire v_1294;
wire v_1295;
wire v_1296;
wire v_1297;
wire v_1298;
wire v_1299;
wire v_1300;
wire v_1301;
wire v_1302;
wire v_1303;
wire v_1304;
wire v_1305;
wire v_1306;
wire v_1307;
wire v_1308;
wire v_1309;
wire v_1310;
wire v_1311;
wire v_1312;
wire v_1313;
wire v_1314;
wire v_1315;
wire v_1316;
wire v_1317;
wire v_1318;
wire v_1319;
wire v_1320;
wire v_1321;
wire v_1322;
wire v_1323;
wire v_1324;
wire v_1325;
wire v_1326;
wire v_1327;
wire v_1328;
wire v_1329;
wire v_1330;
wire v_1331;
wire v_1332;
wire v_1333;
wire v_1334;
wire v_1335;
wire v_1336;
wire v_1337;
wire v_1338;
wire v_1339;
wire v_1340;
wire v_1341;
wire v_1342;
wire v_1343;
wire v_1344;
wire v_1345;
wire v_1346;
wire v_1347;
wire v_1348;
wire v_1349;
wire v_1350;
wire v_1351;
wire v_1352;
wire v_1353;
wire v_1354;
wire v_1355;
wire v_1356;
wire v_1357;
wire v_1358;
wire v_1359;
wire v_1360;
wire v_1361;
wire v_1362;
wire v_1363;
wire v_1364;
wire v_1365;
wire v_1366;
wire v_1367;
wire v_1368;
wire v_1369;
wire v_1370;
wire v_1371;
wire v_1372;
wire v_1373;
wire v_1374;
wire v_1375;
wire v_1376;
wire v_1377;
wire v_1378;
wire v_1379;
wire v_1380;
wire v_1381;
wire v_1382;
wire v_1383;
wire v_1384;
wire v_1385;
wire v_1386;
wire v_1387;
wire v_1388;
wire v_1389;
wire v_1390;
wire v_1391;
wire v_1392;
wire v_1393;
wire v_1394;
wire v_1395;
wire v_1396;
wire v_1397;
wire v_1398;
wire v_1399;
wire v_1400;
wire v_1401;
wire v_1402;
wire v_1403;
wire v_1404;
wire v_1405;
wire v_1406;
wire v_1407;
wire v_1408;
wire v_1409;
wire v_1410;
wire v_1411;
wire v_1412;
wire v_1413;
wire v_1414;
wire v_1415;
wire v_1416;
wire v_1417;
wire v_1418;
wire v_1419;
wire v_1420;
wire v_1421;
wire v_1422;
wire v_1423;
wire v_1424;
wire v_1425;
wire v_1426;
wire v_1427;
wire v_1428;
wire v_1429;
wire v_1430;
wire v_1431;
wire v_1432;
wire v_1433;
wire v_1434;
wire v_1435;
wire v_1436;
wire v_1437;
wire v_1438;
wire v_1439;
wire v_1440;
wire v_1441;
wire v_1442;
wire v_1443;
wire v_1444;
wire v_1445;
wire v_1446;
wire v_1447;
wire v_1448;
wire v_1449;
wire v_1450;
wire v_1451;
wire v_1452;
wire v_1453;
wire v_1454;
wire v_1455;
wire v_1456;
wire v_1457;
wire v_1458;
wire v_1459;
wire v_1460;
wire v_1461;
wire v_1462;
wire v_1463;
wire v_1464;
wire v_1465;
wire v_1466;
wire v_1467;
wire v_1468;
wire v_1469;
wire v_1470;
wire v_1471;
wire v_1472;
wire v_1473;
wire v_1474;
wire v_1475;
wire v_1476;
wire v_1477;
wire v_1478;
wire v_1479;
wire v_1480;
wire v_1481;
wire v_1482;
wire v_1483;
wire v_1484;
wire v_1485;
wire v_1486;
wire v_1487;
wire v_1488;
wire v_1489;
wire v_1490;
wire v_1491;
wire v_1492;
wire v_1493;
wire v_1494;
wire v_1495;
wire v_1496;
wire v_1497;
wire v_1498;
wire v_1499;
wire v_1500;
wire v_1501;
wire v_1502;
wire v_1503;
wire v_1504;
wire v_1505;
wire v_1506;
wire v_1507;
wire v_1508;
wire v_1509;
wire v_1510;
wire v_1511;
wire v_1512;
wire v_1513;
wire v_1514;
wire v_1515;
wire v_1516;
wire v_1517;
wire v_1518;
wire v_1519;
wire v_1520;
wire v_1521;
wire v_1522;
wire v_1523;
wire v_1524;
wire v_1525;
wire v_1526;
wire v_1527;
wire v_1528;
wire v_1529;
wire v_1530;
wire v_1531;
wire v_1532;
wire v_1533;
wire v_1534;
wire v_1535;
wire v_1536;
wire v_1537;
wire v_1538;
wire v_1539;
wire v_1540;
wire v_1541;
wire v_1542;
wire v_1543;
wire v_1544;
wire v_1545;
wire v_1547;
wire v_1548;
wire v_1549;
wire v_1550;
wire v_1551;
wire v_1552;
wire v_1553;
wire v_1554;
wire v_1555;
wire v_1556;
wire v_1557;
wire v_1558;
wire v_1559;
wire v_1560;
wire v_1561;
wire v_1562;
wire v_1563;
wire v_1564;
wire v_1565;
wire v_1566;
wire v_1567;
wire v_1568;
wire v_1569;
wire v_1570;
wire v_1571;
wire v_1572;
wire v_1573;
wire v_1574;
wire v_1575;
wire v_1576;
wire v_1577;
wire v_1578;
wire v_1579;
wire v_1580;
wire v_1581;
wire v_1582;
wire v_1583;
wire v_1584;
wire v_1585;
wire v_1586;
wire v_1587;
wire v_1588;
wire v_1589;
wire v_1590;
wire v_1591;
wire v_1592;
wire v_1593;
wire v_1594;
wire v_1595;
wire v_1596;
wire v_1597;
wire v_1598;
wire v_1599;
wire v_1600;
wire v_1601;
wire v_1602;
wire v_1603;
wire v_1604;
wire v_1605;
wire v_1606;
wire v_1607;
wire v_1608;
wire v_1609;
wire v_1610;
wire v_1611;
wire v_1612;
wire v_1613;
wire v_1614;
wire v_1615;
wire v_1616;
wire v_1617;
wire v_1618;
wire v_1619;
wire v_1620;
wire v_1621;
wire v_1622;
wire v_1623;
wire v_1624;
wire v_1625;
wire v_1626;
wire v_1627;
wire v_1628;
wire v_1629;
wire v_1630;
wire v_1631;
wire v_1632;
wire v_1633;
wire v_1634;
wire v_1635;
wire v_1636;
wire v_1637;
wire v_1638;
wire v_1639;
wire v_1640;
wire v_1641;
wire v_1642;
wire v_1643;
wire v_1644;
wire v_1645;
wire v_1646;
wire v_1647;
wire v_1648;
wire v_1649;
wire v_1650;
wire v_1651;
wire v_1652;
wire v_1653;
wire v_1654;
wire v_1655;
wire v_1656;
wire v_1657;
wire v_1658;
wire v_1659;
wire v_1660;
wire v_1661;
wire v_1662;
wire v_1663;
wire v_1664;
wire v_1665;
wire v_1666;
wire v_1667;
wire v_1668;
wire v_1669;
wire v_1670;
wire v_1671;
wire v_1672;
wire v_1673;
wire v_1674;
wire v_1675;
wire v_1676;
wire v_1677;
wire v_1678;
wire v_1679;
wire v_1680;
wire v_1681;
wire v_1682;
wire v_1683;
wire v_1684;
wire v_1685;
wire v_1686;
wire v_1687;
wire v_1688;
wire v_1689;
wire v_1690;
wire v_1691;
wire v_1692;
wire v_1693;
wire v_1694;
wire v_1695;
wire v_1696;
wire v_1697;
wire v_1698;
wire v_1699;
wire v_1700;
wire v_1701;
wire v_1702;
wire v_1703;
wire v_1704;
wire v_1705;
wire v_1706;
wire v_1707;
wire v_1708;
wire v_1709;
wire v_1710;
wire v_1711;
wire v_1712;
wire v_1713;
wire v_1714;
wire v_1715;
wire v_1716;
wire v_1717;
wire v_1718;
wire v_1719;
wire v_1720;
wire v_1721;
wire v_1722;
wire v_1723;
wire v_1724;
wire v_1725;
wire v_1726;
wire v_1727;
wire v_1728;
wire v_1729;
wire v_1730;
wire v_1731;
wire v_1732;
wire v_1733;
wire v_1734;
wire v_1735;
wire v_1736;
wire v_1737;
wire v_1738;
wire v_1739;
wire v_1740;
wire v_1741;
wire v_1742;
wire v_1743;
wire v_1744;
wire v_1745;
wire v_1746;
wire v_1747;
wire v_1748;
wire v_1749;
wire v_1750;
wire v_1751;
wire v_1752;
wire v_1753;
wire v_1754;
wire v_1755;
wire v_1756;
wire v_1757;
wire v_1758;
wire v_1759;
wire v_1760;
wire v_1761;
wire v_1762;
wire v_1763;
wire v_1764;
wire v_1765;
wire v_1766;
wire v_1767;
wire v_1768;
wire v_1769;
wire v_1770;
wire v_1771;
wire v_1772;
wire v_1773;
wire v_1774;
wire v_1775;
wire v_1776;
wire v_1777;
wire v_1778;
wire v_1779;
wire v_1780;
wire v_1781;
wire v_1782;
wire v_1783;
wire v_1784;
wire v_1785;
wire v_1786;
wire v_1787;
wire v_1788;
wire v_1789;
wire v_1790;
wire v_1791;
wire v_1792;
wire v_1793;
wire v_1794;
wire v_1795;
wire v_1796;
wire v_1797;
wire v_1798;
wire v_1799;
wire v_1800;
wire v_1801;
wire v_1802;
wire v_1803;
wire v_1804;
wire v_1805;
wire v_1806;
wire v_1807;
wire v_1808;
wire v_1809;
wire v_1810;
wire v_1811;
wire v_1812;
wire v_1813;
wire v_1814;
wire v_1815;
wire v_1816;
wire v_1817;
wire v_1818;
wire v_1819;
wire v_1820;
wire v_1821;
wire v_1822;
wire v_1823;
wire v_1824;
wire v_1825;
wire v_1826;
wire v_1827;
wire v_1828;
wire v_1829;
wire v_1830;
wire v_1831;
wire v_1832;
wire v_1833;
wire v_1834;
wire v_1835;
wire v_1836;
wire v_1837;
wire v_1838;
wire v_1839;
wire v_1840;
wire v_1841;
wire v_1842;
wire v_1843;
wire v_1844;
wire v_1845;
wire v_1846;
wire v_1847;
wire v_1848;
wire v_1849;
wire v_1850;
wire v_1851;
wire v_1852;
wire v_1853;
wire v_1854;
wire v_1855;
wire v_1856;
wire v_1857;
wire v_1858;
wire v_1859;
wire v_1860;
wire v_1861;
wire v_1862;
wire v_1863;
wire v_1864;
wire v_1865;
wire v_1866;
wire v_1867;
wire v_1868;
wire v_1869;
wire v_1870;
wire v_1871;
wire v_1872;
wire v_1873;
wire v_1874;
wire v_1875;
wire v_1876;
wire v_1877;
wire v_1878;
wire v_1879;
wire v_1880;
wire v_1881;
wire v_1882;
wire v_1883;
wire v_1884;
wire v_1885;
wire v_1886;
wire v_1887;
wire v_1888;
wire v_1889;
wire v_1890;
wire v_1891;
wire v_1892;
wire v_1893;
wire v_1894;
wire v_1895;
wire v_1896;
wire v_1897;
wire v_1898;
wire v_1899;
wire v_1900;
wire v_1901;
wire v_1902;
wire v_1903;
wire v_1904;
wire v_1905;
wire v_1906;
wire v_1907;
wire v_1908;
wire v_1909;
wire v_1910;
wire v_1911;
wire v_1912;
wire v_1913;
wire v_1914;
wire v_1915;
wire v_1916;
wire v_1917;
wire v_1918;
wire v_1919;
wire v_1920;
wire v_1921;
wire v_1922;
wire v_1923;
wire v_1924;
wire v_1925;
wire v_1926;
wire v_1927;
wire v_1928;
wire v_1929;
wire v_1930;
wire v_1931;
wire v_1932;
wire v_1933;
wire v_1934;
wire v_1935;
wire v_1936;
wire v_1937;
wire v_1938;
wire v_1939;
wire v_1940;
wire v_1941;
wire v_1942;
wire v_1943;
wire v_1944;
wire v_1945;
wire v_1946;
wire v_1947;
wire v_1948;
wire v_1949;
wire v_1950;
wire v_1951;
wire v_1952;
wire v_1953;
wire v_1954;
wire x_1;
wire x_2;
wire x_3;
wire x_4;
wire x_5;
wire x_6;
wire x_7;
wire x_8;
wire x_9;
wire x_10;
wire x_11;
wire x_12;
wire x_13;
assign v_450 = 1;
assign v_518 = 1;
assign v_1163 = 1;
assign v_1547 = 1;
assign v_321 = ~v_257;
assign v_322 = ~v_258 & v_321;
assign v_323 = v_322;
assign v_324 = ~v_259 & v_323;
assign v_325 = v_324;
assign v_326 = ~v_260 & v_325;
assign v_327 = v_326;
assign v_328 = ~v_261 & v_327;
assign v_329 = v_328;
assign v_330 = ~v_262 & v_329;
assign v_331 = v_330;
assign v_332 = ~v_263 & v_331;
assign v_333 = v_332;
assign v_334 = ~v_264 & v_333;
assign v_335 = v_334;
assign v_336 = ~v_265 & v_335;
assign v_337 = v_336;
assign v_338 = ~v_266 & v_337;
assign v_339 = v_338;
assign v_340 = ~v_267 & v_339;
assign v_341 = v_340;
assign v_342 = ~v_268 & v_341;
assign v_343 = v_342;
assign v_344 = ~v_269 & v_343;
assign v_345 = v_344;
assign v_346 = ~v_270 & v_345;
assign v_347 = v_346;
assign v_348 = ~v_271 & v_347;
assign v_349 = v_348;
assign v_350 = ~v_272 & v_349;
assign v_351 = v_350;
assign v_352 = ~v_273 & v_351;
assign v_353 = v_352;
assign v_354 = ~v_274 & v_353;
assign v_355 = v_354;
assign v_356 = ~v_275 & v_355;
assign v_357 = v_356;
assign v_358 = ~v_276 & v_357;
assign v_359 = v_358;
assign v_360 = ~v_277 & v_359;
assign v_361 = v_360;
assign v_362 = ~v_278 & v_361;
assign v_363 = v_362;
assign v_364 = ~v_279 & v_363;
assign v_365 = v_364;
assign v_366 = ~v_280 & v_365;
assign v_367 = v_366;
assign v_368 = ~v_281 & v_367;
assign v_369 = v_368;
assign v_370 = ~v_282 & v_369;
assign v_371 = v_370;
assign v_372 = ~v_283 & v_371;
assign v_373 = v_372;
assign v_374 = ~v_284 & v_373;
assign v_375 = v_374;
assign v_376 = ~v_285 & v_375;
assign v_377 = v_376;
assign v_378 = ~v_286 & v_377;
assign v_379 = v_378;
assign v_380 = ~v_287 & v_379;
assign v_381 = v_380;
assign v_382 = ~v_288 & v_381;
assign v_383 = v_382;
assign v_384 = ~v_289 & v_383;
assign v_385 = v_384;
assign v_386 = ~v_290 & v_385;
assign v_387 = v_386;
assign v_388 = ~v_291 & v_387;
assign v_389 = v_388;
assign v_390 = ~v_292 & v_389;
assign v_391 = v_390;
assign v_392 = ~v_293 & v_391;
assign v_393 = v_392;
assign v_394 = ~v_294 & v_393;
assign v_395 = v_394;
assign v_396 = ~v_295 & v_395;
assign v_397 = v_396;
assign v_398 = ~v_296 & v_397;
assign v_399 = v_398;
assign v_400 = ~v_297 & v_399;
assign v_401 = v_400;
assign v_402 = ~v_298 & v_401;
assign v_403 = v_402;
assign v_404 = ~v_299 & v_403;
assign v_405 = v_404;
assign v_406 = ~v_300 & v_405;
assign v_407 = v_406;
assign v_408 = ~v_301 & v_407;
assign v_409 = v_408;
assign v_410 = ~v_302 & v_409;
assign v_411 = v_410;
assign v_412 = ~v_303 & v_411;
assign v_413 = v_412;
assign v_414 = ~v_304 & v_413;
assign v_415 = v_414;
assign v_416 = ~v_305 & v_415;
assign v_417 = v_416;
assign v_418 = ~v_306 & v_417;
assign v_419 = v_418;
assign v_420 = ~v_307 & v_419;
assign v_421 = v_420;
assign v_422 = ~v_308 & v_421;
assign v_423 = v_422;
assign v_424 = ~v_309 & v_423;
assign v_425 = v_424;
assign v_426 = ~v_310 & v_425;
assign v_427 = v_426;
assign v_428 = ~v_311 & v_427;
assign v_429 = v_428;
assign v_430 = ~v_312 & v_429;
assign v_431 = v_430;
assign v_432 = ~v_313 & v_431;
assign v_433 = v_432;
assign v_434 = ~v_314 & v_433;
assign v_435 = v_434;
assign v_436 = ~v_315 & v_435;
assign v_437 = v_436;
assign v_438 = ~v_316 & v_437;
assign v_439 = v_438;
assign v_440 = ~v_317 & v_439;
assign v_441 = v_440;
assign v_442 = ~v_318 & v_441;
assign v_443 = v_442;
assign v_444 = ~v_319 & v_443;
assign v_445 = v_444;
assign v_446 = ~v_320 & v_445;
assign v_447 = v_446;
assign v_583 = v_1822 & v_1823 & v_1824;
assign v_648 = v_1838 & v_1839 & v_1840;
assign v_713 = v_1854 & v_1855 & v_1856;
assign v_778 = v_1870 & v_1871 & v_1872;
assign v_779 = v_1873 & v_1874;
assign v_908 = ~v_780 & v_844;
assign v_910 = ~v_781 & v_845;
assign v_911 = v_845 & v_909;
assign v_912 = ~v_781 & v_909;
assign v_914 = ~v_782 & v_846;
assign v_915 = v_846 & v_913;
assign v_916 = ~v_782 & v_913;
assign v_918 = ~v_783 & v_847;
assign v_919 = v_847 & v_917;
assign v_920 = ~v_783 & v_917;
assign v_922 = ~v_784 & v_848;
assign v_923 = v_848 & v_921;
assign v_924 = ~v_784 & v_921;
assign v_926 = ~v_785 & v_849;
assign v_927 = v_849 & v_925;
assign v_928 = ~v_785 & v_925;
assign v_930 = ~v_786 & v_850;
assign v_931 = v_850 & v_929;
assign v_932 = ~v_786 & v_929;
assign v_934 = ~v_787 & v_851;
assign v_935 = v_851 & v_933;
assign v_936 = ~v_787 & v_933;
assign v_938 = ~v_788 & v_852;
assign v_939 = v_852 & v_937;
assign v_940 = ~v_788 & v_937;
assign v_942 = ~v_789 & v_853;
assign v_943 = v_853 & v_941;
assign v_944 = ~v_789 & v_941;
assign v_946 = ~v_790 & v_854;
assign v_947 = v_854 & v_945;
assign v_948 = ~v_790 & v_945;
assign v_950 = ~v_791 & v_855;
assign v_951 = v_855 & v_949;
assign v_952 = ~v_791 & v_949;
assign v_954 = ~v_792 & v_856;
assign v_955 = v_856 & v_953;
assign v_956 = ~v_792 & v_953;
assign v_958 = ~v_793 & v_857;
assign v_959 = v_857 & v_957;
assign v_960 = ~v_793 & v_957;
assign v_962 = ~v_794 & v_858;
assign v_963 = v_858 & v_961;
assign v_964 = ~v_794 & v_961;
assign v_966 = ~v_795 & v_859;
assign v_967 = v_859 & v_965;
assign v_968 = ~v_795 & v_965;
assign v_970 = ~v_796 & v_860;
assign v_971 = v_860 & v_969;
assign v_972 = ~v_796 & v_969;
assign v_974 = ~v_797 & v_861;
assign v_975 = v_861 & v_973;
assign v_976 = ~v_797 & v_973;
assign v_978 = ~v_798 & v_862;
assign v_979 = v_862 & v_977;
assign v_980 = ~v_798 & v_977;
assign v_982 = ~v_799 & v_863;
assign v_983 = v_863 & v_981;
assign v_984 = ~v_799 & v_981;
assign v_986 = ~v_800 & v_864;
assign v_987 = v_864 & v_985;
assign v_988 = ~v_800 & v_985;
assign v_990 = ~v_801 & v_865;
assign v_991 = v_865 & v_989;
assign v_992 = ~v_801 & v_989;
assign v_994 = ~v_802 & v_866;
assign v_995 = v_866 & v_993;
assign v_996 = ~v_802 & v_993;
assign v_998 = ~v_803 & v_867;
assign v_999 = v_867 & v_997;
assign v_1000 = ~v_803 & v_997;
assign v_1002 = ~v_804 & v_868;
assign v_1003 = v_868 & v_1001;
assign v_1004 = ~v_804 & v_1001;
assign v_1006 = ~v_805 & v_869;
assign v_1007 = v_869 & v_1005;
assign v_1008 = ~v_805 & v_1005;
assign v_1010 = ~v_806 & v_870;
assign v_1011 = v_870 & v_1009;
assign v_1012 = ~v_806 & v_1009;
assign v_1014 = ~v_807 & v_871;
assign v_1015 = v_871 & v_1013;
assign v_1016 = ~v_807 & v_1013;
assign v_1018 = ~v_808 & v_872;
assign v_1019 = v_872 & v_1017;
assign v_1020 = ~v_808 & v_1017;
assign v_1022 = ~v_809 & v_873;
assign v_1023 = v_873 & v_1021;
assign v_1024 = ~v_809 & v_1021;
assign v_1026 = ~v_810 & v_874;
assign v_1027 = v_874 & v_1025;
assign v_1028 = ~v_810 & v_1025;
assign v_1030 = ~v_811 & v_875;
assign v_1031 = v_875 & v_1029;
assign v_1032 = ~v_811 & v_1029;
assign v_1034 = ~v_812 & v_876;
assign v_1035 = v_876 & v_1033;
assign v_1036 = ~v_812 & v_1033;
assign v_1038 = ~v_813 & v_877;
assign v_1039 = v_877 & v_1037;
assign v_1040 = ~v_813 & v_1037;
assign v_1042 = ~v_814 & v_878;
assign v_1043 = v_878 & v_1041;
assign v_1044 = ~v_814 & v_1041;
assign v_1046 = ~v_815 & v_879;
assign v_1047 = v_879 & v_1045;
assign v_1048 = ~v_815 & v_1045;
assign v_1050 = ~v_816 & v_880;
assign v_1051 = v_880 & v_1049;
assign v_1052 = ~v_816 & v_1049;
assign v_1054 = ~v_817 & v_881;
assign v_1055 = v_881 & v_1053;
assign v_1056 = ~v_817 & v_1053;
assign v_1058 = ~v_818 & v_882;
assign v_1059 = v_882 & v_1057;
assign v_1060 = ~v_818 & v_1057;
assign v_1062 = ~v_819 & v_883;
assign v_1063 = v_883 & v_1061;
assign v_1064 = ~v_819 & v_1061;
assign v_1066 = ~v_820 & v_884;
assign v_1067 = v_884 & v_1065;
assign v_1068 = ~v_820 & v_1065;
assign v_1070 = ~v_821 & v_885;
assign v_1071 = v_885 & v_1069;
assign v_1072 = ~v_821 & v_1069;
assign v_1074 = ~v_822 & v_886;
assign v_1075 = v_886 & v_1073;
assign v_1076 = ~v_822 & v_1073;
assign v_1078 = ~v_823 & v_887;
assign v_1079 = v_887 & v_1077;
assign v_1080 = ~v_823 & v_1077;
assign v_1082 = ~v_824 & v_888;
assign v_1083 = v_888 & v_1081;
assign v_1084 = ~v_824 & v_1081;
assign v_1086 = ~v_825 & v_889;
assign v_1087 = v_889 & v_1085;
assign v_1088 = ~v_825 & v_1085;
assign v_1090 = ~v_826 & v_890;
assign v_1091 = v_890 & v_1089;
assign v_1092 = ~v_826 & v_1089;
assign v_1094 = ~v_827 & v_891;
assign v_1095 = v_891 & v_1093;
assign v_1096 = ~v_827 & v_1093;
assign v_1098 = ~v_828 & v_892;
assign v_1099 = v_892 & v_1097;
assign v_1100 = ~v_828 & v_1097;
assign v_1102 = ~v_829 & v_893;
assign v_1103 = v_893 & v_1101;
assign v_1104 = ~v_829 & v_1101;
assign v_1106 = ~v_830 & v_894;
assign v_1107 = v_894 & v_1105;
assign v_1108 = ~v_830 & v_1105;
assign v_1110 = ~v_831 & v_895;
assign v_1111 = v_895 & v_1109;
assign v_1112 = ~v_831 & v_1109;
assign v_1114 = ~v_832 & v_896;
assign v_1115 = v_896 & v_1113;
assign v_1116 = ~v_832 & v_1113;
assign v_1118 = ~v_833 & v_897;
assign v_1119 = v_897 & v_1117;
assign v_1120 = ~v_833 & v_1117;
assign v_1122 = ~v_834 & v_898;
assign v_1123 = v_898 & v_1121;
assign v_1124 = ~v_834 & v_1121;
assign v_1126 = ~v_835 & v_899;
assign v_1127 = v_899 & v_1125;
assign v_1128 = ~v_835 & v_1125;
assign v_1130 = ~v_836 & v_900;
assign v_1131 = v_900 & v_1129;
assign v_1132 = ~v_836 & v_1129;
assign v_1134 = ~v_837 & v_901;
assign v_1135 = v_901 & v_1133;
assign v_1136 = ~v_837 & v_1133;
assign v_1138 = ~v_838 & v_902;
assign v_1139 = v_902 & v_1137;
assign v_1140 = ~v_838 & v_1137;
assign v_1142 = ~v_839 & v_903;
assign v_1143 = v_903 & v_1141;
assign v_1144 = ~v_839 & v_1141;
assign v_1146 = ~v_840 & v_904;
assign v_1147 = v_904 & v_1145;
assign v_1148 = ~v_840 & v_1145;
assign v_1150 = ~v_841 & v_905;
assign v_1151 = v_905 & v_1149;
assign v_1152 = ~v_841 & v_1149;
assign v_1154 = ~v_842 & v_906;
assign v_1155 = v_906 & v_1153;
assign v_1156 = ~v_842 & v_1153;
assign v_1158 = ~v_843 & v_907;
assign v_1159 = v_907 & v_1157;
assign v_1160 = ~v_843 & v_1157;
assign v_1292 = ~v_1164 & v_1228;
assign v_1294 = ~v_1165 & v_1229;
assign v_1295 = v_1229 & v_1293;
assign v_1296 = ~v_1165 & v_1293;
assign v_1298 = ~v_1166 & v_1230;
assign v_1299 = v_1230 & v_1297;
assign v_1300 = ~v_1166 & v_1297;
assign v_1302 = ~v_1167 & v_1231;
assign v_1303 = v_1231 & v_1301;
assign v_1304 = ~v_1167 & v_1301;
assign v_1306 = ~v_1168 & v_1232;
assign v_1307 = v_1232 & v_1305;
assign v_1308 = ~v_1168 & v_1305;
assign v_1310 = ~v_1169 & v_1233;
assign v_1311 = v_1233 & v_1309;
assign v_1312 = ~v_1169 & v_1309;
assign v_1314 = ~v_1170 & v_1234;
assign v_1315 = v_1234 & v_1313;
assign v_1316 = ~v_1170 & v_1313;
assign v_1318 = ~v_1171 & v_1235;
assign v_1319 = v_1235 & v_1317;
assign v_1320 = ~v_1171 & v_1317;
assign v_1322 = ~v_1172 & v_1236;
assign v_1323 = v_1236 & v_1321;
assign v_1324 = ~v_1172 & v_1321;
assign v_1326 = ~v_1173 & v_1237;
assign v_1327 = v_1237 & v_1325;
assign v_1328 = ~v_1173 & v_1325;
assign v_1330 = ~v_1174 & v_1238;
assign v_1331 = v_1238 & v_1329;
assign v_1332 = ~v_1174 & v_1329;
assign v_1334 = ~v_1175 & v_1239;
assign v_1335 = v_1239 & v_1333;
assign v_1336 = ~v_1175 & v_1333;
assign v_1338 = ~v_1176 & v_1240;
assign v_1339 = v_1240 & v_1337;
assign v_1340 = ~v_1176 & v_1337;
assign v_1342 = ~v_1177 & v_1241;
assign v_1343 = v_1241 & v_1341;
assign v_1344 = ~v_1177 & v_1341;
assign v_1346 = ~v_1178 & v_1242;
assign v_1347 = v_1242 & v_1345;
assign v_1348 = ~v_1178 & v_1345;
assign v_1350 = ~v_1179 & v_1243;
assign v_1351 = v_1243 & v_1349;
assign v_1352 = ~v_1179 & v_1349;
assign v_1354 = ~v_1180 & v_1244;
assign v_1355 = v_1244 & v_1353;
assign v_1356 = ~v_1180 & v_1353;
assign v_1358 = ~v_1181 & v_1245;
assign v_1359 = v_1245 & v_1357;
assign v_1360 = ~v_1181 & v_1357;
assign v_1362 = ~v_1182 & v_1246;
assign v_1363 = v_1246 & v_1361;
assign v_1364 = ~v_1182 & v_1361;
assign v_1366 = ~v_1183 & v_1247;
assign v_1367 = v_1247 & v_1365;
assign v_1368 = ~v_1183 & v_1365;
assign v_1370 = ~v_1184 & v_1248;
assign v_1371 = v_1248 & v_1369;
assign v_1372 = ~v_1184 & v_1369;
assign v_1374 = ~v_1185 & v_1249;
assign v_1375 = v_1249 & v_1373;
assign v_1376 = ~v_1185 & v_1373;
assign v_1378 = ~v_1186 & v_1250;
assign v_1379 = v_1250 & v_1377;
assign v_1380 = ~v_1186 & v_1377;
assign v_1382 = ~v_1187 & v_1251;
assign v_1383 = v_1251 & v_1381;
assign v_1384 = ~v_1187 & v_1381;
assign v_1386 = ~v_1188 & v_1252;
assign v_1387 = v_1252 & v_1385;
assign v_1388 = ~v_1188 & v_1385;
assign v_1390 = ~v_1189 & v_1253;
assign v_1391 = v_1253 & v_1389;
assign v_1392 = ~v_1189 & v_1389;
assign v_1394 = ~v_1190 & v_1254;
assign v_1395 = v_1254 & v_1393;
assign v_1396 = ~v_1190 & v_1393;
assign v_1398 = ~v_1191 & v_1255;
assign v_1399 = v_1255 & v_1397;
assign v_1400 = ~v_1191 & v_1397;
assign v_1402 = ~v_1192 & v_1256;
assign v_1403 = v_1256 & v_1401;
assign v_1404 = ~v_1192 & v_1401;
assign v_1406 = ~v_1193 & v_1257;
assign v_1407 = v_1257 & v_1405;
assign v_1408 = ~v_1193 & v_1405;
assign v_1410 = ~v_1194 & v_1258;
assign v_1411 = v_1258 & v_1409;
assign v_1412 = ~v_1194 & v_1409;
assign v_1414 = ~v_1195 & v_1259;
assign v_1415 = v_1259 & v_1413;
assign v_1416 = ~v_1195 & v_1413;
assign v_1418 = ~v_1196 & v_1260;
assign v_1419 = v_1260 & v_1417;
assign v_1420 = ~v_1196 & v_1417;
assign v_1422 = ~v_1197 & v_1261;
assign v_1423 = v_1261 & v_1421;
assign v_1424 = ~v_1197 & v_1421;
assign v_1426 = ~v_1198 & v_1262;
assign v_1427 = v_1262 & v_1425;
assign v_1428 = ~v_1198 & v_1425;
assign v_1430 = ~v_1199 & v_1263;
assign v_1431 = v_1263 & v_1429;
assign v_1432 = ~v_1199 & v_1429;
assign v_1434 = ~v_1200 & v_1264;
assign v_1435 = v_1264 & v_1433;
assign v_1436 = ~v_1200 & v_1433;
assign v_1438 = ~v_1201 & v_1265;
assign v_1439 = v_1265 & v_1437;
assign v_1440 = ~v_1201 & v_1437;
assign v_1442 = ~v_1202 & v_1266;
assign v_1443 = v_1266 & v_1441;
assign v_1444 = ~v_1202 & v_1441;
assign v_1446 = ~v_1203 & v_1267;
assign v_1447 = v_1267 & v_1445;
assign v_1448 = ~v_1203 & v_1445;
assign v_1450 = ~v_1204 & v_1268;
assign v_1451 = v_1268 & v_1449;
assign v_1452 = ~v_1204 & v_1449;
assign v_1454 = ~v_1205 & v_1269;
assign v_1455 = v_1269 & v_1453;
assign v_1456 = ~v_1205 & v_1453;
assign v_1458 = ~v_1206 & v_1270;
assign v_1459 = v_1270 & v_1457;
assign v_1460 = ~v_1206 & v_1457;
assign v_1462 = ~v_1207 & v_1271;
assign v_1463 = v_1271 & v_1461;
assign v_1464 = ~v_1207 & v_1461;
assign v_1466 = ~v_1208 & v_1272;
assign v_1467 = v_1272 & v_1465;
assign v_1468 = ~v_1208 & v_1465;
assign v_1470 = ~v_1209 & v_1273;
assign v_1471 = v_1273 & v_1469;
assign v_1472 = ~v_1209 & v_1469;
assign v_1474 = ~v_1210 & v_1274;
assign v_1475 = v_1274 & v_1473;
assign v_1476 = ~v_1210 & v_1473;
assign v_1478 = ~v_1211 & v_1275;
assign v_1479 = v_1275 & v_1477;
assign v_1480 = ~v_1211 & v_1477;
assign v_1482 = ~v_1212 & v_1276;
assign v_1483 = v_1276 & v_1481;
assign v_1484 = ~v_1212 & v_1481;
assign v_1486 = ~v_1213 & v_1277;
assign v_1487 = v_1277 & v_1485;
assign v_1488 = ~v_1213 & v_1485;
assign v_1490 = ~v_1214 & v_1278;
assign v_1491 = v_1278 & v_1489;
assign v_1492 = ~v_1214 & v_1489;
assign v_1494 = ~v_1215 & v_1279;
assign v_1495 = v_1279 & v_1493;
assign v_1496 = ~v_1215 & v_1493;
assign v_1498 = ~v_1216 & v_1280;
assign v_1499 = v_1280 & v_1497;
assign v_1500 = ~v_1216 & v_1497;
assign v_1502 = ~v_1217 & v_1281;
assign v_1503 = v_1281 & v_1501;
assign v_1504 = ~v_1217 & v_1501;
assign v_1506 = ~v_1218 & v_1282;
assign v_1507 = v_1282 & v_1505;
assign v_1508 = ~v_1218 & v_1505;
assign v_1510 = ~v_1219 & v_1283;
assign v_1511 = v_1283 & v_1509;
assign v_1512 = ~v_1219 & v_1509;
assign v_1514 = ~v_1220 & v_1284;
assign v_1515 = v_1284 & v_1513;
assign v_1516 = ~v_1220 & v_1513;
assign v_1518 = ~v_1221 & v_1285;
assign v_1519 = v_1285 & v_1517;
assign v_1520 = ~v_1221 & v_1517;
assign v_1522 = ~v_1222 & v_1286;
assign v_1523 = v_1286 & v_1521;
assign v_1524 = ~v_1222 & v_1521;
assign v_1526 = ~v_1223 & v_1287;
assign v_1527 = v_1287 & v_1525;
assign v_1528 = ~v_1223 & v_1525;
assign v_1530 = ~v_1224 & v_1288;
assign v_1531 = v_1288 & v_1529;
assign v_1532 = ~v_1224 & v_1529;
assign v_1534 = ~v_1225 & v_1289;
assign v_1535 = v_1289 & v_1533;
assign v_1536 = ~v_1225 & v_1533;
assign v_1538 = ~v_1226 & v_1290;
assign v_1539 = v_1290 & v_1537;
assign v_1540 = ~v_1226 & v_1537;
assign v_1542 = ~v_1227 & v_1291;
assign v_1543 = v_1291 & v_1541;
assign v_1544 = ~v_1227 & v_1541;
assign v_1548 = ~v_1161 & ~v_1545;
assign v_1613 = v_1888 & v_1889 & v_1890;
assign v_1678 = v_1904 & v_1905 & v_1906;
assign v_1743 = v_1920 & v_1921 & v_1922;
assign v_1808 = v_1936 & v_1937 & v_1938;
assign v_1809 = ~v_519 & ~v_520 & ~v_521 & ~v_522 & ~v_523;
assign v_1810 = ~v_524 & ~v_525 & ~v_526 & ~v_527 & ~v_528;
assign v_1811 = ~v_529 & ~v_530 & ~v_531 & ~v_532 & ~v_533;
assign v_1812 = ~v_534 & ~v_535 & ~v_536 & ~v_537 & ~v_538;
assign v_1813 = ~v_539 & ~v_540 & ~v_541 & ~v_542 & ~v_543;
assign v_1814 = ~v_544 & ~v_545 & ~v_546 & ~v_547 & ~v_548;
assign v_1815 = ~v_549 & ~v_550 & ~v_551 & ~v_552 & ~v_553;
assign v_1816 = ~v_554 & ~v_555 & ~v_556 & ~v_557 & ~v_558;
assign v_1817 = ~v_559 & ~v_560 & ~v_561 & ~v_562 & ~v_563;
assign v_1818 = ~v_564 & ~v_565 & ~v_566 & ~v_567 & ~v_568;
assign v_1819 = ~v_569 & ~v_570 & ~v_571 & ~v_572 & ~v_573;
assign v_1820 = ~v_574 & ~v_575 & ~v_576 & ~v_577 & ~v_578;
assign v_1821 = ~v_579 & ~v_580 & ~v_581 & ~v_582;
assign v_1822 = v_1809 & v_1810 & v_1811 & v_1812 & v_1813;
assign v_1823 = v_1814 & v_1815 & v_1816 & v_1817 & v_1818;
assign v_1824 = v_1819 & v_1820 & v_1821;
assign v_1825 = ~v_584 & ~v_585 & ~v_586 & ~v_587 & ~v_588;
assign v_1826 = ~v_589 & ~v_590 & ~v_591 & ~v_592 & ~v_593;
assign v_1827 = ~v_594 & ~v_595 & ~v_596 & ~v_597 & ~v_598;
assign v_1828 = ~v_599 & ~v_600 & ~v_601 & ~v_602 & ~v_603;
assign v_1829 = ~v_604 & ~v_605 & ~v_606 & ~v_607 & ~v_608;
assign v_1830 = ~v_609 & ~v_610 & ~v_611 & ~v_612 & ~v_613;
assign v_1831 = ~v_614 & ~v_615 & ~v_616 & ~v_617 & ~v_618;
assign v_1832 = ~v_619 & ~v_620 & ~v_621 & ~v_622 & ~v_623;
assign v_1833 = ~v_624 & ~v_625 & ~v_626 & ~v_627 & ~v_628;
assign v_1834 = ~v_629 & ~v_630 & ~v_631 & ~v_632 & ~v_633;
assign v_1835 = ~v_634 & ~v_635 & ~v_636 & ~v_637 & ~v_638;
assign v_1836 = ~v_639 & ~v_640 & ~v_641 & ~v_642 & ~v_643;
assign v_1837 = ~v_644 & ~v_645 & ~v_646 & ~v_647;
assign v_1838 = v_1825 & v_1826 & v_1827 & v_1828 & v_1829;
assign v_1839 = v_1830 & v_1831 & v_1832 & v_1833 & v_1834;
assign v_1840 = v_1835 & v_1836 & v_1837;
assign v_1841 = ~v_649 & ~v_650 & ~v_651 & ~v_652 & ~v_653;
assign v_1842 = ~v_654 & ~v_655 & ~v_656 & ~v_657 & ~v_658;
assign v_1843 = ~v_659 & ~v_660 & ~v_661 & ~v_662 & ~v_663;
assign v_1844 = ~v_664 & ~v_665 & ~v_666 & ~v_667 & ~v_668;
assign v_1845 = ~v_669 & ~v_670 & ~v_671 & ~v_672 & ~v_673;
assign v_1846 = ~v_674 & ~v_675 & ~v_676 & ~v_677 & ~v_678;
assign v_1847 = ~v_679 & ~v_680 & ~v_681 & ~v_682 & ~v_683;
assign v_1848 = ~v_684 & ~v_685 & ~v_686 & ~v_687 & ~v_688;
assign v_1849 = ~v_689 & ~v_690 & ~v_691 & ~v_692 & ~v_693;
assign v_1850 = ~v_694 & ~v_695 & ~v_696 & ~v_697 & ~v_698;
assign v_1851 = ~v_699 & ~v_700 & ~v_701 & ~v_702 & ~v_703;
assign v_1852 = ~v_704 & ~v_705 & ~v_706 & ~v_707 & ~v_708;
assign v_1853 = ~v_709 & ~v_710 & ~v_711 & ~v_712;
assign v_1854 = v_1841 & v_1842 & v_1843 & v_1844 & v_1845;
assign v_1855 = v_1846 & v_1847 & v_1848 & v_1849 & v_1850;
assign v_1856 = v_1851 & v_1852 & v_1853;
assign v_1857 = ~v_714 & ~v_715 & ~v_716 & ~v_717 & ~v_718;
assign v_1858 = ~v_719 & ~v_720 & ~v_721 & ~v_722 & ~v_723;
assign v_1859 = ~v_724 & ~v_725 & ~v_726 & ~v_727 & ~v_728;
assign v_1860 = ~v_729 & ~v_730 & ~v_731 & ~v_732 & ~v_733;
assign v_1861 = ~v_734 & ~v_735 & ~v_736 & ~v_737 & ~v_738;
assign v_1862 = ~v_739 & ~v_740 & ~v_741 & ~v_742 & ~v_743;
assign v_1863 = ~v_744 & ~v_745 & ~v_746 & ~v_747 & ~v_748;
assign v_1864 = ~v_749 & ~v_750 & ~v_751 & ~v_752 & ~v_753;
assign v_1865 = ~v_754 & ~v_755 & ~v_756 & ~v_757 & ~v_758;
assign v_1866 = ~v_759 & ~v_760 & ~v_761 & ~v_762 & ~v_763;
assign v_1867 = ~v_764 & ~v_765 & ~v_766 & ~v_767 & ~v_768;
assign v_1868 = ~v_769 & ~v_770 & ~v_771 & ~v_772 & ~v_773;
assign v_1869 = ~v_774 & ~v_775 & ~v_776 & ~v_777;
assign v_1870 = v_1857 & v_1858 & v_1859 & v_1860 & v_1861;
assign v_1871 = v_1862 & v_1863 & v_1864 & v_1865 & v_1866;
assign v_1872 = v_1867 & v_1868 & v_1869;
assign v_1873 = v_448 & v_516 & v_583 & v_648 & v_713;
assign v_1874 = v_778;
assign v_1875 = ~v_1549 & ~v_1550 & ~v_1551 & ~v_1552 & ~v_1553;
assign v_1876 = ~v_1554 & ~v_1555 & ~v_1556 & ~v_1557 & ~v_1558;
assign v_1877 = ~v_1559 & ~v_1560 & ~v_1561 & ~v_1562 & ~v_1563;
assign v_1878 = ~v_1564 & ~v_1565 & ~v_1566 & ~v_1567 & ~v_1568;
assign v_1879 = ~v_1569 & ~v_1570 & ~v_1571 & ~v_1572 & ~v_1573;
assign v_1880 = ~v_1574 & ~v_1575 & ~v_1576 & ~v_1577 & ~v_1578;
assign v_1881 = ~v_1579 & ~v_1580 & ~v_1581 & ~v_1582 & ~v_1583;
assign v_1882 = ~v_1584 & ~v_1585 & ~v_1586 & ~v_1587 & ~v_1588;
assign v_1883 = ~v_1589 & ~v_1590 & ~v_1591 & ~v_1592 & ~v_1593;
assign v_1884 = ~v_1594 & ~v_1595 & ~v_1596 & ~v_1597 & ~v_1598;
assign v_1885 = ~v_1599 & ~v_1600 & ~v_1601 & ~v_1602 & ~v_1603;
assign v_1886 = ~v_1604 & ~v_1605 & ~v_1606 & ~v_1607 & ~v_1608;
assign v_1887 = ~v_1609 & ~v_1610 & ~v_1611 & ~v_1612;
assign v_1888 = v_1875 & v_1876 & v_1877 & v_1878 & v_1879;
assign v_1889 = v_1880 & v_1881 & v_1882 & v_1883 & v_1884;
assign v_1890 = v_1885 & v_1886 & v_1887;
assign v_1891 = ~v_1614 & ~v_1615 & ~v_1616 & ~v_1617 & ~v_1618;
assign v_1892 = ~v_1619 & ~v_1620 & ~v_1621 & ~v_1622 & ~v_1623;
assign v_1893 = ~v_1624 & ~v_1625 & ~v_1626 & ~v_1627 & ~v_1628;
assign v_1894 = ~v_1629 & ~v_1630 & ~v_1631 & ~v_1632 & ~v_1633;
assign v_1895 = ~v_1634 & ~v_1635 & ~v_1636 & ~v_1637 & ~v_1638;
assign v_1896 = ~v_1639 & ~v_1640 & ~v_1641 & ~v_1642 & ~v_1643;
assign v_1897 = ~v_1644 & ~v_1645 & ~v_1646 & ~v_1647 & ~v_1648;
assign v_1898 = ~v_1649 & ~v_1650 & ~v_1651 & ~v_1652 & ~v_1653;
assign v_1899 = ~v_1654 & ~v_1655 & ~v_1656 & ~v_1657 & ~v_1658;
assign v_1900 = ~v_1659 & ~v_1660 & ~v_1661 & ~v_1662 & ~v_1663;
assign v_1901 = ~v_1664 & ~v_1665 & ~v_1666 & ~v_1667 & ~v_1668;
assign v_1902 = ~v_1669 & ~v_1670 & ~v_1671 & ~v_1672 & ~v_1673;
assign v_1903 = ~v_1674 & ~v_1675 & ~v_1676 & ~v_1677;
assign v_1904 = v_1891 & v_1892 & v_1893 & v_1894 & v_1895;
assign v_1905 = v_1896 & v_1897 & v_1898 & v_1899 & v_1900;
assign v_1906 = v_1901 & v_1902 & v_1903;
assign v_1907 = ~v_1679 & ~v_1680 & ~v_1681 & ~v_1682 & ~v_1683;
assign v_1908 = ~v_1684 & ~v_1685 & ~v_1686 & ~v_1687 & ~v_1688;
assign v_1909 = ~v_1689 & ~v_1690 & ~v_1691 & ~v_1692 & ~v_1693;
assign v_1910 = ~v_1694 & ~v_1695 & ~v_1696 & ~v_1697 & ~v_1698;
assign v_1911 = ~v_1699 & ~v_1700 & ~v_1701 & ~v_1702 & ~v_1703;
assign v_1912 = ~v_1704 & ~v_1705 & ~v_1706 & ~v_1707 & ~v_1708;
assign v_1913 = ~v_1709 & ~v_1710 & ~v_1711 & ~v_1712 & ~v_1713;
assign v_1914 = ~v_1714 & ~v_1715 & ~v_1716 & ~v_1717 & ~v_1718;
assign v_1915 = ~v_1719 & ~v_1720 & ~v_1721 & ~v_1722 & ~v_1723;
assign v_1916 = ~v_1724 & ~v_1725 & ~v_1726 & ~v_1727 & ~v_1728;
assign v_1917 = ~v_1729 & ~v_1730 & ~v_1731 & ~v_1732 & ~v_1733;
assign v_1918 = ~v_1734 & ~v_1735 & ~v_1736 & ~v_1737 & ~v_1738;
assign v_1919 = ~v_1739 & ~v_1740 & ~v_1741 & ~v_1742;
assign v_1920 = v_1907 & v_1908 & v_1909 & v_1910 & v_1911;
assign v_1921 = v_1912 & v_1913 & v_1914 & v_1915 & v_1916;
assign v_1922 = v_1917 & v_1918 & v_1919;
assign v_1923 = ~v_1744 & ~v_1745 & ~v_1746 & ~v_1747 & ~v_1748;
assign v_1924 = ~v_1749 & ~v_1750 & ~v_1751 & ~v_1752 & ~v_1753;
assign v_1925 = ~v_1754 & ~v_1755 & ~v_1756 & ~v_1757 & ~v_1758;
assign v_1926 = ~v_1759 & ~v_1760 & ~v_1761 & ~v_1762 & ~v_1763;
assign v_1927 = ~v_1764 & ~v_1765 & ~v_1766 & ~v_1767 & ~v_1768;
assign v_1928 = ~v_1769 & ~v_1770 & ~v_1771 & ~v_1772 & ~v_1773;
assign v_1929 = ~v_1774 & ~v_1775 & ~v_1776 & ~v_1777 & ~v_1778;
assign v_1930 = ~v_1779 & ~v_1780 & ~v_1781 & ~v_1782 & ~v_1783;
assign v_1931 = ~v_1784 & ~v_1785 & ~v_1786 & ~v_1787 & ~v_1788;
assign v_1932 = ~v_1789 & ~v_1790 & ~v_1791 & ~v_1792 & ~v_1793;
assign v_1933 = ~v_1794 & ~v_1795 & ~v_1796 & ~v_1797 & ~v_1798;
assign v_1934 = ~v_1799 & ~v_1800 & ~v_1801 & ~v_1802 & ~v_1803;
assign v_1935 = ~v_1804 & ~v_1805 & ~v_1806 & ~v_1807;
assign v_1936 = v_1923 & v_1924 & v_1925 & v_1926 & v_1927;
assign v_1937 = v_1928 & v_1929 & v_1930 & v_1931 & v_1932;
assign v_1938 = v_1933 & v_1934 & v_1935;
assign v_515 = v_1952 | v_1953 | v_1954;
assign v_516 = v_514 | ~v_515;
assign v_909 = ~v_780 | v_844 | v_908;
assign v_913 = v_910 | v_911 | v_912;
assign v_917 = v_914 | v_915 | v_916;
assign v_921 = v_918 | v_919 | v_920;
assign v_925 = v_922 | v_923 | v_924;
assign v_929 = v_926 | v_927 | v_928;
assign v_933 = v_930 | v_931 | v_932;
assign v_937 = v_934 | v_935 | v_936;
assign v_941 = v_938 | v_939 | v_940;
assign v_945 = v_942 | v_943 | v_944;
assign v_949 = v_946 | v_947 | v_948;
assign v_953 = v_950 | v_951 | v_952;
assign v_957 = v_954 | v_955 | v_956;
assign v_961 = v_958 | v_959 | v_960;
assign v_965 = v_962 | v_963 | v_964;
assign v_969 = v_966 | v_967 | v_968;
assign v_973 = v_970 | v_971 | v_972;
assign v_977 = v_974 | v_975 | v_976;
assign v_981 = v_978 | v_979 | v_980;
assign v_985 = v_982 | v_983 | v_984;
assign v_989 = v_986 | v_987 | v_988;
assign v_993 = v_990 | v_991 | v_992;
assign v_997 = v_994 | v_995 | v_996;
assign v_1001 = v_998 | v_999 | v_1000;
assign v_1005 = v_1002 | v_1003 | v_1004;
assign v_1009 = v_1006 | v_1007 | v_1008;
assign v_1013 = v_1010 | v_1011 | v_1012;
assign v_1017 = v_1014 | v_1015 | v_1016;
assign v_1021 = v_1018 | v_1019 | v_1020;
assign v_1025 = v_1022 | v_1023 | v_1024;
assign v_1029 = v_1026 | v_1027 | v_1028;
assign v_1033 = v_1030 | v_1031 | v_1032;
assign v_1037 = v_1034 | v_1035 | v_1036;
assign v_1041 = v_1038 | v_1039 | v_1040;
assign v_1045 = v_1042 | v_1043 | v_1044;
assign v_1049 = v_1046 | v_1047 | v_1048;
assign v_1053 = v_1050 | v_1051 | v_1052;
assign v_1057 = v_1054 | v_1055 | v_1056;
assign v_1061 = v_1058 | v_1059 | v_1060;
assign v_1065 = v_1062 | v_1063 | v_1064;
assign v_1069 = v_1066 | v_1067 | v_1068;
assign v_1073 = v_1070 | v_1071 | v_1072;
assign v_1077 = v_1074 | v_1075 | v_1076;
assign v_1081 = v_1078 | v_1079 | v_1080;
assign v_1085 = v_1082 | v_1083 | v_1084;
assign v_1089 = v_1086 | v_1087 | v_1088;
assign v_1093 = v_1090 | v_1091 | v_1092;
assign v_1097 = v_1094 | v_1095 | v_1096;
assign v_1101 = v_1098 | v_1099 | v_1100;
assign v_1105 = v_1102 | v_1103 | v_1104;
assign v_1109 = v_1106 | v_1107 | v_1108;
assign v_1113 = v_1110 | v_1111 | v_1112;
assign v_1117 = v_1114 | v_1115 | v_1116;
assign v_1121 = v_1118 | v_1119 | v_1120;
assign v_1125 = v_1122 | v_1123 | v_1124;
assign v_1129 = v_1126 | v_1127 | v_1128;
assign v_1133 = v_1130 | v_1131 | v_1132;
assign v_1137 = v_1134 | v_1135 | v_1136;
assign v_1141 = v_1138 | v_1139 | v_1140;
assign v_1145 = v_1142 | v_1143 | v_1144;
assign v_1149 = v_1146 | v_1147 | v_1148;
assign v_1153 = v_1150 | v_1151 | v_1152;
assign v_1157 = v_1154 | v_1155 | v_1156;
assign v_1161 = v_1158 | v_1159 | v_1160;
assign v_1293 = ~v_1164 | v_1228 | v_1292;
assign v_1297 = v_1294 | v_1295 | v_1296;
assign v_1301 = v_1298 | v_1299 | v_1300;
assign v_1305 = v_1302 | v_1303 | v_1304;
assign v_1309 = v_1306 | v_1307 | v_1308;
assign v_1313 = v_1310 | v_1311 | v_1312;
assign v_1317 = v_1314 | v_1315 | v_1316;
assign v_1321 = v_1318 | v_1319 | v_1320;
assign v_1325 = v_1322 | v_1323 | v_1324;
assign v_1329 = v_1326 | v_1327 | v_1328;
assign v_1333 = v_1330 | v_1331 | v_1332;
assign v_1337 = v_1334 | v_1335 | v_1336;
assign v_1341 = v_1338 | v_1339 | v_1340;
assign v_1345 = v_1342 | v_1343 | v_1344;
assign v_1349 = v_1346 | v_1347 | v_1348;
assign v_1353 = v_1350 | v_1351 | v_1352;
assign v_1357 = v_1354 | v_1355 | v_1356;
assign v_1361 = v_1358 | v_1359 | v_1360;
assign v_1365 = v_1362 | v_1363 | v_1364;
assign v_1369 = v_1366 | v_1367 | v_1368;
assign v_1373 = v_1370 | v_1371 | v_1372;
assign v_1377 = v_1374 | v_1375 | v_1376;
assign v_1381 = v_1378 | v_1379 | v_1380;
assign v_1385 = v_1382 | v_1383 | v_1384;
assign v_1389 = v_1386 | v_1387 | v_1388;
assign v_1393 = v_1390 | v_1391 | v_1392;
assign v_1397 = v_1394 | v_1395 | v_1396;
assign v_1401 = v_1398 | v_1399 | v_1400;
assign v_1405 = v_1402 | v_1403 | v_1404;
assign v_1409 = v_1406 | v_1407 | v_1408;
assign v_1413 = v_1410 | v_1411 | v_1412;
assign v_1417 = v_1414 | v_1415 | v_1416;
assign v_1421 = v_1418 | v_1419 | v_1420;
assign v_1425 = v_1422 | v_1423 | v_1424;
assign v_1429 = v_1426 | v_1427 | v_1428;
assign v_1433 = v_1430 | v_1431 | v_1432;
assign v_1437 = v_1434 | v_1435 | v_1436;
assign v_1441 = v_1438 | v_1439 | v_1440;
assign v_1445 = v_1442 | v_1443 | v_1444;
assign v_1449 = v_1446 | v_1447 | v_1448;
assign v_1453 = v_1450 | v_1451 | v_1452;
assign v_1457 = v_1454 | v_1455 | v_1456;
assign v_1461 = v_1458 | v_1459 | v_1460;
assign v_1465 = v_1462 | v_1463 | v_1464;
assign v_1469 = v_1466 | v_1467 | v_1468;
assign v_1473 = v_1470 | v_1471 | v_1472;
assign v_1477 = v_1474 | v_1475 | v_1476;
assign v_1481 = v_1478 | v_1479 | v_1480;
assign v_1485 = v_1482 | v_1483 | v_1484;
assign v_1489 = v_1486 | v_1487 | v_1488;
assign v_1493 = v_1490 | v_1491 | v_1492;
assign v_1497 = v_1494 | v_1495 | v_1496;
assign v_1501 = v_1498 | v_1499 | v_1500;
assign v_1505 = v_1502 | v_1503 | v_1504;
assign v_1509 = v_1506 | v_1507 | v_1508;
assign v_1513 = v_1510 | v_1511 | v_1512;
assign v_1517 = v_1514 | v_1515 | v_1516;
assign v_1521 = v_1518 | v_1519 | v_1520;
assign v_1525 = v_1522 | v_1523 | v_1524;
assign v_1529 = v_1526 | v_1527 | v_1528;
assign v_1533 = v_1530 | v_1531 | v_1532;
assign v_1537 = v_1534 | v_1535 | v_1536;
assign v_1541 = v_1538 | v_1539 | v_1540;
assign v_1545 = v_1542 | v_1543 | v_1544;
assign v_1939 = v_451 | v_452 | v_453 | v_454 | v_455;
assign v_1940 = v_456 | v_457 | v_458 | v_459 | v_460;
assign v_1941 = v_461 | v_462 | v_463 | v_464 | v_465;
assign v_1942 = v_466 | v_467 | v_468 | v_469 | v_470;
assign v_1943 = v_471 | v_472 | v_473 | v_474 | v_475;
assign v_1944 = v_476 | v_477 | v_478 | v_479 | v_480;
assign v_1945 = v_481 | v_482 | v_483 | v_484 | v_485;
assign v_1946 = v_486 | v_487 | v_488 | v_489 | v_490;
assign v_1947 = v_491 | v_492 | v_493 | v_494 | v_495;
assign v_1948 = v_496 | v_497 | v_498 | v_499 | v_500;
assign v_1949 = v_501 | v_502 | v_503 | v_504 | v_505;
assign v_1950 = v_506 | v_507 | v_508 | v_509 | v_510;
assign v_1951 = v_511 | v_512 | v_513 | v_514;
assign v_1952 = v_1939 | v_1940 | v_1941 | v_1942 | v_1943;
assign v_1953 = v_1944 | v_1945 | v_1946 | v_1947 | v_1948;
assign v_1954 = v_1949 | v_1950 | v_1951;
assign v_448 = ~v_320 ^ v_447;
assign v_519 = v_1 ^ v_257;
assign v_520 = v_2 ^ v_258;
assign v_521 = v_3 ^ v_259;
assign v_522 = v_4 ^ v_260;
assign v_523 = v_5 ^ v_261;
assign v_524 = v_6 ^ v_262;
assign v_525 = v_7 ^ v_263;
assign v_526 = v_8 ^ v_264;
assign v_527 = v_9 ^ v_265;
assign v_528 = v_10 ^ v_266;
assign v_529 = v_11 ^ v_267;
assign v_530 = v_12 ^ v_268;
assign v_531 = v_13 ^ v_269;
assign v_532 = v_14 ^ v_270;
assign v_533 = v_15 ^ v_271;
assign v_534 = v_16 ^ v_272;
assign v_535 = v_17 ^ v_273;
assign v_536 = v_18 ^ v_274;
assign v_537 = v_19 ^ v_275;
assign v_538 = v_20 ^ v_276;
assign v_539 = v_21 ^ v_277;
assign v_540 = v_22 ^ v_278;
assign v_541 = v_23 ^ v_279;
assign v_542 = v_24 ^ v_280;
assign v_543 = v_25 ^ v_281;
assign v_544 = v_26 ^ v_282;
assign v_545 = v_27 ^ v_283;
assign v_546 = v_28 ^ v_284;
assign v_547 = v_29 ^ v_285;
assign v_548 = v_30 ^ v_286;
assign v_549 = v_31 ^ v_287;
assign v_550 = v_32 ^ v_288;
assign v_551 = v_33 ^ v_289;
assign v_552 = v_34 ^ v_290;
assign v_553 = v_35 ^ v_291;
assign v_554 = v_36 ^ v_292;
assign v_555 = v_37 ^ v_293;
assign v_556 = v_38 ^ v_294;
assign v_557 = v_39 ^ v_295;
assign v_558 = v_40 ^ v_296;
assign v_559 = v_41 ^ v_297;
assign v_560 = v_42 ^ v_298;
assign v_561 = v_43 ^ v_299;
assign v_562 = v_44 ^ v_300;
assign v_563 = v_45 ^ v_301;
assign v_564 = v_46 ^ v_302;
assign v_565 = v_47 ^ v_303;
assign v_566 = v_48 ^ v_304;
assign v_567 = v_49 ^ v_305;
assign v_568 = v_50 ^ v_306;
assign v_569 = v_51 ^ v_307;
assign v_570 = v_52 ^ v_308;
assign v_571 = v_53 ^ v_309;
assign v_572 = v_54 ^ v_310;
assign v_573 = v_55 ^ v_311;
assign v_574 = v_56 ^ v_312;
assign v_575 = v_57 ^ v_313;
assign v_576 = v_58 ^ v_314;
assign v_577 = v_59 ^ v_315;
assign v_578 = v_60 ^ v_316;
assign v_579 = v_61 ^ v_317;
assign v_580 = v_62 ^ v_318;
assign v_581 = v_63 ^ v_319;
assign v_582 = v_64 ^ v_320;
assign v_584 = v_129 ^ v_257;
assign v_585 = v_130 ^ v_258;
assign v_586 = v_131 ^ v_259;
assign v_587 = v_132 ^ v_260;
assign v_588 = v_133 ^ v_261;
assign v_589 = v_134 ^ v_262;
assign v_590 = v_135 ^ v_263;
assign v_591 = v_136 ^ v_264;
assign v_592 = v_137 ^ v_265;
assign v_593 = v_138 ^ v_266;
assign v_594 = v_139 ^ v_267;
assign v_595 = v_140 ^ v_268;
assign v_596 = v_141 ^ v_269;
assign v_597 = v_142 ^ v_270;
assign v_598 = v_143 ^ v_271;
assign v_599 = v_144 ^ v_272;
assign v_600 = v_145 ^ v_273;
assign v_601 = v_146 ^ v_274;
assign v_602 = v_147 ^ v_275;
assign v_603 = v_148 ^ v_276;
assign v_604 = v_149 ^ v_277;
assign v_605 = v_150 ^ v_278;
assign v_606 = v_151 ^ v_279;
assign v_607 = v_152 ^ v_280;
assign v_608 = v_153 ^ v_281;
assign v_609 = v_154 ^ v_282;
assign v_610 = v_155 ^ v_283;
assign v_611 = v_156 ^ v_284;
assign v_612 = v_157 ^ v_285;
assign v_613 = v_158 ^ v_286;
assign v_614 = v_159 ^ v_287;
assign v_615 = v_160 ^ v_288;
assign v_616 = v_161 ^ v_289;
assign v_617 = v_162 ^ v_290;
assign v_618 = v_163 ^ v_291;
assign v_619 = v_164 ^ v_292;
assign v_620 = v_165 ^ v_293;
assign v_621 = v_166 ^ v_294;
assign v_622 = v_167 ^ v_295;
assign v_623 = v_168 ^ v_296;
assign v_624 = v_169 ^ v_297;
assign v_625 = v_170 ^ v_298;
assign v_626 = v_171 ^ v_299;
assign v_627 = v_172 ^ v_300;
assign v_628 = v_173 ^ v_301;
assign v_629 = v_174 ^ v_302;
assign v_630 = v_175 ^ v_303;
assign v_631 = v_176 ^ v_304;
assign v_632 = v_177 ^ v_305;
assign v_633 = v_178 ^ v_306;
assign v_634 = v_179 ^ v_307;
assign v_635 = v_180 ^ v_308;
assign v_636 = v_181 ^ v_309;
assign v_637 = v_182 ^ v_310;
assign v_638 = v_183 ^ v_311;
assign v_639 = v_184 ^ v_312;
assign v_640 = v_185 ^ v_313;
assign v_641 = v_186 ^ v_314;
assign v_642 = v_187 ^ v_315;
assign v_643 = v_188 ^ v_316;
assign v_644 = v_189 ^ v_317;
assign v_645 = v_190 ^ v_318;
assign v_646 = v_191 ^ v_319;
assign v_647 = v_192 ^ v_320;
assign v_649 = v_65 ^ v_451;
assign v_650 = v_66 ^ v_452;
assign v_651 = v_67 ^ v_453;
assign v_652 = v_68 ^ v_454;
assign v_653 = v_69 ^ v_455;
assign v_654 = v_70 ^ v_456;
assign v_655 = v_71 ^ v_457;
assign v_656 = v_72 ^ v_458;
assign v_657 = v_73 ^ v_459;
assign v_658 = v_74 ^ v_460;
assign v_659 = v_75 ^ v_461;
assign v_660 = v_76 ^ v_462;
assign v_661 = v_77 ^ v_463;
assign v_662 = v_78 ^ v_464;
assign v_663 = v_79 ^ v_465;
assign v_664 = v_80 ^ v_466;
assign v_665 = v_81 ^ v_467;
assign v_666 = v_82 ^ v_468;
assign v_667 = v_83 ^ v_469;
assign v_668 = v_84 ^ v_470;
assign v_669 = v_85 ^ v_471;
assign v_670 = v_86 ^ v_472;
assign v_671 = v_87 ^ v_473;
assign v_672 = v_88 ^ v_474;
assign v_673 = v_89 ^ v_475;
assign v_674 = v_90 ^ v_476;
assign v_675 = v_91 ^ v_477;
assign v_676 = v_92 ^ v_478;
assign v_677 = v_93 ^ v_479;
assign v_678 = v_94 ^ v_480;
assign v_679 = v_95 ^ v_481;
assign v_680 = v_96 ^ v_482;
assign v_681 = v_97 ^ v_483;
assign v_682 = v_98 ^ v_484;
assign v_683 = v_99 ^ v_485;
assign v_684 = v_100 ^ v_486;
assign v_685 = v_101 ^ v_487;
assign v_686 = v_102 ^ v_488;
assign v_687 = v_103 ^ v_489;
assign v_688 = v_104 ^ v_490;
assign v_689 = v_105 ^ v_491;
assign v_690 = v_106 ^ v_492;
assign v_691 = v_107 ^ v_493;
assign v_692 = v_108 ^ v_494;
assign v_693 = v_109 ^ v_495;
assign v_694 = v_110 ^ v_496;
assign v_695 = v_111 ^ v_497;
assign v_696 = v_112 ^ v_498;
assign v_697 = v_113 ^ v_499;
assign v_698 = v_114 ^ v_500;
assign v_699 = v_115 ^ v_501;
assign v_700 = v_116 ^ v_502;
assign v_701 = v_117 ^ v_503;
assign v_702 = v_118 ^ v_504;
assign v_703 = v_119 ^ v_505;
assign v_704 = v_120 ^ v_506;
assign v_705 = v_121 ^ v_507;
assign v_706 = v_122 ^ v_508;
assign v_707 = v_123 ^ v_509;
assign v_708 = v_124 ^ v_510;
assign v_709 = v_125 ^ v_511;
assign v_710 = v_126 ^ v_512;
assign v_711 = v_127 ^ v_513;
assign v_712 = v_128 ^ v_514;
assign v_714 = v_193 ^ v_451;
assign v_715 = v_194 ^ v_452;
assign v_716 = v_195 ^ v_453;
assign v_717 = v_196 ^ v_454;
assign v_718 = v_197 ^ v_455;
assign v_719 = v_198 ^ v_456;
assign v_720 = v_199 ^ v_457;
assign v_721 = v_200 ^ v_458;
assign v_722 = v_201 ^ v_459;
assign v_723 = v_202 ^ v_460;
assign v_724 = v_203 ^ v_461;
assign v_725 = v_204 ^ v_462;
assign v_726 = v_205 ^ v_463;
assign v_727 = v_206 ^ v_464;
assign v_728 = v_207 ^ v_465;
assign v_729 = v_208 ^ v_466;
assign v_730 = v_209 ^ v_467;
assign v_731 = v_210 ^ v_468;
assign v_732 = v_211 ^ v_469;
assign v_733 = v_212 ^ v_470;
assign v_734 = v_213 ^ v_471;
assign v_735 = v_214 ^ v_472;
assign v_736 = v_215 ^ v_473;
assign v_737 = v_216 ^ v_474;
assign v_738 = v_217 ^ v_475;
assign v_739 = v_218 ^ v_476;
assign v_740 = v_219 ^ v_477;
assign v_741 = v_220 ^ v_478;
assign v_742 = v_221 ^ v_479;
assign v_743 = v_222 ^ v_480;
assign v_744 = v_223 ^ v_481;
assign v_745 = v_224 ^ v_482;
assign v_746 = v_225 ^ v_483;
assign v_747 = v_226 ^ v_484;
assign v_748 = v_227 ^ v_485;
assign v_749 = v_228 ^ v_486;
assign v_750 = v_229 ^ v_487;
assign v_751 = v_230 ^ v_488;
assign v_752 = v_231 ^ v_489;
assign v_753 = v_232 ^ v_490;
assign v_754 = v_233 ^ v_491;
assign v_755 = v_234 ^ v_492;
assign v_756 = v_235 ^ v_493;
assign v_757 = v_236 ^ v_494;
assign v_758 = v_237 ^ v_495;
assign v_759 = v_238 ^ v_496;
assign v_760 = v_239 ^ v_497;
assign v_761 = v_240 ^ v_498;
assign v_762 = v_241 ^ v_499;
assign v_763 = v_242 ^ v_500;
assign v_764 = v_243 ^ v_501;
assign v_765 = v_244 ^ v_502;
assign v_766 = v_245 ^ v_503;
assign v_767 = v_246 ^ v_504;
assign v_768 = v_247 ^ v_505;
assign v_769 = v_248 ^ v_506;
assign v_770 = v_249 ^ v_507;
assign v_771 = v_250 ^ v_508;
assign v_772 = v_251 ^ v_509;
assign v_773 = v_252 ^ v_510;
assign v_774 = v_253 ^ v_511;
assign v_775 = v_254 ^ v_512;
assign v_776 = v_255 ^ v_513;
assign v_777 = v_256 ^ v_514;
assign v_1549 = v_1 ^ v_129;
assign v_1550 = v_2 ^ v_130;
assign v_1551 = v_3 ^ v_131;
assign v_1552 = v_4 ^ v_132;
assign v_1553 = v_5 ^ v_133;
assign v_1554 = v_6 ^ v_134;
assign v_1555 = v_7 ^ v_135;
assign v_1556 = v_8 ^ v_136;
assign v_1557 = v_9 ^ v_137;
assign v_1558 = v_10 ^ v_138;
assign v_1559 = v_11 ^ v_139;
assign v_1560 = v_12 ^ v_140;
assign v_1561 = v_13 ^ v_141;
assign v_1562 = v_14 ^ v_142;
assign v_1563 = v_15 ^ v_143;
assign v_1564 = v_16 ^ v_144;
assign v_1565 = v_17 ^ v_145;
assign v_1566 = v_18 ^ v_146;
assign v_1567 = v_19 ^ v_147;
assign v_1568 = v_20 ^ v_148;
assign v_1569 = v_21 ^ v_149;
assign v_1570 = v_22 ^ v_150;
assign v_1571 = v_23 ^ v_151;
assign v_1572 = v_24 ^ v_152;
assign v_1573 = v_25 ^ v_153;
assign v_1574 = v_26 ^ v_154;
assign v_1575 = v_27 ^ v_155;
assign v_1576 = v_28 ^ v_156;
assign v_1577 = v_29 ^ v_157;
assign v_1578 = v_30 ^ v_158;
assign v_1579 = v_31 ^ v_159;
assign v_1580 = v_32 ^ v_160;
assign v_1581 = v_33 ^ v_161;
assign v_1582 = v_34 ^ v_162;
assign v_1583 = v_35 ^ v_163;
assign v_1584 = v_36 ^ v_164;
assign v_1585 = v_37 ^ v_165;
assign v_1586 = v_38 ^ v_166;
assign v_1587 = v_39 ^ v_167;
assign v_1588 = v_40 ^ v_168;
assign v_1589 = v_41 ^ v_169;
assign v_1590 = v_42 ^ v_170;
assign v_1591 = v_43 ^ v_171;
assign v_1592 = v_44 ^ v_172;
assign v_1593 = v_45 ^ v_173;
assign v_1594 = v_46 ^ v_174;
assign v_1595 = v_47 ^ v_175;
assign v_1596 = v_48 ^ v_176;
assign v_1597 = v_49 ^ v_177;
assign v_1598 = v_50 ^ v_178;
assign v_1599 = v_51 ^ v_179;
assign v_1600 = v_52 ^ v_180;
assign v_1601 = v_53 ^ v_181;
assign v_1602 = v_54 ^ v_182;
assign v_1603 = v_55 ^ v_183;
assign v_1604 = v_56 ^ v_184;
assign v_1605 = v_57 ^ v_185;
assign v_1606 = v_58 ^ v_186;
assign v_1607 = v_59 ^ v_187;
assign v_1608 = v_60 ^ v_188;
assign v_1609 = v_61 ^ v_189;
assign v_1610 = v_62 ^ v_190;
assign v_1611 = v_63 ^ v_191;
assign v_1612 = v_64 ^ v_192;
assign v_1614 = v_780 ^ v_844;
assign v_1615 = v_781 ^ v_845;
assign v_1616 = v_782 ^ v_846;
assign v_1617 = v_783 ^ v_847;
assign v_1618 = v_784 ^ v_848;
assign v_1619 = v_785 ^ v_849;
assign v_1620 = v_786 ^ v_850;
assign v_1621 = v_787 ^ v_851;
assign v_1622 = v_788 ^ v_852;
assign v_1623 = v_789 ^ v_853;
assign v_1624 = v_790 ^ v_854;
assign v_1625 = v_791 ^ v_855;
assign v_1626 = v_792 ^ v_856;
assign v_1627 = v_793 ^ v_857;
assign v_1628 = v_794 ^ v_858;
assign v_1629 = v_795 ^ v_859;
assign v_1630 = v_796 ^ v_860;
assign v_1631 = v_797 ^ v_861;
assign v_1632 = v_798 ^ v_862;
assign v_1633 = v_799 ^ v_863;
assign v_1634 = v_800 ^ v_864;
assign v_1635 = v_801 ^ v_865;
assign v_1636 = v_802 ^ v_866;
assign v_1637 = v_803 ^ v_867;
assign v_1638 = v_804 ^ v_868;
assign v_1639 = v_805 ^ v_869;
assign v_1640 = v_806 ^ v_870;
assign v_1641 = v_807 ^ v_871;
assign v_1642 = v_808 ^ v_872;
assign v_1643 = v_809 ^ v_873;
assign v_1644 = v_810 ^ v_874;
assign v_1645 = v_811 ^ v_875;
assign v_1646 = v_812 ^ v_876;
assign v_1647 = v_813 ^ v_877;
assign v_1648 = v_814 ^ v_878;
assign v_1649 = v_815 ^ v_879;
assign v_1650 = v_816 ^ v_880;
assign v_1651 = v_817 ^ v_881;
assign v_1652 = v_818 ^ v_882;
assign v_1653 = v_819 ^ v_883;
assign v_1654 = v_820 ^ v_884;
assign v_1655 = v_821 ^ v_885;
assign v_1656 = v_822 ^ v_886;
assign v_1657 = v_823 ^ v_887;
assign v_1658 = v_824 ^ v_888;
assign v_1659 = v_825 ^ v_889;
assign v_1660 = v_826 ^ v_890;
assign v_1661 = v_827 ^ v_891;
assign v_1662 = v_828 ^ v_892;
assign v_1663 = v_829 ^ v_893;
assign v_1664 = v_830 ^ v_894;
assign v_1665 = v_831 ^ v_895;
assign v_1666 = v_832 ^ v_896;
assign v_1667 = v_833 ^ v_897;
assign v_1668 = v_834 ^ v_898;
assign v_1669 = v_835 ^ v_899;
assign v_1670 = v_836 ^ v_900;
assign v_1671 = v_837 ^ v_901;
assign v_1672 = v_838 ^ v_902;
assign v_1673 = v_839 ^ v_903;
assign v_1674 = v_840 ^ v_904;
assign v_1675 = v_841 ^ v_905;
assign v_1676 = v_842 ^ v_906;
assign v_1677 = v_843 ^ v_907;
assign v_1679 = v_65 ^ v_193;
assign v_1680 = v_66 ^ v_194;
assign v_1681 = v_67 ^ v_195;
assign v_1682 = v_68 ^ v_196;
assign v_1683 = v_69 ^ v_197;
assign v_1684 = v_70 ^ v_198;
assign v_1685 = v_71 ^ v_199;
assign v_1686 = v_72 ^ v_200;
assign v_1687 = v_73 ^ v_201;
assign v_1688 = v_74 ^ v_202;
assign v_1689 = v_75 ^ v_203;
assign v_1690 = v_76 ^ v_204;
assign v_1691 = v_77 ^ v_205;
assign v_1692 = v_78 ^ v_206;
assign v_1693 = v_79 ^ v_207;
assign v_1694 = v_80 ^ v_208;
assign v_1695 = v_81 ^ v_209;
assign v_1696 = v_82 ^ v_210;
assign v_1697 = v_83 ^ v_211;
assign v_1698 = v_84 ^ v_212;
assign v_1699 = v_85 ^ v_213;
assign v_1700 = v_86 ^ v_214;
assign v_1701 = v_87 ^ v_215;
assign v_1702 = v_88 ^ v_216;
assign v_1703 = v_89 ^ v_217;
assign v_1704 = v_90 ^ v_218;
assign v_1705 = v_91 ^ v_219;
assign v_1706 = v_92 ^ v_220;
assign v_1707 = v_93 ^ v_221;
assign v_1708 = v_94 ^ v_222;
assign v_1709 = v_95 ^ v_223;
assign v_1710 = v_96 ^ v_224;
assign v_1711 = v_97 ^ v_225;
assign v_1712 = v_98 ^ v_226;
assign v_1713 = v_99 ^ v_227;
assign v_1714 = v_100 ^ v_228;
assign v_1715 = v_101 ^ v_229;
assign v_1716 = v_102 ^ v_230;
assign v_1717 = v_103 ^ v_231;
assign v_1718 = v_104 ^ v_232;
assign v_1719 = v_105 ^ v_233;
assign v_1720 = v_106 ^ v_234;
assign v_1721 = v_107 ^ v_235;
assign v_1722 = v_108 ^ v_236;
assign v_1723 = v_109 ^ v_237;
assign v_1724 = v_110 ^ v_238;
assign v_1725 = v_111 ^ v_239;
assign v_1726 = v_112 ^ v_240;
assign v_1727 = v_113 ^ v_241;
assign v_1728 = v_114 ^ v_242;
assign v_1729 = v_115 ^ v_243;
assign v_1730 = v_116 ^ v_244;
assign v_1731 = v_117 ^ v_245;
assign v_1732 = v_118 ^ v_246;
assign v_1733 = v_119 ^ v_247;
assign v_1734 = v_120 ^ v_248;
assign v_1735 = v_121 ^ v_249;
assign v_1736 = v_122 ^ v_250;
assign v_1737 = v_123 ^ v_251;
assign v_1738 = v_124 ^ v_252;
assign v_1739 = v_125 ^ v_253;
assign v_1740 = v_126 ^ v_254;
assign v_1741 = v_127 ^ v_255;
assign v_1742 = v_128 ^ v_256;
assign v_1744 = v_1164 ^ v_1228;
assign v_1745 = v_1165 ^ v_1229;
assign v_1746 = v_1166 ^ v_1230;
assign v_1747 = v_1167 ^ v_1231;
assign v_1748 = v_1168 ^ v_1232;
assign v_1749 = v_1169 ^ v_1233;
assign v_1750 = v_1170 ^ v_1234;
assign v_1751 = v_1171 ^ v_1235;
assign v_1752 = v_1172 ^ v_1236;
assign v_1753 = v_1173 ^ v_1237;
assign v_1754 = v_1174 ^ v_1238;
assign v_1755 = v_1175 ^ v_1239;
assign v_1756 = v_1176 ^ v_1240;
assign v_1757 = v_1177 ^ v_1241;
assign v_1758 = v_1178 ^ v_1242;
assign v_1759 = v_1179 ^ v_1243;
assign v_1760 = v_1180 ^ v_1244;
assign v_1761 = v_1181 ^ v_1245;
assign v_1762 = v_1182 ^ v_1246;
assign v_1763 = v_1183 ^ v_1247;
assign v_1764 = v_1184 ^ v_1248;
assign v_1765 = v_1185 ^ v_1249;
assign v_1766 = v_1186 ^ v_1250;
assign v_1767 = v_1187 ^ v_1251;
assign v_1768 = v_1188 ^ v_1252;
assign v_1769 = v_1189 ^ v_1253;
assign v_1770 = v_1190 ^ v_1254;
assign v_1771 = v_1191 ^ v_1255;
assign v_1772 = v_1192 ^ v_1256;
assign v_1773 = v_1193 ^ v_1257;
assign v_1774 = v_1194 ^ v_1258;
assign v_1775 = v_1195 ^ v_1259;
assign v_1776 = v_1196 ^ v_1260;
assign v_1777 = v_1197 ^ v_1261;
assign v_1778 = v_1198 ^ v_1262;
assign v_1779 = v_1199 ^ v_1263;
assign v_1780 = v_1200 ^ v_1264;
assign v_1781 = v_1201 ^ v_1265;
assign v_1782 = v_1202 ^ v_1266;
assign v_1783 = v_1203 ^ v_1267;
assign v_1784 = v_1204 ^ v_1268;
assign v_1785 = v_1205 ^ v_1269;
assign v_1786 = v_1206 ^ v_1270;
assign v_1787 = v_1207 ^ v_1271;
assign v_1788 = v_1208 ^ v_1272;
assign v_1789 = v_1209 ^ v_1273;
assign v_1790 = v_1210 ^ v_1274;
assign v_1791 = v_1211 ^ v_1275;
assign v_1792 = v_1212 ^ v_1276;
assign v_1793 = v_1213 ^ v_1277;
assign v_1794 = v_1214 ^ v_1278;
assign v_1795 = v_1215 ^ v_1279;
assign v_1796 = v_1216 ^ v_1280;
assign v_1797 = v_1217 ^ v_1281;
assign v_1798 = v_1218 ^ v_1282;
assign v_1799 = v_1219 ^ v_1283;
assign v_1800 = v_1220 ^ v_1284;
assign v_1801 = v_1221 ^ v_1285;
assign v_1802 = v_1222 ^ v_1286;
assign v_1803 = v_1223 ^ v_1287;
assign v_1804 = v_1224 ^ v_1288;
assign v_1805 = v_1225 ^ v_1289;
assign v_1806 = v_1226 ^ v_1290;
assign v_1807 = v_1227 ^ v_1291;
assign x_1 = ~v_449 | ~v_448;
assign x_2 = ~v_517 | v_516;
assign x_3 = ~v_1162 | v_1161;
assign x_4 = ~v_1546 | v_1545;
assign x_5 = v_1548 | ~v_779;
assign x_6 = v_1678 | ~v_1613;
assign x_7 = v_1808 | ~v_1743;
assign x_8 = x_2 & x_3;
assign x_9 = x_1 & x_8;
assign x_10 = x_4 & x_5;
assign x_11 = x_6 & x_7;
assign x_12 = x_10 & x_11;
assign x_13 = x_9 & x_12;
assign o_1 = x_13;
endmodule
