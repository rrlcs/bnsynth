// skolem function for order file variables
// Generated using findDep.cpp 
module sortnetsort7.AE.stepl.005 (v_49, v_50, v_51, v_52, v_53, v_54, v_55, v_56, v_57, v_58, v_59, v_60, v_61, v_62, v_63, v_64, v_65, v_66, v_67, v_68, v_69, v_70, v_71, v_72, v_73, v_74, v_75, v_76, v_77, v_78, v_79, v_80, v_81, v_82, v_83, v_84, v_85, v_86, v_87, v_88, v_89, v_90, v_91, v_92, v_93, v_94, v_95, v_96, v_97, v_98, v_99, v_100, v_101, v_102, v_103, v_104, v_105, v_106, v_107, v_108, v_109, v_110, v_111, v_112, v_113, v_114, v_115, v_116, v_117, v_118, v_119, v_120, v_121, v_122, v_123, v_124, v_125, v_126, v_127, v_128, v_129, v_130, v_131, v_132, v_133, v_134, v_135, v_136, v_137, v_138, v_139, v_140, v_141, v_142, v_143, v_144, v_145, v_146, v_147, v_148, v_149, v_150, v_151, v_152, v_153, v_154, v_155, v_156, v_157, v_158, v_159, v_160, v_161, v_162, v_163, v_164, v_165, v_166, v_167, v_168, v_169, v_170, v_171, v_172, v_173, v_174, v_175, v_176, v_177, v_178, v_179, v_180, v_181, v_182, v_183, v_184, v_185, v_186, v_187, v_188, v_189, v_190, v_191, v_192, v_193, v_194, v_195, v_196, v_197, v_198, v_199, v_200, v_201, v_202, v_203, v_204, v_205, v_206, v_207, v_208, v_209, v_210, v_211, v_212, v_213, v_1843, v_1844, v_1845, v_1846, v_1847, v_1848, v_1849, v_1850, v_1851, v_1852, v_1853, v_1854, v_1855, v_1856, v_1857, v_1858, v_1859, v_1860, v_1861, v_1862, v_1863, v_1864, v_1865, v_1866, v_1867, v_1868, v_1869, v_1870, v_1871, v_1872, v_1873, v_1874, v_1875, v_1876, v_1877, v_1878, v_1879, v_1880, v_1881, v_1882, v_1883, v_1884, v_1885, v_1886, v_1887, v_1888, v_1889, v_1890, v_1891, v_1892, v_1893, v_1894, v_1895, v_1896, v_1897, v_1898, v_1899, v_1900, v_1901, v_1902, v_1945, v_1946, v_1947, v_1948, v_1949, v_1950, v_1951, v_1952, v_1953, v_1954, v_1955, v_1956, v_1957, v_1958, v_1959, v_1960, v_1961, v_1962, v_1963, v_1964, v_1965, v_1966, v_1967, v_1968, v_1969, v_1970, v_1971, v_1972, v_1973, v_1974, v_1975, v_1976, v_1977, v_1978, v_1979, v_1980, v_1981, v_1982, v_1983, v_1984, v_1985, v_1986, v_1987, v_1988, v_1989, v_1990, v_1991, v_1992, v_1993, v_1994, v_1995, v_1996, v_1997, v_1998, v_1999, v_2000, v_2001, v_2002, v_2003, v_2004, v_2047, v_2048, v_2049, v_2050, v_2051, v_2052, v_2053, v_2054, v_2055, v_2056, v_2057, v_2058, v_2059, v_2060, v_2061, v_2062, v_2063, v_2064, v_2065, v_2066, v_2067, v_2068, v_2069, v_2070, v_2071, v_2072, v_2073, v_2074, v_2075, v_2076, v_2077, v_2078, v_2079, v_2080, v_2081, v_2082, v_2083, v_2084, v_2085, v_2086, v_2087, v_2088, v_2089, v_2090, v_2091, v_2092, v_2093, v_2094, v_2095, v_2096, v_2097, v_2098, v_2099, v_2100, v_2101, v_2102, v_2103, v_2104, v_2105, v_2106, v_2149, v_2150, v_2151, v_2152, v_2153, v_2154, v_2155, v_2156, v_2157, v_2158, v_2159, v_2160, v_2161, v_2162, v_2163, v_2164, v_2165, v_2166, v_2167, v_2168, v_2169, v_2170, v_2171, v_2172, v_2173, v_2174, v_2175, v_2176, v_2177, v_2178, v_2179, v_2180, v_2181, v_2182, v_2183, v_2184, v_2185, v_2186, v_2187, v_2188, v_2189, v_2190, v_2191, v_2192, v_2193, v_2194, v_2195, v_2196, v_2197, v_2198, v_2199, v_2200, v_2201, v_2202, v_2203, v_2204, v_2205, v_2206, v_2207, v_2208, v_1, v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_12, v_13, v_14, v_15, v_16, v_17, v_18, v_19, v_20, v_21, v_22, v_23, v_24, v_25, v_26, v_27, v_28, v_29, v_30, v_31, v_32, v_33, v_34, v_35, v_36, v_37, v_38, v_39, v_40, v_41, v_42, v_43, v_44, v_45, v_46, v_47, v_48, v_214, v_215, v_216, v_217, v_218, v_219, v_220, v_221, v_222, v_223, v_224, v_225, v_226, v_227, v_228, v_229, v_230, v_231, v_232, v_233, v_234, v_235, v_236, v_237, v_238, v_239, v_240, v_241, v_242, v_243, v_244, v_245, v_246, v_247, v_248, v_249, v_250, v_251, v_252, v_253, v_254, v_255, v_256, v_257, v_258, v_259, v_260, v_261, v_262, v_263, v_264, v_265, v_266, v_267, v_268, v_269, v_270, v_271, v_272, v_273, v_274, v_275, v_276, v_277, v_278, v_279, v_280, v_281, v_282, v_283, v_284, v_285, v_286, v_287, v_288, v_289, v_290, v_291, v_292, v_293, v_294, v_295, v_296, v_297, v_298, v_299, v_300, v_301, v_302, v_303, v_304, v_305, v_306, v_307, v_308, v_309, v_310, v_311, v_312, v_313, v_314, v_315, v_316, v_317, v_318, v_319, v_320, v_321, v_322, v_323, v_324, v_325, v_326, v_327, v_328, v_329, v_330, v_331, v_332, v_333, v_334, v_335, v_336, v_337, v_338, v_339, v_340, v_341, v_342, v_343, v_344, v_345, v_346, v_368, v_369, v_370, v_371, v_372, v_373, v_374, v_375, v_376, v_377, v_378, v_379, v_380, v_381, v_382, v_383, v_384, v_385, v_386, v_387, v_388, v_389, v_390, v_391, v_392, v_393, v_394, v_395, v_396, v_397, v_398, v_399, v_400, v_401, v_402, v_403, v_404, v_405, v_406, v_407, v_408, v_409, v_410, v_411, v_412, v_413, v_414, v_415, v_416, v_417, v_418, v_419, v_420, v_421, v_422, v_423, v_424, v_425, v_426, v_427, v_428, v_429, v_430, v_431, v_432, v_433, v_434, v_435, v_436, v_437, v_438, v_439, v_440, v_441, v_442, v_443, v_444, v_445, v_446, v_447, v_448, v_449, v_450, v_451, v_452, v_474, v_475, v_476, v_477, v_478, v_479, v_480, v_481, v_482, v_483, v_484, v_485, v_486, v_487, v_488, v_489, v_490, v_491, v_492, v_493, v_494, v_495, v_496, v_497, v_498, v_499, v_500, v_501, v_502, v_503, v_504, v_505, v_506, v_507, v_508, v_509, v_510, v_511, v_512, v_513, v_514, v_515, v_516, v_517, v_518, v_519, v_520, v_521, v_522, v_523, v_524, v_525, v_526, v_527, v_528, v_529, v_530, v_531, v_532, v_533, v_534, v_535, v_536, v_537, v_538, v_539, v_540, v_541, v_542, v_543, v_544, v_545, v_546, v_547, v_548, v_549, v_550, v_551, v_552, v_553, v_554, v_555, v_556, v_557, v_558, v_580, v_581, v_582, v_583, v_584, v_585, v_586, v_587, v_588, v_589, v_590, v_591, v_592, v_593, v_594, v_595, v_596, v_597, v_598, v_599, v_600, v_601, v_602, v_603, v_604, v_605, v_606, v_607, v_608, v_609, v_610, v_611, v_612, v_613, v_614, v_615, v_616, v_617, v_618, v_619, v_620, v_621, v_622, v_623, v_624, v_625, v_626, v_627, v_628, v_629, v_630, v_631, v_632, v_633, v_634, v_635, v_636, v_637, v_638, v_639, v_640, v_641, v_642, v_643, v_644, v_645, v_646, v_647, v_648, v_649, v_650, v_651, v_652, v_653, v_654, v_655, v_656, v_657, v_658, v_659, v_660, v_661, v_662, v_663, v_664, v_686, v_687, v_688, v_689, v_690, v_691, v_692, v_693, v_694, v_695, v_696, v_697, v_698, v_699, v_700, v_701, v_702, v_703, v_704, v_705, v_706, v_707, v_708, v_709, v_710, v_711, v_712, v_713, v_714, v_715, v_716, v_717, v_718, v_719, v_720, v_721, v_722, v_723, v_724, v_725, v_726, v_727, v_728, v_729, v_730, v_731, v_732, v_733, v_734, v_735, v_736, v_737, v_738, v_739, v_740, v_741, v_742, v_743, v_744, v_745, v_746, v_747, v_748, v_749, v_750, v_751, v_752, v_753, v_754, v_755, v_756, v_757, v_758, v_759, v_760, v_761, v_762, v_763, v_764, v_765, v_766, v_767, v_768, v_769, v_770, v_792, v_793, v_794, v_795, v_796, v_797, v_798, v_799, v_800, v_801, v_802, v_803, v_804, v_805, v_806, v_807, v_808, v_809, v_810, v_811, v_812, v_813, v_814, v_815, v_816, v_817, v_818, v_819, v_820, v_821, v_822, v_823, v_824, v_825, v_826, v_827, v_828, v_829, v_830, v_831, v_832, v_833, v_834, v_835, v_836, v_837, v_838, v_839, v_840, v_841, v_842, v_843, v_844, v_845, v_846, v_847, v_848, v_849, v_850, v_851, v_852, v_853, v_854, v_855, v_856, v_857, v_858, v_859, v_860, v_861, v_862, v_863, v_864, v_865, v_866, v_867, v_868, v_869, v_870, v_871, v_872, v_873, v_874, v_875, v_876, v_877, v_878, v_879, v_880, v_881, v_882, v_883, v_884, v_885, v_886, v_887, v_888, v_889, v_890, v_891, v_892, v_893, v_894, v_895, v_896, v_897, v_898, v_899, v_900, v_901, v_902, v_903, v_904, v_905, v_906, v_907, v_908, v_909, v_910, v_911, v_912, v_913, v_914, v_915, v_916, v_917, v_918, v_919, v_920, v_921, v_922, v_923, v_924, v_925, v_926, v_927, v_928, v_929, v_930, v_931, v_932, v_933, v_934, v_935, v_936, v_937, v_938, v_939, v_940, v_941, v_942, v_943, v_944, v_945, v_946, v_947, v_948, v_949, v_950, v_951, v_952, v_953, v_954, v_955, v_956, v_957, v_958, v_959, v_960, v_961, v_962, v_963, v_964, v_965, v_966, v_967, v_968, v_969, v_970, v_971, v_972, v_973, v_974, v_975, v_976, v_977, v_978, v_979, v_980, v_981, v_982, v_983, v_984, v_985, v_986, v_987, v_988, v_989, v_990, v_991, v_992, v_993, v_994, v_995, v_996, v_997, v_998, v_999, v_1000, v_1001, v_1002, v_1003, v_1004, v_1005, v_1006, v_1007, v_1008, v_1009, v_1010, v_1011, v_1012, v_1013, v_1014, v_1015, v_1016, v_1017, v_1018, v_1019, v_1020, v_1021, v_1022, v_1023, v_1024, v_1025, v_1026, v_1027, v_1028, v_1029, v_1030, v_1031, v_1032, v_1033, v_1034, v_1035, v_1036, v_1037, v_1038, v_1039, v_1040, v_1041, v_1042, v_1043, v_1044, v_1045, v_1046, v_1047, v_1048, v_1049, v_1050, v_1051, v_1052, v_1053, v_1054, v_1055, v_1056, v_1057, v_1058, v_1059, v_1060, v_1061, v_1062, v_1063, v_1064, v_1065, v_1066, v_1067, v_1068, v_1069, v_1070, v_1071, v_1072, v_1073, v_1074, v_1075, v_1076, v_1077, v_1078, v_1079, v_1080, v_1081, v_1082, v_1083, v_1084, v_1085, v_1086, v_1087, v_1088, v_1089, v_1090, v_1091, v_1092, v_1093, v_1094, v_1095, v_1096, v_1097, v_1098, v_1099, v_1100, v_1101, v_1102, v_1103, v_1104, v_1105, v_1106, v_1107, v_1108, v_1109, v_1110, v_1111, v_1112, v_1113, v_1114, v_1115, v_1116, v_1117, v_1118, v_1119, v_1120, v_1121, v_1122, v_1123, v_1124, v_1125, v_1126, v_1127, v_1128, v_1129, v_1130, v_1131, v_1132, v_1133, v_1134, v_1135, v_1136, v_1137, v_1138, v_1139, v_1140, v_1141, v_1142, v_1143, v_1144, v_1145, v_1146, v_1147, v_1148, v_1149, v_1150, v_1151, v_1152, v_1153, v_1154, v_1155, v_1156, v_1157, v_1158, v_1159, v_1160, v_1161, v_1162, v_1163, v_1164, v_1165, v_1166, v_1167, v_1168, v_1169, v_1170, v_1171, v_1172, v_1173, v_1174, v_1175, v_1176, v_1177, v_1178, v_1179, v_1180, v_1181, v_1182, v_1183, v_1184, v_1185, v_1186, v_1187, v_1188, v_1189, v_1190, v_1191, v_1192, v_1193, v_1194, v_1195, v_1196, v_1197, v_1198, v_1199, v_1200, v_1201, v_1202, v_1203, v_1204, v_1205, v_1206, v_1207, v_1208, v_1209, v_1210, v_1211, v_1212, v_1213, v_1214, v_1215, v_1216, v_1217, v_1218, v_1219, v_1220, v_1221, v_1222, v_1223, v_1224, v_1225, v_1226, v_1227, v_1228, v_1229, v_1230, v_1231, v_1232, v_1233, v_1234, v_1235, v_1236, v_1237, v_1238, v_1239, v_1240, v_1241, v_1242, v_1243, v_1244, v_1245, v_1246, v_1247, v_1248, v_1249, v_1250, v_1251, v_1252, v_1253, v_1254, v_1255, v_1256, v_1257, v_1258, v_1259, v_1260, v_1261, v_1262, v_1263, v_1264, v_1265, v_1266, v_1267, v_1268, v_1269, v_1270, v_1271, v_1272, v_1273, v_1274, v_1275, v_1276, v_1277, v_1278, v_1279, v_1280, v_1281, v_1282, v_1283, v_1284, v_1285, v_1286, v_1287, v_1288, v_1289, v_1290, v_1291, v_1292, v_1293, v_1294, v_1295, v_1296, v_1297, v_1298, v_1299, v_1300, v_1301, v_1302, v_1303, v_1304, v_1305, v_1306, v_1307, v_1308, v_1309, v_1310, v_1311, v_1312, v_1313, v_1314, v_1315, v_1316, v_1317, v_1318, v_1319, v_1320, v_1321, v_1322, v_1323, v_1324, v_1325, v_1326, v_1327, v_1328, v_1329, v_1330, v_1331, v_1332, v_1333, v_1334, v_1335, v_1336, v_1337, v_1338, v_1339, v_1340, v_1341, v_1342, v_1343, v_1344, v_1345, v_1346, v_1347, v_1348, v_1349, v_1350, v_1351, v_1352, v_1353, v_1354, v_1355, v_1356, v_1357, v_1358, v_1359, v_1360, v_1361, v_1362, v_1363, v_1364, v_1365, v_1366, v_1367, v_1368, v_1369, v_1370, v_1371, v_1372, v_1373, v_1374, v_1375, v_1376, v_1377, v_1378, v_1379, v_1380, v_1381, v_1382, v_1383, v_1384, v_1385, v_1386, v_1387, v_1388, v_1389, v_1390, v_1391, v_1392, v_1393, v_1394, v_1395, v_1396, v_1397, v_1398, v_1399, v_1400, v_1401, v_1402, v_1403, v_1404, v_1405, v_1406, v_1407, v_1408, v_1409, v_1410, v_1411, v_1412, v_1413, v_1414, v_1415, v_1416, v_1417, v_1418, v_1419, v_1420, v_1421, v_1422, v_1423, v_1424, v_1425, v_1426, v_1427, v_1428, v_1429, v_1430, v_1431, v_1432, v_1433, v_1434, v_1435, v_1436, v_1437, v_1438, v_1439, v_1440, v_1441, v_1442, v_1443, v_1444, v_1445, v_1446, v_1447, v_1448, v_1449, v_1450, v_1451, v_1452, v_1453, v_1454, v_1455, v_1456, v_1457, v_1458, v_1459, v_1460, v_1461, v_1462, v_1463, v_1464, v_1465, v_1466, v_1467, v_1468, v_1469, v_1470, v_1471, v_1472, v_1473, v_1474, v_1475, v_1476, v_1477, v_1478, v_1479, v_1480, v_1481, v_1482, v_1483, v_1484, v_1485, v_1486, v_1487, v_1488, v_1489, v_1490, v_1491, v_1492, v_1493, v_1494, v_1495, v_1496, v_1497, v_1498, v_1499, v_1500, v_1501, v_1502, v_1503, v_1504, v_1505, v_1506, v_1507, v_1508, v_1509, v_1510, v_1511, v_1512, v_1513, v_1514, v_1515, v_1516, v_1517, v_1518, v_1519, v_1520, v_1521, v_1522, v_1523, v_1524, v_1525, v_1526, v_1527, v_1528, v_1529, v_1530, v_1531, v_1532, v_1533, v_1534, v_1535, v_1536, v_1537, v_1538, v_1539, v_1540, v_1541, v_1542, v_1543, v_1544, v_1545, v_1546, v_1547, v_1548, v_1549, v_1550, v_1551, v_1552, v_1553, v_1554, v_1555, v_1556, v_1557, v_1558, v_1559, v_1560, v_1561, v_1562, v_1563, v_1564, v_1565, v_1566, v_1567, v_1568, v_1569, v_1570, v_1571, v_1572, v_1573, v_1574, v_1575, v_1576, v_1577, v_1578, v_1579, v_1580, v_1581, v_1582, v_1583, v_1584, v_1585, v_1586, v_1587, v_1588, v_1589, v_1590, v_1591, v_1592, v_1593, v_1594, v_1595, v_1596, v_1597, v_1598, v_1599, v_1600, v_1601, v_1602, v_1603, v_1604, v_1605, v_1606, v_1607, v_1608, v_1609, v_1610, v_1611, v_1612, v_1613, v_1614, v_1615, v_1616, v_1617, v_1618, v_1619, v_1620, v_1621, v_1622, v_1623, v_1624, v_1625, v_1626, v_1627, v_1628, v_1629, v_1630, v_1631, v_1632, v_1633, v_1634, v_1635, v_1636, v_1637, v_1638, v_1639, v_1640, v_1641, v_1642, v_1643, v_1644, v_1645, v_1646, v_1647, v_1648, v_1649, v_1650, v_1651, v_1652, v_1653, v_1654, v_1655, v_1656, v_1657, v_1658, v_1659, v_1660, v_1661, v_1662, v_1663, v_1664, v_1665, v_1666, v_1667, v_1668, v_1669, v_1670, v_1671, v_1672, v_1673, v_1674, v_1675, v_1676, v_1677, v_1678, v_1679, v_1680, v_1681, v_1682, v_1683, v_1684, v_1685, v_1686, v_1687, v_1688, v_1689, v_1690, v_1691, v_1692, v_1693, v_1694, v_1695, v_1696, v_1697, v_1698, v_1699, v_1700, v_1701, v_1702, v_1703, v_1704, v_1705, v_1706, v_1707, v_1708, v_1709, v_1710, v_1711, v_1712, v_1713, v_1714, v_1715, v_1716, v_1717, v_1718, v_1719, v_1720, v_1721, v_1722, v_1723, v_1724, v_1725, v_1726, v_1727, v_1728, v_1729, v_1730, v_1731, v_1732, v_1733, v_1734, v_1735, v_1736, v_1737, v_1738, v_1739, v_1740, v_1741, v_1742, v_1743, v_1744, v_1745, v_1746, v_1747, v_1748, v_1749, v_1750, v_1751, v_1752, v_1753, v_1754, v_1755, v_1756, v_1757, v_1758, v_1759, v_1760, v_1761, v_1762, v_1763, v_1764, v_1765, v_1766, v_1767, v_1768, v_1769, v_1770, v_1771, v_1772, v_1773, v_1774, v_1775, v_1776, v_1777, v_1778, v_1779, v_1780, v_1781, v_1782, v_1783, v_1784, v_1785, v_1786, v_1787, v_1788, v_1789, v_1790, v_1791, v_1792, v_1793, v_1794, v_1795, v_1796, v_1797, v_1798, v_1799, v_1800, v_1801, v_1802, v_1803, v_1804, v_1805, v_1806, v_1807, v_1808, v_1809, v_1810, v_1811, v_1812, v_1813, v_1814, v_1815, v_1816, v_1817, v_1818, v_1819, v_1820, v_1821, v_1822, v_1823, v_1824, v_1825, v_1826, v_1827, v_1828, v_1829, v_1830, v_1831, v_1832, v_1833, v_1834, v_1835, v_1836, v_1837, v_1838, v_1839, v_1840, v_1841, v_1842, v_1903, v_1904, v_1905, v_1906, v_1907, v_1908, v_1909, v_1910, v_1911, v_1912, v_1913, v_1914, v_1915, v_1916, v_1917, v_1918, v_1919, v_1920, v_1921, v_1922, v_1923, v_1924, v_1925, v_1926, v_1927, v_1928, v_1929, v_1930, v_1931, v_1932, v_1933, v_1934, v_1935, v_1936, v_1937, v_1938, v_1939, v_1940, v_1941, v_1942, v_1943, v_1944, v_2005, v_2006, v_2007, v_2008, v_2009, v_2010, v_2011, v_2012, v_2013, v_2014, v_2015, v_2016, v_2017, v_2018, v_2019, v_2020, v_2021, v_2022, v_2023, v_2024, v_2025, v_2026, v_2027, v_2028, v_2029, v_2030, v_2031, v_2032, v_2033, v_2034, v_2035, v_2036, v_2037, v_2038, v_2039, v_2040, v_2041, v_2042, v_2043, v_2044, v_2045, v_2046, v_2107, v_2108, v_2109, v_2110, v_2111, v_2112, v_2113, v_2114, v_2115, v_2116, v_2117, v_2118, v_2119, v_2120, v_2121, v_2122, v_2123, v_2124, v_2125, v_2126, v_2127, v_2128, v_2129, v_2130, v_2131, v_2132, v_2133, v_2134, v_2135, v_2136, v_2137, v_2138, v_2139, v_2140, v_2141, v_2142, v_2143, v_2144, v_2145, v_2146, v_2147, v_2148, v_2209, v_2210, v_2211, v_2212, v_2213, v_2214, v_2215, v_2216, v_2217, v_2218, v_2219, v_2220, v_2221, v_2222, v_2223, v_2224, v_2225, v_2226, v_2227, v_2228, v_2229, v_2230, v_2231, v_2232, v_2233, v_2234, v_2235, v_2236, v_2237, v_2238, v_2239, v_2240, v_2241, v_2242, v_2243, v_2244, v_2245, v_2246, v_2247, v_2248, v_2249, v_2250, o_1);
input v_49;
input v_50;
input v_51;
input v_52;
input v_53;
input v_54;
input v_55;
input v_56;
input v_57;
input v_58;
input v_59;
input v_60;
input v_61;
input v_62;
input v_63;
input v_64;
input v_65;
input v_66;
input v_67;
input v_68;
input v_69;
input v_70;
input v_71;
input v_72;
input v_73;
input v_74;
input v_75;
input v_76;
input v_77;
input v_78;
input v_79;
input v_80;
input v_81;
input v_82;
input v_83;
input v_84;
input v_85;
input v_86;
input v_87;
input v_88;
input v_89;
input v_90;
input v_91;
input v_92;
input v_93;
input v_94;
input v_95;
input v_96;
input v_97;
input v_98;
input v_99;
input v_100;
input v_101;
input v_102;
input v_103;
input v_104;
input v_105;
input v_106;
input v_107;
input v_108;
input v_109;
input v_110;
input v_111;
input v_112;
input v_113;
input v_114;
input v_115;
input v_116;
input v_117;
input v_118;
input v_119;
input v_120;
input v_121;
input v_122;
input v_123;
input v_124;
input v_125;
input v_126;
input v_127;
input v_128;
input v_129;
input v_130;
input v_131;
input v_132;
input v_133;
input v_134;
input v_135;
input v_136;
input v_137;
input v_138;
input v_139;
input v_140;
input v_141;
input v_142;
input v_143;
input v_144;
input v_145;
input v_146;
input v_147;
input v_148;
input v_149;
input v_150;
input v_151;
input v_152;
input v_153;
input v_154;
input v_155;
input v_156;
input v_157;
input v_158;
input v_159;
input v_160;
input v_161;
input v_162;
input v_163;
input v_164;
input v_165;
input v_166;
input v_167;
input v_168;
input v_169;
input v_170;
input v_171;
input v_172;
input v_173;
input v_174;
input v_175;
input v_176;
input v_177;
input v_178;
input v_179;
input v_180;
input v_181;
input v_182;
input v_183;
input v_184;
input v_185;
input v_186;
input v_187;
input v_188;
input v_189;
input v_190;
input v_191;
input v_192;
input v_193;
input v_194;
input v_195;
input v_196;
input v_197;
input v_198;
input v_199;
input v_200;
input v_201;
input v_202;
input v_203;
input v_204;
input v_205;
input v_206;
input v_207;
input v_208;
input v_209;
input v_210;
input v_211;
input v_212;
input v_213;
input v_1843;
input v_1844;
input v_1845;
input v_1846;
input v_1847;
input v_1848;
input v_1849;
input v_1850;
input v_1851;
input v_1852;
input v_1853;
input v_1854;
input v_1855;
input v_1856;
input v_1857;
input v_1858;
input v_1859;
input v_1860;
input v_1861;
input v_1862;
input v_1863;
input v_1864;
input v_1865;
input v_1866;
input v_1867;
input v_1868;
input v_1869;
input v_1870;
input v_1871;
input v_1872;
input v_1873;
input v_1874;
input v_1875;
input v_1876;
input v_1877;
input v_1878;
input v_1879;
input v_1880;
input v_1881;
input v_1882;
input v_1883;
input v_1884;
input v_1885;
input v_1886;
input v_1887;
input v_1888;
input v_1889;
input v_1890;
input v_1891;
input v_1892;
input v_1893;
input v_1894;
input v_1895;
input v_1896;
input v_1897;
input v_1898;
input v_1899;
input v_1900;
input v_1901;
input v_1902;
input v_1945;
input v_1946;
input v_1947;
input v_1948;
input v_1949;
input v_1950;
input v_1951;
input v_1952;
input v_1953;
input v_1954;
input v_1955;
input v_1956;
input v_1957;
input v_1958;
input v_1959;
input v_1960;
input v_1961;
input v_1962;
input v_1963;
input v_1964;
input v_1965;
input v_1966;
input v_1967;
input v_1968;
input v_1969;
input v_1970;
input v_1971;
input v_1972;
input v_1973;
input v_1974;
input v_1975;
input v_1976;
input v_1977;
input v_1978;
input v_1979;
input v_1980;
input v_1981;
input v_1982;
input v_1983;
input v_1984;
input v_1985;
input v_1986;
input v_1987;
input v_1988;
input v_1989;
input v_1990;
input v_1991;
input v_1992;
input v_1993;
input v_1994;
input v_1995;
input v_1996;
input v_1997;
input v_1998;
input v_1999;
input v_2000;
input v_2001;
input v_2002;
input v_2003;
input v_2004;
input v_2047;
input v_2048;
input v_2049;
input v_2050;
input v_2051;
input v_2052;
input v_2053;
input v_2054;
input v_2055;
input v_2056;
input v_2057;
input v_2058;
input v_2059;
input v_2060;
input v_2061;
input v_2062;
input v_2063;
input v_2064;
input v_2065;
input v_2066;
input v_2067;
input v_2068;
input v_2069;
input v_2070;
input v_2071;
input v_2072;
input v_2073;
input v_2074;
input v_2075;
input v_2076;
input v_2077;
input v_2078;
input v_2079;
input v_2080;
input v_2081;
input v_2082;
input v_2083;
input v_2084;
input v_2085;
input v_2086;
input v_2087;
input v_2088;
input v_2089;
input v_2090;
input v_2091;
input v_2092;
input v_2093;
input v_2094;
input v_2095;
input v_2096;
input v_2097;
input v_2098;
input v_2099;
input v_2100;
input v_2101;
input v_2102;
input v_2103;
input v_2104;
input v_2105;
input v_2106;
input v_2149;
input v_2150;
input v_2151;
input v_2152;
input v_2153;
input v_2154;
input v_2155;
input v_2156;
input v_2157;
input v_2158;
input v_2159;
input v_2160;
input v_2161;
input v_2162;
input v_2163;
input v_2164;
input v_2165;
input v_2166;
input v_2167;
input v_2168;
input v_2169;
input v_2170;
input v_2171;
input v_2172;
input v_2173;
input v_2174;
input v_2175;
input v_2176;
input v_2177;
input v_2178;
input v_2179;
input v_2180;
input v_2181;
input v_2182;
input v_2183;
input v_2184;
input v_2185;
input v_2186;
input v_2187;
input v_2188;
input v_2189;
input v_2190;
input v_2191;
input v_2192;
input v_2193;
input v_2194;
input v_2195;
input v_2196;
input v_2197;
input v_2198;
input v_2199;
input v_2200;
input v_2201;
input v_2202;
input v_2203;
input v_2204;
input v_2205;
input v_2206;
input v_2207;
input v_2208;
input v_1;
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_13;
input v_14;
input v_15;
input v_16;
input v_17;
input v_18;
input v_19;
input v_20;
input v_21;
input v_22;
input v_23;
input v_24;
input v_25;
input v_26;
input v_27;
input v_28;
input v_29;
input v_30;
input v_31;
input v_32;
input v_33;
input v_34;
input v_35;
input v_36;
input v_37;
input v_38;
input v_39;
input v_40;
input v_41;
input v_42;
input v_43;
input v_44;
input v_45;
input v_46;
input v_47;
input v_48;
input v_214;
input v_215;
input v_216;
input v_217;
input v_218;
input v_219;
input v_220;
input v_221;
input v_222;
input v_223;
input v_224;
input v_225;
input v_226;
input v_227;
input v_228;
input v_229;
input v_230;
input v_231;
input v_232;
input v_233;
input v_234;
input v_235;
input v_236;
input v_237;
input v_238;
input v_239;
input v_240;
input v_241;
input v_242;
input v_243;
input v_244;
input v_245;
input v_246;
input v_247;
input v_248;
input v_249;
input v_250;
input v_251;
input v_252;
input v_253;
input v_254;
input v_255;
input v_256;
input v_257;
input v_258;
input v_259;
input v_260;
input v_261;
input v_262;
input v_263;
input v_264;
input v_265;
input v_266;
input v_267;
input v_268;
input v_269;
input v_270;
input v_271;
input v_272;
input v_273;
input v_274;
input v_275;
input v_276;
input v_277;
input v_278;
input v_279;
input v_280;
input v_281;
input v_282;
input v_283;
input v_284;
input v_285;
input v_286;
input v_287;
input v_288;
input v_289;
input v_290;
input v_291;
input v_292;
input v_293;
input v_294;
input v_295;
input v_296;
input v_297;
input v_298;
input v_299;
input v_300;
input v_301;
input v_302;
input v_303;
input v_304;
input v_305;
input v_306;
input v_307;
input v_308;
input v_309;
input v_310;
input v_311;
input v_312;
input v_313;
input v_314;
input v_315;
input v_316;
input v_317;
input v_318;
input v_319;
input v_320;
input v_321;
input v_322;
input v_323;
input v_324;
input v_325;
input v_326;
input v_327;
input v_328;
input v_329;
input v_330;
input v_331;
input v_332;
input v_333;
input v_334;
input v_335;
input v_336;
input v_337;
input v_338;
input v_339;
input v_340;
input v_341;
input v_342;
input v_343;
input v_344;
input v_345;
input v_346;
input v_368;
input v_369;
input v_370;
input v_371;
input v_372;
input v_373;
input v_374;
input v_375;
input v_376;
input v_377;
input v_378;
input v_379;
input v_380;
input v_381;
input v_382;
input v_383;
input v_384;
input v_385;
input v_386;
input v_387;
input v_388;
input v_389;
input v_390;
input v_391;
input v_392;
input v_393;
input v_394;
input v_395;
input v_396;
input v_397;
input v_398;
input v_399;
input v_400;
input v_401;
input v_402;
input v_403;
input v_404;
input v_405;
input v_406;
input v_407;
input v_408;
input v_409;
input v_410;
input v_411;
input v_412;
input v_413;
input v_414;
input v_415;
input v_416;
input v_417;
input v_418;
input v_419;
input v_420;
input v_421;
input v_422;
input v_423;
input v_424;
input v_425;
input v_426;
input v_427;
input v_428;
input v_429;
input v_430;
input v_431;
input v_432;
input v_433;
input v_434;
input v_435;
input v_436;
input v_437;
input v_438;
input v_439;
input v_440;
input v_441;
input v_442;
input v_443;
input v_444;
input v_445;
input v_446;
input v_447;
input v_448;
input v_449;
input v_450;
input v_451;
input v_452;
input v_474;
input v_475;
input v_476;
input v_477;
input v_478;
input v_479;
input v_480;
input v_481;
input v_482;
input v_483;
input v_484;
input v_485;
input v_486;
input v_487;
input v_488;
input v_489;
input v_490;
input v_491;
input v_492;
input v_493;
input v_494;
input v_495;
input v_496;
input v_497;
input v_498;
input v_499;
input v_500;
input v_501;
input v_502;
input v_503;
input v_504;
input v_505;
input v_506;
input v_507;
input v_508;
input v_509;
input v_510;
input v_511;
input v_512;
input v_513;
input v_514;
input v_515;
input v_516;
input v_517;
input v_518;
input v_519;
input v_520;
input v_521;
input v_522;
input v_523;
input v_524;
input v_525;
input v_526;
input v_527;
input v_528;
input v_529;
input v_530;
input v_531;
input v_532;
input v_533;
input v_534;
input v_535;
input v_536;
input v_537;
input v_538;
input v_539;
input v_540;
input v_541;
input v_542;
input v_543;
input v_544;
input v_545;
input v_546;
input v_547;
input v_548;
input v_549;
input v_550;
input v_551;
input v_552;
input v_553;
input v_554;
input v_555;
input v_556;
input v_557;
input v_558;
input v_580;
input v_581;
input v_582;
input v_583;
input v_584;
input v_585;
input v_586;
input v_587;
input v_588;
input v_589;
input v_590;
input v_591;
input v_592;
input v_593;
input v_594;
input v_595;
input v_596;
input v_597;
input v_598;
input v_599;
input v_600;
input v_601;
input v_602;
input v_603;
input v_604;
input v_605;
input v_606;
input v_607;
input v_608;
input v_609;
input v_610;
input v_611;
input v_612;
input v_613;
input v_614;
input v_615;
input v_616;
input v_617;
input v_618;
input v_619;
input v_620;
input v_621;
input v_622;
input v_623;
input v_624;
input v_625;
input v_626;
input v_627;
input v_628;
input v_629;
input v_630;
input v_631;
input v_632;
input v_633;
input v_634;
input v_635;
input v_636;
input v_637;
input v_638;
input v_639;
input v_640;
input v_641;
input v_642;
input v_643;
input v_644;
input v_645;
input v_646;
input v_647;
input v_648;
input v_649;
input v_650;
input v_651;
input v_652;
input v_653;
input v_654;
input v_655;
input v_656;
input v_657;
input v_658;
input v_659;
input v_660;
input v_661;
input v_662;
input v_663;
input v_664;
input v_686;
input v_687;
input v_688;
input v_689;
input v_690;
input v_691;
input v_692;
input v_693;
input v_694;
input v_695;
input v_696;
input v_697;
input v_698;
input v_699;
input v_700;
input v_701;
input v_702;
input v_703;
input v_704;
input v_705;
input v_706;
input v_707;
input v_708;
input v_709;
input v_710;
input v_711;
input v_712;
input v_713;
input v_714;
input v_715;
input v_716;
input v_717;
input v_718;
input v_719;
input v_720;
input v_721;
input v_722;
input v_723;
input v_724;
input v_725;
input v_726;
input v_727;
input v_728;
input v_729;
input v_730;
input v_731;
input v_732;
input v_733;
input v_734;
input v_735;
input v_736;
input v_737;
input v_738;
input v_739;
input v_740;
input v_741;
input v_742;
input v_743;
input v_744;
input v_745;
input v_746;
input v_747;
input v_748;
input v_749;
input v_750;
input v_751;
input v_752;
input v_753;
input v_754;
input v_755;
input v_756;
input v_757;
input v_758;
input v_759;
input v_760;
input v_761;
input v_762;
input v_763;
input v_764;
input v_765;
input v_766;
input v_767;
input v_768;
input v_769;
input v_770;
input v_792;
input v_793;
input v_794;
input v_795;
input v_796;
input v_797;
input v_798;
input v_799;
input v_800;
input v_801;
input v_802;
input v_803;
input v_804;
input v_805;
input v_806;
input v_807;
input v_808;
input v_809;
input v_810;
input v_811;
input v_812;
input v_813;
input v_814;
input v_815;
input v_816;
input v_817;
input v_818;
input v_819;
input v_820;
input v_821;
input v_822;
input v_823;
input v_824;
input v_825;
input v_826;
input v_827;
input v_828;
input v_829;
input v_830;
input v_831;
input v_832;
input v_833;
input v_834;
input v_835;
input v_836;
input v_837;
input v_838;
input v_839;
input v_840;
input v_841;
input v_842;
input v_843;
input v_844;
input v_845;
input v_846;
input v_847;
input v_848;
input v_849;
input v_850;
input v_851;
input v_852;
input v_853;
input v_854;
input v_855;
input v_856;
input v_857;
input v_858;
input v_859;
input v_860;
input v_861;
input v_862;
input v_863;
input v_864;
input v_865;
input v_866;
input v_867;
input v_868;
input v_869;
input v_870;
input v_871;
input v_872;
input v_873;
input v_874;
input v_875;
input v_876;
input v_877;
input v_878;
input v_879;
input v_880;
input v_881;
input v_882;
input v_883;
input v_884;
input v_885;
input v_886;
input v_887;
input v_888;
input v_889;
input v_890;
input v_891;
input v_892;
input v_893;
input v_894;
input v_895;
input v_896;
input v_897;
input v_898;
input v_899;
input v_900;
input v_901;
input v_902;
input v_903;
input v_904;
input v_905;
input v_906;
input v_907;
input v_908;
input v_909;
input v_910;
input v_911;
input v_912;
input v_913;
input v_914;
input v_915;
input v_916;
input v_917;
input v_918;
input v_919;
input v_920;
input v_921;
input v_922;
input v_923;
input v_924;
input v_925;
input v_926;
input v_927;
input v_928;
input v_929;
input v_930;
input v_931;
input v_932;
input v_933;
input v_934;
input v_935;
input v_936;
input v_937;
input v_938;
input v_939;
input v_940;
input v_941;
input v_942;
input v_943;
input v_944;
input v_945;
input v_946;
input v_947;
input v_948;
input v_949;
input v_950;
input v_951;
input v_952;
input v_953;
input v_954;
input v_955;
input v_956;
input v_957;
input v_958;
input v_959;
input v_960;
input v_961;
input v_962;
input v_963;
input v_964;
input v_965;
input v_966;
input v_967;
input v_968;
input v_969;
input v_970;
input v_971;
input v_972;
input v_973;
input v_974;
input v_975;
input v_976;
input v_977;
input v_978;
input v_979;
input v_980;
input v_981;
input v_982;
input v_983;
input v_984;
input v_985;
input v_986;
input v_987;
input v_988;
input v_989;
input v_990;
input v_991;
input v_992;
input v_993;
input v_994;
input v_995;
input v_996;
input v_997;
input v_998;
input v_999;
input v_1000;
input v_1001;
input v_1002;
input v_1003;
input v_1004;
input v_1005;
input v_1006;
input v_1007;
input v_1008;
input v_1009;
input v_1010;
input v_1011;
input v_1012;
input v_1013;
input v_1014;
input v_1015;
input v_1016;
input v_1017;
input v_1018;
input v_1019;
input v_1020;
input v_1021;
input v_1022;
input v_1023;
input v_1024;
input v_1025;
input v_1026;
input v_1027;
input v_1028;
input v_1029;
input v_1030;
input v_1031;
input v_1032;
input v_1033;
input v_1034;
input v_1035;
input v_1036;
input v_1037;
input v_1038;
input v_1039;
input v_1040;
input v_1041;
input v_1042;
input v_1043;
input v_1044;
input v_1045;
input v_1046;
input v_1047;
input v_1048;
input v_1049;
input v_1050;
input v_1051;
input v_1052;
input v_1053;
input v_1054;
input v_1055;
input v_1056;
input v_1057;
input v_1058;
input v_1059;
input v_1060;
input v_1061;
input v_1062;
input v_1063;
input v_1064;
input v_1065;
input v_1066;
input v_1067;
input v_1068;
input v_1069;
input v_1070;
input v_1071;
input v_1072;
input v_1073;
input v_1074;
input v_1075;
input v_1076;
input v_1077;
input v_1078;
input v_1079;
input v_1080;
input v_1081;
input v_1082;
input v_1083;
input v_1084;
input v_1085;
input v_1086;
input v_1087;
input v_1088;
input v_1089;
input v_1090;
input v_1091;
input v_1092;
input v_1093;
input v_1094;
input v_1095;
input v_1096;
input v_1097;
input v_1098;
input v_1099;
input v_1100;
input v_1101;
input v_1102;
input v_1103;
input v_1104;
input v_1105;
input v_1106;
input v_1107;
input v_1108;
input v_1109;
input v_1110;
input v_1111;
input v_1112;
input v_1113;
input v_1114;
input v_1115;
input v_1116;
input v_1117;
input v_1118;
input v_1119;
input v_1120;
input v_1121;
input v_1122;
input v_1123;
input v_1124;
input v_1125;
input v_1126;
input v_1127;
input v_1128;
input v_1129;
input v_1130;
input v_1131;
input v_1132;
input v_1133;
input v_1134;
input v_1135;
input v_1136;
input v_1137;
input v_1138;
input v_1139;
input v_1140;
input v_1141;
input v_1142;
input v_1143;
input v_1144;
input v_1145;
input v_1146;
input v_1147;
input v_1148;
input v_1149;
input v_1150;
input v_1151;
input v_1152;
input v_1153;
input v_1154;
input v_1155;
input v_1156;
input v_1157;
input v_1158;
input v_1159;
input v_1160;
input v_1161;
input v_1162;
input v_1163;
input v_1164;
input v_1165;
input v_1166;
input v_1167;
input v_1168;
input v_1169;
input v_1170;
input v_1171;
input v_1172;
input v_1173;
input v_1174;
input v_1175;
input v_1176;
input v_1177;
input v_1178;
input v_1179;
input v_1180;
input v_1181;
input v_1182;
input v_1183;
input v_1184;
input v_1185;
input v_1186;
input v_1187;
input v_1188;
input v_1189;
input v_1190;
input v_1191;
input v_1192;
input v_1193;
input v_1194;
input v_1195;
input v_1196;
input v_1197;
input v_1198;
input v_1199;
input v_1200;
input v_1201;
input v_1202;
input v_1203;
input v_1204;
input v_1205;
input v_1206;
input v_1207;
input v_1208;
input v_1209;
input v_1210;
input v_1211;
input v_1212;
input v_1213;
input v_1214;
input v_1215;
input v_1216;
input v_1217;
input v_1218;
input v_1219;
input v_1220;
input v_1221;
input v_1222;
input v_1223;
input v_1224;
input v_1225;
input v_1226;
input v_1227;
input v_1228;
input v_1229;
input v_1230;
input v_1231;
input v_1232;
input v_1233;
input v_1234;
input v_1235;
input v_1236;
input v_1237;
input v_1238;
input v_1239;
input v_1240;
input v_1241;
input v_1242;
input v_1243;
input v_1244;
input v_1245;
input v_1246;
input v_1247;
input v_1248;
input v_1249;
input v_1250;
input v_1251;
input v_1252;
input v_1253;
input v_1254;
input v_1255;
input v_1256;
input v_1257;
input v_1258;
input v_1259;
input v_1260;
input v_1261;
input v_1262;
input v_1263;
input v_1264;
input v_1265;
input v_1266;
input v_1267;
input v_1268;
input v_1269;
input v_1270;
input v_1271;
input v_1272;
input v_1273;
input v_1274;
input v_1275;
input v_1276;
input v_1277;
input v_1278;
input v_1279;
input v_1280;
input v_1281;
input v_1282;
input v_1283;
input v_1284;
input v_1285;
input v_1286;
input v_1287;
input v_1288;
input v_1289;
input v_1290;
input v_1291;
input v_1292;
input v_1293;
input v_1294;
input v_1295;
input v_1296;
input v_1297;
input v_1298;
input v_1299;
input v_1300;
input v_1301;
input v_1302;
input v_1303;
input v_1304;
input v_1305;
input v_1306;
input v_1307;
input v_1308;
input v_1309;
input v_1310;
input v_1311;
input v_1312;
input v_1313;
input v_1314;
input v_1315;
input v_1316;
input v_1317;
input v_1318;
input v_1319;
input v_1320;
input v_1321;
input v_1322;
input v_1323;
input v_1324;
input v_1325;
input v_1326;
input v_1327;
input v_1328;
input v_1329;
input v_1330;
input v_1331;
input v_1332;
input v_1333;
input v_1334;
input v_1335;
input v_1336;
input v_1337;
input v_1338;
input v_1339;
input v_1340;
input v_1341;
input v_1342;
input v_1343;
input v_1344;
input v_1345;
input v_1346;
input v_1347;
input v_1348;
input v_1349;
input v_1350;
input v_1351;
input v_1352;
input v_1353;
input v_1354;
input v_1355;
input v_1356;
input v_1357;
input v_1358;
input v_1359;
input v_1360;
input v_1361;
input v_1362;
input v_1363;
input v_1364;
input v_1365;
input v_1366;
input v_1367;
input v_1368;
input v_1369;
input v_1370;
input v_1371;
input v_1372;
input v_1373;
input v_1374;
input v_1375;
input v_1376;
input v_1377;
input v_1378;
input v_1379;
input v_1380;
input v_1381;
input v_1382;
input v_1383;
input v_1384;
input v_1385;
input v_1386;
input v_1387;
input v_1388;
input v_1389;
input v_1390;
input v_1391;
input v_1392;
input v_1393;
input v_1394;
input v_1395;
input v_1396;
input v_1397;
input v_1398;
input v_1399;
input v_1400;
input v_1401;
input v_1402;
input v_1403;
input v_1404;
input v_1405;
input v_1406;
input v_1407;
input v_1408;
input v_1409;
input v_1410;
input v_1411;
input v_1412;
input v_1413;
input v_1414;
input v_1415;
input v_1416;
input v_1417;
input v_1418;
input v_1419;
input v_1420;
input v_1421;
input v_1422;
input v_1423;
input v_1424;
input v_1425;
input v_1426;
input v_1427;
input v_1428;
input v_1429;
input v_1430;
input v_1431;
input v_1432;
input v_1433;
input v_1434;
input v_1435;
input v_1436;
input v_1437;
input v_1438;
input v_1439;
input v_1440;
input v_1441;
input v_1442;
input v_1443;
input v_1444;
input v_1445;
input v_1446;
input v_1447;
input v_1448;
input v_1449;
input v_1450;
input v_1451;
input v_1452;
input v_1453;
input v_1454;
input v_1455;
input v_1456;
input v_1457;
input v_1458;
input v_1459;
input v_1460;
input v_1461;
input v_1462;
input v_1463;
input v_1464;
input v_1465;
input v_1466;
input v_1467;
input v_1468;
input v_1469;
input v_1470;
input v_1471;
input v_1472;
input v_1473;
input v_1474;
input v_1475;
input v_1476;
input v_1477;
input v_1478;
input v_1479;
input v_1480;
input v_1481;
input v_1482;
input v_1483;
input v_1484;
input v_1485;
input v_1486;
input v_1487;
input v_1488;
input v_1489;
input v_1490;
input v_1491;
input v_1492;
input v_1493;
input v_1494;
input v_1495;
input v_1496;
input v_1497;
input v_1498;
input v_1499;
input v_1500;
input v_1501;
input v_1502;
input v_1503;
input v_1504;
input v_1505;
input v_1506;
input v_1507;
input v_1508;
input v_1509;
input v_1510;
input v_1511;
input v_1512;
input v_1513;
input v_1514;
input v_1515;
input v_1516;
input v_1517;
input v_1518;
input v_1519;
input v_1520;
input v_1521;
input v_1522;
input v_1523;
input v_1524;
input v_1525;
input v_1526;
input v_1527;
input v_1528;
input v_1529;
input v_1530;
input v_1531;
input v_1532;
input v_1533;
input v_1534;
input v_1535;
input v_1536;
input v_1537;
input v_1538;
input v_1539;
input v_1540;
input v_1541;
input v_1542;
input v_1543;
input v_1544;
input v_1545;
input v_1546;
input v_1547;
input v_1548;
input v_1549;
input v_1550;
input v_1551;
input v_1552;
input v_1553;
input v_1554;
input v_1555;
input v_1556;
input v_1557;
input v_1558;
input v_1559;
input v_1560;
input v_1561;
input v_1562;
input v_1563;
input v_1564;
input v_1565;
input v_1566;
input v_1567;
input v_1568;
input v_1569;
input v_1570;
input v_1571;
input v_1572;
input v_1573;
input v_1574;
input v_1575;
input v_1576;
input v_1577;
input v_1578;
input v_1579;
input v_1580;
input v_1581;
input v_1582;
input v_1583;
input v_1584;
input v_1585;
input v_1586;
input v_1587;
input v_1588;
input v_1589;
input v_1590;
input v_1591;
input v_1592;
input v_1593;
input v_1594;
input v_1595;
input v_1596;
input v_1597;
input v_1598;
input v_1599;
input v_1600;
input v_1601;
input v_1602;
input v_1603;
input v_1604;
input v_1605;
input v_1606;
input v_1607;
input v_1608;
input v_1609;
input v_1610;
input v_1611;
input v_1612;
input v_1613;
input v_1614;
input v_1615;
input v_1616;
input v_1617;
input v_1618;
input v_1619;
input v_1620;
input v_1621;
input v_1622;
input v_1623;
input v_1624;
input v_1625;
input v_1626;
input v_1627;
input v_1628;
input v_1629;
input v_1630;
input v_1631;
input v_1632;
input v_1633;
input v_1634;
input v_1635;
input v_1636;
input v_1637;
input v_1638;
input v_1639;
input v_1640;
input v_1641;
input v_1642;
input v_1643;
input v_1644;
input v_1645;
input v_1646;
input v_1647;
input v_1648;
input v_1649;
input v_1650;
input v_1651;
input v_1652;
input v_1653;
input v_1654;
input v_1655;
input v_1656;
input v_1657;
input v_1658;
input v_1659;
input v_1660;
input v_1661;
input v_1662;
input v_1663;
input v_1664;
input v_1665;
input v_1666;
input v_1667;
input v_1668;
input v_1669;
input v_1670;
input v_1671;
input v_1672;
input v_1673;
input v_1674;
input v_1675;
input v_1676;
input v_1677;
input v_1678;
input v_1679;
input v_1680;
input v_1681;
input v_1682;
input v_1683;
input v_1684;
input v_1685;
input v_1686;
input v_1687;
input v_1688;
input v_1689;
input v_1690;
input v_1691;
input v_1692;
input v_1693;
input v_1694;
input v_1695;
input v_1696;
input v_1697;
input v_1698;
input v_1699;
input v_1700;
input v_1701;
input v_1702;
input v_1703;
input v_1704;
input v_1705;
input v_1706;
input v_1707;
input v_1708;
input v_1709;
input v_1710;
input v_1711;
input v_1712;
input v_1713;
input v_1714;
input v_1715;
input v_1716;
input v_1717;
input v_1718;
input v_1719;
input v_1720;
input v_1721;
input v_1722;
input v_1723;
input v_1724;
input v_1725;
input v_1726;
input v_1727;
input v_1728;
input v_1729;
input v_1730;
input v_1731;
input v_1732;
input v_1733;
input v_1734;
input v_1735;
input v_1736;
input v_1737;
input v_1738;
input v_1739;
input v_1740;
input v_1741;
input v_1742;
input v_1743;
input v_1744;
input v_1745;
input v_1746;
input v_1747;
input v_1748;
input v_1749;
input v_1750;
input v_1751;
input v_1752;
input v_1753;
input v_1754;
input v_1755;
input v_1756;
input v_1757;
input v_1758;
input v_1759;
input v_1760;
input v_1761;
input v_1762;
input v_1763;
input v_1764;
input v_1765;
input v_1766;
input v_1767;
input v_1768;
input v_1769;
input v_1770;
input v_1771;
input v_1772;
input v_1773;
input v_1774;
input v_1775;
input v_1776;
input v_1777;
input v_1778;
input v_1779;
input v_1780;
input v_1781;
input v_1782;
input v_1783;
input v_1784;
input v_1785;
input v_1786;
input v_1787;
input v_1788;
input v_1789;
input v_1790;
input v_1791;
input v_1792;
input v_1793;
input v_1794;
input v_1795;
input v_1796;
input v_1797;
input v_1798;
input v_1799;
input v_1800;
input v_1801;
input v_1802;
input v_1803;
input v_1804;
input v_1805;
input v_1806;
input v_1807;
input v_1808;
input v_1809;
input v_1810;
input v_1811;
input v_1812;
input v_1813;
input v_1814;
input v_1815;
input v_1816;
input v_1817;
input v_1818;
input v_1819;
input v_1820;
input v_1821;
input v_1822;
input v_1823;
input v_1824;
input v_1825;
input v_1826;
input v_1827;
input v_1828;
input v_1829;
input v_1830;
input v_1831;
input v_1832;
input v_1833;
input v_1834;
input v_1835;
input v_1836;
input v_1837;
input v_1838;
input v_1839;
input v_1840;
input v_1841;
input v_1842;
input v_1903;
input v_1904;
input v_1905;
input v_1906;
input v_1907;
input v_1908;
input v_1909;
input v_1910;
input v_1911;
input v_1912;
input v_1913;
input v_1914;
input v_1915;
input v_1916;
input v_1917;
input v_1918;
input v_1919;
input v_1920;
input v_1921;
input v_1922;
input v_1923;
input v_1924;
input v_1925;
input v_1926;
input v_1927;
input v_1928;
input v_1929;
input v_1930;
input v_1931;
input v_1932;
input v_1933;
input v_1934;
input v_1935;
input v_1936;
input v_1937;
input v_1938;
input v_1939;
input v_1940;
input v_1941;
input v_1942;
input v_1943;
input v_1944;
input v_2005;
input v_2006;
input v_2007;
input v_2008;
input v_2009;
input v_2010;
input v_2011;
input v_2012;
input v_2013;
input v_2014;
input v_2015;
input v_2016;
input v_2017;
input v_2018;
input v_2019;
input v_2020;
input v_2021;
input v_2022;
input v_2023;
input v_2024;
input v_2025;
input v_2026;
input v_2027;
input v_2028;
input v_2029;
input v_2030;
input v_2031;
input v_2032;
input v_2033;
input v_2034;
input v_2035;
input v_2036;
input v_2037;
input v_2038;
input v_2039;
input v_2040;
input v_2041;
input v_2042;
input v_2043;
input v_2044;
input v_2045;
input v_2046;
input v_2107;
input v_2108;
input v_2109;
input v_2110;
input v_2111;
input v_2112;
input v_2113;
input v_2114;
input v_2115;
input v_2116;
input v_2117;
input v_2118;
input v_2119;
input v_2120;
input v_2121;
input v_2122;
input v_2123;
input v_2124;
input v_2125;
input v_2126;
input v_2127;
input v_2128;
input v_2129;
input v_2130;
input v_2131;
input v_2132;
input v_2133;
input v_2134;
input v_2135;
input v_2136;
input v_2137;
input v_2138;
input v_2139;
input v_2140;
input v_2141;
input v_2142;
input v_2143;
input v_2144;
input v_2145;
input v_2146;
input v_2147;
input v_2148;
input v_2209;
input v_2210;
input v_2211;
input v_2212;
input v_2213;
input v_2214;
input v_2215;
input v_2216;
input v_2217;
input v_2218;
input v_2219;
input v_2220;
input v_2221;
input v_2222;
input v_2223;
input v_2224;
input v_2225;
input v_2226;
input v_2227;
input v_2228;
input v_2229;
input v_2230;
input v_2231;
input v_2232;
input v_2233;
input v_2234;
input v_2235;
input v_2236;
input v_2237;
input v_2238;
input v_2239;
input v_2240;
input v_2241;
input v_2242;
input v_2243;
input v_2244;
input v_2245;
input v_2246;
input v_2247;
input v_2248;
input v_2249;
input v_2250;
output o_1;
wire v_347;
wire v_348;
wire v_349;
wire v_350;
wire v_351;
wire v_352;
wire v_353;
wire v_354;
wire v_355;
wire v_356;
wire v_357;
wire v_358;
wire v_359;
wire v_360;
wire v_361;
wire v_362;
wire v_363;
wire v_364;
wire v_365;
wire v_366;
wire v_367;
wire v_453;
wire v_454;
wire v_455;
wire v_456;
wire v_457;
wire v_458;
wire v_459;
wire v_460;
wire v_461;
wire v_462;
wire v_463;
wire v_464;
wire v_465;
wire v_466;
wire v_467;
wire v_468;
wire v_469;
wire v_470;
wire v_471;
wire v_472;
wire v_473;
wire v_559;
wire v_560;
wire v_561;
wire v_562;
wire v_563;
wire v_564;
wire v_565;
wire v_566;
wire v_567;
wire v_568;
wire v_569;
wire v_570;
wire v_571;
wire v_572;
wire v_573;
wire v_574;
wire v_575;
wire v_576;
wire v_577;
wire v_578;
wire v_579;
wire v_665;
wire v_666;
wire v_667;
wire v_668;
wire v_669;
wire v_670;
wire v_671;
wire v_672;
wire v_673;
wire v_674;
wire v_675;
wire v_676;
wire v_677;
wire v_678;
wire v_679;
wire v_680;
wire v_681;
wire v_682;
wire v_683;
wire v_684;
wire v_685;
wire v_771;
wire v_772;
wire v_773;
wire v_774;
wire v_775;
wire v_776;
wire v_777;
wire v_778;
wire v_779;
wire v_780;
wire v_781;
wire v_782;
wire v_783;
wire v_784;
wire v_785;
wire v_786;
wire v_787;
wire v_788;
wire v_789;
wire v_790;
wire v_791;
wire x_1;
wire x_2;
wire x_3;
wire x_4;
wire x_5;
wire x_6;
wire x_7;
wire x_8;
wire x_9;
wire x_10;
wire x_11;
wire x_12;
wire x_13;
wire x_14;
wire x_15;
wire x_16;
wire x_17;
wire x_18;
wire x_19;
wire x_20;
wire x_21;
wire x_22;
wire x_23;
wire x_24;
wire x_25;
wire x_26;
wire x_27;
wire x_28;
wire x_29;
wire x_30;
wire x_31;
wire x_32;
wire x_33;
wire x_34;
wire x_35;
wire x_36;
wire x_37;
wire x_38;
wire x_39;
wire x_40;
wire x_41;
wire x_42;
wire x_43;
wire x_44;
wire x_45;
wire x_46;
wire x_47;
wire x_48;
wire x_49;
wire x_50;
wire x_51;
wire x_52;
wire x_53;
wire x_54;
wire x_55;
wire x_56;
wire x_57;
wire x_58;
wire x_59;
wire x_60;
wire x_61;
wire x_62;
wire x_63;
wire x_64;
wire x_65;
wire x_66;
wire x_67;
wire x_68;
wire x_69;
wire x_70;
wire x_71;
wire x_72;
wire x_73;
wire x_74;
wire x_75;
wire x_76;
wire x_77;
wire x_78;
wire x_79;
wire x_80;
wire x_81;
wire x_82;
wire x_83;
wire x_84;
wire x_85;
wire x_86;
wire x_87;
wire x_88;
wire x_89;
wire x_90;
wire x_91;
wire x_92;
wire x_93;
wire x_94;
wire x_95;
wire x_96;
wire x_97;
wire x_98;
wire x_99;
wire x_100;
wire x_101;
wire x_102;
wire x_103;
wire x_104;
wire x_105;
wire x_106;
wire x_107;
wire x_108;
wire x_109;
wire x_110;
wire x_111;
wire x_112;
wire x_113;
wire x_114;
wire x_115;
wire x_116;
wire x_117;
wire x_118;
wire x_119;
wire x_120;
wire x_121;
wire x_122;
wire x_123;
wire x_124;
wire x_125;
wire x_126;
wire x_127;
wire x_128;
wire x_129;
wire x_130;
wire x_131;
wire x_132;
wire x_133;
wire x_134;
wire x_135;
wire x_136;
wire x_137;
wire x_138;
wire x_139;
wire x_140;
wire x_141;
wire x_142;
wire x_143;
wire x_144;
wire x_145;
wire x_146;
wire x_147;
wire x_148;
wire x_149;
wire x_150;
wire x_151;
wire x_152;
wire x_153;
wire x_154;
wire x_155;
wire x_156;
wire x_157;
wire x_158;
wire x_159;
wire x_160;
wire x_161;
wire x_162;
wire x_163;
wire x_164;
wire x_165;
wire x_166;
wire x_167;
wire x_168;
wire x_169;
wire x_170;
wire x_171;
wire x_172;
wire x_173;
wire x_174;
wire x_175;
wire x_176;
wire x_177;
wire x_178;
wire x_179;
wire x_180;
wire x_181;
wire x_182;
wire x_183;
wire x_184;
wire x_185;
wire x_186;
wire x_187;
wire x_188;
wire x_189;
wire x_190;
wire x_191;
wire x_192;
wire x_193;
wire x_194;
wire x_195;
wire x_196;
wire x_197;
wire x_198;
wire x_199;
wire x_200;
wire x_201;
wire x_202;
wire x_203;
wire x_204;
wire x_205;
wire x_206;
wire x_207;
wire x_208;
wire x_209;
wire x_210;
wire x_211;
wire x_212;
wire x_213;
wire x_214;
wire x_215;
wire x_216;
wire x_217;
wire x_218;
wire x_219;
wire x_220;
wire x_221;
wire x_222;
wire x_223;
wire x_224;
wire x_225;
wire x_226;
wire x_227;
wire x_228;
wire x_229;
wire x_230;
wire x_231;
wire x_232;
wire x_233;
wire x_234;
wire x_235;
wire x_236;
wire x_237;
wire x_238;
wire x_239;
wire x_240;
wire x_241;
wire x_242;
wire x_243;
wire x_244;
wire x_245;
wire x_246;
wire x_247;
wire x_248;
wire x_249;
wire x_250;
wire x_251;
wire x_252;
wire x_253;
wire x_254;
wire x_255;
wire x_256;
wire x_257;
wire x_258;
wire x_259;
wire x_260;
wire x_261;
wire x_262;
wire x_263;
wire x_264;
wire x_265;
wire x_266;
wire x_267;
wire x_268;
wire x_269;
wire x_270;
wire x_271;
wire x_272;
wire x_273;
wire x_274;
wire x_275;
wire x_276;
wire x_277;
wire x_278;
wire x_279;
wire x_280;
wire x_281;
wire x_282;
wire x_283;
wire x_284;
wire x_285;
wire x_286;
wire x_287;
wire x_288;
wire x_289;
wire x_290;
wire x_291;
wire x_292;
wire x_293;
wire x_294;
wire x_295;
wire x_296;
wire x_297;
wire x_298;
wire x_299;
wire x_300;
wire x_301;
wire x_302;
wire x_303;
wire x_304;
wire x_305;
wire x_306;
wire x_307;
wire x_308;
wire x_309;
wire x_310;
wire x_311;
wire x_312;
wire x_313;
wire x_314;
wire x_315;
wire x_316;
wire x_317;
wire x_318;
wire x_319;
wire x_320;
wire x_321;
wire x_322;
wire x_323;
wire x_324;
wire x_325;
wire x_326;
wire x_327;
wire x_328;
wire x_329;
wire x_330;
wire x_331;
wire x_332;
wire x_333;
wire x_334;
wire x_335;
wire x_336;
wire x_337;
wire x_338;
wire x_339;
wire x_340;
wire x_341;
wire x_342;
wire x_343;
wire x_344;
wire x_345;
wire x_346;
wire x_347;
wire x_348;
wire x_349;
wire x_350;
wire x_351;
wire x_352;
wire x_353;
wire x_354;
wire x_355;
wire x_356;
wire x_357;
wire x_358;
wire x_359;
wire x_360;
wire x_361;
wire x_362;
wire x_363;
wire x_364;
wire x_365;
wire x_366;
wire x_367;
wire x_368;
wire x_369;
wire x_370;
wire x_371;
wire x_372;
wire x_373;
wire x_374;
wire x_375;
wire x_376;
wire x_377;
wire x_378;
wire x_379;
wire x_380;
wire x_381;
wire x_382;
wire x_383;
wire x_384;
wire x_385;
wire x_386;
wire x_387;
wire x_388;
wire x_389;
wire x_390;
wire x_391;
wire x_392;
wire x_393;
wire x_394;
wire x_395;
wire x_396;
wire x_397;
wire x_398;
wire x_399;
wire x_400;
wire x_401;
wire x_402;
wire x_403;
wire x_404;
wire x_405;
wire x_406;
wire x_407;
wire x_408;
wire x_409;
wire x_410;
wire x_411;
wire x_412;
wire x_413;
wire x_414;
wire x_415;
wire x_416;
wire x_417;
wire x_418;
wire x_419;
wire x_420;
wire x_421;
wire x_422;
wire x_423;
wire x_424;
wire x_425;
wire x_426;
wire x_427;
wire x_428;
wire x_429;
wire x_430;
wire x_431;
wire x_432;
wire x_433;
wire x_434;
wire x_435;
wire x_436;
wire x_437;
wire x_438;
wire x_439;
wire x_440;
wire x_441;
wire x_442;
wire x_443;
wire x_444;
wire x_445;
wire x_446;
wire x_447;
wire x_448;
wire x_449;
wire x_450;
wire x_451;
wire x_452;
wire x_453;
wire x_454;
wire x_455;
wire x_456;
wire x_457;
wire x_458;
wire x_459;
wire x_460;
wire x_461;
wire x_462;
wire x_463;
wire x_464;
wire x_465;
wire x_466;
wire x_467;
wire x_468;
wire x_469;
wire x_470;
wire x_471;
wire x_472;
wire x_473;
wire x_474;
wire x_475;
wire x_476;
wire x_477;
wire x_478;
wire x_479;
wire x_480;
wire x_481;
wire x_482;
wire x_483;
wire x_484;
wire x_485;
wire x_486;
wire x_487;
wire x_488;
wire x_489;
wire x_490;
wire x_491;
wire x_492;
wire x_493;
wire x_494;
wire x_495;
wire x_496;
wire x_497;
wire x_498;
wire x_499;
wire x_500;
wire x_501;
wire x_502;
wire x_503;
wire x_504;
wire x_505;
wire x_506;
wire x_507;
wire x_508;
wire x_509;
wire x_510;
wire x_511;
wire x_512;
wire x_513;
wire x_514;
wire x_515;
wire x_516;
wire x_517;
wire x_518;
wire x_519;
wire x_520;
wire x_521;
wire x_522;
wire x_523;
wire x_524;
wire x_525;
wire x_526;
wire x_527;
wire x_528;
wire x_529;
wire x_530;
wire x_531;
wire x_532;
wire x_533;
wire x_534;
wire x_535;
wire x_536;
wire x_537;
wire x_538;
wire x_539;
wire x_540;
wire x_541;
wire x_542;
wire x_543;
wire x_544;
wire x_545;
wire x_546;
wire x_547;
wire x_548;
wire x_549;
wire x_550;
wire x_551;
wire x_552;
wire x_553;
wire x_554;
wire x_555;
wire x_556;
wire x_557;
wire x_558;
wire x_559;
wire x_560;
wire x_561;
wire x_562;
wire x_563;
wire x_564;
wire x_565;
wire x_566;
wire x_567;
wire x_568;
wire x_569;
wire x_570;
wire x_571;
wire x_572;
wire x_573;
wire x_574;
wire x_575;
wire x_576;
wire x_577;
wire x_578;
wire x_579;
wire x_580;
wire x_581;
wire x_582;
wire x_583;
wire x_584;
wire x_585;
wire x_586;
wire x_587;
wire x_588;
wire x_589;
wire x_590;
wire x_591;
wire x_592;
wire x_593;
wire x_594;
wire x_595;
wire x_596;
wire x_597;
wire x_598;
wire x_599;
wire x_600;
wire x_601;
wire x_602;
wire x_603;
wire x_604;
wire x_605;
wire x_606;
wire x_607;
wire x_608;
wire x_609;
wire x_610;
wire x_611;
wire x_612;
wire x_613;
wire x_614;
wire x_615;
wire x_616;
wire x_617;
wire x_618;
wire x_619;
wire x_620;
wire x_621;
wire x_622;
wire x_623;
wire x_624;
wire x_625;
wire x_626;
wire x_627;
wire x_628;
wire x_629;
wire x_630;
wire x_631;
wire x_632;
wire x_633;
wire x_634;
wire x_635;
wire x_636;
wire x_637;
wire x_638;
wire x_639;
wire x_640;
wire x_641;
wire x_642;
wire x_643;
wire x_644;
wire x_645;
wire x_646;
wire x_647;
wire x_648;
wire x_649;
wire x_650;
wire x_651;
wire x_652;
wire x_653;
wire x_654;
wire x_655;
wire x_656;
wire x_657;
wire x_658;
wire x_659;
wire x_660;
wire x_661;
wire x_662;
wire x_663;
wire x_664;
wire x_665;
wire x_666;
wire x_667;
wire x_668;
wire x_669;
wire x_670;
wire x_671;
wire x_672;
wire x_673;
wire x_674;
wire x_675;
wire x_676;
wire x_677;
wire x_678;
wire x_679;
wire x_680;
wire x_681;
wire x_682;
wire x_683;
wire x_684;
wire x_685;
wire x_686;
wire x_687;
wire x_688;
wire x_689;
wire x_690;
wire x_691;
wire x_692;
wire x_693;
wire x_694;
wire x_695;
wire x_696;
wire x_697;
wire x_698;
wire x_699;
wire x_700;
wire x_701;
wire x_702;
wire x_703;
wire x_704;
wire x_705;
wire x_706;
wire x_707;
wire x_708;
wire x_709;
wire x_710;
wire x_711;
wire x_712;
wire x_713;
wire x_714;
wire x_715;
wire x_716;
wire x_717;
wire x_718;
wire x_719;
wire x_720;
wire x_721;
wire x_722;
wire x_723;
wire x_724;
wire x_725;
wire x_726;
wire x_727;
wire x_728;
wire x_729;
wire x_730;
wire x_731;
wire x_732;
wire x_733;
wire x_734;
wire x_735;
wire x_736;
wire x_737;
wire x_738;
wire x_739;
wire x_740;
wire x_741;
wire x_742;
wire x_743;
wire x_744;
wire x_745;
wire x_746;
wire x_747;
wire x_748;
wire x_749;
wire x_750;
wire x_751;
wire x_752;
wire x_753;
wire x_754;
wire x_755;
wire x_756;
wire x_757;
wire x_758;
wire x_759;
wire x_760;
wire x_761;
wire x_762;
wire x_763;
wire x_764;
wire x_765;
wire x_766;
wire x_767;
wire x_768;
wire x_769;
wire x_770;
wire x_771;
wire x_772;
wire x_773;
wire x_774;
wire x_775;
wire x_776;
wire x_777;
wire x_778;
wire x_779;
wire x_780;
wire x_781;
wire x_782;
wire x_783;
wire x_784;
wire x_785;
wire x_786;
wire x_787;
wire x_788;
wire x_789;
wire x_790;
wire x_791;
wire x_792;
wire x_793;
wire x_794;
wire x_795;
wire x_796;
wire x_797;
wire x_798;
wire x_799;
wire x_800;
wire x_801;
wire x_802;
wire x_803;
wire x_804;
wire x_805;
wire x_806;
wire x_807;
wire x_808;
wire x_809;
wire x_810;
wire x_811;
wire x_812;
wire x_813;
wire x_814;
wire x_815;
wire x_816;
wire x_817;
wire x_818;
wire x_819;
wire x_820;
wire x_821;
wire x_822;
wire x_823;
wire x_824;
wire x_825;
wire x_826;
wire x_827;
wire x_828;
wire x_829;
wire x_830;
wire x_831;
wire x_832;
wire x_833;
wire x_834;
wire x_835;
wire x_836;
wire x_837;
wire x_838;
wire x_839;
wire x_840;
wire x_841;
wire x_842;
wire x_843;
wire x_844;
wire x_845;
wire x_846;
wire x_847;
wire x_848;
wire x_849;
wire x_850;
wire x_851;
wire x_852;
wire x_853;
wire x_854;
wire x_855;
wire x_856;
wire x_857;
wire x_858;
wire x_859;
wire x_860;
wire x_861;
wire x_862;
wire x_863;
wire x_864;
wire x_865;
wire x_866;
wire x_867;
wire x_868;
wire x_869;
wire x_870;
wire x_871;
wire x_872;
wire x_873;
wire x_874;
wire x_875;
wire x_876;
wire x_877;
wire x_878;
wire x_879;
wire x_880;
wire x_881;
wire x_882;
wire x_883;
wire x_884;
wire x_885;
wire x_886;
wire x_887;
wire x_888;
wire x_889;
wire x_890;
wire x_891;
wire x_892;
wire x_893;
wire x_894;
wire x_895;
wire x_896;
wire x_897;
wire x_898;
wire x_899;
wire x_900;
wire x_901;
wire x_902;
wire x_903;
wire x_904;
wire x_905;
wire x_906;
wire x_907;
wire x_908;
wire x_909;
wire x_910;
wire x_911;
wire x_912;
wire x_913;
wire x_914;
wire x_915;
wire x_916;
wire x_917;
wire x_918;
wire x_919;
wire x_920;
wire x_921;
wire x_922;
wire x_923;
wire x_924;
wire x_925;
wire x_926;
wire x_927;
wire x_928;
wire x_929;
wire x_930;
wire x_931;
wire x_932;
wire x_933;
wire x_934;
wire x_935;
wire x_936;
wire x_937;
wire x_938;
wire x_939;
wire x_940;
wire x_941;
wire x_942;
wire x_943;
wire x_944;
wire x_945;
wire x_946;
wire x_947;
wire x_948;
wire x_949;
wire x_950;
wire x_951;
wire x_952;
wire x_953;
wire x_954;
wire x_955;
wire x_956;
wire x_957;
wire x_958;
wire x_959;
wire x_960;
wire x_961;
wire x_962;
wire x_963;
wire x_964;
wire x_965;
wire x_966;
wire x_967;
wire x_968;
wire x_969;
wire x_970;
wire x_971;
wire x_972;
wire x_973;
wire x_974;
wire x_975;
wire x_976;
wire x_977;
wire x_978;
wire x_979;
wire x_980;
wire x_981;
wire x_982;
wire x_983;
wire x_984;
wire x_985;
wire x_986;
wire x_987;
wire x_988;
wire x_989;
wire x_990;
wire x_991;
wire x_992;
wire x_993;
wire x_994;
wire x_995;
wire x_996;
wire x_997;
wire x_998;
wire x_999;
wire x_1000;
wire x_1001;
wire x_1002;
wire x_1003;
wire x_1004;
wire x_1005;
wire x_1006;
wire x_1007;
wire x_1008;
wire x_1009;
wire x_1010;
wire x_1011;
wire x_1012;
wire x_1013;
wire x_1014;
wire x_1015;
wire x_1016;
wire x_1017;
wire x_1018;
wire x_1019;
wire x_1020;
wire x_1021;
wire x_1022;
wire x_1023;
wire x_1024;
wire x_1025;
wire x_1026;
wire x_1027;
wire x_1028;
wire x_1029;
wire x_1030;
wire x_1031;
wire x_1032;
wire x_1033;
wire x_1034;
wire x_1035;
wire x_1036;
wire x_1037;
wire x_1038;
wire x_1039;
wire x_1040;
wire x_1041;
wire x_1042;
wire x_1043;
wire x_1044;
wire x_1045;
wire x_1046;
wire x_1047;
wire x_1048;
wire x_1049;
wire x_1050;
wire x_1051;
wire x_1052;
wire x_1053;
wire x_1054;
wire x_1055;
wire x_1056;
wire x_1057;
wire x_1058;
wire x_1059;
wire x_1060;
wire x_1061;
wire x_1062;
wire x_1063;
wire x_1064;
wire x_1065;
wire x_1066;
wire x_1067;
wire x_1068;
wire x_1069;
wire x_1070;
wire x_1071;
wire x_1072;
wire x_1073;
wire x_1074;
wire x_1075;
wire x_1076;
wire x_1077;
wire x_1078;
wire x_1079;
wire x_1080;
wire x_1081;
wire x_1082;
wire x_1083;
wire x_1084;
wire x_1085;
wire x_1086;
wire x_1087;
wire x_1088;
wire x_1089;
wire x_1090;
wire x_1091;
wire x_1092;
wire x_1093;
wire x_1094;
wire x_1095;
wire x_1096;
wire x_1097;
wire x_1098;
wire x_1099;
wire x_1100;
wire x_1101;
wire x_1102;
wire x_1103;
wire x_1104;
wire x_1105;
wire x_1106;
wire x_1107;
wire x_1108;
wire x_1109;
wire x_1110;
wire x_1111;
wire x_1112;
wire x_1113;
wire x_1114;
wire x_1115;
wire x_1116;
wire x_1117;
wire x_1118;
wire x_1119;
wire x_1120;
wire x_1121;
wire x_1122;
wire x_1123;
wire x_1124;
wire x_1125;
wire x_1126;
wire x_1127;
wire x_1128;
wire x_1129;
wire x_1130;
wire x_1131;
wire x_1132;
wire x_1133;
wire x_1134;
wire x_1135;
wire x_1136;
wire x_1137;
wire x_1138;
wire x_1139;
wire x_1140;
wire x_1141;
wire x_1142;
wire x_1143;
wire x_1144;
wire x_1145;
wire x_1146;
wire x_1147;
wire x_1148;
wire x_1149;
wire x_1150;
wire x_1151;
wire x_1152;
wire x_1153;
wire x_1154;
wire x_1155;
wire x_1156;
wire x_1157;
wire x_1158;
wire x_1159;
wire x_1160;
wire x_1161;
wire x_1162;
wire x_1163;
wire x_1164;
wire x_1165;
wire x_1166;
wire x_1167;
wire x_1168;
wire x_1169;
wire x_1170;
wire x_1171;
wire x_1172;
wire x_1173;
wire x_1174;
wire x_1175;
wire x_1176;
wire x_1177;
wire x_1178;
wire x_1179;
wire x_1180;
wire x_1181;
wire x_1182;
wire x_1183;
wire x_1184;
wire x_1185;
wire x_1186;
wire x_1187;
wire x_1188;
wire x_1189;
wire x_1190;
wire x_1191;
wire x_1192;
wire x_1193;
wire x_1194;
wire x_1195;
wire x_1196;
wire x_1197;
wire x_1198;
wire x_1199;
wire x_1200;
wire x_1201;
wire x_1202;
wire x_1203;
wire x_1204;
wire x_1205;
wire x_1206;
wire x_1207;
wire x_1208;
wire x_1209;
wire x_1210;
wire x_1211;
wire x_1212;
wire x_1213;
wire x_1214;
wire x_1215;
wire x_1216;
wire x_1217;
wire x_1218;
wire x_1219;
wire x_1220;
wire x_1221;
wire x_1222;
wire x_1223;
wire x_1224;
wire x_1225;
wire x_1226;
wire x_1227;
wire x_1228;
wire x_1229;
wire x_1230;
wire x_1231;
wire x_1232;
wire x_1233;
wire x_1234;
wire x_1235;
wire x_1236;
wire x_1237;
wire x_1238;
wire x_1239;
wire x_1240;
wire x_1241;
wire x_1242;
wire x_1243;
wire x_1244;
wire x_1245;
wire x_1246;
wire x_1247;
wire x_1248;
wire x_1249;
wire x_1250;
wire x_1251;
wire x_1252;
wire x_1253;
wire x_1254;
wire x_1255;
wire x_1256;
wire x_1257;
wire x_1258;
wire x_1259;
wire x_1260;
wire x_1261;
wire x_1262;
wire x_1263;
wire x_1264;
wire x_1265;
wire x_1266;
wire x_1267;
wire x_1268;
wire x_1269;
wire x_1270;
wire x_1271;
wire x_1272;
wire x_1273;
wire x_1274;
wire x_1275;
wire x_1276;
wire x_1277;
wire x_1278;
wire x_1279;
wire x_1280;
wire x_1281;
wire x_1282;
wire x_1283;
wire x_1284;
wire x_1285;
wire x_1286;
wire x_1287;
wire x_1288;
wire x_1289;
wire x_1290;
wire x_1291;
wire x_1292;
wire x_1293;
wire x_1294;
wire x_1295;
wire x_1296;
wire x_1297;
wire x_1298;
wire x_1299;
wire x_1300;
wire x_1301;
wire x_1302;
wire x_1303;
wire x_1304;
wire x_1305;
wire x_1306;
wire x_1307;
wire x_1308;
wire x_1309;
wire x_1310;
wire x_1311;
wire x_1312;
wire x_1313;
wire x_1314;
wire x_1315;
wire x_1316;
wire x_1317;
wire x_1318;
wire x_1319;
wire x_1320;
wire x_1321;
wire x_1322;
wire x_1323;
wire x_1324;
wire x_1325;
wire x_1326;
wire x_1327;
wire x_1328;
wire x_1329;
wire x_1330;
wire x_1331;
wire x_1332;
wire x_1333;
wire x_1334;
wire x_1335;
wire x_1336;
wire x_1337;
wire x_1338;
wire x_1339;
wire x_1340;
wire x_1341;
wire x_1342;
wire x_1343;
wire x_1344;
wire x_1345;
wire x_1346;
wire x_1347;
wire x_1348;
wire x_1349;
wire x_1350;
wire x_1351;
wire x_1352;
wire x_1353;
wire x_1354;
wire x_1355;
wire x_1356;
wire x_1357;
wire x_1358;
wire x_1359;
wire x_1360;
wire x_1361;
wire x_1362;
wire x_1363;
wire x_1364;
wire x_1365;
wire x_1366;
wire x_1367;
wire x_1368;
wire x_1369;
wire x_1370;
wire x_1371;
wire x_1372;
wire x_1373;
wire x_1374;
wire x_1375;
wire x_1376;
wire x_1377;
wire x_1378;
wire x_1379;
wire x_1380;
wire x_1381;
wire x_1382;
wire x_1383;
wire x_1384;
wire x_1385;
wire x_1386;
wire x_1387;
wire x_1388;
wire x_1389;
wire x_1390;
wire x_1391;
wire x_1392;
wire x_1393;
wire x_1394;
wire x_1395;
wire x_1396;
wire x_1397;
wire x_1398;
wire x_1399;
wire x_1400;
wire x_1401;
wire x_1402;
wire x_1403;
wire x_1404;
wire x_1405;
wire x_1406;
wire x_1407;
wire x_1408;
wire x_1409;
wire x_1410;
wire x_1411;
wire x_1412;
wire x_1413;
wire x_1414;
wire x_1415;
wire x_1416;
wire x_1417;
wire x_1418;
wire x_1419;
wire x_1420;
wire x_1421;
wire x_1422;
wire x_1423;
wire x_1424;
wire x_1425;
wire x_1426;
wire x_1427;
wire x_1428;
wire x_1429;
wire x_1430;
wire x_1431;
wire x_1432;
wire x_1433;
wire x_1434;
wire x_1435;
wire x_1436;
wire x_1437;
wire x_1438;
wire x_1439;
wire x_1440;
wire x_1441;
wire x_1442;
wire x_1443;
wire x_1444;
wire x_1445;
wire x_1446;
wire x_1447;
wire x_1448;
wire x_1449;
wire x_1450;
wire x_1451;
wire x_1452;
wire x_1453;
wire x_1454;
wire x_1455;
wire x_1456;
wire x_1457;
wire x_1458;
wire x_1459;
wire x_1460;
wire x_1461;
wire x_1462;
wire x_1463;
wire x_1464;
wire x_1465;
wire x_1466;
wire x_1467;
wire x_1468;
wire x_1469;
wire x_1470;
wire x_1471;
wire x_1472;
wire x_1473;
wire x_1474;
wire x_1475;
wire x_1476;
wire x_1477;
wire x_1478;
wire x_1479;
wire x_1480;
wire x_1481;
wire x_1482;
wire x_1483;
wire x_1484;
wire x_1485;
wire x_1486;
wire x_1487;
wire x_1488;
wire x_1489;
wire x_1490;
wire x_1491;
wire x_1492;
wire x_1493;
wire x_1494;
wire x_1495;
wire x_1496;
wire x_1497;
wire x_1498;
wire x_1499;
wire x_1500;
wire x_1501;
wire x_1502;
wire x_1503;
wire x_1504;
wire x_1505;
wire x_1506;
wire x_1507;
wire x_1508;
wire x_1509;
wire x_1510;
wire x_1511;
wire x_1512;
wire x_1513;
wire x_1514;
wire x_1515;
wire x_1516;
wire x_1517;
wire x_1518;
wire x_1519;
wire x_1520;
wire x_1521;
wire x_1522;
wire x_1523;
wire x_1524;
wire x_1525;
wire x_1526;
wire x_1527;
wire x_1528;
wire x_1529;
wire x_1530;
wire x_1531;
wire x_1532;
wire x_1533;
wire x_1534;
wire x_1535;
wire x_1536;
wire x_1537;
wire x_1538;
wire x_1539;
wire x_1540;
wire x_1541;
wire x_1542;
wire x_1543;
wire x_1544;
wire x_1545;
wire x_1546;
wire x_1547;
wire x_1548;
wire x_1549;
wire x_1550;
wire x_1551;
wire x_1552;
wire x_1553;
wire x_1554;
wire x_1555;
wire x_1556;
wire x_1557;
wire x_1558;
wire x_1559;
wire x_1560;
wire x_1561;
wire x_1562;
wire x_1563;
wire x_1564;
wire x_1565;
wire x_1566;
wire x_1567;
wire x_1568;
wire x_1569;
wire x_1570;
wire x_1571;
wire x_1572;
wire x_1573;
wire x_1574;
wire x_1575;
wire x_1576;
wire x_1577;
wire x_1578;
wire x_1579;
wire x_1580;
wire x_1581;
wire x_1582;
wire x_1583;
wire x_1584;
wire x_1585;
wire x_1586;
wire x_1587;
wire x_1588;
wire x_1589;
wire x_1590;
wire x_1591;
wire x_1592;
wire x_1593;
wire x_1594;
wire x_1595;
wire x_1596;
wire x_1597;
wire x_1598;
wire x_1599;
wire x_1600;
wire x_1601;
wire x_1602;
wire x_1603;
wire x_1604;
wire x_1605;
wire x_1606;
wire x_1607;
wire x_1608;
wire x_1609;
wire x_1610;
wire x_1611;
wire x_1612;
wire x_1613;
wire x_1614;
wire x_1615;
wire x_1616;
wire x_1617;
wire x_1618;
wire x_1619;
wire x_1620;
wire x_1621;
wire x_1622;
wire x_1623;
wire x_1624;
wire x_1625;
wire x_1626;
wire x_1627;
wire x_1628;
wire x_1629;
wire x_1630;
wire x_1631;
wire x_1632;
wire x_1633;
wire x_1634;
wire x_1635;
wire x_1636;
wire x_1637;
wire x_1638;
wire x_1639;
wire x_1640;
wire x_1641;
wire x_1642;
wire x_1643;
wire x_1644;
wire x_1645;
wire x_1646;
wire x_1647;
wire x_1648;
wire x_1649;
wire x_1650;
wire x_1651;
wire x_1652;
wire x_1653;
wire x_1654;
wire x_1655;
wire x_1656;
wire x_1657;
wire x_1658;
wire x_1659;
wire x_1660;
wire x_1661;
wire x_1662;
wire x_1663;
wire x_1664;
wire x_1665;
wire x_1666;
wire x_1667;
wire x_1668;
wire x_1669;
wire x_1670;
wire x_1671;
wire x_1672;
wire x_1673;
wire x_1674;
wire x_1675;
wire x_1676;
wire x_1677;
wire x_1678;
wire x_1679;
wire x_1680;
wire x_1681;
wire x_1682;
wire x_1683;
wire x_1684;
wire x_1685;
wire x_1686;
wire x_1687;
wire x_1688;
wire x_1689;
wire x_1690;
wire x_1691;
wire x_1692;
wire x_1693;
wire x_1694;
wire x_1695;
wire x_1696;
wire x_1697;
wire x_1698;
wire x_1699;
wire x_1700;
wire x_1701;
wire x_1702;
wire x_1703;
wire x_1704;
wire x_1705;
wire x_1706;
wire x_1707;
wire x_1708;
wire x_1709;
wire x_1710;
wire x_1711;
wire x_1712;
wire x_1713;
wire x_1714;
wire x_1715;
wire x_1716;
wire x_1717;
wire x_1718;
wire x_1719;
wire x_1720;
wire x_1721;
wire x_1722;
wire x_1723;
wire x_1724;
wire x_1725;
wire x_1726;
wire x_1727;
wire x_1728;
wire x_1729;
wire x_1730;
wire x_1731;
wire x_1732;
wire x_1733;
wire x_1734;
wire x_1735;
wire x_1736;
wire x_1737;
wire x_1738;
wire x_1739;
wire x_1740;
wire x_1741;
wire x_1742;
wire x_1743;
wire x_1744;
wire x_1745;
wire x_1746;
wire x_1747;
wire x_1748;
wire x_1749;
wire x_1750;
wire x_1751;
wire x_1752;
wire x_1753;
wire x_1754;
wire x_1755;
wire x_1756;
wire x_1757;
wire x_1758;
wire x_1759;
wire x_1760;
wire x_1761;
wire x_1762;
wire x_1763;
wire x_1764;
wire x_1765;
wire x_1766;
wire x_1767;
wire x_1768;
wire x_1769;
wire x_1770;
wire x_1771;
wire x_1772;
wire x_1773;
wire x_1774;
wire x_1775;
wire x_1776;
wire x_1777;
wire x_1778;
wire x_1779;
wire x_1780;
wire x_1781;
wire x_1782;
wire x_1783;
wire x_1784;
wire x_1785;
wire x_1786;
wire x_1787;
wire x_1788;
wire x_1789;
wire x_1790;
wire x_1791;
wire x_1792;
wire x_1793;
wire x_1794;
wire x_1795;
wire x_1796;
wire x_1797;
wire x_1798;
wire x_1799;
wire x_1800;
wire x_1801;
wire x_1802;
wire x_1803;
wire x_1804;
wire x_1805;
wire x_1806;
wire x_1807;
wire x_1808;
wire x_1809;
wire x_1810;
wire x_1811;
wire x_1812;
wire x_1813;
wire x_1814;
wire x_1815;
wire x_1816;
wire x_1817;
wire x_1818;
wire x_1819;
wire x_1820;
wire x_1821;
wire x_1822;
wire x_1823;
wire x_1824;
wire x_1825;
wire x_1826;
wire x_1827;
wire x_1828;
wire x_1829;
wire x_1830;
wire x_1831;
wire x_1832;
wire x_1833;
wire x_1834;
wire x_1835;
wire x_1836;
wire x_1837;
wire x_1838;
wire x_1839;
wire x_1840;
wire x_1841;
wire x_1842;
wire x_1843;
wire x_1844;
wire x_1845;
wire x_1846;
wire x_1847;
wire x_1848;
wire x_1849;
wire x_1850;
wire x_1851;
wire x_1852;
wire x_1853;
wire x_1854;
wire x_1855;
wire x_1856;
wire x_1857;
wire x_1858;
wire x_1859;
wire x_1860;
wire x_1861;
wire x_1862;
wire x_1863;
wire x_1864;
wire x_1865;
wire x_1866;
wire x_1867;
wire x_1868;
wire x_1869;
wire x_1870;
wire x_1871;
wire x_1872;
wire x_1873;
wire x_1874;
wire x_1875;
wire x_1876;
wire x_1877;
wire x_1878;
wire x_1879;
wire x_1880;
wire x_1881;
wire x_1882;
wire x_1883;
wire x_1884;
wire x_1885;
wire x_1886;
wire x_1887;
wire x_1888;
wire x_1889;
wire x_1890;
wire x_1891;
wire x_1892;
wire x_1893;
wire x_1894;
wire x_1895;
wire x_1896;
wire x_1897;
wire x_1898;
wire x_1899;
wire x_1900;
wire x_1901;
wire x_1902;
wire x_1903;
wire x_1904;
wire x_1905;
wire x_1906;
wire x_1907;
wire x_1908;
wire x_1909;
wire x_1910;
wire x_1911;
wire x_1912;
wire x_1913;
wire x_1914;
wire x_1915;
wire x_1916;
wire x_1917;
wire x_1918;
wire x_1919;
wire x_1920;
wire x_1921;
wire x_1922;
wire x_1923;
wire x_1924;
wire x_1925;
wire x_1926;
wire x_1927;
wire x_1928;
wire x_1929;
wire x_1930;
wire x_1931;
wire x_1932;
wire x_1933;
wire x_1934;
wire x_1935;
wire x_1936;
wire x_1937;
wire x_1938;
wire x_1939;
wire x_1940;
wire x_1941;
wire x_1942;
wire x_1943;
wire x_1944;
wire x_1945;
wire x_1946;
wire x_1947;
wire x_1948;
wire x_1949;
wire x_1950;
wire x_1951;
wire x_1952;
wire x_1953;
wire x_1954;
wire x_1955;
wire x_1956;
wire x_1957;
wire x_1958;
wire x_1959;
wire x_1960;
wire x_1961;
wire x_1962;
wire x_1963;
wire x_1964;
wire x_1965;
wire x_1966;
wire x_1967;
wire x_1968;
wire x_1969;
wire x_1970;
wire x_1971;
wire x_1972;
wire x_1973;
wire x_1974;
wire x_1975;
wire x_1976;
wire x_1977;
wire x_1978;
wire x_1979;
wire x_1980;
wire x_1981;
wire x_1982;
wire x_1983;
wire x_1984;
wire x_1985;
wire x_1986;
wire x_1987;
wire x_1988;
wire x_1989;
wire x_1990;
wire x_1991;
wire x_1992;
wire x_1993;
wire x_1994;
wire x_1995;
wire x_1996;
wire x_1997;
wire x_1998;
wire x_1999;
wire x_2000;
wire x_2001;
wire x_2002;
wire x_2003;
wire x_2004;
wire x_2005;
wire x_2006;
wire x_2007;
wire x_2008;
wire x_2009;
wire x_2010;
wire x_2011;
wire x_2012;
wire x_2013;
wire x_2014;
wire x_2015;
wire x_2016;
wire x_2017;
wire x_2018;
wire x_2019;
wire x_2020;
wire x_2021;
wire x_2022;
wire x_2023;
wire x_2024;
wire x_2025;
wire x_2026;
wire x_2027;
wire x_2028;
wire x_2029;
wire x_2030;
wire x_2031;
wire x_2032;
wire x_2033;
wire x_2034;
wire x_2035;
wire x_2036;
wire x_2037;
wire x_2038;
wire x_2039;
wire x_2040;
wire x_2041;
wire x_2042;
wire x_2043;
wire x_2044;
wire x_2045;
wire x_2046;
wire x_2047;
wire x_2048;
wire x_2049;
wire x_2050;
wire x_2051;
wire x_2052;
wire x_2053;
wire x_2054;
wire x_2055;
wire x_2056;
wire x_2057;
wire x_2058;
wire x_2059;
wire x_2060;
wire x_2061;
wire x_2062;
wire x_2063;
wire x_2064;
wire x_2065;
wire x_2066;
wire x_2067;
wire x_2068;
wire x_2069;
wire x_2070;
wire x_2071;
wire x_2072;
wire x_2073;
wire x_2074;
wire x_2075;
wire x_2076;
wire x_2077;
wire x_2078;
wire x_2079;
wire x_2080;
wire x_2081;
wire x_2082;
wire x_2083;
wire x_2084;
wire x_2085;
wire x_2086;
wire x_2087;
wire x_2088;
wire x_2089;
wire x_2090;
wire x_2091;
wire x_2092;
wire x_2093;
wire x_2094;
wire x_2095;
wire x_2096;
wire x_2097;
wire x_2098;
wire x_2099;
wire x_2100;
wire x_2101;
wire x_2102;
wire x_2103;
wire x_2104;
wire x_2105;
wire x_2106;
wire x_2107;
wire x_2108;
wire x_2109;
wire x_2110;
wire x_2111;
wire x_2112;
wire x_2113;
wire x_2114;
wire x_2115;
wire x_2116;
wire x_2117;
wire x_2118;
wire x_2119;
wire x_2120;
wire x_2121;
wire x_2122;
wire x_2123;
wire x_2124;
wire x_2125;
wire x_2126;
wire x_2127;
wire x_2128;
wire x_2129;
wire x_2130;
wire x_2131;
wire x_2132;
wire x_2133;
wire x_2134;
wire x_2135;
wire x_2136;
wire x_2137;
wire x_2138;
wire x_2139;
wire x_2140;
wire x_2141;
wire x_2142;
wire x_2143;
wire x_2144;
wire x_2145;
wire x_2146;
wire x_2147;
wire x_2148;
wire x_2149;
wire x_2150;
wire x_2151;
wire x_2152;
wire x_2153;
wire x_2154;
wire x_2155;
wire x_2156;
wire x_2157;
wire x_2158;
wire x_2159;
wire x_2160;
wire x_2161;
wire x_2162;
wire x_2163;
wire x_2164;
wire x_2165;
wire x_2166;
wire x_2167;
wire x_2168;
wire x_2169;
wire x_2170;
wire x_2171;
wire x_2172;
wire x_2173;
wire x_2174;
wire x_2175;
wire x_2176;
wire x_2177;
wire x_2178;
wire x_2179;
wire x_2180;
wire x_2181;
wire x_2182;
wire x_2183;
wire x_2184;
wire x_2185;
wire x_2186;
wire x_2187;
wire x_2188;
wire x_2189;
wire x_2190;
wire x_2191;
wire x_2192;
wire x_2193;
wire x_2194;
wire x_2195;
wire x_2196;
wire x_2197;
wire x_2198;
wire x_2199;
wire x_2200;
wire x_2201;
wire x_2202;
wire x_2203;
wire x_2204;
wire x_2205;
wire x_2206;
wire x_2207;
wire x_2208;
wire x_2209;
wire x_2210;
wire x_2211;
wire x_2212;
wire x_2213;
wire x_2214;
wire x_2215;
wire x_2216;
wire x_2217;
wire x_2218;
wire x_2219;
wire x_2220;
wire x_2221;
wire x_2222;
wire x_2223;
wire x_2224;
wire x_2225;
wire x_2226;
wire x_2227;
wire x_2228;
wire x_2229;
wire x_2230;
wire x_2231;
wire x_2232;
wire x_2233;
wire x_2234;
wire x_2235;
wire x_2236;
wire x_2237;
wire x_2238;
wire x_2239;
wire x_2240;
wire x_2241;
wire x_2242;
wire x_2243;
wire x_2244;
wire x_2245;
wire x_2246;
wire x_2247;
wire x_2248;
wire x_2249;
wire x_2250;
wire x_2251;
wire x_2252;
wire x_2253;
wire x_2254;
wire x_2255;
wire x_2256;
wire x_2257;
wire x_2258;
wire x_2259;
wire x_2260;
wire x_2261;
wire x_2262;
wire x_2263;
wire x_2264;
wire x_2265;
wire x_2266;
wire x_2267;
wire x_2268;
wire x_2269;
wire x_2270;
wire x_2271;
wire x_2272;
wire x_2273;
wire x_2274;
wire x_2275;
wire x_2276;
wire x_2277;
wire x_2278;
wire x_2279;
wire x_2280;
wire x_2281;
wire x_2282;
wire x_2283;
wire x_2284;
wire x_2285;
wire x_2286;
wire x_2287;
wire x_2288;
wire x_2289;
wire x_2290;
wire x_2291;
wire x_2292;
wire x_2293;
wire x_2294;
wire x_2295;
wire x_2296;
wire x_2297;
wire x_2298;
wire x_2299;
wire x_2300;
wire x_2301;
wire x_2302;
wire x_2303;
wire x_2304;
wire x_2305;
wire x_2306;
wire x_2307;
wire x_2308;
wire x_2309;
wire x_2310;
wire x_2311;
wire x_2312;
wire x_2313;
wire x_2314;
wire x_2315;
wire x_2316;
wire x_2317;
wire x_2318;
wire x_2319;
wire x_2320;
wire x_2321;
wire x_2322;
wire x_2323;
wire x_2324;
wire x_2325;
wire x_2326;
wire x_2327;
wire x_2328;
wire x_2329;
wire x_2330;
wire x_2331;
wire x_2332;
wire x_2333;
wire x_2334;
wire x_2335;
wire x_2336;
wire x_2337;
wire x_2338;
wire x_2339;
wire x_2340;
wire x_2341;
wire x_2342;
wire x_2343;
wire x_2344;
wire x_2345;
wire x_2346;
wire x_2347;
wire x_2348;
wire x_2349;
wire x_2350;
wire x_2351;
wire x_2352;
wire x_2353;
wire x_2354;
wire x_2355;
wire x_2356;
wire x_2357;
wire x_2358;
wire x_2359;
wire x_2360;
wire x_2361;
wire x_2362;
wire x_2363;
wire x_2364;
wire x_2365;
wire x_2366;
wire x_2367;
wire x_2368;
wire x_2369;
wire x_2370;
wire x_2371;
wire x_2372;
wire x_2373;
wire x_2374;
wire x_2375;
wire x_2376;
wire x_2377;
wire x_2378;
wire x_2379;
wire x_2380;
wire x_2381;
wire x_2382;
wire x_2383;
wire x_2384;
wire x_2385;
wire x_2386;
wire x_2387;
wire x_2388;
wire x_2389;
wire x_2390;
wire x_2391;
wire x_2392;
wire x_2393;
wire x_2394;
wire x_2395;
wire x_2396;
wire x_2397;
wire x_2398;
wire x_2399;
wire x_2400;
wire x_2401;
wire x_2402;
wire x_2403;
wire x_2404;
wire x_2405;
wire x_2406;
wire x_2407;
wire x_2408;
wire x_2409;
wire x_2410;
wire x_2411;
wire x_2412;
wire x_2413;
wire x_2414;
wire x_2415;
wire x_2416;
wire x_2417;
wire x_2418;
wire x_2419;
wire x_2420;
wire x_2421;
wire x_2422;
wire x_2423;
wire x_2424;
wire x_2425;
wire x_2426;
wire x_2427;
wire x_2428;
wire x_2429;
wire x_2430;
wire x_2431;
wire x_2432;
wire x_2433;
wire x_2434;
wire x_2435;
wire x_2436;
wire x_2437;
wire x_2438;
wire x_2439;
wire x_2440;
wire x_2441;
wire x_2442;
wire x_2443;
wire x_2444;
wire x_2445;
wire x_2446;
wire x_2447;
wire x_2448;
wire x_2449;
wire x_2450;
wire x_2451;
wire x_2452;
wire x_2453;
wire x_2454;
wire x_2455;
wire x_2456;
wire x_2457;
wire x_2458;
wire x_2459;
wire x_2460;
wire x_2461;
wire x_2462;
wire x_2463;
wire x_2464;
wire x_2465;
wire x_2466;
wire x_2467;
wire x_2468;
wire x_2469;
wire x_2470;
wire x_2471;
wire x_2472;
wire x_2473;
wire x_2474;
wire x_2475;
wire x_2476;
wire x_2477;
wire x_2478;
wire x_2479;
wire x_2480;
wire x_2481;
wire x_2482;
wire x_2483;
wire x_2484;
wire x_2485;
wire x_2486;
wire x_2487;
wire x_2488;
wire x_2489;
wire x_2490;
wire x_2491;
wire x_2492;
wire x_2493;
wire x_2494;
wire x_2495;
wire x_2496;
wire x_2497;
wire x_2498;
wire x_2499;
wire x_2500;
wire x_2501;
wire x_2502;
wire x_2503;
wire x_2504;
wire x_2505;
wire x_2506;
wire x_2507;
wire x_2508;
wire x_2509;
wire x_2510;
wire x_2511;
wire x_2512;
wire x_2513;
wire x_2514;
wire x_2515;
wire x_2516;
wire x_2517;
wire x_2518;
wire x_2519;
wire x_2520;
wire x_2521;
wire x_2522;
wire x_2523;
wire x_2524;
wire x_2525;
wire x_2526;
wire x_2527;
wire x_2528;
wire x_2529;
wire x_2530;
wire x_2531;
wire x_2532;
wire x_2533;
wire x_2534;
wire x_2535;
wire x_2536;
wire x_2537;
wire x_2538;
wire x_2539;
wire x_2540;
wire x_2541;
wire x_2542;
wire x_2543;
wire x_2544;
wire x_2545;
wire x_2546;
wire x_2547;
wire x_2548;
wire x_2549;
wire x_2550;
wire x_2551;
wire x_2552;
wire x_2553;
wire x_2554;
wire x_2555;
wire x_2556;
wire x_2557;
wire x_2558;
wire x_2559;
wire x_2560;
wire x_2561;
wire x_2562;
wire x_2563;
wire x_2564;
wire x_2565;
wire x_2566;
wire x_2567;
wire x_2568;
wire x_2569;
wire x_2570;
wire x_2571;
wire x_2572;
wire x_2573;
wire x_2574;
wire x_2575;
wire x_2576;
wire x_2577;
wire x_2578;
wire x_2579;
wire x_2580;
wire x_2581;
wire x_2582;
wire x_2583;
wire x_2584;
wire x_2585;
wire x_2586;
wire x_2587;
wire x_2588;
wire x_2589;
wire x_2590;
wire x_2591;
wire x_2592;
wire x_2593;
wire x_2594;
wire x_2595;
wire x_2596;
wire x_2597;
wire x_2598;
wire x_2599;
wire x_2600;
wire x_2601;
wire x_2602;
wire x_2603;
wire x_2604;
wire x_2605;
wire x_2606;
wire x_2607;
wire x_2608;
wire x_2609;
wire x_2610;
wire x_2611;
wire x_2612;
wire x_2613;
wire x_2614;
wire x_2615;
wire x_2616;
wire x_2617;
wire x_2618;
wire x_2619;
wire x_2620;
wire x_2621;
wire x_2622;
wire x_2623;
wire x_2624;
wire x_2625;
wire x_2626;
wire x_2627;
wire x_2628;
wire x_2629;
wire x_2630;
wire x_2631;
wire x_2632;
wire x_2633;
wire x_2634;
wire x_2635;
wire x_2636;
wire x_2637;
wire x_2638;
wire x_2639;
wire x_2640;
wire x_2641;
wire x_2642;
wire x_2643;
wire x_2644;
wire x_2645;
wire x_2646;
wire x_2647;
wire x_2648;
wire x_2649;
wire x_2650;
wire x_2651;
wire x_2652;
wire x_2653;
wire x_2654;
wire x_2655;
wire x_2656;
wire x_2657;
wire x_2658;
wire x_2659;
wire x_2660;
wire x_2661;
wire x_2662;
wire x_2663;
wire x_2664;
wire x_2665;
wire x_2666;
wire x_2667;
wire x_2668;
wire x_2669;
wire x_2670;
wire x_2671;
wire x_2672;
wire x_2673;
wire x_2674;
wire x_2675;
wire x_2676;
wire x_2677;
wire x_2678;
wire x_2679;
wire x_2680;
wire x_2681;
wire x_2682;
wire x_2683;
wire x_2684;
wire x_2685;
wire x_2686;
wire x_2687;
wire x_2688;
wire x_2689;
wire x_2690;
wire x_2691;
wire x_2692;
wire x_2693;
wire x_2694;
wire x_2695;
wire x_2696;
wire x_2697;
wire x_2698;
wire x_2699;
wire x_2700;
wire x_2701;
wire x_2702;
wire x_2703;
wire x_2704;
wire x_2705;
wire x_2706;
wire x_2707;
wire x_2708;
wire x_2709;
wire x_2710;
wire x_2711;
wire x_2712;
wire x_2713;
wire x_2714;
wire x_2715;
wire x_2716;
wire x_2717;
wire x_2718;
wire x_2719;
wire x_2720;
wire x_2721;
wire x_2722;
wire x_2723;
wire x_2724;
wire x_2725;
wire x_2726;
wire x_2727;
wire x_2728;
wire x_2729;
wire x_2730;
wire x_2731;
wire x_2732;
wire x_2733;
wire x_2734;
wire x_2735;
wire x_2736;
wire x_2737;
wire x_2738;
wire x_2739;
wire x_2740;
wire x_2741;
wire x_2742;
wire x_2743;
wire x_2744;
wire x_2745;
wire x_2746;
wire x_2747;
wire x_2748;
wire x_2749;
wire x_2750;
wire x_2751;
wire x_2752;
wire x_2753;
wire x_2754;
wire x_2755;
wire x_2756;
wire x_2757;
wire x_2758;
wire x_2759;
wire x_2760;
wire x_2761;
wire x_2762;
wire x_2763;
wire x_2764;
wire x_2765;
wire x_2766;
wire x_2767;
wire x_2768;
wire x_2769;
wire x_2770;
wire x_2771;
wire x_2772;
wire x_2773;
wire x_2774;
wire x_2775;
wire x_2776;
wire x_2777;
wire x_2778;
wire x_2779;
wire x_2780;
wire x_2781;
wire x_2782;
wire x_2783;
wire x_2784;
wire x_2785;
wire x_2786;
wire x_2787;
wire x_2788;
wire x_2789;
wire x_2790;
wire x_2791;
wire x_2792;
wire x_2793;
wire x_2794;
wire x_2795;
wire x_2796;
wire x_2797;
wire x_2798;
wire x_2799;
wire x_2800;
wire x_2801;
wire x_2802;
wire x_2803;
wire x_2804;
wire x_2805;
wire x_2806;
wire x_2807;
wire x_2808;
wire x_2809;
wire x_2810;
wire x_2811;
wire x_2812;
wire x_2813;
wire x_2814;
wire x_2815;
wire x_2816;
wire x_2817;
wire x_2818;
wire x_2819;
wire x_2820;
wire x_2821;
wire x_2822;
wire x_2823;
wire x_2824;
wire x_2825;
wire x_2826;
wire x_2827;
wire x_2828;
wire x_2829;
wire x_2830;
wire x_2831;
wire x_2832;
wire x_2833;
wire x_2834;
wire x_2835;
wire x_2836;
wire x_2837;
wire x_2838;
wire x_2839;
wire x_2840;
wire x_2841;
wire x_2842;
wire x_2843;
wire x_2844;
wire x_2845;
wire x_2846;
wire x_2847;
wire x_2848;
wire x_2849;
wire x_2850;
wire x_2851;
wire x_2852;
wire x_2853;
wire x_2854;
wire x_2855;
wire x_2856;
wire x_2857;
wire x_2858;
wire x_2859;
wire x_2860;
wire x_2861;
wire x_2862;
wire x_2863;
wire x_2864;
wire x_2865;
wire x_2866;
wire x_2867;
wire x_2868;
wire x_2869;
wire x_2870;
wire x_2871;
wire x_2872;
wire x_2873;
wire x_2874;
wire x_2875;
wire x_2876;
wire x_2877;
wire x_2878;
wire x_2879;
wire x_2880;
wire x_2881;
wire x_2882;
wire x_2883;
wire x_2884;
wire x_2885;
wire x_2886;
wire x_2887;
wire x_2888;
wire x_2889;
wire x_2890;
wire x_2891;
wire x_2892;
wire x_2893;
wire x_2894;
wire x_2895;
wire x_2896;
wire x_2897;
wire x_2898;
wire x_2899;
wire x_2900;
wire x_2901;
wire x_2902;
wire x_2903;
wire x_2904;
wire x_2905;
wire x_2906;
wire x_2907;
wire x_2908;
wire x_2909;
wire x_2910;
wire x_2911;
wire x_2912;
wire x_2913;
wire x_2914;
wire x_2915;
wire x_2916;
wire x_2917;
wire x_2918;
wire x_2919;
wire x_2920;
wire x_2921;
wire x_2922;
wire x_2923;
wire x_2924;
wire x_2925;
wire x_2926;
wire x_2927;
wire x_2928;
wire x_2929;
wire x_2930;
wire x_2931;
wire x_2932;
wire x_2933;
wire x_2934;
wire x_2935;
wire x_2936;
wire x_2937;
wire x_2938;
wire x_2939;
wire x_2940;
wire x_2941;
wire x_2942;
wire x_2943;
wire x_2944;
wire x_2945;
wire x_2946;
wire x_2947;
wire x_2948;
wire x_2949;
wire x_2950;
wire x_2951;
wire x_2952;
wire x_2953;
wire x_2954;
wire x_2955;
wire x_2956;
wire x_2957;
wire x_2958;
wire x_2959;
wire x_2960;
wire x_2961;
wire x_2962;
wire x_2963;
wire x_2964;
wire x_2965;
wire x_2966;
wire x_2967;
wire x_2968;
wire x_2969;
wire x_2970;
wire x_2971;
wire x_2972;
wire x_2973;
wire x_2974;
wire x_2975;
wire x_2976;
wire x_2977;
wire x_2978;
wire x_2979;
wire x_2980;
wire x_2981;
wire x_2982;
wire x_2983;
wire x_2984;
wire x_2985;
wire x_2986;
wire x_2987;
wire x_2988;
wire x_2989;
wire x_2990;
wire x_2991;
wire x_2992;
wire x_2993;
wire x_2994;
wire x_2995;
wire x_2996;
wire x_2997;
wire x_2998;
wire x_2999;
wire x_3000;
wire x_3001;
wire x_3002;
wire x_3003;
wire x_3004;
wire x_3005;
wire x_3006;
wire x_3007;
wire x_3008;
wire x_3009;
wire x_3010;
wire x_3011;
wire x_3012;
wire x_3013;
wire x_3014;
wire x_3015;
wire x_3016;
wire x_3017;
wire x_3018;
wire x_3019;
wire x_3020;
wire x_3021;
wire x_3022;
wire x_3023;
wire x_3024;
wire x_3025;
wire x_3026;
wire x_3027;
wire x_3028;
wire x_3029;
wire x_3030;
wire x_3031;
wire x_3032;
wire x_3033;
wire x_3034;
wire x_3035;
wire x_3036;
wire x_3037;
wire x_3038;
wire x_3039;
wire x_3040;
wire x_3041;
wire x_3042;
wire x_3043;
wire x_3044;
wire x_3045;
wire x_3046;
wire x_3047;
wire x_3048;
wire x_3049;
wire x_3050;
wire x_3051;
wire x_3052;
wire x_3053;
wire x_3054;
wire x_3055;
wire x_3056;
wire x_3057;
wire x_3058;
wire x_3059;
wire x_3060;
wire x_3061;
wire x_3062;
wire x_3063;
wire x_3064;
wire x_3065;
wire x_3066;
wire x_3067;
wire x_3068;
wire x_3069;
wire x_3070;
wire x_3071;
wire x_3072;
wire x_3073;
wire x_3074;
wire x_3075;
wire x_3076;
wire x_3077;
wire x_3078;
wire x_3079;
wire x_3080;
wire x_3081;
wire x_3082;
wire x_3083;
wire x_3084;
wire x_3085;
wire x_3086;
wire x_3087;
wire x_3088;
wire x_3089;
wire x_3090;
wire x_3091;
wire x_3092;
wire x_3093;
wire x_3094;
wire x_3095;
wire x_3096;
wire x_3097;
wire x_3098;
wire x_3099;
wire x_3100;
wire x_3101;
wire x_3102;
wire x_3103;
wire x_3104;
wire x_3105;
wire x_3106;
wire x_3107;
wire x_3108;
wire x_3109;
wire x_3110;
wire x_3111;
wire x_3112;
wire x_3113;
wire x_3114;
wire x_3115;
wire x_3116;
wire x_3117;
wire x_3118;
wire x_3119;
wire x_3120;
wire x_3121;
wire x_3122;
wire x_3123;
wire x_3124;
wire x_3125;
wire x_3126;
wire x_3127;
wire x_3128;
wire x_3129;
wire x_3130;
wire x_3131;
wire x_3132;
wire x_3133;
wire x_3134;
wire x_3135;
wire x_3136;
wire x_3137;
wire x_3138;
wire x_3139;
wire x_3140;
wire x_3141;
wire x_3142;
wire x_3143;
wire x_3144;
wire x_3145;
wire x_3146;
wire x_3147;
wire x_3148;
wire x_3149;
wire x_3150;
wire x_3151;
wire x_3152;
wire x_3153;
wire x_3154;
wire x_3155;
wire x_3156;
wire x_3157;
wire x_3158;
wire x_3159;
wire x_3160;
wire x_3161;
wire x_3162;
wire x_3163;
wire x_3164;
wire x_3165;
wire x_3166;
wire x_3167;
wire x_3168;
wire x_3169;
wire x_3170;
wire x_3171;
wire x_3172;
wire x_3173;
wire x_3174;
wire x_3175;
wire x_3176;
wire x_3177;
wire x_3178;
wire x_3179;
wire x_3180;
wire x_3181;
wire x_3182;
wire x_3183;
wire x_3184;
wire x_3185;
wire x_3186;
wire x_3187;
wire x_3188;
wire x_3189;
wire x_3190;
wire x_3191;
wire x_3192;
wire x_3193;
wire x_3194;
wire x_3195;
wire x_3196;
wire x_3197;
wire x_3198;
wire x_3199;
wire x_3200;
wire x_3201;
wire x_3202;
wire x_3203;
wire x_3204;
wire x_3205;
wire x_3206;
wire x_3207;
wire x_3208;
wire x_3209;
wire x_3210;
wire x_3211;
wire x_3212;
wire x_3213;
wire x_3214;
wire x_3215;
wire x_3216;
wire x_3217;
wire x_3218;
wire x_3219;
wire x_3220;
wire x_3221;
wire x_3222;
wire x_3223;
wire x_3224;
wire x_3225;
wire x_3226;
wire x_3227;
wire x_3228;
wire x_3229;
wire x_3230;
wire x_3231;
wire x_3232;
wire x_3233;
wire x_3234;
wire x_3235;
wire x_3236;
wire x_3237;
wire x_3238;
wire x_3239;
wire x_3240;
wire x_3241;
wire x_3242;
wire x_3243;
wire x_3244;
wire x_3245;
wire x_3246;
wire x_3247;
wire x_3248;
wire x_3249;
wire x_3250;
wire x_3251;
wire x_3252;
wire x_3253;
wire x_3254;
wire x_3255;
wire x_3256;
wire x_3257;
wire x_3258;
wire x_3259;
wire x_3260;
wire x_3261;
wire x_3262;
wire x_3263;
wire x_3264;
wire x_3265;
wire x_3266;
wire x_3267;
wire x_3268;
wire x_3269;
wire x_3270;
wire x_3271;
wire x_3272;
wire x_3273;
wire x_3274;
wire x_3275;
wire x_3276;
wire x_3277;
wire x_3278;
wire x_3279;
wire x_3280;
wire x_3281;
wire x_3282;
wire x_3283;
wire x_3284;
wire x_3285;
wire x_3286;
wire x_3287;
wire x_3288;
wire x_3289;
wire x_3290;
wire x_3291;
wire x_3292;
wire x_3293;
wire x_3294;
wire x_3295;
wire x_3296;
wire x_3297;
wire x_3298;
wire x_3299;
wire x_3300;
wire x_3301;
wire x_3302;
wire x_3303;
wire x_3304;
wire x_3305;
wire x_3306;
wire x_3307;
wire x_3308;
wire x_3309;
wire x_3310;
wire x_3311;
wire x_3312;
wire x_3313;
wire x_3314;
wire x_3315;
wire x_3316;
wire x_3317;
wire x_3318;
wire x_3319;
wire x_3320;
wire x_3321;
wire x_3322;
wire x_3323;
wire x_3324;
wire x_3325;
wire x_3326;
wire x_3327;
wire x_3328;
wire x_3329;
wire x_3330;
wire x_3331;
wire x_3332;
wire x_3333;
wire x_3334;
wire x_3335;
wire x_3336;
wire x_3337;
wire x_3338;
wire x_3339;
wire x_3340;
wire x_3341;
wire x_3342;
wire x_3343;
wire x_3344;
wire x_3345;
wire x_3346;
wire x_3347;
wire x_3348;
wire x_3349;
wire x_3350;
wire x_3351;
wire x_3352;
wire x_3353;
wire x_3354;
wire x_3355;
wire x_3356;
wire x_3357;
wire x_3358;
wire x_3359;
wire x_3360;
wire x_3361;
wire x_3362;
wire x_3363;
wire x_3364;
wire x_3365;
wire x_3366;
wire x_3367;
wire x_3368;
wire x_3369;
wire x_3370;
wire x_3371;
wire x_3372;
wire x_3373;
wire x_3374;
wire x_3375;
wire x_3376;
wire x_3377;
wire x_3378;
wire x_3379;
wire x_3380;
wire x_3381;
wire x_3382;
wire x_3383;
wire x_3384;
wire x_3385;
wire x_3386;
wire x_3387;
wire x_3388;
wire x_3389;
wire x_3390;
wire x_3391;
wire x_3392;
wire x_3393;
wire x_3394;
wire x_3395;
wire x_3396;
wire x_3397;
wire x_3398;
wire x_3399;
wire x_3400;
wire x_3401;
wire x_3402;
wire x_3403;
wire x_3404;
wire x_3405;
wire x_3406;
wire x_3407;
wire x_3408;
wire x_3409;
wire x_3410;
wire x_3411;
wire x_3412;
wire x_3413;
wire x_3414;
wire x_3415;
wire x_3416;
wire x_3417;
wire x_3418;
wire x_3419;
wire x_3420;
wire x_3421;
wire x_3422;
wire x_3423;
wire x_3424;
wire x_3425;
wire x_3426;
wire x_3427;
wire x_3428;
wire x_3429;
wire x_3430;
wire x_3431;
wire x_3432;
wire x_3433;
wire x_3434;
wire x_3435;
wire x_3436;
wire x_3437;
wire x_3438;
wire x_3439;
wire x_3440;
wire x_3441;
wire x_3442;
wire x_3443;
wire x_3444;
wire x_3445;
wire x_3446;
wire x_3447;
wire x_3448;
wire x_3449;
wire x_3450;
wire x_3451;
wire x_3452;
wire x_3453;
wire x_3454;
wire x_3455;
wire x_3456;
wire x_3457;
wire x_3458;
wire x_3459;
wire x_3460;
wire x_3461;
wire x_3462;
wire x_3463;
wire x_3464;
wire x_3465;
wire x_3466;
wire x_3467;
wire x_3468;
wire x_3469;
wire x_3470;
wire x_3471;
wire x_3472;
wire x_3473;
wire x_3474;
wire x_3475;
wire x_3476;
wire x_3477;
wire x_3478;
wire x_3479;
wire x_3480;
wire x_3481;
wire x_3482;
wire x_3483;
wire x_3484;
wire x_3485;
wire x_3486;
wire x_3487;
wire x_3488;
wire x_3489;
wire x_3490;
wire x_3491;
wire x_3492;
wire x_3493;
wire x_3494;
wire x_3495;
wire x_3496;
wire x_3497;
wire x_3498;
wire x_3499;
wire x_3500;
wire x_3501;
wire x_3502;
wire x_3503;
wire x_3504;
wire x_3505;
wire x_3506;
wire x_3507;
wire x_3508;
wire x_3509;
wire x_3510;
wire x_3511;
wire x_3512;
wire x_3513;
wire x_3514;
wire x_3515;
wire x_3516;
wire x_3517;
wire x_3518;
wire x_3519;
wire x_3520;
wire x_3521;
wire x_3522;
wire x_3523;
wire x_3524;
wire x_3525;
wire x_3526;
wire x_3527;
wire x_3528;
wire x_3529;
wire x_3530;
wire x_3531;
wire x_3532;
wire x_3533;
wire x_3534;
wire x_3535;
wire x_3536;
wire x_3537;
wire x_3538;
wire x_3539;
wire x_3540;
wire x_3541;
wire x_3542;
wire x_3543;
wire x_3544;
wire x_3545;
wire x_3546;
wire x_3547;
wire x_3548;
wire x_3549;
wire x_3550;
wire x_3551;
wire x_3552;
wire x_3553;
wire x_3554;
wire x_3555;
wire x_3556;
wire x_3557;
wire x_3558;
wire x_3559;
wire x_3560;
wire x_3561;
wire x_3562;
wire x_3563;
wire x_3564;
wire x_3565;
wire x_3566;
wire x_3567;
wire x_3568;
wire x_3569;
wire x_3570;
wire x_3571;
wire x_3572;
wire x_3573;
wire x_3574;
wire x_3575;
wire x_3576;
wire x_3577;
wire x_3578;
wire x_3579;
wire x_3580;
wire x_3581;
wire x_3582;
wire x_3583;
wire x_3584;
wire x_3585;
wire x_3586;
wire x_3587;
wire x_3588;
wire x_3589;
wire x_3590;
wire x_3591;
wire x_3592;
wire x_3593;
wire x_3594;
wire x_3595;
wire x_3596;
wire x_3597;
wire x_3598;
wire x_3599;
wire x_3600;
wire x_3601;
wire x_3602;
wire x_3603;
wire x_3604;
wire x_3605;
wire x_3606;
wire x_3607;
wire x_3608;
wire x_3609;
wire x_3610;
wire x_3611;
wire x_3612;
wire x_3613;
wire x_3614;
wire x_3615;
wire x_3616;
wire x_3617;
wire x_3618;
wire x_3619;
wire x_3620;
wire x_3621;
wire x_3622;
wire x_3623;
wire x_3624;
wire x_3625;
wire x_3626;
wire x_3627;
wire x_3628;
wire x_3629;
wire x_3630;
wire x_3631;
wire x_3632;
wire x_3633;
wire x_3634;
wire x_3635;
wire x_3636;
wire x_3637;
wire x_3638;
wire x_3639;
wire x_3640;
wire x_3641;
wire x_3642;
wire x_3643;
wire x_3644;
wire x_3645;
wire x_3646;
wire x_3647;
wire x_3648;
wire x_3649;
wire x_3650;
wire x_3651;
wire x_3652;
wire x_3653;
wire x_3654;
wire x_3655;
wire x_3656;
wire x_3657;
wire x_3658;
wire x_3659;
wire x_3660;
wire x_3661;
wire x_3662;
wire x_3663;
wire x_3664;
wire x_3665;
wire x_3666;
wire x_3667;
wire x_3668;
wire x_3669;
wire x_3670;
wire x_3671;
wire x_3672;
wire x_3673;
wire x_3674;
wire x_3675;
wire x_3676;
wire x_3677;
wire x_3678;
wire x_3679;
wire x_3680;
wire x_3681;
wire x_3682;
wire x_3683;
wire x_3684;
wire x_3685;
wire x_3686;
wire x_3687;
wire x_3688;
wire x_3689;
wire x_3690;
wire x_3691;
wire x_3692;
wire x_3693;
wire x_3694;
wire x_3695;
wire x_3696;
wire x_3697;
wire x_3698;
wire x_3699;
wire x_3700;
wire x_3701;
wire x_3702;
wire x_3703;
wire x_3704;
wire x_3705;
wire x_3706;
wire x_3707;
wire x_3708;
wire x_3709;
wire x_3710;
wire x_3711;
wire x_3712;
wire x_3713;
wire x_3714;
wire x_3715;
wire x_3716;
wire x_3717;
wire x_3718;
wire x_3719;
wire x_3720;
wire x_3721;
wire x_3722;
wire x_3723;
wire x_3724;
wire x_3725;
wire x_3726;
wire x_3727;
wire x_3728;
wire x_3729;
wire x_3730;
wire x_3731;
wire x_3732;
wire x_3733;
wire x_3734;
wire x_3735;
wire x_3736;
wire x_3737;
wire x_3738;
wire x_3739;
wire x_3740;
wire x_3741;
wire x_3742;
wire x_3743;
wire x_3744;
wire x_3745;
wire x_3746;
wire x_3747;
wire x_3748;
wire x_3749;
wire x_3750;
wire x_3751;
wire x_3752;
wire x_3753;
wire x_3754;
wire x_3755;
wire x_3756;
wire x_3757;
wire x_3758;
wire x_3759;
wire x_3760;
wire x_3761;
wire x_3762;
wire x_3763;
wire x_3764;
wire x_3765;
wire x_3766;
wire x_3767;
wire x_3768;
wire x_3769;
wire x_3770;
wire x_3771;
wire x_3772;
wire x_3773;
wire x_3774;
wire x_3775;
wire x_3776;
wire x_3777;
wire x_3778;
wire x_3779;
wire x_3780;
wire x_3781;
wire x_3782;
wire x_3783;
wire x_3784;
wire x_3785;
wire x_3786;
wire x_3787;
wire x_3788;
wire x_3789;
wire x_3790;
wire x_3791;
wire x_3792;
wire x_3793;
wire x_3794;
wire x_3795;
wire x_3796;
wire x_3797;
wire x_3798;
wire x_3799;
wire x_3800;
wire x_3801;
wire x_3802;
wire x_3803;
wire x_3804;
wire x_3805;
wire x_3806;
wire x_3807;
wire x_3808;
wire x_3809;
wire x_3810;
wire x_3811;
wire x_3812;
wire x_3813;
wire x_3814;
wire x_3815;
wire x_3816;
wire x_3817;
wire x_3818;
wire x_3819;
wire x_3820;
wire x_3821;
wire x_3822;
wire x_3823;
wire x_3824;
wire x_3825;
wire x_3826;
wire x_3827;
wire x_3828;
wire x_3829;
wire x_3830;
wire x_3831;
wire x_3832;
wire x_3833;
wire x_3834;
wire x_3835;
wire x_3836;
wire x_3837;
wire x_3838;
wire x_3839;
wire x_3840;
wire x_3841;
wire x_3842;
wire x_3843;
wire x_3844;
wire x_3845;
wire x_3846;
wire x_3847;
wire x_3848;
wire x_3849;
wire x_3850;
wire x_3851;
wire x_3852;
wire x_3853;
wire x_3854;
wire x_3855;
wire x_3856;
wire x_3857;
wire x_3858;
wire x_3859;
wire x_3860;
wire x_3861;
wire x_3862;
wire x_3863;
wire x_3864;
wire x_3865;
wire x_3866;
wire x_3867;
wire x_3868;
wire x_3869;
wire x_3870;
wire x_3871;
wire x_3872;
wire x_3873;
wire x_3874;
wire x_3875;
wire x_3876;
wire x_3877;
wire x_3878;
wire x_3879;
wire x_3880;
wire x_3881;
wire x_3882;
wire x_3883;
wire x_3884;
wire x_3885;
wire x_3886;
wire x_3887;
wire x_3888;
wire x_3889;
wire x_3890;
wire x_3891;
wire x_3892;
wire x_3893;
wire x_3894;
wire x_3895;
wire x_3896;
wire x_3897;
wire x_3898;
wire x_3899;
wire x_3900;
wire x_3901;
wire x_3902;
wire x_3903;
wire x_3904;
wire x_3905;
wire x_3906;
wire x_3907;
wire x_3908;
wire x_3909;
wire x_3910;
wire x_3911;
wire x_3912;
wire x_3913;
wire x_3914;
wire x_3915;
wire x_3916;
wire x_3917;
wire x_3918;
wire x_3919;
wire x_3920;
wire x_3921;
wire x_3922;
wire x_3923;
wire x_3924;
wire x_3925;
wire x_3926;
wire x_3927;
wire x_3928;
wire x_3929;
wire x_3930;
wire x_3931;
wire x_3932;
wire x_3933;
wire x_3934;
wire x_3935;
wire x_3936;
wire x_3937;
wire x_3938;
wire x_3939;
wire x_3940;
wire x_3941;
wire x_3942;
wire x_3943;
wire x_3944;
wire x_3945;
wire x_3946;
wire x_3947;
wire x_3948;
wire x_3949;
wire x_3950;
wire x_3951;
wire x_3952;
wire x_3953;
wire x_3954;
wire x_3955;
wire x_3956;
wire x_3957;
wire x_3958;
wire x_3959;
wire x_3960;
wire x_3961;
wire x_3962;
wire x_3963;
wire x_3964;
wire x_3965;
wire x_3966;
wire x_3967;
wire x_3968;
wire x_3969;
wire x_3970;
wire x_3971;
wire x_3972;
wire x_3973;
wire x_3974;
wire x_3975;
wire x_3976;
wire x_3977;
wire x_3978;
wire x_3979;
wire x_3980;
wire x_3981;
wire x_3982;
wire x_3983;
wire x_3984;
wire x_3985;
wire x_3986;
wire x_3987;
wire x_3988;
wire x_3989;
wire x_3990;
wire x_3991;
wire x_3992;
wire x_3993;
wire x_3994;
wire x_3995;
wire x_3996;
wire x_3997;
wire x_3998;
wire x_3999;
wire x_4000;
wire x_4001;
wire x_4002;
wire x_4003;
wire x_4004;
wire x_4005;
wire x_4006;
wire x_4007;
wire x_4008;
wire x_4009;
wire x_4010;
wire x_4011;
wire x_4012;
wire x_4013;
wire x_4014;
wire x_4015;
wire x_4016;
wire x_4017;
wire x_4018;
wire x_4019;
wire x_4020;
wire x_4021;
wire x_4022;
wire x_4023;
wire x_4024;
wire x_4025;
wire x_4026;
wire x_4027;
wire x_4028;
wire x_4029;
wire x_4030;
wire x_4031;
wire x_4032;
wire x_4033;
wire x_4034;
wire x_4035;
wire x_4036;
wire x_4037;
wire x_4038;
wire x_4039;
wire x_4040;
wire x_4041;
wire x_4042;
wire x_4043;
wire x_4044;
wire x_4045;
wire x_4046;
wire x_4047;
wire x_4048;
wire x_4049;
wire x_4050;
wire x_4051;
wire x_4052;
wire x_4053;
wire x_4054;
wire x_4055;
wire x_4056;
wire x_4057;
wire x_4058;
wire x_4059;
wire x_4060;
wire x_4061;
wire x_4062;
wire x_4063;
wire x_4064;
wire x_4065;
wire x_4066;
wire x_4067;
wire x_4068;
wire x_4069;
wire x_4070;
wire x_4071;
wire x_4072;
wire x_4073;
wire x_4074;
wire x_4075;
wire x_4076;
wire x_4077;
wire x_4078;
wire x_4079;
wire x_4080;
wire x_4081;
wire x_4082;
wire x_4083;
wire x_4084;
wire x_4085;
wire x_4086;
wire x_4087;
wire x_4088;
wire x_4089;
wire x_4090;
wire x_4091;
wire x_4092;
wire x_4093;
wire x_4094;
wire x_4095;
wire x_4096;
wire x_4097;
wire x_4098;
wire x_4099;
wire x_4100;
wire x_4101;
wire x_4102;
wire x_4103;
wire x_4104;
wire x_4105;
wire x_4106;
wire x_4107;
wire x_4108;
wire x_4109;
wire x_4110;
wire x_4111;
wire x_4112;
wire x_4113;
wire x_4114;
wire x_4115;
wire x_4116;
wire x_4117;
wire x_4118;
wire x_4119;
wire x_4120;
wire x_4121;
wire x_4122;
wire x_4123;
wire x_4124;
wire x_4125;
wire x_4126;
wire x_4127;
wire x_4128;
wire x_4129;
wire x_4130;
wire x_4131;
wire x_4132;
wire x_4133;
wire x_4134;
wire x_4135;
wire x_4136;
wire x_4137;
wire x_4138;
wire x_4139;
wire x_4140;
wire x_4141;
wire x_4142;
wire x_4143;
wire x_4144;
wire x_4145;
wire x_4146;
wire x_4147;
wire x_4148;
wire x_4149;
wire x_4150;
wire x_4151;
wire x_4152;
wire x_4153;
wire x_4154;
wire x_4155;
wire x_4156;
wire x_4157;
wire x_4158;
wire x_4159;
wire x_4160;
wire x_4161;
wire x_4162;
wire x_4163;
wire x_4164;
wire x_4165;
wire x_4166;
wire x_4167;
wire x_4168;
wire x_4169;
wire x_4170;
wire x_4171;
wire x_4172;
wire x_4173;
wire x_4174;
wire x_4175;
wire x_4176;
wire x_4177;
wire x_4178;
wire x_4179;
wire x_4180;
wire x_4181;
wire x_4182;
wire x_4183;
wire x_4184;
wire x_4185;
wire x_4186;
wire x_4187;
wire x_4188;
wire x_4189;
wire x_4190;
wire x_4191;
wire x_4192;
wire x_4193;
wire x_4194;
wire x_4195;
wire x_4196;
wire x_4197;
wire x_4198;
wire x_4199;
wire x_4200;
wire x_4201;
wire x_4202;
wire x_4203;
wire x_4204;
wire x_4205;
wire x_4206;
wire x_4207;
wire x_4208;
wire x_4209;
wire x_4210;
wire x_4211;
wire x_4212;
wire x_4213;
wire x_4214;
wire x_4215;
wire x_4216;
wire x_4217;
wire x_4218;
wire x_4219;
wire x_4220;
wire x_4221;
wire x_4222;
wire x_4223;
wire x_4224;
wire x_4225;
wire x_4226;
wire x_4227;
wire x_4228;
wire x_4229;
wire x_4230;
wire x_4231;
wire x_4232;
wire x_4233;
wire x_4234;
wire x_4235;
wire x_4236;
wire x_4237;
wire x_4238;
wire x_4239;
wire x_4240;
wire x_4241;
wire x_4242;
wire x_4243;
wire x_4244;
wire x_4245;
wire x_4246;
wire x_4247;
wire x_4248;
wire x_4249;
wire x_4250;
wire x_4251;
wire x_4252;
wire x_4253;
wire x_4254;
wire x_4255;
wire x_4256;
wire x_4257;
wire x_4258;
wire x_4259;
wire x_4260;
wire x_4261;
wire x_4262;
wire x_4263;
wire x_4264;
wire x_4265;
wire x_4266;
wire x_4267;
wire x_4268;
wire x_4269;
wire x_4270;
wire x_4271;
wire x_4272;
wire x_4273;
wire x_4274;
wire x_4275;
wire x_4276;
wire x_4277;
wire x_4278;
wire x_4279;
wire x_4280;
wire x_4281;
wire x_4282;
wire x_4283;
wire x_4284;
wire x_4285;
wire x_4286;
wire x_4287;
wire x_4288;
wire x_4289;
wire x_4290;
wire x_4291;
wire x_4292;
wire x_4293;
wire x_4294;
wire x_4295;
wire x_4296;
wire x_4297;
wire x_4298;
wire x_4299;
wire x_4300;
wire x_4301;
wire x_4302;
wire x_4303;
wire x_4304;
wire x_4305;
wire x_4306;
wire x_4307;
wire x_4308;
wire x_4309;
wire x_4310;
wire x_4311;
wire x_4312;
wire x_4313;
wire x_4314;
wire x_4315;
wire x_4316;
wire x_4317;
wire x_4318;
wire x_4319;
wire x_4320;
wire x_4321;
wire x_4322;
wire x_4323;
wire x_4324;
wire x_4325;
wire x_4326;
wire x_4327;
wire x_4328;
wire x_4329;
wire x_4330;
wire x_4331;
wire x_4332;
wire x_4333;
wire x_4334;
wire x_4335;
wire x_4336;
wire x_4337;
wire x_4338;
wire x_4339;
wire x_4340;
wire x_4341;
wire x_4342;
wire x_4343;
wire x_4344;
wire x_4345;
wire x_4346;
wire x_4347;
wire x_4348;
wire x_4349;
wire x_4350;
wire x_4351;
wire x_4352;
wire x_4353;
wire x_4354;
wire x_4355;
wire x_4356;
wire x_4357;
wire x_4358;
wire x_4359;
wire x_4360;
wire x_4361;
wire x_4362;
wire x_4363;
wire x_4364;
wire x_4365;
wire x_4366;
wire x_4367;
wire x_4368;
wire x_4369;
wire x_4370;
wire x_4371;
wire x_4372;
wire x_4373;
wire x_4374;
wire x_4375;
wire x_4376;
wire x_4377;
wire x_4378;
wire x_4379;
wire x_4380;
wire x_4381;
wire x_4382;
wire x_4383;
wire x_4384;
wire x_4385;
wire x_4386;
wire x_4387;
wire x_4388;
wire x_4389;
wire x_4390;
wire x_4391;
wire x_4392;
wire x_4393;
wire x_4394;
wire x_4395;
wire x_4396;
wire x_4397;
wire x_4398;
wire x_4399;
wire x_4400;
wire x_4401;
wire x_4402;
wire x_4403;
wire x_4404;
wire x_4405;
wire x_4406;
wire x_4407;
wire x_4408;
wire x_4409;
wire x_4410;
wire x_4411;
wire x_4412;
wire x_4413;
wire x_4414;
wire x_4415;
wire x_4416;
wire x_4417;
wire x_4418;
wire x_4419;
wire x_4420;
wire x_4421;
wire x_4422;
wire x_4423;
wire x_4424;
wire x_4425;
wire x_4426;
wire x_4427;
wire x_4428;
wire x_4429;
wire x_4430;
wire x_4431;
wire x_4432;
wire x_4433;
wire x_4434;
wire x_4435;
wire x_4436;
wire x_4437;
wire x_4438;
wire x_4439;
wire x_4440;
wire x_4441;
wire x_4442;
wire x_4443;
wire x_4444;
wire x_4445;
wire x_4446;
wire x_4447;
wire x_4448;
wire x_4449;
wire x_4450;
wire x_4451;
wire x_4452;
wire x_4453;
wire x_4454;
wire x_4455;
wire x_4456;
wire x_4457;
wire x_4458;
wire x_4459;
wire x_4460;
wire x_4461;
wire x_4462;
wire x_4463;
wire x_4464;
wire x_4465;
wire x_4466;
wire x_4467;
wire x_4468;
wire x_4469;
wire x_4470;
wire x_4471;
wire x_4472;
wire x_4473;
wire x_4474;
wire x_4475;
wire x_4476;
wire x_4477;
wire x_4478;
wire x_4479;
wire x_4480;
wire x_4481;
wire x_4482;
wire x_4483;
wire x_4484;
wire x_4485;
wire x_4486;
wire x_4487;
wire x_4488;
wire x_4489;
wire x_4490;
wire x_4491;
wire x_4492;
wire x_4493;
wire x_4494;
wire x_4495;
wire x_4496;
wire x_4497;
wire x_4498;
wire x_4499;
wire x_4500;
wire x_4501;
wire x_4502;
wire x_4503;
wire x_4504;
wire x_4505;
wire x_4506;
wire x_4507;
wire x_4508;
wire x_4509;
wire x_4510;
wire x_4511;
wire x_4512;
wire x_4513;
wire x_4514;
wire x_4515;
wire x_4516;
wire x_4517;
wire x_4518;
wire x_4519;
wire x_4520;
wire x_4521;
wire x_4522;
wire x_4523;
wire x_4524;
wire x_4525;
wire x_4526;
wire x_4527;
wire x_4528;
wire x_4529;
wire x_4530;
wire x_4531;
wire x_4532;
wire x_4533;
wire x_4534;
wire x_4535;
wire x_4536;
wire x_4537;
wire x_4538;
wire x_4539;
wire x_4540;
wire x_4541;
wire x_4542;
wire x_4543;
wire x_4544;
wire x_4545;
wire x_4546;
wire x_4547;
wire x_4548;
wire x_4549;
wire x_4550;
wire x_4551;
wire x_4552;
wire x_4553;
wire x_4554;
wire x_4555;
wire x_4556;
wire x_4557;
wire x_4558;
wire x_4559;
wire x_4560;
wire x_4561;
wire x_4562;
wire x_4563;
wire x_4564;
wire x_4565;
wire x_4566;
wire x_4567;
wire x_4568;
wire x_4569;
wire x_4570;
wire x_4571;
wire x_4572;
wire x_4573;
wire x_4574;
wire x_4575;
wire x_4576;
wire x_4577;
wire x_4578;
wire x_4579;
wire x_4580;
wire x_4581;
wire x_4582;
wire x_4583;
wire x_4584;
wire x_4585;
wire x_4586;
wire x_4587;
wire x_4588;
wire x_4589;
wire x_4590;
wire x_4591;
wire x_4592;
wire x_4593;
wire x_4594;
wire x_4595;
wire x_4596;
wire x_4597;
wire x_4598;
wire x_4599;
wire x_4600;
wire x_4601;
wire x_4602;
wire x_4603;
wire x_4604;
wire x_4605;
wire x_4606;
wire x_4607;
wire x_4608;
wire x_4609;
wire x_4610;
wire x_4611;
wire x_4612;
wire x_4613;
wire x_4614;
wire x_4615;
wire x_4616;
wire x_4617;
wire x_4618;
wire x_4619;
wire x_4620;
wire x_4621;
wire x_4622;
wire x_4623;
wire x_4624;
wire x_4625;
wire x_4626;
wire x_4627;
wire x_4628;
wire x_4629;
wire x_4630;
wire x_4631;
wire x_4632;
wire x_4633;
wire x_4634;
wire x_4635;
wire x_4636;
wire x_4637;
wire x_4638;
wire x_4639;
wire x_4640;
wire x_4641;
wire x_4642;
wire x_4643;
wire x_4644;
wire x_4645;
wire x_4646;
wire x_4647;
wire x_4648;
wire x_4649;
wire x_4650;
wire x_4651;
wire x_4652;
wire x_4653;
wire x_4654;
wire x_4655;
wire x_4656;
wire x_4657;
wire x_4658;
wire x_4659;
wire x_4660;
wire x_4661;
wire x_4662;
wire x_4663;
wire x_4664;
wire x_4665;
wire x_4666;
wire x_4667;
wire x_4668;
wire x_4669;
wire x_4670;
wire x_4671;
wire x_4672;
wire x_4673;
wire x_4674;
wire x_4675;
wire x_4676;
wire x_4677;
wire x_4678;
wire x_4679;
wire x_4680;
wire x_4681;
wire x_4682;
wire x_4683;
wire x_4684;
wire x_4685;
wire x_4686;
wire x_4687;
wire x_4688;
wire x_4689;
wire x_4690;
wire x_4691;
wire x_4692;
wire x_4693;
wire x_4694;
wire x_4695;
wire x_4696;
wire x_4697;
wire x_4698;
wire x_4699;
wire x_4700;
wire x_4701;
wire x_4702;
wire x_4703;
wire x_4704;
wire x_4705;
wire x_4706;
wire x_4707;
wire x_4708;
wire x_4709;
wire x_4710;
wire x_4711;
wire x_4712;
wire x_4713;
wire x_4714;
wire x_4715;
wire x_4716;
wire x_4717;
wire x_4718;
wire x_4719;
wire x_4720;
wire x_4721;
wire x_4722;
wire x_4723;
wire x_4724;
wire x_4725;
wire x_4726;
wire x_4727;
wire x_4728;
wire x_4729;
wire x_4730;
wire x_4731;
wire x_4732;
wire x_4733;
wire x_4734;
wire x_4735;
wire x_4736;
wire x_4737;
wire x_4738;
wire x_4739;
wire x_4740;
wire x_4741;
wire x_4742;
wire x_4743;
wire x_4744;
wire x_4745;
wire x_4746;
wire x_4747;
wire x_4748;
wire x_4749;
wire x_4750;
wire x_4751;
wire x_4752;
wire x_4753;
wire x_4754;
wire x_4755;
wire x_4756;
wire x_4757;
wire x_4758;
wire x_4759;
wire x_4760;
wire x_4761;
wire x_4762;
wire x_4763;
wire x_4764;
wire x_4765;
wire x_4766;
wire x_4767;
wire x_4768;
wire x_4769;
wire x_4770;
wire x_4771;
wire x_4772;
wire x_4773;
wire x_4774;
wire x_4775;
wire x_4776;
wire x_4777;
wire x_4778;
wire x_4779;
wire x_4780;
wire x_4781;
wire x_4782;
wire x_4783;
wire x_4784;
wire x_4785;
wire x_4786;
wire x_4787;
wire x_4788;
wire x_4789;
wire x_4790;
wire x_4791;
wire x_4792;
wire x_4793;
wire x_4794;
wire x_4795;
wire x_4796;
wire x_4797;
wire x_4798;
wire x_4799;
wire x_4800;
wire x_4801;
wire x_4802;
wire x_4803;
wire x_4804;
wire x_4805;
wire x_4806;
wire x_4807;
wire x_4808;
wire x_4809;
wire x_4810;
wire x_4811;
wire x_4812;
wire x_4813;
wire x_4814;
wire x_4815;
wire x_4816;
wire x_4817;
wire x_4818;
wire x_4819;
wire x_4820;
wire x_4821;
wire x_4822;
wire x_4823;
wire x_4824;
wire x_4825;
wire x_4826;
wire x_4827;
wire x_4828;
wire x_4829;
wire x_4830;
wire x_4831;
wire x_4832;
wire x_4833;
wire x_4834;
wire x_4835;
wire x_4836;
wire x_4837;
wire x_4838;
wire x_4839;
wire x_4840;
wire x_4841;
wire x_4842;
wire x_4843;
wire x_4844;
wire x_4845;
wire x_4846;
wire x_4847;
wire x_4848;
wire x_4849;
wire x_4850;
wire x_4851;
wire x_4852;
wire x_4853;
wire x_4854;
wire x_4855;
wire x_4856;
wire x_4857;
wire x_4858;
wire x_4859;
wire x_4860;
wire x_4861;
wire x_4862;
wire x_4863;
wire x_4864;
wire x_4865;
wire x_4866;
wire x_4867;
wire x_4868;
wire x_4869;
wire x_4870;
wire x_4871;
wire x_4872;
wire x_4873;
wire x_4874;
wire x_4875;
wire x_4876;
wire x_4877;
wire x_4878;
wire x_4879;
wire x_4880;
wire x_4881;
wire x_4882;
wire x_4883;
wire x_4884;
wire x_4885;
wire x_4886;
wire x_4887;
wire x_4888;
wire x_4889;
wire x_4890;
wire x_4891;
wire x_4892;
wire x_4893;
wire x_4894;
wire x_4895;
wire x_4896;
wire x_4897;
wire x_4898;
wire x_4899;
wire x_4900;
wire x_4901;
wire x_4902;
wire x_4903;
wire x_4904;
wire x_4905;
wire x_4906;
wire x_4907;
wire x_4908;
wire x_4909;
wire x_4910;
wire x_4911;
wire x_4912;
wire x_4913;
wire x_4914;
wire x_4915;
wire x_4916;
wire x_4917;
wire x_4918;
wire x_4919;
wire x_4920;
wire x_4921;
wire x_4922;
wire x_4923;
wire x_4924;
wire x_4925;
wire x_4926;
wire x_4927;
wire x_4928;
wire x_4929;
wire x_4930;
wire x_4931;
wire x_4932;
wire x_4933;
wire x_4934;
wire x_4935;
wire x_4936;
wire x_4937;
wire x_4938;
wire x_4939;
wire x_4940;
wire x_4941;
wire x_4942;
wire x_4943;
wire x_4944;
wire x_4945;
wire x_4946;
wire x_4947;
wire x_4948;
wire x_4949;
wire x_4950;
wire x_4951;
wire x_4952;
wire x_4953;
wire x_4954;
wire x_4955;
wire x_4956;
wire x_4957;
wire x_4958;
wire x_4959;
wire x_4960;
wire x_4961;
wire x_4962;
wire x_4963;
wire x_4964;
wire x_4965;
wire x_4966;
wire x_4967;
wire x_4968;
wire x_4969;
wire x_4970;
wire x_4971;
wire x_4972;
wire x_4973;
wire x_4974;
wire x_4975;
wire x_4976;
wire x_4977;
wire x_4978;
wire x_4979;
wire x_4980;
wire x_4981;
wire x_4982;
wire x_4983;
wire x_4984;
wire x_4985;
wire x_4986;
wire x_4987;
wire x_4988;
wire x_4989;
wire x_4990;
wire x_4991;
wire x_4992;
wire x_4993;
wire x_4994;
wire x_4995;
wire x_4996;
wire x_4997;
wire x_4998;
wire x_4999;
wire x_5000;
wire x_5001;
wire x_5002;
wire x_5003;
wire x_5004;
wire x_5005;
wire x_5006;
wire x_5007;
wire x_5008;
wire x_5009;
wire x_5010;
wire x_5011;
wire x_5012;
wire x_5013;
wire x_5014;
wire x_5015;
wire x_5016;
wire x_5017;
wire x_5018;
wire x_5019;
wire x_5020;
wire x_5021;
wire x_5022;
wire x_5023;
wire x_5024;
wire x_5025;
wire x_5026;
wire x_5027;
wire x_5028;
wire x_5029;
wire x_5030;
wire x_5031;
wire x_5032;
wire x_5033;
wire x_5034;
wire x_5035;
wire x_5036;
wire x_5037;
wire x_5038;
wire x_5039;
wire x_5040;
wire x_5041;
wire x_5042;
wire x_5043;
wire x_5044;
wire x_5045;
wire x_5046;
wire x_5047;
wire x_5048;
wire x_5049;
wire x_5050;
wire x_5051;
wire x_5052;
wire x_5053;
wire x_5054;
wire x_5055;
wire x_5056;
wire x_5057;
wire x_5058;
wire x_5059;
wire x_5060;
wire x_5061;
wire x_5062;
wire x_5063;
wire x_5064;
wire x_5065;
wire x_5066;
wire x_5067;
wire x_5068;
wire x_5069;
wire x_5070;
wire x_5071;
wire x_5072;
wire x_5073;
wire x_5074;
wire x_5075;
wire x_5076;
wire x_5077;
wire x_5078;
wire x_5079;
wire x_5080;
wire x_5081;
wire x_5082;
wire x_5083;
wire x_5084;
wire x_5085;
wire x_5086;
wire x_5087;
wire x_5088;
wire x_5089;
wire x_5090;
wire x_5091;
wire x_5092;
wire x_5093;
wire x_5094;
wire x_5095;
wire x_5096;
wire x_5097;
wire x_5098;
wire x_5099;
wire x_5100;
wire x_5101;
wire x_5102;
wire x_5103;
wire x_5104;
wire x_5105;
wire x_5106;
wire x_5107;
wire x_5108;
wire x_5109;
wire x_5110;
wire x_5111;
wire x_5112;
wire x_5113;
wire x_5114;
wire x_5115;
wire x_5116;
wire x_5117;
wire x_5118;
wire x_5119;
wire x_5120;
wire x_5121;
wire x_5122;
wire x_5123;
wire x_5124;
wire x_5125;
wire x_5126;
wire x_5127;
wire x_5128;
wire x_5129;
wire x_5130;
wire x_5131;
wire x_5132;
wire x_5133;
wire x_5134;
wire x_5135;
wire x_5136;
wire x_5137;
wire x_5138;
wire x_5139;
wire x_5140;
wire x_5141;
wire x_5142;
wire x_5143;
wire x_5144;
wire x_5145;
wire x_5146;
wire x_5147;
wire x_5148;
wire x_5149;
wire x_5150;
wire x_5151;
wire x_5152;
wire x_5153;
wire x_5154;
wire x_5155;
wire x_5156;
wire x_5157;
wire x_5158;
wire x_5159;
wire x_5160;
wire x_5161;
wire x_5162;
wire x_5163;
wire x_5164;
wire x_5165;
wire x_5166;
wire x_5167;
wire x_5168;
wire x_5169;
wire x_5170;
wire x_5171;
wire x_5172;
wire x_5173;
wire x_5174;
wire x_5175;
wire x_5176;
wire x_5177;
wire x_5178;
wire x_5179;
wire x_5180;
wire x_5181;
wire x_5182;
wire x_5183;
wire x_5184;
wire x_5185;
wire x_5186;
wire x_5187;
wire x_5188;
wire x_5189;
wire x_5190;
wire x_5191;
wire x_5192;
wire x_5193;
wire x_5194;
wire x_5195;
wire x_5196;
wire x_5197;
wire x_5198;
wire x_5199;
wire x_5200;
wire x_5201;
wire x_5202;
wire x_5203;
wire x_5204;
wire x_5205;
wire x_5206;
wire x_5207;
wire x_5208;
wire x_5209;
wire x_5210;
wire x_5211;
wire x_5212;
wire x_5213;
wire x_5214;
wire x_5215;
wire x_5216;
wire x_5217;
wire x_5218;
wire x_5219;
wire x_5220;
wire x_5221;
wire x_5222;
wire x_5223;
wire x_5224;
wire x_5225;
wire x_5226;
wire x_5227;
wire x_5228;
wire x_5229;
wire x_5230;
wire x_5231;
wire x_5232;
wire x_5233;
wire x_5234;
wire x_5235;
wire x_5236;
wire x_5237;
wire x_5238;
wire x_5239;
wire x_5240;
wire x_5241;
wire x_5242;
wire x_5243;
wire x_5244;
wire x_5245;
wire x_5246;
wire x_5247;
wire x_5248;
wire x_5249;
wire x_5250;
wire x_5251;
wire x_5252;
wire x_5253;
wire x_5254;
wire x_5255;
wire x_5256;
wire x_5257;
wire x_5258;
wire x_5259;
wire x_5260;
wire x_5261;
wire x_5262;
wire x_5263;
wire x_5264;
wire x_5265;
wire x_5266;
wire x_5267;
wire x_5268;
wire x_5269;
wire x_5270;
wire x_5271;
wire x_5272;
wire x_5273;
wire x_5274;
wire x_5275;
wire x_5276;
wire x_5277;
wire x_5278;
wire x_5279;
wire x_5280;
wire x_5281;
wire x_5282;
wire x_5283;
wire x_5284;
wire x_5285;
wire x_5286;
wire x_5287;
wire x_5288;
wire x_5289;
wire x_5290;
wire x_5291;
wire x_5292;
wire x_5293;
wire x_5294;
wire x_5295;
wire x_5296;
wire x_5297;
wire x_5298;
wire x_5299;
wire x_5300;
wire x_5301;
wire x_5302;
wire x_5303;
wire x_5304;
wire x_5305;
wire x_5306;
wire x_5307;
wire x_5308;
wire x_5309;
wire x_5310;
wire x_5311;
wire x_5312;
wire x_5313;
wire x_5314;
wire x_5315;
wire x_5316;
wire x_5317;
wire x_5318;
wire x_5319;
wire x_5320;
wire x_5321;
wire x_5322;
wire x_5323;
wire x_5324;
wire x_5325;
wire x_5326;
wire x_5327;
wire x_5328;
wire x_5329;
wire x_5330;
wire x_5331;
wire x_5332;
wire x_5333;
wire x_5334;
wire x_5335;
wire x_5336;
wire x_5337;
wire x_5338;
wire x_5339;
wire x_5340;
wire x_5341;
wire x_5342;
wire x_5343;
wire x_5344;
wire x_5345;
wire x_5346;
wire x_5347;
wire x_5348;
wire x_5349;
wire x_5350;
wire x_5351;
wire x_5352;
wire x_5353;
wire x_5354;
wire x_5355;
wire x_5356;
wire x_5357;
wire x_5358;
wire x_5359;
wire x_5360;
wire x_5361;
wire x_5362;
wire x_5363;
wire x_5364;
wire x_5365;
wire x_5366;
wire x_5367;
wire x_5368;
wire x_5369;
wire x_5370;
wire x_5371;
wire x_5372;
wire x_5373;
wire x_5374;
wire x_5375;
wire x_5376;
wire x_5377;
wire x_5378;
wire x_5379;
wire x_5380;
wire x_5381;
wire x_5382;
wire x_5383;
wire x_5384;
wire x_5385;
wire x_5386;
wire x_5387;
wire x_5388;
wire x_5389;
wire x_5390;
wire x_5391;
wire x_5392;
wire x_5393;
wire x_5394;
wire x_5395;
wire x_5396;
wire x_5397;
wire x_5398;
wire x_5399;
wire x_5400;
wire x_5401;
wire x_5402;
wire x_5403;
wire x_5404;
wire x_5405;
wire x_5406;
wire x_5407;
wire x_5408;
wire x_5409;
wire x_5410;
wire x_5411;
wire x_5412;
wire x_5413;
wire x_5414;
wire x_5415;
wire x_5416;
wire x_5417;
wire x_5418;
wire x_5419;
wire x_5420;
wire x_5421;
wire x_5422;
wire x_5423;
wire x_5424;
wire x_5425;
wire x_5426;
wire x_5427;
wire x_5428;
wire x_5429;
wire x_5430;
wire x_5431;
wire x_5432;
wire x_5433;
wire x_5434;
wire x_5435;
wire x_5436;
wire x_5437;
wire x_5438;
wire x_5439;
wire x_5440;
wire x_5441;
wire x_5442;
wire x_5443;
wire x_5444;
wire x_5445;
wire x_5446;
wire x_5447;
wire x_5448;
wire x_5449;
wire x_5450;
wire x_5451;
wire x_5452;
wire x_5453;
wire x_5454;
wire x_5455;
wire x_5456;
wire x_5457;
wire x_5458;
wire x_5459;
wire x_5460;
wire x_5461;
wire x_5462;
wire x_5463;
wire x_5464;
wire x_5465;
wire x_5466;
wire x_5467;
wire x_5468;
wire x_5469;
wire x_5470;
wire x_5471;
wire x_5472;
wire x_5473;
wire x_5474;
wire x_5475;
wire x_5476;
wire x_5477;
wire x_5478;
wire x_5479;
wire x_5480;
wire x_5481;
wire x_5482;
wire x_5483;
wire x_5484;
wire x_5485;
wire x_5486;
wire x_5487;
wire x_5488;
wire x_5489;
wire x_5490;
wire x_5491;
wire x_5492;
wire x_5493;
wire x_5494;
wire x_5495;
wire x_5496;
wire x_5497;
wire x_5498;
wire x_5499;
wire x_5500;
wire x_5501;
wire x_5502;
wire x_5503;
wire x_5504;
wire x_5505;
wire x_5506;
wire x_5507;
wire x_5508;
wire x_5509;
wire x_5510;
wire x_5511;
wire x_5512;
wire x_5513;
wire x_5514;
wire x_5515;
wire x_5516;
wire x_5517;
wire x_5518;
wire x_5519;
wire x_5520;
wire x_5521;
wire x_5522;
wire x_5523;
wire x_5524;
wire x_5525;
wire x_5526;
wire x_5527;
wire x_5528;
wire x_5529;
wire x_5530;
wire x_5531;
wire x_5532;
wire x_5533;
wire x_5534;
wire x_5535;
wire x_5536;
wire x_5537;
wire x_5538;
wire x_5539;
wire x_5540;
wire x_5541;
wire x_5542;
wire x_5543;
wire x_5544;
wire x_5545;
wire x_5546;
wire x_5547;
wire x_5548;
wire x_5549;
wire x_5550;
wire x_5551;
wire x_5552;
wire x_5553;
wire x_5554;
wire x_5555;
wire x_5556;
wire x_5557;
wire x_5558;
wire x_5559;
wire x_5560;
wire x_5561;
wire x_5562;
wire x_5563;
wire x_5564;
wire x_5565;
wire x_5566;
wire x_5567;
wire x_5568;
wire x_5569;
wire x_5570;
wire x_5571;
wire x_5572;
wire x_5573;
wire x_5574;
wire x_5575;
wire x_5576;
wire x_5577;
wire x_5578;
wire x_5579;
wire x_5580;
wire x_5581;
wire x_5582;
wire x_5583;
wire x_5584;
wire x_5585;
wire x_5586;
wire x_5587;
wire x_5588;
wire x_5589;
wire x_5590;
wire x_5591;
wire x_5592;
wire x_5593;
wire x_5594;
wire x_5595;
wire x_5596;
wire x_5597;
wire x_5598;
wire x_5599;
wire x_5600;
wire x_5601;
wire x_5602;
wire x_5603;
wire x_5604;
wire x_5605;
wire x_5606;
wire x_5607;
wire x_5608;
wire x_5609;
wire x_5610;
wire x_5611;
wire x_5612;
wire x_5613;
wire x_5614;
wire x_5615;
wire x_5616;
wire x_5617;
wire x_5618;
wire x_5619;
wire x_5620;
wire x_5621;
wire x_5622;
wire x_5623;
wire x_5624;
wire x_5625;
wire x_5626;
wire x_5627;
wire x_5628;
wire x_5629;
wire x_5630;
wire x_5631;
wire x_5632;
wire x_5633;
wire x_5634;
wire x_5635;
wire x_5636;
wire x_5637;
wire x_5638;
wire x_5639;
wire x_5640;
wire x_5641;
wire x_5642;
wire x_5643;
wire x_5644;
wire x_5645;
wire x_5646;
wire x_5647;
wire x_5648;
wire x_5649;
wire x_5650;
wire x_5651;
wire x_5652;
wire x_5653;
wire x_5654;
wire x_5655;
wire x_5656;
wire x_5657;
wire x_5658;
wire x_5659;
wire x_5660;
wire x_5661;
wire x_5662;
wire x_5663;
wire x_5664;
wire x_5665;
wire x_5666;
wire x_5667;
wire x_5668;
wire x_5669;
wire x_5670;
wire x_5671;
wire x_5672;
wire x_5673;
wire x_5674;
wire x_5675;
wire x_5676;
wire x_5677;
wire x_5678;
wire x_5679;
wire x_5680;
wire x_5681;
wire x_5682;
wire x_5683;
wire x_5684;
wire x_5685;
wire x_5686;
wire x_5687;
wire x_5688;
wire x_5689;
wire x_5690;
wire x_5691;
wire x_5692;
wire x_5693;
wire x_5694;
wire x_5695;
wire x_5696;
wire x_5697;
wire x_5698;
wire x_5699;
wire x_5700;
wire x_5701;
wire x_5702;
wire x_5703;
wire x_5704;
wire x_5705;
wire x_5706;
wire x_5707;
wire x_5708;
wire x_5709;
wire x_5710;
wire x_5711;
wire x_5712;
wire x_5713;
wire x_5714;
wire x_5715;
wire x_5716;
wire x_5717;
wire x_5718;
wire x_5719;
wire x_5720;
wire x_5721;
wire x_5722;
wire x_5723;
wire x_5724;
wire x_5725;
wire x_5726;
wire x_5727;
wire x_5728;
wire x_5729;
wire x_5730;
wire x_5731;
wire x_5732;
wire x_5733;
wire x_5734;
wire x_5735;
wire x_5736;
wire x_5737;
wire x_5738;
wire x_5739;
wire x_5740;
wire x_5741;
wire x_5742;
wire x_5743;
wire x_5744;
wire x_5745;
wire x_5746;
wire x_5747;
wire x_5748;
wire x_5749;
wire x_5750;
wire x_5751;
wire x_5752;
wire x_5753;
wire x_5754;
wire x_5755;
wire x_5756;
wire x_5757;
wire x_5758;
wire x_5759;
wire x_5760;
wire x_5761;
wire x_5762;
wire x_5763;
wire x_5764;
wire x_5765;
wire x_5766;
wire x_5767;
wire x_5768;
wire x_5769;
wire x_5770;
wire x_5771;
wire x_5772;
wire x_5773;
wire x_5774;
wire x_5775;
wire x_5776;
wire x_5777;
wire x_5778;
wire x_5779;
wire x_5780;
wire x_5781;
wire x_5782;
wire x_5783;
wire x_5784;
wire x_5785;
wire x_5786;
wire x_5787;
wire x_5788;
wire x_5789;
wire x_5790;
wire x_5791;
wire x_5792;
wire x_5793;
wire x_5794;
wire x_5795;
wire x_5796;
wire x_5797;
wire x_5798;
wire x_5799;
wire x_5800;
wire x_5801;
wire x_5802;
wire x_5803;
wire x_5804;
wire x_5805;
wire x_5806;
wire x_5807;
wire x_5808;
wire x_5809;
wire x_5810;
wire x_5811;
wire x_5812;
wire x_5813;
wire x_5814;
wire x_5815;
wire x_5816;
wire x_5817;
wire x_5818;
wire x_5819;
wire x_5820;
wire x_5821;
wire x_5822;
wire x_5823;
wire x_5824;
wire x_5825;
wire x_5826;
wire x_5827;
wire x_5828;
wire x_5829;
wire x_5830;
wire x_5831;
wire x_5832;
wire x_5833;
wire x_5834;
wire x_5835;
wire x_5836;
wire x_5837;
wire x_5838;
wire x_5839;
wire x_5840;
wire x_5841;
wire x_5842;
wire x_5843;
wire x_5844;
wire x_5845;
wire x_5846;
wire x_5847;
wire x_5848;
wire x_5849;
wire x_5850;
wire x_5851;
wire x_5852;
wire x_5853;
wire x_5854;
wire x_5855;
wire x_5856;
wire x_5857;
wire x_5858;
wire x_5859;
wire x_5860;
wire x_5861;
wire x_5862;
wire x_5863;
wire x_5864;
wire x_5865;
wire x_5866;
wire x_5867;
wire x_5868;
wire x_5869;
wire x_5870;
wire x_5871;
wire x_5872;
wire x_5873;
wire x_5874;
wire x_5875;
wire x_5876;
wire x_5877;
wire x_5878;
wire x_5879;
wire x_5880;
wire x_5881;
wire x_5882;
wire x_5883;
wire x_5884;
wire x_5885;
wire x_5886;
wire x_5887;
wire x_5888;
wire x_5889;
wire x_5890;
wire x_5891;
wire x_5892;
wire x_5893;
wire x_5894;
wire x_5895;
wire x_5896;
wire x_5897;
wire x_5898;
wire x_5899;
wire x_5900;
wire x_5901;
wire x_5902;
wire x_5903;
wire x_5904;
wire x_5905;
wire x_5906;
wire x_5907;
wire x_5908;
wire x_5909;
wire x_5910;
wire x_5911;
wire x_5912;
wire x_5913;
wire x_5914;
wire x_5915;
wire x_5916;
wire x_5917;
wire x_5918;
wire x_5919;
wire x_5920;
wire x_5921;
wire x_5922;
wire x_5923;
wire x_5924;
wire x_5925;
wire x_5926;
wire x_5927;
wire x_5928;
wire x_5929;
wire x_5930;
wire x_5931;
wire x_5932;
wire x_5933;
wire x_5934;
wire x_5935;
wire x_5936;
wire x_5937;
wire x_5938;
wire x_5939;
wire x_5940;
wire x_5941;
wire x_5942;
wire x_5943;
wire x_5944;
wire x_5945;
wire x_5946;
wire x_5947;
wire x_5948;
wire x_5949;
wire x_5950;
wire x_5951;
wire x_5952;
wire x_5953;
wire x_5954;
wire x_5955;
wire x_5956;
wire x_5957;
wire x_5958;
wire x_5959;
wire x_5960;
wire x_5961;
wire x_5962;
wire x_5963;
wire x_5964;
wire x_5965;
wire x_5966;
wire x_5967;
wire x_5968;
wire x_5969;
wire x_5970;
wire x_5971;
wire x_5972;
wire x_5973;
wire x_5974;
wire x_5975;
wire x_5976;
wire x_5977;
wire x_5978;
wire x_5979;
wire x_5980;
wire x_5981;
wire x_5982;
wire x_5983;
wire x_5984;
wire x_5985;
wire x_5986;
wire x_5987;
wire x_5988;
wire x_5989;
wire x_5990;
wire x_5991;
wire x_5992;
wire x_5993;
wire x_5994;
wire x_5995;
wire x_5996;
wire x_5997;
wire x_5998;
wire x_5999;
wire x_6000;
wire x_6001;
wire x_6002;
wire x_6003;
wire x_6004;
wire x_6005;
wire x_6006;
wire x_6007;
wire x_6008;
wire x_6009;
wire x_6010;
wire x_6011;
wire x_6012;
wire x_6013;
wire x_6014;
wire x_6015;
wire x_6016;
wire x_6017;
wire x_6018;
wire x_6019;
wire x_6020;
wire x_6021;
wire x_6022;
wire x_6023;
wire x_6024;
wire x_6025;
wire x_6026;
wire x_6027;
wire x_6028;
wire x_6029;
wire x_6030;
wire x_6031;
wire x_6032;
wire x_6033;
wire x_6034;
wire x_6035;
wire x_6036;
wire x_6037;
wire x_6038;
wire x_6039;
wire x_6040;
wire x_6041;
wire x_6042;
wire x_6043;
wire x_6044;
wire x_6045;
wire x_6046;
wire x_6047;
wire x_6048;
wire x_6049;
wire x_6050;
wire x_6051;
wire x_6052;
wire x_6053;
wire x_6054;
wire x_6055;
wire x_6056;
wire x_6057;
wire x_6058;
wire x_6059;
wire x_6060;
wire x_6061;
wire x_6062;
wire x_6063;
wire x_6064;
wire x_6065;
wire x_6066;
wire x_6067;
wire x_6068;
wire x_6069;
wire x_6070;
wire x_6071;
wire x_6072;
wire x_6073;
wire x_6074;
wire x_6075;
wire x_6076;
wire x_6077;
wire x_6078;
wire x_6079;
wire x_6080;
wire x_6081;
wire x_6082;
wire x_6083;
wire x_6084;
wire x_6085;
wire x_6086;
wire x_6087;
wire x_6088;
wire x_6089;
wire x_6090;
wire x_6091;
wire x_6092;
wire x_6093;
wire x_6094;
wire x_6095;
wire x_6096;
wire x_6097;
wire x_6098;
wire x_6099;
wire x_6100;
wire x_6101;
wire x_6102;
wire x_6103;
wire x_6104;
wire x_6105;
wire x_6106;
wire x_6107;
wire x_6108;
wire x_6109;
wire x_6110;
wire x_6111;
wire x_6112;
wire x_6113;
wire x_6114;
wire x_6115;
wire x_6116;
wire x_6117;
wire x_6118;
wire x_6119;
wire x_6120;
wire x_6121;
wire x_6122;
wire x_6123;
wire x_6124;
wire x_6125;
wire x_6126;
wire x_6127;
wire x_6128;
wire x_6129;
wire x_6130;
wire x_6131;
wire x_6132;
wire x_6133;
wire x_6134;
wire x_6135;
wire x_6136;
wire x_6137;
wire x_6138;
wire x_6139;
wire x_6140;
wire x_6141;
wire x_6142;
wire x_6143;
wire x_6144;
wire x_6145;
wire x_6146;
wire x_6147;
wire x_6148;
wire x_6149;
wire x_6150;
wire x_6151;
wire x_6152;
wire x_6153;
wire x_6154;
wire x_6155;
wire x_6156;
wire x_6157;
wire x_6158;
wire x_6159;
wire x_6160;
wire x_6161;
wire x_6162;
wire x_6163;
wire x_6164;
wire x_6165;
wire x_6166;
wire x_6167;
wire x_6168;
wire x_6169;
wire x_6170;
wire x_6171;
wire x_6172;
wire x_6173;
wire x_6174;
wire x_6175;
wire x_6176;
wire x_6177;
wire x_6178;
wire x_6179;
wire x_6180;
wire x_6181;
wire x_6182;
wire x_6183;
wire x_6184;
wire x_6185;
wire x_6186;
wire x_6187;
wire x_6188;
wire x_6189;
wire x_6190;
wire x_6191;
wire x_6192;
wire x_6193;
wire x_6194;
wire x_6195;
wire x_6196;
wire x_6197;
wire x_6198;
wire x_6199;
wire x_6200;
wire x_6201;
wire x_6202;
wire x_6203;
wire x_6204;
wire x_6205;
wire x_6206;
wire x_6207;
wire x_6208;
wire x_6209;
wire x_6210;
wire x_6211;
wire x_6212;
wire x_6213;
wire x_6214;
wire x_6215;
wire x_6216;
wire x_6217;
wire x_6218;
wire x_6219;
wire x_6220;
wire x_6221;
wire x_6222;
wire x_6223;
wire x_6224;
wire x_6225;
wire x_6226;
wire x_6227;
wire x_6228;
wire x_6229;
wire x_6230;
wire x_6231;
wire x_6232;
wire x_6233;
wire x_6234;
wire x_6235;
wire x_6236;
wire x_6237;
wire x_6238;
wire x_6239;
wire x_6240;
wire x_6241;
wire x_6242;
wire x_6243;
wire x_6244;
wire x_6245;
wire x_6246;
wire x_6247;
wire x_6248;
wire x_6249;
wire x_6250;
wire x_6251;
wire x_6252;
wire x_6253;
wire x_6254;
wire x_6255;
wire x_6256;
wire x_6257;
wire x_6258;
wire x_6259;
wire x_6260;
wire x_6261;
wire x_6262;
wire x_6263;
wire x_6264;
wire x_6265;
wire x_6266;
wire x_6267;
wire x_6268;
wire x_6269;
wire x_6270;
wire x_6271;
wire x_6272;
wire x_6273;
wire x_6274;
wire x_6275;
wire x_6276;
wire x_6277;
wire x_6278;
wire x_6279;
wire x_6280;
wire x_6281;
wire x_6282;
wire x_6283;
wire x_6284;
wire x_6285;
wire x_6286;
wire x_6287;
wire x_6288;
wire x_6289;
wire x_6290;
wire x_6291;
wire x_6292;
wire x_6293;
wire x_6294;
wire x_6295;
wire x_6296;
wire x_6297;
wire x_6298;
wire x_6299;
wire x_6300;
wire x_6301;
wire x_6302;
wire x_6303;
wire x_6304;
wire x_6305;
wire x_6306;
wire x_6307;
wire x_6308;
wire x_6309;
wire x_6310;
wire x_6311;
wire x_6312;
wire x_6313;
wire x_6314;
wire x_6315;
wire x_6316;
wire x_6317;
wire x_6318;
wire x_6319;
wire x_6320;
wire x_6321;
wire x_6322;
wire x_6323;
wire x_6324;
wire x_6325;
wire x_6326;
wire x_6327;
wire x_6328;
wire x_6329;
wire x_6330;
wire x_6331;
wire x_6332;
wire x_6333;
wire x_6334;
wire x_6335;
wire x_6336;
wire x_6337;
wire x_6338;
wire x_6339;
wire x_6340;
wire x_6341;
wire x_6342;
wire x_6343;
wire x_6344;
wire x_6345;
wire x_6346;
wire x_6347;
wire x_6348;
wire x_6349;
wire x_6350;
wire x_6351;
wire x_6352;
wire x_6353;
wire x_6354;
wire x_6355;
wire x_6356;
wire x_6357;
wire x_6358;
wire x_6359;
wire x_6360;
wire x_6361;
wire x_6362;
wire x_6363;
wire x_6364;
wire x_6365;
wire x_6366;
wire x_6367;
wire x_6368;
wire x_6369;
wire x_6370;
wire x_6371;
wire x_6372;
wire x_6373;
wire x_6374;
wire x_6375;
wire x_6376;
wire x_6377;
wire x_6378;
wire x_6379;
wire x_6380;
wire x_6381;
wire x_6382;
wire x_6383;
wire x_6384;
wire x_6385;
wire x_6386;
wire x_6387;
wire x_6388;
wire x_6389;
wire x_6390;
wire x_6391;
wire x_6392;
wire x_6393;
wire x_6394;
wire x_6395;
wire x_6396;
wire x_6397;
wire x_6398;
wire x_6399;
wire x_6400;
wire x_6401;
wire x_6402;
wire x_6403;
wire x_6404;
wire x_6405;
wire x_6406;
wire x_6407;
wire x_6408;
wire x_6409;
wire x_6410;
wire x_6411;
wire x_6412;
wire x_6413;
wire x_6414;
wire x_6415;
wire x_6416;
wire x_6417;
wire x_6418;
wire x_6419;
wire x_6420;
wire x_6421;
wire x_6422;
wire x_6423;
wire x_6424;
wire x_6425;
wire x_6426;
wire x_6427;
wire x_6428;
wire x_6429;
wire x_6430;
wire x_6431;
wire x_6432;
wire x_6433;
wire x_6434;
wire x_6435;
wire x_6436;
wire x_6437;
wire x_6438;
wire x_6439;
wire x_6440;
wire x_6441;
wire x_6442;
wire x_6443;
wire x_6444;
wire x_6445;
wire x_6446;
wire x_6447;
wire x_6448;
wire x_6449;
wire x_6450;
wire x_6451;
wire x_6452;
wire x_6453;
wire x_6454;
wire x_6455;
wire x_6456;
wire x_6457;
wire x_6458;
wire x_6459;
wire x_6460;
wire x_6461;
wire x_6462;
wire x_6463;
wire x_6464;
wire x_6465;
wire x_6466;
wire x_6467;
wire x_6468;
wire x_6469;
wire x_6470;
wire x_6471;
wire x_6472;
wire x_6473;
wire x_6474;
wire x_6475;
wire x_6476;
wire x_6477;
wire x_6478;
wire x_6479;
wire x_6480;
wire x_6481;
wire x_6482;
wire x_6483;
wire x_6484;
wire x_6485;
wire x_6486;
wire x_6487;
wire x_6488;
wire x_6489;
wire x_6490;
wire x_6491;
wire x_6492;
wire x_6493;
wire x_6494;
wire x_6495;
wire x_6496;
wire x_6497;
wire x_6498;
wire x_6499;
wire x_6500;
wire x_6501;
wire x_6502;
wire x_6503;
wire x_6504;
wire x_6505;
wire x_6506;
wire x_6507;
wire x_6508;
wire x_6509;
wire x_6510;
wire x_6511;
wire x_6512;
wire x_6513;
wire x_6514;
wire x_6515;
wire x_6516;
wire x_6517;
wire x_6518;
wire x_6519;
wire x_6520;
wire x_6521;
wire x_6522;
wire x_6523;
wire x_6524;
wire x_6525;
wire x_6526;
wire x_6527;
wire x_6528;
wire x_6529;
wire x_6530;
wire x_6531;
wire x_6532;
wire x_6533;
wire x_6534;
wire x_6535;
wire x_6536;
wire x_6537;
wire x_6538;
wire x_6539;
wire x_6540;
wire x_6541;
wire x_6542;
wire x_6543;
wire x_6544;
wire x_6545;
wire x_6546;
wire x_6547;
wire x_6548;
wire x_6549;
wire x_6550;
wire x_6551;
wire x_6552;
wire x_6553;
wire x_6554;
wire x_6555;
wire x_6556;
wire x_6557;
wire x_6558;
wire x_6559;
wire x_6560;
wire x_6561;
wire x_6562;
wire x_6563;
wire x_6564;
wire x_6565;
wire x_6566;
wire x_6567;
wire x_6568;
wire x_6569;
wire x_6570;
wire x_6571;
wire x_6572;
wire x_6573;
wire x_6574;
wire x_6575;
wire x_6576;
wire x_6577;
wire x_6578;
wire x_6579;
wire x_6580;
wire x_6581;
wire x_6582;
wire x_6583;
wire x_6584;
wire x_6585;
wire x_6586;
wire x_6587;
wire x_6588;
wire x_6589;
wire x_6590;
wire x_6591;
wire x_6592;
wire x_6593;
wire x_6594;
wire x_6595;
wire x_6596;
wire x_6597;
wire x_6598;
wire x_6599;
wire x_6600;
wire x_6601;
wire x_6602;
wire x_6603;
wire x_6604;
wire x_6605;
wire x_6606;
wire x_6607;
wire x_6608;
wire x_6609;
wire x_6610;
wire x_6611;
wire x_6612;
wire x_6613;
wire x_6614;
wire x_6615;
wire x_6616;
wire x_6617;
wire x_6618;
wire x_6619;
wire x_6620;
wire x_6621;
wire x_6622;
wire x_6623;
wire x_6624;
wire x_6625;
wire x_6626;
wire x_6627;
wire x_6628;
wire x_6629;
wire x_6630;
wire x_6631;
wire x_6632;
wire x_6633;
wire x_6634;
wire x_6635;
wire x_6636;
wire x_6637;
wire x_6638;
wire x_6639;
wire x_6640;
wire x_6641;
wire x_6642;
wire x_6643;
wire x_6644;
wire x_6645;
wire x_6646;
wire x_6647;
wire x_6648;
wire x_6649;
wire x_6650;
wire x_6651;
wire x_6652;
wire x_6653;
wire x_6654;
wire x_6655;
wire x_6656;
wire x_6657;
wire x_6658;
wire x_6659;
wire x_6660;
wire x_6661;
wire x_6662;
wire x_6663;
wire x_6664;
wire x_6665;
wire x_6666;
wire x_6667;
wire x_6668;
wire x_6669;
wire x_6670;
wire x_6671;
wire x_6672;
wire x_6673;
wire x_6674;
wire x_6675;
wire x_6676;
wire x_6677;
wire x_6678;
wire x_6679;
wire x_6680;
wire x_6681;
wire x_6682;
wire x_6683;
wire x_6684;
wire x_6685;
wire x_6686;
wire x_6687;
wire x_6688;
wire x_6689;
wire x_6690;
wire x_6691;
wire x_6692;
wire x_6693;
wire x_6694;
wire x_6695;
wire x_6696;
wire x_6697;
wire x_6698;
wire x_6699;
wire x_6700;
wire x_6701;
wire x_6702;
wire x_6703;
wire x_6704;
wire x_6705;
wire x_6706;
wire x_6707;
wire x_6708;
wire x_6709;
wire x_6710;
wire x_6711;
wire x_6712;
wire x_6713;
wire x_6714;
wire x_6715;
wire x_6716;
wire x_6717;
wire x_6718;
wire x_6719;
wire x_6720;
wire x_6721;
wire x_6722;
wire x_6723;
wire x_6724;
wire x_6725;
wire x_6726;
wire x_6727;
wire x_6728;
wire x_6729;
wire x_6730;
wire x_6731;
wire x_6732;
wire x_6733;
wire x_6734;
wire x_6735;
wire x_6736;
wire x_6737;
wire x_6738;
wire x_6739;
wire x_6740;
wire x_6741;
wire x_6742;
wire x_6743;
wire x_6744;
wire x_6745;
wire x_6746;
wire x_6747;
wire x_6748;
wire x_6749;
wire x_6750;
wire x_6751;
wire x_6752;
wire x_6753;
wire x_6754;
wire x_6755;
wire x_6756;
wire x_6757;
wire x_6758;
wire x_6759;
wire x_6760;
wire x_6761;
wire x_6762;
wire x_6763;
wire x_6764;
wire x_6765;
wire x_6766;
wire x_6767;
wire x_6768;
wire x_6769;
wire x_6770;
wire x_6771;
wire x_6772;
wire x_6773;
wire x_6774;
wire x_6775;
wire x_6776;
wire x_6777;
wire x_6778;
wire x_6779;
wire x_6780;
wire x_6781;
wire x_6782;
wire x_6783;
wire x_6784;
wire x_6785;
wire x_6786;
wire x_6787;
wire x_6788;
wire x_6789;
wire x_6790;
wire x_6791;
wire x_6792;
wire x_6793;
wire x_6794;
wire x_6795;
wire x_6796;
wire x_6797;
wire x_6798;
wire x_6799;
wire x_6800;
wire x_6801;
wire x_6802;
wire x_6803;
wire x_6804;
wire x_6805;
wire x_6806;
wire x_6807;
wire x_6808;
wire x_6809;
wire x_6810;
wire x_6811;
wire x_6812;
wire x_6813;
wire x_6814;
wire x_6815;
wire x_6816;
wire x_6817;
wire x_6818;
wire x_6819;
wire x_6820;
wire x_6821;
wire x_6822;
wire x_6823;
wire x_6824;
wire x_6825;
wire x_6826;
wire x_6827;
wire x_6828;
wire x_6829;
wire x_6830;
wire x_6831;
wire x_6832;
wire x_6833;
wire x_6834;
wire x_6835;
wire x_6836;
wire x_6837;
wire x_6838;
wire x_6839;
wire x_6840;
wire x_6841;
wire x_6842;
wire x_6843;
wire x_6844;
wire x_6845;
wire x_6846;
wire x_6847;
wire x_6848;
wire x_6849;
wire x_6850;
wire x_6851;
wire x_6852;
wire x_6853;
wire x_6854;
wire x_6855;
wire x_6856;
wire x_6857;
wire x_6858;
wire x_6859;
wire x_6860;
wire x_6861;
wire x_6862;
wire x_6863;
wire x_6864;
wire x_6865;
wire x_6866;
wire x_6867;
wire x_6868;
wire x_6869;
wire x_6870;
wire x_6871;
wire x_6872;
wire x_6873;
wire x_6874;
wire x_6875;
wire x_6876;
wire x_6877;
wire x_6878;
wire x_6879;
wire x_6880;
wire x_6881;
wire x_6882;
wire x_6883;
wire x_6884;
wire x_6885;
wire x_6886;
wire x_6887;
wire x_6888;
wire x_6889;
wire x_6890;
wire x_6891;
wire x_6892;
wire x_6893;
wire x_6894;
wire x_6895;
wire x_6896;
wire x_6897;
wire x_6898;
wire x_6899;
wire x_6900;
wire x_6901;
wire x_6902;
wire x_6903;
wire x_6904;
wire x_6905;
wire x_6906;
wire x_6907;
wire x_6908;
wire x_6909;
wire x_6910;
wire x_6911;
wire x_6912;
wire x_6913;
wire x_6914;
wire x_6915;
wire x_6916;
wire x_6917;
wire x_6918;
wire x_6919;
wire x_6920;
wire x_6921;
wire x_6922;
wire x_6923;
wire x_6924;
wire x_6925;
wire x_6926;
wire x_6927;
wire x_6928;
wire x_6929;
wire x_6930;
wire x_6931;
wire x_6932;
wire x_6933;
wire x_6934;
wire x_6935;
wire x_6936;
wire x_6937;
wire x_6938;
wire x_6939;
wire x_6940;
wire x_6941;
wire x_6942;
wire x_6943;
wire x_6944;
wire x_6945;
wire x_6946;
wire x_6947;
wire x_6948;
wire x_6949;
wire x_6950;
wire x_6951;
wire x_6952;
wire x_6953;
wire x_6954;
wire x_6955;
wire x_6956;
wire x_6957;
wire x_6958;
wire x_6959;
wire x_6960;
wire x_6961;
wire x_6962;
wire x_6963;
wire x_6964;
wire x_6965;
wire x_6966;
wire x_6967;
wire x_6968;
wire x_6969;
wire x_6970;
wire x_6971;
wire x_6972;
wire x_6973;
wire x_6974;
wire x_6975;
wire x_6976;
wire x_6977;
wire x_6978;
wire x_6979;
wire x_6980;
wire x_6981;
wire x_6982;
wire x_6983;
wire x_6984;
wire x_6985;
wire x_6986;
wire x_6987;
wire x_6988;
wire x_6989;
wire x_6990;
wire x_6991;
wire x_6992;
wire x_6993;
wire x_6994;
wire x_6995;
wire x_6996;
wire x_6997;
wire x_6998;
wire x_6999;
wire x_7000;
wire x_7001;
wire x_7002;
wire x_7003;
wire x_7004;
wire x_7005;
wire x_7006;
wire x_7007;
wire x_7008;
wire x_7009;
wire x_7010;
wire x_7011;
wire x_7012;
wire x_7013;
wire x_7014;
wire x_7015;
wire x_7016;
wire x_7017;
wire x_7018;
wire x_7019;
wire x_7020;
wire x_7021;
wire x_7022;
wire x_7023;
wire x_7024;
wire x_7025;
wire x_7026;
wire x_7027;
wire x_7028;
wire x_7029;
wire x_7030;
wire x_7031;
wire x_7032;
wire x_7033;
wire x_7034;
wire x_7035;
wire x_7036;
wire x_7037;
wire x_7038;
wire x_7039;
wire x_7040;
wire x_7041;
wire x_7042;
wire x_7043;
wire x_7044;
wire x_7045;
wire x_7046;
wire x_7047;
wire x_7048;
wire x_7049;
wire x_7050;
wire x_7051;
wire x_7052;
wire x_7053;
wire x_7054;
wire x_7055;
wire x_7056;
wire x_7057;
wire x_7058;
wire x_7059;
wire x_7060;
wire x_7061;
wire x_7062;
wire x_7063;
wire x_7064;
wire x_7065;
wire x_7066;
wire x_7067;
wire x_7068;
wire x_7069;
wire x_7070;
wire x_7071;
wire x_7072;
wire x_7073;
wire x_7074;
wire x_7075;
wire x_7076;
wire x_7077;
wire x_7078;
wire x_7079;
wire x_7080;
wire x_7081;
wire x_7082;
wire x_7083;
wire x_7084;
wire x_7085;
wire x_7086;
wire x_7087;
wire x_7088;
wire x_7089;
wire x_7090;
wire x_7091;
wire x_7092;
wire x_7093;
wire x_7094;
wire x_7095;
wire x_7096;
wire x_7097;
wire x_7098;
wire x_7099;
wire x_7100;
wire x_7101;
wire x_7102;
wire x_7103;
wire x_7104;
wire x_7105;
wire x_7106;
wire x_7107;
wire x_7108;
wire x_7109;
wire x_7110;
wire x_7111;
wire x_7112;
wire x_7113;
wire x_7114;
wire x_7115;
wire x_7116;
wire x_7117;
wire x_7118;
wire x_7119;
wire x_7120;
wire x_7121;
wire x_7122;
wire x_7123;
wire x_7124;
wire x_7125;
wire x_7126;
wire x_7127;
wire x_7128;
wire x_7129;
wire x_7130;
wire x_7131;
wire x_7132;
wire x_7133;
wire x_7134;
wire x_7135;
wire x_7136;
wire x_7137;
wire x_7138;
wire x_7139;
wire x_7140;
wire x_7141;
wire x_7142;
wire x_7143;
wire x_7144;
wire x_7145;
wire x_7146;
wire x_7147;
wire x_7148;
wire x_7149;
wire x_7150;
wire x_7151;
wire x_7152;
wire x_7153;
wire x_7154;
wire x_7155;
wire x_7156;
wire x_7157;
wire x_7158;
wire x_7159;
wire x_7160;
wire x_7161;
wire x_7162;
wire x_7163;
wire x_7164;
wire x_7165;
wire x_7166;
wire x_7167;
wire x_7168;
wire x_7169;
wire x_7170;
wire x_7171;
wire x_7172;
wire x_7173;
wire x_7174;
wire x_7175;
wire x_7176;
wire x_7177;
wire x_7178;
wire x_7179;
wire x_7180;
wire x_7181;
wire x_7182;
wire x_7183;
wire x_7184;
wire x_7185;
wire x_7186;
wire x_7187;
wire x_7188;
wire x_7189;
wire x_7190;
wire x_7191;
wire x_7192;
wire x_7193;
wire x_7194;
wire x_7195;
wire x_7196;
wire x_7197;
wire x_7198;
wire x_7199;
wire x_7200;
wire x_7201;
wire x_7202;
wire x_7203;
wire x_7204;
wire x_7205;
wire x_7206;
wire x_7207;
wire x_7208;
wire x_7209;
wire x_7210;
wire x_7211;
wire x_7212;
wire x_7213;
wire x_7214;
wire x_7215;
wire x_7216;
wire x_7217;
wire x_7218;
wire x_7219;
wire x_7220;
wire x_7221;
wire x_7222;
wire x_7223;
wire x_7224;
wire x_7225;
wire x_7226;
wire x_7227;
wire x_7228;
wire x_7229;
wire x_7230;
wire x_7231;
wire x_7232;
wire x_7233;
wire x_7234;
wire x_7235;
wire x_7236;
wire x_7237;
wire x_7238;
wire x_7239;
wire x_7240;
wire x_7241;
wire x_7242;
wire x_7243;
wire x_7244;
wire x_7245;
wire x_7246;
wire x_7247;
wire x_7248;
wire x_7249;
wire x_7250;
wire x_7251;
wire x_7252;
wire x_7253;
wire x_7254;
wire x_7255;
wire x_7256;
wire x_7257;
wire x_7258;
wire x_7259;
wire x_7260;
wire x_7261;
wire x_7262;
wire x_7263;
wire x_7264;
wire x_7265;
wire x_7266;
wire x_7267;
wire x_7268;
wire x_7269;
wire x_7270;
wire x_7271;
wire x_7272;
wire x_7273;
wire x_7274;
wire x_7275;
wire x_7276;
wire x_7277;
wire x_7278;
wire x_7279;
wire x_7280;
wire x_7281;
wire x_7282;
wire x_7283;
wire x_7284;
wire x_7285;
wire x_7286;
wire x_7287;
wire x_7288;
wire x_7289;
wire x_7290;
wire x_7291;
wire x_7292;
wire x_7293;
wire x_7294;
wire x_7295;
wire x_7296;
wire x_7297;
wire x_7298;
wire x_7299;
wire x_7300;
wire x_7301;
wire x_7302;
wire x_7303;
wire x_7304;
wire x_7305;
wire x_7306;
wire x_7307;
wire x_7308;
wire x_7309;
wire x_7310;
wire x_7311;
wire x_7312;
wire x_7313;
wire x_7314;
wire x_7315;
wire x_7316;
wire x_7317;
wire x_7318;
wire x_7319;
wire x_7320;
wire x_7321;
wire x_7322;
wire x_7323;
wire x_7324;
wire x_7325;
wire x_7326;
wire x_7327;
wire x_7328;
wire x_7329;
wire x_7330;
wire x_7331;
wire x_7332;
wire x_7333;
wire x_7334;
wire x_7335;
wire x_7336;
wire x_7337;
assign v_791 = 0;
assign v_790 = 0;
assign v_789 = 0;
assign v_788 = 0;
assign v_787 = 0;
assign v_786 = 0;
assign v_785 = 0;
assign v_784 = 0;
assign v_783 = 0;
assign v_782 = 0;
assign v_781 = 0;
assign v_780 = 0;
assign v_779 = 0;
assign v_778 = 0;
assign v_777 = 0;
assign v_776 = 0;
assign v_775 = 0;
assign v_774 = 0;
assign v_773 = 0;
assign v_772 = 0;
assign v_771 = 0;
assign v_685 = 0;
assign v_684 = 0;
assign v_683 = 0;
assign v_682 = 0;
assign v_681 = 0;
assign v_680 = 0;
assign v_679 = 0;
assign v_678 = 0;
assign v_677 = 0;
assign v_676 = 0;
assign v_675 = 0;
assign v_674 = 0;
assign v_673 = 0;
assign v_672 = 0;
assign v_671 = 0;
assign v_670 = 0;
assign v_669 = 0;
assign v_668 = 0;
assign v_667 = 0;
assign v_666 = 0;
assign v_665 = 0;
assign v_579 = 0;
assign v_578 = 0;
assign v_577 = 0;
assign v_576 = 0;
assign v_575 = 0;
assign v_574 = 0;
assign v_573 = 0;
assign v_572 = 0;
assign v_571 = 0;
assign v_570 = 0;
assign v_569 = 0;
assign v_568 = 0;
assign v_567 = 0;
assign v_566 = 0;
assign v_565 = 0;
assign v_564 = 0;
assign v_563 = 0;
assign v_562 = 0;
assign v_561 = 0;
assign v_560 = 0;
assign v_559 = 0;
assign v_473 = 0;
assign v_472 = 0;
assign v_471 = 0;
assign v_470 = 0;
assign v_469 = 0;
assign v_468 = 0;
assign v_467 = 0;
assign v_466 = 0;
assign v_465 = 0;
assign v_464 = 0;
assign v_463 = 0;
assign v_462 = 0;
assign v_461 = 0;
assign v_460 = 0;
assign v_459 = 0;
assign v_458 = 0;
assign v_457 = 0;
assign v_456 = 0;
assign v_455 = 0;
assign v_454 = 0;
assign v_453 = 0;
assign v_367 = 0;
assign v_366 = 0;
assign v_365 = 0;
assign v_364 = 0;
assign v_363 = 0;
assign v_362 = 0;
assign v_361 = 0;
assign v_360 = 0;
assign v_359 = 0;
assign v_358 = 0;
assign v_357 = 0;
assign v_356 = 0;
assign v_355 = 0;
assign v_354 = 0;
assign v_353 = 0;
assign v_352 = 0;
assign v_351 = 0;
assign v_350 = 0;
assign v_349 = 0;
assign v_348 = 0;
assign v_347 = 0;
assign x_1 = v_792 | v_793 | v_794 | v_795 | v_796 | v_797 | v_798 | v_799 | v_800 | v_801 | v_802 | v_803 | v_804 | v_805 | v_806 | v_807 | v_808 | v_809 | v_810 | v_811 | v_812 | v_813 | v_814 | v_815 | v_816 | v_817 | v_818 | v_819 | v_820 | v_821 | v_822 | v_823 | v_824 | v_825 | v_826 | v_827 | v_828 | v_829 | v_830 | v_831 | v_832 | v_833 | v_834 | v_835 | v_836 | v_837 | v_838 | v_839 | v_840 | v_841 | v_842 | v_843 | v_844 | v_845 | v_846 | v_847 | v_848 | v_849 | v_850 | v_851 | v_852 | v_853 | v_854 | v_855 | v_856 | v_857 | v_858 | v_859 | v_860 | v_861 | v_862 | v_863 | v_864 | v_865 | v_866 | v_867 | v_868 | v_869 | v_870 | v_871 | v_872 | v_873 | v_874 | v_875 | v_876 | v_877 | v_878 | v_879 | v_880 | v_881 | v_882 | v_883 | v_884 | v_885 | v_886 | v_887 | v_888 | v_889 | v_890 | v_891 | v_892 | v_893 | v_894 | v_895 | v_896 | v_897 | v_898 | v_899 | v_900 | v_901 | v_902 | v_903 | v_904 | v_905 | v_906 | v_907 | v_908 | v_909 | v_910 | v_911 | v_912 | v_913 | v_914 | v_915 | v_916 | v_917 | v_918 | v_919 | v_920 | v_921 | v_922 | v_923 | v_924 | v_925 | v_926 | v_927 | v_928 | v_929 | v_930 | v_931 | v_932 | v_933 | v_934 | v_935 | v_936 | v_937 | v_938 | v_939 | v_940 | v_941 | v_942 | v_943 | v_944 | v_945 | v_946 | v_947 | v_948 | v_949 | v_950 | v_951 | v_952 | v_953 | v_954 | v_955 | v_956 | v_957 | v_958 | v_959 | v_960 | v_961 | v_962 | v_963 | v_964 | v_965 | v_966 | v_967 | v_968 | v_969 | v_970 | v_971 | v_972 | v_973 | v_974 | v_975 | v_976 | v_977 | v_978 | v_979 | v_980 | v_981 | v_982 | v_983 | v_984 | v_985 | v_986 | v_987 | v_988 | v_989 | v_990 | v_991 | v_992 | v_993 | v_994 | v_995 | v_996 | v_997 | v_998 | v_999 | v_1000 | v_1001 | v_1002 | v_1003 | v_1004 | v_1005 | v_1006 | v_1007 | v_1008 | v_1009 | v_1010 | v_1011 | v_1012 | v_1013 | v_1014 | v_1015 | v_1016 | v_1017 | v_1018 | v_1019 | v_1020 | v_1021 | v_1022 | v_1023 | v_1024 | v_1025 | v_1026 | v_1027 | v_1028 | v_1029 | v_1030 | v_1031 | v_1032 | v_1033 | v_1034 | v_1035 | v_1036 | v_1037 | v_1038 | v_1039 | v_1040 | v_1041 | v_1042 | v_1043 | v_1044 | v_1045 | v_1046 | v_1047 | v_1048 | v_1049 | v_1050 | v_1051 | v_1052 | v_1053 | v_1054 | v_1055 | v_1056 | v_1057 | v_1058 | v_1059 | v_1060 | v_1061 | v_1062 | v_1063 | v_1064 | v_1065 | v_1066 | v_1067 | v_1068 | v_1069 | v_1070 | v_1071 | v_1072 | v_1073 | v_1074 | v_1075 | v_1076 | v_1077 | v_1078 | v_1079 | v_1080 | v_1081 | v_1082 | v_1083 | v_1084 | v_1085 | v_1086 | v_1087 | v_1088 | v_1089 | v_1090 | v_1091 | v_1092 | v_1093 | v_1094 | v_1095 | v_1096 | v_1097 | v_1098 | v_1099 | v_1100 | v_1101 | v_1102 | v_1103 | v_1104 | v_1105 | v_1106 | v_1107 | v_1108 | v_1109 | v_1110 | v_1111 | v_1112 | v_1113 | v_1114 | v_1115 | v_1116 | v_1117 | v_1118 | v_1119 | v_1120 | v_1121 | v_1122 | v_1123 | v_1124 | v_1125 | v_1126 | v_1127 | v_1128 | v_1129 | v_1130 | v_1131 | v_1132 | v_1133 | v_1134 | v_1135 | v_1136 | v_1137 | v_1138 | v_1139 | v_1140 | v_1141 | v_1142 | v_1143 | v_1144 | v_1145 | v_1146 | v_1147 | v_1148 | v_1149 | v_1150 | v_1151 | v_1152 | v_1153 | v_1154 | v_1155 | v_1156 | v_1157 | v_1158 | v_1159 | v_1160 | v_1161 | v_1162 | v_1163 | v_1164 | v_1165 | v_1166 | v_1167 | v_1168 | v_1169 | v_1170 | v_1171 | v_1172 | v_1173 | v_1174 | v_1175 | v_1176 | v_1177 | v_1178 | v_1179 | v_1180 | v_1181 | v_1182 | v_1183 | v_1184 | v_1185 | v_1186 | v_1187 | v_1188 | v_1189 | v_1190 | v_1191 | v_1192 | v_1193 | v_1194 | v_1195 | v_1196 | v_1197 | v_1198 | v_1199 | v_1200 | v_1201 | v_1202 | v_1203 | v_1204 | v_1205 | v_1206 | v_1207 | v_1208 | v_1209 | v_1210 | v_1211 | v_1212 | v_1213 | v_1214 | v_1215 | v_1216 | v_1217 | v_1218 | v_1219 | v_1220 | v_1221 | v_1222 | v_1223 | v_1224 | v_1225 | v_1226 | v_1227 | v_1228 | v_1229 | v_1230 | v_1231 | v_1232 | v_1233 | v_1234 | v_1235 | v_1236 | v_1237 | v_1238 | v_1239 | v_1240 | v_1241 | v_1242 | v_1243 | v_1244 | v_1245 | v_1246 | v_1247 | v_1248 | v_1249 | v_1250 | v_1251 | v_1252 | v_1253 | v_1254 | v_1255 | v_1256 | v_1257 | v_1258 | v_1259 | v_1260 | v_1261 | v_1262 | v_1263 | v_1264 | v_1265 | v_1266 | v_1267 | v_1268 | v_1269 | v_1270 | v_1271 | v_1272 | v_1273 | v_1274 | v_1275 | v_1276 | v_1277 | v_1278 | v_1279 | v_1280 | v_1281 | v_1282 | v_1283 | v_1284 | v_1285 | v_1286 | v_1287 | v_1288 | v_1289 | v_1290 | v_1291 | v_1292 | v_1293 | v_1294 | v_1295 | v_1296 | v_1297 | v_1298 | v_1299 | v_1300 | v_1301 | v_1302 | v_1303 | v_1304 | v_1305 | v_1306 | v_1307 | v_1308 | v_1309 | v_1310 | v_1311 | v_1312 | v_1313 | v_1314 | v_1315 | v_1316 | v_1317 | v_1318 | v_1319 | v_1320 | v_1321 | v_1322 | v_1323 | v_1324 | v_1325 | v_1326 | v_1327 | v_1328 | v_1329 | v_1330 | v_1331 | v_1332 | v_1333 | v_1334 | v_1335 | v_1336 | v_1337 | v_1338 | v_1339 | v_1340 | v_1341 | v_1342 | v_1343 | v_1344 | v_1345 | v_1346 | v_1347 | v_1348 | v_1349 | v_1350 | v_1351 | v_1352 | v_1353 | v_1354 | v_1355 | v_1356 | v_1357 | v_1358 | v_1359 | v_1360 | v_1361 | v_1362 | v_1363 | v_1364 | v_1365 | v_1366 | v_1367 | v_1368 | v_1369 | v_1370 | v_1371 | v_1372 | v_1373 | v_1374 | v_1375 | v_1376 | v_1377 | v_1378 | v_1379 | v_1380 | v_1381 | v_1382 | v_1383 | v_1384 | v_1385 | v_1386 | v_1387 | v_1388 | v_1389 | v_1390 | v_1391 | v_1392 | v_1393 | v_1394 | v_1395 | v_1396 | v_1397 | v_1398 | v_1399 | v_1400 | v_1401 | v_1402 | v_1403 | v_1404 | v_1405 | v_1406 | v_1407 | v_1408 | v_1409 | v_1410 | v_1411 | v_1412 | v_1413 | v_1414 | v_1415 | v_1416 | v_1417 | v_1418 | v_1419 | v_1420 | v_1421 | v_1422 | v_1423 | v_1424 | v_1425 | v_1426 | v_1427 | v_1428 | v_1429 | v_1430 | v_1431 | v_1432 | v_1433 | v_1434 | v_1435 | v_1436 | v_1437 | v_1438 | v_1439 | v_1440 | v_1441 | v_1442 | v_1443 | v_1444 | v_1445 | v_1446 | v_1447 | v_1448 | v_1449 | v_1450 | v_1451 | v_1452 | v_1453 | v_1454 | v_1455 | v_1456 | v_1457 | v_1458 | v_1459 | v_1460 | v_1461 | v_1462 | v_1463 | v_1464 | v_1465 | v_1466 | v_1467 | v_1468 | v_1469 | v_1470 | v_1471 | v_1472 | v_1473 | v_1474 | v_1475 | v_1476 | v_1477 | v_1478 | v_1479 | v_1480 | v_1481 | v_1482 | v_1483 | v_1484 | v_1485 | v_1486 | v_1487 | v_1488 | v_1489 | v_1490 | v_1491 | v_1492 | v_1493 | v_1494 | v_1495 | v_1496 | v_1497 | v_1498 | v_1499 | v_1500 | v_1501 | v_1502 | v_1503 | v_1504 | v_1505 | v_1506 | v_1507 | v_1508 | v_1509 | v_1510 | v_1511 | v_1512 | v_1513 | v_1514 | v_1515 | v_1516 | v_1517 | v_1518 | v_1519 | v_1520 | v_1521 | v_1522 | v_1523 | v_1524 | v_1525 | v_1526 | v_1527 | v_1528 | v_1529 | v_1530 | v_1531 | v_1532 | v_1533 | v_1534 | v_1535 | v_1536 | v_1537 | v_1538 | v_1539 | v_1540 | v_1541 | v_1542 | v_1543 | v_1544 | v_1545 | v_1546 | v_1547 | v_1548 | v_1549 | v_1550 | v_1551 | v_1552 | v_1553 | v_1554 | v_1555 | v_1556 | v_1557 | v_1558 | v_1559 | v_1560 | v_1561 | v_1562 | v_1563 | v_1564 | v_1565 | v_1566 | v_1567 | v_1568 | v_1569 | v_1570 | v_1571 | v_1572 | v_1573 | v_1574 | v_1575 | v_1576 | v_1577 | v_1578 | v_1579 | v_1580 | v_1581 | v_1582 | v_1583 | v_1584 | v_1585 | v_1586 | v_1587 | v_1588 | v_1589 | v_1590 | v_1591 | v_1592 | v_1593 | v_1594 | v_1595 | v_1596 | v_1597 | v_1598 | v_1599 | v_1600 | v_1601 | v_1602 | v_1603 | v_1604 | v_1605 | v_1606 | v_1607 | v_1608 | v_1609 | v_1610 | v_1611 | v_1612 | v_1613 | v_1614 | v_1615 | v_1616 | v_1617 | v_1618 | v_1619 | v_1620 | v_1621 | v_1622 | v_1623 | v_1624 | v_1625 | v_1626 | v_1627 | v_1628 | v_1629 | v_1630 | v_1631 | v_1632 | v_1633 | v_1634 | v_1635 | v_1636 | v_1637 | v_1638 | v_1639 | v_1640 | v_1641 | v_1642 | v_1643 | v_1644 | v_1645 | v_1646 | v_1647 | v_1648 | v_1649 | v_1650 | v_1651 | v_1652 | v_1653 | v_1654 | v_1655 | v_1656 | v_1657 | v_1658 | v_1659 | v_1660 | v_1661 | v_1662 | v_1663 | v_1664 | v_1665 | v_1666 | v_1667 | v_1668 | v_1669 | v_1670 | v_1671 | v_1672 | v_1673 | v_1674 | v_1675 | v_1676 | v_1677 | v_1678 | v_1679 | v_1680 | v_1681 | v_1682 | v_1683 | v_1684 | v_1685 | v_1686 | v_1687 | v_1688 | v_1689 | v_1690 | v_1691 | v_1692 | v_1693 | v_1694 | v_1695 | v_1696 | v_1697 | v_1698 | v_1699 | v_1700 | v_1701 | v_1702 | v_1703 | v_1704 | v_1705 | v_1706 | v_1707 | v_1708 | v_1709 | v_1710 | v_1711 | v_1712 | v_1713 | v_1714 | v_1715 | v_1716 | v_1717 | v_1718 | v_1719 | v_1720 | v_1721 | v_1722 | v_1723 | v_1724 | v_1725 | v_1726 | v_1727 | v_1728 | v_1729 | v_1730 | v_1731 | v_1732 | v_1733 | v_1734 | v_1735 | v_1736 | v_1737 | v_1738 | v_1739 | v_1740 | v_1741 | v_1742 | v_1743 | v_1744 | v_1745 | v_1746 | v_1747 | v_1748 | v_1749 | v_1750 | v_1751 | v_1752 | v_1753 | v_1754 | v_1755 | v_1756 | v_1757 | v_1758 | v_1759 | v_1760 | v_1761 | v_1762 | v_1763 | v_1764 | v_1765 | v_1766 | v_1767 | v_1768 | v_1769 | v_1770 | v_1771 | v_1772 | v_1773 | v_1774 | v_1775 | v_1776 | v_1777 | v_1778 | v_1779 | v_1780 | v_1781 | v_1782 | v_1783 | v_1784 | v_1785 | v_1786 | v_1787 | v_1788 | v_1789 | v_1790 | v_1791 | v_1792 | v_1793 | v_1794 | v_1795 | v_1796 | v_1797 | v_1798 | v_1799 | v_1800 | v_1801 | v_1802 | v_1803 | v_1804 | v_1805 | v_1806 | v_1807 | v_1808 | v_1809 | v_1810 | v_1811 | v_1812 | v_1813 | v_1814 | v_1815 | v_1816 | v_1817 | v_1818 | v_1819 | v_1820 | v_1821 | v_1822 | v_1823 | v_1824 | v_1825 | v_1826 | v_1827 | v_1828 | v_1829 | v_1830 | v_1831 | v_1832 | v_1833 | v_1834 | v_1835 | v_1836 | v_1837 | v_1838 | v_1839 | v_1840 | v_1841 | v_1842;
assign x_2 = ~v_792 | v_770;
assign x_3 = ~v_793 | v_182;
assign x_4 = ~v_793 | ~v_183;
assign x_5 = ~v_794 | v_54;
assign x_6 = ~v_794 | ~v_183;
assign x_7 = ~v_795 | v_182;
assign x_8 = ~v_795 | v_54;
assign x_9 = ~v_796 | v_181;
assign x_10 = ~v_796 | ~v_182;
assign x_11 = ~v_797 | v_53;
assign x_12 = ~v_797 | ~v_182;
assign x_13 = ~v_798 | v_181;
assign x_14 = ~v_798 | v_53;
assign x_15 = ~v_799 | v_180;
assign x_16 = ~v_799 | ~v_181;
assign x_17 = ~v_800 | v_52;
assign x_18 = ~v_800 | ~v_181;
assign x_19 = ~v_801 | v_180;
assign x_20 = ~v_801 | v_52;
assign x_21 = ~v_802 | v_179;
assign x_22 = ~v_802 | ~v_180;
assign x_23 = ~v_803 | v_51;
assign x_24 = ~v_803 | ~v_180;
assign x_25 = ~v_804 | v_179;
assign x_26 = ~v_804 | v_51;
assign x_27 = ~v_805 | v_49;
assign x_28 = ~v_805 | ~v_179;
assign x_29 = ~v_806 | v_50;
assign x_30 = ~v_806 | ~v_179;
assign x_31 = ~v_807 | v_49;
assign x_32 = ~v_807 | v_50;
assign x_33 = ~v_808 | v_177;
assign x_34 = ~v_808 | ~v_178;
assign x_35 = ~v_809 | v_59;
assign x_36 = ~v_809 | ~v_178;
assign x_37 = ~v_810 | v_177;
assign x_38 = ~v_810 | v_59;
assign x_39 = ~v_811 | v_176;
assign x_40 = ~v_811 | ~v_177;
assign x_41 = ~v_812 | v_58;
assign x_42 = ~v_812 | ~v_177;
assign x_43 = ~v_813 | v_176;
assign x_44 = ~v_813 | v_58;
assign x_45 = ~v_814 | v_175;
assign x_46 = ~v_814 | ~v_176;
assign x_47 = ~v_815 | v_57;
assign x_48 = ~v_815 | ~v_176;
assign x_49 = ~v_816 | v_175;
assign x_50 = ~v_816 | v_57;
assign x_51 = ~v_817 | v_55;
assign x_52 = ~v_817 | ~v_175;
assign x_53 = ~v_818 | v_56;
assign x_54 = ~v_818 | ~v_175;
assign x_55 = ~v_819 | v_55;
assign x_56 = ~v_819 | v_56;
assign x_57 = ~v_820 | v_49;
assign x_58 = ~v_820 | v_59;
assign x_59 = ~v_821 | v_49;
assign x_60 = ~v_821 | v_58;
assign x_61 = ~v_822 | v_49;
assign x_62 = ~v_822 | v_57;
assign x_63 = ~v_823 | v_49;
assign x_64 = ~v_823 | v_56;
assign x_65 = ~v_824 | v_49;
assign x_66 = ~v_824 | v_55;
assign x_67 = ~v_825 | v_173;
assign x_68 = ~v_825 | ~v_174;
assign x_69 = ~v_826 | v_63;
assign x_70 = ~v_826 | ~v_174;
assign x_71 = ~v_827 | v_173;
assign x_72 = ~v_827 | v_63;
assign x_73 = ~v_828 | v_172;
assign x_74 = ~v_828 | ~v_173;
assign x_75 = ~v_829 | v_62;
assign x_76 = ~v_829 | ~v_173;
assign x_77 = ~v_830 | v_172;
assign x_78 = ~v_830 | v_62;
assign x_79 = ~v_831 | v_60;
assign x_80 = ~v_831 | ~v_172;
assign x_81 = ~v_832 | v_61;
assign x_82 = ~v_832 | ~v_172;
assign x_83 = ~v_833 | v_60;
assign x_84 = ~v_833 | v_61;
assign x_85 = ~v_834 | v_171;
assign x_86 = ~v_834 | v_63;
assign x_87 = ~v_835 | v_171;
assign x_88 = ~v_835 | v_62;
assign x_89 = ~v_836 | v_171;
assign x_90 = ~v_836 | v_61;
assign x_91 = ~v_837 | v_171;
assign x_92 = ~v_837 | v_60;
assign x_93 = ~v_838 | v_50;
assign x_94 = ~v_838 | ~v_171;
assign x_95 = ~v_839 | v_55;
assign x_96 = ~v_839 | ~v_171;
assign x_97 = ~v_840 | v_50;
assign x_98 = ~v_840 | v_55;
assign x_99 = ~v_841 | v_169;
assign x_100 = ~v_841 | ~v_170;
assign x_101 = ~v_842 | v_66;
assign x_102 = ~v_842 | ~v_170;
assign x_103 = ~v_843 | v_169;
assign x_104 = ~v_843 | v_66;
assign x_105 = ~v_844 | v_64;
assign x_106 = ~v_844 | ~v_169;
assign x_107 = ~v_845 | v_65;
assign x_108 = ~v_845 | ~v_169;
assign x_109 = ~v_846 | v_64;
assign x_110 = ~v_846 | v_65;
assign x_111 = ~v_847 | v_168;
assign x_112 = ~v_847 | v_66;
assign x_113 = ~v_848 | v_168;
assign x_114 = ~v_848 | v_65;
assign x_115 = ~v_849 | v_168;
assign x_116 = ~v_849 | v_64;
assign x_117 = ~v_850 | v_167;
assign x_118 = ~v_850 | ~v_168;
assign x_119 = ~v_851 | v_60;
assign x_120 = ~v_851 | ~v_168;
assign x_121 = ~v_852 | v_167;
assign x_122 = ~v_852 | v_60;
assign x_123 = ~v_853 | v_51;
assign x_124 = ~v_853 | ~v_167;
assign x_125 = ~v_854 | v_56;
assign x_126 = ~v_854 | ~v_167;
assign x_127 = ~v_855 | v_51;
assign x_128 = ~v_855 | v_56;
assign x_129 = ~v_856 | v_67;
assign x_130 = ~v_856 | ~v_166;
assign x_131 = ~v_857 | v_68;
assign x_132 = ~v_857 | ~v_166;
assign x_133 = ~v_858 | v_67;
assign x_134 = ~v_858 | v_68;
assign x_135 = ~v_859 | v_165;
assign x_136 = ~v_859 | v_68;
assign x_137 = ~v_860 | v_165;
assign x_138 = ~v_860 | v_67;
assign x_139 = ~v_861 | v_164;
assign x_140 = ~v_861 | ~v_165;
assign x_141 = ~v_862 | v_64;
assign x_142 = ~v_862 | ~v_165;
assign x_143 = ~v_863 | v_164;
assign x_144 = ~v_863 | v_64;
assign x_145 = ~v_864 | v_163;
assign x_146 = ~v_864 | ~v_164;
assign x_147 = ~v_865 | v_61;
assign x_148 = ~v_865 | ~v_164;
assign x_149 = ~v_866 | v_163;
assign x_150 = ~v_866 | v_61;
assign x_151 = ~v_867 | v_52;
assign x_152 = ~v_867 | ~v_163;
assign x_153 = ~v_868 | v_57;
assign x_154 = ~v_868 | ~v_163;
assign x_155 = ~v_869 | v_52;
assign x_156 = ~v_869 | v_57;
assign x_157 = ~v_870 | v_162;
assign x_158 = ~v_870 | v_69;
assign x_159 = ~v_871 | v_161;
assign x_160 = ~v_871 | ~v_162;
assign x_161 = ~v_872 | v_67;
assign x_162 = ~v_872 | ~v_162;
assign x_163 = ~v_873 | v_161;
assign x_164 = ~v_873 | v_67;
assign x_165 = ~v_874 | v_160;
assign x_166 = ~v_874 | ~v_161;
assign x_167 = ~v_875 | v_65;
assign x_168 = ~v_875 | ~v_161;
assign x_169 = ~v_876 | v_160;
assign x_170 = ~v_876 | v_65;
assign x_171 = ~v_877 | v_159;
assign x_172 = ~v_877 | ~v_160;
assign x_173 = ~v_878 | v_62;
assign x_174 = ~v_878 | ~v_160;
assign x_175 = ~v_879 | v_159;
assign x_176 = ~v_879 | v_62;
assign x_177 = ~v_880 | v_53;
assign x_178 = ~v_880 | ~v_159;
assign x_179 = ~v_881 | v_58;
assign x_180 = ~v_881 | ~v_159;
assign x_181 = ~v_882 | v_53;
assign x_182 = ~v_882 | v_58;
assign x_183 = ~v_883 | v_157;
assign x_184 = ~v_883 | ~v_158;
assign x_185 = ~v_884 | v_69;
assign x_186 = ~v_884 | ~v_158;
assign x_187 = ~v_885 | v_157;
assign x_188 = ~v_885 | v_69;
assign x_189 = ~v_886 | v_156;
assign x_190 = ~v_886 | ~v_157;
assign x_191 = ~v_887 | v_68;
assign x_192 = ~v_887 | ~v_157;
assign x_193 = ~v_888 | v_156;
assign x_194 = ~v_888 | v_68;
assign x_195 = ~v_889 | v_155;
assign x_196 = ~v_889 | ~v_156;
assign x_197 = ~v_890 | v_66;
assign x_198 = ~v_890 | ~v_156;
assign x_199 = ~v_891 | v_155;
assign x_200 = ~v_891 | v_66;
assign x_201 = ~v_892 | v_154;
assign x_202 = ~v_892 | ~v_155;
assign x_203 = ~v_893 | v_63;
assign x_204 = ~v_893 | ~v_155;
assign x_205 = ~v_894 | v_154;
assign x_206 = ~v_894 | v_63;
assign x_207 = ~v_895 | v_54;
assign x_208 = ~v_895 | ~v_154;
assign x_209 = ~v_896 | v_59;
assign x_210 = ~v_896 | ~v_154;
assign x_211 = ~v_897 | v_54;
assign x_212 = ~v_897 | v_59;
assign x_213 = ~v_898 | v_212;
assign x_214 = ~v_898 | ~v_213;
assign x_215 = ~v_899 | v_49;
assign x_216 = ~v_899 | ~v_213;
assign x_217 = ~v_900 | v_212;
assign x_218 = ~v_900 | v_49;
assign x_219 = ~v_901 | v_211;
assign x_220 = ~v_901 | ~v_212;
assign x_221 = ~v_902 | v_50;
assign x_222 = ~v_902 | ~v_212;
assign x_223 = ~v_903 | v_211;
assign x_224 = ~v_903 | v_50;
assign x_225 = ~v_904 | v_210;
assign x_226 = ~v_904 | ~v_211;
assign x_227 = ~v_905 | v_51;
assign x_228 = ~v_905 | ~v_211;
assign x_229 = ~v_906 | v_210;
assign x_230 = ~v_906 | v_51;
assign x_231 = ~v_907 | v_209;
assign x_232 = ~v_907 | ~v_210;
assign x_233 = ~v_908 | v_52;
assign x_234 = ~v_908 | ~v_210;
assign x_235 = ~v_909 | v_209;
assign x_236 = ~v_909 | v_52;
assign x_237 = ~v_910 | v_54;
assign x_238 = ~v_910 | ~v_209;
assign x_239 = ~v_911 | v_53;
assign x_240 = ~v_911 | ~v_209;
assign x_241 = ~v_912 | v_54;
assign x_242 = ~v_912 | v_53;
assign x_243 = ~v_913 | v_208;
assign x_244 = ~v_913 | v_49;
assign x_245 = ~v_914 | v_207;
assign x_246 = ~v_914 | ~v_208;
assign x_247 = ~v_915 | v_55;
assign x_248 = ~v_915 | ~v_208;
assign x_249 = ~v_916 | v_207;
assign x_250 = ~v_916 | v_55;
assign x_251 = ~v_917 | v_206;
assign x_252 = ~v_917 | ~v_207;
assign x_253 = ~v_918 | v_56;
assign x_254 = ~v_918 | ~v_207;
assign x_255 = ~v_919 | v_206;
assign x_256 = ~v_919 | v_56;
assign x_257 = ~v_920 | v_205;
assign x_258 = ~v_920 | ~v_206;
assign x_259 = ~v_921 | v_57;
assign x_260 = ~v_921 | ~v_206;
assign x_261 = ~v_922 | v_205;
assign x_262 = ~v_922 | v_57;
assign x_263 = ~v_923 | v_59;
assign x_264 = ~v_923 | ~v_205;
assign x_265 = ~v_924 | v_58;
assign x_266 = ~v_924 | ~v_205;
assign x_267 = ~v_925 | v_59;
assign x_268 = ~v_925 | v_58;
assign x_269 = ~v_926 | v_204;
assign x_270 = ~v_926 | v_50;
assign x_271 = ~v_927 | v_204;
assign x_272 = ~v_927 | v_55;
assign x_273 = ~v_928 | v_203;
assign x_274 = ~v_928 | ~v_204;
assign x_275 = ~v_929 | v_60;
assign x_276 = ~v_929 | ~v_204;
assign x_277 = ~v_930 | v_203;
assign x_278 = ~v_930 | v_60;
assign x_279 = ~v_931 | v_202;
assign x_280 = ~v_931 | ~v_203;
assign x_281 = ~v_932 | v_61;
assign x_282 = ~v_932 | ~v_203;
assign x_283 = ~v_933 | v_202;
assign x_284 = ~v_933 | v_61;
assign x_285 = ~v_934 | v_63;
assign x_286 = ~v_934 | ~v_202;
assign x_287 = ~v_935 | v_62;
assign x_288 = ~v_935 | ~v_202;
assign x_289 = ~v_936 | v_63;
assign x_290 = ~v_936 | v_62;
assign x_291 = ~v_937 | v_55;
assign x_292 = ~v_937 | ~v_201;
assign x_293 = ~v_938 | v_50;
assign x_294 = ~v_938 | ~v_201;
assign x_295 = ~v_939 | v_55;
assign x_296 = ~v_939 | v_50;
assign x_297 = ~v_940 | v_200;
assign x_298 = ~v_940 | v_51;
assign x_299 = ~v_941 | v_200;
assign x_300 = ~v_941 | v_56;
assign x_301 = ~v_942 | v_200;
assign x_302 = ~v_942 | v_60;
assign x_303 = ~v_943 | v_199;
assign x_304 = ~v_943 | ~v_200;
assign x_305 = ~v_944 | v_64;
assign x_306 = ~v_944 | ~v_200;
assign x_307 = ~v_945 | v_199;
assign x_308 = ~v_945 | v_64;
assign x_309 = ~v_946 | v_66;
assign x_310 = ~v_946 | ~v_199;
assign x_311 = ~v_947 | v_65;
assign x_312 = ~v_947 | ~v_199;
assign x_313 = ~v_948 | v_66;
assign x_314 = ~v_948 | v_65;
assign x_315 = ~v_949 | v_197;
assign x_316 = ~v_949 | ~v_198;
assign x_317 = ~v_950 | v_51;
assign x_318 = ~v_950 | ~v_198;
assign x_319 = ~v_951 | v_197;
assign x_320 = ~v_951 | v_51;
assign x_321 = ~v_952 | v_60;
assign x_322 = ~v_952 | ~v_197;
assign x_323 = ~v_953 | v_56;
assign x_324 = ~v_953 | ~v_197;
assign x_325 = ~v_954 | v_60;
assign x_326 = ~v_954 | v_56;
assign x_327 = ~v_955 | v_196;
assign x_328 = ~v_955 | v_52;
assign x_329 = ~v_956 | v_196;
assign x_330 = ~v_956 | v_57;
assign x_331 = ~v_957 | v_196;
assign x_332 = ~v_957 | v_61;
assign x_333 = ~v_958 | v_196;
assign x_334 = ~v_958 | v_64;
assign x_335 = ~v_959 | v_68;
assign x_336 = ~v_959 | ~v_196;
assign x_337 = ~v_960 | v_67;
assign x_338 = ~v_960 | ~v_196;
assign x_339 = ~v_961 | v_68;
assign x_340 = ~v_961 | v_67;
assign x_341 = ~v_962 | v_194;
assign x_342 = ~v_962 | ~v_195;
assign x_343 = ~v_963 | v_52;
assign x_344 = ~v_963 | ~v_195;
assign x_345 = ~v_964 | v_194;
assign x_346 = ~v_964 | v_52;
assign x_347 = ~v_965 | v_193;
assign x_348 = ~v_965 | ~v_194;
assign x_349 = ~v_966 | v_57;
assign x_350 = ~v_966 | ~v_194;
assign x_351 = ~v_967 | v_193;
assign x_352 = ~v_967 | v_57;
assign x_353 = ~v_968 | v_64;
assign x_354 = ~v_968 | ~v_193;
assign x_355 = ~v_969 | v_61;
assign x_356 = ~v_969 | ~v_193;
assign x_357 = ~v_970 | v_64;
assign x_358 = ~v_970 | v_61;
assign x_359 = ~v_971 | v_69;
assign x_360 = ~v_971 | v_53;
assign x_361 = ~v_972 | v_69;
assign x_362 = ~v_972 | v_58;
assign x_363 = ~v_973 | v_69;
assign x_364 = ~v_973 | v_62;
assign x_365 = ~v_974 | v_69;
assign x_366 = ~v_974 | v_65;
assign x_367 = ~v_975 | v_69;
assign x_368 = ~v_975 | v_67;
assign x_369 = ~v_976 | v_191;
assign x_370 = ~v_976 | ~v_192;
assign x_371 = ~v_977 | v_53;
assign x_372 = ~v_977 | ~v_192;
assign x_373 = ~v_978 | v_191;
assign x_374 = ~v_978 | v_53;
assign x_375 = ~v_979 | v_190;
assign x_376 = ~v_979 | ~v_191;
assign x_377 = ~v_980 | v_58;
assign x_378 = ~v_980 | ~v_191;
assign x_379 = ~v_981 | v_190;
assign x_380 = ~v_981 | v_58;
assign x_381 = ~v_982 | v_189;
assign x_382 = ~v_982 | ~v_190;
assign x_383 = ~v_983 | v_62;
assign x_384 = ~v_983 | ~v_190;
assign x_385 = ~v_984 | v_189;
assign x_386 = ~v_984 | v_62;
assign x_387 = ~v_985 | v_67;
assign x_388 = ~v_985 | ~v_189;
assign x_389 = ~v_986 | v_65;
assign x_390 = ~v_986 | ~v_189;
assign x_391 = ~v_987 | v_67;
assign x_392 = ~v_987 | v_65;
assign x_393 = ~v_988 | v_187;
assign x_394 = ~v_988 | ~v_188;
assign x_395 = ~v_989 | v_54;
assign x_396 = ~v_989 | ~v_188;
assign x_397 = ~v_990 | v_187;
assign x_398 = ~v_990 | v_54;
assign x_399 = ~v_991 | v_186;
assign x_400 = ~v_991 | ~v_187;
assign x_401 = ~v_992 | v_59;
assign x_402 = ~v_992 | ~v_187;
assign x_403 = ~v_993 | v_186;
assign x_404 = ~v_993 | v_59;
assign x_405 = ~v_994 | v_185;
assign x_406 = ~v_994 | ~v_186;
assign x_407 = ~v_995 | v_63;
assign x_408 = ~v_995 | ~v_186;
assign x_409 = ~v_996 | v_185;
assign x_410 = ~v_996 | v_63;
assign x_411 = ~v_997 | v_184;
assign x_412 = ~v_997 | ~v_185;
assign x_413 = ~v_998 | v_66;
assign x_414 = ~v_998 | ~v_185;
assign x_415 = ~v_999 | v_184;
assign x_416 = ~v_999 | v_66;
assign x_417 = ~v_1000 | v_69;
assign x_418 = ~v_1000 | ~v_184;
assign x_419 = ~v_1001 | v_68;
assign x_420 = ~v_1001 | ~v_184;
assign x_421 = ~v_1002 | v_69;
assign x_422 = ~v_1002 | v_68;
assign x_423 = ~v_1003 | v_1871;
assign x_424 = ~v_1003 | ~v_1872;
assign x_425 = ~v_1004 | v_75;
assign x_426 = ~v_1004 | ~v_1872;
assign x_427 = ~v_1005 | v_1871;
assign x_428 = ~v_1005 | v_75;
assign x_429 = ~v_1006 | v_1870;
assign x_430 = ~v_1006 | ~v_1871;
assign x_431 = ~v_1007 | v_74;
assign x_432 = ~v_1007 | ~v_1871;
assign x_433 = ~v_1008 | v_1870;
assign x_434 = ~v_1008 | v_74;
assign x_435 = ~v_1009 | v_1869;
assign x_436 = ~v_1009 | ~v_1870;
assign x_437 = ~v_1010 | v_73;
assign x_438 = ~v_1010 | ~v_1870;
assign x_439 = ~v_1011 | v_1869;
assign x_440 = ~v_1011 | v_73;
assign x_441 = ~v_1012 | v_1868;
assign x_442 = ~v_1012 | ~v_1869;
assign x_443 = ~v_1013 | v_72;
assign x_444 = ~v_1013 | ~v_1869;
assign x_445 = ~v_1014 | v_1868;
assign x_446 = ~v_1014 | v_72;
assign x_447 = ~v_1015 | v_70;
assign x_448 = ~v_1015 | ~v_1868;
assign x_449 = ~v_1016 | v_71;
assign x_450 = ~v_1016 | ~v_1868;
assign x_451 = ~v_1017 | v_70;
assign x_452 = ~v_1017 | v_71;
assign x_453 = ~v_1018 | v_1866;
assign x_454 = ~v_1018 | ~v_1867;
assign x_455 = ~v_1019 | v_80;
assign x_456 = ~v_1019 | ~v_1867;
assign x_457 = ~v_1020 | v_1866;
assign x_458 = ~v_1020 | v_80;
assign x_459 = ~v_1021 | v_1865;
assign x_460 = ~v_1021 | ~v_1866;
assign x_461 = ~v_1022 | v_79;
assign x_462 = ~v_1022 | ~v_1866;
assign x_463 = ~v_1023 | v_1865;
assign x_464 = ~v_1023 | v_79;
assign x_465 = ~v_1024 | v_1864;
assign x_466 = ~v_1024 | ~v_1865;
assign x_467 = ~v_1025 | v_78;
assign x_468 = ~v_1025 | ~v_1865;
assign x_469 = ~v_1026 | v_1864;
assign x_470 = ~v_1026 | v_78;
assign x_471 = ~v_1027 | v_76;
assign x_472 = ~v_1027 | ~v_1864;
assign x_473 = ~v_1028 | v_77;
assign x_474 = ~v_1028 | ~v_1864;
assign x_475 = ~v_1029 | v_76;
assign x_476 = ~v_1029 | v_77;
assign x_477 = ~v_1030 | v_70;
assign x_478 = ~v_1030 | v_80;
assign x_479 = ~v_1031 | v_70;
assign x_480 = ~v_1031 | v_79;
assign x_481 = ~v_1032 | v_70;
assign x_482 = ~v_1032 | v_78;
assign x_483 = ~v_1033 | v_70;
assign x_484 = ~v_1033 | v_77;
assign x_485 = ~v_1034 | v_70;
assign x_486 = ~v_1034 | v_76;
assign x_487 = ~v_1035 | v_1862;
assign x_488 = ~v_1035 | ~v_1863;
assign x_489 = ~v_1036 | v_84;
assign x_490 = ~v_1036 | ~v_1863;
assign x_491 = ~v_1037 | v_1862;
assign x_492 = ~v_1037 | v_84;
assign x_493 = ~v_1038 | v_1861;
assign x_494 = ~v_1038 | ~v_1862;
assign x_495 = ~v_1039 | v_83;
assign x_496 = ~v_1039 | ~v_1862;
assign x_497 = ~v_1040 | v_1861;
assign x_498 = ~v_1040 | v_83;
assign x_499 = ~v_1041 | v_81;
assign x_500 = ~v_1041 | ~v_1861;
assign x_501 = ~v_1042 | v_82;
assign x_502 = ~v_1042 | ~v_1861;
assign x_503 = ~v_1043 | v_81;
assign x_504 = ~v_1043 | v_82;
assign x_505 = ~v_1044 | v_1860;
assign x_506 = ~v_1044 | v_84;
assign x_507 = ~v_1045 | v_1860;
assign x_508 = ~v_1045 | v_83;
assign x_509 = ~v_1046 | v_1860;
assign x_510 = ~v_1046 | v_82;
assign x_511 = ~v_1047 | v_1860;
assign x_512 = ~v_1047 | v_81;
assign x_513 = ~v_1048 | v_71;
assign x_514 = ~v_1048 | ~v_1860;
assign x_515 = ~v_1049 | v_76;
assign x_516 = ~v_1049 | ~v_1860;
assign x_517 = ~v_1050 | v_71;
assign x_518 = ~v_1050 | v_76;
assign x_519 = ~v_1051 | v_1858;
assign x_520 = ~v_1051 | ~v_1859;
assign x_521 = ~v_1052 | v_87;
assign x_522 = ~v_1052 | ~v_1859;
assign x_523 = ~v_1053 | v_1858;
assign x_524 = ~v_1053 | v_87;
assign x_525 = ~v_1054 | v_85;
assign x_526 = ~v_1054 | ~v_1858;
assign x_527 = ~v_1055 | v_86;
assign x_528 = ~v_1055 | ~v_1858;
assign x_529 = ~v_1056 | v_85;
assign x_530 = ~v_1056 | v_86;
assign x_531 = ~v_1057 | v_1857;
assign x_532 = ~v_1057 | v_87;
assign x_533 = ~v_1058 | v_1857;
assign x_534 = ~v_1058 | v_86;
assign x_535 = ~v_1059 | v_1857;
assign x_536 = ~v_1059 | v_85;
assign x_537 = ~v_1060 | v_1856;
assign x_538 = ~v_1060 | ~v_1857;
assign x_539 = ~v_1061 | v_81;
assign x_540 = ~v_1061 | ~v_1857;
assign x_541 = ~v_1062 | v_1856;
assign x_542 = ~v_1062 | v_81;
assign x_543 = ~v_1063 | v_72;
assign x_544 = ~v_1063 | ~v_1856;
assign x_545 = ~v_1064 | v_77;
assign x_546 = ~v_1064 | ~v_1856;
assign x_547 = ~v_1065 | v_72;
assign x_548 = ~v_1065 | v_77;
assign x_549 = ~v_1066 | v_88;
assign x_550 = ~v_1066 | ~v_1855;
assign x_551 = ~v_1067 | v_89;
assign x_552 = ~v_1067 | ~v_1855;
assign x_553 = ~v_1068 | v_88;
assign x_554 = ~v_1068 | v_89;
assign x_555 = ~v_1069 | v_1854;
assign x_556 = ~v_1069 | v_89;
assign x_557 = ~v_1070 | v_1854;
assign x_558 = ~v_1070 | v_88;
assign x_559 = ~v_1071 | v_1853;
assign x_560 = ~v_1071 | ~v_1854;
assign x_561 = ~v_1072 | v_85;
assign x_562 = ~v_1072 | ~v_1854;
assign x_563 = ~v_1073 | v_1853;
assign x_564 = ~v_1073 | v_85;
assign x_565 = ~v_1074 | v_1852;
assign x_566 = ~v_1074 | ~v_1853;
assign x_567 = ~v_1075 | v_82;
assign x_568 = ~v_1075 | ~v_1853;
assign x_569 = ~v_1076 | v_1852;
assign x_570 = ~v_1076 | v_82;
assign x_571 = ~v_1077 | v_73;
assign x_572 = ~v_1077 | ~v_1852;
assign x_573 = ~v_1078 | v_78;
assign x_574 = ~v_1078 | ~v_1852;
assign x_575 = ~v_1079 | v_73;
assign x_576 = ~v_1079 | v_78;
assign x_577 = ~v_1080 | v_1851;
assign x_578 = ~v_1080 | v_90;
assign x_579 = ~v_1081 | v_1850;
assign x_580 = ~v_1081 | ~v_1851;
assign x_581 = ~v_1082 | v_88;
assign x_582 = ~v_1082 | ~v_1851;
assign x_583 = ~v_1083 | v_1850;
assign x_584 = ~v_1083 | v_88;
assign x_585 = ~v_1084 | v_1849;
assign x_586 = ~v_1084 | ~v_1850;
assign x_587 = ~v_1085 | v_86;
assign x_588 = ~v_1085 | ~v_1850;
assign x_589 = ~v_1086 | v_1849;
assign x_590 = ~v_1086 | v_86;
assign x_591 = ~v_1087 | v_1848;
assign x_592 = ~v_1087 | ~v_1849;
assign x_593 = ~v_1088 | v_83;
assign x_594 = ~v_1088 | ~v_1849;
assign x_595 = ~v_1089 | v_1848;
assign x_596 = ~v_1089 | v_83;
assign x_597 = ~v_1090 | v_74;
assign x_598 = ~v_1090 | ~v_1848;
assign x_599 = ~v_1091 | v_79;
assign x_600 = ~v_1091 | ~v_1848;
assign x_601 = ~v_1092 | v_74;
assign x_602 = ~v_1092 | v_79;
assign x_603 = ~v_1093 | v_1846;
assign x_604 = ~v_1093 | ~v_1847;
assign x_605 = ~v_1094 | v_90;
assign x_606 = ~v_1094 | ~v_1847;
assign x_607 = ~v_1095 | v_1846;
assign x_608 = ~v_1095 | v_90;
assign x_609 = ~v_1096 | v_1845;
assign x_610 = ~v_1096 | ~v_1846;
assign x_611 = ~v_1097 | v_89;
assign x_612 = ~v_1097 | ~v_1846;
assign x_613 = ~v_1098 | v_1845;
assign x_614 = ~v_1098 | v_89;
assign x_615 = ~v_1099 | v_1844;
assign x_616 = ~v_1099 | ~v_1845;
assign x_617 = ~v_1100 | v_87;
assign x_618 = ~v_1100 | ~v_1845;
assign x_619 = ~v_1101 | v_1844;
assign x_620 = ~v_1101 | v_87;
assign x_621 = ~v_1102 | v_1843;
assign x_622 = ~v_1102 | ~v_1844;
assign x_623 = ~v_1103 | v_84;
assign x_624 = ~v_1103 | ~v_1844;
assign x_625 = ~v_1104 | v_1843;
assign x_626 = ~v_1104 | v_84;
assign x_627 = ~v_1105 | v_75;
assign x_628 = ~v_1105 | ~v_1843;
assign x_629 = ~v_1106 | v_80;
assign x_630 = ~v_1106 | ~v_1843;
assign x_631 = ~v_1107 | v_75;
assign x_632 = ~v_1107 | v_80;
assign x_633 = ~v_1108 | v_1901;
assign x_634 = ~v_1108 | ~v_1902;
assign x_635 = ~v_1109 | v_70;
assign x_636 = ~v_1109 | ~v_1902;
assign x_637 = ~v_1110 | v_1901;
assign x_638 = ~v_1110 | v_70;
assign x_639 = ~v_1111 | v_1900;
assign x_640 = ~v_1111 | ~v_1901;
assign x_641 = ~v_1112 | v_71;
assign x_642 = ~v_1112 | ~v_1901;
assign x_643 = ~v_1113 | v_1900;
assign x_644 = ~v_1113 | v_71;
assign x_645 = ~v_1114 | v_1899;
assign x_646 = ~v_1114 | ~v_1900;
assign x_647 = ~v_1115 | v_72;
assign x_648 = ~v_1115 | ~v_1900;
assign x_649 = ~v_1116 | v_1899;
assign x_650 = ~v_1116 | v_72;
assign x_651 = ~v_1117 | v_1898;
assign x_652 = ~v_1117 | ~v_1899;
assign x_653 = ~v_1118 | v_73;
assign x_654 = ~v_1118 | ~v_1899;
assign x_655 = ~v_1119 | v_1898;
assign x_656 = ~v_1119 | v_73;
assign x_657 = ~v_1120 | v_75;
assign x_658 = ~v_1120 | ~v_1898;
assign x_659 = ~v_1121 | v_74;
assign x_660 = ~v_1121 | ~v_1898;
assign x_661 = ~v_1122 | v_75;
assign x_662 = ~v_1122 | v_74;
assign x_663 = ~v_1123 | v_1897;
assign x_664 = ~v_1123 | v_70;
assign x_665 = ~v_1124 | v_1896;
assign x_666 = ~v_1124 | ~v_1897;
assign x_667 = ~v_1125 | v_76;
assign x_668 = ~v_1125 | ~v_1897;
assign x_669 = ~v_1126 | v_1896;
assign x_670 = ~v_1126 | v_76;
assign x_671 = ~v_1127 | v_1895;
assign x_672 = ~v_1127 | ~v_1896;
assign x_673 = ~v_1128 | v_77;
assign x_674 = ~v_1128 | ~v_1896;
assign x_675 = ~v_1129 | v_1895;
assign x_676 = ~v_1129 | v_77;
assign x_677 = ~v_1130 | v_1894;
assign x_678 = ~v_1130 | ~v_1895;
assign x_679 = ~v_1131 | v_78;
assign x_680 = ~v_1131 | ~v_1895;
assign x_681 = ~v_1132 | v_1894;
assign x_682 = ~v_1132 | v_78;
assign x_683 = ~v_1133 | v_80;
assign x_684 = ~v_1133 | ~v_1894;
assign x_685 = ~v_1134 | v_79;
assign x_686 = ~v_1134 | ~v_1894;
assign x_687 = ~v_1135 | v_80;
assign x_688 = ~v_1135 | v_79;
assign x_689 = ~v_1136 | v_1893;
assign x_690 = ~v_1136 | v_71;
assign x_691 = ~v_1137 | v_1893;
assign x_692 = ~v_1137 | v_76;
assign x_693 = ~v_1138 | v_1892;
assign x_694 = ~v_1138 | ~v_1893;
assign x_695 = ~v_1139 | v_81;
assign x_696 = ~v_1139 | ~v_1893;
assign x_697 = ~v_1140 | v_1892;
assign x_698 = ~v_1140 | v_81;
assign x_699 = ~v_1141 | v_1891;
assign x_700 = ~v_1141 | ~v_1892;
assign x_701 = ~v_1142 | v_82;
assign x_702 = ~v_1142 | ~v_1892;
assign x_703 = ~v_1143 | v_1891;
assign x_704 = ~v_1143 | v_82;
assign x_705 = ~v_1144 | v_84;
assign x_706 = ~v_1144 | ~v_1891;
assign x_707 = ~v_1145 | v_83;
assign x_708 = ~v_1145 | ~v_1891;
assign x_709 = ~v_1146 | v_84;
assign x_710 = ~v_1146 | v_83;
assign x_711 = ~v_1147 | v_76;
assign x_712 = ~v_1147 | ~v_1890;
assign x_713 = ~v_1148 | v_71;
assign x_714 = ~v_1148 | ~v_1890;
assign x_715 = ~v_1149 | v_76;
assign x_716 = ~v_1149 | v_71;
assign x_717 = ~v_1150 | v_1889;
assign x_718 = ~v_1150 | v_72;
assign x_719 = ~v_1151 | v_1889;
assign x_720 = ~v_1151 | v_77;
assign x_721 = ~v_1152 | v_1889;
assign x_722 = ~v_1152 | v_81;
assign x_723 = ~v_1153 | v_1888;
assign x_724 = ~v_1153 | ~v_1889;
assign x_725 = ~v_1154 | v_85;
assign x_726 = ~v_1154 | ~v_1889;
assign x_727 = ~v_1155 | v_1888;
assign x_728 = ~v_1155 | v_85;
assign x_729 = ~v_1156 | v_87;
assign x_730 = ~v_1156 | ~v_1888;
assign x_731 = ~v_1157 | v_86;
assign x_732 = ~v_1157 | ~v_1888;
assign x_733 = ~v_1158 | v_87;
assign x_734 = ~v_1158 | v_86;
assign x_735 = ~v_1159 | v_1886;
assign x_736 = ~v_1159 | ~v_1887;
assign x_737 = ~v_1160 | v_72;
assign x_738 = ~v_1160 | ~v_1887;
assign x_739 = ~v_1161 | v_1886;
assign x_740 = ~v_1161 | v_72;
assign x_741 = ~v_1162 | v_81;
assign x_742 = ~v_1162 | ~v_1886;
assign x_743 = ~v_1163 | v_77;
assign x_744 = ~v_1163 | ~v_1886;
assign x_745 = ~v_1164 | v_81;
assign x_746 = ~v_1164 | v_77;
assign x_747 = ~v_1165 | v_1885;
assign x_748 = ~v_1165 | v_73;
assign x_749 = ~v_1166 | v_1885;
assign x_750 = ~v_1166 | v_78;
assign x_751 = ~v_1167 | v_1885;
assign x_752 = ~v_1167 | v_82;
assign x_753 = ~v_1168 | v_1885;
assign x_754 = ~v_1168 | v_85;
assign x_755 = ~v_1169 | v_89;
assign x_756 = ~v_1169 | ~v_1885;
assign x_757 = ~v_1170 | v_88;
assign x_758 = ~v_1170 | ~v_1885;
assign x_759 = ~v_1171 | v_89;
assign x_760 = ~v_1171 | v_88;
assign x_761 = ~v_1172 | v_1883;
assign x_762 = ~v_1172 | ~v_1884;
assign x_763 = ~v_1173 | v_73;
assign x_764 = ~v_1173 | ~v_1884;
assign x_765 = ~v_1174 | v_1883;
assign x_766 = ~v_1174 | v_73;
assign x_767 = ~v_1175 | v_1882;
assign x_768 = ~v_1175 | ~v_1883;
assign x_769 = ~v_1176 | v_78;
assign x_770 = ~v_1176 | ~v_1883;
assign x_771 = ~v_1177 | v_1882;
assign x_772 = ~v_1177 | v_78;
assign x_773 = ~v_1178 | v_85;
assign x_774 = ~v_1178 | ~v_1882;
assign x_775 = ~v_1179 | v_82;
assign x_776 = ~v_1179 | ~v_1882;
assign x_777 = ~v_1180 | v_85;
assign x_778 = ~v_1180 | v_82;
assign x_779 = ~v_1181 | v_90;
assign x_780 = ~v_1181 | v_74;
assign x_781 = ~v_1182 | v_90;
assign x_782 = ~v_1182 | v_79;
assign x_783 = ~v_1183 | v_90;
assign x_784 = ~v_1183 | v_83;
assign x_785 = ~v_1184 | v_90;
assign x_786 = ~v_1184 | v_86;
assign x_787 = ~v_1185 | v_90;
assign x_788 = ~v_1185 | v_88;
assign x_789 = ~v_1186 | v_1880;
assign x_790 = ~v_1186 | ~v_1881;
assign x_791 = ~v_1187 | v_74;
assign x_792 = ~v_1187 | ~v_1881;
assign x_793 = ~v_1188 | v_1880;
assign x_794 = ~v_1188 | v_74;
assign x_795 = ~v_1189 | v_1879;
assign x_796 = ~v_1189 | ~v_1880;
assign x_797 = ~v_1190 | v_79;
assign x_798 = ~v_1190 | ~v_1880;
assign x_799 = ~v_1191 | v_1879;
assign x_800 = ~v_1191 | v_79;
assign x_801 = ~v_1192 | v_1878;
assign x_802 = ~v_1192 | ~v_1879;
assign x_803 = ~v_1193 | v_83;
assign x_804 = ~v_1193 | ~v_1879;
assign x_805 = ~v_1194 | v_1878;
assign x_806 = ~v_1194 | v_83;
assign x_807 = ~v_1195 | v_88;
assign x_808 = ~v_1195 | ~v_1878;
assign x_809 = ~v_1196 | v_86;
assign x_810 = ~v_1196 | ~v_1878;
assign x_811 = ~v_1197 | v_88;
assign x_812 = ~v_1197 | v_86;
assign x_813 = ~v_1198 | v_1876;
assign x_814 = ~v_1198 | ~v_1877;
assign x_815 = ~v_1199 | v_75;
assign x_816 = ~v_1199 | ~v_1877;
assign x_817 = ~v_1200 | v_1876;
assign x_818 = ~v_1200 | v_75;
assign x_819 = ~v_1201 | v_1875;
assign x_820 = ~v_1201 | ~v_1876;
assign x_821 = ~v_1202 | v_80;
assign x_822 = ~v_1202 | ~v_1876;
assign x_823 = ~v_1203 | v_1875;
assign x_824 = ~v_1203 | v_80;
assign x_825 = ~v_1204 | v_1874;
assign x_826 = ~v_1204 | ~v_1875;
assign x_827 = ~v_1205 | v_84;
assign x_828 = ~v_1205 | ~v_1875;
assign x_829 = ~v_1206 | v_1874;
assign x_830 = ~v_1206 | v_84;
assign x_831 = ~v_1207 | v_1873;
assign x_832 = ~v_1207 | ~v_1874;
assign x_833 = ~v_1208 | v_87;
assign x_834 = ~v_1208 | ~v_1874;
assign x_835 = ~v_1209 | v_1873;
assign x_836 = ~v_1209 | v_87;
assign x_837 = ~v_1210 | v_90;
assign x_838 = ~v_1210 | ~v_1873;
assign x_839 = ~v_1211 | v_89;
assign x_840 = ~v_1211 | ~v_1873;
assign x_841 = ~v_1212 | v_90;
assign x_842 = ~v_1212 | v_89;
assign x_843 = ~v_1213 | v_1973;
assign x_844 = ~v_1213 | ~v_1974;
assign x_845 = ~v_1214 | v_96;
assign x_846 = ~v_1214 | ~v_1974;
assign x_847 = ~v_1215 | v_1973;
assign x_848 = ~v_1215 | v_96;
assign x_849 = ~v_1216 | v_1972;
assign x_850 = ~v_1216 | ~v_1973;
assign x_851 = ~v_1217 | v_95;
assign x_852 = ~v_1217 | ~v_1973;
assign x_853 = ~v_1218 | v_1972;
assign x_854 = ~v_1218 | v_95;
assign x_855 = ~v_1219 | v_1971;
assign x_856 = ~v_1219 | ~v_1972;
assign x_857 = ~v_1220 | v_94;
assign x_858 = ~v_1220 | ~v_1972;
assign x_859 = ~v_1221 | v_1971;
assign x_860 = ~v_1221 | v_94;
assign x_861 = ~v_1222 | v_1970;
assign x_862 = ~v_1222 | ~v_1971;
assign x_863 = ~v_1223 | v_93;
assign x_864 = ~v_1223 | ~v_1971;
assign x_865 = ~v_1224 | v_1970;
assign x_866 = ~v_1224 | v_93;
assign x_867 = ~v_1225 | v_91;
assign x_868 = ~v_1225 | ~v_1970;
assign x_869 = ~v_1226 | v_92;
assign x_870 = ~v_1226 | ~v_1970;
assign x_871 = ~v_1227 | v_91;
assign x_872 = ~v_1227 | v_92;
assign x_873 = ~v_1228 | v_1968;
assign x_874 = ~v_1228 | ~v_1969;
assign x_875 = ~v_1229 | v_101;
assign x_876 = ~v_1229 | ~v_1969;
assign x_877 = ~v_1230 | v_1968;
assign x_878 = ~v_1230 | v_101;
assign x_879 = ~v_1231 | v_1967;
assign x_880 = ~v_1231 | ~v_1968;
assign x_881 = ~v_1232 | v_100;
assign x_882 = ~v_1232 | ~v_1968;
assign x_883 = ~v_1233 | v_1967;
assign x_884 = ~v_1233 | v_100;
assign x_885 = ~v_1234 | v_1966;
assign x_886 = ~v_1234 | ~v_1967;
assign x_887 = ~v_1235 | v_99;
assign x_888 = ~v_1235 | ~v_1967;
assign x_889 = ~v_1236 | v_1966;
assign x_890 = ~v_1236 | v_99;
assign x_891 = ~v_1237 | v_97;
assign x_892 = ~v_1237 | ~v_1966;
assign x_893 = ~v_1238 | v_98;
assign x_894 = ~v_1238 | ~v_1966;
assign x_895 = ~v_1239 | v_97;
assign x_896 = ~v_1239 | v_98;
assign x_897 = ~v_1240 | v_91;
assign x_898 = ~v_1240 | v_101;
assign x_899 = ~v_1241 | v_91;
assign x_900 = ~v_1241 | v_100;
assign x_901 = ~v_1242 | v_91;
assign x_902 = ~v_1242 | v_99;
assign x_903 = ~v_1243 | v_91;
assign x_904 = ~v_1243 | v_98;
assign x_905 = ~v_1244 | v_91;
assign x_906 = ~v_1244 | v_97;
assign x_907 = ~v_1245 | v_1964;
assign x_908 = ~v_1245 | ~v_1965;
assign x_909 = ~v_1246 | v_105;
assign x_910 = ~v_1246 | ~v_1965;
assign x_911 = ~v_1247 | v_1964;
assign x_912 = ~v_1247 | v_105;
assign x_913 = ~v_1248 | v_1963;
assign x_914 = ~v_1248 | ~v_1964;
assign x_915 = ~v_1249 | v_104;
assign x_916 = ~v_1249 | ~v_1964;
assign x_917 = ~v_1250 | v_1963;
assign x_918 = ~v_1250 | v_104;
assign x_919 = ~v_1251 | v_102;
assign x_920 = ~v_1251 | ~v_1963;
assign x_921 = ~v_1252 | v_103;
assign x_922 = ~v_1252 | ~v_1963;
assign x_923 = ~v_1253 | v_102;
assign x_924 = ~v_1253 | v_103;
assign x_925 = ~v_1254 | v_1962;
assign x_926 = ~v_1254 | v_105;
assign x_927 = ~v_1255 | v_1962;
assign x_928 = ~v_1255 | v_104;
assign x_929 = ~v_1256 | v_1962;
assign x_930 = ~v_1256 | v_103;
assign x_931 = ~v_1257 | v_1962;
assign x_932 = ~v_1257 | v_102;
assign x_933 = ~v_1258 | v_92;
assign x_934 = ~v_1258 | ~v_1962;
assign x_935 = ~v_1259 | v_97;
assign x_936 = ~v_1259 | ~v_1962;
assign x_937 = ~v_1260 | v_92;
assign x_938 = ~v_1260 | v_97;
assign x_939 = ~v_1261 | v_1960;
assign x_940 = ~v_1261 | ~v_1961;
assign x_941 = ~v_1262 | v_108;
assign x_942 = ~v_1262 | ~v_1961;
assign x_943 = ~v_1263 | v_1960;
assign x_944 = ~v_1263 | v_108;
assign x_945 = ~v_1264 | v_106;
assign x_946 = ~v_1264 | ~v_1960;
assign x_947 = ~v_1265 | v_107;
assign x_948 = ~v_1265 | ~v_1960;
assign x_949 = ~v_1266 | v_106;
assign x_950 = ~v_1266 | v_107;
assign x_951 = ~v_1267 | v_1959;
assign x_952 = ~v_1267 | v_108;
assign x_953 = ~v_1268 | v_1959;
assign x_954 = ~v_1268 | v_107;
assign x_955 = ~v_1269 | v_1959;
assign x_956 = ~v_1269 | v_106;
assign x_957 = ~v_1270 | v_1958;
assign x_958 = ~v_1270 | ~v_1959;
assign x_959 = ~v_1271 | v_102;
assign x_960 = ~v_1271 | ~v_1959;
assign x_961 = ~v_1272 | v_1958;
assign x_962 = ~v_1272 | v_102;
assign x_963 = ~v_1273 | v_93;
assign x_964 = ~v_1273 | ~v_1958;
assign x_965 = ~v_1274 | v_98;
assign x_966 = ~v_1274 | ~v_1958;
assign x_967 = ~v_1275 | v_93;
assign x_968 = ~v_1275 | v_98;
assign x_969 = ~v_1276 | v_109;
assign x_970 = ~v_1276 | ~v_1957;
assign x_971 = ~v_1277 | v_110;
assign x_972 = ~v_1277 | ~v_1957;
assign x_973 = ~v_1278 | v_109;
assign x_974 = ~v_1278 | v_110;
assign x_975 = ~v_1279 | v_1956;
assign x_976 = ~v_1279 | v_110;
assign x_977 = ~v_1280 | v_1956;
assign x_978 = ~v_1280 | v_109;
assign x_979 = ~v_1281 | v_1955;
assign x_980 = ~v_1281 | ~v_1956;
assign x_981 = ~v_1282 | v_106;
assign x_982 = ~v_1282 | ~v_1956;
assign x_983 = ~v_1283 | v_1955;
assign x_984 = ~v_1283 | v_106;
assign x_985 = ~v_1284 | v_1954;
assign x_986 = ~v_1284 | ~v_1955;
assign x_987 = ~v_1285 | v_103;
assign x_988 = ~v_1285 | ~v_1955;
assign x_989 = ~v_1286 | v_1954;
assign x_990 = ~v_1286 | v_103;
assign x_991 = ~v_1287 | v_94;
assign x_992 = ~v_1287 | ~v_1954;
assign x_993 = ~v_1288 | v_99;
assign x_994 = ~v_1288 | ~v_1954;
assign x_995 = ~v_1289 | v_94;
assign x_996 = ~v_1289 | v_99;
assign x_997 = ~v_1290 | v_1953;
assign x_998 = ~v_1290 | v_111;
assign x_999 = ~v_1291 | v_1952;
assign x_1000 = ~v_1291 | ~v_1953;
assign x_1001 = ~v_1292 | v_109;
assign x_1002 = ~v_1292 | ~v_1953;
assign x_1003 = ~v_1293 | v_1952;
assign x_1004 = ~v_1293 | v_109;
assign x_1005 = ~v_1294 | v_1951;
assign x_1006 = ~v_1294 | ~v_1952;
assign x_1007 = ~v_1295 | v_107;
assign x_1008 = ~v_1295 | ~v_1952;
assign x_1009 = ~v_1296 | v_1951;
assign x_1010 = ~v_1296 | v_107;
assign x_1011 = ~v_1297 | v_1950;
assign x_1012 = ~v_1297 | ~v_1951;
assign x_1013 = ~v_1298 | v_104;
assign x_1014 = ~v_1298 | ~v_1951;
assign x_1015 = ~v_1299 | v_1950;
assign x_1016 = ~v_1299 | v_104;
assign x_1017 = ~v_1300 | v_95;
assign x_1018 = ~v_1300 | ~v_1950;
assign x_1019 = ~v_1301 | v_100;
assign x_1020 = ~v_1301 | ~v_1950;
assign x_1021 = ~v_1302 | v_95;
assign x_1022 = ~v_1302 | v_100;
assign x_1023 = ~v_1303 | v_1948;
assign x_1024 = ~v_1303 | ~v_1949;
assign x_1025 = ~v_1304 | v_111;
assign x_1026 = ~v_1304 | ~v_1949;
assign x_1027 = ~v_1305 | v_1948;
assign x_1028 = ~v_1305 | v_111;
assign x_1029 = ~v_1306 | v_1947;
assign x_1030 = ~v_1306 | ~v_1948;
assign x_1031 = ~v_1307 | v_110;
assign x_1032 = ~v_1307 | ~v_1948;
assign x_1033 = ~v_1308 | v_1947;
assign x_1034 = ~v_1308 | v_110;
assign x_1035 = ~v_1309 | v_1946;
assign x_1036 = ~v_1309 | ~v_1947;
assign x_1037 = ~v_1310 | v_108;
assign x_1038 = ~v_1310 | ~v_1947;
assign x_1039 = ~v_1311 | v_1946;
assign x_1040 = ~v_1311 | v_108;
assign x_1041 = ~v_1312 | v_1945;
assign x_1042 = ~v_1312 | ~v_1946;
assign x_1043 = ~v_1313 | v_105;
assign x_1044 = ~v_1313 | ~v_1946;
assign x_1045 = ~v_1314 | v_1945;
assign x_1046 = ~v_1314 | v_105;
assign x_1047 = ~v_1315 | v_96;
assign x_1048 = ~v_1315 | ~v_1945;
assign x_1049 = ~v_1316 | v_101;
assign x_1050 = ~v_1316 | ~v_1945;
assign x_1051 = ~v_1317 | v_96;
assign x_1052 = ~v_1317 | v_101;
assign x_1053 = ~v_1318 | v_2003;
assign x_1054 = ~v_1318 | ~v_2004;
assign x_1055 = ~v_1319 | v_91;
assign x_1056 = ~v_1319 | ~v_2004;
assign x_1057 = ~v_1320 | v_2003;
assign x_1058 = ~v_1320 | v_91;
assign x_1059 = ~v_1321 | v_2002;
assign x_1060 = ~v_1321 | ~v_2003;
assign x_1061 = ~v_1322 | v_92;
assign x_1062 = ~v_1322 | ~v_2003;
assign x_1063 = ~v_1323 | v_2002;
assign x_1064 = ~v_1323 | v_92;
assign x_1065 = ~v_1324 | v_2001;
assign x_1066 = ~v_1324 | ~v_2002;
assign x_1067 = ~v_1325 | v_93;
assign x_1068 = ~v_1325 | ~v_2002;
assign x_1069 = ~v_1326 | v_2001;
assign x_1070 = ~v_1326 | v_93;
assign x_1071 = ~v_1327 | v_2000;
assign x_1072 = ~v_1327 | ~v_2001;
assign x_1073 = ~v_1328 | v_94;
assign x_1074 = ~v_1328 | ~v_2001;
assign x_1075 = ~v_1329 | v_2000;
assign x_1076 = ~v_1329 | v_94;
assign x_1077 = ~v_1330 | v_96;
assign x_1078 = ~v_1330 | ~v_2000;
assign x_1079 = ~v_1331 | v_95;
assign x_1080 = ~v_1331 | ~v_2000;
assign x_1081 = ~v_1332 | v_96;
assign x_1082 = ~v_1332 | v_95;
assign x_1083 = ~v_1333 | v_1999;
assign x_1084 = ~v_1333 | v_91;
assign x_1085 = ~v_1334 | v_1998;
assign x_1086 = ~v_1334 | ~v_1999;
assign x_1087 = ~v_1335 | v_97;
assign x_1088 = ~v_1335 | ~v_1999;
assign x_1089 = ~v_1336 | v_1998;
assign x_1090 = ~v_1336 | v_97;
assign x_1091 = ~v_1337 | v_1997;
assign x_1092 = ~v_1337 | ~v_1998;
assign x_1093 = ~v_1338 | v_98;
assign x_1094 = ~v_1338 | ~v_1998;
assign x_1095 = ~v_1339 | v_1997;
assign x_1096 = ~v_1339 | v_98;
assign x_1097 = ~v_1340 | v_1996;
assign x_1098 = ~v_1340 | ~v_1997;
assign x_1099 = ~v_1341 | v_99;
assign x_1100 = ~v_1341 | ~v_1997;
assign x_1101 = ~v_1342 | v_1996;
assign x_1102 = ~v_1342 | v_99;
assign x_1103 = ~v_1343 | v_101;
assign x_1104 = ~v_1343 | ~v_1996;
assign x_1105 = ~v_1344 | v_100;
assign x_1106 = ~v_1344 | ~v_1996;
assign x_1107 = ~v_1345 | v_101;
assign x_1108 = ~v_1345 | v_100;
assign x_1109 = ~v_1346 | v_1995;
assign x_1110 = ~v_1346 | v_92;
assign x_1111 = ~v_1347 | v_1995;
assign x_1112 = ~v_1347 | v_97;
assign x_1113 = ~v_1348 | v_1994;
assign x_1114 = ~v_1348 | ~v_1995;
assign x_1115 = ~v_1349 | v_102;
assign x_1116 = ~v_1349 | ~v_1995;
assign x_1117 = ~v_1350 | v_1994;
assign x_1118 = ~v_1350 | v_102;
assign x_1119 = ~v_1351 | v_1993;
assign x_1120 = ~v_1351 | ~v_1994;
assign x_1121 = ~v_1352 | v_103;
assign x_1122 = ~v_1352 | ~v_1994;
assign x_1123 = ~v_1353 | v_1993;
assign x_1124 = ~v_1353 | v_103;
assign x_1125 = ~v_1354 | v_105;
assign x_1126 = ~v_1354 | ~v_1993;
assign x_1127 = ~v_1355 | v_104;
assign x_1128 = ~v_1355 | ~v_1993;
assign x_1129 = ~v_1356 | v_105;
assign x_1130 = ~v_1356 | v_104;
assign x_1131 = ~v_1357 | v_97;
assign x_1132 = ~v_1357 | ~v_1992;
assign x_1133 = ~v_1358 | v_92;
assign x_1134 = ~v_1358 | ~v_1992;
assign x_1135 = ~v_1359 | v_97;
assign x_1136 = ~v_1359 | v_92;
assign x_1137 = ~v_1360 | v_1991;
assign x_1138 = ~v_1360 | v_93;
assign x_1139 = ~v_1361 | v_1991;
assign x_1140 = ~v_1361 | v_98;
assign x_1141 = ~v_1362 | v_1991;
assign x_1142 = ~v_1362 | v_102;
assign x_1143 = ~v_1363 | v_1990;
assign x_1144 = ~v_1363 | ~v_1991;
assign x_1145 = ~v_1364 | v_106;
assign x_1146 = ~v_1364 | ~v_1991;
assign x_1147 = ~v_1365 | v_1990;
assign x_1148 = ~v_1365 | v_106;
assign x_1149 = ~v_1366 | v_108;
assign x_1150 = ~v_1366 | ~v_1990;
assign x_1151 = ~v_1367 | v_107;
assign x_1152 = ~v_1367 | ~v_1990;
assign x_1153 = ~v_1368 | v_108;
assign x_1154 = ~v_1368 | v_107;
assign x_1155 = ~v_1369 | v_1988;
assign x_1156 = ~v_1369 | ~v_1989;
assign x_1157 = ~v_1370 | v_93;
assign x_1158 = ~v_1370 | ~v_1989;
assign x_1159 = ~v_1371 | v_1988;
assign x_1160 = ~v_1371 | v_93;
assign x_1161 = ~v_1372 | v_102;
assign x_1162 = ~v_1372 | ~v_1988;
assign x_1163 = ~v_1373 | v_98;
assign x_1164 = ~v_1373 | ~v_1988;
assign x_1165 = ~v_1374 | v_102;
assign x_1166 = ~v_1374 | v_98;
assign x_1167 = ~v_1375 | v_1987;
assign x_1168 = ~v_1375 | v_94;
assign x_1169 = ~v_1376 | v_1987;
assign x_1170 = ~v_1376 | v_99;
assign x_1171 = ~v_1377 | v_1987;
assign x_1172 = ~v_1377 | v_103;
assign x_1173 = ~v_1378 | v_1987;
assign x_1174 = ~v_1378 | v_106;
assign x_1175 = ~v_1379 | v_110;
assign x_1176 = ~v_1379 | ~v_1987;
assign x_1177 = ~v_1380 | v_109;
assign x_1178 = ~v_1380 | ~v_1987;
assign x_1179 = ~v_1381 | v_110;
assign x_1180 = ~v_1381 | v_109;
assign x_1181 = ~v_1382 | v_1985;
assign x_1182 = ~v_1382 | ~v_1986;
assign x_1183 = ~v_1383 | v_94;
assign x_1184 = ~v_1383 | ~v_1986;
assign x_1185 = ~v_1384 | v_1985;
assign x_1186 = ~v_1384 | v_94;
assign x_1187 = ~v_1385 | v_1984;
assign x_1188 = ~v_1385 | ~v_1985;
assign x_1189 = ~v_1386 | v_99;
assign x_1190 = ~v_1386 | ~v_1985;
assign x_1191 = ~v_1387 | v_1984;
assign x_1192 = ~v_1387 | v_99;
assign x_1193 = ~v_1388 | v_106;
assign x_1194 = ~v_1388 | ~v_1984;
assign x_1195 = ~v_1389 | v_103;
assign x_1196 = ~v_1389 | ~v_1984;
assign x_1197 = ~v_1390 | v_106;
assign x_1198 = ~v_1390 | v_103;
assign x_1199 = ~v_1391 | v_111;
assign x_1200 = ~v_1391 | v_95;
assign x_1201 = ~v_1392 | v_111;
assign x_1202 = ~v_1392 | v_100;
assign x_1203 = ~v_1393 | v_111;
assign x_1204 = ~v_1393 | v_104;
assign x_1205 = ~v_1394 | v_111;
assign x_1206 = ~v_1394 | v_107;
assign x_1207 = ~v_1395 | v_111;
assign x_1208 = ~v_1395 | v_109;
assign x_1209 = ~v_1396 | v_1982;
assign x_1210 = ~v_1396 | ~v_1983;
assign x_1211 = ~v_1397 | v_95;
assign x_1212 = ~v_1397 | ~v_1983;
assign x_1213 = ~v_1398 | v_1982;
assign x_1214 = ~v_1398 | v_95;
assign x_1215 = ~v_1399 | v_1981;
assign x_1216 = ~v_1399 | ~v_1982;
assign x_1217 = ~v_1400 | v_100;
assign x_1218 = ~v_1400 | ~v_1982;
assign x_1219 = ~v_1401 | v_1981;
assign x_1220 = ~v_1401 | v_100;
assign x_1221 = ~v_1402 | v_1980;
assign x_1222 = ~v_1402 | ~v_1981;
assign x_1223 = ~v_1403 | v_104;
assign x_1224 = ~v_1403 | ~v_1981;
assign x_1225 = ~v_1404 | v_1980;
assign x_1226 = ~v_1404 | v_104;
assign x_1227 = ~v_1405 | v_109;
assign x_1228 = ~v_1405 | ~v_1980;
assign x_1229 = ~v_1406 | v_107;
assign x_1230 = ~v_1406 | ~v_1980;
assign x_1231 = ~v_1407 | v_109;
assign x_1232 = ~v_1407 | v_107;
assign x_1233 = ~v_1408 | v_1978;
assign x_1234 = ~v_1408 | ~v_1979;
assign x_1235 = ~v_1409 | v_96;
assign x_1236 = ~v_1409 | ~v_1979;
assign x_1237 = ~v_1410 | v_1978;
assign x_1238 = ~v_1410 | v_96;
assign x_1239 = ~v_1411 | v_1977;
assign x_1240 = ~v_1411 | ~v_1978;
assign x_1241 = ~v_1412 | v_101;
assign x_1242 = ~v_1412 | ~v_1978;
assign x_1243 = ~v_1413 | v_1977;
assign x_1244 = ~v_1413 | v_101;
assign x_1245 = ~v_1414 | v_1976;
assign x_1246 = ~v_1414 | ~v_1977;
assign x_1247 = ~v_1415 | v_105;
assign x_1248 = ~v_1415 | ~v_1977;
assign x_1249 = ~v_1416 | v_1976;
assign x_1250 = ~v_1416 | v_105;
assign x_1251 = ~v_1417 | v_1975;
assign x_1252 = ~v_1417 | ~v_1976;
assign x_1253 = ~v_1418 | v_108;
assign x_1254 = ~v_1418 | ~v_1976;
assign x_1255 = ~v_1419 | v_1975;
assign x_1256 = ~v_1419 | v_108;
assign x_1257 = ~v_1420 | v_111;
assign x_1258 = ~v_1420 | ~v_1975;
assign x_1259 = ~v_1421 | v_110;
assign x_1260 = ~v_1421 | ~v_1975;
assign x_1261 = ~v_1422 | v_111;
assign x_1262 = ~v_1422 | v_110;
assign x_1263 = ~v_1423 | v_2075;
assign x_1264 = ~v_1423 | ~v_2076;
assign x_1265 = ~v_1424 | v_117;
assign x_1266 = ~v_1424 | ~v_2076;
assign x_1267 = ~v_1425 | v_2075;
assign x_1268 = ~v_1425 | v_117;
assign x_1269 = ~v_1426 | v_2074;
assign x_1270 = ~v_1426 | ~v_2075;
assign x_1271 = ~v_1427 | v_116;
assign x_1272 = ~v_1427 | ~v_2075;
assign x_1273 = ~v_1428 | v_2074;
assign x_1274 = ~v_1428 | v_116;
assign x_1275 = ~v_1429 | v_2073;
assign x_1276 = ~v_1429 | ~v_2074;
assign x_1277 = ~v_1430 | v_115;
assign x_1278 = ~v_1430 | ~v_2074;
assign x_1279 = ~v_1431 | v_2073;
assign x_1280 = ~v_1431 | v_115;
assign x_1281 = ~v_1432 | v_2072;
assign x_1282 = ~v_1432 | ~v_2073;
assign x_1283 = ~v_1433 | v_114;
assign x_1284 = ~v_1433 | ~v_2073;
assign x_1285 = ~v_1434 | v_2072;
assign x_1286 = ~v_1434 | v_114;
assign x_1287 = ~v_1435 | v_112;
assign x_1288 = ~v_1435 | ~v_2072;
assign x_1289 = ~v_1436 | v_113;
assign x_1290 = ~v_1436 | ~v_2072;
assign x_1291 = ~v_1437 | v_112;
assign x_1292 = ~v_1437 | v_113;
assign x_1293 = ~v_1438 | v_2070;
assign x_1294 = ~v_1438 | ~v_2071;
assign x_1295 = ~v_1439 | v_122;
assign x_1296 = ~v_1439 | ~v_2071;
assign x_1297 = ~v_1440 | v_2070;
assign x_1298 = ~v_1440 | v_122;
assign x_1299 = ~v_1441 | v_2069;
assign x_1300 = ~v_1441 | ~v_2070;
assign x_1301 = ~v_1442 | v_121;
assign x_1302 = ~v_1442 | ~v_2070;
assign x_1303 = ~v_1443 | v_2069;
assign x_1304 = ~v_1443 | v_121;
assign x_1305 = ~v_1444 | v_2068;
assign x_1306 = ~v_1444 | ~v_2069;
assign x_1307 = ~v_1445 | v_120;
assign x_1308 = ~v_1445 | ~v_2069;
assign x_1309 = ~v_1446 | v_2068;
assign x_1310 = ~v_1446 | v_120;
assign x_1311 = ~v_1447 | v_118;
assign x_1312 = ~v_1447 | ~v_2068;
assign x_1313 = ~v_1448 | v_119;
assign x_1314 = ~v_1448 | ~v_2068;
assign x_1315 = ~v_1449 | v_118;
assign x_1316 = ~v_1449 | v_119;
assign x_1317 = ~v_1450 | v_112;
assign x_1318 = ~v_1450 | v_122;
assign x_1319 = ~v_1451 | v_112;
assign x_1320 = ~v_1451 | v_121;
assign x_1321 = ~v_1452 | v_112;
assign x_1322 = ~v_1452 | v_120;
assign x_1323 = ~v_1453 | v_112;
assign x_1324 = ~v_1453 | v_119;
assign x_1325 = ~v_1454 | v_112;
assign x_1326 = ~v_1454 | v_118;
assign x_1327 = ~v_1455 | v_2066;
assign x_1328 = ~v_1455 | ~v_2067;
assign x_1329 = ~v_1456 | v_126;
assign x_1330 = ~v_1456 | ~v_2067;
assign x_1331 = ~v_1457 | v_2066;
assign x_1332 = ~v_1457 | v_126;
assign x_1333 = ~v_1458 | v_2065;
assign x_1334 = ~v_1458 | ~v_2066;
assign x_1335 = ~v_1459 | v_125;
assign x_1336 = ~v_1459 | ~v_2066;
assign x_1337 = ~v_1460 | v_2065;
assign x_1338 = ~v_1460 | v_125;
assign x_1339 = ~v_1461 | v_123;
assign x_1340 = ~v_1461 | ~v_2065;
assign x_1341 = ~v_1462 | v_124;
assign x_1342 = ~v_1462 | ~v_2065;
assign x_1343 = ~v_1463 | v_123;
assign x_1344 = ~v_1463 | v_124;
assign x_1345 = ~v_1464 | v_2064;
assign x_1346 = ~v_1464 | v_126;
assign x_1347 = ~v_1465 | v_2064;
assign x_1348 = ~v_1465 | v_125;
assign x_1349 = ~v_1466 | v_2064;
assign x_1350 = ~v_1466 | v_124;
assign x_1351 = ~v_1467 | v_2064;
assign x_1352 = ~v_1467 | v_123;
assign x_1353 = ~v_1468 | v_113;
assign x_1354 = ~v_1468 | ~v_2064;
assign x_1355 = ~v_1469 | v_118;
assign x_1356 = ~v_1469 | ~v_2064;
assign x_1357 = ~v_1470 | v_113;
assign x_1358 = ~v_1470 | v_118;
assign x_1359 = ~v_1471 | v_2062;
assign x_1360 = ~v_1471 | ~v_2063;
assign x_1361 = ~v_1472 | v_129;
assign x_1362 = ~v_1472 | ~v_2063;
assign x_1363 = ~v_1473 | v_2062;
assign x_1364 = ~v_1473 | v_129;
assign x_1365 = ~v_1474 | v_127;
assign x_1366 = ~v_1474 | ~v_2062;
assign x_1367 = ~v_1475 | v_128;
assign x_1368 = ~v_1475 | ~v_2062;
assign x_1369 = ~v_1476 | v_127;
assign x_1370 = ~v_1476 | v_128;
assign x_1371 = ~v_1477 | v_2061;
assign x_1372 = ~v_1477 | v_129;
assign x_1373 = ~v_1478 | v_2061;
assign x_1374 = ~v_1478 | v_128;
assign x_1375 = ~v_1479 | v_2061;
assign x_1376 = ~v_1479 | v_127;
assign x_1377 = ~v_1480 | v_2060;
assign x_1378 = ~v_1480 | ~v_2061;
assign x_1379 = ~v_1481 | v_123;
assign x_1380 = ~v_1481 | ~v_2061;
assign x_1381 = ~v_1482 | v_2060;
assign x_1382 = ~v_1482 | v_123;
assign x_1383 = ~v_1483 | v_114;
assign x_1384 = ~v_1483 | ~v_2060;
assign x_1385 = ~v_1484 | v_119;
assign x_1386 = ~v_1484 | ~v_2060;
assign x_1387 = ~v_1485 | v_114;
assign x_1388 = ~v_1485 | v_119;
assign x_1389 = ~v_1486 | v_130;
assign x_1390 = ~v_1486 | ~v_2059;
assign x_1391 = ~v_1487 | v_131;
assign x_1392 = ~v_1487 | ~v_2059;
assign x_1393 = ~v_1488 | v_130;
assign x_1394 = ~v_1488 | v_131;
assign x_1395 = ~v_1489 | v_2058;
assign x_1396 = ~v_1489 | v_131;
assign x_1397 = ~v_1490 | v_2058;
assign x_1398 = ~v_1490 | v_130;
assign x_1399 = ~v_1491 | v_2057;
assign x_1400 = ~v_1491 | ~v_2058;
assign x_1401 = ~v_1492 | v_127;
assign x_1402 = ~v_1492 | ~v_2058;
assign x_1403 = ~v_1493 | v_2057;
assign x_1404 = ~v_1493 | v_127;
assign x_1405 = ~v_1494 | v_2056;
assign x_1406 = ~v_1494 | ~v_2057;
assign x_1407 = ~v_1495 | v_124;
assign x_1408 = ~v_1495 | ~v_2057;
assign x_1409 = ~v_1496 | v_2056;
assign x_1410 = ~v_1496 | v_124;
assign x_1411 = ~v_1497 | v_115;
assign x_1412 = ~v_1497 | ~v_2056;
assign x_1413 = ~v_1498 | v_120;
assign x_1414 = ~v_1498 | ~v_2056;
assign x_1415 = ~v_1499 | v_115;
assign x_1416 = ~v_1499 | v_120;
assign x_1417 = ~v_1500 | v_2055;
assign x_1418 = ~v_1500 | v_132;
assign x_1419 = ~v_1501 | v_2054;
assign x_1420 = ~v_1501 | ~v_2055;
assign x_1421 = ~v_1502 | v_130;
assign x_1422 = ~v_1502 | ~v_2055;
assign x_1423 = ~v_1503 | v_2054;
assign x_1424 = ~v_1503 | v_130;
assign x_1425 = ~v_1504 | v_2053;
assign x_1426 = ~v_1504 | ~v_2054;
assign x_1427 = ~v_1505 | v_128;
assign x_1428 = ~v_1505 | ~v_2054;
assign x_1429 = ~v_1506 | v_2053;
assign x_1430 = ~v_1506 | v_128;
assign x_1431 = ~v_1507 | v_2052;
assign x_1432 = ~v_1507 | ~v_2053;
assign x_1433 = ~v_1508 | v_125;
assign x_1434 = ~v_1508 | ~v_2053;
assign x_1435 = ~v_1509 | v_2052;
assign x_1436 = ~v_1509 | v_125;
assign x_1437 = ~v_1510 | v_116;
assign x_1438 = ~v_1510 | ~v_2052;
assign x_1439 = ~v_1511 | v_121;
assign x_1440 = ~v_1511 | ~v_2052;
assign x_1441 = ~v_1512 | v_116;
assign x_1442 = ~v_1512 | v_121;
assign x_1443 = ~v_1513 | v_2050;
assign x_1444 = ~v_1513 | ~v_2051;
assign x_1445 = ~v_1514 | v_132;
assign x_1446 = ~v_1514 | ~v_2051;
assign x_1447 = ~v_1515 | v_2050;
assign x_1448 = ~v_1515 | v_132;
assign x_1449 = ~v_1516 | v_2049;
assign x_1450 = ~v_1516 | ~v_2050;
assign x_1451 = ~v_1517 | v_131;
assign x_1452 = ~v_1517 | ~v_2050;
assign x_1453 = ~v_1518 | v_2049;
assign x_1454 = ~v_1518 | v_131;
assign x_1455 = ~v_1519 | v_2048;
assign x_1456 = ~v_1519 | ~v_2049;
assign x_1457 = ~v_1520 | v_129;
assign x_1458 = ~v_1520 | ~v_2049;
assign x_1459 = ~v_1521 | v_2048;
assign x_1460 = ~v_1521 | v_129;
assign x_1461 = ~v_1522 | v_2047;
assign x_1462 = ~v_1522 | ~v_2048;
assign x_1463 = ~v_1523 | v_126;
assign x_1464 = ~v_1523 | ~v_2048;
assign x_1465 = ~v_1524 | v_2047;
assign x_1466 = ~v_1524 | v_126;
assign x_1467 = ~v_1525 | v_117;
assign x_1468 = ~v_1525 | ~v_2047;
assign x_1469 = ~v_1526 | v_122;
assign x_1470 = ~v_1526 | ~v_2047;
assign x_1471 = ~v_1527 | v_117;
assign x_1472 = ~v_1527 | v_122;
assign x_1473 = ~v_1528 | v_2105;
assign x_1474 = ~v_1528 | ~v_2106;
assign x_1475 = ~v_1529 | v_112;
assign x_1476 = ~v_1529 | ~v_2106;
assign x_1477 = ~v_1530 | v_2105;
assign x_1478 = ~v_1530 | v_112;
assign x_1479 = ~v_1531 | v_2104;
assign x_1480 = ~v_1531 | ~v_2105;
assign x_1481 = ~v_1532 | v_113;
assign x_1482 = ~v_1532 | ~v_2105;
assign x_1483 = ~v_1533 | v_2104;
assign x_1484 = ~v_1533 | v_113;
assign x_1485 = ~v_1534 | v_2103;
assign x_1486 = ~v_1534 | ~v_2104;
assign x_1487 = ~v_1535 | v_114;
assign x_1488 = ~v_1535 | ~v_2104;
assign x_1489 = ~v_1536 | v_2103;
assign x_1490 = ~v_1536 | v_114;
assign x_1491 = ~v_1537 | v_2102;
assign x_1492 = ~v_1537 | ~v_2103;
assign x_1493 = ~v_1538 | v_115;
assign x_1494 = ~v_1538 | ~v_2103;
assign x_1495 = ~v_1539 | v_2102;
assign x_1496 = ~v_1539 | v_115;
assign x_1497 = ~v_1540 | v_117;
assign x_1498 = ~v_1540 | ~v_2102;
assign x_1499 = ~v_1541 | v_116;
assign x_1500 = ~v_1541 | ~v_2102;
assign x_1501 = ~v_1542 | v_117;
assign x_1502 = ~v_1542 | v_116;
assign x_1503 = ~v_1543 | v_2101;
assign x_1504 = ~v_1543 | v_112;
assign x_1505 = ~v_1544 | v_2100;
assign x_1506 = ~v_1544 | ~v_2101;
assign x_1507 = ~v_1545 | v_118;
assign x_1508 = ~v_1545 | ~v_2101;
assign x_1509 = ~v_1546 | v_2100;
assign x_1510 = ~v_1546 | v_118;
assign x_1511 = ~v_1547 | v_2099;
assign x_1512 = ~v_1547 | ~v_2100;
assign x_1513 = ~v_1548 | v_119;
assign x_1514 = ~v_1548 | ~v_2100;
assign x_1515 = ~v_1549 | v_2099;
assign x_1516 = ~v_1549 | v_119;
assign x_1517 = ~v_1550 | v_2098;
assign x_1518 = ~v_1550 | ~v_2099;
assign x_1519 = ~v_1551 | v_120;
assign x_1520 = ~v_1551 | ~v_2099;
assign x_1521 = ~v_1552 | v_2098;
assign x_1522 = ~v_1552 | v_120;
assign x_1523 = ~v_1553 | v_122;
assign x_1524 = ~v_1553 | ~v_2098;
assign x_1525 = ~v_1554 | v_121;
assign x_1526 = ~v_1554 | ~v_2098;
assign x_1527 = ~v_1555 | v_122;
assign x_1528 = ~v_1555 | v_121;
assign x_1529 = ~v_1556 | v_2097;
assign x_1530 = ~v_1556 | v_113;
assign x_1531 = ~v_1557 | v_2097;
assign x_1532 = ~v_1557 | v_118;
assign x_1533 = ~v_1558 | v_2096;
assign x_1534 = ~v_1558 | ~v_2097;
assign x_1535 = ~v_1559 | v_123;
assign x_1536 = ~v_1559 | ~v_2097;
assign x_1537 = ~v_1560 | v_2096;
assign x_1538 = ~v_1560 | v_123;
assign x_1539 = ~v_1561 | v_2095;
assign x_1540 = ~v_1561 | ~v_2096;
assign x_1541 = ~v_1562 | v_124;
assign x_1542 = ~v_1562 | ~v_2096;
assign x_1543 = ~v_1563 | v_2095;
assign x_1544 = ~v_1563 | v_124;
assign x_1545 = ~v_1564 | v_126;
assign x_1546 = ~v_1564 | ~v_2095;
assign x_1547 = ~v_1565 | v_125;
assign x_1548 = ~v_1565 | ~v_2095;
assign x_1549 = ~v_1566 | v_126;
assign x_1550 = ~v_1566 | v_125;
assign x_1551 = ~v_1567 | v_118;
assign x_1552 = ~v_1567 | ~v_2094;
assign x_1553 = ~v_1568 | v_113;
assign x_1554 = ~v_1568 | ~v_2094;
assign x_1555 = ~v_1569 | v_118;
assign x_1556 = ~v_1569 | v_113;
assign x_1557 = ~v_1570 | v_2093;
assign x_1558 = ~v_1570 | v_114;
assign x_1559 = ~v_1571 | v_2093;
assign x_1560 = ~v_1571 | v_119;
assign x_1561 = ~v_1572 | v_2093;
assign x_1562 = ~v_1572 | v_123;
assign x_1563 = ~v_1573 | v_2092;
assign x_1564 = ~v_1573 | ~v_2093;
assign x_1565 = ~v_1574 | v_127;
assign x_1566 = ~v_1574 | ~v_2093;
assign x_1567 = ~v_1575 | v_2092;
assign x_1568 = ~v_1575 | v_127;
assign x_1569 = ~v_1576 | v_129;
assign x_1570 = ~v_1576 | ~v_2092;
assign x_1571 = ~v_1577 | v_128;
assign x_1572 = ~v_1577 | ~v_2092;
assign x_1573 = ~v_1578 | v_129;
assign x_1574 = ~v_1578 | v_128;
assign x_1575 = ~v_1579 | v_2090;
assign x_1576 = ~v_1579 | ~v_2091;
assign x_1577 = ~v_1580 | v_114;
assign x_1578 = ~v_1580 | ~v_2091;
assign x_1579 = ~v_1581 | v_2090;
assign x_1580 = ~v_1581 | v_114;
assign x_1581 = ~v_1582 | v_123;
assign x_1582 = ~v_1582 | ~v_2090;
assign x_1583 = ~v_1583 | v_119;
assign x_1584 = ~v_1583 | ~v_2090;
assign x_1585 = ~v_1584 | v_123;
assign x_1586 = ~v_1584 | v_119;
assign x_1587 = ~v_1585 | v_2089;
assign x_1588 = ~v_1585 | v_115;
assign x_1589 = ~v_1586 | v_2089;
assign x_1590 = ~v_1586 | v_120;
assign x_1591 = ~v_1587 | v_2089;
assign x_1592 = ~v_1587 | v_124;
assign x_1593 = ~v_1588 | v_2089;
assign x_1594 = ~v_1588 | v_127;
assign x_1595 = ~v_1589 | v_131;
assign x_1596 = ~v_1589 | ~v_2089;
assign x_1597 = ~v_1590 | v_130;
assign x_1598 = ~v_1590 | ~v_2089;
assign x_1599 = ~v_1591 | v_131;
assign x_1600 = ~v_1591 | v_130;
assign x_1601 = ~v_1592 | v_2087;
assign x_1602 = ~v_1592 | ~v_2088;
assign x_1603 = ~v_1593 | v_115;
assign x_1604 = ~v_1593 | ~v_2088;
assign x_1605 = ~v_1594 | v_2087;
assign x_1606 = ~v_1594 | v_115;
assign x_1607 = ~v_1595 | v_2086;
assign x_1608 = ~v_1595 | ~v_2087;
assign x_1609 = ~v_1596 | v_120;
assign x_1610 = ~v_1596 | ~v_2087;
assign x_1611 = ~v_1597 | v_2086;
assign x_1612 = ~v_1597 | v_120;
assign x_1613 = ~v_1598 | v_127;
assign x_1614 = ~v_1598 | ~v_2086;
assign x_1615 = ~v_1599 | v_124;
assign x_1616 = ~v_1599 | ~v_2086;
assign x_1617 = ~v_1600 | v_127;
assign x_1618 = ~v_1600 | v_124;
assign x_1619 = ~v_1601 | v_132;
assign x_1620 = ~v_1601 | v_116;
assign x_1621 = ~v_1602 | v_132;
assign x_1622 = ~v_1602 | v_121;
assign x_1623 = ~v_1603 | v_132;
assign x_1624 = ~v_1603 | v_125;
assign x_1625 = ~v_1604 | v_132;
assign x_1626 = ~v_1604 | v_128;
assign x_1627 = ~v_1605 | v_132;
assign x_1628 = ~v_1605 | v_130;
assign x_1629 = ~v_1606 | v_2084;
assign x_1630 = ~v_1606 | ~v_2085;
assign x_1631 = ~v_1607 | v_116;
assign x_1632 = ~v_1607 | ~v_2085;
assign x_1633 = ~v_1608 | v_2084;
assign x_1634 = ~v_1608 | v_116;
assign x_1635 = ~v_1609 | v_2083;
assign x_1636 = ~v_1609 | ~v_2084;
assign x_1637 = ~v_1610 | v_121;
assign x_1638 = ~v_1610 | ~v_2084;
assign x_1639 = ~v_1611 | v_2083;
assign x_1640 = ~v_1611 | v_121;
assign x_1641 = ~v_1612 | v_2082;
assign x_1642 = ~v_1612 | ~v_2083;
assign x_1643 = ~v_1613 | v_125;
assign x_1644 = ~v_1613 | ~v_2083;
assign x_1645 = ~v_1614 | v_2082;
assign x_1646 = ~v_1614 | v_125;
assign x_1647 = ~v_1615 | v_130;
assign x_1648 = ~v_1615 | ~v_2082;
assign x_1649 = ~v_1616 | v_128;
assign x_1650 = ~v_1616 | ~v_2082;
assign x_1651 = ~v_1617 | v_130;
assign x_1652 = ~v_1617 | v_128;
assign x_1653 = ~v_1618 | v_2080;
assign x_1654 = ~v_1618 | ~v_2081;
assign x_1655 = ~v_1619 | v_117;
assign x_1656 = ~v_1619 | ~v_2081;
assign x_1657 = ~v_1620 | v_2080;
assign x_1658 = ~v_1620 | v_117;
assign x_1659 = ~v_1621 | v_2079;
assign x_1660 = ~v_1621 | ~v_2080;
assign x_1661 = ~v_1622 | v_122;
assign x_1662 = ~v_1622 | ~v_2080;
assign x_1663 = ~v_1623 | v_2079;
assign x_1664 = ~v_1623 | v_122;
assign x_1665 = ~v_1624 | v_2078;
assign x_1666 = ~v_1624 | ~v_2079;
assign x_1667 = ~v_1625 | v_126;
assign x_1668 = ~v_1625 | ~v_2079;
assign x_1669 = ~v_1626 | v_2078;
assign x_1670 = ~v_1626 | v_126;
assign x_1671 = ~v_1627 | v_2077;
assign x_1672 = ~v_1627 | ~v_2078;
assign x_1673 = ~v_1628 | v_129;
assign x_1674 = ~v_1628 | ~v_2078;
assign x_1675 = ~v_1629 | v_2077;
assign x_1676 = ~v_1629 | v_129;
assign x_1677 = ~v_1630 | v_132;
assign x_1678 = ~v_1630 | ~v_2077;
assign x_1679 = ~v_1631 | v_131;
assign x_1680 = ~v_1631 | ~v_2077;
assign x_1681 = ~v_1632 | v_132;
assign x_1682 = ~v_1632 | v_131;
assign x_1683 = ~v_1633 | v_2177;
assign x_1684 = ~v_1633 | ~v_2178;
assign x_1685 = ~v_1634 | v_138;
assign x_1686 = ~v_1634 | ~v_2178;
assign x_1687 = ~v_1635 | v_2177;
assign x_1688 = ~v_1635 | v_138;
assign x_1689 = ~v_1636 | v_2176;
assign x_1690 = ~v_1636 | ~v_2177;
assign x_1691 = ~v_1637 | v_137;
assign x_1692 = ~v_1637 | ~v_2177;
assign x_1693 = ~v_1638 | v_2176;
assign x_1694 = ~v_1638 | v_137;
assign x_1695 = ~v_1639 | v_2175;
assign x_1696 = ~v_1639 | ~v_2176;
assign x_1697 = ~v_1640 | v_136;
assign x_1698 = ~v_1640 | ~v_2176;
assign x_1699 = ~v_1641 | v_2175;
assign x_1700 = ~v_1641 | v_136;
assign x_1701 = ~v_1642 | v_2174;
assign x_1702 = ~v_1642 | ~v_2175;
assign x_1703 = ~v_1643 | v_135;
assign x_1704 = ~v_1643 | ~v_2175;
assign x_1705 = ~v_1644 | v_2174;
assign x_1706 = ~v_1644 | v_135;
assign x_1707 = ~v_1645 | v_133;
assign x_1708 = ~v_1645 | ~v_2174;
assign x_1709 = ~v_1646 | v_134;
assign x_1710 = ~v_1646 | ~v_2174;
assign x_1711 = ~v_1647 | v_133;
assign x_1712 = ~v_1647 | v_134;
assign x_1713 = ~v_1648 | v_2172;
assign x_1714 = ~v_1648 | ~v_2173;
assign x_1715 = ~v_1649 | v_143;
assign x_1716 = ~v_1649 | ~v_2173;
assign x_1717 = ~v_1650 | v_2172;
assign x_1718 = ~v_1650 | v_143;
assign x_1719 = ~v_1651 | v_2171;
assign x_1720 = ~v_1651 | ~v_2172;
assign x_1721 = ~v_1652 | v_142;
assign x_1722 = ~v_1652 | ~v_2172;
assign x_1723 = ~v_1653 | v_2171;
assign x_1724 = ~v_1653 | v_142;
assign x_1725 = ~v_1654 | v_2170;
assign x_1726 = ~v_1654 | ~v_2171;
assign x_1727 = ~v_1655 | v_141;
assign x_1728 = ~v_1655 | ~v_2171;
assign x_1729 = ~v_1656 | v_2170;
assign x_1730 = ~v_1656 | v_141;
assign x_1731 = ~v_1657 | v_139;
assign x_1732 = ~v_1657 | ~v_2170;
assign x_1733 = ~v_1658 | v_140;
assign x_1734 = ~v_1658 | ~v_2170;
assign x_1735 = ~v_1659 | v_139;
assign x_1736 = ~v_1659 | v_140;
assign x_1737 = ~v_1660 | v_133;
assign x_1738 = ~v_1660 | v_143;
assign x_1739 = ~v_1661 | v_133;
assign x_1740 = ~v_1661 | v_142;
assign x_1741 = ~v_1662 | v_133;
assign x_1742 = ~v_1662 | v_141;
assign x_1743 = ~v_1663 | v_133;
assign x_1744 = ~v_1663 | v_140;
assign x_1745 = ~v_1664 | v_133;
assign x_1746 = ~v_1664 | v_139;
assign x_1747 = ~v_1665 | v_2168;
assign x_1748 = ~v_1665 | ~v_2169;
assign x_1749 = ~v_1666 | v_147;
assign x_1750 = ~v_1666 | ~v_2169;
assign x_1751 = ~v_1667 | v_2168;
assign x_1752 = ~v_1667 | v_147;
assign x_1753 = ~v_1668 | v_2167;
assign x_1754 = ~v_1668 | ~v_2168;
assign x_1755 = ~v_1669 | v_146;
assign x_1756 = ~v_1669 | ~v_2168;
assign x_1757 = ~v_1670 | v_2167;
assign x_1758 = ~v_1670 | v_146;
assign x_1759 = ~v_1671 | v_144;
assign x_1760 = ~v_1671 | ~v_2167;
assign x_1761 = ~v_1672 | v_145;
assign x_1762 = ~v_1672 | ~v_2167;
assign x_1763 = ~v_1673 | v_144;
assign x_1764 = ~v_1673 | v_145;
assign x_1765 = ~v_1674 | v_2166;
assign x_1766 = ~v_1674 | v_147;
assign x_1767 = ~v_1675 | v_2166;
assign x_1768 = ~v_1675 | v_146;
assign x_1769 = ~v_1676 | v_2166;
assign x_1770 = ~v_1676 | v_145;
assign x_1771 = ~v_1677 | v_2166;
assign x_1772 = ~v_1677 | v_144;
assign x_1773 = ~v_1678 | v_134;
assign x_1774 = ~v_1678 | ~v_2166;
assign x_1775 = ~v_1679 | v_139;
assign x_1776 = ~v_1679 | ~v_2166;
assign x_1777 = ~v_1680 | v_134;
assign x_1778 = ~v_1680 | v_139;
assign x_1779 = ~v_1681 | v_2164;
assign x_1780 = ~v_1681 | ~v_2165;
assign x_1781 = ~v_1682 | v_150;
assign x_1782 = ~v_1682 | ~v_2165;
assign x_1783 = ~v_1683 | v_2164;
assign x_1784 = ~v_1683 | v_150;
assign x_1785 = ~v_1684 | v_148;
assign x_1786 = ~v_1684 | ~v_2164;
assign x_1787 = ~v_1685 | v_149;
assign x_1788 = ~v_1685 | ~v_2164;
assign x_1789 = ~v_1686 | v_148;
assign x_1790 = ~v_1686 | v_149;
assign x_1791 = ~v_1687 | v_2163;
assign x_1792 = ~v_1687 | v_150;
assign x_1793 = ~v_1688 | v_2163;
assign x_1794 = ~v_1688 | v_149;
assign x_1795 = ~v_1689 | v_2163;
assign x_1796 = ~v_1689 | v_148;
assign x_1797 = ~v_1690 | v_2162;
assign x_1798 = ~v_1690 | ~v_2163;
assign x_1799 = ~v_1691 | v_144;
assign x_1800 = ~v_1691 | ~v_2163;
assign x_1801 = ~v_1692 | v_2162;
assign x_1802 = ~v_1692 | v_144;
assign x_1803 = ~v_1693 | v_135;
assign x_1804 = ~v_1693 | ~v_2162;
assign x_1805 = ~v_1694 | v_140;
assign x_1806 = ~v_1694 | ~v_2162;
assign x_1807 = ~v_1695 | v_135;
assign x_1808 = ~v_1695 | v_140;
assign x_1809 = ~v_1696 | v_151;
assign x_1810 = ~v_1696 | ~v_2161;
assign x_1811 = ~v_1697 | v_152;
assign x_1812 = ~v_1697 | ~v_2161;
assign x_1813 = ~v_1698 | v_151;
assign x_1814 = ~v_1698 | v_152;
assign x_1815 = ~v_1699 | v_2160;
assign x_1816 = ~v_1699 | v_152;
assign x_1817 = ~v_1700 | v_2160;
assign x_1818 = ~v_1700 | v_151;
assign x_1819 = ~v_1701 | v_2159;
assign x_1820 = ~v_1701 | ~v_2160;
assign x_1821 = ~v_1702 | v_148;
assign x_1822 = ~v_1702 | ~v_2160;
assign x_1823 = ~v_1703 | v_2159;
assign x_1824 = ~v_1703 | v_148;
assign x_1825 = ~v_1704 | v_2158;
assign x_1826 = ~v_1704 | ~v_2159;
assign x_1827 = ~v_1705 | v_145;
assign x_1828 = ~v_1705 | ~v_2159;
assign x_1829 = ~v_1706 | v_2158;
assign x_1830 = ~v_1706 | v_145;
assign x_1831 = ~v_1707 | v_136;
assign x_1832 = ~v_1707 | ~v_2158;
assign x_1833 = ~v_1708 | v_141;
assign x_1834 = ~v_1708 | ~v_2158;
assign x_1835 = ~v_1709 | v_136;
assign x_1836 = ~v_1709 | v_141;
assign x_1837 = ~v_1710 | v_2157;
assign x_1838 = ~v_1710 | v_153;
assign x_1839 = ~v_1711 | v_2156;
assign x_1840 = ~v_1711 | ~v_2157;
assign x_1841 = ~v_1712 | v_151;
assign x_1842 = ~v_1712 | ~v_2157;
assign x_1843 = ~v_1713 | v_2156;
assign x_1844 = ~v_1713 | v_151;
assign x_1845 = ~v_1714 | v_2155;
assign x_1846 = ~v_1714 | ~v_2156;
assign x_1847 = ~v_1715 | v_149;
assign x_1848 = ~v_1715 | ~v_2156;
assign x_1849 = ~v_1716 | v_2155;
assign x_1850 = ~v_1716 | v_149;
assign x_1851 = ~v_1717 | v_2154;
assign x_1852 = ~v_1717 | ~v_2155;
assign x_1853 = ~v_1718 | v_146;
assign x_1854 = ~v_1718 | ~v_2155;
assign x_1855 = ~v_1719 | v_2154;
assign x_1856 = ~v_1719 | v_146;
assign x_1857 = ~v_1720 | v_137;
assign x_1858 = ~v_1720 | ~v_2154;
assign x_1859 = ~v_1721 | v_142;
assign x_1860 = ~v_1721 | ~v_2154;
assign x_1861 = ~v_1722 | v_137;
assign x_1862 = ~v_1722 | v_142;
assign x_1863 = ~v_1723 | v_2152;
assign x_1864 = ~v_1723 | ~v_2153;
assign x_1865 = ~v_1724 | v_153;
assign x_1866 = ~v_1724 | ~v_2153;
assign x_1867 = ~v_1725 | v_2152;
assign x_1868 = ~v_1725 | v_153;
assign x_1869 = ~v_1726 | v_2151;
assign x_1870 = ~v_1726 | ~v_2152;
assign x_1871 = ~v_1727 | v_152;
assign x_1872 = ~v_1727 | ~v_2152;
assign x_1873 = ~v_1728 | v_2151;
assign x_1874 = ~v_1728 | v_152;
assign x_1875 = ~v_1729 | v_2150;
assign x_1876 = ~v_1729 | ~v_2151;
assign x_1877 = ~v_1730 | v_150;
assign x_1878 = ~v_1730 | ~v_2151;
assign x_1879 = ~v_1731 | v_2150;
assign x_1880 = ~v_1731 | v_150;
assign x_1881 = ~v_1732 | v_2149;
assign x_1882 = ~v_1732 | ~v_2150;
assign x_1883 = ~v_1733 | v_147;
assign x_1884 = ~v_1733 | ~v_2150;
assign x_1885 = ~v_1734 | v_2149;
assign x_1886 = ~v_1734 | v_147;
assign x_1887 = ~v_1735 | v_138;
assign x_1888 = ~v_1735 | ~v_2149;
assign x_1889 = ~v_1736 | v_143;
assign x_1890 = ~v_1736 | ~v_2149;
assign x_1891 = ~v_1737 | v_138;
assign x_1892 = ~v_1737 | v_143;
assign x_1893 = ~v_1738 | v_2207;
assign x_1894 = ~v_1738 | ~v_2208;
assign x_1895 = ~v_1739 | v_133;
assign x_1896 = ~v_1739 | ~v_2208;
assign x_1897 = ~v_1740 | v_2207;
assign x_1898 = ~v_1740 | v_133;
assign x_1899 = ~v_1741 | v_2206;
assign x_1900 = ~v_1741 | ~v_2207;
assign x_1901 = ~v_1742 | v_134;
assign x_1902 = ~v_1742 | ~v_2207;
assign x_1903 = ~v_1743 | v_2206;
assign x_1904 = ~v_1743 | v_134;
assign x_1905 = ~v_1744 | v_2205;
assign x_1906 = ~v_1744 | ~v_2206;
assign x_1907 = ~v_1745 | v_135;
assign x_1908 = ~v_1745 | ~v_2206;
assign x_1909 = ~v_1746 | v_2205;
assign x_1910 = ~v_1746 | v_135;
assign x_1911 = ~v_1747 | v_2204;
assign x_1912 = ~v_1747 | ~v_2205;
assign x_1913 = ~v_1748 | v_136;
assign x_1914 = ~v_1748 | ~v_2205;
assign x_1915 = ~v_1749 | v_2204;
assign x_1916 = ~v_1749 | v_136;
assign x_1917 = ~v_1750 | v_138;
assign x_1918 = ~v_1750 | ~v_2204;
assign x_1919 = ~v_1751 | v_137;
assign x_1920 = ~v_1751 | ~v_2204;
assign x_1921 = ~v_1752 | v_138;
assign x_1922 = ~v_1752 | v_137;
assign x_1923 = ~v_1753 | v_2203;
assign x_1924 = ~v_1753 | v_133;
assign x_1925 = ~v_1754 | v_2202;
assign x_1926 = ~v_1754 | ~v_2203;
assign x_1927 = ~v_1755 | v_139;
assign x_1928 = ~v_1755 | ~v_2203;
assign x_1929 = ~v_1756 | v_2202;
assign x_1930 = ~v_1756 | v_139;
assign x_1931 = ~v_1757 | v_2201;
assign x_1932 = ~v_1757 | ~v_2202;
assign x_1933 = ~v_1758 | v_140;
assign x_1934 = ~v_1758 | ~v_2202;
assign x_1935 = ~v_1759 | v_2201;
assign x_1936 = ~v_1759 | v_140;
assign x_1937 = ~v_1760 | v_2200;
assign x_1938 = ~v_1760 | ~v_2201;
assign x_1939 = ~v_1761 | v_141;
assign x_1940 = ~v_1761 | ~v_2201;
assign x_1941 = ~v_1762 | v_2200;
assign x_1942 = ~v_1762 | v_141;
assign x_1943 = ~v_1763 | v_143;
assign x_1944 = ~v_1763 | ~v_2200;
assign x_1945 = ~v_1764 | v_142;
assign x_1946 = ~v_1764 | ~v_2200;
assign x_1947 = ~v_1765 | v_143;
assign x_1948 = ~v_1765 | v_142;
assign x_1949 = ~v_1766 | v_2199;
assign x_1950 = ~v_1766 | v_134;
assign x_1951 = ~v_1767 | v_2199;
assign x_1952 = ~v_1767 | v_139;
assign x_1953 = ~v_1768 | v_2198;
assign x_1954 = ~v_1768 | ~v_2199;
assign x_1955 = ~v_1769 | v_144;
assign x_1956 = ~v_1769 | ~v_2199;
assign x_1957 = ~v_1770 | v_2198;
assign x_1958 = ~v_1770 | v_144;
assign x_1959 = ~v_1771 | v_2197;
assign x_1960 = ~v_1771 | ~v_2198;
assign x_1961 = ~v_1772 | v_145;
assign x_1962 = ~v_1772 | ~v_2198;
assign x_1963 = ~v_1773 | v_2197;
assign x_1964 = ~v_1773 | v_145;
assign x_1965 = ~v_1774 | v_147;
assign x_1966 = ~v_1774 | ~v_2197;
assign x_1967 = ~v_1775 | v_146;
assign x_1968 = ~v_1775 | ~v_2197;
assign x_1969 = ~v_1776 | v_147;
assign x_1970 = ~v_1776 | v_146;
assign x_1971 = ~v_1777 | v_139;
assign x_1972 = ~v_1777 | ~v_2196;
assign x_1973 = ~v_1778 | v_134;
assign x_1974 = ~v_1778 | ~v_2196;
assign x_1975 = ~v_1779 | v_139;
assign x_1976 = ~v_1779 | v_134;
assign x_1977 = ~v_1780 | v_2195;
assign x_1978 = ~v_1780 | v_135;
assign x_1979 = ~v_1781 | v_2195;
assign x_1980 = ~v_1781 | v_140;
assign x_1981 = ~v_1782 | v_2195;
assign x_1982 = ~v_1782 | v_144;
assign x_1983 = ~v_1783 | v_2194;
assign x_1984 = ~v_1783 | ~v_2195;
assign x_1985 = ~v_1784 | v_148;
assign x_1986 = ~v_1784 | ~v_2195;
assign x_1987 = ~v_1785 | v_2194;
assign x_1988 = ~v_1785 | v_148;
assign x_1989 = ~v_1786 | v_150;
assign x_1990 = ~v_1786 | ~v_2194;
assign x_1991 = ~v_1787 | v_149;
assign x_1992 = ~v_1787 | ~v_2194;
assign x_1993 = ~v_1788 | v_150;
assign x_1994 = ~v_1788 | v_149;
assign x_1995 = ~v_1789 | v_2192;
assign x_1996 = ~v_1789 | ~v_2193;
assign x_1997 = ~v_1790 | v_135;
assign x_1998 = ~v_1790 | ~v_2193;
assign x_1999 = ~v_1791 | v_2192;
assign x_2000 = ~v_1791 | v_135;
assign x_2001 = ~v_1792 | v_144;
assign x_2002 = ~v_1792 | ~v_2192;
assign x_2003 = ~v_1793 | v_140;
assign x_2004 = ~v_1793 | ~v_2192;
assign x_2005 = ~v_1794 | v_144;
assign x_2006 = ~v_1794 | v_140;
assign x_2007 = ~v_1795 | v_2191;
assign x_2008 = ~v_1795 | v_136;
assign x_2009 = ~v_1796 | v_2191;
assign x_2010 = ~v_1796 | v_141;
assign x_2011 = ~v_1797 | v_2191;
assign x_2012 = ~v_1797 | v_145;
assign x_2013 = ~v_1798 | v_2191;
assign x_2014 = ~v_1798 | v_148;
assign x_2015 = ~v_1799 | v_152;
assign x_2016 = ~v_1799 | ~v_2191;
assign x_2017 = ~v_1800 | v_151;
assign x_2018 = ~v_1800 | ~v_2191;
assign x_2019 = ~v_1801 | v_152;
assign x_2020 = ~v_1801 | v_151;
assign x_2021 = ~v_1802 | v_2189;
assign x_2022 = ~v_1802 | ~v_2190;
assign x_2023 = ~v_1803 | v_136;
assign x_2024 = ~v_1803 | ~v_2190;
assign x_2025 = ~v_1804 | v_2189;
assign x_2026 = ~v_1804 | v_136;
assign x_2027 = ~v_1805 | v_2188;
assign x_2028 = ~v_1805 | ~v_2189;
assign x_2029 = ~v_1806 | v_141;
assign x_2030 = ~v_1806 | ~v_2189;
assign x_2031 = ~v_1807 | v_2188;
assign x_2032 = ~v_1807 | v_141;
assign x_2033 = ~v_1808 | v_148;
assign x_2034 = ~v_1808 | ~v_2188;
assign x_2035 = ~v_1809 | v_145;
assign x_2036 = ~v_1809 | ~v_2188;
assign x_2037 = ~v_1810 | v_148;
assign x_2038 = ~v_1810 | v_145;
assign x_2039 = ~v_1811 | v_153;
assign x_2040 = ~v_1811 | v_137;
assign x_2041 = ~v_1812 | v_153;
assign x_2042 = ~v_1812 | v_142;
assign x_2043 = ~v_1813 | v_153;
assign x_2044 = ~v_1813 | v_146;
assign x_2045 = ~v_1814 | v_153;
assign x_2046 = ~v_1814 | v_149;
assign x_2047 = ~v_1815 | v_153;
assign x_2048 = ~v_1815 | v_151;
assign x_2049 = ~v_1816 | v_2186;
assign x_2050 = ~v_1816 | ~v_2187;
assign x_2051 = ~v_1817 | v_137;
assign x_2052 = ~v_1817 | ~v_2187;
assign x_2053 = ~v_1818 | v_2186;
assign x_2054 = ~v_1818 | v_137;
assign x_2055 = ~v_1819 | v_2185;
assign x_2056 = ~v_1819 | ~v_2186;
assign x_2057 = ~v_1820 | v_142;
assign x_2058 = ~v_1820 | ~v_2186;
assign x_2059 = ~v_1821 | v_2185;
assign x_2060 = ~v_1821 | v_142;
assign x_2061 = ~v_1822 | v_2184;
assign x_2062 = ~v_1822 | ~v_2185;
assign x_2063 = ~v_1823 | v_146;
assign x_2064 = ~v_1823 | ~v_2185;
assign x_2065 = ~v_1824 | v_2184;
assign x_2066 = ~v_1824 | v_146;
assign x_2067 = ~v_1825 | v_151;
assign x_2068 = ~v_1825 | ~v_2184;
assign x_2069 = ~v_1826 | v_149;
assign x_2070 = ~v_1826 | ~v_2184;
assign x_2071 = ~v_1827 | v_151;
assign x_2072 = ~v_1827 | v_149;
assign x_2073 = ~v_1828 | v_2182;
assign x_2074 = ~v_1828 | ~v_2183;
assign x_2075 = ~v_1829 | v_138;
assign x_2076 = ~v_1829 | ~v_2183;
assign x_2077 = ~v_1830 | v_2182;
assign x_2078 = ~v_1830 | v_138;
assign x_2079 = ~v_1831 | v_2181;
assign x_2080 = ~v_1831 | ~v_2182;
assign x_2081 = ~v_1832 | v_143;
assign x_2082 = ~v_1832 | ~v_2182;
assign x_2083 = ~v_1833 | v_2181;
assign x_2084 = ~v_1833 | v_143;
assign x_2085 = ~v_1834 | v_2180;
assign x_2086 = ~v_1834 | ~v_2181;
assign x_2087 = ~v_1835 | v_147;
assign x_2088 = ~v_1835 | ~v_2181;
assign x_2089 = ~v_1836 | v_2180;
assign x_2090 = ~v_1836 | v_147;
assign x_2091 = ~v_1837 | v_2179;
assign x_2092 = ~v_1837 | ~v_2180;
assign x_2093 = ~v_1838 | v_150;
assign x_2094 = ~v_1838 | ~v_2180;
assign x_2095 = ~v_1839 | v_2179;
assign x_2096 = ~v_1839 | v_150;
assign x_2097 = ~v_1840 | v_153;
assign x_2098 = ~v_1840 | ~v_2179;
assign x_2099 = ~v_1841 | v_152;
assign x_2100 = ~v_1841 | ~v_2179;
assign x_2101 = ~v_1842 | v_153;
assign x_2102 = ~v_1842 | v_152;
assign x_2103 = ~v_770 | v_1 | ~v_9;
assign x_2104 = ~v_770 | ~v_1 | v_9 | v_219 | v_218 | v_217 | v_216 | v_215 | v_214;
assign x_2105 = ~v_770 | ~v_219 | v_769;
assign x_2106 = ~v_770 | ~v_49 | ~v_1 | v_2 | v_219;
assign x_2107 = ~v_770 | ~v_218 | v_768;
assign x_2108 = ~v_770 | ~v_50 | ~v_1 | v_3 | v_218;
assign x_2109 = ~v_770 | ~v_217 | v_767;
assign x_2110 = ~v_770 | ~v_51 | ~v_1 | v_4 | v_217;
assign x_2111 = ~v_770 | ~v_216 | v_766;
assign x_2112 = ~v_770 | ~v_52 | ~v_1 | v_5 | v_216;
assign x_2113 = ~v_770 | ~v_215 | v_765;
assign x_2114 = ~v_770 | ~v_53 | ~v_1 | v_6 | v_215;
assign x_2115 = ~v_770 | ~v_214 | v_764;
assign x_2116 = ~v_770 | ~v_54 | ~v_1 | v_7 | v_214;
assign x_2117 = ~v_770 | v_2 | ~v_10 | v_220;
assign x_2118 = ~v_770 | ~v_2 | v_10 | v_225 | v_224 | v_223 | v_222 | v_221;
assign x_2119 = ~v_770 | ~v_220 | v_763;
assign x_2120 = ~v_770 | ~v_49 | ~v_1 | v_2 | v_220;
assign x_2121 = ~v_770 | ~v_225 | v_762;
assign x_2122 = ~v_770 | ~v_55 | ~v_2 | v_3 | v_225;
assign x_2123 = ~v_770 | ~v_224 | v_761;
assign x_2124 = ~v_770 | ~v_56 | ~v_2 | v_4 | v_224;
assign x_2125 = ~v_770 | ~v_223 | v_760;
assign x_2126 = ~v_770 | ~v_57 | ~v_2 | v_5 | v_223;
assign x_2127 = ~v_770 | ~v_222 | v_759;
assign x_2128 = ~v_770 | ~v_58 | ~v_2 | v_6 | v_222;
assign x_2129 = ~v_770 | ~v_221 | v_758;
assign x_2130 = ~v_770 | ~v_59 | ~v_2 | v_7 | v_221;
assign x_2131 = ~v_770 | v_3 | ~v_11 | v_227 | v_226;
assign x_2132 = ~v_770 | ~v_3 | v_11 | v_231 | v_230 | v_229 | v_228;
assign x_2133 = ~v_770 | ~v_227 | v_757;
assign x_2134 = ~v_770 | ~v_50 | ~v_1 | v_3 | v_227;
assign x_2135 = ~v_770 | ~v_226 | v_756;
assign x_2136 = ~v_770 | ~v_55 | ~v_2 | v_3 | v_226;
assign x_2137 = ~v_770 | ~v_231 | v_755;
assign x_2138 = ~v_770 | ~v_60 | ~v_3 | v_4 | v_231;
assign x_2139 = ~v_770 | ~v_230 | v_754;
assign x_2140 = ~v_770 | ~v_61 | ~v_3 | v_5 | v_230;
assign x_2141 = ~v_770 | ~v_229 | v_753;
assign x_2142 = ~v_770 | ~v_62 | ~v_3 | v_6 | v_229;
assign x_2143 = ~v_770 | ~v_228 | v_752;
assign x_2144 = ~v_770 | ~v_63 | ~v_3 | v_7 | v_228;
assign x_2145 = ~v_770 | v_4 | ~v_12 | v_234 | v_233 | v_232;
assign x_2146 = ~v_770 | ~v_4 | v_12 | v_237 | v_236 | v_235;
assign x_2147 = ~v_770 | ~v_234 | v_751;
assign x_2148 = ~v_770 | ~v_51 | ~v_1 | v_4 | v_234;
assign x_2149 = ~v_770 | ~v_233 | v_750;
assign x_2150 = ~v_770 | ~v_56 | ~v_2 | v_4 | v_233;
assign x_2151 = ~v_770 | ~v_232 | v_749;
assign x_2152 = ~v_770 | ~v_60 | ~v_3 | v_4 | v_232;
assign x_2153 = ~v_770 | ~v_237 | v_748;
assign x_2154 = ~v_770 | ~v_64 | ~v_4 | v_5 | v_237;
assign x_2155 = ~v_770 | ~v_236 | v_747;
assign x_2156 = ~v_770 | ~v_65 | ~v_4 | v_6 | v_236;
assign x_2157 = ~v_770 | ~v_235 | v_746;
assign x_2158 = ~v_770 | ~v_66 | ~v_4 | v_7 | v_235;
assign x_2159 = ~v_770 | v_5 | ~v_13 | v_241 | v_240 | v_239 | v_238;
assign x_2160 = ~v_770 | ~v_5 | v_13 | v_243 | v_242;
assign x_2161 = ~v_770 | ~v_241 | v_745;
assign x_2162 = ~v_770 | ~v_52 | ~v_1 | v_5 | v_241;
assign x_2163 = ~v_770 | ~v_240 | v_744;
assign x_2164 = ~v_770 | ~v_57 | ~v_2 | v_5 | v_240;
assign x_2165 = ~v_770 | ~v_239 | v_743;
assign x_2166 = ~v_770 | ~v_61 | ~v_3 | v_5 | v_239;
assign x_2167 = ~v_770 | ~v_238 | v_742;
assign x_2168 = ~v_770 | ~v_64 | ~v_4 | v_5 | v_238;
assign x_2169 = ~v_770 | ~v_243 | v_741;
assign x_2170 = ~v_770 | ~v_67 | ~v_5 | v_6 | v_243;
assign x_2171 = ~v_770 | ~v_242 | v_740;
assign x_2172 = ~v_770 | ~v_68 | ~v_5 | v_7 | v_242;
assign x_2173 = ~v_770 | v_6 | ~v_14 | v_248 | v_247 | v_246 | v_245 | v_244;
assign x_2174 = ~v_770 | ~v_6 | v_14 | v_249;
assign x_2175 = ~v_770 | ~v_248 | v_739;
assign x_2176 = ~v_770 | ~v_53 | ~v_1 | v_6 | v_248;
assign x_2177 = ~v_770 | ~v_247 | v_738;
assign x_2178 = ~v_770 | ~v_58 | ~v_2 | v_6 | v_247;
assign x_2179 = ~v_770 | ~v_246 | v_737;
assign x_2180 = ~v_770 | ~v_62 | ~v_3 | v_6 | v_246;
assign x_2181 = ~v_770 | ~v_245 | v_736;
assign x_2182 = ~v_770 | ~v_65 | ~v_4 | v_6 | v_245;
assign x_2183 = ~v_770 | ~v_244 | v_735;
assign x_2184 = ~v_770 | ~v_67 | ~v_5 | v_6 | v_244;
assign x_2185 = ~v_770 | ~v_249 | v_734;
assign x_2186 = ~v_770 | ~v_69 | ~v_6 | v_7 | v_249;
assign x_2187 = ~v_770 | v_7 | ~v_15 | v_255 | v_254 | v_253 | v_252 | v_251 | v_250;
assign x_2188 = ~v_770 | ~v_7 | v_15;
assign x_2189 = ~v_770 | ~v_255 | v_733;
assign x_2190 = ~v_770 | ~v_54 | ~v_1 | v_7 | v_255;
assign x_2191 = ~v_770 | ~v_254 | v_732;
assign x_2192 = ~v_770 | ~v_59 | ~v_2 | v_7 | v_254;
assign x_2193 = ~v_770 | ~v_253 | v_731;
assign x_2194 = ~v_770 | ~v_63 | ~v_3 | v_7 | v_253;
assign x_2195 = ~v_770 | ~v_252 | v_730;
assign x_2196 = ~v_770 | ~v_66 | ~v_4 | v_7 | v_252;
assign x_2197 = ~v_770 | ~v_251 | v_729;
assign x_2198 = ~v_770 | ~v_68 | ~v_5 | v_7 | v_251;
assign x_2199 = ~v_770 | ~v_250 | v_728;
assign x_2200 = ~v_770 | ~v_69 | ~v_6 | v_7 | v_250;
assign x_2201 = ~v_770 | v_8 | ~v_16;
assign x_2202 = ~v_770 | ~v_8 | v_16;
assign x_2203 = ~v_770 | v_726 | v_727;
assign x_2204 = ~v_770 | v_724 | v_725;
assign x_2205 = ~v_770 | v_722 | v_723;
assign x_2206 = ~v_770 | v_720 | v_721;
assign x_2207 = ~v_770 | v_718 | v_719;
assign x_2208 = ~v_770 | v_716 | v_717;
assign x_2209 = ~v_770 | v_714 | v_715;
assign x_2210 = ~v_770 | v_712 | v_713;
assign x_2211 = ~v_770 | v_710 | v_711;
assign x_2212 = ~v_770 | v_708 | v_709;
assign x_2213 = ~v_770 | v_706 | v_707;
assign x_2214 = ~v_770 | v_704 | v_705;
assign x_2215 = ~v_770 | v_702 | v_703;
assign x_2216 = ~v_770 | v_700 | v_701;
assign x_2217 = ~v_770 | v_698 | v_699;
assign x_2218 = ~v_770 | v_696 | v_697;
assign x_2219 = ~v_770 | v_694 | v_695;
assign x_2220 = ~v_770 | v_692 | v_693;
assign x_2221 = ~v_770 | v_690 | v_691;
assign x_2222 = ~v_770 | v_688 | v_689;
assign x_2223 = ~v_770 | v_686 | v_687;
assign x_2224 = ~v_770 | v_664;
assign x_2225 = ~v_769 | v_49;
assign x_2226 = ~v_769 | v_1;
assign x_2227 = ~v_769 | ~v_2;
assign x_2228 = ~v_768 | v_50;
assign x_2229 = ~v_768 | v_1;
assign x_2230 = ~v_768 | ~v_3;
assign x_2231 = ~v_767 | v_51;
assign x_2232 = ~v_767 | v_1;
assign x_2233 = ~v_767 | ~v_4;
assign x_2234 = ~v_766 | v_52;
assign x_2235 = ~v_766 | v_1;
assign x_2236 = ~v_766 | ~v_5;
assign x_2237 = ~v_765 | v_53;
assign x_2238 = ~v_765 | v_1;
assign x_2239 = ~v_765 | ~v_6;
assign x_2240 = ~v_764 | v_54;
assign x_2241 = ~v_764 | v_1;
assign x_2242 = ~v_764 | ~v_7;
assign x_2243 = ~v_763 | v_49;
assign x_2244 = ~v_763 | v_1;
assign x_2245 = ~v_763 | ~v_2;
assign x_2246 = ~v_762 | v_55;
assign x_2247 = ~v_762 | v_2;
assign x_2248 = ~v_762 | ~v_3;
assign x_2249 = ~v_761 | v_56;
assign x_2250 = ~v_761 | v_2;
assign x_2251 = ~v_761 | ~v_4;
assign x_2252 = ~v_760 | v_57;
assign x_2253 = ~v_760 | v_2;
assign x_2254 = ~v_760 | ~v_5;
assign x_2255 = ~v_759 | v_58;
assign x_2256 = ~v_759 | v_2;
assign x_2257 = ~v_759 | ~v_6;
assign x_2258 = ~v_758 | v_59;
assign x_2259 = ~v_758 | v_2;
assign x_2260 = ~v_758 | ~v_7;
assign x_2261 = ~v_757 | v_50;
assign x_2262 = ~v_757 | v_1;
assign x_2263 = ~v_757 | ~v_3;
assign x_2264 = ~v_756 | v_55;
assign x_2265 = ~v_756 | v_2;
assign x_2266 = ~v_756 | ~v_3;
assign x_2267 = ~v_755 | v_60;
assign x_2268 = ~v_755 | v_3;
assign x_2269 = ~v_755 | ~v_4;
assign x_2270 = ~v_754 | v_61;
assign x_2271 = ~v_754 | v_3;
assign x_2272 = ~v_754 | ~v_5;
assign x_2273 = ~v_753 | v_62;
assign x_2274 = ~v_753 | v_3;
assign x_2275 = ~v_753 | ~v_6;
assign x_2276 = ~v_752 | v_63;
assign x_2277 = ~v_752 | v_3;
assign x_2278 = ~v_752 | ~v_7;
assign x_2279 = ~v_751 | v_51;
assign x_2280 = ~v_751 | v_1;
assign x_2281 = ~v_751 | ~v_4;
assign x_2282 = ~v_750 | v_56;
assign x_2283 = ~v_750 | v_2;
assign x_2284 = ~v_750 | ~v_4;
assign x_2285 = ~v_749 | v_60;
assign x_2286 = ~v_749 | v_3;
assign x_2287 = ~v_749 | ~v_4;
assign x_2288 = ~v_748 | v_64;
assign x_2289 = ~v_748 | v_4;
assign x_2290 = ~v_748 | ~v_5;
assign x_2291 = ~v_747 | v_65;
assign x_2292 = ~v_747 | v_4;
assign x_2293 = ~v_747 | ~v_6;
assign x_2294 = ~v_746 | v_66;
assign x_2295 = ~v_746 | v_4;
assign x_2296 = ~v_746 | ~v_7;
assign x_2297 = ~v_745 | v_52;
assign x_2298 = ~v_745 | v_1;
assign x_2299 = ~v_745 | ~v_5;
assign x_2300 = ~v_744 | v_57;
assign x_2301 = ~v_744 | v_2;
assign x_2302 = ~v_744 | ~v_5;
assign x_2303 = ~v_743 | v_61;
assign x_2304 = ~v_743 | v_3;
assign x_2305 = ~v_743 | ~v_5;
assign x_2306 = ~v_742 | v_64;
assign x_2307 = ~v_742 | v_4;
assign x_2308 = ~v_742 | ~v_5;
assign x_2309 = ~v_741 | v_67;
assign x_2310 = ~v_741 | v_5;
assign x_2311 = ~v_741 | ~v_6;
assign x_2312 = ~v_740 | v_68;
assign x_2313 = ~v_740 | v_5;
assign x_2314 = ~v_740 | ~v_7;
assign x_2315 = ~v_739 | v_53;
assign x_2316 = ~v_739 | v_1;
assign x_2317 = ~v_739 | ~v_6;
assign x_2318 = ~v_738 | v_58;
assign x_2319 = ~v_738 | v_2;
assign x_2320 = ~v_738 | ~v_6;
assign x_2321 = ~v_737 | v_62;
assign x_2322 = ~v_737 | v_3;
assign x_2323 = ~v_737 | ~v_6;
assign x_2324 = ~v_736 | v_65;
assign x_2325 = ~v_736 | v_4;
assign x_2326 = ~v_736 | ~v_6;
assign x_2327 = ~v_735 | v_67;
assign x_2328 = ~v_735 | v_5;
assign x_2329 = ~v_735 | ~v_6;
assign x_2330 = ~v_734 | v_69;
assign x_2331 = ~v_734 | v_6;
assign x_2332 = ~v_734 | ~v_7;
assign x_2333 = ~v_733 | v_54;
assign x_2334 = ~v_733 | v_1;
assign x_2335 = ~v_733 | ~v_7;
assign x_2336 = ~v_732 | v_59;
assign x_2337 = ~v_732 | v_2;
assign x_2338 = ~v_732 | ~v_7;
assign x_2339 = ~v_731 | v_63;
assign x_2340 = ~v_731 | v_3;
assign x_2341 = ~v_731 | ~v_7;
assign x_2342 = ~v_730 | v_66;
assign x_2343 = ~v_730 | v_4;
assign x_2344 = ~v_730 | ~v_7;
assign x_2345 = ~v_729 | v_68;
assign x_2346 = ~v_729 | v_5;
assign x_2347 = ~v_729 | ~v_7;
assign x_2348 = ~v_728 | v_69;
assign x_2349 = ~v_728 | v_6;
assign x_2350 = ~v_728 | ~v_7;
assign x_2351 = ~v_726 | ~v_49 | ~v_1 | v_2;
assign x_2352 = ~v_727 | ~v_9;
assign x_2353 = ~v_727 | v_10;
assign x_2354 = ~v_724 | ~v_50 | ~v_1 | v_3;
assign x_2355 = ~v_725 | ~v_9;
assign x_2356 = ~v_725 | v_11;
assign x_2357 = ~v_722 | ~v_51 | ~v_1 | v_4;
assign x_2358 = ~v_723 | ~v_9;
assign x_2359 = ~v_723 | v_12;
assign x_2360 = ~v_720 | ~v_52 | ~v_1 | v_5;
assign x_2361 = ~v_721 | ~v_9;
assign x_2362 = ~v_721 | v_13;
assign x_2363 = ~v_718 | ~v_53 | ~v_1 | v_6;
assign x_2364 = ~v_719 | ~v_9;
assign x_2365 = ~v_719 | v_14;
assign x_2366 = ~v_716 | ~v_54 | ~v_1 | v_7;
assign x_2367 = ~v_717 | ~v_9;
assign x_2368 = ~v_717 | v_15;
assign x_2369 = ~v_714 | ~v_55 | ~v_2 | v_3;
assign x_2370 = ~v_715 | ~v_10;
assign x_2371 = ~v_715 | v_11;
assign x_2372 = ~v_712 | ~v_56 | ~v_2 | v_4;
assign x_2373 = ~v_713 | ~v_10;
assign x_2374 = ~v_713 | v_12;
assign x_2375 = ~v_710 | ~v_57 | ~v_2 | v_5;
assign x_2376 = ~v_711 | ~v_10;
assign x_2377 = ~v_711 | v_13;
assign x_2378 = ~v_708 | ~v_58 | ~v_2 | v_6;
assign x_2379 = ~v_709 | ~v_10;
assign x_2380 = ~v_709 | v_14;
assign x_2381 = ~v_706 | ~v_59 | ~v_2 | v_7;
assign x_2382 = ~v_707 | ~v_10;
assign x_2383 = ~v_707 | v_15;
assign x_2384 = ~v_704 | ~v_60 | ~v_3 | v_4;
assign x_2385 = ~v_705 | ~v_11;
assign x_2386 = ~v_705 | v_12;
assign x_2387 = ~v_702 | ~v_61 | ~v_3 | v_5;
assign x_2388 = ~v_703 | ~v_11;
assign x_2389 = ~v_703 | v_13;
assign x_2390 = ~v_700 | ~v_62 | ~v_3 | v_6;
assign x_2391 = ~v_701 | ~v_11;
assign x_2392 = ~v_701 | v_14;
assign x_2393 = ~v_698 | ~v_63 | ~v_3 | v_7;
assign x_2394 = ~v_699 | ~v_11;
assign x_2395 = ~v_699 | v_15;
assign x_2396 = ~v_696 | ~v_64 | ~v_4 | v_5;
assign x_2397 = ~v_697 | ~v_12;
assign x_2398 = ~v_697 | v_13;
assign x_2399 = ~v_694 | ~v_65 | ~v_4 | v_6;
assign x_2400 = ~v_695 | ~v_12;
assign x_2401 = ~v_695 | v_14;
assign x_2402 = ~v_692 | ~v_66 | ~v_4 | v_7;
assign x_2403 = ~v_693 | ~v_12;
assign x_2404 = ~v_693 | v_15;
assign x_2405 = ~v_690 | ~v_67 | ~v_5 | v_6;
assign x_2406 = ~v_691 | ~v_13;
assign x_2407 = ~v_691 | v_14;
assign x_2408 = ~v_688 | ~v_68 | ~v_5 | v_7;
assign x_2409 = ~v_689 | ~v_13;
assign x_2410 = ~v_689 | v_15;
assign x_2411 = ~v_686 | ~v_69 | ~v_6 | v_7;
assign x_2412 = ~v_687 | ~v_14;
assign x_2413 = ~v_687 | v_15;
assign x_2414 = ~v_664 | v_9 | ~v_17;
assign x_2415 = ~v_664 | ~v_9 | v_17 | v_1908 | v_1907 | v_1906 | v_1905 | v_1904 | v_1903;
assign x_2416 = ~v_664 | ~v_1908 | v_663;
assign x_2417 = ~v_664 | ~v_70 | ~v_9 | v_10 | v_1908;
assign x_2418 = ~v_664 | ~v_1907 | v_662;
assign x_2419 = ~v_664 | ~v_71 | ~v_9 | v_11 | v_1907;
assign x_2420 = ~v_664 | ~v_1906 | v_661;
assign x_2421 = ~v_664 | ~v_72 | ~v_9 | v_12 | v_1906;
assign x_2422 = ~v_664 | ~v_1905 | v_660;
assign x_2423 = ~v_664 | ~v_73 | ~v_9 | v_13 | v_1905;
assign x_2424 = ~v_664 | ~v_1904 | v_659;
assign x_2425 = ~v_664 | ~v_74 | ~v_9 | v_14 | v_1904;
assign x_2426 = ~v_664 | ~v_1903 | v_658;
assign x_2427 = ~v_664 | ~v_75 | ~v_9 | v_15 | v_1903;
assign x_2428 = ~v_664 | v_10 | ~v_18 | v_1909;
assign x_2429 = ~v_664 | ~v_10 | v_18 | v_1914 | v_1913 | v_1912 | v_1911 | v_1910;
assign x_2430 = ~v_664 | ~v_1909 | v_657;
assign x_2431 = ~v_664 | ~v_70 | ~v_9 | v_10 | v_1909;
assign x_2432 = ~v_664 | ~v_1914 | v_656;
assign x_2433 = ~v_664 | ~v_76 | ~v_10 | v_11 | v_1914;
assign x_2434 = ~v_664 | ~v_1913 | v_655;
assign x_2435 = ~v_664 | ~v_77 | ~v_10 | v_12 | v_1913;
assign x_2436 = ~v_664 | ~v_1912 | v_654;
assign x_2437 = ~v_664 | ~v_78 | ~v_10 | v_13 | v_1912;
assign x_2438 = ~v_664 | ~v_1911 | v_653;
assign x_2439 = ~v_664 | ~v_79 | ~v_10 | v_14 | v_1911;
assign x_2440 = ~v_664 | ~v_1910 | v_652;
assign x_2441 = ~v_664 | ~v_80 | ~v_10 | v_15 | v_1910;
assign x_2442 = ~v_664 | v_11 | ~v_19 | v_1916 | v_1915;
assign x_2443 = ~v_664 | ~v_11 | v_19 | v_1920 | v_1919 | v_1918 | v_1917;
assign x_2444 = ~v_664 | ~v_1916 | v_651;
assign x_2445 = ~v_664 | ~v_71 | ~v_9 | v_11 | v_1916;
assign x_2446 = ~v_664 | ~v_1915 | v_650;
assign x_2447 = ~v_664 | ~v_76 | ~v_10 | v_11 | v_1915;
assign x_2448 = ~v_664 | ~v_1920 | v_649;
assign x_2449 = ~v_664 | ~v_81 | ~v_11 | v_12 | v_1920;
assign x_2450 = ~v_664 | ~v_1919 | v_648;
assign x_2451 = ~v_664 | ~v_82 | ~v_11 | v_13 | v_1919;
assign x_2452 = ~v_664 | ~v_1918 | v_647;
assign x_2453 = ~v_664 | ~v_83 | ~v_11 | v_14 | v_1918;
assign x_2454 = ~v_664 | ~v_1917 | v_646;
assign x_2455 = ~v_664 | ~v_84 | ~v_11 | v_15 | v_1917;
assign x_2456 = ~v_664 | v_12 | ~v_20 | v_1923 | v_1922 | v_1921;
assign x_2457 = ~v_664 | ~v_12 | v_20 | v_1926 | v_1925 | v_1924;
assign x_2458 = ~v_664 | ~v_1923 | v_645;
assign x_2459 = ~v_664 | ~v_72 | ~v_9 | v_12 | v_1923;
assign x_2460 = ~v_664 | ~v_1922 | v_644;
assign x_2461 = ~v_664 | ~v_77 | ~v_10 | v_12 | v_1922;
assign x_2462 = ~v_664 | ~v_1921 | v_643;
assign x_2463 = ~v_664 | ~v_81 | ~v_11 | v_12 | v_1921;
assign x_2464 = ~v_664 | ~v_1926 | v_642;
assign x_2465 = ~v_664 | ~v_85 | ~v_12 | v_13 | v_1926;
assign x_2466 = ~v_664 | ~v_1925 | v_641;
assign x_2467 = ~v_664 | ~v_86 | ~v_12 | v_14 | v_1925;
assign x_2468 = ~v_664 | ~v_1924 | v_640;
assign x_2469 = ~v_664 | ~v_87 | ~v_12 | v_15 | v_1924;
assign x_2470 = ~v_664 | v_13 | ~v_21 | v_1930 | v_1929 | v_1928 | v_1927;
assign x_2471 = ~v_664 | ~v_13 | v_21 | v_1932 | v_1931;
assign x_2472 = ~v_664 | ~v_1930 | v_639;
assign x_2473 = ~v_664 | ~v_73 | ~v_9 | v_13 | v_1930;
assign x_2474 = ~v_664 | ~v_1929 | v_638;
assign x_2475 = ~v_664 | ~v_78 | ~v_10 | v_13 | v_1929;
assign x_2476 = ~v_664 | ~v_1928 | v_637;
assign x_2477 = ~v_664 | ~v_82 | ~v_11 | v_13 | v_1928;
assign x_2478 = ~v_664 | ~v_1927 | v_636;
assign x_2479 = ~v_664 | ~v_85 | ~v_12 | v_13 | v_1927;
assign x_2480 = ~v_664 | ~v_1932 | v_635;
assign x_2481 = ~v_664 | ~v_88 | ~v_13 | v_14 | v_1932;
assign x_2482 = ~v_664 | ~v_1931 | v_634;
assign x_2483 = ~v_664 | ~v_89 | ~v_13 | v_15 | v_1931;
assign x_2484 = ~v_664 | v_14 | ~v_22 | v_1937 | v_1936 | v_1935 | v_1934 | v_1933;
assign x_2485 = ~v_664 | ~v_14 | v_22 | v_1938;
assign x_2486 = ~v_664 | ~v_1937 | v_633;
assign x_2487 = ~v_664 | ~v_74 | ~v_9 | v_14 | v_1937;
assign x_2488 = ~v_664 | ~v_1936 | v_632;
assign x_2489 = ~v_664 | ~v_79 | ~v_10 | v_14 | v_1936;
assign x_2490 = ~v_664 | ~v_1935 | v_631;
assign x_2491 = ~v_664 | ~v_83 | ~v_11 | v_14 | v_1935;
assign x_2492 = ~v_664 | ~v_1934 | v_630;
assign x_2493 = ~v_664 | ~v_86 | ~v_12 | v_14 | v_1934;
assign x_2494 = ~v_664 | ~v_1933 | v_629;
assign x_2495 = ~v_664 | ~v_88 | ~v_13 | v_14 | v_1933;
assign x_2496 = ~v_664 | ~v_1938 | v_628;
assign x_2497 = ~v_664 | ~v_90 | ~v_14 | v_15 | v_1938;
assign x_2498 = ~v_664 | v_15 | ~v_23 | v_1944 | v_1943 | v_1942 | v_1941 | v_1940 | v_1939;
assign x_2499 = ~v_664 | ~v_15 | v_23;
assign x_2500 = ~v_664 | ~v_1944 | v_627;
assign x_2501 = ~v_664 | ~v_75 | ~v_9 | v_15 | v_1944;
assign x_2502 = ~v_664 | ~v_1943 | v_626;
assign x_2503 = ~v_664 | ~v_80 | ~v_10 | v_15 | v_1943;
assign x_2504 = ~v_664 | ~v_1942 | v_625;
assign x_2505 = ~v_664 | ~v_84 | ~v_11 | v_15 | v_1942;
assign x_2506 = ~v_664 | ~v_1941 | v_624;
assign x_2507 = ~v_664 | ~v_87 | ~v_12 | v_15 | v_1941;
assign x_2508 = ~v_664 | ~v_1940 | v_623;
assign x_2509 = ~v_664 | ~v_89 | ~v_13 | v_15 | v_1940;
assign x_2510 = ~v_664 | ~v_1939 | v_622;
assign x_2511 = ~v_664 | ~v_90 | ~v_14 | v_15 | v_1939;
assign x_2512 = ~v_664 | v_16 | ~v_24;
assign x_2513 = ~v_664 | ~v_16 | v_24;
assign x_2514 = ~v_664 | v_620 | v_621;
assign x_2515 = ~v_664 | v_618 | v_619;
assign x_2516 = ~v_664 | v_616 | v_617;
assign x_2517 = ~v_664 | v_614 | v_615;
assign x_2518 = ~v_664 | v_612 | v_613;
assign x_2519 = ~v_664 | v_610 | v_611;
assign x_2520 = ~v_664 | v_608 | v_609;
assign x_2521 = ~v_664 | v_606 | v_607;
assign x_2522 = ~v_664 | v_604 | v_605;
assign x_2523 = ~v_664 | v_602 | v_603;
assign x_2524 = ~v_664 | v_600 | v_601;
assign x_2525 = ~v_664 | v_598 | v_599;
assign x_2526 = ~v_664 | v_596 | v_597;
assign x_2527 = ~v_664 | v_594 | v_595;
assign x_2528 = ~v_664 | v_592 | v_593;
assign x_2529 = ~v_664 | v_590 | v_591;
assign x_2530 = ~v_664 | v_588 | v_589;
assign x_2531 = ~v_664 | v_586 | v_587;
assign x_2532 = ~v_664 | v_584 | v_585;
assign x_2533 = ~v_664 | v_582 | v_583;
assign x_2534 = ~v_664 | v_580 | v_581;
assign x_2535 = ~v_664 | v_558;
assign x_2536 = ~v_663 | v_70;
assign x_2537 = ~v_663 | v_9;
assign x_2538 = ~v_663 | ~v_10;
assign x_2539 = ~v_662 | v_71;
assign x_2540 = ~v_662 | v_9;
assign x_2541 = ~v_662 | ~v_11;
assign x_2542 = ~v_661 | v_72;
assign x_2543 = ~v_661 | v_9;
assign x_2544 = ~v_661 | ~v_12;
assign x_2545 = ~v_660 | v_73;
assign x_2546 = ~v_660 | v_9;
assign x_2547 = ~v_660 | ~v_13;
assign x_2548 = ~v_659 | v_74;
assign x_2549 = ~v_659 | v_9;
assign x_2550 = ~v_659 | ~v_14;
assign x_2551 = ~v_658 | v_75;
assign x_2552 = ~v_658 | v_9;
assign x_2553 = ~v_658 | ~v_15;
assign x_2554 = ~v_657 | v_70;
assign x_2555 = ~v_657 | v_9;
assign x_2556 = ~v_657 | ~v_10;
assign x_2557 = ~v_656 | v_76;
assign x_2558 = ~v_656 | v_10;
assign x_2559 = ~v_656 | ~v_11;
assign x_2560 = ~v_655 | v_77;
assign x_2561 = ~v_655 | v_10;
assign x_2562 = ~v_655 | ~v_12;
assign x_2563 = ~v_654 | v_78;
assign x_2564 = ~v_654 | v_10;
assign x_2565 = ~v_654 | ~v_13;
assign x_2566 = ~v_653 | v_79;
assign x_2567 = ~v_653 | v_10;
assign x_2568 = ~v_653 | ~v_14;
assign x_2569 = ~v_652 | v_80;
assign x_2570 = ~v_652 | v_10;
assign x_2571 = ~v_652 | ~v_15;
assign x_2572 = ~v_651 | v_71;
assign x_2573 = ~v_651 | v_9;
assign x_2574 = ~v_651 | ~v_11;
assign x_2575 = ~v_650 | v_76;
assign x_2576 = ~v_650 | v_10;
assign x_2577 = ~v_650 | ~v_11;
assign x_2578 = ~v_649 | v_81;
assign x_2579 = ~v_649 | v_11;
assign x_2580 = ~v_649 | ~v_12;
assign x_2581 = ~v_648 | v_82;
assign x_2582 = ~v_648 | v_11;
assign x_2583 = ~v_648 | ~v_13;
assign x_2584 = ~v_647 | v_83;
assign x_2585 = ~v_647 | v_11;
assign x_2586 = ~v_647 | ~v_14;
assign x_2587 = ~v_646 | v_84;
assign x_2588 = ~v_646 | v_11;
assign x_2589 = ~v_646 | ~v_15;
assign x_2590 = ~v_645 | v_72;
assign x_2591 = ~v_645 | v_9;
assign x_2592 = ~v_645 | ~v_12;
assign x_2593 = ~v_644 | v_77;
assign x_2594 = ~v_644 | v_10;
assign x_2595 = ~v_644 | ~v_12;
assign x_2596 = ~v_643 | v_81;
assign x_2597 = ~v_643 | v_11;
assign x_2598 = ~v_643 | ~v_12;
assign x_2599 = ~v_642 | v_85;
assign x_2600 = ~v_642 | v_12;
assign x_2601 = ~v_642 | ~v_13;
assign x_2602 = ~v_641 | v_86;
assign x_2603 = ~v_641 | v_12;
assign x_2604 = ~v_641 | ~v_14;
assign x_2605 = ~v_640 | v_87;
assign x_2606 = ~v_640 | v_12;
assign x_2607 = ~v_640 | ~v_15;
assign x_2608 = ~v_639 | v_73;
assign x_2609 = ~v_639 | v_9;
assign x_2610 = ~v_639 | ~v_13;
assign x_2611 = ~v_638 | v_78;
assign x_2612 = ~v_638 | v_10;
assign x_2613 = ~v_638 | ~v_13;
assign x_2614 = ~v_637 | v_82;
assign x_2615 = ~v_637 | v_11;
assign x_2616 = ~v_637 | ~v_13;
assign x_2617 = ~v_636 | v_85;
assign x_2618 = ~v_636 | v_12;
assign x_2619 = ~v_636 | ~v_13;
assign x_2620 = ~v_635 | v_88;
assign x_2621 = ~v_635 | v_13;
assign x_2622 = ~v_635 | ~v_14;
assign x_2623 = ~v_634 | v_89;
assign x_2624 = ~v_634 | v_13;
assign x_2625 = ~v_634 | ~v_15;
assign x_2626 = ~v_633 | v_74;
assign x_2627 = ~v_633 | v_9;
assign x_2628 = ~v_633 | ~v_14;
assign x_2629 = ~v_632 | v_79;
assign x_2630 = ~v_632 | v_10;
assign x_2631 = ~v_632 | ~v_14;
assign x_2632 = ~v_631 | v_83;
assign x_2633 = ~v_631 | v_11;
assign x_2634 = ~v_631 | ~v_14;
assign x_2635 = ~v_630 | v_86;
assign x_2636 = ~v_630 | v_12;
assign x_2637 = ~v_630 | ~v_14;
assign x_2638 = ~v_629 | v_88;
assign x_2639 = ~v_629 | v_13;
assign x_2640 = ~v_629 | ~v_14;
assign x_2641 = ~v_628 | v_90;
assign x_2642 = ~v_628 | v_14;
assign x_2643 = ~v_628 | ~v_15;
assign x_2644 = ~v_627 | v_75;
assign x_2645 = ~v_627 | v_9;
assign x_2646 = ~v_627 | ~v_15;
assign x_2647 = ~v_626 | v_80;
assign x_2648 = ~v_626 | v_10;
assign x_2649 = ~v_626 | ~v_15;
assign x_2650 = ~v_625 | v_84;
assign x_2651 = ~v_625 | v_11;
assign x_2652 = ~v_625 | ~v_15;
assign x_2653 = ~v_624 | v_87;
assign x_2654 = ~v_624 | v_12;
assign x_2655 = ~v_624 | ~v_15;
assign x_2656 = ~v_623 | v_89;
assign x_2657 = ~v_623 | v_13;
assign x_2658 = ~v_623 | ~v_15;
assign x_2659 = ~v_622 | v_90;
assign x_2660 = ~v_622 | v_14;
assign x_2661 = ~v_622 | ~v_15;
assign x_2662 = ~v_620 | ~v_70 | ~v_9 | v_10;
assign x_2663 = ~v_621 | ~v_17;
assign x_2664 = ~v_621 | v_18;
assign x_2665 = ~v_618 | ~v_71 | ~v_9 | v_11;
assign x_2666 = ~v_619 | ~v_17;
assign x_2667 = ~v_619 | v_19;
assign x_2668 = ~v_616 | ~v_72 | ~v_9 | v_12;
assign x_2669 = ~v_617 | ~v_17;
assign x_2670 = ~v_617 | v_20;
assign x_2671 = ~v_614 | ~v_73 | ~v_9 | v_13;
assign x_2672 = ~v_615 | ~v_17;
assign x_2673 = ~v_615 | v_21;
assign x_2674 = ~v_612 | ~v_74 | ~v_9 | v_14;
assign x_2675 = ~v_613 | ~v_17;
assign x_2676 = ~v_613 | v_22;
assign x_2677 = ~v_610 | ~v_75 | ~v_9 | v_15;
assign x_2678 = ~v_611 | ~v_17;
assign x_2679 = ~v_611 | v_23;
assign x_2680 = ~v_608 | ~v_76 | ~v_10 | v_11;
assign x_2681 = ~v_609 | ~v_18;
assign x_2682 = ~v_609 | v_19;
assign x_2683 = ~v_606 | ~v_77 | ~v_10 | v_12;
assign x_2684 = ~v_607 | ~v_18;
assign x_2685 = ~v_607 | v_20;
assign x_2686 = ~v_604 | ~v_78 | ~v_10 | v_13;
assign x_2687 = ~v_605 | ~v_18;
assign x_2688 = ~v_605 | v_21;
assign x_2689 = ~v_602 | ~v_79 | ~v_10 | v_14;
assign x_2690 = ~v_603 | ~v_18;
assign x_2691 = ~v_603 | v_22;
assign x_2692 = ~v_600 | ~v_80 | ~v_10 | v_15;
assign x_2693 = ~v_601 | ~v_18;
assign x_2694 = ~v_601 | v_23;
assign x_2695 = ~v_598 | ~v_81 | ~v_11 | v_12;
assign x_2696 = ~v_599 | ~v_19;
assign x_2697 = ~v_599 | v_20;
assign x_2698 = ~v_596 | ~v_82 | ~v_11 | v_13;
assign x_2699 = ~v_597 | ~v_19;
assign x_2700 = ~v_597 | v_21;
assign x_2701 = ~v_594 | ~v_83 | ~v_11 | v_14;
assign x_2702 = ~v_595 | ~v_19;
assign x_2703 = ~v_595 | v_22;
assign x_2704 = ~v_592 | ~v_84 | ~v_11 | v_15;
assign x_2705 = ~v_593 | ~v_19;
assign x_2706 = ~v_593 | v_23;
assign x_2707 = ~v_590 | ~v_85 | ~v_12 | v_13;
assign x_2708 = ~v_591 | ~v_20;
assign x_2709 = ~v_591 | v_21;
assign x_2710 = ~v_588 | ~v_86 | ~v_12 | v_14;
assign x_2711 = ~v_589 | ~v_20;
assign x_2712 = ~v_589 | v_22;
assign x_2713 = ~v_586 | ~v_87 | ~v_12 | v_15;
assign x_2714 = ~v_587 | ~v_20;
assign x_2715 = ~v_587 | v_23;
assign x_2716 = ~v_584 | ~v_88 | ~v_13 | v_14;
assign x_2717 = ~v_585 | ~v_21;
assign x_2718 = ~v_585 | v_22;
assign x_2719 = ~v_582 | ~v_89 | ~v_13 | v_15;
assign x_2720 = ~v_583 | ~v_21;
assign x_2721 = ~v_583 | v_23;
assign x_2722 = ~v_580 | ~v_90 | ~v_14 | v_15;
assign x_2723 = ~v_581 | ~v_22;
assign x_2724 = ~v_581 | v_23;
assign x_2725 = ~v_558 | v_17 | ~v_25;
assign x_2726 = ~v_558 | ~v_17 | v_25 | v_2010 | v_2009 | v_2008 | v_2007 | v_2006 | v_2005;
assign x_2727 = ~v_558 | ~v_2010 | v_557;
assign x_2728 = ~v_558 | ~v_91 | ~v_17 | v_18 | v_2010;
assign x_2729 = ~v_558 | ~v_2009 | v_556;
assign x_2730 = ~v_558 | ~v_92 | ~v_17 | v_19 | v_2009;
assign x_2731 = ~v_558 | ~v_2008 | v_555;
assign x_2732 = ~v_558 | ~v_93 | ~v_17 | v_20 | v_2008;
assign x_2733 = ~v_558 | ~v_2007 | v_554;
assign x_2734 = ~v_558 | ~v_94 | ~v_17 | v_21 | v_2007;
assign x_2735 = ~v_558 | ~v_2006 | v_553;
assign x_2736 = ~v_558 | ~v_95 | ~v_17 | v_22 | v_2006;
assign x_2737 = ~v_558 | ~v_2005 | v_552;
assign x_2738 = ~v_558 | ~v_96 | ~v_17 | v_23 | v_2005;
assign x_2739 = ~v_558 | v_18 | ~v_26 | v_2011;
assign x_2740 = ~v_558 | ~v_18 | v_26 | v_2016 | v_2015 | v_2014 | v_2013 | v_2012;
assign x_2741 = ~v_558 | ~v_2011 | v_551;
assign x_2742 = ~v_558 | ~v_91 | ~v_17 | v_18 | v_2011;
assign x_2743 = ~v_558 | ~v_2016 | v_550;
assign x_2744 = ~v_558 | ~v_97 | ~v_18 | v_19 | v_2016;
assign x_2745 = ~v_558 | ~v_2015 | v_549;
assign x_2746 = ~v_558 | ~v_98 | ~v_18 | v_20 | v_2015;
assign x_2747 = ~v_558 | ~v_2014 | v_548;
assign x_2748 = ~v_558 | ~v_99 | ~v_18 | v_21 | v_2014;
assign x_2749 = ~v_558 | ~v_2013 | v_547;
assign x_2750 = ~v_558 | ~v_100 | ~v_18 | v_22 | v_2013;
assign x_2751 = ~v_558 | ~v_2012 | v_546;
assign x_2752 = ~v_558 | ~v_101 | ~v_18 | v_23 | v_2012;
assign x_2753 = ~v_558 | v_19 | ~v_27 | v_2018 | v_2017;
assign x_2754 = ~v_558 | ~v_19 | v_27 | v_2022 | v_2021 | v_2020 | v_2019;
assign x_2755 = ~v_558 | ~v_2018 | v_545;
assign x_2756 = ~v_558 | ~v_92 | ~v_17 | v_19 | v_2018;
assign x_2757 = ~v_558 | ~v_2017 | v_544;
assign x_2758 = ~v_558 | ~v_97 | ~v_18 | v_19 | v_2017;
assign x_2759 = ~v_558 | ~v_2022 | v_543;
assign x_2760 = ~v_558 | ~v_102 | ~v_19 | v_20 | v_2022;
assign x_2761 = ~v_558 | ~v_2021 | v_542;
assign x_2762 = ~v_558 | ~v_103 | ~v_19 | v_21 | v_2021;
assign x_2763 = ~v_558 | ~v_2020 | v_541;
assign x_2764 = ~v_558 | ~v_104 | ~v_19 | v_22 | v_2020;
assign x_2765 = ~v_558 | ~v_2019 | v_540;
assign x_2766 = ~v_558 | ~v_105 | ~v_19 | v_23 | v_2019;
assign x_2767 = ~v_558 | v_20 | ~v_28 | v_2025 | v_2024 | v_2023;
assign x_2768 = ~v_558 | ~v_20 | v_28 | v_2028 | v_2027 | v_2026;
assign x_2769 = ~v_558 | ~v_2025 | v_539;
assign x_2770 = ~v_558 | ~v_93 | ~v_17 | v_20 | v_2025;
assign x_2771 = ~v_558 | ~v_2024 | v_538;
assign x_2772 = ~v_558 | ~v_98 | ~v_18 | v_20 | v_2024;
assign x_2773 = ~v_558 | ~v_2023 | v_537;
assign x_2774 = ~v_558 | ~v_102 | ~v_19 | v_20 | v_2023;
assign x_2775 = ~v_558 | ~v_2028 | v_536;
assign x_2776 = ~v_558 | ~v_106 | ~v_20 | v_21 | v_2028;
assign x_2777 = ~v_558 | ~v_2027 | v_535;
assign x_2778 = ~v_558 | ~v_107 | ~v_20 | v_22 | v_2027;
assign x_2779 = ~v_558 | ~v_2026 | v_534;
assign x_2780 = ~v_558 | ~v_108 | ~v_20 | v_23 | v_2026;
assign x_2781 = ~v_558 | v_21 | ~v_29 | v_2032 | v_2031 | v_2030 | v_2029;
assign x_2782 = ~v_558 | ~v_21 | v_29 | v_2034 | v_2033;
assign x_2783 = ~v_558 | ~v_2032 | v_533;
assign x_2784 = ~v_558 | ~v_94 | ~v_17 | v_21 | v_2032;
assign x_2785 = ~v_558 | ~v_2031 | v_532;
assign x_2786 = ~v_558 | ~v_99 | ~v_18 | v_21 | v_2031;
assign x_2787 = ~v_558 | ~v_2030 | v_531;
assign x_2788 = ~v_558 | ~v_103 | ~v_19 | v_21 | v_2030;
assign x_2789 = ~v_558 | ~v_2029 | v_530;
assign x_2790 = ~v_558 | ~v_106 | ~v_20 | v_21 | v_2029;
assign x_2791 = ~v_558 | ~v_2034 | v_529;
assign x_2792 = ~v_558 | ~v_109 | ~v_21 | v_22 | v_2034;
assign x_2793 = ~v_558 | ~v_2033 | v_528;
assign x_2794 = ~v_558 | ~v_110 | ~v_21 | v_23 | v_2033;
assign x_2795 = ~v_558 | v_22 | ~v_30 | v_2039 | v_2038 | v_2037 | v_2036 | v_2035;
assign x_2796 = ~v_558 | ~v_22 | v_30 | v_2040;
assign x_2797 = ~v_558 | ~v_2039 | v_527;
assign x_2798 = ~v_558 | ~v_95 | ~v_17 | v_22 | v_2039;
assign x_2799 = ~v_558 | ~v_2038 | v_526;
assign x_2800 = ~v_558 | ~v_100 | ~v_18 | v_22 | v_2038;
assign x_2801 = ~v_558 | ~v_2037 | v_525;
assign x_2802 = ~v_558 | ~v_104 | ~v_19 | v_22 | v_2037;
assign x_2803 = ~v_558 | ~v_2036 | v_524;
assign x_2804 = ~v_558 | ~v_107 | ~v_20 | v_22 | v_2036;
assign x_2805 = ~v_558 | ~v_2035 | v_523;
assign x_2806 = ~v_558 | ~v_109 | ~v_21 | v_22 | v_2035;
assign x_2807 = ~v_558 | ~v_2040 | v_522;
assign x_2808 = ~v_558 | ~v_111 | ~v_22 | v_23 | v_2040;
assign x_2809 = ~v_558 | v_23 | ~v_31 | v_2046 | v_2045 | v_2044 | v_2043 | v_2042 | v_2041;
assign x_2810 = ~v_558 | ~v_23 | v_31;
assign x_2811 = ~v_558 | ~v_2046 | v_521;
assign x_2812 = ~v_558 | ~v_96 | ~v_17 | v_23 | v_2046;
assign x_2813 = ~v_558 | ~v_2045 | v_520;
assign x_2814 = ~v_558 | ~v_101 | ~v_18 | v_23 | v_2045;
assign x_2815 = ~v_558 | ~v_2044 | v_519;
assign x_2816 = ~v_558 | ~v_105 | ~v_19 | v_23 | v_2044;
assign x_2817 = ~v_558 | ~v_2043 | v_518;
assign x_2818 = ~v_558 | ~v_108 | ~v_20 | v_23 | v_2043;
assign x_2819 = ~v_558 | ~v_2042 | v_517;
assign x_2820 = ~v_558 | ~v_110 | ~v_21 | v_23 | v_2042;
assign x_2821 = ~v_558 | ~v_2041 | v_516;
assign x_2822 = ~v_558 | ~v_111 | ~v_22 | v_23 | v_2041;
assign x_2823 = ~v_558 | v_24 | ~v_32;
assign x_2824 = ~v_558 | ~v_24 | v_32;
assign x_2825 = ~v_558 | v_514 | v_515;
assign x_2826 = ~v_558 | v_512 | v_513;
assign x_2827 = ~v_558 | v_510 | v_511;
assign x_2828 = ~v_558 | v_508 | v_509;
assign x_2829 = ~v_558 | v_506 | v_507;
assign x_2830 = ~v_558 | v_504 | v_505;
assign x_2831 = ~v_558 | v_502 | v_503;
assign x_2832 = ~v_558 | v_500 | v_501;
assign x_2833 = ~v_558 | v_498 | v_499;
assign x_2834 = ~v_558 | v_496 | v_497;
assign x_2835 = ~v_558 | v_494 | v_495;
assign x_2836 = ~v_558 | v_492 | v_493;
assign x_2837 = ~v_558 | v_490 | v_491;
assign x_2838 = ~v_558 | v_488 | v_489;
assign x_2839 = ~v_558 | v_486 | v_487;
assign x_2840 = ~v_558 | v_484 | v_485;
assign x_2841 = ~v_558 | v_482 | v_483;
assign x_2842 = ~v_558 | v_480 | v_481;
assign x_2843 = ~v_558 | v_478 | v_479;
assign x_2844 = ~v_558 | v_476 | v_477;
assign x_2845 = ~v_558 | v_474 | v_475;
assign x_2846 = ~v_558 | v_452;
assign x_2847 = ~v_557 | v_91;
assign x_2848 = ~v_557 | v_17;
assign x_2849 = ~v_557 | ~v_18;
assign x_2850 = ~v_556 | v_92;
assign x_2851 = ~v_556 | v_17;
assign x_2852 = ~v_556 | ~v_19;
assign x_2853 = ~v_555 | v_93;
assign x_2854 = ~v_555 | v_17;
assign x_2855 = ~v_555 | ~v_20;
assign x_2856 = ~v_554 | v_94;
assign x_2857 = ~v_554 | v_17;
assign x_2858 = ~v_554 | ~v_21;
assign x_2859 = ~v_553 | v_95;
assign x_2860 = ~v_553 | v_17;
assign x_2861 = ~v_553 | ~v_22;
assign x_2862 = ~v_552 | v_96;
assign x_2863 = ~v_552 | v_17;
assign x_2864 = ~v_552 | ~v_23;
assign x_2865 = ~v_551 | v_91;
assign x_2866 = ~v_551 | v_17;
assign x_2867 = ~v_551 | ~v_18;
assign x_2868 = ~v_550 | v_97;
assign x_2869 = ~v_550 | v_18;
assign x_2870 = ~v_550 | ~v_19;
assign x_2871 = ~v_549 | v_98;
assign x_2872 = ~v_549 | v_18;
assign x_2873 = ~v_549 | ~v_20;
assign x_2874 = ~v_548 | v_99;
assign x_2875 = ~v_548 | v_18;
assign x_2876 = ~v_548 | ~v_21;
assign x_2877 = ~v_547 | v_100;
assign x_2878 = ~v_547 | v_18;
assign x_2879 = ~v_547 | ~v_22;
assign x_2880 = ~v_546 | v_101;
assign x_2881 = ~v_546 | v_18;
assign x_2882 = ~v_546 | ~v_23;
assign x_2883 = ~v_545 | v_92;
assign x_2884 = ~v_545 | v_17;
assign x_2885 = ~v_545 | ~v_19;
assign x_2886 = ~v_544 | v_97;
assign x_2887 = ~v_544 | v_18;
assign x_2888 = ~v_544 | ~v_19;
assign x_2889 = ~v_543 | v_102;
assign x_2890 = ~v_543 | v_19;
assign x_2891 = ~v_543 | ~v_20;
assign x_2892 = ~v_542 | v_103;
assign x_2893 = ~v_542 | v_19;
assign x_2894 = ~v_542 | ~v_21;
assign x_2895 = ~v_541 | v_104;
assign x_2896 = ~v_541 | v_19;
assign x_2897 = ~v_541 | ~v_22;
assign x_2898 = ~v_540 | v_105;
assign x_2899 = ~v_540 | v_19;
assign x_2900 = ~v_540 | ~v_23;
assign x_2901 = ~v_539 | v_93;
assign x_2902 = ~v_539 | v_17;
assign x_2903 = ~v_539 | ~v_20;
assign x_2904 = ~v_538 | v_98;
assign x_2905 = ~v_538 | v_18;
assign x_2906 = ~v_538 | ~v_20;
assign x_2907 = ~v_537 | v_102;
assign x_2908 = ~v_537 | v_19;
assign x_2909 = ~v_537 | ~v_20;
assign x_2910 = ~v_536 | v_106;
assign x_2911 = ~v_536 | v_20;
assign x_2912 = ~v_536 | ~v_21;
assign x_2913 = ~v_535 | v_107;
assign x_2914 = ~v_535 | v_20;
assign x_2915 = ~v_535 | ~v_22;
assign x_2916 = ~v_534 | v_108;
assign x_2917 = ~v_534 | v_20;
assign x_2918 = ~v_534 | ~v_23;
assign x_2919 = ~v_533 | v_94;
assign x_2920 = ~v_533 | v_17;
assign x_2921 = ~v_533 | ~v_21;
assign x_2922 = ~v_532 | v_99;
assign x_2923 = ~v_532 | v_18;
assign x_2924 = ~v_532 | ~v_21;
assign x_2925 = ~v_531 | v_103;
assign x_2926 = ~v_531 | v_19;
assign x_2927 = ~v_531 | ~v_21;
assign x_2928 = ~v_530 | v_106;
assign x_2929 = ~v_530 | v_20;
assign x_2930 = ~v_530 | ~v_21;
assign x_2931 = ~v_529 | v_109;
assign x_2932 = ~v_529 | v_21;
assign x_2933 = ~v_529 | ~v_22;
assign x_2934 = ~v_528 | v_110;
assign x_2935 = ~v_528 | v_21;
assign x_2936 = ~v_528 | ~v_23;
assign x_2937 = ~v_527 | v_95;
assign x_2938 = ~v_527 | v_17;
assign x_2939 = ~v_527 | ~v_22;
assign x_2940 = ~v_526 | v_100;
assign x_2941 = ~v_526 | v_18;
assign x_2942 = ~v_526 | ~v_22;
assign x_2943 = ~v_525 | v_104;
assign x_2944 = ~v_525 | v_19;
assign x_2945 = ~v_525 | ~v_22;
assign x_2946 = ~v_524 | v_107;
assign x_2947 = ~v_524 | v_20;
assign x_2948 = ~v_524 | ~v_22;
assign x_2949 = ~v_523 | v_109;
assign x_2950 = ~v_523 | v_21;
assign x_2951 = ~v_523 | ~v_22;
assign x_2952 = ~v_522 | v_111;
assign x_2953 = ~v_522 | v_22;
assign x_2954 = ~v_522 | ~v_23;
assign x_2955 = ~v_521 | v_96;
assign x_2956 = ~v_521 | v_17;
assign x_2957 = ~v_521 | ~v_23;
assign x_2958 = ~v_520 | v_101;
assign x_2959 = ~v_520 | v_18;
assign x_2960 = ~v_520 | ~v_23;
assign x_2961 = ~v_519 | v_105;
assign x_2962 = ~v_519 | v_19;
assign x_2963 = ~v_519 | ~v_23;
assign x_2964 = ~v_518 | v_108;
assign x_2965 = ~v_518 | v_20;
assign x_2966 = ~v_518 | ~v_23;
assign x_2967 = ~v_517 | v_110;
assign x_2968 = ~v_517 | v_21;
assign x_2969 = ~v_517 | ~v_23;
assign x_2970 = ~v_516 | v_111;
assign x_2971 = ~v_516 | v_22;
assign x_2972 = ~v_516 | ~v_23;
assign x_2973 = ~v_514 | ~v_91 | ~v_17 | v_18;
assign x_2974 = ~v_515 | ~v_25;
assign x_2975 = ~v_515 | v_26;
assign x_2976 = ~v_512 | ~v_92 | ~v_17 | v_19;
assign x_2977 = ~v_513 | ~v_25;
assign x_2978 = ~v_513 | v_27;
assign x_2979 = ~v_510 | ~v_93 | ~v_17 | v_20;
assign x_2980 = ~v_511 | ~v_25;
assign x_2981 = ~v_511 | v_28;
assign x_2982 = ~v_508 | ~v_94 | ~v_17 | v_21;
assign x_2983 = ~v_509 | ~v_25;
assign x_2984 = ~v_509 | v_29;
assign x_2985 = ~v_506 | ~v_95 | ~v_17 | v_22;
assign x_2986 = ~v_507 | ~v_25;
assign x_2987 = ~v_507 | v_30;
assign x_2988 = ~v_504 | ~v_96 | ~v_17 | v_23;
assign x_2989 = ~v_505 | ~v_25;
assign x_2990 = ~v_505 | v_31;
assign x_2991 = ~v_502 | ~v_97 | ~v_18 | v_19;
assign x_2992 = ~v_503 | ~v_26;
assign x_2993 = ~v_503 | v_27;
assign x_2994 = ~v_500 | ~v_98 | ~v_18 | v_20;
assign x_2995 = ~v_501 | ~v_26;
assign x_2996 = ~v_501 | v_28;
assign x_2997 = ~v_498 | ~v_99 | ~v_18 | v_21;
assign x_2998 = ~v_499 | ~v_26;
assign x_2999 = ~v_499 | v_29;
assign x_3000 = ~v_496 | ~v_100 | ~v_18 | v_22;
assign x_3001 = ~v_497 | ~v_26;
assign x_3002 = ~v_497 | v_30;
assign x_3003 = ~v_494 | ~v_101 | ~v_18 | v_23;
assign x_3004 = ~v_495 | ~v_26;
assign x_3005 = ~v_495 | v_31;
assign x_3006 = ~v_492 | ~v_102 | ~v_19 | v_20;
assign x_3007 = ~v_493 | ~v_27;
assign x_3008 = ~v_493 | v_28;
assign x_3009 = ~v_490 | ~v_103 | ~v_19 | v_21;
assign x_3010 = ~v_491 | ~v_27;
assign x_3011 = ~v_491 | v_29;
assign x_3012 = ~v_488 | ~v_104 | ~v_19 | v_22;
assign x_3013 = ~v_489 | ~v_27;
assign x_3014 = ~v_489 | v_30;
assign x_3015 = ~v_486 | ~v_105 | ~v_19 | v_23;
assign x_3016 = ~v_487 | ~v_27;
assign x_3017 = ~v_487 | v_31;
assign x_3018 = ~v_484 | ~v_106 | ~v_20 | v_21;
assign x_3019 = ~v_485 | ~v_28;
assign x_3020 = ~v_485 | v_29;
assign x_3021 = ~v_482 | ~v_107 | ~v_20 | v_22;
assign x_3022 = ~v_483 | ~v_28;
assign x_3023 = ~v_483 | v_30;
assign x_3024 = ~v_480 | ~v_108 | ~v_20 | v_23;
assign x_3025 = ~v_481 | ~v_28;
assign x_3026 = ~v_481 | v_31;
assign x_3027 = ~v_478 | ~v_109 | ~v_21 | v_22;
assign x_3028 = ~v_479 | ~v_29;
assign x_3029 = ~v_479 | v_30;
assign x_3030 = ~v_476 | ~v_110 | ~v_21 | v_23;
assign x_3031 = ~v_477 | ~v_29;
assign x_3032 = ~v_477 | v_31;
assign x_3033 = ~v_474 | ~v_111 | ~v_22 | v_23;
assign x_3034 = ~v_475 | ~v_30;
assign x_3035 = ~v_475 | v_31;
assign x_3036 = ~v_452 | v_25 | ~v_33;
assign x_3037 = ~v_452 | ~v_25 | v_33 | v_2112 | v_2111 | v_2110 | v_2109 | v_2108 | v_2107;
assign x_3038 = ~v_452 | ~v_2112 | v_451;
assign x_3039 = ~v_452 | ~v_112 | ~v_25 | v_26 | v_2112;
assign x_3040 = ~v_452 | ~v_2111 | v_450;
assign x_3041 = ~v_452 | ~v_113 | ~v_25 | v_27 | v_2111;
assign x_3042 = ~v_452 | ~v_2110 | v_449;
assign x_3043 = ~v_452 | ~v_114 | ~v_25 | v_28 | v_2110;
assign x_3044 = ~v_452 | ~v_2109 | v_448;
assign x_3045 = ~v_452 | ~v_115 | ~v_25 | v_29 | v_2109;
assign x_3046 = ~v_452 | ~v_2108 | v_447;
assign x_3047 = ~v_452 | ~v_116 | ~v_25 | v_30 | v_2108;
assign x_3048 = ~v_452 | ~v_2107 | v_446;
assign x_3049 = ~v_452 | ~v_117 | ~v_25 | v_31 | v_2107;
assign x_3050 = ~v_452 | v_26 | ~v_34 | v_2113;
assign x_3051 = ~v_452 | ~v_26 | v_34 | v_2118 | v_2117 | v_2116 | v_2115 | v_2114;
assign x_3052 = ~v_452 | ~v_2113 | v_445;
assign x_3053 = ~v_452 | ~v_112 | ~v_25 | v_26 | v_2113;
assign x_3054 = ~v_452 | ~v_2118 | v_444;
assign x_3055 = ~v_452 | ~v_118 | ~v_26 | v_27 | v_2118;
assign x_3056 = ~v_452 | ~v_2117 | v_443;
assign x_3057 = ~v_452 | ~v_119 | ~v_26 | v_28 | v_2117;
assign x_3058 = ~v_452 | ~v_2116 | v_442;
assign x_3059 = ~v_452 | ~v_120 | ~v_26 | v_29 | v_2116;
assign x_3060 = ~v_452 | ~v_2115 | v_441;
assign x_3061 = ~v_452 | ~v_121 | ~v_26 | v_30 | v_2115;
assign x_3062 = ~v_452 | ~v_2114 | v_440;
assign x_3063 = ~v_452 | ~v_122 | ~v_26 | v_31 | v_2114;
assign x_3064 = ~v_452 | v_27 | ~v_35 | v_2120 | v_2119;
assign x_3065 = ~v_452 | ~v_27 | v_35 | v_2124 | v_2123 | v_2122 | v_2121;
assign x_3066 = ~v_452 | ~v_2120 | v_439;
assign x_3067 = ~v_452 | ~v_113 | ~v_25 | v_27 | v_2120;
assign x_3068 = ~v_452 | ~v_2119 | v_438;
assign x_3069 = ~v_452 | ~v_118 | ~v_26 | v_27 | v_2119;
assign x_3070 = ~v_452 | ~v_2124 | v_437;
assign x_3071 = ~v_452 | ~v_123 | ~v_27 | v_28 | v_2124;
assign x_3072 = ~v_452 | ~v_2123 | v_436;
assign x_3073 = ~v_452 | ~v_124 | ~v_27 | v_29 | v_2123;
assign x_3074 = ~v_452 | ~v_2122 | v_435;
assign x_3075 = ~v_452 | ~v_125 | ~v_27 | v_30 | v_2122;
assign x_3076 = ~v_452 | ~v_2121 | v_434;
assign x_3077 = ~v_452 | ~v_126 | ~v_27 | v_31 | v_2121;
assign x_3078 = ~v_452 | v_28 | ~v_36 | v_2127 | v_2126 | v_2125;
assign x_3079 = ~v_452 | ~v_28 | v_36 | v_2130 | v_2129 | v_2128;
assign x_3080 = ~v_452 | ~v_2127 | v_433;
assign x_3081 = ~v_452 | ~v_114 | ~v_25 | v_28 | v_2127;
assign x_3082 = ~v_452 | ~v_2126 | v_432;
assign x_3083 = ~v_452 | ~v_119 | ~v_26 | v_28 | v_2126;
assign x_3084 = ~v_452 | ~v_2125 | v_431;
assign x_3085 = ~v_452 | ~v_123 | ~v_27 | v_28 | v_2125;
assign x_3086 = ~v_452 | ~v_2130 | v_430;
assign x_3087 = ~v_452 | ~v_127 | ~v_28 | v_29 | v_2130;
assign x_3088 = ~v_452 | ~v_2129 | v_429;
assign x_3089 = ~v_452 | ~v_128 | ~v_28 | v_30 | v_2129;
assign x_3090 = ~v_452 | ~v_2128 | v_428;
assign x_3091 = ~v_452 | ~v_129 | ~v_28 | v_31 | v_2128;
assign x_3092 = ~v_452 | v_29 | ~v_37 | v_2134 | v_2133 | v_2132 | v_2131;
assign x_3093 = ~v_452 | ~v_29 | v_37 | v_2136 | v_2135;
assign x_3094 = ~v_452 | ~v_2134 | v_427;
assign x_3095 = ~v_452 | ~v_115 | ~v_25 | v_29 | v_2134;
assign x_3096 = ~v_452 | ~v_2133 | v_426;
assign x_3097 = ~v_452 | ~v_120 | ~v_26 | v_29 | v_2133;
assign x_3098 = ~v_452 | ~v_2132 | v_425;
assign x_3099 = ~v_452 | ~v_124 | ~v_27 | v_29 | v_2132;
assign x_3100 = ~v_452 | ~v_2131 | v_424;
assign x_3101 = ~v_452 | ~v_127 | ~v_28 | v_29 | v_2131;
assign x_3102 = ~v_452 | ~v_2136 | v_423;
assign x_3103 = ~v_452 | ~v_130 | ~v_29 | v_30 | v_2136;
assign x_3104 = ~v_452 | ~v_2135 | v_422;
assign x_3105 = ~v_452 | ~v_131 | ~v_29 | v_31 | v_2135;
assign x_3106 = ~v_452 | v_30 | ~v_38 | v_2141 | v_2140 | v_2139 | v_2138 | v_2137;
assign x_3107 = ~v_452 | ~v_30 | v_38 | v_2142;
assign x_3108 = ~v_452 | ~v_2141 | v_421;
assign x_3109 = ~v_452 | ~v_116 | ~v_25 | v_30 | v_2141;
assign x_3110 = ~v_452 | ~v_2140 | v_420;
assign x_3111 = ~v_452 | ~v_121 | ~v_26 | v_30 | v_2140;
assign x_3112 = ~v_452 | ~v_2139 | v_419;
assign x_3113 = ~v_452 | ~v_125 | ~v_27 | v_30 | v_2139;
assign x_3114 = ~v_452 | ~v_2138 | v_418;
assign x_3115 = ~v_452 | ~v_128 | ~v_28 | v_30 | v_2138;
assign x_3116 = ~v_452 | ~v_2137 | v_417;
assign x_3117 = ~v_452 | ~v_130 | ~v_29 | v_30 | v_2137;
assign x_3118 = ~v_452 | ~v_2142 | v_416;
assign x_3119 = ~v_452 | ~v_132 | ~v_30 | v_31 | v_2142;
assign x_3120 = ~v_452 | v_31 | ~v_39 | v_2148 | v_2147 | v_2146 | v_2145 | v_2144 | v_2143;
assign x_3121 = ~v_452 | ~v_31 | v_39;
assign x_3122 = ~v_452 | ~v_2148 | v_415;
assign x_3123 = ~v_452 | ~v_117 | ~v_25 | v_31 | v_2148;
assign x_3124 = ~v_452 | ~v_2147 | v_414;
assign x_3125 = ~v_452 | ~v_122 | ~v_26 | v_31 | v_2147;
assign x_3126 = ~v_452 | ~v_2146 | v_413;
assign x_3127 = ~v_452 | ~v_126 | ~v_27 | v_31 | v_2146;
assign x_3128 = ~v_452 | ~v_2145 | v_412;
assign x_3129 = ~v_452 | ~v_129 | ~v_28 | v_31 | v_2145;
assign x_3130 = ~v_452 | ~v_2144 | v_411;
assign x_3131 = ~v_452 | ~v_131 | ~v_29 | v_31 | v_2144;
assign x_3132 = ~v_452 | ~v_2143 | v_410;
assign x_3133 = ~v_452 | ~v_132 | ~v_30 | v_31 | v_2143;
assign x_3134 = ~v_452 | v_32 | ~v_40;
assign x_3135 = ~v_452 | ~v_32 | v_40;
assign x_3136 = ~v_452 | v_408 | v_409;
assign x_3137 = ~v_452 | v_406 | v_407;
assign x_3138 = ~v_452 | v_404 | v_405;
assign x_3139 = ~v_452 | v_402 | v_403;
assign x_3140 = ~v_452 | v_400 | v_401;
assign x_3141 = ~v_452 | v_398 | v_399;
assign x_3142 = ~v_452 | v_396 | v_397;
assign x_3143 = ~v_452 | v_394 | v_395;
assign x_3144 = ~v_452 | v_392 | v_393;
assign x_3145 = ~v_452 | v_390 | v_391;
assign x_3146 = ~v_452 | v_388 | v_389;
assign x_3147 = ~v_452 | v_386 | v_387;
assign x_3148 = ~v_452 | v_384 | v_385;
assign x_3149 = ~v_452 | v_382 | v_383;
assign x_3150 = ~v_452 | v_380 | v_381;
assign x_3151 = ~v_452 | v_378 | v_379;
assign x_3152 = ~v_452 | v_376 | v_377;
assign x_3153 = ~v_452 | v_374 | v_375;
assign x_3154 = ~v_452 | v_372 | v_373;
assign x_3155 = ~v_452 | v_370 | v_371;
assign x_3156 = ~v_452 | v_368 | v_369;
assign x_3157 = ~v_452 | v_346;
assign x_3158 = ~v_451 | v_112;
assign x_3159 = ~v_451 | v_25;
assign x_3160 = ~v_451 | ~v_26;
assign x_3161 = ~v_450 | v_113;
assign x_3162 = ~v_450 | v_25;
assign x_3163 = ~v_450 | ~v_27;
assign x_3164 = ~v_449 | v_114;
assign x_3165 = ~v_449 | v_25;
assign x_3166 = ~v_449 | ~v_28;
assign x_3167 = ~v_448 | v_115;
assign x_3168 = ~v_448 | v_25;
assign x_3169 = ~v_448 | ~v_29;
assign x_3170 = ~v_447 | v_116;
assign x_3171 = ~v_447 | v_25;
assign x_3172 = ~v_447 | ~v_30;
assign x_3173 = ~v_446 | v_117;
assign x_3174 = ~v_446 | v_25;
assign x_3175 = ~v_446 | ~v_31;
assign x_3176 = ~v_445 | v_112;
assign x_3177 = ~v_445 | v_25;
assign x_3178 = ~v_445 | ~v_26;
assign x_3179 = ~v_444 | v_118;
assign x_3180 = ~v_444 | v_26;
assign x_3181 = ~v_444 | ~v_27;
assign x_3182 = ~v_443 | v_119;
assign x_3183 = ~v_443 | v_26;
assign x_3184 = ~v_443 | ~v_28;
assign x_3185 = ~v_442 | v_120;
assign x_3186 = ~v_442 | v_26;
assign x_3187 = ~v_442 | ~v_29;
assign x_3188 = ~v_441 | v_121;
assign x_3189 = ~v_441 | v_26;
assign x_3190 = ~v_441 | ~v_30;
assign x_3191 = ~v_440 | v_122;
assign x_3192 = ~v_440 | v_26;
assign x_3193 = ~v_440 | ~v_31;
assign x_3194 = ~v_439 | v_113;
assign x_3195 = ~v_439 | v_25;
assign x_3196 = ~v_439 | ~v_27;
assign x_3197 = ~v_438 | v_118;
assign x_3198 = ~v_438 | v_26;
assign x_3199 = ~v_438 | ~v_27;
assign x_3200 = ~v_437 | v_123;
assign x_3201 = ~v_437 | v_27;
assign x_3202 = ~v_437 | ~v_28;
assign x_3203 = ~v_436 | v_124;
assign x_3204 = ~v_436 | v_27;
assign x_3205 = ~v_436 | ~v_29;
assign x_3206 = ~v_435 | v_125;
assign x_3207 = ~v_435 | v_27;
assign x_3208 = ~v_435 | ~v_30;
assign x_3209 = ~v_434 | v_126;
assign x_3210 = ~v_434 | v_27;
assign x_3211 = ~v_434 | ~v_31;
assign x_3212 = ~v_433 | v_114;
assign x_3213 = ~v_433 | v_25;
assign x_3214 = ~v_433 | ~v_28;
assign x_3215 = ~v_432 | v_119;
assign x_3216 = ~v_432 | v_26;
assign x_3217 = ~v_432 | ~v_28;
assign x_3218 = ~v_431 | v_123;
assign x_3219 = ~v_431 | v_27;
assign x_3220 = ~v_431 | ~v_28;
assign x_3221 = ~v_430 | v_127;
assign x_3222 = ~v_430 | v_28;
assign x_3223 = ~v_430 | ~v_29;
assign x_3224 = ~v_429 | v_128;
assign x_3225 = ~v_429 | v_28;
assign x_3226 = ~v_429 | ~v_30;
assign x_3227 = ~v_428 | v_129;
assign x_3228 = ~v_428 | v_28;
assign x_3229 = ~v_428 | ~v_31;
assign x_3230 = ~v_427 | v_115;
assign x_3231 = ~v_427 | v_25;
assign x_3232 = ~v_427 | ~v_29;
assign x_3233 = ~v_426 | v_120;
assign x_3234 = ~v_426 | v_26;
assign x_3235 = ~v_426 | ~v_29;
assign x_3236 = ~v_425 | v_124;
assign x_3237 = ~v_425 | v_27;
assign x_3238 = ~v_425 | ~v_29;
assign x_3239 = ~v_424 | v_127;
assign x_3240 = ~v_424 | v_28;
assign x_3241 = ~v_424 | ~v_29;
assign x_3242 = ~v_423 | v_130;
assign x_3243 = ~v_423 | v_29;
assign x_3244 = ~v_423 | ~v_30;
assign x_3245 = ~v_422 | v_131;
assign x_3246 = ~v_422 | v_29;
assign x_3247 = ~v_422 | ~v_31;
assign x_3248 = ~v_421 | v_116;
assign x_3249 = ~v_421 | v_25;
assign x_3250 = ~v_421 | ~v_30;
assign x_3251 = ~v_420 | v_121;
assign x_3252 = ~v_420 | v_26;
assign x_3253 = ~v_420 | ~v_30;
assign x_3254 = ~v_419 | v_125;
assign x_3255 = ~v_419 | v_27;
assign x_3256 = ~v_419 | ~v_30;
assign x_3257 = ~v_418 | v_128;
assign x_3258 = ~v_418 | v_28;
assign x_3259 = ~v_418 | ~v_30;
assign x_3260 = ~v_417 | v_130;
assign x_3261 = ~v_417 | v_29;
assign x_3262 = ~v_417 | ~v_30;
assign x_3263 = ~v_416 | v_132;
assign x_3264 = ~v_416 | v_30;
assign x_3265 = ~v_416 | ~v_31;
assign x_3266 = ~v_415 | v_117;
assign x_3267 = ~v_415 | v_25;
assign x_3268 = ~v_415 | ~v_31;
assign x_3269 = ~v_414 | v_122;
assign x_3270 = ~v_414 | v_26;
assign x_3271 = ~v_414 | ~v_31;
assign x_3272 = ~v_413 | v_126;
assign x_3273 = ~v_413 | v_27;
assign x_3274 = ~v_413 | ~v_31;
assign x_3275 = ~v_412 | v_129;
assign x_3276 = ~v_412 | v_28;
assign x_3277 = ~v_412 | ~v_31;
assign x_3278 = ~v_411 | v_131;
assign x_3279 = ~v_411 | v_29;
assign x_3280 = ~v_411 | ~v_31;
assign x_3281 = ~v_410 | v_132;
assign x_3282 = ~v_410 | v_30;
assign x_3283 = ~v_410 | ~v_31;
assign x_3284 = ~v_408 | ~v_112 | ~v_25 | v_26;
assign x_3285 = ~v_409 | ~v_33;
assign x_3286 = ~v_409 | v_34;
assign x_3287 = ~v_406 | ~v_113 | ~v_25 | v_27;
assign x_3288 = ~v_407 | ~v_33;
assign x_3289 = ~v_407 | v_35;
assign x_3290 = ~v_404 | ~v_114 | ~v_25 | v_28;
assign x_3291 = ~v_405 | ~v_33;
assign x_3292 = ~v_405 | v_36;
assign x_3293 = ~v_402 | ~v_115 | ~v_25 | v_29;
assign x_3294 = ~v_403 | ~v_33;
assign x_3295 = ~v_403 | v_37;
assign x_3296 = ~v_400 | ~v_116 | ~v_25 | v_30;
assign x_3297 = ~v_401 | ~v_33;
assign x_3298 = ~v_401 | v_38;
assign x_3299 = ~v_398 | ~v_117 | ~v_25 | v_31;
assign x_3300 = ~v_399 | ~v_33;
assign x_3301 = ~v_399 | v_39;
assign x_3302 = ~v_396 | ~v_118 | ~v_26 | v_27;
assign x_3303 = ~v_397 | ~v_34;
assign x_3304 = ~v_397 | v_35;
assign x_3305 = ~v_394 | ~v_119 | ~v_26 | v_28;
assign x_3306 = ~v_395 | ~v_34;
assign x_3307 = ~v_395 | v_36;
assign x_3308 = ~v_392 | ~v_120 | ~v_26 | v_29;
assign x_3309 = ~v_393 | ~v_34;
assign x_3310 = ~v_393 | v_37;
assign x_3311 = ~v_390 | ~v_121 | ~v_26 | v_30;
assign x_3312 = ~v_391 | ~v_34;
assign x_3313 = ~v_391 | v_38;
assign x_3314 = ~v_388 | ~v_122 | ~v_26 | v_31;
assign x_3315 = ~v_389 | ~v_34;
assign x_3316 = ~v_389 | v_39;
assign x_3317 = ~v_386 | ~v_123 | ~v_27 | v_28;
assign x_3318 = ~v_387 | ~v_35;
assign x_3319 = ~v_387 | v_36;
assign x_3320 = ~v_384 | ~v_124 | ~v_27 | v_29;
assign x_3321 = ~v_385 | ~v_35;
assign x_3322 = ~v_385 | v_37;
assign x_3323 = ~v_382 | ~v_125 | ~v_27 | v_30;
assign x_3324 = ~v_383 | ~v_35;
assign x_3325 = ~v_383 | v_38;
assign x_3326 = ~v_380 | ~v_126 | ~v_27 | v_31;
assign x_3327 = ~v_381 | ~v_35;
assign x_3328 = ~v_381 | v_39;
assign x_3329 = ~v_378 | ~v_127 | ~v_28 | v_29;
assign x_3330 = ~v_379 | ~v_36;
assign x_3331 = ~v_379 | v_37;
assign x_3332 = ~v_376 | ~v_128 | ~v_28 | v_30;
assign x_3333 = ~v_377 | ~v_36;
assign x_3334 = ~v_377 | v_38;
assign x_3335 = ~v_374 | ~v_129 | ~v_28 | v_31;
assign x_3336 = ~v_375 | ~v_36;
assign x_3337 = ~v_375 | v_39;
assign x_3338 = ~v_372 | ~v_130 | ~v_29 | v_30;
assign x_3339 = ~v_373 | ~v_37;
assign x_3340 = ~v_373 | v_38;
assign x_3341 = ~v_370 | ~v_131 | ~v_29 | v_31;
assign x_3342 = ~v_371 | ~v_37;
assign x_3343 = ~v_371 | v_39;
assign x_3344 = ~v_368 | ~v_132 | ~v_30 | v_31;
assign x_3345 = ~v_369 | ~v_38;
assign x_3346 = ~v_369 | v_39;
assign x_3347 = ~v_346 | v_33 | ~v_41;
assign x_3348 = ~v_346 | ~v_33 | v_41 | v_2214 | v_2213 | v_2212 | v_2211 | v_2210 | v_2209;
assign x_3349 = ~v_346 | ~v_2214 | v_345;
assign x_3350 = ~v_346 | ~v_133 | ~v_33 | v_34 | v_2214;
assign x_3351 = ~v_346 | ~v_2213 | v_344;
assign x_3352 = ~v_346 | ~v_134 | ~v_33 | v_35 | v_2213;
assign x_3353 = ~v_346 | ~v_2212 | v_343;
assign x_3354 = ~v_346 | ~v_135 | ~v_33 | v_36 | v_2212;
assign x_3355 = ~v_346 | ~v_2211 | v_342;
assign x_3356 = ~v_346 | ~v_136 | ~v_33 | v_37 | v_2211;
assign x_3357 = ~v_346 | ~v_2210 | v_341;
assign x_3358 = ~v_346 | ~v_137 | ~v_33 | v_38 | v_2210;
assign x_3359 = ~v_346 | ~v_2209 | v_340;
assign x_3360 = ~v_346 | ~v_138 | ~v_33 | v_39 | v_2209;
assign x_3361 = ~v_346 | v_34 | ~v_42 | v_2215;
assign x_3362 = ~v_346 | ~v_34 | v_42 | v_2220 | v_2219 | v_2218 | v_2217 | v_2216;
assign x_3363 = ~v_346 | ~v_2215 | v_339;
assign x_3364 = ~v_346 | ~v_133 | ~v_33 | v_34 | v_2215;
assign x_3365 = ~v_346 | ~v_2220 | v_338;
assign x_3366 = ~v_346 | ~v_139 | ~v_34 | v_35 | v_2220;
assign x_3367 = ~v_346 | ~v_2219 | v_337;
assign x_3368 = ~v_346 | ~v_140 | ~v_34 | v_36 | v_2219;
assign x_3369 = ~v_346 | ~v_2218 | v_336;
assign x_3370 = ~v_346 | ~v_141 | ~v_34 | v_37 | v_2218;
assign x_3371 = ~v_346 | ~v_2217 | v_335;
assign x_3372 = ~v_346 | ~v_142 | ~v_34 | v_38 | v_2217;
assign x_3373 = ~v_346 | ~v_2216 | v_334;
assign x_3374 = ~v_346 | ~v_143 | ~v_34 | v_39 | v_2216;
assign x_3375 = ~v_346 | v_35 | ~v_43 | v_2222 | v_2221;
assign x_3376 = ~v_346 | ~v_35 | v_43 | v_2226 | v_2225 | v_2224 | v_2223;
assign x_3377 = ~v_346 | ~v_2222 | v_333;
assign x_3378 = ~v_346 | ~v_134 | ~v_33 | v_35 | v_2222;
assign x_3379 = ~v_346 | ~v_2221 | v_332;
assign x_3380 = ~v_346 | ~v_139 | ~v_34 | v_35 | v_2221;
assign x_3381 = ~v_346 | ~v_2226 | v_331;
assign x_3382 = ~v_346 | ~v_144 | ~v_35 | v_36 | v_2226;
assign x_3383 = ~v_346 | ~v_2225 | v_330;
assign x_3384 = ~v_346 | ~v_145 | ~v_35 | v_37 | v_2225;
assign x_3385 = ~v_346 | ~v_2224 | v_329;
assign x_3386 = ~v_346 | ~v_146 | ~v_35 | v_38 | v_2224;
assign x_3387 = ~v_346 | ~v_2223 | v_328;
assign x_3388 = ~v_346 | ~v_147 | ~v_35 | v_39 | v_2223;
assign x_3389 = ~v_346 | v_36 | ~v_44 | v_2229 | v_2228 | v_2227;
assign x_3390 = ~v_346 | ~v_36 | v_44 | v_2232 | v_2231 | v_2230;
assign x_3391 = ~v_346 | ~v_2229 | v_327;
assign x_3392 = ~v_346 | ~v_135 | ~v_33 | v_36 | v_2229;
assign x_3393 = ~v_346 | ~v_2228 | v_326;
assign x_3394 = ~v_346 | ~v_140 | ~v_34 | v_36 | v_2228;
assign x_3395 = ~v_346 | ~v_2227 | v_325;
assign x_3396 = ~v_346 | ~v_144 | ~v_35 | v_36 | v_2227;
assign x_3397 = ~v_346 | ~v_2232 | v_324;
assign x_3398 = ~v_346 | ~v_148 | ~v_36 | v_37 | v_2232;
assign x_3399 = ~v_346 | ~v_2231 | v_323;
assign x_3400 = ~v_346 | ~v_149 | ~v_36 | v_38 | v_2231;
assign x_3401 = ~v_346 | ~v_2230 | v_322;
assign x_3402 = ~v_346 | ~v_150 | ~v_36 | v_39 | v_2230;
assign x_3403 = ~v_346 | v_37 | ~v_45 | v_2236 | v_2235 | v_2234 | v_2233;
assign x_3404 = ~v_346 | ~v_37 | v_45 | v_2238 | v_2237;
assign x_3405 = ~v_346 | ~v_2236 | v_321;
assign x_3406 = ~v_346 | ~v_136 | ~v_33 | v_37 | v_2236;
assign x_3407 = ~v_346 | ~v_2235 | v_320;
assign x_3408 = ~v_346 | ~v_141 | ~v_34 | v_37 | v_2235;
assign x_3409 = ~v_346 | ~v_2234 | v_319;
assign x_3410 = ~v_346 | ~v_145 | ~v_35 | v_37 | v_2234;
assign x_3411 = ~v_346 | ~v_2233 | v_318;
assign x_3412 = ~v_346 | ~v_148 | ~v_36 | v_37 | v_2233;
assign x_3413 = ~v_346 | ~v_2238 | v_317;
assign x_3414 = ~v_346 | ~v_151 | ~v_37 | v_38 | v_2238;
assign x_3415 = ~v_346 | ~v_2237 | v_316;
assign x_3416 = ~v_346 | ~v_152 | ~v_37 | v_39 | v_2237;
assign x_3417 = ~v_346 | v_38 | ~v_46 | v_2243 | v_2242 | v_2241 | v_2240 | v_2239;
assign x_3418 = ~v_346 | ~v_38 | v_46 | v_2244;
assign x_3419 = ~v_346 | ~v_2243 | v_315;
assign x_3420 = ~v_346 | ~v_137 | ~v_33 | v_38 | v_2243;
assign x_3421 = ~v_346 | ~v_2242 | v_314;
assign x_3422 = ~v_346 | ~v_142 | ~v_34 | v_38 | v_2242;
assign x_3423 = ~v_346 | ~v_2241 | v_313;
assign x_3424 = ~v_346 | ~v_146 | ~v_35 | v_38 | v_2241;
assign x_3425 = ~v_346 | ~v_2240 | v_312;
assign x_3426 = ~v_346 | ~v_149 | ~v_36 | v_38 | v_2240;
assign x_3427 = ~v_346 | ~v_2239 | v_311;
assign x_3428 = ~v_346 | ~v_151 | ~v_37 | v_38 | v_2239;
assign x_3429 = ~v_346 | ~v_2244 | v_310;
assign x_3430 = ~v_346 | ~v_153 | ~v_38 | v_39 | v_2244;
assign x_3431 = ~v_346 | v_39 | ~v_47 | v_2250 | v_2249 | v_2248 | v_2247 | v_2246 | v_2245;
assign x_3432 = ~v_346 | ~v_39 | v_47;
assign x_3433 = ~v_346 | ~v_2250 | v_309;
assign x_3434 = ~v_346 | ~v_138 | ~v_33 | v_39 | v_2250;
assign x_3435 = ~v_346 | ~v_2249 | v_308;
assign x_3436 = ~v_346 | ~v_143 | ~v_34 | v_39 | v_2249;
assign x_3437 = ~v_346 | ~v_2248 | v_307;
assign x_3438 = ~v_346 | ~v_147 | ~v_35 | v_39 | v_2248;
assign x_3439 = ~v_346 | ~v_2247 | v_306;
assign x_3440 = ~v_346 | ~v_150 | ~v_36 | v_39 | v_2247;
assign x_3441 = ~v_346 | ~v_2246 | v_305;
assign x_3442 = ~v_346 | ~v_152 | ~v_37 | v_39 | v_2246;
assign x_3443 = ~v_346 | ~v_2245 | v_304;
assign x_3444 = ~v_346 | ~v_153 | ~v_38 | v_39 | v_2245;
assign x_3445 = ~v_346 | v_40 | ~v_48;
assign x_3446 = ~v_346 | ~v_40 | v_48;
assign x_3447 = ~v_346 | v_302 | v_303;
assign x_3448 = ~v_346 | v_300 | v_301;
assign x_3449 = ~v_346 | v_298 | v_299;
assign x_3450 = ~v_346 | v_296 | v_297;
assign x_3451 = ~v_346 | v_294 | v_295;
assign x_3452 = ~v_346 | v_292 | v_293;
assign x_3453 = ~v_346 | v_290 | v_291;
assign x_3454 = ~v_346 | v_288 | v_289;
assign x_3455 = ~v_346 | v_286 | v_287;
assign x_3456 = ~v_346 | v_284 | v_285;
assign x_3457 = ~v_346 | v_282 | v_283;
assign x_3458 = ~v_346 | v_280 | v_281;
assign x_3459 = ~v_346 | v_278 | v_279;
assign x_3460 = ~v_346 | v_276 | v_277;
assign x_3461 = ~v_346 | v_274 | v_275;
assign x_3462 = ~v_346 | v_272 | v_273;
assign x_3463 = ~v_346 | v_270 | v_271;
assign x_3464 = ~v_346 | v_268 | v_269;
assign x_3465 = ~v_346 | v_266 | v_267;
assign x_3466 = ~v_346 | v_264 | v_265;
assign x_3467 = ~v_346 | v_262 | v_263;
assign x_3468 = ~v_346 | v_256 | v_257 | v_258 | v_259 | v_260 | v_261;
assign x_3469 = ~v_345 | v_133;
assign x_3470 = ~v_345 | v_33;
assign x_3471 = ~v_345 | ~v_34;
assign x_3472 = ~v_344 | v_134;
assign x_3473 = ~v_344 | v_33;
assign x_3474 = ~v_344 | ~v_35;
assign x_3475 = ~v_343 | v_135;
assign x_3476 = ~v_343 | v_33;
assign x_3477 = ~v_343 | ~v_36;
assign x_3478 = ~v_342 | v_136;
assign x_3479 = ~v_342 | v_33;
assign x_3480 = ~v_342 | ~v_37;
assign x_3481 = ~v_341 | v_137;
assign x_3482 = ~v_341 | v_33;
assign x_3483 = ~v_341 | ~v_38;
assign x_3484 = ~v_340 | v_138;
assign x_3485 = ~v_340 | v_33;
assign x_3486 = ~v_340 | ~v_39;
assign x_3487 = ~v_339 | v_133;
assign x_3488 = ~v_339 | v_33;
assign x_3489 = ~v_339 | ~v_34;
assign x_3490 = ~v_338 | v_139;
assign x_3491 = ~v_338 | v_34;
assign x_3492 = ~v_338 | ~v_35;
assign x_3493 = ~v_337 | v_140;
assign x_3494 = ~v_337 | v_34;
assign x_3495 = ~v_337 | ~v_36;
assign x_3496 = ~v_336 | v_141;
assign x_3497 = ~v_336 | v_34;
assign x_3498 = ~v_336 | ~v_37;
assign x_3499 = ~v_335 | v_142;
assign x_3500 = ~v_335 | v_34;
assign x_3501 = ~v_335 | ~v_38;
assign x_3502 = ~v_334 | v_143;
assign x_3503 = ~v_334 | v_34;
assign x_3504 = ~v_334 | ~v_39;
assign x_3505 = ~v_333 | v_134;
assign x_3506 = ~v_333 | v_33;
assign x_3507 = ~v_333 | ~v_35;
assign x_3508 = ~v_332 | v_139;
assign x_3509 = ~v_332 | v_34;
assign x_3510 = ~v_332 | ~v_35;
assign x_3511 = ~v_331 | v_144;
assign x_3512 = ~v_331 | v_35;
assign x_3513 = ~v_331 | ~v_36;
assign x_3514 = ~v_330 | v_145;
assign x_3515 = ~v_330 | v_35;
assign x_3516 = ~v_330 | ~v_37;
assign x_3517 = ~v_329 | v_146;
assign x_3518 = ~v_329 | v_35;
assign x_3519 = ~v_329 | ~v_38;
assign x_3520 = ~v_328 | v_147;
assign x_3521 = ~v_328 | v_35;
assign x_3522 = ~v_328 | ~v_39;
assign x_3523 = ~v_327 | v_135;
assign x_3524 = ~v_327 | v_33;
assign x_3525 = ~v_327 | ~v_36;
assign x_3526 = ~v_326 | v_140;
assign x_3527 = ~v_326 | v_34;
assign x_3528 = ~v_326 | ~v_36;
assign x_3529 = ~v_325 | v_144;
assign x_3530 = ~v_325 | v_35;
assign x_3531 = ~v_325 | ~v_36;
assign x_3532 = ~v_324 | v_148;
assign x_3533 = ~v_324 | v_36;
assign x_3534 = ~v_324 | ~v_37;
assign x_3535 = ~v_323 | v_149;
assign x_3536 = ~v_323 | v_36;
assign x_3537 = ~v_323 | ~v_38;
assign x_3538 = ~v_322 | v_150;
assign x_3539 = ~v_322 | v_36;
assign x_3540 = ~v_322 | ~v_39;
assign x_3541 = ~v_321 | v_136;
assign x_3542 = ~v_321 | v_33;
assign x_3543 = ~v_321 | ~v_37;
assign x_3544 = ~v_320 | v_141;
assign x_3545 = ~v_320 | v_34;
assign x_3546 = ~v_320 | ~v_37;
assign x_3547 = ~v_319 | v_145;
assign x_3548 = ~v_319 | v_35;
assign x_3549 = ~v_319 | ~v_37;
assign x_3550 = ~v_318 | v_148;
assign x_3551 = ~v_318 | v_36;
assign x_3552 = ~v_318 | ~v_37;
assign x_3553 = ~v_317 | v_151;
assign x_3554 = ~v_317 | v_37;
assign x_3555 = ~v_317 | ~v_38;
assign x_3556 = ~v_316 | v_152;
assign x_3557 = ~v_316 | v_37;
assign x_3558 = ~v_316 | ~v_39;
assign x_3559 = ~v_315 | v_137;
assign x_3560 = ~v_315 | v_33;
assign x_3561 = ~v_315 | ~v_38;
assign x_3562 = ~v_314 | v_142;
assign x_3563 = ~v_314 | v_34;
assign x_3564 = ~v_314 | ~v_38;
assign x_3565 = ~v_313 | v_146;
assign x_3566 = ~v_313 | v_35;
assign x_3567 = ~v_313 | ~v_38;
assign x_3568 = ~v_312 | v_149;
assign x_3569 = ~v_312 | v_36;
assign x_3570 = ~v_312 | ~v_38;
assign x_3571 = ~v_311 | v_151;
assign x_3572 = ~v_311 | v_37;
assign x_3573 = ~v_311 | ~v_38;
assign x_3574 = ~v_310 | v_153;
assign x_3575 = ~v_310 | v_38;
assign x_3576 = ~v_310 | ~v_39;
assign x_3577 = ~v_309 | v_138;
assign x_3578 = ~v_309 | v_33;
assign x_3579 = ~v_309 | ~v_39;
assign x_3580 = ~v_308 | v_143;
assign x_3581 = ~v_308 | v_34;
assign x_3582 = ~v_308 | ~v_39;
assign x_3583 = ~v_307 | v_147;
assign x_3584 = ~v_307 | v_35;
assign x_3585 = ~v_307 | ~v_39;
assign x_3586 = ~v_306 | v_150;
assign x_3587 = ~v_306 | v_36;
assign x_3588 = ~v_306 | ~v_39;
assign x_3589 = ~v_305 | v_152;
assign x_3590 = ~v_305 | v_37;
assign x_3591 = ~v_305 | ~v_39;
assign x_3592 = ~v_304 | v_153;
assign x_3593 = ~v_304 | v_38;
assign x_3594 = ~v_304 | ~v_39;
assign x_3595 = ~v_302 | ~v_133 | ~v_33 | v_34;
assign x_3596 = ~v_303 | ~v_41;
assign x_3597 = ~v_303 | v_42;
assign x_3598 = ~v_300 | ~v_134 | ~v_33 | v_35;
assign x_3599 = ~v_301 | ~v_41;
assign x_3600 = ~v_301 | v_43;
assign x_3601 = ~v_298 | ~v_135 | ~v_33 | v_36;
assign x_3602 = ~v_299 | ~v_41;
assign x_3603 = ~v_299 | v_44;
assign x_3604 = ~v_296 | ~v_136 | ~v_33 | v_37;
assign x_3605 = ~v_297 | ~v_41;
assign x_3606 = ~v_297 | v_45;
assign x_3607 = ~v_294 | ~v_137 | ~v_33 | v_38;
assign x_3608 = ~v_295 | ~v_41;
assign x_3609 = ~v_295 | v_46;
assign x_3610 = ~v_292 | ~v_138 | ~v_33 | v_39;
assign x_3611 = ~v_293 | ~v_41;
assign x_3612 = ~v_293 | v_47;
assign x_3613 = ~v_290 | ~v_139 | ~v_34 | v_35;
assign x_3614 = ~v_291 | ~v_42;
assign x_3615 = ~v_291 | v_43;
assign x_3616 = ~v_288 | ~v_140 | ~v_34 | v_36;
assign x_3617 = ~v_289 | ~v_42;
assign x_3618 = ~v_289 | v_44;
assign x_3619 = ~v_286 | ~v_141 | ~v_34 | v_37;
assign x_3620 = ~v_287 | ~v_42;
assign x_3621 = ~v_287 | v_45;
assign x_3622 = ~v_284 | ~v_142 | ~v_34 | v_38;
assign x_3623 = ~v_285 | ~v_42;
assign x_3624 = ~v_285 | v_46;
assign x_3625 = ~v_282 | ~v_143 | ~v_34 | v_39;
assign x_3626 = ~v_283 | ~v_42;
assign x_3627 = ~v_283 | v_47;
assign x_3628 = ~v_280 | ~v_144 | ~v_35 | v_36;
assign x_3629 = ~v_281 | ~v_43;
assign x_3630 = ~v_281 | v_44;
assign x_3631 = ~v_278 | ~v_145 | ~v_35 | v_37;
assign x_3632 = ~v_279 | ~v_43;
assign x_3633 = ~v_279 | v_45;
assign x_3634 = ~v_276 | ~v_146 | ~v_35 | v_38;
assign x_3635 = ~v_277 | ~v_43;
assign x_3636 = ~v_277 | v_46;
assign x_3637 = ~v_274 | ~v_147 | ~v_35 | v_39;
assign x_3638 = ~v_275 | ~v_43;
assign x_3639 = ~v_275 | v_47;
assign x_3640 = ~v_272 | ~v_148 | ~v_36 | v_37;
assign x_3641 = ~v_273 | ~v_44;
assign x_3642 = ~v_273 | v_45;
assign x_3643 = ~v_270 | ~v_149 | ~v_36 | v_38;
assign x_3644 = ~v_271 | ~v_44;
assign x_3645 = ~v_271 | v_46;
assign x_3646 = ~v_268 | ~v_150 | ~v_36 | v_39;
assign x_3647 = ~v_269 | ~v_44;
assign x_3648 = ~v_269 | v_47;
assign x_3649 = ~v_266 | ~v_151 | ~v_37 | v_38;
assign x_3650 = ~v_267 | ~v_45;
assign x_3651 = ~v_267 | v_46;
assign x_3652 = ~v_264 | ~v_152 | ~v_37 | v_39;
assign x_3653 = ~v_265 | ~v_45;
assign x_3654 = ~v_265 | v_47;
assign x_3655 = ~v_262 | ~v_153 | ~v_38 | v_39;
assign x_3656 = ~v_263 | ~v_46;
assign x_3657 = ~v_263 | v_47;
assign x_3658 = ~v_256 | v_41;
assign x_3659 = ~v_256 | ~v_42;
assign x_3660 = ~v_257 | v_42;
assign x_3661 = ~v_257 | ~v_43;
assign x_3662 = ~v_258 | v_43;
assign x_3663 = ~v_258 | ~v_44;
assign x_3664 = ~v_259 | v_44;
assign x_3665 = ~v_259 | ~v_45;
assign x_3666 = ~v_260 | v_45;
assign x_3667 = ~v_260 | ~v_46;
assign x_3668 = ~v_261 | v_46;
assign x_3669 = ~v_261 | ~v_47;
assign x_3670 = x_2 & x_3;
assign x_3671 = x_1 & x_3670;
assign x_3672 = x_4 & x_5;
assign x_3673 = x_6 & x_7;
assign x_3674 = x_3672 & x_3673;
assign x_3675 = x_3671 & x_3674;
assign x_3676 = x_9 & x_10;
assign x_3677 = x_8 & x_3676;
assign x_3678 = x_11 & x_12;
assign x_3679 = x_13 & x_14;
assign x_3680 = x_3678 & x_3679;
assign x_3681 = x_3677 & x_3680;
assign x_3682 = x_3675 & x_3681;
assign x_3683 = x_16 & x_17;
assign x_3684 = x_15 & x_3683;
assign x_3685 = x_18 & x_19;
assign x_3686 = x_20 & x_21;
assign x_3687 = x_3685 & x_3686;
assign x_3688 = x_3684 & x_3687;
assign x_3689 = x_23 & x_24;
assign x_3690 = x_22 & x_3689;
assign x_3691 = x_25 & x_26;
assign x_3692 = x_27 & x_28;
assign x_3693 = x_3691 & x_3692;
assign x_3694 = x_3690 & x_3693;
assign x_3695 = x_3688 & x_3694;
assign x_3696 = x_3682 & x_3695;
assign x_3697 = x_30 & x_31;
assign x_3698 = x_29 & x_3697;
assign x_3699 = x_32 & x_33;
assign x_3700 = x_34 & x_35;
assign x_3701 = x_3699 & x_3700;
assign x_3702 = x_3698 & x_3701;
assign x_3703 = x_37 & x_38;
assign x_3704 = x_36 & x_3703;
assign x_3705 = x_39 & x_40;
assign x_3706 = x_41 & x_42;
assign x_3707 = x_3705 & x_3706;
assign x_3708 = x_3704 & x_3707;
assign x_3709 = x_3702 & x_3708;
assign x_3710 = x_44 & x_45;
assign x_3711 = x_43 & x_3710;
assign x_3712 = x_46 & x_47;
assign x_3713 = x_48 & x_49;
assign x_3714 = x_3712 & x_3713;
assign x_3715 = x_3711 & x_3714;
assign x_3716 = x_50 & x_51;
assign x_3717 = x_52 & x_53;
assign x_3718 = x_3716 & x_3717;
assign x_3719 = x_54 & x_55;
assign x_3720 = x_56 & x_57;
assign x_3721 = x_3719 & x_3720;
assign x_3722 = x_3718 & x_3721;
assign x_3723 = x_3715 & x_3722;
assign x_3724 = x_3709 & x_3723;
assign x_3725 = x_3696 & x_3724;
assign x_3726 = x_59 & x_60;
assign x_3727 = x_58 & x_3726;
assign x_3728 = x_61 & x_62;
assign x_3729 = x_63 & x_64;
assign x_3730 = x_3728 & x_3729;
assign x_3731 = x_3727 & x_3730;
assign x_3732 = x_66 & x_67;
assign x_3733 = x_65 & x_3732;
assign x_3734 = x_68 & x_69;
assign x_3735 = x_70 & x_71;
assign x_3736 = x_3734 & x_3735;
assign x_3737 = x_3733 & x_3736;
assign x_3738 = x_3731 & x_3737;
assign x_3739 = x_73 & x_74;
assign x_3740 = x_72 & x_3739;
assign x_3741 = x_75 & x_76;
assign x_3742 = x_77 & x_78;
assign x_3743 = x_3741 & x_3742;
assign x_3744 = x_3740 & x_3743;
assign x_3745 = x_80 & x_81;
assign x_3746 = x_79 & x_3745;
assign x_3747 = x_82 & x_83;
assign x_3748 = x_84 & x_85;
assign x_3749 = x_3747 & x_3748;
assign x_3750 = x_3746 & x_3749;
assign x_3751 = x_3744 & x_3750;
assign x_3752 = x_3738 & x_3751;
assign x_3753 = x_87 & x_88;
assign x_3754 = x_86 & x_3753;
assign x_3755 = x_89 & x_90;
assign x_3756 = x_91 & x_92;
assign x_3757 = x_3755 & x_3756;
assign x_3758 = x_3754 & x_3757;
assign x_3759 = x_94 & x_95;
assign x_3760 = x_93 & x_3759;
assign x_3761 = x_96 & x_97;
assign x_3762 = x_98 & x_99;
assign x_3763 = x_3761 & x_3762;
assign x_3764 = x_3760 & x_3763;
assign x_3765 = x_3758 & x_3764;
assign x_3766 = x_101 & x_102;
assign x_3767 = x_100 & x_3766;
assign x_3768 = x_103 & x_104;
assign x_3769 = x_105 & x_106;
assign x_3770 = x_3768 & x_3769;
assign x_3771 = x_3767 & x_3770;
assign x_3772 = x_107 & x_108;
assign x_3773 = x_109 & x_110;
assign x_3774 = x_3772 & x_3773;
assign x_3775 = x_111 & x_112;
assign x_3776 = x_113 & x_114;
assign x_3777 = x_3775 & x_3776;
assign x_3778 = x_3774 & x_3777;
assign x_3779 = x_3771 & x_3778;
assign x_3780 = x_3765 & x_3779;
assign x_3781 = x_3752 & x_3780;
assign x_3782 = x_3725 & x_3781;
assign x_3783 = x_116 & x_117;
assign x_3784 = x_115 & x_3783;
assign x_3785 = x_118 & x_119;
assign x_3786 = x_120 & x_121;
assign x_3787 = x_3785 & x_3786;
assign x_3788 = x_3784 & x_3787;
assign x_3789 = x_123 & x_124;
assign x_3790 = x_122 & x_3789;
assign x_3791 = x_125 & x_126;
assign x_3792 = x_127 & x_128;
assign x_3793 = x_3791 & x_3792;
assign x_3794 = x_3790 & x_3793;
assign x_3795 = x_3788 & x_3794;
assign x_3796 = x_130 & x_131;
assign x_3797 = x_129 & x_3796;
assign x_3798 = x_132 & x_133;
assign x_3799 = x_134 & x_135;
assign x_3800 = x_3798 & x_3799;
assign x_3801 = x_3797 & x_3800;
assign x_3802 = x_137 & x_138;
assign x_3803 = x_136 & x_3802;
assign x_3804 = x_139 & x_140;
assign x_3805 = x_141 & x_142;
assign x_3806 = x_3804 & x_3805;
assign x_3807 = x_3803 & x_3806;
assign x_3808 = x_3801 & x_3807;
assign x_3809 = x_3795 & x_3808;
assign x_3810 = x_144 & x_145;
assign x_3811 = x_143 & x_3810;
assign x_3812 = x_146 & x_147;
assign x_3813 = x_148 & x_149;
assign x_3814 = x_3812 & x_3813;
assign x_3815 = x_3811 & x_3814;
assign x_3816 = x_151 & x_152;
assign x_3817 = x_150 & x_3816;
assign x_3818 = x_153 & x_154;
assign x_3819 = x_155 & x_156;
assign x_3820 = x_3818 & x_3819;
assign x_3821 = x_3817 & x_3820;
assign x_3822 = x_3815 & x_3821;
assign x_3823 = x_158 & x_159;
assign x_3824 = x_157 & x_3823;
assign x_3825 = x_160 & x_161;
assign x_3826 = x_162 & x_163;
assign x_3827 = x_3825 & x_3826;
assign x_3828 = x_3824 & x_3827;
assign x_3829 = x_164 & x_165;
assign x_3830 = x_166 & x_167;
assign x_3831 = x_3829 & x_3830;
assign x_3832 = x_168 & x_169;
assign x_3833 = x_170 & x_171;
assign x_3834 = x_3832 & x_3833;
assign x_3835 = x_3831 & x_3834;
assign x_3836 = x_3828 & x_3835;
assign x_3837 = x_3822 & x_3836;
assign x_3838 = x_3809 & x_3837;
assign x_3839 = x_173 & x_174;
assign x_3840 = x_172 & x_3839;
assign x_3841 = x_175 & x_176;
assign x_3842 = x_177 & x_178;
assign x_3843 = x_3841 & x_3842;
assign x_3844 = x_3840 & x_3843;
assign x_3845 = x_180 & x_181;
assign x_3846 = x_179 & x_3845;
assign x_3847 = x_182 & x_183;
assign x_3848 = x_184 & x_185;
assign x_3849 = x_3847 & x_3848;
assign x_3850 = x_3846 & x_3849;
assign x_3851 = x_3844 & x_3850;
assign x_3852 = x_187 & x_188;
assign x_3853 = x_186 & x_3852;
assign x_3854 = x_189 & x_190;
assign x_3855 = x_191 & x_192;
assign x_3856 = x_3854 & x_3855;
assign x_3857 = x_3853 & x_3856;
assign x_3858 = x_193 & x_194;
assign x_3859 = x_195 & x_196;
assign x_3860 = x_3858 & x_3859;
assign x_3861 = x_197 & x_198;
assign x_3862 = x_199 & x_200;
assign x_3863 = x_3861 & x_3862;
assign x_3864 = x_3860 & x_3863;
assign x_3865 = x_3857 & x_3864;
assign x_3866 = x_3851 & x_3865;
assign x_3867 = x_202 & x_203;
assign x_3868 = x_201 & x_3867;
assign x_3869 = x_204 & x_205;
assign x_3870 = x_206 & x_207;
assign x_3871 = x_3869 & x_3870;
assign x_3872 = x_3868 & x_3871;
assign x_3873 = x_209 & x_210;
assign x_3874 = x_208 & x_3873;
assign x_3875 = x_211 & x_212;
assign x_3876 = x_213 & x_214;
assign x_3877 = x_3875 & x_3876;
assign x_3878 = x_3874 & x_3877;
assign x_3879 = x_3872 & x_3878;
assign x_3880 = x_216 & x_217;
assign x_3881 = x_215 & x_3880;
assign x_3882 = x_218 & x_219;
assign x_3883 = x_220 & x_221;
assign x_3884 = x_3882 & x_3883;
assign x_3885 = x_3881 & x_3884;
assign x_3886 = x_222 & x_223;
assign x_3887 = x_224 & x_225;
assign x_3888 = x_3886 & x_3887;
assign x_3889 = x_226 & x_227;
assign x_3890 = x_228 & x_229;
assign x_3891 = x_3889 & x_3890;
assign x_3892 = x_3888 & x_3891;
assign x_3893 = x_3885 & x_3892;
assign x_3894 = x_3879 & x_3893;
assign x_3895 = x_3866 & x_3894;
assign x_3896 = x_3838 & x_3895;
assign x_3897 = x_3782 & x_3896;
assign x_3898 = x_231 & x_232;
assign x_3899 = x_230 & x_3898;
assign x_3900 = x_233 & x_234;
assign x_3901 = x_235 & x_236;
assign x_3902 = x_3900 & x_3901;
assign x_3903 = x_3899 & x_3902;
assign x_3904 = x_238 & x_239;
assign x_3905 = x_237 & x_3904;
assign x_3906 = x_240 & x_241;
assign x_3907 = x_242 & x_243;
assign x_3908 = x_3906 & x_3907;
assign x_3909 = x_3905 & x_3908;
assign x_3910 = x_3903 & x_3909;
assign x_3911 = x_245 & x_246;
assign x_3912 = x_244 & x_3911;
assign x_3913 = x_247 & x_248;
assign x_3914 = x_249 & x_250;
assign x_3915 = x_3913 & x_3914;
assign x_3916 = x_3912 & x_3915;
assign x_3917 = x_252 & x_253;
assign x_3918 = x_251 & x_3917;
assign x_3919 = x_254 & x_255;
assign x_3920 = x_256 & x_257;
assign x_3921 = x_3919 & x_3920;
assign x_3922 = x_3918 & x_3921;
assign x_3923 = x_3916 & x_3922;
assign x_3924 = x_3910 & x_3923;
assign x_3925 = x_259 & x_260;
assign x_3926 = x_258 & x_3925;
assign x_3927 = x_261 & x_262;
assign x_3928 = x_263 & x_264;
assign x_3929 = x_3927 & x_3928;
assign x_3930 = x_3926 & x_3929;
assign x_3931 = x_266 & x_267;
assign x_3932 = x_265 & x_3931;
assign x_3933 = x_268 & x_269;
assign x_3934 = x_270 & x_271;
assign x_3935 = x_3933 & x_3934;
assign x_3936 = x_3932 & x_3935;
assign x_3937 = x_3930 & x_3936;
assign x_3938 = x_273 & x_274;
assign x_3939 = x_272 & x_3938;
assign x_3940 = x_275 & x_276;
assign x_3941 = x_277 & x_278;
assign x_3942 = x_3940 & x_3941;
assign x_3943 = x_3939 & x_3942;
assign x_3944 = x_279 & x_280;
assign x_3945 = x_281 & x_282;
assign x_3946 = x_3944 & x_3945;
assign x_3947 = x_283 & x_284;
assign x_3948 = x_285 & x_286;
assign x_3949 = x_3947 & x_3948;
assign x_3950 = x_3946 & x_3949;
assign x_3951 = x_3943 & x_3950;
assign x_3952 = x_3937 & x_3951;
assign x_3953 = x_3924 & x_3952;
assign x_3954 = x_288 & x_289;
assign x_3955 = x_287 & x_3954;
assign x_3956 = x_290 & x_291;
assign x_3957 = x_292 & x_293;
assign x_3958 = x_3956 & x_3957;
assign x_3959 = x_3955 & x_3958;
assign x_3960 = x_295 & x_296;
assign x_3961 = x_294 & x_3960;
assign x_3962 = x_297 & x_298;
assign x_3963 = x_299 & x_300;
assign x_3964 = x_3962 & x_3963;
assign x_3965 = x_3961 & x_3964;
assign x_3966 = x_3959 & x_3965;
assign x_3967 = x_302 & x_303;
assign x_3968 = x_301 & x_3967;
assign x_3969 = x_304 & x_305;
assign x_3970 = x_306 & x_307;
assign x_3971 = x_3969 & x_3970;
assign x_3972 = x_3968 & x_3971;
assign x_3973 = x_309 & x_310;
assign x_3974 = x_308 & x_3973;
assign x_3975 = x_311 & x_312;
assign x_3976 = x_313 & x_314;
assign x_3977 = x_3975 & x_3976;
assign x_3978 = x_3974 & x_3977;
assign x_3979 = x_3972 & x_3978;
assign x_3980 = x_3966 & x_3979;
assign x_3981 = x_316 & x_317;
assign x_3982 = x_315 & x_3981;
assign x_3983 = x_318 & x_319;
assign x_3984 = x_320 & x_321;
assign x_3985 = x_3983 & x_3984;
assign x_3986 = x_3982 & x_3985;
assign x_3987 = x_323 & x_324;
assign x_3988 = x_322 & x_3987;
assign x_3989 = x_325 & x_326;
assign x_3990 = x_327 & x_328;
assign x_3991 = x_3989 & x_3990;
assign x_3992 = x_3988 & x_3991;
assign x_3993 = x_3986 & x_3992;
assign x_3994 = x_330 & x_331;
assign x_3995 = x_329 & x_3994;
assign x_3996 = x_332 & x_333;
assign x_3997 = x_334 & x_335;
assign x_3998 = x_3996 & x_3997;
assign x_3999 = x_3995 & x_3998;
assign x_4000 = x_336 & x_337;
assign x_4001 = x_338 & x_339;
assign x_4002 = x_4000 & x_4001;
assign x_4003 = x_340 & x_341;
assign x_4004 = x_342 & x_343;
assign x_4005 = x_4003 & x_4004;
assign x_4006 = x_4002 & x_4005;
assign x_4007 = x_3999 & x_4006;
assign x_4008 = x_3993 & x_4007;
assign x_4009 = x_3980 & x_4008;
assign x_4010 = x_3953 & x_4009;
assign x_4011 = x_345 & x_346;
assign x_4012 = x_344 & x_4011;
assign x_4013 = x_347 & x_348;
assign x_4014 = x_349 & x_350;
assign x_4015 = x_4013 & x_4014;
assign x_4016 = x_4012 & x_4015;
assign x_4017 = x_352 & x_353;
assign x_4018 = x_351 & x_4017;
assign x_4019 = x_354 & x_355;
assign x_4020 = x_356 & x_357;
assign x_4021 = x_4019 & x_4020;
assign x_4022 = x_4018 & x_4021;
assign x_4023 = x_4016 & x_4022;
assign x_4024 = x_359 & x_360;
assign x_4025 = x_358 & x_4024;
assign x_4026 = x_361 & x_362;
assign x_4027 = x_363 & x_364;
assign x_4028 = x_4026 & x_4027;
assign x_4029 = x_4025 & x_4028;
assign x_4030 = x_366 & x_367;
assign x_4031 = x_365 & x_4030;
assign x_4032 = x_368 & x_369;
assign x_4033 = x_370 & x_371;
assign x_4034 = x_4032 & x_4033;
assign x_4035 = x_4031 & x_4034;
assign x_4036 = x_4029 & x_4035;
assign x_4037 = x_4023 & x_4036;
assign x_4038 = x_373 & x_374;
assign x_4039 = x_372 & x_4038;
assign x_4040 = x_375 & x_376;
assign x_4041 = x_377 & x_378;
assign x_4042 = x_4040 & x_4041;
assign x_4043 = x_4039 & x_4042;
assign x_4044 = x_380 & x_381;
assign x_4045 = x_379 & x_4044;
assign x_4046 = x_382 & x_383;
assign x_4047 = x_384 & x_385;
assign x_4048 = x_4046 & x_4047;
assign x_4049 = x_4045 & x_4048;
assign x_4050 = x_4043 & x_4049;
assign x_4051 = x_387 & x_388;
assign x_4052 = x_386 & x_4051;
assign x_4053 = x_389 & x_390;
assign x_4054 = x_391 & x_392;
assign x_4055 = x_4053 & x_4054;
assign x_4056 = x_4052 & x_4055;
assign x_4057 = x_393 & x_394;
assign x_4058 = x_395 & x_396;
assign x_4059 = x_4057 & x_4058;
assign x_4060 = x_397 & x_398;
assign x_4061 = x_399 & x_400;
assign x_4062 = x_4060 & x_4061;
assign x_4063 = x_4059 & x_4062;
assign x_4064 = x_4056 & x_4063;
assign x_4065 = x_4050 & x_4064;
assign x_4066 = x_4037 & x_4065;
assign x_4067 = x_402 & x_403;
assign x_4068 = x_401 & x_4067;
assign x_4069 = x_404 & x_405;
assign x_4070 = x_406 & x_407;
assign x_4071 = x_4069 & x_4070;
assign x_4072 = x_4068 & x_4071;
assign x_4073 = x_409 & x_410;
assign x_4074 = x_408 & x_4073;
assign x_4075 = x_411 & x_412;
assign x_4076 = x_413 & x_414;
assign x_4077 = x_4075 & x_4076;
assign x_4078 = x_4074 & x_4077;
assign x_4079 = x_4072 & x_4078;
assign x_4080 = x_416 & x_417;
assign x_4081 = x_415 & x_4080;
assign x_4082 = x_418 & x_419;
assign x_4083 = x_420 & x_421;
assign x_4084 = x_4082 & x_4083;
assign x_4085 = x_4081 & x_4084;
assign x_4086 = x_422 & x_423;
assign x_4087 = x_424 & x_425;
assign x_4088 = x_4086 & x_4087;
assign x_4089 = x_426 & x_427;
assign x_4090 = x_428 & x_429;
assign x_4091 = x_4089 & x_4090;
assign x_4092 = x_4088 & x_4091;
assign x_4093 = x_4085 & x_4092;
assign x_4094 = x_4079 & x_4093;
assign x_4095 = x_431 & x_432;
assign x_4096 = x_430 & x_4095;
assign x_4097 = x_433 & x_434;
assign x_4098 = x_435 & x_436;
assign x_4099 = x_4097 & x_4098;
assign x_4100 = x_4096 & x_4099;
assign x_4101 = x_438 & x_439;
assign x_4102 = x_437 & x_4101;
assign x_4103 = x_440 & x_441;
assign x_4104 = x_442 & x_443;
assign x_4105 = x_4103 & x_4104;
assign x_4106 = x_4102 & x_4105;
assign x_4107 = x_4100 & x_4106;
assign x_4108 = x_445 & x_446;
assign x_4109 = x_444 & x_4108;
assign x_4110 = x_447 & x_448;
assign x_4111 = x_449 & x_450;
assign x_4112 = x_4110 & x_4111;
assign x_4113 = x_4109 & x_4112;
assign x_4114 = x_451 & x_452;
assign x_4115 = x_453 & x_454;
assign x_4116 = x_4114 & x_4115;
assign x_4117 = x_455 & x_456;
assign x_4118 = x_457 & x_458;
assign x_4119 = x_4117 & x_4118;
assign x_4120 = x_4116 & x_4119;
assign x_4121 = x_4113 & x_4120;
assign x_4122 = x_4107 & x_4121;
assign x_4123 = x_4094 & x_4122;
assign x_4124 = x_4066 & x_4123;
assign x_4125 = x_4010 & x_4124;
assign x_4126 = x_3897 & x_4125;
assign x_4127 = x_460 & x_461;
assign x_4128 = x_459 & x_4127;
assign x_4129 = x_462 & x_463;
assign x_4130 = x_464 & x_465;
assign x_4131 = x_4129 & x_4130;
assign x_4132 = x_4128 & x_4131;
assign x_4133 = x_467 & x_468;
assign x_4134 = x_466 & x_4133;
assign x_4135 = x_469 & x_470;
assign x_4136 = x_471 & x_472;
assign x_4137 = x_4135 & x_4136;
assign x_4138 = x_4134 & x_4137;
assign x_4139 = x_4132 & x_4138;
assign x_4140 = x_474 & x_475;
assign x_4141 = x_473 & x_4140;
assign x_4142 = x_476 & x_477;
assign x_4143 = x_478 & x_479;
assign x_4144 = x_4142 & x_4143;
assign x_4145 = x_4141 & x_4144;
assign x_4146 = x_481 & x_482;
assign x_4147 = x_480 & x_4146;
assign x_4148 = x_483 & x_484;
assign x_4149 = x_485 & x_486;
assign x_4150 = x_4148 & x_4149;
assign x_4151 = x_4147 & x_4150;
assign x_4152 = x_4145 & x_4151;
assign x_4153 = x_4139 & x_4152;
assign x_4154 = x_488 & x_489;
assign x_4155 = x_487 & x_4154;
assign x_4156 = x_490 & x_491;
assign x_4157 = x_492 & x_493;
assign x_4158 = x_4156 & x_4157;
assign x_4159 = x_4155 & x_4158;
assign x_4160 = x_495 & x_496;
assign x_4161 = x_494 & x_4160;
assign x_4162 = x_497 & x_498;
assign x_4163 = x_499 & x_500;
assign x_4164 = x_4162 & x_4163;
assign x_4165 = x_4161 & x_4164;
assign x_4166 = x_4159 & x_4165;
assign x_4167 = x_502 & x_503;
assign x_4168 = x_501 & x_4167;
assign x_4169 = x_504 & x_505;
assign x_4170 = x_506 & x_507;
assign x_4171 = x_4169 & x_4170;
assign x_4172 = x_4168 & x_4171;
assign x_4173 = x_508 & x_509;
assign x_4174 = x_510 & x_511;
assign x_4175 = x_4173 & x_4174;
assign x_4176 = x_512 & x_513;
assign x_4177 = x_514 & x_515;
assign x_4178 = x_4176 & x_4177;
assign x_4179 = x_4175 & x_4178;
assign x_4180 = x_4172 & x_4179;
assign x_4181 = x_4166 & x_4180;
assign x_4182 = x_4153 & x_4181;
assign x_4183 = x_517 & x_518;
assign x_4184 = x_516 & x_4183;
assign x_4185 = x_519 & x_520;
assign x_4186 = x_521 & x_522;
assign x_4187 = x_4185 & x_4186;
assign x_4188 = x_4184 & x_4187;
assign x_4189 = x_524 & x_525;
assign x_4190 = x_523 & x_4189;
assign x_4191 = x_526 & x_527;
assign x_4192 = x_528 & x_529;
assign x_4193 = x_4191 & x_4192;
assign x_4194 = x_4190 & x_4193;
assign x_4195 = x_4188 & x_4194;
assign x_4196 = x_531 & x_532;
assign x_4197 = x_530 & x_4196;
assign x_4198 = x_533 & x_534;
assign x_4199 = x_535 & x_536;
assign x_4200 = x_4198 & x_4199;
assign x_4201 = x_4197 & x_4200;
assign x_4202 = x_538 & x_539;
assign x_4203 = x_537 & x_4202;
assign x_4204 = x_540 & x_541;
assign x_4205 = x_542 & x_543;
assign x_4206 = x_4204 & x_4205;
assign x_4207 = x_4203 & x_4206;
assign x_4208 = x_4201 & x_4207;
assign x_4209 = x_4195 & x_4208;
assign x_4210 = x_545 & x_546;
assign x_4211 = x_544 & x_4210;
assign x_4212 = x_547 & x_548;
assign x_4213 = x_549 & x_550;
assign x_4214 = x_4212 & x_4213;
assign x_4215 = x_4211 & x_4214;
assign x_4216 = x_552 & x_553;
assign x_4217 = x_551 & x_4216;
assign x_4218 = x_554 & x_555;
assign x_4219 = x_556 & x_557;
assign x_4220 = x_4218 & x_4219;
assign x_4221 = x_4217 & x_4220;
assign x_4222 = x_4215 & x_4221;
assign x_4223 = x_559 & x_560;
assign x_4224 = x_558 & x_4223;
assign x_4225 = x_561 & x_562;
assign x_4226 = x_563 & x_564;
assign x_4227 = x_4225 & x_4226;
assign x_4228 = x_4224 & x_4227;
assign x_4229 = x_565 & x_566;
assign x_4230 = x_567 & x_568;
assign x_4231 = x_4229 & x_4230;
assign x_4232 = x_569 & x_570;
assign x_4233 = x_571 & x_572;
assign x_4234 = x_4232 & x_4233;
assign x_4235 = x_4231 & x_4234;
assign x_4236 = x_4228 & x_4235;
assign x_4237 = x_4222 & x_4236;
assign x_4238 = x_4209 & x_4237;
assign x_4239 = x_4182 & x_4238;
assign x_4240 = x_574 & x_575;
assign x_4241 = x_573 & x_4240;
assign x_4242 = x_576 & x_577;
assign x_4243 = x_578 & x_579;
assign x_4244 = x_4242 & x_4243;
assign x_4245 = x_4241 & x_4244;
assign x_4246 = x_581 & x_582;
assign x_4247 = x_580 & x_4246;
assign x_4248 = x_583 & x_584;
assign x_4249 = x_585 & x_586;
assign x_4250 = x_4248 & x_4249;
assign x_4251 = x_4247 & x_4250;
assign x_4252 = x_4245 & x_4251;
assign x_4253 = x_588 & x_589;
assign x_4254 = x_587 & x_4253;
assign x_4255 = x_590 & x_591;
assign x_4256 = x_592 & x_593;
assign x_4257 = x_4255 & x_4256;
assign x_4258 = x_4254 & x_4257;
assign x_4259 = x_595 & x_596;
assign x_4260 = x_594 & x_4259;
assign x_4261 = x_597 & x_598;
assign x_4262 = x_599 & x_600;
assign x_4263 = x_4261 & x_4262;
assign x_4264 = x_4260 & x_4263;
assign x_4265 = x_4258 & x_4264;
assign x_4266 = x_4252 & x_4265;
assign x_4267 = x_602 & x_603;
assign x_4268 = x_601 & x_4267;
assign x_4269 = x_604 & x_605;
assign x_4270 = x_606 & x_607;
assign x_4271 = x_4269 & x_4270;
assign x_4272 = x_4268 & x_4271;
assign x_4273 = x_609 & x_610;
assign x_4274 = x_608 & x_4273;
assign x_4275 = x_611 & x_612;
assign x_4276 = x_613 & x_614;
assign x_4277 = x_4275 & x_4276;
assign x_4278 = x_4274 & x_4277;
assign x_4279 = x_4272 & x_4278;
assign x_4280 = x_616 & x_617;
assign x_4281 = x_615 & x_4280;
assign x_4282 = x_618 & x_619;
assign x_4283 = x_620 & x_621;
assign x_4284 = x_4282 & x_4283;
assign x_4285 = x_4281 & x_4284;
assign x_4286 = x_622 & x_623;
assign x_4287 = x_624 & x_625;
assign x_4288 = x_4286 & x_4287;
assign x_4289 = x_626 & x_627;
assign x_4290 = x_628 & x_629;
assign x_4291 = x_4289 & x_4290;
assign x_4292 = x_4288 & x_4291;
assign x_4293 = x_4285 & x_4292;
assign x_4294 = x_4279 & x_4293;
assign x_4295 = x_4266 & x_4294;
assign x_4296 = x_631 & x_632;
assign x_4297 = x_630 & x_4296;
assign x_4298 = x_633 & x_634;
assign x_4299 = x_635 & x_636;
assign x_4300 = x_4298 & x_4299;
assign x_4301 = x_4297 & x_4300;
assign x_4302 = x_638 & x_639;
assign x_4303 = x_637 & x_4302;
assign x_4304 = x_640 & x_641;
assign x_4305 = x_642 & x_643;
assign x_4306 = x_4304 & x_4305;
assign x_4307 = x_4303 & x_4306;
assign x_4308 = x_4301 & x_4307;
assign x_4309 = x_645 & x_646;
assign x_4310 = x_644 & x_4309;
assign x_4311 = x_647 & x_648;
assign x_4312 = x_649 & x_650;
assign x_4313 = x_4311 & x_4312;
assign x_4314 = x_4310 & x_4313;
assign x_4315 = x_651 & x_652;
assign x_4316 = x_653 & x_654;
assign x_4317 = x_4315 & x_4316;
assign x_4318 = x_655 & x_656;
assign x_4319 = x_657 & x_658;
assign x_4320 = x_4318 & x_4319;
assign x_4321 = x_4317 & x_4320;
assign x_4322 = x_4314 & x_4321;
assign x_4323 = x_4308 & x_4322;
assign x_4324 = x_660 & x_661;
assign x_4325 = x_659 & x_4324;
assign x_4326 = x_662 & x_663;
assign x_4327 = x_664 & x_665;
assign x_4328 = x_4326 & x_4327;
assign x_4329 = x_4325 & x_4328;
assign x_4330 = x_667 & x_668;
assign x_4331 = x_666 & x_4330;
assign x_4332 = x_669 & x_670;
assign x_4333 = x_671 & x_672;
assign x_4334 = x_4332 & x_4333;
assign x_4335 = x_4331 & x_4334;
assign x_4336 = x_4329 & x_4335;
assign x_4337 = x_674 & x_675;
assign x_4338 = x_673 & x_4337;
assign x_4339 = x_676 & x_677;
assign x_4340 = x_678 & x_679;
assign x_4341 = x_4339 & x_4340;
assign x_4342 = x_4338 & x_4341;
assign x_4343 = x_680 & x_681;
assign x_4344 = x_682 & x_683;
assign x_4345 = x_4343 & x_4344;
assign x_4346 = x_684 & x_685;
assign x_4347 = x_686 & x_687;
assign x_4348 = x_4346 & x_4347;
assign x_4349 = x_4345 & x_4348;
assign x_4350 = x_4342 & x_4349;
assign x_4351 = x_4336 & x_4350;
assign x_4352 = x_4323 & x_4351;
assign x_4353 = x_4295 & x_4352;
assign x_4354 = x_4239 & x_4353;
assign x_4355 = x_689 & x_690;
assign x_4356 = x_688 & x_4355;
assign x_4357 = x_691 & x_692;
assign x_4358 = x_693 & x_694;
assign x_4359 = x_4357 & x_4358;
assign x_4360 = x_4356 & x_4359;
assign x_4361 = x_696 & x_697;
assign x_4362 = x_695 & x_4361;
assign x_4363 = x_698 & x_699;
assign x_4364 = x_700 & x_701;
assign x_4365 = x_4363 & x_4364;
assign x_4366 = x_4362 & x_4365;
assign x_4367 = x_4360 & x_4366;
assign x_4368 = x_703 & x_704;
assign x_4369 = x_702 & x_4368;
assign x_4370 = x_705 & x_706;
assign x_4371 = x_707 & x_708;
assign x_4372 = x_4370 & x_4371;
assign x_4373 = x_4369 & x_4372;
assign x_4374 = x_710 & x_711;
assign x_4375 = x_709 & x_4374;
assign x_4376 = x_712 & x_713;
assign x_4377 = x_714 & x_715;
assign x_4378 = x_4376 & x_4377;
assign x_4379 = x_4375 & x_4378;
assign x_4380 = x_4373 & x_4379;
assign x_4381 = x_4367 & x_4380;
assign x_4382 = x_717 & x_718;
assign x_4383 = x_716 & x_4382;
assign x_4384 = x_719 & x_720;
assign x_4385 = x_721 & x_722;
assign x_4386 = x_4384 & x_4385;
assign x_4387 = x_4383 & x_4386;
assign x_4388 = x_724 & x_725;
assign x_4389 = x_723 & x_4388;
assign x_4390 = x_726 & x_727;
assign x_4391 = x_728 & x_729;
assign x_4392 = x_4390 & x_4391;
assign x_4393 = x_4389 & x_4392;
assign x_4394 = x_4387 & x_4393;
assign x_4395 = x_731 & x_732;
assign x_4396 = x_730 & x_4395;
assign x_4397 = x_733 & x_734;
assign x_4398 = x_735 & x_736;
assign x_4399 = x_4397 & x_4398;
assign x_4400 = x_4396 & x_4399;
assign x_4401 = x_737 & x_738;
assign x_4402 = x_739 & x_740;
assign x_4403 = x_4401 & x_4402;
assign x_4404 = x_741 & x_742;
assign x_4405 = x_743 & x_744;
assign x_4406 = x_4404 & x_4405;
assign x_4407 = x_4403 & x_4406;
assign x_4408 = x_4400 & x_4407;
assign x_4409 = x_4394 & x_4408;
assign x_4410 = x_4381 & x_4409;
assign x_4411 = x_746 & x_747;
assign x_4412 = x_745 & x_4411;
assign x_4413 = x_748 & x_749;
assign x_4414 = x_750 & x_751;
assign x_4415 = x_4413 & x_4414;
assign x_4416 = x_4412 & x_4415;
assign x_4417 = x_753 & x_754;
assign x_4418 = x_752 & x_4417;
assign x_4419 = x_755 & x_756;
assign x_4420 = x_757 & x_758;
assign x_4421 = x_4419 & x_4420;
assign x_4422 = x_4418 & x_4421;
assign x_4423 = x_4416 & x_4422;
assign x_4424 = x_760 & x_761;
assign x_4425 = x_759 & x_4424;
assign x_4426 = x_762 & x_763;
assign x_4427 = x_764 & x_765;
assign x_4428 = x_4426 & x_4427;
assign x_4429 = x_4425 & x_4428;
assign x_4430 = x_766 & x_767;
assign x_4431 = x_768 & x_769;
assign x_4432 = x_4430 & x_4431;
assign x_4433 = x_770 & x_771;
assign x_4434 = x_772 & x_773;
assign x_4435 = x_4433 & x_4434;
assign x_4436 = x_4432 & x_4435;
assign x_4437 = x_4429 & x_4436;
assign x_4438 = x_4423 & x_4437;
assign x_4439 = x_775 & x_776;
assign x_4440 = x_774 & x_4439;
assign x_4441 = x_777 & x_778;
assign x_4442 = x_779 & x_780;
assign x_4443 = x_4441 & x_4442;
assign x_4444 = x_4440 & x_4443;
assign x_4445 = x_782 & x_783;
assign x_4446 = x_781 & x_4445;
assign x_4447 = x_784 & x_785;
assign x_4448 = x_786 & x_787;
assign x_4449 = x_4447 & x_4448;
assign x_4450 = x_4446 & x_4449;
assign x_4451 = x_4444 & x_4450;
assign x_4452 = x_789 & x_790;
assign x_4453 = x_788 & x_4452;
assign x_4454 = x_791 & x_792;
assign x_4455 = x_793 & x_794;
assign x_4456 = x_4454 & x_4455;
assign x_4457 = x_4453 & x_4456;
assign x_4458 = x_795 & x_796;
assign x_4459 = x_797 & x_798;
assign x_4460 = x_4458 & x_4459;
assign x_4461 = x_799 & x_800;
assign x_4462 = x_801 & x_802;
assign x_4463 = x_4461 & x_4462;
assign x_4464 = x_4460 & x_4463;
assign x_4465 = x_4457 & x_4464;
assign x_4466 = x_4451 & x_4465;
assign x_4467 = x_4438 & x_4466;
assign x_4468 = x_4410 & x_4467;
assign x_4469 = x_804 & x_805;
assign x_4470 = x_803 & x_4469;
assign x_4471 = x_806 & x_807;
assign x_4472 = x_808 & x_809;
assign x_4473 = x_4471 & x_4472;
assign x_4474 = x_4470 & x_4473;
assign x_4475 = x_811 & x_812;
assign x_4476 = x_810 & x_4475;
assign x_4477 = x_813 & x_814;
assign x_4478 = x_815 & x_816;
assign x_4479 = x_4477 & x_4478;
assign x_4480 = x_4476 & x_4479;
assign x_4481 = x_4474 & x_4480;
assign x_4482 = x_818 & x_819;
assign x_4483 = x_817 & x_4482;
assign x_4484 = x_820 & x_821;
assign x_4485 = x_822 & x_823;
assign x_4486 = x_4484 & x_4485;
assign x_4487 = x_4483 & x_4486;
assign x_4488 = x_825 & x_826;
assign x_4489 = x_824 & x_4488;
assign x_4490 = x_827 & x_828;
assign x_4491 = x_829 & x_830;
assign x_4492 = x_4490 & x_4491;
assign x_4493 = x_4489 & x_4492;
assign x_4494 = x_4487 & x_4493;
assign x_4495 = x_4481 & x_4494;
assign x_4496 = x_832 & x_833;
assign x_4497 = x_831 & x_4496;
assign x_4498 = x_834 & x_835;
assign x_4499 = x_836 & x_837;
assign x_4500 = x_4498 & x_4499;
assign x_4501 = x_4497 & x_4500;
assign x_4502 = x_839 & x_840;
assign x_4503 = x_838 & x_4502;
assign x_4504 = x_841 & x_842;
assign x_4505 = x_843 & x_844;
assign x_4506 = x_4504 & x_4505;
assign x_4507 = x_4503 & x_4506;
assign x_4508 = x_4501 & x_4507;
assign x_4509 = x_846 & x_847;
assign x_4510 = x_845 & x_4509;
assign x_4511 = x_848 & x_849;
assign x_4512 = x_850 & x_851;
assign x_4513 = x_4511 & x_4512;
assign x_4514 = x_4510 & x_4513;
assign x_4515 = x_852 & x_853;
assign x_4516 = x_854 & x_855;
assign x_4517 = x_4515 & x_4516;
assign x_4518 = x_856 & x_857;
assign x_4519 = x_858 & x_859;
assign x_4520 = x_4518 & x_4519;
assign x_4521 = x_4517 & x_4520;
assign x_4522 = x_4514 & x_4521;
assign x_4523 = x_4508 & x_4522;
assign x_4524 = x_4495 & x_4523;
assign x_4525 = x_861 & x_862;
assign x_4526 = x_860 & x_4525;
assign x_4527 = x_863 & x_864;
assign x_4528 = x_865 & x_866;
assign x_4529 = x_4527 & x_4528;
assign x_4530 = x_4526 & x_4529;
assign x_4531 = x_868 & x_869;
assign x_4532 = x_867 & x_4531;
assign x_4533 = x_870 & x_871;
assign x_4534 = x_872 & x_873;
assign x_4535 = x_4533 & x_4534;
assign x_4536 = x_4532 & x_4535;
assign x_4537 = x_4530 & x_4536;
assign x_4538 = x_875 & x_876;
assign x_4539 = x_874 & x_4538;
assign x_4540 = x_877 & x_878;
assign x_4541 = x_879 & x_880;
assign x_4542 = x_4540 & x_4541;
assign x_4543 = x_4539 & x_4542;
assign x_4544 = x_881 & x_882;
assign x_4545 = x_883 & x_884;
assign x_4546 = x_4544 & x_4545;
assign x_4547 = x_885 & x_886;
assign x_4548 = x_887 & x_888;
assign x_4549 = x_4547 & x_4548;
assign x_4550 = x_4546 & x_4549;
assign x_4551 = x_4543 & x_4550;
assign x_4552 = x_4537 & x_4551;
assign x_4553 = x_890 & x_891;
assign x_4554 = x_889 & x_4553;
assign x_4555 = x_892 & x_893;
assign x_4556 = x_894 & x_895;
assign x_4557 = x_4555 & x_4556;
assign x_4558 = x_4554 & x_4557;
assign x_4559 = x_897 & x_898;
assign x_4560 = x_896 & x_4559;
assign x_4561 = x_899 & x_900;
assign x_4562 = x_901 & x_902;
assign x_4563 = x_4561 & x_4562;
assign x_4564 = x_4560 & x_4563;
assign x_4565 = x_4558 & x_4564;
assign x_4566 = x_904 & x_905;
assign x_4567 = x_903 & x_4566;
assign x_4568 = x_906 & x_907;
assign x_4569 = x_908 & x_909;
assign x_4570 = x_4568 & x_4569;
assign x_4571 = x_4567 & x_4570;
assign x_4572 = x_910 & x_911;
assign x_4573 = x_912 & x_913;
assign x_4574 = x_4572 & x_4573;
assign x_4575 = x_914 & x_915;
assign x_4576 = x_916 & x_917;
assign x_4577 = x_4575 & x_4576;
assign x_4578 = x_4574 & x_4577;
assign x_4579 = x_4571 & x_4578;
assign x_4580 = x_4565 & x_4579;
assign x_4581 = x_4552 & x_4580;
assign x_4582 = x_4524 & x_4581;
assign x_4583 = x_4468 & x_4582;
assign x_4584 = x_4354 & x_4583;
assign x_4585 = x_4126 & x_4584;
assign x_4586 = x_919 & x_920;
assign x_4587 = x_918 & x_4586;
assign x_4588 = x_921 & x_922;
assign x_4589 = x_923 & x_924;
assign x_4590 = x_4588 & x_4589;
assign x_4591 = x_4587 & x_4590;
assign x_4592 = x_926 & x_927;
assign x_4593 = x_925 & x_4592;
assign x_4594 = x_928 & x_929;
assign x_4595 = x_930 & x_931;
assign x_4596 = x_4594 & x_4595;
assign x_4597 = x_4593 & x_4596;
assign x_4598 = x_4591 & x_4597;
assign x_4599 = x_933 & x_934;
assign x_4600 = x_932 & x_4599;
assign x_4601 = x_935 & x_936;
assign x_4602 = x_937 & x_938;
assign x_4603 = x_4601 & x_4602;
assign x_4604 = x_4600 & x_4603;
assign x_4605 = x_940 & x_941;
assign x_4606 = x_939 & x_4605;
assign x_4607 = x_942 & x_943;
assign x_4608 = x_944 & x_945;
assign x_4609 = x_4607 & x_4608;
assign x_4610 = x_4606 & x_4609;
assign x_4611 = x_4604 & x_4610;
assign x_4612 = x_4598 & x_4611;
assign x_4613 = x_947 & x_948;
assign x_4614 = x_946 & x_4613;
assign x_4615 = x_949 & x_950;
assign x_4616 = x_951 & x_952;
assign x_4617 = x_4615 & x_4616;
assign x_4618 = x_4614 & x_4617;
assign x_4619 = x_954 & x_955;
assign x_4620 = x_953 & x_4619;
assign x_4621 = x_956 & x_957;
assign x_4622 = x_958 & x_959;
assign x_4623 = x_4621 & x_4622;
assign x_4624 = x_4620 & x_4623;
assign x_4625 = x_4618 & x_4624;
assign x_4626 = x_961 & x_962;
assign x_4627 = x_960 & x_4626;
assign x_4628 = x_963 & x_964;
assign x_4629 = x_965 & x_966;
assign x_4630 = x_4628 & x_4629;
assign x_4631 = x_4627 & x_4630;
assign x_4632 = x_967 & x_968;
assign x_4633 = x_969 & x_970;
assign x_4634 = x_4632 & x_4633;
assign x_4635 = x_971 & x_972;
assign x_4636 = x_973 & x_974;
assign x_4637 = x_4635 & x_4636;
assign x_4638 = x_4634 & x_4637;
assign x_4639 = x_4631 & x_4638;
assign x_4640 = x_4625 & x_4639;
assign x_4641 = x_4612 & x_4640;
assign x_4642 = x_976 & x_977;
assign x_4643 = x_975 & x_4642;
assign x_4644 = x_978 & x_979;
assign x_4645 = x_980 & x_981;
assign x_4646 = x_4644 & x_4645;
assign x_4647 = x_4643 & x_4646;
assign x_4648 = x_983 & x_984;
assign x_4649 = x_982 & x_4648;
assign x_4650 = x_985 & x_986;
assign x_4651 = x_987 & x_988;
assign x_4652 = x_4650 & x_4651;
assign x_4653 = x_4649 & x_4652;
assign x_4654 = x_4647 & x_4653;
assign x_4655 = x_990 & x_991;
assign x_4656 = x_989 & x_4655;
assign x_4657 = x_992 & x_993;
assign x_4658 = x_994 & x_995;
assign x_4659 = x_4657 & x_4658;
assign x_4660 = x_4656 & x_4659;
assign x_4661 = x_997 & x_998;
assign x_4662 = x_996 & x_4661;
assign x_4663 = x_999 & x_1000;
assign x_4664 = x_1001 & x_1002;
assign x_4665 = x_4663 & x_4664;
assign x_4666 = x_4662 & x_4665;
assign x_4667 = x_4660 & x_4666;
assign x_4668 = x_4654 & x_4667;
assign x_4669 = x_1004 & x_1005;
assign x_4670 = x_1003 & x_4669;
assign x_4671 = x_1006 & x_1007;
assign x_4672 = x_1008 & x_1009;
assign x_4673 = x_4671 & x_4672;
assign x_4674 = x_4670 & x_4673;
assign x_4675 = x_1011 & x_1012;
assign x_4676 = x_1010 & x_4675;
assign x_4677 = x_1013 & x_1014;
assign x_4678 = x_1015 & x_1016;
assign x_4679 = x_4677 & x_4678;
assign x_4680 = x_4676 & x_4679;
assign x_4681 = x_4674 & x_4680;
assign x_4682 = x_1018 & x_1019;
assign x_4683 = x_1017 & x_4682;
assign x_4684 = x_1020 & x_1021;
assign x_4685 = x_1022 & x_1023;
assign x_4686 = x_4684 & x_4685;
assign x_4687 = x_4683 & x_4686;
assign x_4688 = x_1024 & x_1025;
assign x_4689 = x_1026 & x_1027;
assign x_4690 = x_4688 & x_4689;
assign x_4691 = x_1028 & x_1029;
assign x_4692 = x_1030 & x_1031;
assign x_4693 = x_4691 & x_4692;
assign x_4694 = x_4690 & x_4693;
assign x_4695 = x_4687 & x_4694;
assign x_4696 = x_4681 & x_4695;
assign x_4697 = x_4668 & x_4696;
assign x_4698 = x_4641 & x_4697;
assign x_4699 = x_1033 & x_1034;
assign x_4700 = x_1032 & x_4699;
assign x_4701 = x_1035 & x_1036;
assign x_4702 = x_1037 & x_1038;
assign x_4703 = x_4701 & x_4702;
assign x_4704 = x_4700 & x_4703;
assign x_4705 = x_1040 & x_1041;
assign x_4706 = x_1039 & x_4705;
assign x_4707 = x_1042 & x_1043;
assign x_4708 = x_1044 & x_1045;
assign x_4709 = x_4707 & x_4708;
assign x_4710 = x_4706 & x_4709;
assign x_4711 = x_4704 & x_4710;
assign x_4712 = x_1047 & x_1048;
assign x_4713 = x_1046 & x_4712;
assign x_4714 = x_1049 & x_1050;
assign x_4715 = x_1051 & x_1052;
assign x_4716 = x_4714 & x_4715;
assign x_4717 = x_4713 & x_4716;
assign x_4718 = x_1054 & x_1055;
assign x_4719 = x_1053 & x_4718;
assign x_4720 = x_1056 & x_1057;
assign x_4721 = x_1058 & x_1059;
assign x_4722 = x_4720 & x_4721;
assign x_4723 = x_4719 & x_4722;
assign x_4724 = x_4717 & x_4723;
assign x_4725 = x_4711 & x_4724;
assign x_4726 = x_1061 & x_1062;
assign x_4727 = x_1060 & x_4726;
assign x_4728 = x_1063 & x_1064;
assign x_4729 = x_1065 & x_1066;
assign x_4730 = x_4728 & x_4729;
assign x_4731 = x_4727 & x_4730;
assign x_4732 = x_1068 & x_1069;
assign x_4733 = x_1067 & x_4732;
assign x_4734 = x_1070 & x_1071;
assign x_4735 = x_1072 & x_1073;
assign x_4736 = x_4734 & x_4735;
assign x_4737 = x_4733 & x_4736;
assign x_4738 = x_4731 & x_4737;
assign x_4739 = x_1075 & x_1076;
assign x_4740 = x_1074 & x_4739;
assign x_4741 = x_1077 & x_1078;
assign x_4742 = x_1079 & x_1080;
assign x_4743 = x_4741 & x_4742;
assign x_4744 = x_4740 & x_4743;
assign x_4745 = x_1081 & x_1082;
assign x_4746 = x_1083 & x_1084;
assign x_4747 = x_4745 & x_4746;
assign x_4748 = x_1085 & x_1086;
assign x_4749 = x_1087 & x_1088;
assign x_4750 = x_4748 & x_4749;
assign x_4751 = x_4747 & x_4750;
assign x_4752 = x_4744 & x_4751;
assign x_4753 = x_4738 & x_4752;
assign x_4754 = x_4725 & x_4753;
assign x_4755 = x_1090 & x_1091;
assign x_4756 = x_1089 & x_4755;
assign x_4757 = x_1092 & x_1093;
assign x_4758 = x_1094 & x_1095;
assign x_4759 = x_4757 & x_4758;
assign x_4760 = x_4756 & x_4759;
assign x_4761 = x_1097 & x_1098;
assign x_4762 = x_1096 & x_4761;
assign x_4763 = x_1099 & x_1100;
assign x_4764 = x_1101 & x_1102;
assign x_4765 = x_4763 & x_4764;
assign x_4766 = x_4762 & x_4765;
assign x_4767 = x_4760 & x_4766;
assign x_4768 = x_1104 & x_1105;
assign x_4769 = x_1103 & x_4768;
assign x_4770 = x_1106 & x_1107;
assign x_4771 = x_1108 & x_1109;
assign x_4772 = x_4770 & x_4771;
assign x_4773 = x_4769 & x_4772;
assign x_4774 = x_1110 & x_1111;
assign x_4775 = x_1112 & x_1113;
assign x_4776 = x_4774 & x_4775;
assign x_4777 = x_1114 & x_1115;
assign x_4778 = x_1116 & x_1117;
assign x_4779 = x_4777 & x_4778;
assign x_4780 = x_4776 & x_4779;
assign x_4781 = x_4773 & x_4780;
assign x_4782 = x_4767 & x_4781;
assign x_4783 = x_1119 & x_1120;
assign x_4784 = x_1118 & x_4783;
assign x_4785 = x_1121 & x_1122;
assign x_4786 = x_1123 & x_1124;
assign x_4787 = x_4785 & x_4786;
assign x_4788 = x_4784 & x_4787;
assign x_4789 = x_1126 & x_1127;
assign x_4790 = x_1125 & x_4789;
assign x_4791 = x_1128 & x_1129;
assign x_4792 = x_1130 & x_1131;
assign x_4793 = x_4791 & x_4792;
assign x_4794 = x_4790 & x_4793;
assign x_4795 = x_4788 & x_4794;
assign x_4796 = x_1133 & x_1134;
assign x_4797 = x_1132 & x_4796;
assign x_4798 = x_1135 & x_1136;
assign x_4799 = x_1137 & x_1138;
assign x_4800 = x_4798 & x_4799;
assign x_4801 = x_4797 & x_4800;
assign x_4802 = x_1139 & x_1140;
assign x_4803 = x_1141 & x_1142;
assign x_4804 = x_4802 & x_4803;
assign x_4805 = x_1143 & x_1144;
assign x_4806 = x_1145 & x_1146;
assign x_4807 = x_4805 & x_4806;
assign x_4808 = x_4804 & x_4807;
assign x_4809 = x_4801 & x_4808;
assign x_4810 = x_4795 & x_4809;
assign x_4811 = x_4782 & x_4810;
assign x_4812 = x_4754 & x_4811;
assign x_4813 = x_4698 & x_4812;
assign x_4814 = x_1148 & x_1149;
assign x_4815 = x_1147 & x_4814;
assign x_4816 = x_1150 & x_1151;
assign x_4817 = x_1152 & x_1153;
assign x_4818 = x_4816 & x_4817;
assign x_4819 = x_4815 & x_4818;
assign x_4820 = x_1155 & x_1156;
assign x_4821 = x_1154 & x_4820;
assign x_4822 = x_1157 & x_1158;
assign x_4823 = x_1159 & x_1160;
assign x_4824 = x_4822 & x_4823;
assign x_4825 = x_4821 & x_4824;
assign x_4826 = x_4819 & x_4825;
assign x_4827 = x_1162 & x_1163;
assign x_4828 = x_1161 & x_4827;
assign x_4829 = x_1164 & x_1165;
assign x_4830 = x_1166 & x_1167;
assign x_4831 = x_4829 & x_4830;
assign x_4832 = x_4828 & x_4831;
assign x_4833 = x_1169 & x_1170;
assign x_4834 = x_1168 & x_4833;
assign x_4835 = x_1171 & x_1172;
assign x_4836 = x_1173 & x_1174;
assign x_4837 = x_4835 & x_4836;
assign x_4838 = x_4834 & x_4837;
assign x_4839 = x_4832 & x_4838;
assign x_4840 = x_4826 & x_4839;
assign x_4841 = x_1176 & x_1177;
assign x_4842 = x_1175 & x_4841;
assign x_4843 = x_1178 & x_1179;
assign x_4844 = x_1180 & x_1181;
assign x_4845 = x_4843 & x_4844;
assign x_4846 = x_4842 & x_4845;
assign x_4847 = x_1183 & x_1184;
assign x_4848 = x_1182 & x_4847;
assign x_4849 = x_1185 & x_1186;
assign x_4850 = x_1187 & x_1188;
assign x_4851 = x_4849 & x_4850;
assign x_4852 = x_4848 & x_4851;
assign x_4853 = x_4846 & x_4852;
assign x_4854 = x_1190 & x_1191;
assign x_4855 = x_1189 & x_4854;
assign x_4856 = x_1192 & x_1193;
assign x_4857 = x_1194 & x_1195;
assign x_4858 = x_4856 & x_4857;
assign x_4859 = x_4855 & x_4858;
assign x_4860 = x_1196 & x_1197;
assign x_4861 = x_1198 & x_1199;
assign x_4862 = x_4860 & x_4861;
assign x_4863 = x_1200 & x_1201;
assign x_4864 = x_1202 & x_1203;
assign x_4865 = x_4863 & x_4864;
assign x_4866 = x_4862 & x_4865;
assign x_4867 = x_4859 & x_4866;
assign x_4868 = x_4853 & x_4867;
assign x_4869 = x_4840 & x_4868;
assign x_4870 = x_1205 & x_1206;
assign x_4871 = x_1204 & x_4870;
assign x_4872 = x_1207 & x_1208;
assign x_4873 = x_1209 & x_1210;
assign x_4874 = x_4872 & x_4873;
assign x_4875 = x_4871 & x_4874;
assign x_4876 = x_1212 & x_1213;
assign x_4877 = x_1211 & x_4876;
assign x_4878 = x_1214 & x_1215;
assign x_4879 = x_1216 & x_1217;
assign x_4880 = x_4878 & x_4879;
assign x_4881 = x_4877 & x_4880;
assign x_4882 = x_4875 & x_4881;
assign x_4883 = x_1219 & x_1220;
assign x_4884 = x_1218 & x_4883;
assign x_4885 = x_1221 & x_1222;
assign x_4886 = x_1223 & x_1224;
assign x_4887 = x_4885 & x_4886;
assign x_4888 = x_4884 & x_4887;
assign x_4889 = x_1226 & x_1227;
assign x_4890 = x_1225 & x_4889;
assign x_4891 = x_1228 & x_1229;
assign x_4892 = x_1230 & x_1231;
assign x_4893 = x_4891 & x_4892;
assign x_4894 = x_4890 & x_4893;
assign x_4895 = x_4888 & x_4894;
assign x_4896 = x_4882 & x_4895;
assign x_4897 = x_1233 & x_1234;
assign x_4898 = x_1232 & x_4897;
assign x_4899 = x_1235 & x_1236;
assign x_4900 = x_1237 & x_1238;
assign x_4901 = x_4899 & x_4900;
assign x_4902 = x_4898 & x_4901;
assign x_4903 = x_1240 & x_1241;
assign x_4904 = x_1239 & x_4903;
assign x_4905 = x_1242 & x_1243;
assign x_4906 = x_1244 & x_1245;
assign x_4907 = x_4905 & x_4906;
assign x_4908 = x_4904 & x_4907;
assign x_4909 = x_4902 & x_4908;
assign x_4910 = x_1247 & x_1248;
assign x_4911 = x_1246 & x_4910;
assign x_4912 = x_1249 & x_1250;
assign x_4913 = x_1251 & x_1252;
assign x_4914 = x_4912 & x_4913;
assign x_4915 = x_4911 & x_4914;
assign x_4916 = x_1253 & x_1254;
assign x_4917 = x_1255 & x_1256;
assign x_4918 = x_4916 & x_4917;
assign x_4919 = x_1257 & x_1258;
assign x_4920 = x_1259 & x_1260;
assign x_4921 = x_4919 & x_4920;
assign x_4922 = x_4918 & x_4921;
assign x_4923 = x_4915 & x_4922;
assign x_4924 = x_4909 & x_4923;
assign x_4925 = x_4896 & x_4924;
assign x_4926 = x_4869 & x_4925;
assign x_4927 = x_1262 & x_1263;
assign x_4928 = x_1261 & x_4927;
assign x_4929 = x_1264 & x_1265;
assign x_4930 = x_1266 & x_1267;
assign x_4931 = x_4929 & x_4930;
assign x_4932 = x_4928 & x_4931;
assign x_4933 = x_1269 & x_1270;
assign x_4934 = x_1268 & x_4933;
assign x_4935 = x_1271 & x_1272;
assign x_4936 = x_1273 & x_1274;
assign x_4937 = x_4935 & x_4936;
assign x_4938 = x_4934 & x_4937;
assign x_4939 = x_4932 & x_4938;
assign x_4940 = x_1276 & x_1277;
assign x_4941 = x_1275 & x_4940;
assign x_4942 = x_1278 & x_1279;
assign x_4943 = x_1280 & x_1281;
assign x_4944 = x_4942 & x_4943;
assign x_4945 = x_4941 & x_4944;
assign x_4946 = x_1283 & x_1284;
assign x_4947 = x_1282 & x_4946;
assign x_4948 = x_1285 & x_1286;
assign x_4949 = x_1287 & x_1288;
assign x_4950 = x_4948 & x_4949;
assign x_4951 = x_4947 & x_4950;
assign x_4952 = x_4945 & x_4951;
assign x_4953 = x_4939 & x_4952;
assign x_4954 = x_1290 & x_1291;
assign x_4955 = x_1289 & x_4954;
assign x_4956 = x_1292 & x_1293;
assign x_4957 = x_1294 & x_1295;
assign x_4958 = x_4956 & x_4957;
assign x_4959 = x_4955 & x_4958;
assign x_4960 = x_1297 & x_1298;
assign x_4961 = x_1296 & x_4960;
assign x_4962 = x_1299 & x_1300;
assign x_4963 = x_1301 & x_1302;
assign x_4964 = x_4962 & x_4963;
assign x_4965 = x_4961 & x_4964;
assign x_4966 = x_4959 & x_4965;
assign x_4967 = x_1304 & x_1305;
assign x_4968 = x_1303 & x_4967;
assign x_4969 = x_1306 & x_1307;
assign x_4970 = x_1308 & x_1309;
assign x_4971 = x_4969 & x_4970;
assign x_4972 = x_4968 & x_4971;
assign x_4973 = x_1310 & x_1311;
assign x_4974 = x_1312 & x_1313;
assign x_4975 = x_4973 & x_4974;
assign x_4976 = x_1314 & x_1315;
assign x_4977 = x_1316 & x_1317;
assign x_4978 = x_4976 & x_4977;
assign x_4979 = x_4975 & x_4978;
assign x_4980 = x_4972 & x_4979;
assign x_4981 = x_4966 & x_4980;
assign x_4982 = x_4953 & x_4981;
assign x_4983 = x_1319 & x_1320;
assign x_4984 = x_1318 & x_4983;
assign x_4985 = x_1321 & x_1322;
assign x_4986 = x_1323 & x_1324;
assign x_4987 = x_4985 & x_4986;
assign x_4988 = x_4984 & x_4987;
assign x_4989 = x_1326 & x_1327;
assign x_4990 = x_1325 & x_4989;
assign x_4991 = x_1328 & x_1329;
assign x_4992 = x_1330 & x_1331;
assign x_4993 = x_4991 & x_4992;
assign x_4994 = x_4990 & x_4993;
assign x_4995 = x_4988 & x_4994;
assign x_4996 = x_1333 & x_1334;
assign x_4997 = x_1332 & x_4996;
assign x_4998 = x_1335 & x_1336;
assign x_4999 = x_1337 & x_1338;
assign x_5000 = x_4998 & x_4999;
assign x_5001 = x_4997 & x_5000;
assign x_5002 = x_1339 & x_1340;
assign x_5003 = x_1341 & x_1342;
assign x_5004 = x_5002 & x_5003;
assign x_5005 = x_1343 & x_1344;
assign x_5006 = x_1345 & x_1346;
assign x_5007 = x_5005 & x_5006;
assign x_5008 = x_5004 & x_5007;
assign x_5009 = x_5001 & x_5008;
assign x_5010 = x_4995 & x_5009;
assign x_5011 = x_1348 & x_1349;
assign x_5012 = x_1347 & x_5011;
assign x_5013 = x_1350 & x_1351;
assign x_5014 = x_1352 & x_1353;
assign x_5015 = x_5013 & x_5014;
assign x_5016 = x_5012 & x_5015;
assign x_5017 = x_1355 & x_1356;
assign x_5018 = x_1354 & x_5017;
assign x_5019 = x_1357 & x_1358;
assign x_5020 = x_1359 & x_1360;
assign x_5021 = x_5019 & x_5020;
assign x_5022 = x_5018 & x_5021;
assign x_5023 = x_5016 & x_5022;
assign x_5024 = x_1362 & x_1363;
assign x_5025 = x_1361 & x_5024;
assign x_5026 = x_1364 & x_1365;
assign x_5027 = x_1366 & x_1367;
assign x_5028 = x_5026 & x_5027;
assign x_5029 = x_5025 & x_5028;
assign x_5030 = x_1368 & x_1369;
assign x_5031 = x_1370 & x_1371;
assign x_5032 = x_5030 & x_5031;
assign x_5033 = x_1372 & x_1373;
assign x_5034 = x_1374 & x_1375;
assign x_5035 = x_5033 & x_5034;
assign x_5036 = x_5032 & x_5035;
assign x_5037 = x_5029 & x_5036;
assign x_5038 = x_5023 & x_5037;
assign x_5039 = x_5010 & x_5038;
assign x_5040 = x_4982 & x_5039;
assign x_5041 = x_4926 & x_5040;
assign x_5042 = x_4813 & x_5041;
assign x_5043 = x_1377 & x_1378;
assign x_5044 = x_1376 & x_5043;
assign x_5045 = x_1379 & x_1380;
assign x_5046 = x_1381 & x_1382;
assign x_5047 = x_5045 & x_5046;
assign x_5048 = x_5044 & x_5047;
assign x_5049 = x_1384 & x_1385;
assign x_5050 = x_1383 & x_5049;
assign x_5051 = x_1386 & x_1387;
assign x_5052 = x_1388 & x_1389;
assign x_5053 = x_5051 & x_5052;
assign x_5054 = x_5050 & x_5053;
assign x_5055 = x_5048 & x_5054;
assign x_5056 = x_1391 & x_1392;
assign x_5057 = x_1390 & x_5056;
assign x_5058 = x_1393 & x_1394;
assign x_5059 = x_1395 & x_1396;
assign x_5060 = x_5058 & x_5059;
assign x_5061 = x_5057 & x_5060;
assign x_5062 = x_1398 & x_1399;
assign x_5063 = x_1397 & x_5062;
assign x_5064 = x_1400 & x_1401;
assign x_5065 = x_1402 & x_1403;
assign x_5066 = x_5064 & x_5065;
assign x_5067 = x_5063 & x_5066;
assign x_5068 = x_5061 & x_5067;
assign x_5069 = x_5055 & x_5068;
assign x_5070 = x_1405 & x_1406;
assign x_5071 = x_1404 & x_5070;
assign x_5072 = x_1407 & x_1408;
assign x_5073 = x_1409 & x_1410;
assign x_5074 = x_5072 & x_5073;
assign x_5075 = x_5071 & x_5074;
assign x_5076 = x_1412 & x_1413;
assign x_5077 = x_1411 & x_5076;
assign x_5078 = x_1414 & x_1415;
assign x_5079 = x_1416 & x_1417;
assign x_5080 = x_5078 & x_5079;
assign x_5081 = x_5077 & x_5080;
assign x_5082 = x_5075 & x_5081;
assign x_5083 = x_1419 & x_1420;
assign x_5084 = x_1418 & x_5083;
assign x_5085 = x_1421 & x_1422;
assign x_5086 = x_1423 & x_1424;
assign x_5087 = x_5085 & x_5086;
assign x_5088 = x_5084 & x_5087;
assign x_5089 = x_1425 & x_1426;
assign x_5090 = x_1427 & x_1428;
assign x_5091 = x_5089 & x_5090;
assign x_5092 = x_1429 & x_1430;
assign x_5093 = x_1431 & x_1432;
assign x_5094 = x_5092 & x_5093;
assign x_5095 = x_5091 & x_5094;
assign x_5096 = x_5088 & x_5095;
assign x_5097 = x_5082 & x_5096;
assign x_5098 = x_5069 & x_5097;
assign x_5099 = x_1434 & x_1435;
assign x_5100 = x_1433 & x_5099;
assign x_5101 = x_1436 & x_1437;
assign x_5102 = x_1438 & x_1439;
assign x_5103 = x_5101 & x_5102;
assign x_5104 = x_5100 & x_5103;
assign x_5105 = x_1441 & x_1442;
assign x_5106 = x_1440 & x_5105;
assign x_5107 = x_1443 & x_1444;
assign x_5108 = x_1445 & x_1446;
assign x_5109 = x_5107 & x_5108;
assign x_5110 = x_5106 & x_5109;
assign x_5111 = x_5104 & x_5110;
assign x_5112 = x_1448 & x_1449;
assign x_5113 = x_1447 & x_5112;
assign x_5114 = x_1450 & x_1451;
assign x_5115 = x_1452 & x_1453;
assign x_5116 = x_5114 & x_5115;
assign x_5117 = x_5113 & x_5116;
assign x_5118 = x_1455 & x_1456;
assign x_5119 = x_1454 & x_5118;
assign x_5120 = x_1457 & x_1458;
assign x_5121 = x_1459 & x_1460;
assign x_5122 = x_5120 & x_5121;
assign x_5123 = x_5119 & x_5122;
assign x_5124 = x_5117 & x_5123;
assign x_5125 = x_5111 & x_5124;
assign x_5126 = x_1462 & x_1463;
assign x_5127 = x_1461 & x_5126;
assign x_5128 = x_1464 & x_1465;
assign x_5129 = x_1466 & x_1467;
assign x_5130 = x_5128 & x_5129;
assign x_5131 = x_5127 & x_5130;
assign x_5132 = x_1469 & x_1470;
assign x_5133 = x_1468 & x_5132;
assign x_5134 = x_1471 & x_1472;
assign x_5135 = x_1473 & x_1474;
assign x_5136 = x_5134 & x_5135;
assign x_5137 = x_5133 & x_5136;
assign x_5138 = x_5131 & x_5137;
assign x_5139 = x_1476 & x_1477;
assign x_5140 = x_1475 & x_5139;
assign x_5141 = x_1478 & x_1479;
assign x_5142 = x_1480 & x_1481;
assign x_5143 = x_5141 & x_5142;
assign x_5144 = x_5140 & x_5143;
assign x_5145 = x_1482 & x_1483;
assign x_5146 = x_1484 & x_1485;
assign x_5147 = x_5145 & x_5146;
assign x_5148 = x_1486 & x_1487;
assign x_5149 = x_1488 & x_1489;
assign x_5150 = x_5148 & x_5149;
assign x_5151 = x_5147 & x_5150;
assign x_5152 = x_5144 & x_5151;
assign x_5153 = x_5138 & x_5152;
assign x_5154 = x_5125 & x_5153;
assign x_5155 = x_5098 & x_5154;
assign x_5156 = x_1491 & x_1492;
assign x_5157 = x_1490 & x_5156;
assign x_5158 = x_1493 & x_1494;
assign x_5159 = x_1495 & x_1496;
assign x_5160 = x_5158 & x_5159;
assign x_5161 = x_5157 & x_5160;
assign x_5162 = x_1498 & x_1499;
assign x_5163 = x_1497 & x_5162;
assign x_5164 = x_1500 & x_1501;
assign x_5165 = x_1502 & x_1503;
assign x_5166 = x_5164 & x_5165;
assign x_5167 = x_5163 & x_5166;
assign x_5168 = x_5161 & x_5167;
assign x_5169 = x_1505 & x_1506;
assign x_5170 = x_1504 & x_5169;
assign x_5171 = x_1507 & x_1508;
assign x_5172 = x_1509 & x_1510;
assign x_5173 = x_5171 & x_5172;
assign x_5174 = x_5170 & x_5173;
assign x_5175 = x_1512 & x_1513;
assign x_5176 = x_1511 & x_5175;
assign x_5177 = x_1514 & x_1515;
assign x_5178 = x_1516 & x_1517;
assign x_5179 = x_5177 & x_5178;
assign x_5180 = x_5176 & x_5179;
assign x_5181 = x_5174 & x_5180;
assign x_5182 = x_5168 & x_5181;
assign x_5183 = x_1519 & x_1520;
assign x_5184 = x_1518 & x_5183;
assign x_5185 = x_1521 & x_1522;
assign x_5186 = x_1523 & x_1524;
assign x_5187 = x_5185 & x_5186;
assign x_5188 = x_5184 & x_5187;
assign x_5189 = x_1526 & x_1527;
assign x_5190 = x_1525 & x_5189;
assign x_5191 = x_1528 & x_1529;
assign x_5192 = x_1530 & x_1531;
assign x_5193 = x_5191 & x_5192;
assign x_5194 = x_5190 & x_5193;
assign x_5195 = x_5188 & x_5194;
assign x_5196 = x_1533 & x_1534;
assign x_5197 = x_1532 & x_5196;
assign x_5198 = x_1535 & x_1536;
assign x_5199 = x_1537 & x_1538;
assign x_5200 = x_5198 & x_5199;
assign x_5201 = x_5197 & x_5200;
assign x_5202 = x_1539 & x_1540;
assign x_5203 = x_1541 & x_1542;
assign x_5204 = x_5202 & x_5203;
assign x_5205 = x_1543 & x_1544;
assign x_5206 = x_1545 & x_1546;
assign x_5207 = x_5205 & x_5206;
assign x_5208 = x_5204 & x_5207;
assign x_5209 = x_5201 & x_5208;
assign x_5210 = x_5195 & x_5209;
assign x_5211 = x_5182 & x_5210;
assign x_5212 = x_1548 & x_1549;
assign x_5213 = x_1547 & x_5212;
assign x_5214 = x_1550 & x_1551;
assign x_5215 = x_1552 & x_1553;
assign x_5216 = x_5214 & x_5215;
assign x_5217 = x_5213 & x_5216;
assign x_5218 = x_1555 & x_1556;
assign x_5219 = x_1554 & x_5218;
assign x_5220 = x_1557 & x_1558;
assign x_5221 = x_1559 & x_1560;
assign x_5222 = x_5220 & x_5221;
assign x_5223 = x_5219 & x_5222;
assign x_5224 = x_5217 & x_5223;
assign x_5225 = x_1562 & x_1563;
assign x_5226 = x_1561 & x_5225;
assign x_5227 = x_1564 & x_1565;
assign x_5228 = x_1566 & x_1567;
assign x_5229 = x_5227 & x_5228;
assign x_5230 = x_5226 & x_5229;
assign x_5231 = x_1568 & x_1569;
assign x_5232 = x_1570 & x_1571;
assign x_5233 = x_5231 & x_5232;
assign x_5234 = x_1572 & x_1573;
assign x_5235 = x_1574 & x_1575;
assign x_5236 = x_5234 & x_5235;
assign x_5237 = x_5233 & x_5236;
assign x_5238 = x_5230 & x_5237;
assign x_5239 = x_5224 & x_5238;
assign x_5240 = x_1577 & x_1578;
assign x_5241 = x_1576 & x_5240;
assign x_5242 = x_1579 & x_1580;
assign x_5243 = x_1581 & x_1582;
assign x_5244 = x_5242 & x_5243;
assign x_5245 = x_5241 & x_5244;
assign x_5246 = x_1584 & x_1585;
assign x_5247 = x_1583 & x_5246;
assign x_5248 = x_1586 & x_1587;
assign x_5249 = x_1588 & x_1589;
assign x_5250 = x_5248 & x_5249;
assign x_5251 = x_5247 & x_5250;
assign x_5252 = x_5245 & x_5251;
assign x_5253 = x_1591 & x_1592;
assign x_5254 = x_1590 & x_5253;
assign x_5255 = x_1593 & x_1594;
assign x_5256 = x_1595 & x_1596;
assign x_5257 = x_5255 & x_5256;
assign x_5258 = x_5254 & x_5257;
assign x_5259 = x_1597 & x_1598;
assign x_5260 = x_1599 & x_1600;
assign x_5261 = x_5259 & x_5260;
assign x_5262 = x_1601 & x_1602;
assign x_5263 = x_1603 & x_1604;
assign x_5264 = x_5262 & x_5263;
assign x_5265 = x_5261 & x_5264;
assign x_5266 = x_5258 & x_5265;
assign x_5267 = x_5252 & x_5266;
assign x_5268 = x_5239 & x_5267;
assign x_5269 = x_5211 & x_5268;
assign x_5270 = x_5155 & x_5269;
assign x_5271 = x_1606 & x_1607;
assign x_5272 = x_1605 & x_5271;
assign x_5273 = x_1608 & x_1609;
assign x_5274 = x_1610 & x_1611;
assign x_5275 = x_5273 & x_5274;
assign x_5276 = x_5272 & x_5275;
assign x_5277 = x_1613 & x_1614;
assign x_5278 = x_1612 & x_5277;
assign x_5279 = x_1615 & x_1616;
assign x_5280 = x_1617 & x_1618;
assign x_5281 = x_5279 & x_5280;
assign x_5282 = x_5278 & x_5281;
assign x_5283 = x_5276 & x_5282;
assign x_5284 = x_1620 & x_1621;
assign x_5285 = x_1619 & x_5284;
assign x_5286 = x_1622 & x_1623;
assign x_5287 = x_1624 & x_1625;
assign x_5288 = x_5286 & x_5287;
assign x_5289 = x_5285 & x_5288;
assign x_5290 = x_1627 & x_1628;
assign x_5291 = x_1626 & x_5290;
assign x_5292 = x_1629 & x_1630;
assign x_5293 = x_1631 & x_1632;
assign x_5294 = x_5292 & x_5293;
assign x_5295 = x_5291 & x_5294;
assign x_5296 = x_5289 & x_5295;
assign x_5297 = x_5283 & x_5296;
assign x_5298 = x_1634 & x_1635;
assign x_5299 = x_1633 & x_5298;
assign x_5300 = x_1636 & x_1637;
assign x_5301 = x_1638 & x_1639;
assign x_5302 = x_5300 & x_5301;
assign x_5303 = x_5299 & x_5302;
assign x_5304 = x_1641 & x_1642;
assign x_5305 = x_1640 & x_5304;
assign x_5306 = x_1643 & x_1644;
assign x_5307 = x_1645 & x_1646;
assign x_5308 = x_5306 & x_5307;
assign x_5309 = x_5305 & x_5308;
assign x_5310 = x_5303 & x_5309;
assign x_5311 = x_1648 & x_1649;
assign x_5312 = x_1647 & x_5311;
assign x_5313 = x_1650 & x_1651;
assign x_5314 = x_1652 & x_1653;
assign x_5315 = x_5313 & x_5314;
assign x_5316 = x_5312 & x_5315;
assign x_5317 = x_1654 & x_1655;
assign x_5318 = x_1656 & x_1657;
assign x_5319 = x_5317 & x_5318;
assign x_5320 = x_1658 & x_1659;
assign x_5321 = x_1660 & x_1661;
assign x_5322 = x_5320 & x_5321;
assign x_5323 = x_5319 & x_5322;
assign x_5324 = x_5316 & x_5323;
assign x_5325 = x_5310 & x_5324;
assign x_5326 = x_5297 & x_5325;
assign x_5327 = x_1663 & x_1664;
assign x_5328 = x_1662 & x_5327;
assign x_5329 = x_1665 & x_1666;
assign x_5330 = x_1667 & x_1668;
assign x_5331 = x_5329 & x_5330;
assign x_5332 = x_5328 & x_5331;
assign x_5333 = x_1670 & x_1671;
assign x_5334 = x_1669 & x_5333;
assign x_5335 = x_1672 & x_1673;
assign x_5336 = x_1674 & x_1675;
assign x_5337 = x_5335 & x_5336;
assign x_5338 = x_5334 & x_5337;
assign x_5339 = x_5332 & x_5338;
assign x_5340 = x_1677 & x_1678;
assign x_5341 = x_1676 & x_5340;
assign x_5342 = x_1679 & x_1680;
assign x_5343 = x_1681 & x_1682;
assign x_5344 = x_5342 & x_5343;
assign x_5345 = x_5341 & x_5344;
assign x_5346 = x_1683 & x_1684;
assign x_5347 = x_1685 & x_1686;
assign x_5348 = x_5346 & x_5347;
assign x_5349 = x_1687 & x_1688;
assign x_5350 = x_1689 & x_1690;
assign x_5351 = x_5349 & x_5350;
assign x_5352 = x_5348 & x_5351;
assign x_5353 = x_5345 & x_5352;
assign x_5354 = x_5339 & x_5353;
assign x_5355 = x_1692 & x_1693;
assign x_5356 = x_1691 & x_5355;
assign x_5357 = x_1694 & x_1695;
assign x_5358 = x_1696 & x_1697;
assign x_5359 = x_5357 & x_5358;
assign x_5360 = x_5356 & x_5359;
assign x_5361 = x_1699 & x_1700;
assign x_5362 = x_1698 & x_5361;
assign x_5363 = x_1701 & x_1702;
assign x_5364 = x_1703 & x_1704;
assign x_5365 = x_5363 & x_5364;
assign x_5366 = x_5362 & x_5365;
assign x_5367 = x_5360 & x_5366;
assign x_5368 = x_1706 & x_1707;
assign x_5369 = x_1705 & x_5368;
assign x_5370 = x_1708 & x_1709;
assign x_5371 = x_1710 & x_1711;
assign x_5372 = x_5370 & x_5371;
assign x_5373 = x_5369 & x_5372;
assign x_5374 = x_1712 & x_1713;
assign x_5375 = x_1714 & x_1715;
assign x_5376 = x_5374 & x_5375;
assign x_5377 = x_1716 & x_1717;
assign x_5378 = x_1718 & x_1719;
assign x_5379 = x_5377 & x_5378;
assign x_5380 = x_5376 & x_5379;
assign x_5381 = x_5373 & x_5380;
assign x_5382 = x_5367 & x_5381;
assign x_5383 = x_5354 & x_5382;
assign x_5384 = x_5326 & x_5383;
assign x_5385 = x_1721 & x_1722;
assign x_5386 = x_1720 & x_5385;
assign x_5387 = x_1723 & x_1724;
assign x_5388 = x_1725 & x_1726;
assign x_5389 = x_5387 & x_5388;
assign x_5390 = x_5386 & x_5389;
assign x_5391 = x_1728 & x_1729;
assign x_5392 = x_1727 & x_5391;
assign x_5393 = x_1730 & x_1731;
assign x_5394 = x_1732 & x_1733;
assign x_5395 = x_5393 & x_5394;
assign x_5396 = x_5392 & x_5395;
assign x_5397 = x_5390 & x_5396;
assign x_5398 = x_1735 & x_1736;
assign x_5399 = x_1734 & x_5398;
assign x_5400 = x_1737 & x_1738;
assign x_5401 = x_1739 & x_1740;
assign x_5402 = x_5400 & x_5401;
assign x_5403 = x_5399 & x_5402;
assign x_5404 = x_1742 & x_1743;
assign x_5405 = x_1741 & x_5404;
assign x_5406 = x_1744 & x_1745;
assign x_5407 = x_1746 & x_1747;
assign x_5408 = x_5406 & x_5407;
assign x_5409 = x_5405 & x_5408;
assign x_5410 = x_5403 & x_5409;
assign x_5411 = x_5397 & x_5410;
assign x_5412 = x_1749 & x_1750;
assign x_5413 = x_1748 & x_5412;
assign x_5414 = x_1751 & x_1752;
assign x_5415 = x_1753 & x_1754;
assign x_5416 = x_5414 & x_5415;
assign x_5417 = x_5413 & x_5416;
assign x_5418 = x_1756 & x_1757;
assign x_5419 = x_1755 & x_5418;
assign x_5420 = x_1758 & x_1759;
assign x_5421 = x_1760 & x_1761;
assign x_5422 = x_5420 & x_5421;
assign x_5423 = x_5419 & x_5422;
assign x_5424 = x_5417 & x_5423;
assign x_5425 = x_1763 & x_1764;
assign x_5426 = x_1762 & x_5425;
assign x_5427 = x_1765 & x_1766;
assign x_5428 = x_1767 & x_1768;
assign x_5429 = x_5427 & x_5428;
assign x_5430 = x_5426 & x_5429;
assign x_5431 = x_1769 & x_1770;
assign x_5432 = x_1771 & x_1772;
assign x_5433 = x_5431 & x_5432;
assign x_5434 = x_1773 & x_1774;
assign x_5435 = x_1775 & x_1776;
assign x_5436 = x_5434 & x_5435;
assign x_5437 = x_5433 & x_5436;
assign x_5438 = x_5430 & x_5437;
assign x_5439 = x_5424 & x_5438;
assign x_5440 = x_5411 & x_5439;
assign x_5441 = x_1778 & x_1779;
assign x_5442 = x_1777 & x_5441;
assign x_5443 = x_1780 & x_1781;
assign x_5444 = x_1782 & x_1783;
assign x_5445 = x_5443 & x_5444;
assign x_5446 = x_5442 & x_5445;
assign x_5447 = x_1785 & x_1786;
assign x_5448 = x_1784 & x_5447;
assign x_5449 = x_1787 & x_1788;
assign x_5450 = x_1789 & x_1790;
assign x_5451 = x_5449 & x_5450;
assign x_5452 = x_5448 & x_5451;
assign x_5453 = x_5446 & x_5452;
assign x_5454 = x_1792 & x_1793;
assign x_5455 = x_1791 & x_5454;
assign x_5456 = x_1794 & x_1795;
assign x_5457 = x_1796 & x_1797;
assign x_5458 = x_5456 & x_5457;
assign x_5459 = x_5455 & x_5458;
assign x_5460 = x_1798 & x_1799;
assign x_5461 = x_1800 & x_1801;
assign x_5462 = x_5460 & x_5461;
assign x_5463 = x_1802 & x_1803;
assign x_5464 = x_1804 & x_1805;
assign x_5465 = x_5463 & x_5464;
assign x_5466 = x_5462 & x_5465;
assign x_5467 = x_5459 & x_5466;
assign x_5468 = x_5453 & x_5467;
assign x_5469 = x_1807 & x_1808;
assign x_5470 = x_1806 & x_5469;
assign x_5471 = x_1809 & x_1810;
assign x_5472 = x_1811 & x_1812;
assign x_5473 = x_5471 & x_5472;
assign x_5474 = x_5470 & x_5473;
assign x_5475 = x_1814 & x_1815;
assign x_5476 = x_1813 & x_5475;
assign x_5477 = x_1816 & x_1817;
assign x_5478 = x_1818 & x_1819;
assign x_5479 = x_5477 & x_5478;
assign x_5480 = x_5476 & x_5479;
assign x_5481 = x_5474 & x_5480;
assign x_5482 = x_1821 & x_1822;
assign x_5483 = x_1820 & x_5482;
assign x_5484 = x_1823 & x_1824;
assign x_5485 = x_1825 & x_1826;
assign x_5486 = x_5484 & x_5485;
assign x_5487 = x_5483 & x_5486;
assign x_5488 = x_1827 & x_1828;
assign x_5489 = x_1829 & x_1830;
assign x_5490 = x_5488 & x_5489;
assign x_5491 = x_1831 & x_1832;
assign x_5492 = x_1833 & x_1834;
assign x_5493 = x_5491 & x_5492;
assign x_5494 = x_5490 & x_5493;
assign x_5495 = x_5487 & x_5494;
assign x_5496 = x_5481 & x_5495;
assign x_5497 = x_5468 & x_5496;
assign x_5498 = x_5440 & x_5497;
assign x_5499 = x_5384 & x_5498;
assign x_5500 = x_5270 & x_5499;
assign x_5501 = x_5042 & x_5500;
assign x_5502 = x_4585 & x_5501;
assign x_5503 = x_1836 & x_1837;
assign x_5504 = x_1835 & x_5503;
assign x_5505 = x_1838 & x_1839;
assign x_5506 = x_1840 & x_1841;
assign x_5507 = x_5505 & x_5506;
assign x_5508 = x_5504 & x_5507;
assign x_5509 = x_1843 & x_1844;
assign x_5510 = x_1842 & x_5509;
assign x_5511 = x_1845 & x_1846;
assign x_5512 = x_1847 & x_1848;
assign x_5513 = x_5511 & x_5512;
assign x_5514 = x_5510 & x_5513;
assign x_5515 = x_5508 & x_5514;
assign x_5516 = x_1850 & x_1851;
assign x_5517 = x_1849 & x_5516;
assign x_5518 = x_1852 & x_1853;
assign x_5519 = x_1854 & x_1855;
assign x_5520 = x_5518 & x_5519;
assign x_5521 = x_5517 & x_5520;
assign x_5522 = x_1857 & x_1858;
assign x_5523 = x_1856 & x_5522;
assign x_5524 = x_1859 & x_1860;
assign x_5525 = x_1861 & x_1862;
assign x_5526 = x_5524 & x_5525;
assign x_5527 = x_5523 & x_5526;
assign x_5528 = x_5521 & x_5527;
assign x_5529 = x_5515 & x_5528;
assign x_5530 = x_1864 & x_1865;
assign x_5531 = x_1863 & x_5530;
assign x_5532 = x_1866 & x_1867;
assign x_5533 = x_1868 & x_1869;
assign x_5534 = x_5532 & x_5533;
assign x_5535 = x_5531 & x_5534;
assign x_5536 = x_1871 & x_1872;
assign x_5537 = x_1870 & x_5536;
assign x_5538 = x_1873 & x_1874;
assign x_5539 = x_1875 & x_1876;
assign x_5540 = x_5538 & x_5539;
assign x_5541 = x_5537 & x_5540;
assign x_5542 = x_5535 & x_5541;
assign x_5543 = x_1878 & x_1879;
assign x_5544 = x_1877 & x_5543;
assign x_5545 = x_1880 & x_1881;
assign x_5546 = x_1882 & x_1883;
assign x_5547 = x_5545 & x_5546;
assign x_5548 = x_5544 & x_5547;
assign x_5549 = x_1884 & x_1885;
assign x_5550 = x_1886 & x_1887;
assign x_5551 = x_5549 & x_5550;
assign x_5552 = x_1888 & x_1889;
assign x_5553 = x_1890 & x_1891;
assign x_5554 = x_5552 & x_5553;
assign x_5555 = x_5551 & x_5554;
assign x_5556 = x_5548 & x_5555;
assign x_5557 = x_5542 & x_5556;
assign x_5558 = x_5529 & x_5557;
assign x_5559 = x_1893 & x_1894;
assign x_5560 = x_1892 & x_5559;
assign x_5561 = x_1895 & x_1896;
assign x_5562 = x_1897 & x_1898;
assign x_5563 = x_5561 & x_5562;
assign x_5564 = x_5560 & x_5563;
assign x_5565 = x_1900 & x_1901;
assign x_5566 = x_1899 & x_5565;
assign x_5567 = x_1902 & x_1903;
assign x_5568 = x_1904 & x_1905;
assign x_5569 = x_5567 & x_5568;
assign x_5570 = x_5566 & x_5569;
assign x_5571 = x_5564 & x_5570;
assign x_5572 = x_1907 & x_1908;
assign x_5573 = x_1906 & x_5572;
assign x_5574 = x_1909 & x_1910;
assign x_5575 = x_1911 & x_1912;
assign x_5576 = x_5574 & x_5575;
assign x_5577 = x_5573 & x_5576;
assign x_5578 = x_1914 & x_1915;
assign x_5579 = x_1913 & x_5578;
assign x_5580 = x_1916 & x_1917;
assign x_5581 = x_1918 & x_1919;
assign x_5582 = x_5580 & x_5581;
assign x_5583 = x_5579 & x_5582;
assign x_5584 = x_5577 & x_5583;
assign x_5585 = x_5571 & x_5584;
assign x_5586 = x_1921 & x_1922;
assign x_5587 = x_1920 & x_5586;
assign x_5588 = x_1923 & x_1924;
assign x_5589 = x_1925 & x_1926;
assign x_5590 = x_5588 & x_5589;
assign x_5591 = x_5587 & x_5590;
assign x_5592 = x_1928 & x_1929;
assign x_5593 = x_1927 & x_5592;
assign x_5594 = x_1930 & x_1931;
assign x_5595 = x_1932 & x_1933;
assign x_5596 = x_5594 & x_5595;
assign x_5597 = x_5593 & x_5596;
assign x_5598 = x_5591 & x_5597;
assign x_5599 = x_1935 & x_1936;
assign x_5600 = x_1934 & x_5599;
assign x_5601 = x_1937 & x_1938;
assign x_5602 = x_1939 & x_1940;
assign x_5603 = x_5601 & x_5602;
assign x_5604 = x_5600 & x_5603;
assign x_5605 = x_1941 & x_1942;
assign x_5606 = x_1943 & x_1944;
assign x_5607 = x_5605 & x_5606;
assign x_5608 = x_1945 & x_1946;
assign x_5609 = x_1947 & x_1948;
assign x_5610 = x_5608 & x_5609;
assign x_5611 = x_5607 & x_5610;
assign x_5612 = x_5604 & x_5611;
assign x_5613 = x_5598 & x_5612;
assign x_5614 = x_5585 & x_5613;
assign x_5615 = x_5558 & x_5614;
assign x_5616 = x_1950 & x_1951;
assign x_5617 = x_1949 & x_5616;
assign x_5618 = x_1952 & x_1953;
assign x_5619 = x_1954 & x_1955;
assign x_5620 = x_5618 & x_5619;
assign x_5621 = x_5617 & x_5620;
assign x_5622 = x_1957 & x_1958;
assign x_5623 = x_1956 & x_5622;
assign x_5624 = x_1959 & x_1960;
assign x_5625 = x_1961 & x_1962;
assign x_5626 = x_5624 & x_5625;
assign x_5627 = x_5623 & x_5626;
assign x_5628 = x_5621 & x_5627;
assign x_5629 = x_1964 & x_1965;
assign x_5630 = x_1963 & x_5629;
assign x_5631 = x_1966 & x_1967;
assign x_5632 = x_1968 & x_1969;
assign x_5633 = x_5631 & x_5632;
assign x_5634 = x_5630 & x_5633;
assign x_5635 = x_1971 & x_1972;
assign x_5636 = x_1970 & x_5635;
assign x_5637 = x_1973 & x_1974;
assign x_5638 = x_1975 & x_1976;
assign x_5639 = x_5637 & x_5638;
assign x_5640 = x_5636 & x_5639;
assign x_5641 = x_5634 & x_5640;
assign x_5642 = x_5628 & x_5641;
assign x_5643 = x_1978 & x_1979;
assign x_5644 = x_1977 & x_5643;
assign x_5645 = x_1980 & x_1981;
assign x_5646 = x_1982 & x_1983;
assign x_5647 = x_5645 & x_5646;
assign x_5648 = x_5644 & x_5647;
assign x_5649 = x_1985 & x_1986;
assign x_5650 = x_1984 & x_5649;
assign x_5651 = x_1987 & x_1988;
assign x_5652 = x_1989 & x_1990;
assign x_5653 = x_5651 & x_5652;
assign x_5654 = x_5650 & x_5653;
assign x_5655 = x_5648 & x_5654;
assign x_5656 = x_1992 & x_1993;
assign x_5657 = x_1991 & x_5656;
assign x_5658 = x_1994 & x_1995;
assign x_5659 = x_1996 & x_1997;
assign x_5660 = x_5658 & x_5659;
assign x_5661 = x_5657 & x_5660;
assign x_5662 = x_1998 & x_1999;
assign x_5663 = x_2000 & x_2001;
assign x_5664 = x_5662 & x_5663;
assign x_5665 = x_2002 & x_2003;
assign x_5666 = x_2004 & x_2005;
assign x_5667 = x_5665 & x_5666;
assign x_5668 = x_5664 & x_5667;
assign x_5669 = x_5661 & x_5668;
assign x_5670 = x_5655 & x_5669;
assign x_5671 = x_5642 & x_5670;
assign x_5672 = x_2007 & x_2008;
assign x_5673 = x_2006 & x_5672;
assign x_5674 = x_2009 & x_2010;
assign x_5675 = x_2011 & x_2012;
assign x_5676 = x_5674 & x_5675;
assign x_5677 = x_5673 & x_5676;
assign x_5678 = x_2014 & x_2015;
assign x_5679 = x_2013 & x_5678;
assign x_5680 = x_2016 & x_2017;
assign x_5681 = x_2018 & x_2019;
assign x_5682 = x_5680 & x_5681;
assign x_5683 = x_5679 & x_5682;
assign x_5684 = x_5677 & x_5683;
assign x_5685 = x_2021 & x_2022;
assign x_5686 = x_2020 & x_5685;
assign x_5687 = x_2023 & x_2024;
assign x_5688 = x_2025 & x_2026;
assign x_5689 = x_5687 & x_5688;
assign x_5690 = x_5686 & x_5689;
assign x_5691 = x_2027 & x_2028;
assign x_5692 = x_2029 & x_2030;
assign x_5693 = x_5691 & x_5692;
assign x_5694 = x_2031 & x_2032;
assign x_5695 = x_2033 & x_2034;
assign x_5696 = x_5694 & x_5695;
assign x_5697 = x_5693 & x_5696;
assign x_5698 = x_5690 & x_5697;
assign x_5699 = x_5684 & x_5698;
assign x_5700 = x_2036 & x_2037;
assign x_5701 = x_2035 & x_5700;
assign x_5702 = x_2038 & x_2039;
assign x_5703 = x_2040 & x_2041;
assign x_5704 = x_5702 & x_5703;
assign x_5705 = x_5701 & x_5704;
assign x_5706 = x_2043 & x_2044;
assign x_5707 = x_2042 & x_5706;
assign x_5708 = x_2045 & x_2046;
assign x_5709 = x_2047 & x_2048;
assign x_5710 = x_5708 & x_5709;
assign x_5711 = x_5707 & x_5710;
assign x_5712 = x_5705 & x_5711;
assign x_5713 = x_2050 & x_2051;
assign x_5714 = x_2049 & x_5713;
assign x_5715 = x_2052 & x_2053;
assign x_5716 = x_2054 & x_2055;
assign x_5717 = x_5715 & x_5716;
assign x_5718 = x_5714 & x_5717;
assign x_5719 = x_2056 & x_2057;
assign x_5720 = x_2058 & x_2059;
assign x_5721 = x_5719 & x_5720;
assign x_5722 = x_2060 & x_2061;
assign x_5723 = x_2062 & x_2063;
assign x_5724 = x_5722 & x_5723;
assign x_5725 = x_5721 & x_5724;
assign x_5726 = x_5718 & x_5725;
assign x_5727 = x_5712 & x_5726;
assign x_5728 = x_5699 & x_5727;
assign x_5729 = x_5671 & x_5728;
assign x_5730 = x_5615 & x_5729;
assign x_5731 = x_2065 & x_2066;
assign x_5732 = x_2064 & x_5731;
assign x_5733 = x_2067 & x_2068;
assign x_5734 = x_2069 & x_2070;
assign x_5735 = x_5733 & x_5734;
assign x_5736 = x_5732 & x_5735;
assign x_5737 = x_2072 & x_2073;
assign x_5738 = x_2071 & x_5737;
assign x_5739 = x_2074 & x_2075;
assign x_5740 = x_2076 & x_2077;
assign x_5741 = x_5739 & x_5740;
assign x_5742 = x_5738 & x_5741;
assign x_5743 = x_5736 & x_5742;
assign x_5744 = x_2079 & x_2080;
assign x_5745 = x_2078 & x_5744;
assign x_5746 = x_2081 & x_2082;
assign x_5747 = x_2083 & x_2084;
assign x_5748 = x_5746 & x_5747;
assign x_5749 = x_5745 & x_5748;
assign x_5750 = x_2086 & x_2087;
assign x_5751 = x_2085 & x_5750;
assign x_5752 = x_2088 & x_2089;
assign x_5753 = x_2090 & x_2091;
assign x_5754 = x_5752 & x_5753;
assign x_5755 = x_5751 & x_5754;
assign x_5756 = x_5749 & x_5755;
assign x_5757 = x_5743 & x_5756;
assign x_5758 = x_2093 & x_2094;
assign x_5759 = x_2092 & x_5758;
assign x_5760 = x_2095 & x_2096;
assign x_5761 = x_2097 & x_2098;
assign x_5762 = x_5760 & x_5761;
assign x_5763 = x_5759 & x_5762;
assign x_5764 = x_2100 & x_2101;
assign x_5765 = x_2099 & x_5764;
assign x_5766 = x_2102 & x_2103;
assign x_5767 = x_2104 & x_2105;
assign x_5768 = x_5766 & x_5767;
assign x_5769 = x_5765 & x_5768;
assign x_5770 = x_5763 & x_5769;
assign x_5771 = x_2107 & x_2108;
assign x_5772 = x_2106 & x_5771;
assign x_5773 = x_2109 & x_2110;
assign x_5774 = x_2111 & x_2112;
assign x_5775 = x_5773 & x_5774;
assign x_5776 = x_5772 & x_5775;
assign x_5777 = x_2113 & x_2114;
assign x_5778 = x_2115 & x_2116;
assign x_5779 = x_5777 & x_5778;
assign x_5780 = x_2117 & x_2118;
assign x_5781 = x_2119 & x_2120;
assign x_5782 = x_5780 & x_5781;
assign x_5783 = x_5779 & x_5782;
assign x_5784 = x_5776 & x_5783;
assign x_5785 = x_5770 & x_5784;
assign x_5786 = x_5757 & x_5785;
assign x_5787 = x_2122 & x_2123;
assign x_5788 = x_2121 & x_5787;
assign x_5789 = x_2124 & x_2125;
assign x_5790 = x_2126 & x_2127;
assign x_5791 = x_5789 & x_5790;
assign x_5792 = x_5788 & x_5791;
assign x_5793 = x_2129 & x_2130;
assign x_5794 = x_2128 & x_5793;
assign x_5795 = x_2131 & x_2132;
assign x_5796 = x_2133 & x_2134;
assign x_5797 = x_5795 & x_5796;
assign x_5798 = x_5794 & x_5797;
assign x_5799 = x_5792 & x_5798;
assign x_5800 = x_2136 & x_2137;
assign x_5801 = x_2135 & x_5800;
assign x_5802 = x_2138 & x_2139;
assign x_5803 = x_2140 & x_2141;
assign x_5804 = x_5802 & x_5803;
assign x_5805 = x_5801 & x_5804;
assign x_5806 = x_2143 & x_2144;
assign x_5807 = x_2142 & x_5806;
assign x_5808 = x_2145 & x_2146;
assign x_5809 = x_2147 & x_2148;
assign x_5810 = x_5808 & x_5809;
assign x_5811 = x_5807 & x_5810;
assign x_5812 = x_5805 & x_5811;
assign x_5813 = x_5799 & x_5812;
assign x_5814 = x_2150 & x_2151;
assign x_5815 = x_2149 & x_5814;
assign x_5816 = x_2152 & x_2153;
assign x_5817 = x_2154 & x_2155;
assign x_5818 = x_5816 & x_5817;
assign x_5819 = x_5815 & x_5818;
assign x_5820 = x_2157 & x_2158;
assign x_5821 = x_2156 & x_5820;
assign x_5822 = x_2159 & x_2160;
assign x_5823 = x_2161 & x_2162;
assign x_5824 = x_5822 & x_5823;
assign x_5825 = x_5821 & x_5824;
assign x_5826 = x_5819 & x_5825;
assign x_5827 = x_2164 & x_2165;
assign x_5828 = x_2163 & x_5827;
assign x_5829 = x_2166 & x_2167;
assign x_5830 = x_2168 & x_2169;
assign x_5831 = x_5829 & x_5830;
assign x_5832 = x_5828 & x_5831;
assign x_5833 = x_2170 & x_2171;
assign x_5834 = x_2172 & x_2173;
assign x_5835 = x_5833 & x_5834;
assign x_5836 = x_2174 & x_2175;
assign x_5837 = x_2176 & x_2177;
assign x_5838 = x_5836 & x_5837;
assign x_5839 = x_5835 & x_5838;
assign x_5840 = x_5832 & x_5839;
assign x_5841 = x_5826 & x_5840;
assign x_5842 = x_5813 & x_5841;
assign x_5843 = x_5786 & x_5842;
assign x_5844 = x_2179 & x_2180;
assign x_5845 = x_2178 & x_5844;
assign x_5846 = x_2181 & x_2182;
assign x_5847 = x_2183 & x_2184;
assign x_5848 = x_5846 & x_5847;
assign x_5849 = x_5845 & x_5848;
assign x_5850 = x_2186 & x_2187;
assign x_5851 = x_2185 & x_5850;
assign x_5852 = x_2188 & x_2189;
assign x_5853 = x_2190 & x_2191;
assign x_5854 = x_5852 & x_5853;
assign x_5855 = x_5851 & x_5854;
assign x_5856 = x_5849 & x_5855;
assign x_5857 = x_2193 & x_2194;
assign x_5858 = x_2192 & x_5857;
assign x_5859 = x_2195 & x_2196;
assign x_5860 = x_2197 & x_2198;
assign x_5861 = x_5859 & x_5860;
assign x_5862 = x_5858 & x_5861;
assign x_5863 = x_2200 & x_2201;
assign x_5864 = x_2199 & x_5863;
assign x_5865 = x_2202 & x_2203;
assign x_5866 = x_2204 & x_2205;
assign x_5867 = x_5865 & x_5866;
assign x_5868 = x_5864 & x_5867;
assign x_5869 = x_5862 & x_5868;
assign x_5870 = x_5856 & x_5869;
assign x_5871 = x_2207 & x_2208;
assign x_5872 = x_2206 & x_5871;
assign x_5873 = x_2209 & x_2210;
assign x_5874 = x_2211 & x_2212;
assign x_5875 = x_5873 & x_5874;
assign x_5876 = x_5872 & x_5875;
assign x_5877 = x_2214 & x_2215;
assign x_5878 = x_2213 & x_5877;
assign x_5879 = x_2216 & x_2217;
assign x_5880 = x_2218 & x_2219;
assign x_5881 = x_5879 & x_5880;
assign x_5882 = x_5878 & x_5881;
assign x_5883 = x_5876 & x_5882;
assign x_5884 = x_2221 & x_2222;
assign x_5885 = x_2220 & x_5884;
assign x_5886 = x_2223 & x_2224;
assign x_5887 = x_2225 & x_2226;
assign x_5888 = x_5886 & x_5887;
assign x_5889 = x_5885 & x_5888;
assign x_5890 = x_2227 & x_2228;
assign x_5891 = x_2229 & x_2230;
assign x_5892 = x_5890 & x_5891;
assign x_5893 = x_2231 & x_2232;
assign x_5894 = x_2233 & x_2234;
assign x_5895 = x_5893 & x_5894;
assign x_5896 = x_5892 & x_5895;
assign x_5897 = x_5889 & x_5896;
assign x_5898 = x_5883 & x_5897;
assign x_5899 = x_5870 & x_5898;
assign x_5900 = x_2236 & x_2237;
assign x_5901 = x_2235 & x_5900;
assign x_5902 = x_2238 & x_2239;
assign x_5903 = x_2240 & x_2241;
assign x_5904 = x_5902 & x_5903;
assign x_5905 = x_5901 & x_5904;
assign x_5906 = x_2243 & x_2244;
assign x_5907 = x_2242 & x_5906;
assign x_5908 = x_2245 & x_2246;
assign x_5909 = x_2247 & x_2248;
assign x_5910 = x_5908 & x_5909;
assign x_5911 = x_5907 & x_5910;
assign x_5912 = x_5905 & x_5911;
assign x_5913 = x_2250 & x_2251;
assign x_5914 = x_2249 & x_5913;
assign x_5915 = x_2252 & x_2253;
assign x_5916 = x_2254 & x_2255;
assign x_5917 = x_5915 & x_5916;
assign x_5918 = x_5914 & x_5917;
assign x_5919 = x_2256 & x_2257;
assign x_5920 = x_2258 & x_2259;
assign x_5921 = x_5919 & x_5920;
assign x_5922 = x_2260 & x_2261;
assign x_5923 = x_2262 & x_2263;
assign x_5924 = x_5922 & x_5923;
assign x_5925 = x_5921 & x_5924;
assign x_5926 = x_5918 & x_5925;
assign x_5927 = x_5912 & x_5926;
assign x_5928 = x_2265 & x_2266;
assign x_5929 = x_2264 & x_5928;
assign x_5930 = x_2267 & x_2268;
assign x_5931 = x_2269 & x_2270;
assign x_5932 = x_5930 & x_5931;
assign x_5933 = x_5929 & x_5932;
assign x_5934 = x_2272 & x_2273;
assign x_5935 = x_2271 & x_5934;
assign x_5936 = x_2274 & x_2275;
assign x_5937 = x_2276 & x_2277;
assign x_5938 = x_5936 & x_5937;
assign x_5939 = x_5935 & x_5938;
assign x_5940 = x_5933 & x_5939;
assign x_5941 = x_2279 & x_2280;
assign x_5942 = x_2278 & x_5941;
assign x_5943 = x_2281 & x_2282;
assign x_5944 = x_2283 & x_2284;
assign x_5945 = x_5943 & x_5944;
assign x_5946 = x_5942 & x_5945;
assign x_5947 = x_2285 & x_2286;
assign x_5948 = x_2287 & x_2288;
assign x_5949 = x_5947 & x_5948;
assign x_5950 = x_2289 & x_2290;
assign x_5951 = x_2291 & x_2292;
assign x_5952 = x_5950 & x_5951;
assign x_5953 = x_5949 & x_5952;
assign x_5954 = x_5946 & x_5953;
assign x_5955 = x_5940 & x_5954;
assign x_5956 = x_5927 & x_5955;
assign x_5957 = x_5899 & x_5956;
assign x_5958 = x_5843 & x_5957;
assign x_5959 = x_5730 & x_5958;
assign x_5960 = x_2294 & x_2295;
assign x_5961 = x_2293 & x_5960;
assign x_5962 = x_2296 & x_2297;
assign x_5963 = x_2298 & x_2299;
assign x_5964 = x_5962 & x_5963;
assign x_5965 = x_5961 & x_5964;
assign x_5966 = x_2301 & x_2302;
assign x_5967 = x_2300 & x_5966;
assign x_5968 = x_2303 & x_2304;
assign x_5969 = x_2305 & x_2306;
assign x_5970 = x_5968 & x_5969;
assign x_5971 = x_5967 & x_5970;
assign x_5972 = x_5965 & x_5971;
assign x_5973 = x_2308 & x_2309;
assign x_5974 = x_2307 & x_5973;
assign x_5975 = x_2310 & x_2311;
assign x_5976 = x_2312 & x_2313;
assign x_5977 = x_5975 & x_5976;
assign x_5978 = x_5974 & x_5977;
assign x_5979 = x_2315 & x_2316;
assign x_5980 = x_2314 & x_5979;
assign x_5981 = x_2317 & x_2318;
assign x_5982 = x_2319 & x_2320;
assign x_5983 = x_5981 & x_5982;
assign x_5984 = x_5980 & x_5983;
assign x_5985 = x_5978 & x_5984;
assign x_5986 = x_5972 & x_5985;
assign x_5987 = x_2322 & x_2323;
assign x_5988 = x_2321 & x_5987;
assign x_5989 = x_2324 & x_2325;
assign x_5990 = x_2326 & x_2327;
assign x_5991 = x_5989 & x_5990;
assign x_5992 = x_5988 & x_5991;
assign x_5993 = x_2329 & x_2330;
assign x_5994 = x_2328 & x_5993;
assign x_5995 = x_2331 & x_2332;
assign x_5996 = x_2333 & x_2334;
assign x_5997 = x_5995 & x_5996;
assign x_5998 = x_5994 & x_5997;
assign x_5999 = x_5992 & x_5998;
assign x_6000 = x_2336 & x_2337;
assign x_6001 = x_2335 & x_6000;
assign x_6002 = x_2338 & x_2339;
assign x_6003 = x_2340 & x_2341;
assign x_6004 = x_6002 & x_6003;
assign x_6005 = x_6001 & x_6004;
assign x_6006 = x_2342 & x_2343;
assign x_6007 = x_2344 & x_2345;
assign x_6008 = x_6006 & x_6007;
assign x_6009 = x_2346 & x_2347;
assign x_6010 = x_2348 & x_2349;
assign x_6011 = x_6009 & x_6010;
assign x_6012 = x_6008 & x_6011;
assign x_6013 = x_6005 & x_6012;
assign x_6014 = x_5999 & x_6013;
assign x_6015 = x_5986 & x_6014;
assign x_6016 = x_2351 & x_2352;
assign x_6017 = x_2350 & x_6016;
assign x_6018 = x_2353 & x_2354;
assign x_6019 = x_2355 & x_2356;
assign x_6020 = x_6018 & x_6019;
assign x_6021 = x_6017 & x_6020;
assign x_6022 = x_2358 & x_2359;
assign x_6023 = x_2357 & x_6022;
assign x_6024 = x_2360 & x_2361;
assign x_6025 = x_2362 & x_2363;
assign x_6026 = x_6024 & x_6025;
assign x_6027 = x_6023 & x_6026;
assign x_6028 = x_6021 & x_6027;
assign x_6029 = x_2365 & x_2366;
assign x_6030 = x_2364 & x_6029;
assign x_6031 = x_2367 & x_2368;
assign x_6032 = x_2369 & x_2370;
assign x_6033 = x_6031 & x_6032;
assign x_6034 = x_6030 & x_6033;
assign x_6035 = x_2372 & x_2373;
assign x_6036 = x_2371 & x_6035;
assign x_6037 = x_2374 & x_2375;
assign x_6038 = x_2376 & x_2377;
assign x_6039 = x_6037 & x_6038;
assign x_6040 = x_6036 & x_6039;
assign x_6041 = x_6034 & x_6040;
assign x_6042 = x_6028 & x_6041;
assign x_6043 = x_2379 & x_2380;
assign x_6044 = x_2378 & x_6043;
assign x_6045 = x_2381 & x_2382;
assign x_6046 = x_2383 & x_2384;
assign x_6047 = x_6045 & x_6046;
assign x_6048 = x_6044 & x_6047;
assign x_6049 = x_2386 & x_2387;
assign x_6050 = x_2385 & x_6049;
assign x_6051 = x_2388 & x_2389;
assign x_6052 = x_2390 & x_2391;
assign x_6053 = x_6051 & x_6052;
assign x_6054 = x_6050 & x_6053;
assign x_6055 = x_6048 & x_6054;
assign x_6056 = x_2393 & x_2394;
assign x_6057 = x_2392 & x_6056;
assign x_6058 = x_2395 & x_2396;
assign x_6059 = x_2397 & x_2398;
assign x_6060 = x_6058 & x_6059;
assign x_6061 = x_6057 & x_6060;
assign x_6062 = x_2399 & x_2400;
assign x_6063 = x_2401 & x_2402;
assign x_6064 = x_6062 & x_6063;
assign x_6065 = x_2403 & x_2404;
assign x_6066 = x_2405 & x_2406;
assign x_6067 = x_6065 & x_6066;
assign x_6068 = x_6064 & x_6067;
assign x_6069 = x_6061 & x_6068;
assign x_6070 = x_6055 & x_6069;
assign x_6071 = x_6042 & x_6070;
assign x_6072 = x_6015 & x_6071;
assign x_6073 = x_2408 & x_2409;
assign x_6074 = x_2407 & x_6073;
assign x_6075 = x_2410 & x_2411;
assign x_6076 = x_2412 & x_2413;
assign x_6077 = x_6075 & x_6076;
assign x_6078 = x_6074 & x_6077;
assign x_6079 = x_2415 & x_2416;
assign x_6080 = x_2414 & x_6079;
assign x_6081 = x_2417 & x_2418;
assign x_6082 = x_2419 & x_2420;
assign x_6083 = x_6081 & x_6082;
assign x_6084 = x_6080 & x_6083;
assign x_6085 = x_6078 & x_6084;
assign x_6086 = x_2422 & x_2423;
assign x_6087 = x_2421 & x_6086;
assign x_6088 = x_2424 & x_2425;
assign x_6089 = x_2426 & x_2427;
assign x_6090 = x_6088 & x_6089;
assign x_6091 = x_6087 & x_6090;
assign x_6092 = x_2429 & x_2430;
assign x_6093 = x_2428 & x_6092;
assign x_6094 = x_2431 & x_2432;
assign x_6095 = x_2433 & x_2434;
assign x_6096 = x_6094 & x_6095;
assign x_6097 = x_6093 & x_6096;
assign x_6098 = x_6091 & x_6097;
assign x_6099 = x_6085 & x_6098;
assign x_6100 = x_2436 & x_2437;
assign x_6101 = x_2435 & x_6100;
assign x_6102 = x_2438 & x_2439;
assign x_6103 = x_2440 & x_2441;
assign x_6104 = x_6102 & x_6103;
assign x_6105 = x_6101 & x_6104;
assign x_6106 = x_2443 & x_2444;
assign x_6107 = x_2442 & x_6106;
assign x_6108 = x_2445 & x_2446;
assign x_6109 = x_2447 & x_2448;
assign x_6110 = x_6108 & x_6109;
assign x_6111 = x_6107 & x_6110;
assign x_6112 = x_6105 & x_6111;
assign x_6113 = x_2450 & x_2451;
assign x_6114 = x_2449 & x_6113;
assign x_6115 = x_2452 & x_2453;
assign x_6116 = x_2454 & x_2455;
assign x_6117 = x_6115 & x_6116;
assign x_6118 = x_6114 & x_6117;
assign x_6119 = x_2456 & x_2457;
assign x_6120 = x_2458 & x_2459;
assign x_6121 = x_6119 & x_6120;
assign x_6122 = x_2460 & x_2461;
assign x_6123 = x_2462 & x_2463;
assign x_6124 = x_6122 & x_6123;
assign x_6125 = x_6121 & x_6124;
assign x_6126 = x_6118 & x_6125;
assign x_6127 = x_6112 & x_6126;
assign x_6128 = x_6099 & x_6127;
assign x_6129 = x_2465 & x_2466;
assign x_6130 = x_2464 & x_6129;
assign x_6131 = x_2467 & x_2468;
assign x_6132 = x_2469 & x_2470;
assign x_6133 = x_6131 & x_6132;
assign x_6134 = x_6130 & x_6133;
assign x_6135 = x_2472 & x_2473;
assign x_6136 = x_2471 & x_6135;
assign x_6137 = x_2474 & x_2475;
assign x_6138 = x_2476 & x_2477;
assign x_6139 = x_6137 & x_6138;
assign x_6140 = x_6136 & x_6139;
assign x_6141 = x_6134 & x_6140;
assign x_6142 = x_2479 & x_2480;
assign x_6143 = x_2478 & x_6142;
assign x_6144 = x_2481 & x_2482;
assign x_6145 = x_2483 & x_2484;
assign x_6146 = x_6144 & x_6145;
assign x_6147 = x_6143 & x_6146;
assign x_6148 = x_2485 & x_2486;
assign x_6149 = x_2487 & x_2488;
assign x_6150 = x_6148 & x_6149;
assign x_6151 = x_2489 & x_2490;
assign x_6152 = x_2491 & x_2492;
assign x_6153 = x_6151 & x_6152;
assign x_6154 = x_6150 & x_6153;
assign x_6155 = x_6147 & x_6154;
assign x_6156 = x_6141 & x_6155;
assign x_6157 = x_2494 & x_2495;
assign x_6158 = x_2493 & x_6157;
assign x_6159 = x_2496 & x_2497;
assign x_6160 = x_2498 & x_2499;
assign x_6161 = x_6159 & x_6160;
assign x_6162 = x_6158 & x_6161;
assign x_6163 = x_2501 & x_2502;
assign x_6164 = x_2500 & x_6163;
assign x_6165 = x_2503 & x_2504;
assign x_6166 = x_2505 & x_2506;
assign x_6167 = x_6165 & x_6166;
assign x_6168 = x_6164 & x_6167;
assign x_6169 = x_6162 & x_6168;
assign x_6170 = x_2508 & x_2509;
assign x_6171 = x_2507 & x_6170;
assign x_6172 = x_2510 & x_2511;
assign x_6173 = x_2512 & x_2513;
assign x_6174 = x_6172 & x_6173;
assign x_6175 = x_6171 & x_6174;
assign x_6176 = x_2514 & x_2515;
assign x_6177 = x_2516 & x_2517;
assign x_6178 = x_6176 & x_6177;
assign x_6179 = x_2518 & x_2519;
assign x_6180 = x_2520 & x_2521;
assign x_6181 = x_6179 & x_6180;
assign x_6182 = x_6178 & x_6181;
assign x_6183 = x_6175 & x_6182;
assign x_6184 = x_6169 & x_6183;
assign x_6185 = x_6156 & x_6184;
assign x_6186 = x_6128 & x_6185;
assign x_6187 = x_6072 & x_6186;
assign x_6188 = x_2523 & x_2524;
assign x_6189 = x_2522 & x_6188;
assign x_6190 = x_2525 & x_2526;
assign x_6191 = x_2527 & x_2528;
assign x_6192 = x_6190 & x_6191;
assign x_6193 = x_6189 & x_6192;
assign x_6194 = x_2530 & x_2531;
assign x_6195 = x_2529 & x_6194;
assign x_6196 = x_2532 & x_2533;
assign x_6197 = x_2534 & x_2535;
assign x_6198 = x_6196 & x_6197;
assign x_6199 = x_6195 & x_6198;
assign x_6200 = x_6193 & x_6199;
assign x_6201 = x_2537 & x_2538;
assign x_6202 = x_2536 & x_6201;
assign x_6203 = x_2539 & x_2540;
assign x_6204 = x_2541 & x_2542;
assign x_6205 = x_6203 & x_6204;
assign x_6206 = x_6202 & x_6205;
assign x_6207 = x_2544 & x_2545;
assign x_6208 = x_2543 & x_6207;
assign x_6209 = x_2546 & x_2547;
assign x_6210 = x_2548 & x_2549;
assign x_6211 = x_6209 & x_6210;
assign x_6212 = x_6208 & x_6211;
assign x_6213 = x_6206 & x_6212;
assign x_6214 = x_6200 & x_6213;
assign x_6215 = x_2551 & x_2552;
assign x_6216 = x_2550 & x_6215;
assign x_6217 = x_2553 & x_2554;
assign x_6218 = x_2555 & x_2556;
assign x_6219 = x_6217 & x_6218;
assign x_6220 = x_6216 & x_6219;
assign x_6221 = x_2558 & x_2559;
assign x_6222 = x_2557 & x_6221;
assign x_6223 = x_2560 & x_2561;
assign x_6224 = x_2562 & x_2563;
assign x_6225 = x_6223 & x_6224;
assign x_6226 = x_6222 & x_6225;
assign x_6227 = x_6220 & x_6226;
assign x_6228 = x_2565 & x_2566;
assign x_6229 = x_2564 & x_6228;
assign x_6230 = x_2567 & x_2568;
assign x_6231 = x_2569 & x_2570;
assign x_6232 = x_6230 & x_6231;
assign x_6233 = x_6229 & x_6232;
assign x_6234 = x_2571 & x_2572;
assign x_6235 = x_2573 & x_2574;
assign x_6236 = x_6234 & x_6235;
assign x_6237 = x_2575 & x_2576;
assign x_6238 = x_2577 & x_2578;
assign x_6239 = x_6237 & x_6238;
assign x_6240 = x_6236 & x_6239;
assign x_6241 = x_6233 & x_6240;
assign x_6242 = x_6227 & x_6241;
assign x_6243 = x_6214 & x_6242;
assign x_6244 = x_2580 & x_2581;
assign x_6245 = x_2579 & x_6244;
assign x_6246 = x_2582 & x_2583;
assign x_6247 = x_2584 & x_2585;
assign x_6248 = x_6246 & x_6247;
assign x_6249 = x_6245 & x_6248;
assign x_6250 = x_2587 & x_2588;
assign x_6251 = x_2586 & x_6250;
assign x_6252 = x_2589 & x_2590;
assign x_6253 = x_2591 & x_2592;
assign x_6254 = x_6252 & x_6253;
assign x_6255 = x_6251 & x_6254;
assign x_6256 = x_6249 & x_6255;
assign x_6257 = x_2594 & x_2595;
assign x_6258 = x_2593 & x_6257;
assign x_6259 = x_2596 & x_2597;
assign x_6260 = x_2598 & x_2599;
assign x_6261 = x_6259 & x_6260;
assign x_6262 = x_6258 & x_6261;
assign x_6263 = x_2600 & x_2601;
assign x_6264 = x_2602 & x_2603;
assign x_6265 = x_6263 & x_6264;
assign x_6266 = x_2604 & x_2605;
assign x_6267 = x_2606 & x_2607;
assign x_6268 = x_6266 & x_6267;
assign x_6269 = x_6265 & x_6268;
assign x_6270 = x_6262 & x_6269;
assign x_6271 = x_6256 & x_6270;
assign x_6272 = x_2609 & x_2610;
assign x_6273 = x_2608 & x_6272;
assign x_6274 = x_2611 & x_2612;
assign x_6275 = x_2613 & x_2614;
assign x_6276 = x_6274 & x_6275;
assign x_6277 = x_6273 & x_6276;
assign x_6278 = x_2616 & x_2617;
assign x_6279 = x_2615 & x_6278;
assign x_6280 = x_2618 & x_2619;
assign x_6281 = x_2620 & x_2621;
assign x_6282 = x_6280 & x_6281;
assign x_6283 = x_6279 & x_6282;
assign x_6284 = x_6277 & x_6283;
assign x_6285 = x_2623 & x_2624;
assign x_6286 = x_2622 & x_6285;
assign x_6287 = x_2625 & x_2626;
assign x_6288 = x_2627 & x_2628;
assign x_6289 = x_6287 & x_6288;
assign x_6290 = x_6286 & x_6289;
assign x_6291 = x_2629 & x_2630;
assign x_6292 = x_2631 & x_2632;
assign x_6293 = x_6291 & x_6292;
assign x_6294 = x_2633 & x_2634;
assign x_6295 = x_2635 & x_2636;
assign x_6296 = x_6294 & x_6295;
assign x_6297 = x_6293 & x_6296;
assign x_6298 = x_6290 & x_6297;
assign x_6299 = x_6284 & x_6298;
assign x_6300 = x_6271 & x_6299;
assign x_6301 = x_6243 & x_6300;
assign x_6302 = x_2638 & x_2639;
assign x_6303 = x_2637 & x_6302;
assign x_6304 = x_2640 & x_2641;
assign x_6305 = x_2642 & x_2643;
assign x_6306 = x_6304 & x_6305;
assign x_6307 = x_6303 & x_6306;
assign x_6308 = x_2645 & x_2646;
assign x_6309 = x_2644 & x_6308;
assign x_6310 = x_2647 & x_2648;
assign x_6311 = x_2649 & x_2650;
assign x_6312 = x_6310 & x_6311;
assign x_6313 = x_6309 & x_6312;
assign x_6314 = x_6307 & x_6313;
assign x_6315 = x_2652 & x_2653;
assign x_6316 = x_2651 & x_6315;
assign x_6317 = x_2654 & x_2655;
assign x_6318 = x_2656 & x_2657;
assign x_6319 = x_6317 & x_6318;
assign x_6320 = x_6316 & x_6319;
assign x_6321 = x_2659 & x_2660;
assign x_6322 = x_2658 & x_6321;
assign x_6323 = x_2661 & x_2662;
assign x_6324 = x_2663 & x_2664;
assign x_6325 = x_6323 & x_6324;
assign x_6326 = x_6322 & x_6325;
assign x_6327 = x_6320 & x_6326;
assign x_6328 = x_6314 & x_6327;
assign x_6329 = x_2666 & x_2667;
assign x_6330 = x_2665 & x_6329;
assign x_6331 = x_2668 & x_2669;
assign x_6332 = x_2670 & x_2671;
assign x_6333 = x_6331 & x_6332;
assign x_6334 = x_6330 & x_6333;
assign x_6335 = x_2673 & x_2674;
assign x_6336 = x_2672 & x_6335;
assign x_6337 = x_2675 & x_2676;
assign x_6338 = x_2677 & x_2678;
assign x_6339 = x_6337 & x_6338;
assign x_6340 = x_6336 & x_6339;
assign x_6341 = x_6334 & x_6340;
assign x_6342 = x_2680 & x_2681;
assign x_6343 = x_2679 & x_6342;
assign x_6344 = x_2682 & x_2683;
assign x_6345 = x_2684 & x_2685;
assign x_6346 = x_6344 & x_6345;
assign x_6347 = x_6343 & x_6346;
assign x_6348 = x_2686 & x_2687;
assign x_6349 = x_2688 & x_2689;
assign x_6350 = x_6348 & x_6349;
assign x_6351 = x_2690 & x_2691;
assign x_6352 = x_2692 & x_2693;
assign x_6353 = x_6351 & x_6352;
assign x_6354 = x_6350 & x_6353;
assign x_6355 = x_6347 & x_6354;
assign x_6356 = x_6341 & x_6355;
assign x_6357 = x_6328 & x_6356;
assign x_6358 = x_2695 & x_2696;
assign x_6359 = x_2694 & x_6358;
assign x_6360 = x_2697 & x_2698;
assign x_6361 = x_2699 & x_2700;
assign x_6362 = x_6360 & x_6361;
assign x_6363 = x_6359 & x_6362;
assign x_6364 = x_2702 & x_2703;
assign x_6365 = x_2701 & x_6364;
assign x_6366 = x_2704 & x_2705;
assign x_6367 = x_2706 & x_2707;
assign x_6368 = x_6366 & x_6367;
assign x_6369 = x_6365 & x_6368;
assign x_6370 = x_6363 & x_6369;
assign x_6371 = x_2709 & x_2710;
assign x_6372 = x_2708 & x_6371;
assign x_6373 = x_2711 & x_2712;
assign x_6374 = x_2713 & x_2714;
assign x_6375 = x_6373 & x_6374;
assign x_6376 = x_6372 & x_6375;
assign x_6377 = x_2715 & x_2716;
assign x_6378 = x_2717 & x_2718;
assign x_6379 = x_6377 & x_6378;
assign x_6380 = x_2719 & x_2720;
assign x_6381 = x_2721 & x_2722;
assign x_6382 = x_6380 & x_6381;
assign x_6383 = x_6379 & x_6382;
assign x_6384 = x_6376 & x_6383;
assign x_6385 = x_6370 & x_6384;
assign x_6386 = x_2724 & x_2725;
assign x_6387 = x_2723 & x_6386;
assign x_6388 = x_2726 & x_2727;
assign x_6389 = x_2728 & x_2729;
assign x_6390 = x_6388 & x_6389;
assign x_6391 = x_6387 & x_6390;
assign x_6392 = x_2731 & x_2732;
assign x_6393 = x_2730 & x_6392;
assign x_6394 = x_2733 & x_2734;
assign x_6395 = x_2735 & x_2736;
assign x_6396 = x_6394 & x_6395;
assign x_6397 = x_6393 & x_6396;
assign x_6398 = x_6391 & x_6397;
assign x_6399 = x_2738 & x_2739;
assign x_6400 = x_2737 & x_6399;
assign x_6401 = x_2740 & x_2741;
assign x_6402 = x_2742 & x_2743;
assign x_6403 = x_6401 & x_6402;
assign x_6404 = x_6400 & x_6403;
assign x_6405 = x_2744 & x_2745;
assign x_6406 = x_2746 & x_2747;
assign x_6407 = x_6405 & x_6406;
assign x_6408 = x_2748 & x_2749;
assign x_6409 = x_2750 & x_2751;
assign x_6410 = x_6408 & x_6409;
assign x_6411 = x_6407 & x_6410;
assign x_6412 = x_6404 & x_6411;
assign x_6413 = x_6398 & x_6412;
assign x_6414 = x_6385 & x_6413;
assign x_6415 = x_6357 & x_6414;
assign x_6416 = x_6301 & x_6415;
assign x_6417 = x_6187 & x_6416;
assign x_6418 = x_5959 & x_6417;
assign x_6419 = x_2753 & x_2754;
assign x_6420 = x_2752 & x_6419;
assign x_6421 = x_2755 & x_2756;
assign x_6422 = x_2757 & x_2758;
assign x_6423 = x_6421 & x_6422;
assign x_6424 = x_6420 & x_6423;
assign x_6425 = x_2760 & x_2761;
assign x_6426 = x_2759 & x_6425;
assign x_6427 = x_2762 & x_2763;
assign x_6428 = x_2764 & x_2765;
assign x_6429 = x_6427 & x_6428;
assign x_6430 = x_6426 & x_6429;
assign x_6431 = x_6424 & x_6430;
assign x_6432 = x_2767 & x_2768;
assign x_6433 = x_2766 & x_6432;
assign x_6434 = x_2769 & x_2770;
assign x_6435 = x_2771 & x_2772;
assign x_6436 = x_6434 & x_6435;
assign x_6437 = x_6433 & x_6436;
assign x_6438 = x_2774 & x_2775;
assign x_6439 = x_2773 & x_6438;
assign x_6440 = x_2776 & x_2777;
assign x_6441 = x_2778 & x_2779;
assign x_6442 = x_6440 & x_6441;
assign x_6443 = x_6439 & x_6442;
assign x_6444 = x_6437 & x_6443;
assign x_6445 = x_6431 & x_6444;
assign x_6446 = x_2781 & x_2782;
assign x_6447 = x_2780 & x_6446;
assign x_6448 = x_2783 & x_2784;
assign x_6449 = x_2785 & x_2786;
assign x_6450 = x_6448 & x_6449;
assign x_6451 = x_6447 & x_6450;
assign x_6452 = x_2788 & x_2789;
assign x_6453 = x_2787 & x_6452;
assign x_6454 = x_2790 & x_2791;
assign x_6455 = x_2792 & x_2793;
assign x_6456 = x_6454 & x_6455;
assign x_6457 = x_6453 & x_6456;
assign x_6458 = x_6451 & x_6457;
assign x_6459 = x_2795 & x_2796;
assign x_6460 = x_2794 & x_6459;
assign x_6461 = x_2797 & x_2798;
assign x_6462 = x_2799 & x_2800;
assign x_6463 = x_6461 & x_6462;
assign x_6464 = x_6460 & x_6463;
assign x_6465 = x_2801 & x_2802;
assign x_6466 = x_2803 & x_2804;
assign x_6467 = x_6465 & x_6466;
assign x_6468 = x_2805 & x_2806;
assign x_6469 = x_2807 & x_2808;
assign x_6470 = x_6468 & x_6469;
assign x_6471 = x_6467 & x_6470;
assign x_6472 = x_6464 & x_6471;
assign x_6473 = x_6458 & x_6472;
assign x_6474 = x_6445 & x_6473;
assign x_6475 = x_2810 & x_2811;
assign x_6476 = x_2809 & x_6475;
assign x_6477 = x_2812 & x_2813;
assign x_6478 = x_2814 & x_2815;
assign x_6479 = x_6477 & x_6478;
assign x_6480 = x_6476 & x_6479;
assign x_6481 = x_2817 & x_2818;
assign x_6482 = x_2816 & x_6481;
assign x_6483 = x_2819 & x_2820;
assign x_6484 = x_2821 & x_2822;
assign x_6485 = x_6483 & x_6484;
assign x_6486 = x_6482 & x_6485;
assign x_6487 = x_6480 & x_6486;
assign x_6488 = x_2824 & x_2825;
assign x_6489 = x_2823 & x_6488;
assign x_6490 = x_2826 & x_2827;
assign x_6491 = x_2828 & x_2829;
assign x_6492 = x_6490 & x_6491;
assign x_6493 = x_6489 & x_6492;
assign x_6494 = x_2831 & x_2832;
assign x_6495 = x_2830 & x_6494;
assign x_6496 = x_2833 & x_2834;
assign x_6497 = x_2835 & x_2836;
assign x_6498 = x_6496 & x_6497;
assign x_6499 = x_6495 & x_6498;
assign x_6500 = x_6493 & x_6499;
assign x_6501 = x_6487 & x_6500;
assign x_6502 = x_2838 & x_2839;
assign x_6503 = x_2837 & x_6502;
assign x_6504 = x_2840 & x_2841;
assign x_6505 = x_2842 & x_2843;
assign x_6506 = x_6504 & x_6505;
assign x_6507 = x_6503 & x_6506;
assign x_6508 = x_2845 & x_2846;
assign x_6509 = x_2844 & x_6508;
assign x_6510 = x_2847 & x_2848;
assign x_6511 = x_2849 & x_2850;
assign x_6512 = x_6510 & x_6511;
assign x_6513 = x_6509 & x_6512;
assign x_6514 = x_6507 & x_6513;
assign x_6515 = x_2852 & x_2853;
assign x_6516 = x_2851 & x_6515;
assign x_6517 = x_2854 & x_2855;
assign x_6518 = x_2856 & x_2857;
assign x_6519 = x_6517 & x_6518;
assign x_6520 = x_6516 & x_6519;
assign x_6521 = x_2858 & x_2859;
assign x_6522 = x_2860 & x_2861;
assign x_6523 = x_6521 & x_6522;
assign x_6524 = x_2862 & x_2863;
assign x_6525 = x_2864 & x_2865;
assign x_6526 = x_6524 & x_6525;
assign x_6527 = x_6523 & x_6526;
assign x_6528 = x_6520 & x_6527;
assign x_6529 = x_6514 & x_6528;
assign x_6530 = x_6501 & x_6529;
assign x_6531 = x_6474 & x_6530;
assign x_6532 = x_2867 & x_2868;
assign x_6533 = x_2866 & x_6532;
assign x_6534 = x_2869 & x_2870;
assign x_6535 = x_2871 & x_2872;
assign x_6536 = x_6534 & x_6535;
assign x_6537 = x_6533 & x_6536;
assign x_6538 = x_2874 & x_2875;
assign x_6539 = x_2873 & x_6538;
assign x_6540 = x_2876 & x_2877;
assign x_6541 = x_2878 & x_2879;
assign x_6542 = x_6540 & x_6541;
assign x_6543 = x_6539 & x_6542;
assign x_6544 = x_6537 & x_6543;
assign x_6545 = x_2881 & x_2882;
assign x_6546 = x_2880 & x_6545;
assign x_6547 = x_2883 & x_2884;
assign x_6548 = x_2885 & x_2886;
assign x_6549 = x_6547 & x_6548;
assign x_6550 = x_6546 & x_6549;
assign x_6551 = x_2888 & x_2889;
assign x_6552 = x_2887 & x_6551;
assign x_6553 = x_2890 & x_2891;
assign x_6554 = x_2892 & x_2893;
assign x_6555 = x_6553 & x_6554;
assign x_6556 = x_6552 & x_6555;
assign x_6557 = x_6550 & x_6556;
assign x_6558 = x_6544 & x_6557;
assign x_6559 = x_2895 & x_2896;
assign x_6560 = x_2894 & x_6559;
assign x_6561 = x_2897 & x_2898;
assign x_6562 = x_2899 & x_2900;
assign x_6563 = x_6561 & x_6562;
assign x_6564 = x_6560 & x_6563;
assign x_6565 = x_2902 & x_2903;
assign x_6566 = x_2901 & x_6565;
assign x_6567 = x_2904 & x_2905;
assign x_6568 = x_2906 & x_2907;
assign x_6569 = x_6567 & x_6568;
assign x_6570 = x_6566 & x_6569;
assign x_6571 = x_6564 & x_6570;
assign x_6572 = x_2909 & x_2910;
assign x_6573 = x_2908 & x_6572;
assign x_6574 = x_2911 & x_2912;
assign x_6575 = x_2913 & x_2914;
assign x_6576 = x_6574 & x_6575;
assign x_6577 = x_6573 & x_6576;
assign x_6578 = x_2915 & x_2916;
assign x_6579 = x_2917 & x_2918;
assign x_6580 = x_6578 & x_6579;
assign x_6581 = x_2919 & x_2920;
assign x_6582 = x_2921 & x_2922;
assign x_6583 = x_6581 & x_6582;
assign x_6584 = x_6580 & x_6583;
assign x_6585 = x_6577 & x_6584;
assign x_6586 = x_6571 & x_6585;
assign x_6587 = x_6558 & x_6586;
assign x_6588 = x_2924 & x_2925;
assign x_6589 = x_2923 & x_6588;
assign x_6590 = x_2926 & x_2927;
assign x_6591 = x_2928 & x_2929;
assign x_6592 = x_6590 & x_6591;
assign x_6593 = x_6589 & x_6592;
assign x_6594 = x_2931 & x_2932;
assign x_6595 = x_2930 & x_6594;
assign x_6596 = x_2933 & x_2934;
assign x_6597 = x_2935 & x_2936;
assign x_6598 = x_6596 & x_6597;
assign x_6599 = x_6595 & x_6598;
assign x_6600 = x_6593 & x_6599;
assign x_6601 = x_2938 & x_2939;
assign x_6602 = x_2937 & x_6601;
assign x_6603 = x_2940 & x_2941;
assign x_6604 = x_2942 & x_2943;
assign x_6605 = x_6603 & x_6604;
assign x_6606 = x_6602 & x_6605;
assign x_6607 = x_2944 & x_2945;
assign x_6608 = x_2946 & x_2947;
assign x_6609 = x_6607 & x_6608;
assign x_6610 = x_2948 & x_2949;
assign x_6611 = x_2950 & x_2951;
assign x_6612 = x_6610 & x_6611;
assign x_6613 = x_6609 & x_6612;
assign x_6614 = x_6606 & x_6613;
assign x_6615 = x_6600 & x_6614;
assign x_6616 = x_2953 & x_2954;
assign x_6617 = x_2952 & x_6616;
assign x_6618 = x_2955 & x_2956;
assign x_6619 = x_2957 & x_2958;
assign x_6620 = x_6618 & x_6619;
assign x_6621 = x_6617 & x_6620;
assign x_6622 = x_2960 & x_2961;
assign x_6623 = x_2959 & x_6622;
assign x_6624 = x_2962 & x_2963;
assign x_6625 = x_2964 & x_2965;
assign x_6626 = x_6624 & x_6625;
assign x_6627 = x_6623 & x_6626;
assign x_6628 = x_6621 & x_6627;
assign x_6629 = x_2967 & x_2968;
assign x_6630 = x_2966 & x_6629;
assign x_6631 = x_2969 & x_2970;
assign x_6632 = x_2971 & x_2972;
assign x_6633 = x_6631 & x_6632;
assign x_6634 = x_6630 & x_6633;
assign x_6635 = x_2973 & x_2974;
assign x_6636 = x_2975 & x_2976;
assign x_6637 = x_6635 & x_6636;
assign x_6638 = x_2977 & x_2978;
assign x_6639 = x_2979 & x_2980;
assign x_6640 = x_6638 & x_6639;
assign x_6641 = x_6637 & x_6640;
assign x_6642 = x_6634 & x_6641;
assign x_6643 = x_6628 & x_6642;
assign x_6644 = x_6615 & x_6643;
assign x_6645 = x_6587 & x_6644;
assign x_6646 = x_6531 & x_6645;
assign x_6647 = x_2982 & x_2983;
assign x_6648 = x_2981 & x_6647;
assign x_6649 = x_2984 & x_2985;
assign x_6650 = x_2986 & x_2987;
assign x_6651 = x_6649 & x_6650;
assign x_6652 = x_6648 & x_6651;
assign x_6653 = x_2989 & x_2990;
assign x_6654 = x_2988 & x_6653;
assign x_6655 = x_2991 & x_2992;
assign x_6656 = x_2993 & x_2994;
assign x_6657 = x_6655 & x_6656;
assign x_6658 = x_6654 & x_6657;
assign x_6659 = x_6652 & x_6658;
assign x_6660 = x_2996 & x_2997;
assign x_6661 = x_2995 & x_6660;
assign x_6662 = x_2998 & x_2999;
assign x_6663 = x_3000 & x_3001;
assign x_6664 = x_6662 & x_6663;
assign x_6665 = x_6661 & x_6664;
assign x_6666 = x_3003 & x_3004;
assign x_6667 = x_3002 & x_6666;
assign x_6668 = x_3005 & x_3006;
assign x_6669 = x_3007 & x_3008;
assign x_6670 = x_6668 & x_6669;
assign x_6671 = x_6667 & x_6670;
assign x_6672 = x_6665 & x_6671;
assign x_6673 = x_6659 & x_6672;
assign x_6674 = x_3010 & x_3011;
assign x_6675 = x_3009 & x_6674;
assign x_6676 = x_3012 & x_3013;
assign x_6677 = x_3014 & x_3015;
assign x_6678 = x_6676 & x_6677;
assign x_6679 = x_6675 & x_6678;
assign x_6680 = x_3017 & x_3018;
assign x_6681 = x_3016 & x_6680;
assign x_6682 = x_3019 & x_3020;
assign x_6683 = x_3021 & x_3022;
assign x_6684 = x_6682 & x_6683;
assign x_6685 = x_6681 & x_6684;
assign x_6686 = x_6679 & x_6685;
assign x_6687 = x_3024 & x_3025;
assign x_6688 = x_3023 & x_6687;
assign x_6689 = x_3026 & x_3027;
assign x_6690 = x_3028 & x_3029;
assign x_6691 = x_6689 & x_6690;
assign x_6692 = x_6688 & x_6691;
assign x_6693 = x_3030 & x_3031;
assign x_6694 = x_3032 & x_3033;
assign x_6695 = x_6693 & x_6694;
assign x_6696 = x_3034 & x_3035;
assign x_6697 = x_3036 & x_3037;
assign x_6698 = x_6696 & x_6697;
assign x_6699 = x_6695 & x_6698;
assign x_6700 = x_6692 & x_6699;
assign x_6701 = x_6686 & x_6700;
assign x_6702 = x_6673 & x_6701;
assign x_6703 = x_3039 & x_3040;
assign x_6704 = x_3038 & x_6703;
assign x_6705 = x_3041 & x_3042;
assign x_6706 = x_3043 & x_3044;
assign x_6707 = x_6705 & x_6706;
assign x_6708 = x_6704 & x_6707;
assign x_6709 = x_3046 & x_3047;
assign x_6710 = x_3045 & x_6709;
assign x_6711 = x_3048 & x_3049;
assign x_6712 = x_3050 & x_3051;
assign x_6713 = x_6711 & x_6712;
assign x_6714 = x_6710 & x_6713;
assign x_6715 = x_6708 & x_6714;
assign x_6716 = x_3053 & x_3054;
assign x_6717 = x_3052 & x_6716;
assign x_6718 = x_3055 & x_3056;
assign x_6719 = x_3057 & x_3058;
assign x_6720 = x_6718 & x_6719;
assign x_6721 = x_6717 & x_6720;
assign x_6722 = x_3059 & x_3060;
assign x_6723 = x_3061 & x_3062;
assign x_6724 = x_6722 & x_6723;
assign x_6725 = x_3063 & x_3064;
assign x_6726 = x_3065 & x_3066;
assign x_6727 = x_6725 & x_6726;
assign x_6728 = x_6724 & x_6727;
assign x_6729 = x_6721 & x_6728;
assign x_6730 = x_6715 & x_6729;
assign x_6731 = x_3068 & x_3069;
assign x_6732 = x_3067 & x_6731;
assign x_6733 = x_3070 & x_3071;
assign x_6734 = x_3072 & x_3073;
assign x_6735 = x_6733 & x_6734;
assign x_6736 = x_6732 & x_6735;
assign x_6737 = x_3075 & x_3076;
assign x_6738 = x_3074 & x_6737;
assign x_6739 = x_3077 & x_3078;
assign x_6740 = x_3079 & x_3080;
assign x_6741 = x_6739 & x_6740;
assign x_6742 = x_6738 & x_6741;
assign x_6743 = x_6736 & x_6742;
assign x_6744 = x_3082 & x_3083;
assign x_6745 = x_3081 & x_6744;
assign x_6746 = x_3084 & x_3085;
assign x_6747 = x_3086 & x_3087;
assign x_6748 = x_6746 & x_6747;
assign x_6749 = x_6745 & x_6748;
assign x_6750 = x_3088 & x_3089;
assign x_6751 = x_3090 & x_3091;
assign x_6752 = x_6750 & x_6751;
assign x_6753 = x_3092 & x_3093;
assign x_6754 = x_3094 & x_3095;
assign x_6755 = x_6753 & x_6754;
assign x_6756 = x_6752 & x_6755;
assign x_6757 = x_6749 & x_6756;
assign x_6758 = x_6743 & x_6757;
assign x_6759 = x_6730 & x_6758;
assign x_6760 = x_6702 & x_6759;
assign x_6761 = x_3097 & x_3098;
assign x_6762 = x_3096 & x_6761;
assign x_6763 = x_3099 & x_3100;
assign x_6764 = x_3101 & x_3102;
assign x_6765 = x_6763 & x_6764;
assign x_6766 = x_6762 & x_6765;
assign x_6767 = x_3104 & x_3105;
assign x_6768 = x_3103 & x_6767;
assign x_6769 = x_3106 & x_3107;
assign x_6770 = x_3108 & x_3109;
assign x_6771 = x_6769 & x_6770;
assign x_6772 = x_6768 & x_6771;
assign x_6773 = x_6766 & x_6772;
assign x_6774 = x_3111 & x_3112;
assign x_6775 = x_3110 & x_6774;
assign x_6776 = x_3113 & x_3114;
assign x_6777 = x_3115 & x_3116;
assign x_6778 = x_6776 & x_6777;
assign x_6779 = x_6775 & x_6778;
assign x_6780 = x_3118 & x_3119;
assign x_6781 = x_3117 & x_6780;
assign x_6782 = x_3120 & x_3121;
assign x_6783 = x_3122 & x_3123;
assign x_6784 = x_6782 & x_6783;
assign x_6785 = x_6781 & x_6784;
assign x_6786 = x_6779 & x_6785;
assign x_6787 = x_6773 & x_6786;
assign x_6788 = x_3125 & x_3126;
assign x_6789 = x_3124 & x_6788;
assign x_6790 = x_3127 & x_3128;
assign x_6791 = x_3129 & x_3130;
assign x_6792 = x_6790 & x_6791;
assign x_6793 = x_6789 & x_6792;
assign x_6794 = x_3132 & x_3133;
assign x_6795 = x_3131 & x_6794;
assign x_6796 = x_3134 & x_3135;
assign x_6797 = x_3136 & x_3137;
assign x_6798 = x_6796 & x_6797;
assign x_6799 = x_6795 & x_6798;
assign x_6800 = x_6793 & x_6799;
assign x_6801 = x_3139 & x_3140;
assign x_6802 = x_3138 & x_6801;
assign x_6803 = x_3141 & x_3142;
assign x_6804 = x_3143 & x_3144;
assign x_6805 = x_6803 & x_6804;
assign x_6806 = x_6802 & x_6805;
assign x_6807 = x_3145 & x_3146;
assign x_6808 = x_3147 & x_3148;
assign x_6809 = x_6807 & x_6808;
assign x_6810 = x_3149 & x_3150;
assign x_6811 = x_3151 & x_3152;
assign x_6812 = x_6810 & x_6811;
assign x_6813 = x_6809 & x_6812;
assign x_6814 = x_6806 & x_6813;
assign x_6815 = x_6800 & x_6814;
assign x_6816 = x_6787 & x_6815;
assign x_6817 = x_3154 & x_3155;
assign x_6818 = x_3153 & x_6817;
assign x_6819 = x_3156 & x_3157;
assign x_6820 = x_3158 & x_3159;
assign x_6821 = x_6819 & x_6820;
assign x_6822 = x_6818 & x_6821;
assign x_6823 = x_3161 & x_3162;
assign x_6824 = x_3160 & x_6823;
assign x_6825 = x_3163 & x_3164;
assign x_6826 = x_3165 & x_3166;
assign x_6827 = x_6825 & x_6826;
assign x_6828 = x_6824 & x_6827;
assign x_6829 = x_6822 & x_6828;
assign x_6830 = x_3168 & x_3169;
assign x_6831 = x_3167 & x_6830;
assign x_6832 = x_3170 & x_3171;
assign x_6833 = x_3172 & x_3173;
assign x_6834 = x_6832 & x_6833;
assign x_6835 = x_6831 & x_6834;
assign x_6836 = x_3174 & x_3175;
assign x_6837 = x_3176 & x_3177;
assign x_6838 = x_6836 & x_6837;
assign x_6839 = x_3178 & x_3179;
assign x_6840 = x_3180 & x_3181;
assign x_6841 = x_6839 & x_6840;
assign x_6842 = x_6838 & x_6841;
assign x_6843 = x_6835 & x_6842;
assign x_6844 = x_6829 & x_6843;
assign x_6845 = x_3183 & x_3184;
assign x_6846 = x_3182 & x_6845;
assign x_6847 = x_3185 & x_3186;
assign x_6848 = x_3187 & x_3188;
assign x_6849 = x_6847 & x_6848;
assign x_6850 = x_6846 & x_6849;
assign x_6851 = x_3190 & x_3191;
assign x_6852 = x_3189 & x_6851;
assign x_6853 = x_3192 & x_3193;
assign x_6854 = x_3194 & x_3195;
assign x_6855 = x_6853 & x_6854;
assign x_6856 = x_6852 & x_6855;
assign x_6857 = x_6850 & x_6856;
assign x_6858 = x_3197 & x_3198;
assign x_6859 = x_3196 & x_6858;
assign x_6860 = x_3199 & x_3200;
assign x_6861 = x_3201 & x_3202;
assign x_6862 = x_6860 & x_6861;
assign x_6863 = x_6859 & x_6862;
assign x_6864 = x_3203 & x_3204;
assign x_6865 = x_3205 & x_3206;
assign x_6866 = x_6864 & x_6865;
assign x_6867 = x_3207 & x_3208;
assign x_6868 = x_3209 & x_3210;
assign x_6869 = x_6867 & x_6868;
assign x_6870 = x_6866 & x_6869;
assign x_6871 = x_6863 & x_6870;
assign x_6872 = x_6857 & x_6871;
assign x_6873 = x_6844 & x_6872;
assign x_6874 = x_6816 & x_6873;
assign x_6875 = x_6760 & x_6874;
assign x_6876 = x_6646 & x_6875;
assign x_6877 = x_3212 & x_3213;
assign x_6878 = x_3211 & x_6877;
assign x_6879 = x_3214 & x_3215;
assign x_6880 = x_3216 & x_3217;
assign x_6881 = x_6879 & x_6880;
assign x_6882 = x_6878 & x_6881;
assign x_6883 = x_3219 & x_3220;
assign x_6884 = x_3218 & x_6883;
assign x_6885 = x_3221 & x_3222;
assign x_6886 = x_3223 & x_3224;
assign x_6887 = x_6885 & x_6886;
assign x_6888 = x_6884 & x_6887;
assign x_6889 = x_6882 & x_6888;
assign x_6890 = x_3226 & x_3227;
assign x_6891 = x_3225 & x_6890;
assign x_6892 = x_3228 & x_3229;
assign x_6893 = x_3230 & x_3231;
assign x_6894 = x_6892 & x_6893;
assign x_6895 = x_6891 & x_6894;
assign x_6896 = x_3233 & x_3234;
assign x_6897 = x_3232 & x_6896;
assign x_6898 = x_3235 & x_3236;
assign x_6899 = x_3237 & x_3238;
assign x_6900 = x_6898 & x_6899;
assign x_6901 = x_6897 & x_6900;
assign x_6902 = x_6895 & x_6901;
assign x_6903 = x_6889 & x_6902;
assign x_6904 = x_3240 & x_3241;
assign x_6905 = x_3239 & x_6904;
assign x_6906 = x_3242 & x_3243;
assign x_6907 = x_3244 & x_3245;
assign x_6908 = x_6906 & x_6907;
assign x_6909 = x_6905 & x_6908;
assign x_6910 = x_3247 & x_3248;
assign x_6911 = x_3246 & x_6910;
assign x_6912 = x_3249 & x_3250;
assign x_6913 = x_3251 & x_3252;
assign x_6914 = x_6912 & x_6913;
assign x_6915 = x_6911 & x_6914;
assign x_6916 = x_6909 & x_6915;
assign x_6917 = x_3254 & x_3255;
assign x_6918 = x_3253 & x_6917;
assign x_6919 = x_3256 & x_3257;
assign x_6920 = x_3258 & x_3259;
assign x_6921 = x_6919 & x_6920;
assign x_6922 = x_6918 & x_6921;
assign x_6923 = x_3260 & x_3261;
assign x_6924 = x_3262 & x_3263;
assign x_6925 = x_6923 & x_6924;
assign x_6926 = x_3264 & x_3265;
assign x_6927 = x_3266 & x_3267;
assign x_6928 = x_6926 & x_6927;
assign x_6929 = x_6925 & x_6928;
assign x_6930 = x_6922 & x_6929;
assign x_6931 = x_6916 & x_6930;
assign x_6932 = x_6903 & x_6931;
assign x_6933 = x_3269 & x_3270;
assign x_6934 = x_3268 & x_6933;
assign x_6935 = x_3271 & x_3272;
assign x_6936 = x_3273 & x_3274;
assign x_6937 = x_6935 & x_6936;
assign x_6938 = x_6934 & x_6937;
assign x_6939 = x_3276 & x_3277;
assign x_6940 = x_3275 & x_6939;
assign x_6941 = x_3278 & x_3279;
assign x_6942 = x_3280 & x_3281;
assign x_6943 = x_6941 & x_6942;
assign x_6944 = x_6940 & x_6943;
assign x_6945 = x_6938 & x_6944;
assign x_6946 = x_3283 & x_3284;
assign x_6947 = x_3282 & x_6946;
assign x_6948 = x_3285 & x_3286;
assign x_6949 = x_3287 & x_3288;
assign x_6950 = x_6948 & x_6949;
assign x_6951 = x_6947 & x_6950;
assign x_6952 = x_3290 & x_3291;
assign x_6953 = x_3289 & x_6952;
assign x_6954 = x_3292 & x_3293;
assign x_6955 = x_3294 & x_3295;
assign x_6956 = x_6954 & x_6955;
assign x_6957 = x_6953 & x_6956;
assign x_6958 = x_6951 & x_6957;
assign x_6959 = x_6945 & x_6958;
assign x_6960 = x_3297 & x_3298;
assign x_6961 = x_3296 & x_6960;
assign x_6962 = x_3299 & x_3300;
assign x_6963 = x_3301 & x_3302;
assign x_6964 = x_6962 & x_6963;
assign x_6965 = x_6961 & x_6964;
assign x_6966 = x_3304 & x_3305;
assign x_6967 = x_3303 & x_6966;
assign x_6968 = x_3306 & x_3307;
assign x_6969 = x_3308 & x_3309;
assign x_6970 = x_6968 & x_6969;
assign x_6971 = x_6967 & x_6970;
assign x_6972 = x_6965 & x_6971;
assign x_6973 = x_3311 & x_3312;
assign x_6974 = x_3310 & x_6973;
assign x_6975 = x_3313 & x_3314;
assign x_6976 = x_3315 & x_3316;
assign x_6977 = x_6975 & x_6976;
assign x_6978 = x_6974 & x_6977;
assign x_6979 = x_3317 & x_3318;
assign x_6980 = x_3319 & x_3320;
assign x_6981 = x_6979 & x_6980;
assign x_6982 = x_3321 & x_3322;
assign x_6983 = x_3323 & x_3324;
assign x_6984 = x_6982 & x_6983;
assign x_6985 = x_6981 & x_6984;
assign x_6986 = x_6978 & x_6985;
assign x_6987 = x_6972 & x_6986;
assign x_6988 = x_6959 & x_6987;
assign x_6989 = x_6932 & x_6988;
assign x_6990 = x_3326 & x_3327;
assign x_6991 = x_3325 & x_6990;
assign x_6992 = x_3328 & x_3329;
assign x_6993 = x_3330 & x_3331;
assign x_6994 = x_6992 & x_6993;
assign x_6995 = x_6991 & x_6994;
assign x_6996 = x_3333 & x_3334;
assign x_6997 = x_3332 & x_6996;
assign x_6998 = x_3335 & x_3336;
assign x_6999 = x_3337 & x_3338;
assign x_7000 = x_6998 & x_6999;
assign x_7001 = x_6997 & x_7000;
assign x_7002 = x_6995 & x_7001;
assign x_7003 = x_3340 & x_3341;
assign x_7004 = x_3339 & x_7003;
assign x_7005 = x_3342 & x_3343;
assign x_7006 = x_3344 & x_3345;
assign x_7007 = x_7005 & x_7006;
assign x_7008 = x_7004 & x_7007;
assign x_7009 = x_3347 & x_3348;
assign x_7010 = x_3346 & x_7009;
assign x_7011 = x_3349 & x_3350;
assign x_7012 = x_3351 & x_3352;
assign x_7013 = x_7011 & x_7012;
assign x_7014 = x_7010 & x_7013;
assign x_7015 = x_7008 & x_7014;
assign x_7016 = x_7002 & x_7015;
assign x_7017 = x_3354 & x_3355;
assign x_7018 = x_3353 & x_7017;
assign x_7019 = x_3356 & x_3357;
assign x_7020 = x_3358 & x_3359;
assign x_7021 = x_7019 & x_7020;
assign x_7022 = x_7018 & x_7021;
assign x_7023 = x_3361 & x_3362;
assign x_7024 = x_3360 & x_7023;
assign x_7025 = x_3363 & x_3364;
assign x_7026 = x_3365 & x_3366;
assign x_7027 = x_7025 & x_7026;
assign x_7028 = x_7024 & x_7027;
assign x_7029 = x_7022 & x_7028;
assign x_7030 = x_3368 & x_3369;
assign x_7031 = x_3367 & x_7030;
assign x_7032 = x_3370 & x_3371;
assign x_7033 = x_3372 & x_3373;
assign x_7034 = x_7032 & x_7033;
assign x_7035 = x_7031 & x_7034;
assign x_7036 = x_3374 & x_3375;
assign x_7037 = x_3376 & x_3377;
assign x_7038 = x_7036 & x_7037;
assign x_7039 = x_3378 & x_3379;
assign x_7040 = x_3380 & x_3381;
assign x_7041 = x_7039 & x_7040;
assign x_7042 = x_7038 & x_7041;
assign x_7043 = x_7035 & x_7042;
assign x_7044 = x_7029 & x_7043;
assign x_7045 = x_7016 & x_7044;
assign x_7046 = x_3383 & x_3384;
assign x_7047 = x_3382 & x_7046;
assign x_7048 = x_3385 & x_3386;
assign x_7049 = x_3387 & x_3388;
assign x_7050 = x_7048 & x_7049;
assign x_7051 = x_7047 & x_7050;
assign x_7052 = x_3390 & x_3391;
assign x_7053 = x_3389 & x_7052;
assign x_7054 = x_3392 & x_3393;
assign x_7055 = x_3394 & x_3395;
assign x_7056 = x_7054 & x_7055;
assign x_7057 = x_7053 & x_7056;
assign x_7058 = x_7051 & x_7057;
assign x_7059 = x_3397 & x_3398;
assign x_7060 = x_3396 & x_7059;
assign x_7061 = x_3399 & x_3400;
assign x_7062 = x_3401 & x_3402;
assign x_7063 = x_7061 & x_7062;
assign x_7064 = x_7060 & x_7063;
assign x_7065 = x_3403 & x_3404;
assign x_7066 = x_3405 & x_3406;
assign x_7067 = x_7065 & x_7066;
assign x_7068 = x_3407 & x_3408;
assign x_7069 = x_3409 & x_3410;
assign x_7070 = x_7068 & x_7069;
assign x_7071 = x_7067 & x_7070;
assign x_7072 = x_7064 & x_7071;
assign x_7073 = x_7058 & x_7072;
assign x_7074 = x_3412 & x_3413;
assign x_7075 = x_3411 & x_7074;
assign x_7076 = x_3414 & x_3415;
assign x_7077 = x_3416 & x_3417;
assign x_7078 = x_7076 & x_7077;
assign x_7079 = x_7075 & x_7078;
assign x_7080 = x_3419 & x_3420;
assign x_7081 = x_3418 & x_7080;
assign x_7082 = x_3421 & x_3422;
assign x_7083 = x_3423 & x_3424;
assign x_7084 = x_7082 & x_7083;
assign x_7085 = x_7081 & x_7084;
assign x_7086 = x_7079 & x_7085;
assign x_7087 = x_3426 & x_3427;
assign x_7088 = x_3425 & x_7087;
assign x_7089 = x_3428 & x_3429;
assign x_7090 = x_3430 & x_3431;
assign x_7091 = x_7089 & x_7090;
assign x_7092 = x_7088 & x_7091;
assign x_7093 = x_3432 & x_3433;
assign x_7094 = x_3434 & x_3435;
assign x_7095 = x_7093 & x_7094;
assign x_7096 = x_3436 & x_3437;
assign x_7097 = x_3438 & x_3439;
assign x_7098 = x_7096 & x_7097;
assign x_7099 = x_7095 & x_7098;
assign x_7100 = x_7092 & x_7099;
assign x_7101 = x_7086 & x_7100;
assign x_7102 = x_7073 & x_7101;
assign x_7103 = x_7045 & x_7102;
assign x_7104 = x_6989 & x_7103;
assign x_7105 = x_3441 & x_3442;
assign x_7106 = x_3440 & x_7105;
assign x_7107 = x_3443 & x_3444;
assign x_7108 = x_3445 & x_3446;
assign x_7109 = x_7107 & x_7108;
assign x_7110 = x_7106 & x_7109;
assign x_7111 = x_3448 & x_3449;
assign x_7112 = x_3447 & x_7111;
assign x_7113 = x_3450 & x_3451;
assign x_7114 = x_3452 & x_3453;
assign x_7115 = x_7113 & x_7114;
assign x_7116 = x_7112 & x_7115;
assign x_7117 = x_7110 & x_7116;
assign x_7118 = x_3455 & x_3456;
assign x_7119 = x_3454 & x_7118;
assign x_7120 = x_3457 & x_3458;
assign x_7121 = x_3459 & x_3460;
assign x_7122 = x_7120 & x_7121;
assign x_7123 = x_7119 & x_7122;
assign x_7124 = x_3462 & x_3463;
assign x_7125 = x_3461 & x_7124;
assign x_7126 = x_3464 & x_3465;
assign x_7127 = x_3466 & x_3467;
assign x_7128 = x_7126 & x_7127;
assign x_7129 = x_7125 & x_7128;
assign x_7130 = x_7123 & x_7129;
assign x_7131 = x_7117 & x_7130;
assign x_7132 = x_3469 & x_3470;
assign x_7133 = x_3468 & x_7132;
assign x_7134 = x_3471 & x_3472;
assign x_7135 = x_3473 & x_3474;
assign x_7136 = x_7134 & x_7135;
assign x_7137 = x_7133 & x_7136;
assign x_7138 = x_3476 & x_3477;
assign x_7139 = x_3475 & x_7138;
assign x_7140 = x_3478 & x_3479;
assign x_7141 = x_3480 & x_3481;
assign x_7142 = x_7140 & x_7141;
assign x_7143 = x_7139 & x_7142;
assign x_7144 = x_7137 & x_7143;
assign x_7145 = x_3483 & x_3484;
assign x_7146 = x_3482 & x_7145;
assign x_7147 = x_3485 & x_3486;
assign x_7148 = x_3487 & x_3488;
assign x_7149 = x_7147 & x_7148;
assign x_7150 = x_7146 & x_7149;
assign x_7151 = x_3489 & x_3490;
assign x_7152 = x_3491 & x_3492;
assign x_7153 = x_7151 & x_7152;
assign x_7154 = x_3493 & x_3494;
assign x_7155 = x_3495 & x_3496;
assign x_7156 = x_7154 & x_7155;
assign x_7157 = x_7153 & x_7156;
assign x_7158 = x_7150 & x_7157;
assign x_7159 = x_7144 & x_7158;
assign x_7160 = x_7131 & x_7159;
assign x_7161 = x_3498 & x_3499;
assign x_7162 = x_3497 & x_7161;
assign x_7163 = x_3500 & x_3501;
assign x_7164 = x_3502 & x_3503;
assign x_7165 = x_7163 & x_7164;
assign x_7166 = x_7162 & x_7165;
assign x_7167 = x_3505 & x_3506;
assign x_7168 = x_3504 & x_7167;
assign x_7169 = x_3507 & x_3508;
assign x_7170 = x_3509 & x_3510;
assign x_7171 = x_7169 & x_7170;
assign x_7172 = x_7168 & x_7171;
assign x_7173 = x_7166 & x_7172;
assign x_7174 = x_3512 & x_3513;
assign x_7175 = x_3511 & x_7174;
assign x_7176 = x_3514 & x_3515;
assign x_7177 = x_3516 & x_3517;
assign x_7178 = x_7176 & x_7177;
assign x_7179 = x_7175 & x_7178;
assign x_7180 = x_3518 & x_3519;
assign x_7181 = x_3520 & x_3521;
assign x_7182 = x_7180 & x_7181;
assign x_7183 = x_3522 & x_3523;
assign x_7184 = x_3524 & x_3525;
assign x_7185 = x_7183 & x_7184;
assign x_7186 = x_7182 & x_7185;
assign x_7187 = x_7179 & x_7186;
assign x_7188 = x_7173 & x_7187;
assign x_7189 = x_3527 & x_3528;
assign x_7190 = x_3526 & x_7189;
assign x_7191 = x_3529 & x_3530;
assign x_7192 = x_3531 & x_3532;
assign x_7193 = x_7191 & x_7192;
assign x_7194 = x_7190 & x_7193;
assign x_7195 = x_3534 & x_3535;
assign x_7196 = x_3533 & x_7195;
assign x_7197 = x_3536 & x_3537;
assign x_7198 = x_3538 & x_3539;
assign x_7199 = x_7197 & x_7198;
assign x_7200 = x_7196 & x_7199;
assign x_7201 = x_7194 & x_7200;
assign x_7202 = x_3541 & x_3542;
assign x_7203 = x_3540 & x_7202;
assign x_7204 = x_3543 & x_3544;
assign x_7205 = x_3545 & x_3546;
assign x_7206 = x_7204 & x_7205;
assign x_7207 = x_7203 & x_7206;
assign x_7208 = x_3547 & x_3548;
assign x_7209 = x_3549 & x_3550;
assign x_7210 = x_7208 & x_7209;
assign x_7211 = x_3551 & x_3552;
assign x_7212 = x_3553 & x_3554;
assign x_7213 = x_7211 & x_7212;
assign x_7214 = x_7210 & x_7213;
assign x_7215 = x_7207 & x_7214;
assign x_7216 = x_7201 & x_7215;
assign x_7217 = x_7188 & x_7216;
assign x_7218 = x_7160 & x_7217;
assign x_7219 = x_3556 & x_3557;
assign x_7220 = x_3555 & x_7219;
assign x_7221 = x_3558 & x_3559;
assign x_7222 = x_3560 & x_3561;
assign x_7223 = x_7221 & x_7222;
assign x_7224 = x_7220 & x_7223;
assign x_7225 = x_3563 & x_3564;
assign x_7226 = x_3562 & x_7225;
assign x_7227 = x_3565 & x_3566;
assign x_7228 = x_3567 & x_3568;
assign x_7229 = x_7227 & x_7228;
assign x_7230 = x_7226 & x_7229;
assign x_7231 = x_7224 & x_7230;
assign x_7232 = x_3570 & x_3571;
assign x_7233 = x_3569 & x_7232;
assign x_7234 = x_3572 & x_3573;
assign x_7235 = x_3574 & x_3575;
assign x_7236 = x_7234 & x_7235;
assign x_7237 = x_7233 & x_7236;
assign x_7238 = x_3577 & x_3578;
assign x_7239 = x_3576 & x_7238;
assign x_7240 = x_3579 & x_3580;
assign x_7241 = x_3581 & x_3582;
assign x_7242 = x_7240 & x_7241;
assign x_7243 = x_7239 & x_7242;
assign x_7244 = x_7237 & x_7243;
assign x_7245 = x_7231 & x_7244;
assign x_7246 = x_3584 & x_3585;
assign x_7247 = x_3583 & x_7246;
assign x_7248 = x_3586 & x_3587;
assign x_7249 = x_3588 & x_3589;
assign x_7250 = x_7248 & x_7249;
assign x_7251 = x_7247 & x_7250;
assign x_7252 = x_3591 & x_3592;
assign x_7253 = x_3590 & x_7252;
assign x_7254 = x_3593 & x_3594;
assign x_7255 = x_3595 & x_3596;
assign x_7256 = x_7254 & x_7255;
assign x_7257 = x_7253 & x_7256;
assign x_7258 = x_7251 & x_7257;
assign x_7259 = x_3598 & x_3599;
assign x_7260 = x_3597 & x_7259;
assign x_7261 = x_3600 & x_3601;
assign x_7262 = x_3602 & x_3603;
assign x_7263 = x_7261 & x_7262;
assign x_7264 = x_7260 & x_7263;
assign x_7265 = x_3604 & x_3605;
assign x_7266 = x_3606 & x_3607;
assign x_7267 = x_7265 & x_7266;
assign x_7268 = x_3608 & x_3609;
assign x_7269 = x_3610 & x_3611;
assign x_7270 = x_7268 & x_7269;
assign x_7271 = x_7267 & x_7270;
assign x_7272 = x_7264 & x_7271;
assign x_7273 = x_7258 & x_7272;
assign x_7274 = x_7245 & x_7273;
assign x_7275 = x_3613 & x_3614;
assign x_7276 = x_3612 & x_7275;
assign x_7277 = x_3615 & x_3616;
assign x_7278 = x_3617 & x_3618;
assign x_7279 = x_7277 & x_7278;
assign x_7280 = x_7276 & x_7279;
assign x_7281 = x_3620 & x_3621;
assign x_7282 = x_3619 & x_7281;
assign x_7283 = x_3622 & x_3623;
assign x_7284 = x_3624 & x_3625;
assign x_7285 = x_7283 & x_7284;
assign x_7286 = x_7282 & x_7285;
assign x_7287 = x_7280 & x_7286;
assign x_7288 = x_3627 & x_3628;
assign x_7289 = x_3626 & x_7288;
assign x_7290 = x_3629 & x_3630;
assign x_7291 = x_3631 & x_3632;
assign x_7292 = x_7290 & x_7291;
assign x_7293 = x_7289 & x_7292;
assign x_7294 = x_3633 & x_3634;
assign x_7295 = x_3635 & x_3636;
assign x_7296 = x_7294 & x_7295;
assign x_7297 = x_3637 & x_3638;
assign x_7298 = x_3639 & x_3640;
assign x_7299 = x_7297 & x_7298;
assign x_7300 = x_7296 & x_7299;
assign x_7301 = x_7293 & x_7300;
assign x_7302 = x_7287 & x_7301;
assign x_7303 = x_3642 & x_3643;
assign x_7304 = x_3641 & x_7303;
assign x_7305 = x_3644 & x_3645;
assign x_7306 = x_3646 & x_3647;
assign x_7307 = x_7305 & x_7306;
assign x_7308 = x_7304 & x_7307;
assign x_7309 = x_3649 & x_3650;
assign x_7310 = x_3648 & x_7309;
assign x_7311 = x_3651 & x_3652;
assign x_7312 = x_3653 & x_3654;
assign x_7313 = x_7311 & x_7312;
assign x_7314 = x_7310 & x_7313;
assign x_7315 = x_7308 & x_7314;
assign x_7316 = x_3656 & x_3657;
assign x_7317 = x_3655 & x_7316;
assign x_7318 = x_3658 & x_3659;
assign x_7319 = x_3660 & x_3661;
assign x_7320 = x_7318 & x_7319;
assign x_7321 = x_7317 & x_7320;
assign x_7322 = x_3662 & x_3663;
assign x_7323 = x_3664 & x_3665;
assign x_7324 = x_7322 & x_7323;
assign x_7325 = x_3666 & x_3667;
assign x_7326 = x_3668 & x_3669;
assign x_7327 = x_7325 & x_7326;
assign x_7328 = x_7324 & x_7327;
assign x_7329 = x_7321 & x_7328;
assign x_7330 = x_7315 & x_7329;
assign x_7331 = x_7302 & x_7330;
assign x_7332 = x_7274 & x_7331;
assign x_7333 = x_7218 & x_7332;
assign x_7334 = x_7104 & x_7333;
assign x_7335 = x_6876 & x_7334;
assign x_7336 = x_6418 & x_7335;
assign x_7337 = x_5502 & x_7336;
assign o_1 = x_7337;
endmodule
