// Benchmark "SKOLEMFORMULA" written by ABC on Sun May 22 05:53:57 2022

module SKOLEMFORMULA ( 
    i0,
    i1, i2, i3, i4  );
  input  i0;
  output i1, i2, i3, i4;
  assign i1 = 1'b0;
  assign i2 = 1'b1;
  assign i3 = 1'b1;
  assign i4 = ~i0;
endmodule


