module formula(i_12,i_33,out);
	input i_12 ,i_33;

	output out;
	assign out = i_12;
endmodule
