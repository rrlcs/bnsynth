// skolem function for order file variables
// Generated using findDep.cpp 
module kenflashp12 (v_338, v_339, v_340, v_341, v_342, v_343, v_344, v_345, v_346, v_347, v_348, v_349, v_350, v_351, v_352, v_353, v_354, v_355, v_356, v_357, v_358, v_359, v_360, v_361, v_362, v_363, v_364, v_365, v_366, v_367, v_368, v_369, v_370, v_371, v_372, v_373, v_374, v_375, v_376, v_377, v_378, v_379, v_380, v_381, v_296, v_297, v_298, v_299, v_300, v_301, v_302, v_303, v_304, v_305, v_306, v_307, v_308, v_309, v_310, v_311, v_312, v_313, v_314, v_315, v_316, v_317, v_318, v_319, v_320, v_321, v_322, v_323, v_324, v_325, v_326, v_327, v_328, v_329, v_330, v_331, v_332, v_333, v_334, v_335, v_336, v_337, v_5, v_7, v_8, v_10, v_12, v_15, v_16, v_18, v_24, v_26, v_27, v_30, v_31, v_40, v_42, v_45, v_51, v_53, v_55, v_57, v_59, v_63, v_66, v_67, v_70, v_71, v_72, v_74, v_77, v_78, v_79, v_81, v_82, v_87, v_88, v_89, v_94, v_95, v_97, v_99, v_100, v_101, v_102, v_105, v_106, v_107, v_108, v_109, v_112, v_114, v_116, v_119, v_121, v_122, v_123, v_124, v_126, v_128, v_130, v_131, v_132, v_133, v_136, v_138, v_139, v_140, v_141, v_143, v_145, v_146, v_147, v_148, v_151, v_154, v_155, v_157, v_159, v_161, v_163, v_166, v_167, v_169, v_172, v_173, v_175, v_176, v_177, v_178, v_179, v_180, v_182, v_183, v_184, v_185, v_186, v_187, v_189, v_190, v_191, v_192, v_193, v_194, v_195, v_196, v_197, v_198, v_200, v_201, v_203, v_205, v_206, v_209, v_211, v_212, v_214, v_216, v_217, v_218, v_220, v_221, v_222, v_224, v_226, v_227, v_228, v_230, v_231, v_233, v_234, v_236, v_237, v_238, v_239, v_240, v_242, v_243, v_245, v_246, v_247, v_250, v_251, v_255, v_256, v_259, v_260, v_261, v_267, v_269, v_270, v_271, v_272, v_273, v_275, v_277, v_279, v_280, v_281, v_282, v_284, v_285, v_286, v_291, v_292, v_293, o_1);
input v_338;
input v_339;
input v_340;
input v_341;
input v_342;
input v_343;
input v_344;
input v_345;
input v_346;
input v_347;
input v_348;
input v_349;
input v_350;
input v_351;
input v_352;
input v_353;
input v_354;
input v_355;
input v_356;
input v_357;
input v_358;
input v_359;
input v_360;
input v_361;
input v_362;
input v_363;
input v_364;
input v_365;
input v_366;
input v_367;
input v_368;
input v_369;
input v_370;
input v_371;
input v_372;
input v_373;
input v_374;
input v_375;
input v_376;
input v_377;
input v_378;
input v_379;
input v_380;
input v_381;
input v_296;
input v_297;
input v_298;
input v_299;
input v_300;
input v_301;
input v_302;
input v_303;
input v_304;
input v_305;
input v_306;
input v_307;
input v_308;
input v_309;
input v_310;
input v_311;
input v_312;
input v_313;
input v_314;
input v_315;
input v_316;
input v_317;
input v_318;
input v_319;
input v_320;
input v_321;
input v_322;
input v_323;
input v_324;
input v_325;
input v_326;
input v_327;
input v_328;
input v_329;
input v_330;
input v_331;
input v_332;
input v_333;
input v_334;
input v_335;
input v_336;
input v_337;
input v_5;
input v_7;
input v_8;
input v_10;
input v_12;
input v_15;
input v_16;
input v_18;
input v_24;
input v_26;
input v_27;
input v_30;
input v_31;
input v_40;
input v_42;
input v_45;
input v_51;
input v_53;
input v_55;
input v_57;
input v_59;
input v_63;
input v_66;
input v_67;
input v_70;
input v_71;
input v_72;
input v_74;
input v_77;
input v_78;
input v_79;
input v_81;
input v_82;
input v_87;
input v_88;
input v_89;
input v_94;
input v_95;
input v_97;
input v_99;
input v_100;
input v_101;
input v_102;
input v_105;
input v_106;
input v_107;
input v_108;
input v_109;
input v_112;
input v_114;
input v_116;
input v_119;
input v_121;
input v_122;
input v_123;
input v_124;
input v_126;
input v_128;
input v_130;
input v_131;
input v_132;
input v_133;
input v_136;
input v_138;
input v_139;
input v_140;
input v_141;
input v_143;
input v_145;
input v_146;
input v_147;
input v_148;
input v_151;
input v_154;
input v_155;
input v_157;
input v_159;
input v_161;
input v_163;
input v_166;
input v_167;
input v_169;
input v_172;
input v_173;
input v_175;
input v_176;
input v_177;
input v_178;
input v_179;
input v_180;
input v_182;
input v_183;
input v_184;
input v_185;
input v_186;
input v_187;
input v_189;
input v_190;
input v_191;
input v_192;
input v_193;
input v_194;
input v_195;
input v_196;
input v_197;
input v_198;
input v_200;
input v_201;
input v_203;
input v_205;
input v_206;
input v_209;
input v_211;
input v_212;
input v_214;
input v_216;
input v_217;
input v_218;
input v_220;
input v_221;
input v_222;
input v_224;
input v_226;
input v_227;
input v_228;
input v_230;
input v_231;
input v_233;
input v_234;
input v_236;
input v_237;
input v_238;
input v_239;
input v_240;
input v_242;
input v_243;
input v_245;
input v_246;
input v_247;
input v_250;
input v_251;
input v_255;
input v_256;
input v_259;
input v_260;
input v_261;
input v_267;
input v_269;
input v_270;
input v_271;
input v_272;
input v_273;
input v_275;
input v_277;
input v_279;
input v_280;
input v_281;
input v_282;
input v_284;
input v_285;
input v_286;
input v_291;
input v_292;
input v_293;
output o_1;
wire v_2;
wire v_3;
wire v_4;
wire v_6;
wire v_9;
wire v_11;
wire v_13;
wire v_14;
wire v_17;
wire v_19;
wire v_20;
wire v_21;
wire v_22;
wire v_23;
wire v_25;
wire v_28;
wire v_29;
wire v_32;
wire v_33;
wire v_34;
wire v_35;
wire v_36;
wire v_37;
wire v_38;
wire v_39;
wire v_41;
wire v_43;
wire v_44;
wire v_46;
wire v_47;
wire v_48;
wire v_49;
wire v_50;
wire v_52;
wire v_54;
wire v_56;
wire v_58;
wire v_60;
wire v_61;
wire v_62;
wire v_64;
wire v_65;
wire v_68;
wire v_69;
wire v_73;
wire v_75;
wire v_76;
wire v_80;
wire v_83;
wire v_84;
wire v_85;
wire v_86;
wire v_90;
wire v_91;
wire v_92;
wire v_93;
wire v_96;
wire v_98;
wire v_103;
wire v_104;
wire v_110;
wire v_111;
wire v_113;
wire v_115;
wire v_117;
wire v_118;
wire v_120;
wire v_125;
wire v_127;
wire v_129;
wire v_134;
wire v_135;
wire v_137;
wire v_142;
wire v_144;
wire v_149;
wire v_150;
wire v_152;
wire v_153;
wire v_156;
wire v_158;
wire v_160;
wire v_162;
wire v_164;
wire v_165;
wire v_168;
wire v_170;
wire v_171;
wire v_174;
wire v_181;
wire v_188;
wire v_199;
wire v_202;
wire v_204;
wire v_207;
wire v_208;
wire v_210;
wire v_213;
wire v_215;
wire v_219;
wire v_223;
wire v_225;
wire v_229;
wire v_232;
wire v_235;
wire v_241;
wire v_244;
wire v_248;
wire v_249;
wire v_252;
wire v_253;
wire v_254;
wire v_257;
wire v_258;
wire v_262;
wire v_263;
wire v_264;
wire v_265;
wire v_266;
wire v_268;
wire v_274;
wire v_276;
wire v_278;
wire v_283;
wire v_287;
wire v_288;
wire v_289;
wire v_290;
wire v_294;
wire v_295;
wire v_426;
wire x_1;
wire x_2;
wire x_3;
wire x_4;
wire x_5;
wire x_6;
wire x_7;
wire x_8;
wire x_9;
wire x_10;
wire x_11;
wire x_12;
wire x_13;
wire x_14;
wire x_15;
wire x_16;
wire x_17;
wire x_18;
wire x_19;
wire x_20;
wire x_21;
wire x_22;
wire x_23;
wire x_24;
wire x_25;
wire x_26;
wire x_27;
wire x_28;
wire x_29;
wire x_30;
wire x_31;
wire x_32;
wire x_33;
wire x_34;
wire x_35;
wire x_36;
wire x_37;
wire x_38;
wire x_39;
wire x_40;
wire x_41;
wire x_42;
wire x_43;
wire x_44;
wire x_45;
wire x_46;
wire x_47;
wire x_48;
wire x_49;
wire x_50;
wire x_51;
wire x_52;
wire x_53;
wire x_54;
wire x_55;
wire x_56;
wire x_57;
wire x_58;
wire x_59;
wire x_60;
wire x_61;
wire x_62;
wire x_63;
wire x_64;
wire x_65;
wire x_66;
wire x_67;
wire x_68;
wire x_69;
wire x_70;
wire x_71;
wire x_72;
wire x_73;
wire x_74;
wire x_75;
wire x_76;
wire x_77;
wire x_78;
wire x_79;
wire x_80;
wire x_81;
wire x_82;
wire x_83;
wire x_84;
wire x_85;
wire x_86;
wire x_87;
wire x_88;
wire x_89;
wire x_90;
wire x_91;
wire x_92;
wire x_93;
wire x_94;
wire x_95;
wire x_96;
wire x_97;
wire x_98;
wire x_99;
wire x_100;
wire x_101;
wire x_102;
wire x_103;
wire x_104;
wire x_105;
wire x_106;
wire x_107;
wire x_108;
wire x_109;
wire x_110;
wire x_111;
wire x_112;
wire x_113;
wire x_114;
wire x_115;
wire x_116;
wire x_117;
wire x_118;
wire x_119;
wire x_120;
wire x_121;
wire x_122;
wire x_123;
wire x_124;
wire x_125;
wire x_126;
wire x_127;
wire x_128;
wire x_129;
wire x_130;
wire x_131;
wire x_132;
wire x_133;
wire x_134;
wire x_135;
wire x_136;
wire x_137;
wire x_138;
wire x_139;
wire x_140;
wire x_141;
wire x_142;
wire x_143;
wire x_144;
wire x_145;
wire x_146;
wire x_147;
wire x_148;
wire x_149;
wire x_150;
wire x_151;
wire x_152;
wire x_153;
wire x_154;
wire x_155;
wire x_156;
wire x_157;
wire x_158;
wire x_159;
wire x_160;
wire x_161;
wire x_162;
wire x_163;
wire x_164;
wire x_165;
wire x_166;
wire x_167;
wire x_168;
wire x_169;
wire x_170;
wire x_171;
wire x_172;
wire x_173;
wire x_174;
wire x_175;
wire x_176;
wire x_177;
wire x_178;
wire x_179;
wire x_180;
wire x_181;
wire x_182;
wire x_183;
wire x_184;
wire x_185;
wire x_186;
wire x_187;
wire x_188;
wire x_189;
wire x_190;
wire x_191;
wire x_192;
wire x_193;
wire x_194;
wire x_195;
wire x_196;
wire x_197;
wire x_198;
wire x_199;
wire x_200;
wire x_201;
wire x_202;
wire x_203;
wire x_204;
wire x_205;
wire x_206;
wire x_207;
wire x_208;
wire x_209;
wire x_210;
wire x_211;
wire x_212;
wire x_213;
wire x_214;
wire x_215;
wire x_216;
wire x_217;
wire x_218;
wire x_219;
wire x_220;
wire x_221;
wire x_222;
wire x_223;
wire x_224;
wire x_225;
wire x_226;
wire x_227;
wire x_228;
wire x_229;
wire x_230;
wire x_231;
wire x_232;
wire x_233;
wire x_234;
wire x_235;
wire x_236;
wire x_237;
wire x_238;
wire x_239;
wire x_240;
wire x_241;
wire x_242;
wire x_243;
wire x_244;
wire x_245;
wire x_246;
wire x_247;
wire x_248;
wire x_249;
wire x_250;
wire x_251;
wire x_252;
wire x_253;
wire x_254;
wire x_255;
wire x_256;
wire x_257;
wire x_258;
wire x_259;
wire x_260;
wire x_261;
wire x_262;
wire x_263;
wire x_264;
wire x_265;
wire x_266;
wire x_267;
wire x_268;
wire x_269;
wire x_270;
wire x_271;
wire x_272;
wire x_273;
wire x_274;
wire x_275;
wire x_276;
wire x_277;
wire x_278;
wire x_279;
wire x_280;
wire x_281;
wire x_282;
wire x_283;
wire x_284;
wire x_285;
wire x_286;
wire x_287;
wire x_288;
wire x_289;
wire x_290;
wire x_291;
wire x_292;
wire x_293;
wire x_294;
wire x_295;
wire x_296;
wire x_297;
wire x_298;
wire x_299;
wire x_300;
wire x_301;
wire x_302;
wire x_303;
wire x_304;
wire x_305;
wire x_306;
wire x_307;
wire x_308;
wire x_309;
wire x_310;
wire x_311;
wire x_312;
wire x_313;
wire x_314;
wire x_315;
wire x_316;
wire x_317;
wire x_318;
wire x_319;
wire x_320;
wire x_321;
wire x_322;
wire x_323;
wire x_324;
wire x_325;
wire x_326;
wire x_327;
wire x_328;
wire x_329;
wire x_330;
wire x_331;
wire x_332;
wire x_333;
wire x_334;
wire x_335;
wire x_336;
wire x_337;
wire x_338;
wire x_339;
wire x_340;
wire x_341;
wire x_342;
wire x_343;
wire x_344;
wire x_345;
wire x_346;
wire x_347;
wire x_348;
wire x_349;
wire x_350;
wire x_351;
wire x_352;
wire x_353;
wire x_354;
wire x_355;
wire x_356;
wire x_357;
wire x_358;
wire x_359;
wire x_360;
wire x_361;
wire x_362;
wire x_363;
wire x_364;
wire x_365;
wire x_366;
wire x_367;
wire x_368;
wire x_369;
wire x_370;
wire x_371;
wire x_372;
wire x_373;
wire x_374;
wire x_375;
wire x_376;
wire x_377;
wire x_378;
wire x_379;
wire x_380;
wire x_381;
wire x_382;
wire x_383;
wire x_384;
wire x_385;
wire x_386;
wire x_387;
wire x_388;
wire x_389;
wire x_390;
wire x_391;
wire x_392;
wire x_393;
wire x_394;
wire x_395;
wire x_396;
wire x_397;
wire x_398;
wire x_399;
wire x_400;
wire x_401;
wire x_402;
wire x_403;
wire x_404;
wire x_405;
wire x_406;
wire x_407;
wire x_408;
wire x_409;
wire x_410;
wire x_411;
wire x_412;
wire x_413;
wire x_414;
wire x_415;
wire x_416;
wire x_417;
wire x_418;
wire x_419;
wire x_420;
wire x_421;
wire x_422;
wire x_423;
wire x_424;
wire x_425;
wire x_426;
wire x_427;
wire x_428;
wire x_429;
wire x_430;
wire x_431;
wire x_432;
wire x_433;
wire x_434;
wire x_435;
wire x_436;
wire x_437;
wire x_438;
wire x_439;
wire x_440;
wire x_441;
wire x_442;
wire x_443;
wire x_444;
wire x_445;
wire x_446;
wire x_447;
wire x_448;
wire x_449;
wire x_450;
wire x_451;
wire x_452;
wire x_453;
wire x_454;
wire x_455;
wire x_456;
wire x_457;
wire x_458;
wire x_459;
wire x_460;
wire x_461;
wire x_462;
wire x_463;
wire x_464;
wire x_465;
wire x_466;
wire x_467;
wire x_468;
wire x_469;
wire x_470;
wire x_471;
wire x_472;
wire x_473;
wire x_474;
wire x_475;
wire x_476;
wire x_477;
wire x_478;
wire x_479;
wire x_480;
wire x_481;
wire x_482;
wire x_483;
wire x_484;
wire x_485;
wire x_486;
wire x_487;
wire x_488;
wire x_489;
wire x_490;
wire x_491;
wire x_492;
wire x_493;
wire x_494;
wire x_495;
wire x_496;
wire x_497;
wire x_498;
wire x_499;
wire x_500;
wire x_501;
wire x_502;
wire x_503;
wire x_504;
wire x_505;
wire x_506;
wire x_507;
wire x_508;
wire x_509;
wire x_510;
wire x_511;
wire x_512;
wire x_513;
wire x_514;
wire x_515;
wire x_516;
wire x_517;
wire x_518;
wire x_519;
wire x_520;
wire x_521;
wire x_522;
wire x_523;
wire x_524;
wire x_525;
wire x_526;
wire x_527;
wire x_528;
wire x_529;
wire x_530;
wire x_531;
wire x_532;
wire x_533;
wire x_534;
wire x_535;
wire x_536;
wire x_537;
wire x_538;
wire x_539;
wire x_540;
wire x_541;
wire x_542;
wire x_543;
wire x_544;
wire x_545;
wire x_546;
wire x_547;
wire x_548;
wire x_549;
wire x_550;
wire x_551;
wire x_552;
wire x_553;
wire x_554;
wire x_555;
wire x_556;
wire x_557;
wire x_558;
wire x_559;
wire x_560;
wire x_561;
wire x_562;
wire x_563;
wire x_564;
wire x_565;
wire x_566;
wire x_567;
wire x_568;
wire x_569;
wire x_570;
wire x_571;
wire x_572;
wire x_573;
wire x_574;
wire x_575;
wire x_576;
wire x_577;
wire x_578;
wire x_579;
wire x_580;
wire x_581;
wire x_582;
wire x_583;
wire x_584;
wire x_585;
wire x_586;
wire x_587;
wire x_588;
wire x_589;
wire x_590;
wire x_591;
wire x_592;
wire x_593;
wire x_594;
wire x_595;
wire x_596;
wire x_597;
wire x_598;
wire x_599;
wire x_600;
wire x_601;
wire x_602;
wire x_603;
wire x_604;
wire x_605;
wire x_606;
wire x_607;
wire x_608;
wire x_609;
wire x_610;
wire x_611;
wire x_612;
wire x_613;
wire x_614;
wire x_615;
wire x_616;
wire x_617;
wire x_618;
wire x_619;
wire x_620;
wire x_621;
wire x_622;
wire x_623;
wire x_624;
wire x_625;
wire x_626;
wire x_627;
wire x_628;
wire x_629;
wire x_630;
wire x_631;
wire x_632;
wire x_633;
wire x_634;
wire x_635;
wire x_636;
wire x_637;
wire x_638;
wire x_639;
wire x_640;
wire x_641;
wire x_642;
wire x_643;
wire x_644;
wire x_645;
wire x_646;
wire x_647;
wire x_648;
wire x_649;
wire x_650;
wire x_651;
wire x_652;
wire x_653;
wire x_654;
wire x_655;
wire x_656;
wire x_657;
wire x_658;
wire x_659;
wire x_660;
wire x_661;
wire x_662;
wire x_663;
wire x_664;
wire x_665;
wire x_666;
wire x_667;
wire x_668;
wire x_669;
wire x_670;
wire x_671;
wire x_672;
wire x_673;
wire x_674;
wire x_675;
wire x_676;
wire x_677;
wire x_678;
wire x_679;
wire x_680;
wire x_681;
wire x_682;
wire x_683;
wire x_684;
wire x_685;
wire x_686;
wire x_687;
wire x_688;
wire x_689;
wire x_690;
wire x_691;
wire x_692;
wire x_693;
wire x_694;
wire x_695;
wire x_696;
wire x_697;
wire x_698;
wire x_699;
wire x_700;
wire x_701;
wire x_702;
wire x_703;
wire x_704;
wire x_705;
wire x_706;
wire x_707;
wire x_708;
wire x_709;
wire x_710;
wire x_711;
wire x_712;
wire x_713;
wire x_714;
wire x_715;
wire x_716;
wire x_717;
wire x_718;
wire x_719;
wire x_720;
wire x_721;
wire x_722;
wire x_723;
wire x_724;
wire x_725;
wire x_726;
wire x_727;
wire x_728;
wire x_729;
wire x_730;
wire x_731;
wire x_732;
wire x_733;
wire x_734;
wire x_735;
wire x_736;
wire x_737;
wire x_738;
wire x_739;
wire x_740;
wire x_741;
wire x_742;
wire x_743;
wire x_744;
wire x_745;
wire x_746;
wire x_747;
wire x_748;
wire x_749;
wire x_750;
wire x_751;
wire x_752;
wire x_753;
wire x_754;
wire x_755;
wire x_756;
wire x_757;
wire x_758;
wire x_759;
wire x_760;
wire x_761;
wire x_762;
wire x_763;
wire x_764;
wire x_765;
wire x_766;
wire x_767;
wire x_768;
wire x_769;
wire x_770;
wire x_771;
wire x_772;
wire x_773;
wire x_774;
wire x_775;
wire x_776;
wire x_777;
wire x_778;
wire x_779;
wire x_780;
wire x_781;
wire x_782;
wire x_783;
wire x_784;
wire x_785;
wire x_786;
wire x_787;
wire x_788;
wire x_789;
wire x_790;
wire x_791;
wire x_792;
wire x_793;
wire x_794;
wire x_795;
wire x_796;
wire x_797;
wire x_798;
wire x_799;
wire x_800;
wire x_801;
wire x_802;
wire x_803;
wire x_804;
wire x_805;
wire x_806;
wire x_807;
wire x_808;
wire x_809;
wire x_810;
wire x_811;
wire x_812;
wire x_813;
wire x_814;
wire x_815;
wire x_816;
wire x_817;
wire x_818;
wire x_819;
wire x_820;
wire x_821;
wire x_822;
wire x_823;
wire x_824;
wire x_825;
wire x_826;
wire x_827;
wire x_828;
wire x_829;
wire x_830;
wire x_831;
wire x_832;
wire x_833;
wire x_834;
wire x_835;
wire x_836;
wire x_837;
wire x_838;
wire x_839;
wire x_840;
wire x_841;
wire x_842;
wire x_843;
wire x_844;
wire x_845;
wire x_846;
wire x_847;
wire x_848;
wire x_849;
wire x_850;
wire x_851;
wire x_852;
wire x_853;
wire x_854;
wire x_855;
wire x_856;
wire x_857;
wire x_858;
wire x_859;
wire x_860;
wire x_861;
wire x_862;
wire x_863;
wire x_864;
wire x_865;
wire x_866;
wire x_867;
wire x_868;
wire x_869;
wire x_870;
wire x_871;
wire x_872;
wire x_873;
wire x_874;
wire x_875;
wire x_876;
wire x_877;
wire x_878;
wire x_879;
wire x_880;
wire x_881;
wire x_882;
wire x_883;
wire x_884;
wire x_885;
wire x_886;
wire x_887;
wire x_888;
wire x_889;
wire x_890;
wire x_891;
wire x_892;
wire x_893;
wire x_894;
wire x_895;
wire x_896;
wire x_897;
wire x_898;
wire x_899;
wire x_900;
wire x_901;
wire x_902;
wire x_903;
wire x_904;
wire x_905;
wire x_906;
wire x_907;
wire x_908;
wire x_909;
wire x_910;
wire x_911;
wire x_912;
wire x_913;
wire x_914;
wire x_915;
wire x_916;
wire x_917;
wire x_918;
wire x_919;
wire x_920;
wire x_921;
wire x_922;
wire x_923;
wire x_924;
wire x_925;
wire x_926;
wire x_927;
wire x_928;
wire x_929;
wire x_930;
wire x_931;
wire x_932;
wire x_933;
wire x_934;
wire x_935;
wire x_936;
wire x_937;
wire x_938;
wire x_939;
wire x_940;
wire x_941;
wire x_942;
wire x_943;
wire x_944;
wire x_945;
wire x_946;
wire x_947;
wire x_948;
wire x_949;
wire x_950;
wire x_951;
wire x_952;
wire x_953;
wire x_954;
wire x_955;
wire x_956;
wire x_957;
wire x_958;
wire x_959;
wire x_960;
wire x_961;
wire x_962;
wire x_963;
wire x_964;
wire x_965;
wire x_966;
wire x_967;
wire x_968;
wire x_969;
wire x_970;
wire x_971;
wire x_972;
wire x_973;
wire x_974;
wire x_975;
wire x_976;
wire x_977;
wire x_978;
wire x_979;
wire x_980;
wire x_981;
wire x_982;
wire x_983;
wire x_984;
wire x_985;
wire x_986;
wire x_987;
wire x_988;
wire x_989;
wire x_990;
wire x_991;
wire x_992;
wire x_993;
wire x_994;
wire x_995;
wire x_996;
wire x_997;
wire x_998;
wire x_999;
wire x_1000;
wire x_1001;
wire x_1002;
wire x_1003;
wire x_1004;
wire x_1005;
wire x_1006;
wire x_1007;
wire x_1008;
wire x_1009;
wire x_1010;
wire x_1011;
wire x_1012;
wire x_1013;
wire x_1014;
wire x_1015;
wire x_1016;
wire x_1017;
wire x_1018;
wire x_1019;
wire x_1020;
wire x_1021;
wire x_1022;
wire x_1023;
wire x_1024;
wire x_1025;
wire x_1026;
wire x_1027;
wire x_1028;
wire x_1029;
wire x_1030;
wire x_1031;
wire x_1032;
wire x_1033;
wire x_1034;
wire x_1035;
wire x_1036;
wire x_1037;
wire x_1038;
wire x_1039;
wire x_1040;
wire x_1041;
wire x_1042;
wire x_1043;
wire x_1044;
wire x_1045;
wire x_1046;
wire x_1047;
wire x_1048;
wire x_1049;
wire x_1050;
wire x_1051;
wire x_1052;
wire x_1053;
wire x_1054;
wire x_1055;
wire x_1056;
wire x_1057;
wire x_1058;
wire x_1059;
wire x_1060;
wire x_1061;
wire x_1062;
wire x_1063;
wire x_1064;
wire x_1065;
wire x_1066;
wire x_1067;
wire x_1068;
wire x_1069;
wire x_1070;
wire x_1071;
wire x_1072;
wire x_1073;
wire x_1074;
wire x_1075;
wire x_1076;
wire x_1077;
wire x_1078;
wire x_1079;
wire x_1080;
wire x_1081;
wire x_1082;
wire x_1083;
wire x_1084;
wire x_1085;
wire x_1086;
wire x_1087;
wire x_1088;
wire x_1089;
wire x_1090;
wire x_1091;
wire x_1092;
wire x_1093;
wire x_1094;
wire x_1095;
wire x_1096;
wire x_1097;
wire x_1098;
wire x_1099;
wire x_1100;
wire x_1101;
wire x_1102;
wire x_1103;
wire x_1104;
wire x_1105;
wire x_1106;
wire x_1107;
wire x_1108;
wire x_1109;
wire x_1110;
wire x_1111;
wire x_1112;
wire x_1113;
wire x_1114;
wire x_1115;
wire x_1116;
wire x_1117;
wire x_1118;
wire x_1119;
wire x_1120;
wire x_1121;
wire x_1122;
wire x_1123;
wire x_1124;
wire x_1125;
wire x_1126;
wire x_1127;
wire x_1128;
wire x_1129;
wire x_1130;
wire x_1131;
wire x_1132;
wire x_1133;
wire x_1134;
wire x_1135;
wire x_1136;
wire x_1137;
wire x_1138;
wire x_1139;
wire x_1140;
wire x_1141;
wire x_1142;
wire x_1143;
wire x_1144;
wire x_1145;
wire x_1146;
wire x_1147;
wire x_1148;
wire x_1149;
wire x_1150;
wire x_1151;
wire x_1152;
wire x_1153;
wire x_1154;
wire x_1155;
wire x_1156;
wire x_1157;
wire x_1158;
wire x_1159;
wire x_1160;
wire x_1161;
wire x_1162;
wire x_1163;
wire x_1164;
wire x_1165;
wire x_1166;
wire x_1167;
wire x_1168;
wire x_1169;
wire x_1170;
wire x_1171;
wire x_1172;
wire x_1173;
wire x_1174;
wire x_1175;
wire x_1176;
wire x_1177;
wire x_1178;
wire x_1179;
wire x_1180;
wire x_1181;
wire x_1182;
wire x_1183;
wire x_1184;
wire x_1185;
wire x_1186;
wire x_1187;
wire x_1188;
wire x_1189;
wire x_1190;
wire x_1191;
wire x_1192;
wire x_1193;
wire x_1194;
wire x_1195;
wire x_1196;
wire x_1197;
wire x_1198;
wire x_1199;
wire x_1200;
wire x_1201;
wire x_1202;
wire x_1203;
wire x_1204;
wire x_1205;
wire x_1206;
wire x_1207;
wire x_1208;
wire x_1209;
wire x_1210;
wire x_1211;
wire x_1212;
wire x_1213;
wire x_1214;
wire x_1215;
wire x_1216;
wire x_1217;
wire x_1218;
wire x_1219;
wire x_1220;
wire x_1221;
wire x_1222;
wire x_1223;
wire x_1224;
wire x_1225;
wire x_1226;
wire x_1227;
wire x_1228;
wire x_1229;
wire x_1230;
wire x_1231;
wire x_1232;
wire x_1233;
wire x_1234;
wire x_1235;
wire x_1236;
wire x_1237;
wire x_1238;
wire x_1239;
wire x_1240;
wire x_1241;
wire x_1242;
wire x_1243;
wire x_1244;
wire x_1245;
wire x_1246;
wire x_1247;
wire x_1248;
wire x_1249;
wire x_1250;
wire x_1251;
wire x_1252;
wire x_1253;
wire x_1254;
wire x_1255;
wire x_1256;
wire x_1257;
wire x_1258;
wire x_1259;
wire x_1260;
wire x_1261;
wire x_1262;
wire x_1263;
wire x_1264;
wire x_1265;
wire x_1266;
wire x_1267;
wire x_1268;
wire x_1269;
wire x_1270;
wire x_1271;
wire x_1272;
wire x_1273;
wire x_1274;
wire x_1275;
wire x_1276;
wire x_1277;
wire x_1278;
wire x_1279;
wire x_1280;
wire x_1281;
wire x_1282;
wire x_1283;
wire x_1284;
wire x_1285;
wire x_1286;
wire x_1287;
wire x_1288;
wire x_1289;
wire x_1290;
wire x_1291;
wire x_1292;
wire x_1293;
wire x_1294;
wire x_1295;
wire x_1296;
wire x_1297;
wire x_1298;
wire x_1299;
wire x_1300;
wire x_1301;
wire x_1302;
wire x_1303;
wire x_1304;
wire x_1305;
wire x_1306;
wire x_1307;
wire x_1308;
wire x_1309;
wire x_1310;
wire x_1311;
wire x_1312;
wire x_1313;
wire x_1314;
wire x_1315;
wire x_1316;
wire x_1317;
wire x_1318;
wire x_1319;
wire x_1320;
wire x_1321;
wire x_1322;
wire x_1323;
wire x_1324;
wire x_1325;
wire x_1326;
wire x_1327;
wire x_1328;
wire x_1329;
wire x_1330;
wire x_1331;
wire x_1332;
wire x_1333;
wire x_1334;
wire x_1335;
wire x_1336;
wire x_1337;
wire x_1338;
wire x_1339;
wire x_1340;
wire x_1341;
wire x_1342;
wire x_1343;
wire x_1344;
wire x_1345;
wire x_1346;
wire x_1347;
wire x_1348;
wire x_1349;
wire x_1350;
wire x_1351;
wire x_1352;
wire x_1353;
wire x_1354;
wire x_1355;
wire x_1356;
wire x_1357;
wire x_1358;
wire x_1359;
wire x_1360;
wire x_1361;
wire x_1362;
wire x_1363;
wire x_1364;
wire x_1365;
wire x_1366;
wire x_1367;
wire x_1368;
wire x_1369;
wire x_1370;
wire x_1371;
wire x_1372;
wire x_1373;
wire x_1374;
wire x_1375;
wire x_1376;
wire x_1377;
wire x_1378;
wire x_1379;
wire x_1380;
wire x_1381;
wire x_1382;
wire x_1383;
wire x_1384;
wire x_1385;
wire x_1386;
wire x_1387;
wire x_1388;
wire x_1389;
wire x_1390;
wire x_1391;
wire x_1392;
wire x_1393;
wire x_1394;
wire x_1395;
wire x_1396;
wire x_1397;
wire x_1398;
wire x_1399;
wire x_1400;
wire x_1401;
wire x_1402;
wire x_1403;
wire x_1404;
wire x_1405;
wire x_1406;
wire x_1407;
wire x_1408;
wire x_1409;
wire x_1410;
wire x_1411;
wire x_1412;
wire x_1413;
wire x_1414;
wire x_1415;
wire x_1416;
wire x_1417;
wire x_1418;
wire x_1419;
wire x_1420;
wire x_1421;
wire x_1422;
wire x_1423;
wire x_1424;
wire x_1425;
wire x_1426;
wire x_1427;
wire x_1428;
wire x_1429;
wire x_1430;
wire x_1431;
wire x_1432;
wire x_1433;
wire x_1434;
wire x_1435;
wire x_1436;
wire x_1437;
wire x_1438;
wire x_1439;
wire x_1440;
wire x_1441;
wire x_1442;
wire x_1443;
wire x_1444;
wire x_1445;
wire x_1446;
wire x_1447;
wire x_1448;
wire x_1449;
wire x_1450;
wire x_1451;
wire x_1452;
wire x_1453;
wire x_1454;
wire x_1455;
wire x_1456;
wire x_1457;
wire x_1458;
wire x_1459;
wire x_1460;
wire x_1461;
wire x_1462;
wire x_1463;
wire x_1464;
wire x_1465;
wire x_1466;
wire x_1467;
wire x_1468;
wire x_1469;
wire x_1470;
wire x_1471;
wire x_1472;
wire x_1473;
wire x_1474;
wire x_1475;
wire x_1476;
wire x_1477;
wire x_1478;
wire x_1479;
wire x_1480;
wire x_1481;
wire x_1482;
wire x_1483;
wire x_1484;
wire x_1485;
wire x_1486;
wire x_1487;
wire x_1488;
wire x_1489;
wire x_1490;
wire x_1491;
wire x_1492;
wire x_1493;
wire x_1494;
wire x_1495;
wire x_1496;
wire x_1497;
wire x_1498;
wire x_1499;
wire x_1500;
wire x_1501;
wire x_1502;
wire x_1503;
wire x_1504;
wire x_1505;
wire x_1506;
wire x_1507;
wire x_1508;
wire x_1509;
wire x_1510;
wire x_1511;
wire x_1512;
wire x_1513;
wire x_1514;
wire x_1515;
wire x_1516;
wire x_1517;
wire x_1518;
wire x_1519;
wire x_1520;
wire x_1521;
wire x_1522;
wire x_1523;
wire x_1524;
wire x_1525;
wire x_1526;
wire x_1527;
wire x_1528;
wire x_1529;
wire x_1530;
wire x_1531;
wire x_1532;
wire x_1533;
wire x_1534;
wire x_1535;
wire x_1536;
wire x_1537;
wire x_1538;
wire x_1539;
wire x_1540;
wire x_1541;
wire x_1542;
wire x_1543;
wire x_1544;
wire x_1545;
wire x_1546;
wire x_1547;
wire x_1548;
wire x_1549;
wire x_1550;
wire x_1551;
wire x_1552;
wire x_1553;
wire x_1554;
wire x_1555;
wire x_1556;
wire x_1557;
wire x_1558;
wire x_1559;
wire x_1560;
wire x_1561;
wire x_1562;
wire x_1563;
wire x_1564;
wire x_1565;
wire x_1566;
wire x_1567;
wire x_1568;
wire x_1569;
wire x_1570;
wire x_1571;
wire x_1572;
wire x_1573;
wire x_1574;
wire x_1575;
wire x_1576;
wire x_1577;
wire x_1578;
wire x_1579;
wire x_1580;
wire x_1581;
wire x_1582;
wire x_1583;
wire x_1584;
wire x_1585;
wire x_1586;
wire x_1587;
wire x_1588;
wire x_1589;
wire x_1590;
wire x_1591;
wire x_1592;
wire x_1593;
wire x_1594;
wire x_1595;
wire x_1596;
wire x_1597;
wire x_1598;
wire x_1599;
wire x_1600;
wire x_1601;
wire x_1602;
wire x_1603;
wire x_1604;
wire x_1605;
wire x_1606;
wire x_1607;
wire x_1608;
wire x_1609;
wire x_1610;
wire x_1611;
wire x_1612;
wire x_1613;
wire x_1614;
wire x_1615;
wire x_1616;
wire x_1617;
wire x_1618;
wire x_1619;
wire x_1620;
wire x_1621;
wire x_1622;
wire x_1623;
wire x_1624;
wire x_1625;
wire x_1626;
wire x_1627;
wire x_1628;
wire x_1629;
wire x_1630;
wire x_1631;
wire x_1632;
wire x_1633;
wire x_1634;
wire x_1635;
wire x_1636;
wire x_1637;
wire x_1638;
wire x_1639;
wire x_1640;
wire x_1641;
wire x_1642;
wire x_1643;
wire x_1644;
wire x_1645;
wire x_1646;
wire x_1647;
wire x_1648;
wire x_1649;
wire x_1650;
wire x_1651;
wire x_1652;
wire x_1653;
wire x_1654;
wire x_1655;
wire x_1656;
wire x_1657;
wire x_1658;
wire x_1659;
wire x_1660;
wire x_1661;
wire x_1662;
wire x_1663;
wire x_1664;
wire x_1665;
wire x_1666;
wire x_1667;
wire x_1668;
wire x_1669;
wire x_1670;
wire x_1671;
wire x_1672;
wire x_1673;
wire x_1674;
wire x_1675;
wire x_1676;
wire x_1677;
wire x_1678;
wire x_1679;
wire x_1680;
wire x_1681;
wire x_1682;
wire x_1683;
wire x_1684;
wire x_1685;
wire x_1686;
wire x_1687;
wire x_1688;
wire x_1689;
wire x_1690;
wire x_1691;
wire x_1692;
wire x_1693;
wire x_1694;
wire x_1695;
wire x_1696;
wire x_1697;
wire x_1698;
wire x_1699;
wire x_1700;
wire x_1701;
wire x_1702;
wire x_1703;
wire x_1704;
wire x_1705;
wire x_1706;
wire x_1707;
wire x_1708;
wire x_1709;
wire x_1710;
wire x_1711;
wire x_1712;
wire x_1713;
wire x_1714;
wire x_1715;
wire x_1716;
wire x_1717;
wire x_1718;
wire x_1719;
wire x_1720;
wire x_1721;
wire x_1722;
wire x_1723;
wire x_1724;
wire x_1725;
wire x_1726;
wire x_1727;
wire x_1728;
wire x_1729;
wire x_1730;
wire x_1731;
wire x_1732;
wire x_1733;
wire x_1734;
wire x_1735;
wire x_1736;
wire x_1737;
wire x_1738;
wire x_1739;
wire x_1740;
wire x_1741;
wire x_1742;
wire x_1743;
wire x_1744;
wire x_1745;
wire x_1746;
wire x_1747;
wire x_1748;
wire x_1749;
wire x_1750;
wire x_1751;
wire x_1752;
wire x_1753;
wire x_1754;
wire x_1755;
wire x_1756;
wire x_1757;
wire x_1758;
wire x_1759;
wire x_1760;
wire x_1761;
wire x_1762;
wire x_1763;
wire x_1764;
wire x_1765;
wire x_1766;
wire x_1767;
assign v_4 = 0;
assign v_2 = 1;
assign v_3 = 1;
assign v_426 = 1;
assign v_6 = ~v_7 & v_88 & v_130 & v_174;
assign v_9 = ~v_12 & v_10 & v_14;
assign v_11 = ~v_371 & v_373;
assign v_13 = ~v_369 & ~v_370;
assign v_14 = ~v_15 & v_16;
assign v_17 = v_371 & v_372;
assign v_19 = v_20 & v_21;
assign v_20 = ~v_10 & ~v_12;
assign v_21 = ~v_22 & v_23;
assign v_23 = ~v_24 & ~v_25;
assign v_25 = v_369 & v_26;
assign v_28 = ~v_369 & ~v_370 & ~v_371 & v_29;
assign v_29 = ~v_10 & v_12;
assign v_33 = v_361 & v_34;
assign v_34 = v_35 & v_36;
assign v_35 = v_10 & v_12;
assign v_36 = v_15 & v_16;
assign v_37 = v_22 & v_29 & v_23;
assign v_38 = v_20 & v_39;
assign v_39 = ~v_17 & v_25;
assign v_41 = ~v_361 & v_362;
assign v_43 = ~v_311 & ~v_46 & v_353 & v_44;
assign v_44 = ~v_45 & v_343;
assign v_46 = ~v_47 & v_49;
assign v_47 = ~v_338 & v_339 & v_48;
assign v_48 = ~v_359 & v_360;
assign v_49 = v_344 & v_50;
assign v_50 = v_353 & v_44;
assign v_52 = ~v_47 & v_50;
assign v_54 = ~v_377 & ~v_55 & v_376 & v_378;
assign v_56 = ~v_377 & ~v_57 & v_376 & v_378;
assign v_58 = ~v_359 & ~v_360;
assign v_60 = ~v_376 & ~v_377 & ~v_57 & v_378;
assign v_61 = ~v_376 & ~v_377 & ~v_55 & v_378;
assign v_62 = v_36 & v_29;
assign v_64 = ~v_376 & ~v_378 & v_377 & v_65;
assign v_65 = ~v_47 & ~v_45 & v_66;
assign v_68 = ~v_376 & ~v_378 & v_377 & v_69;
assign v_69 = ~v_45 & ~v_70;
assign v_73 = ~v_354 & v_356;
assign v_75 = ~v_76 & v_356;
assign v_76 = ~v_342 & v_77;
assign v_80 = v_35 & v_21;
assign v_83 = ~v_355 & v_354;
assign v_84 = v_69 & v_85;
assign v_85 = ~v_346 & ~v_377 & ~v_378 & v_376;
assign v_86 = v_65 & v_85;
assign v_90 = v_68 & v_91;
assign v_91 = ~v_353 & ~v_354;
assign v_93 = v_64 & v_91;
assign v_96 = v_29 & v_14;
assign v_98 = ~v_95 & ~v_96;
assign v_104 = ~v_353 & ~v_355 & v_354;
assign v_110 = ~v_353 & ~v_106;
assign v_111 = v_353 & v_103;
assign v_113 = ~v_353 & v_326 & v_75;
assign v_115 = ~v_49 & v_38;
assign v_117 = ~v_46 & v_38;
assign v_118 = ~v_52 & v_103;
assign v_125 = ~v_52 & v_120;
assign v_127 = v_354 & v_355;
assign v_129 = ~v_56 & v_120;
assign v_135 = v_346 & v_364 & v_35 & v_39;
assign v_137 = ~v_136 & v_361;
assign v_142 = ~v_76 & v_73;
assign v_144 = v_363 & v_364;
assign v_150 = v_86 & v_91;
assign v_152 = v_84 & v_91;
assign v_153 = ~v_354 & v_338 & v_356;
assign v_156 = v_338 & v_135;
assign v_158 = v_351 & v_361;
assign v_160 = ~v_93 & v_149;
assign v_164 = v_165 & v_73;
assign v_165 = ~v_338 & ~v_339;
assign v_168 = v_165 & v_135;
assign v_170 = v_361 & v_171;
assign v_171 = ~v_351 & ~v_352;
assign v_174 = ~v_227 & ~v_236 & v_175 & v_216;
assign v_199 = ~v_338 & v_363;
assign v_202 = ~v_319 & ~v_320;
assign v_204 = ~v_205 & ~v_211 & v_206 & v_212;
assign v_207 = ~v_317 & v_318;
assign v_210 = ~v_351 & v_352;
assign v_213 = ~v_165 & v_365;
assign v_215 = ~v_165 & v_367;
assign v_219 = ~v_361 & v_354 & v_362 & v_37;
assign v_223 = v_49 & v_224;
assign v_225 = ~v_338 & v_366;
assign v_232 = v_350 & v_96;
assign v_235 = ~v_93 & v_229;
assign v_241 = ~v_240 & v_361;
assign v_244 = ~v_325 & v_165;
assign v_248 = ~v_357 & ~v_358;
assign v_249 = v_364 & v_365;
assign v_252 = ~v_315 & v_316;
assign v_253 = ~v_323 & ~v_324 & ~v_325 & ~v_326;
assign v_254 = ~v_313 & ~v_314 & ~v_321 & ~v_322;
assign v_257 = ~v_311 & ~v_312 & ~v_319 & ~v_320;
assign v_258 = v_259 & v_260 & v_261 & v_262;
assign v_262 = v_32 & v_263 & v_264 & v_181;
assign v_265 = v_266 & v_278 & v_285 & v_290;
assign v_266 = v_267 & v_270 & v_274 & v_275;
assign v_274 = v_92 & v_149 & v_188 & v_229;
assign v_278 = v_279 & v_280 & v_281 & v_282;
assign v_283 = ~v_303 & v_345;
assign v_287 = ~v_335 & v_377;
assign v_288 = ~v_328 & v_370;
assign v_290 = v_291 & v_292 & v_293;
assign v_294 = ~v_370 & v_328;
assign v_295 = ~v_344 & v_302;
assign v_22 = v_369 ^ v_15;
assign v_32 = ~v_311 ^ v_353;
assign v_92 = ~v_312 ^ v_354;
assign v_103 = ~v_326 ^ v_368;
assign v_120 = ~v_313 ^ v_355;
assign v_134 = ~v_324 ^ v_366;
assign v_149 = ~v_321 ^ v_363;
assign v_162 = ~v_323 ^ v_365;
assign v_181 = ~v_325 ^ v_367;
assign v_188 = ~v_322 ^ v_364;
assign v_208 = ~v_317 ^ v_359;
assign v_229 = ~v_314 ^ v_356;
assign v_263 = ~v_315 ^ v_357;
assign v_264 = ~v_316 ^ v_358;
assign v_268 = v_307 ^ v_349;
assign v_276 = ~v_309 ^ v_351;
assign v_289 = ~v_305 ^ v_347;
assign x_1 = ~v_265 | v_380 | v_5 | ~v_258;
assign x_2 = ~v_265 | ~v_380 | ~v_5 | ~v_258;
assign x_3 = v_5 | ~v_381 | ~v_6;
assign x_4 = v_5 | v_381 | ~v_251 | ~v_255;
assign x_5 = v_381 | v_251 | ~v_5;
assign x_6 = v_6 | ~v_5 | ~v_381;
assign x_7 = v_381 | v_255 | ~v_5;
assign x_8 = v_7 | v_80 | ~v_8;
assign x_9 = v_7 | v_87 | ~v_80;
assign x_10 = v_7 | v_80 | ~v_81;
assign x_11 = ~v_7 | ~v_80 | ~v_87;
assign x_12 = v_8 | v_80 | v_81 | ~v_7;
assign x_13 = v_8 | v_18 | v_62 | ~v_63;
assign x_14 = v_8 | v_9 | v_18 | v_62;
assign x_15 = ~v_8 | ~v_62;
assign x_16 = ~v_8 | ~v_18;
assign x_17 = v_63 | ~v_8 | ~v_9;
assign x_18 = v_10 | v_370 | ~v_372;
assign x_19 = v_10 | v_372 | v_11 | ~v_370;
assign x_20 = v_10 | v_370 | ~v_369 | ~v_11;
assign x_21 = ~v_10 | ~v_370 | ~v_11;
assign x_22 = v_370 | v_372 | v_11 | ~v_10;
assign x_23 = ~v_10 | ~v_370 | ~v_372;
assign x_24 = v_369 | v_372 | ~v_10 | ~v_11;
assign x_25 = v_12 | v_372 | ~v_371 | ~v_373;
assign x_26 = v_12 | v_371 | v_373 | v_13;
assign x_27 = v_12 | v_371 | ~v_372 | ~v_373;
assign x_28 = v_12 | v_372 | ~v_373 | ~v_13;
assign x_29 = ~v_12 | ~v_371 | ~v_372;
assign x_30 = v_371 | v_372 | v_13 | ~v_12 | ~v_373;
assign x_31 = v_373 | ~v_12 | ~v_371;
assign x_32 = v_373 | ~v_12 | ~v_13;
assign x_33 = v_15 | v_371 | ~v_372;
assign x_34 = v_15 | v_370 | v_371;
assign x_35 = v_15 | v_371 | ~v_373;
assign x_36 = v_15 | v_372 | ~v_370 | ~v_371;
assign x_37 = v_370 | ~v_15 | ~v_371;
assign x_38 = ~v_15 | ~v_371 | ~v_372;
assign x_39 = v_371 | v_372 | v_373 | ~v_15 | ~v_370;
assign x_40 = v_16 | v_369 | v_17 | ~v_370;
assign x_41 = v_16 | v_369 | v_370 | ~v_371;
assign x_42 = ~v_16 | ~v_369;
assign x_43 = ~v_16 | ~v_370 | ~v_17;
assign x_44 = v_370 | v_371 | ~v_16;
assign x_45 = v_18 | v_27 | v_9 | v_59;
assign x_46 = v_18 | v_19 | v_27 | v_9;
assign x_47 = ~v_18 | ~v_9;
assign x_48 = ~v_18 | ~v_27;
assign x_49 = ~v_18 | ~v_19 | ~v_59;
assign x_50 = v_24 | v_369 | v_17;
assign x_51 = v_24 | v_369 | v_370;
assign x_52 = ~v_24 | ~v_369;
assign x_53 = ~v_24 | ~v_370 | ~v_17;
assign x_54 = v_26 | ~v_370 | ~v_371;
assign x_55 = v_26 | ~v_370 | ~v_373;
assign x_56 = v_26 | ~v_370 | ~v_372;
assign x_57 = v_370 | ~v_26;
assign x_58 = v_371 | v_372 | v_373 | ~v_26;
assign x_59 = v_27 | v_30 | v_19 | ~v_53;
assign x_60 = v_27 | v_28 | v_30 | v_19;
assign x_61 = ~v_27 | ~v_19;
assign x_62 = ~v_27 | ~v_30;
assign x_63 = v_53 | ~v_27 | ~v_28;
assign x_64 = v_30 | ~v_31 | ~v_42;
assign x_65 = v_30 | ~v_38 | ~v_42;
assign x_66 = v_30 | ~v_40 | ~v_42;
assign x_67 = v_42 | ~v_30;
assign x_68 = v_31 | v_38 | v_40 | ~v_30;
assign x_69 = v_31 | v_311 | v_37 | ~v_33;
assign x_70 = v_31 | v_33 | v_37 | ~v_32;
assign x_71 = ~v_31 | ~v_37;
assign x_72 = ~v_31 | ~v_311 | ~v_33;
assign x_73 = v_32 | v_33 | ~v_31;
assign x_74 = v_40 | v_311 | ~v_37 | ~v_41;
assign x_75 = v_40 | v_41 | ~v_32 | ~v_37;
assign x_76 = v_37 | ~v_40;
assign x_77 = v_32 | v_41 | ~v_40;
assign x_78 = ~v_40 | ~v_311 | ~v_41;
assign x_79 = v_42 | v_28 | ~v_51;
assign x_80 = v_42 | v_28 | ~v_43;
assign x_81 = v_42 | v_38 | v_28;
assign x_82 = ~v_42 | ~v_28;
assign x_83 = v_43 | v_51 | ~v_42 | ~v_38;
assign x_84 = v_45 | ~v_338 | ~v_359;
assign x_85 = v_45 | v_338 | v_339 | v_359 | v_360;
assign x_86 = v_338 | ~v_45 | ~v_339;
assign x_87 = v_359 | ~v_45 | ~v_338;
assign x_88 = v_359 | ~v_45 | ~v_360;
assign x_89 = v_338 | ~v_45 | ~v_359;
assign x_90 = v_51 | ~v_344 | ~v_32;
assign x_91 = v_51 | v_52 | ~v_32;
assign x_92 = v_32 | ~v_51;
assign x_93 = v_344 | ~v_51 | ~v_52;
assign x_94 = v_53 | ~v_311 | ~v_56;
assign x_95 = v_53 | v_32 | v_54;
assign x_96 = v_53 | v_54 | ~v_56;
assign x_97 = v_53 | v_32 | ~v_311;
assign x_98 = v_56 | ~v_53 | ~v_32;
assign x_99 = v_311 | ~v_53 | ~v_54;
assign x_100 = v_55 | v_359 | ~v_347;
assign x_101 = v_55 | v_347 | v_360 | ~v_348;
assign x_102 = v_55 | v_347 | ~v_359;
assign x_103 = v_55 | v_348 | v_359 | ~v_360;
assign x_104 = ~v_55 | ~v_347 | ~v_359;
assign x_105 = v_347 | v_359 | ~v_55 | ~v_348 | ~v_360;
assign x_106 = v_347 | v_348 | v_359 | v_360 | ~v_55;
assign x_107 = v_57 | v_347 | ~v_348;
assign x_108 = v_57 | v_359 | ~v_347;
assign x_109 = v_57 | v_347 | v_58;
assign x_110 = ~v_57 | ~v_347 | ~v_359;
assign x_111 = v_347 | v_348 | ~v_57 | ~v_58;
assign x_112 = v_59 | v_32 | ~v_311;
assign x_113 = v_59 | v_61 | ~v_60;
assign x_114 = v_59 | v_32 | v_61;
assign x_115 = v_59 | ~v_311 | ~v_60;
assign x_116 = v_60 | ~v_59 | ~v_32;
assign x_117 = v_311 | ~v_59 | ~v_61;
assign x_118 = v_63 | v_67 | ~v_64;
assign x_119 = v_63 | v_32 | v_67;
assign x_120 = ~v_63 | ~v_67;
assign x_121 = v_64 | ~v_63 | ~v_32;
assign x_122 = v_66 | ~v_340 | ~v_359;
assign x_123 = v_66 | v_340 | v_341 | v_359 | v_360;
assign x_124 = v_340 | ~v_66 | ~v_341;
assign x_125 = v_359 | ~v_66 | ~v_340;
assign x_126 = v_359 | ~v_66 | ~v_360;
assign x_127 = v_340 | ~v_66 | ~v_359;
assign x_128 = v_67 | ~v_68 | ~v_78;
assign x_129 = v_67 | v_354 | v_71 | ~v_68;
assign x_130 = v_68 | ~v_67;
assign x_131 = v_78 | ~v_67 | ~v_354;
assign x_132 = v_78 | ~v_67 | ~v_71;
assign x_133 = v_70 | v_359 | ~v_340;
assign x_134 = v_70 | v_340 | v_360 | ~v_341;
assign x_135 = v_70 | v_340 | ~v_359;
assign x_136 = v_70 | v_341 | v_359 | ~v_360;
assign x_137 = ~v_70 | ~v_340 | ~v_359;
assign x_138 = v_340 | v_359 | ~v_70 | ~v_341 | ~v_360;
assign x_139 = v_340 | v_341 | v_359 | v_360 | ~v_70;
assign x_140 = v_71 | v_311 | v_32;
assign x_141 = v_71 | v_75 | ~v_72;
assign x_142 = v_71 | v_32 | v_75;
assign x_143 = v_71 | v_311 | ~v_72;
assign x_144 = ~v_71 | ~v_311 | ~v_75;
assign x_145 = v_72 | ~v_71 | ~v_32;
assign x_146 = v_72 | ~v_342 | ~v_73;
assign x_147 = v_72 | ~v_73 | ~v_74;
assign x_148 = v_73 | ~v_72;
assign x_149 = v_342 | v_74 | ~v_72;
assign x_150 = v_74 | v_357 | ~v_338;
assign x_151 = v_74 | v_338 | v_358 | ~v_339;
assign x_152 = v_74 | v_338 | ~v_357;
assign x_153 = v_74 | v_339 | v_357 | ~v_358;
assign x_154 = ~v_74 | ~v_338 | ~v_357;
assign x_155 = v_338 | v_357 | ~v_74 | ~v_339 | ~v_358;
assign x_156 = v_338 | v_339 | v_357 | v_358 | ~v_74;
assign x_157 = v_77 | ~v_338 | ~v_357;
assign x_158 = v_77 | v_338 | v_339 | v_357 | v_358;
assign x_159 = v_338 | ~v_77 | ~v_339;
assign x_160 = v_357 | ~v_77 | ~v_338;
assign x_161 = v_357 | ~v_77 | ~v_358;
assign x_162 = v_338 | ~v_77 | ~v_357;
assign x_163 = v_78 | v_355 | v_79 | ~v_354;
assign x_164 = v_78 | ~v_354 | ~v_355 | ~v_32;
assign x_165 = v_354 | ~v_78;
assign x_166 = v_32 | ~v_78 | ~v_355;
assign x_167 = v_355 | ~v_78 | ~v_79;
assign x_168 = v_79 | v_311 | v_32;
assign x_169 = v_79 | ~v_77 | ~v_74;
assign x_170 = v_79 | v_311 | ~v_74;
assign x_171 = v_79 | v_32 | ~v_77;
assign x_172 = v_77 | ~v_79 | ~v_311;
assign x_173 = v_74 | ~v_79 | ~v_32;
assign x_174 = v_81 | v_32 | v_82 | ~v_62;
assign x_175 = v_81 | v_82 | ~v_62 | ~v_86;
assign x_176 = v_62 | ~v_81;
assign x_177 = ~v_81 | ~v_82;
assign x_178 = v_86 | ~v_81 | ~v_32;
assign x_179 = v_82 | v_83 | ~v_32 | ~v_84;
assign x_180 = v_82 | v_79 | ~v_83 | ~v_84;
assign x_181 = v_84 | ~v_82;
assign x_182 = ~v_82 | ~v_79 | ~v_83;
assign x_183 = v_32 | v_83 | ~v_82;
assign x_184 = v_87 | v_311 | ~v_345;
assign x_185 = v_87 | v_345 | ~v_32;
assign x_186 = ~v_87 | ~v_311 | ~v_345;
assign x_187 = v_345 | v_32 | ~v_87;
assign x_188 = v_88 | ~v_94 | ~v_100;
assign x_189 = v_88 | v_89 | ~v_9 | ~v_100;
assign x_190 = v_100 | ~v_88;
assign x_191 = v_94 | ~v_88 | ~v_89;
assign x_192 = v_9 | v_94 | ~v_88;
assign x_193 = v_89 | v_312 | ~v_93;
assign x_194 = v_89 | v_90 | v_92;
assign x_195 = v_89 | v_90 | ~v_93;
assign x_196 = v_89 | v_312 | v_92;
assign x_197 = ~v_89 | ~v_312 | ~v_90;
assign x_198 = v_93 | ~v_89 | ~v_92;
assign x_199 = v_94 | v_9 | v_99 | ~v_19;
assign x_200 = v_94 | v_19 | v_9 | ~v_95;
assign x_201 = ~v_94 | ~v_9;
assign x_202 = ~v_94 | ~v_19 | ~v_99;
assign x_203 = v_19 | v_95 | ~v_94;
assign x_204 = v_95 | v_97 | v_98;
assign x_205 = ~v_95 | ~v_96 | ~v_97;
assign x_206 = v_97 | ~v_312 | ~v_350;
assign x_207 = v_97 | v_350 | v_92;
assign x_208 = v_312 | ~v_97 | ~v_350;
assign x_209 = v_350 | ~v_97 | ~v_92;
assign x_210 = v_98 | v_96 | ~v_312 | ~v_33;
assign x_211 = v_98 | v_33 | v_92 | v_96;
assign x_212 = v_312 | ~v_98 | ~v_33;
assign x_213 = v_33 | ~v_98 | ~v_92;
assign x_214 = v_99 | v_61 | ~v_60;
assign x_215 = v_99 | v_92 | ~v_312;
assign x_216 = v_99 | ~v_312 | ~v_60;
assign x_217 = v_99 | v_61 | v_92;
assign x_218 = v_60 | ~v_99 | ~v_92;
assign x_219 = v_312 | ~v_99 | ~v_61;
assign x_220 = v_100 | v_9 | v_101 | v_121;
assign x_221 = v_100 | v_101 | v_119 | ~v_9;
assign x_222 = ~v_100 | ~v_101;
assign x_223 = v_9 | ~v_100 | ~v_121;
assign x_224 = ~v_100 | ~v_9 | ~v_119;
assign x_225 = v_101 | ~v_62 | ~v_102;
assign x_226 = v_101 | v_62 | ~v_114;
assign x_227 = v_101 | v_62 | ~v_107;
assign x_228 = v_102 | ~v_101 | ~v_62;
assign x_229 = v_62 | v_107 | v_114 | ~v_101;
assign x_230 = v_102 | v_105 | ~v_86;
assign x_231 = v_102 | v_103 | v_104;
assign x_232 = v_102 | v_103 | v_105;
assign x_233 = v_86 | ~v_102 | ~v_103;
assign x_234 = ~v_102 | ~v_104 | ~v_105;
assign x_235 = ~v_102 | ~v_103 | ~v_105;
assign x_236 = v_105 | ~v_353 | ~v_84;
assign x_237 = v_105 | v_83 | ~v_84;
assign x_238 = v_105 | v_106 | ~v_84;
assign x_239 = v_84 | ~v_105;
assign x_240 = v_353 | ~v_105 | ~v_83 | ~v_106;
assign x_241 = v_106 | ~v_77 | ~v_74;
assign x_242 = v_106 | v_103 | ~v_326;
assign x_243 = v_106 | ~v_326 | ~v_74;
assign x_244 = v_106 | v_103 | ~v_77;
assign x_245 = v_74 | ~v_106 | ~v_103;
assign x_246 = v_326 | v_77 | ~v_106;
assign x_247 = v_107 | v_108 | ~v_9 | ~v_64;
assign x_248 = v_107 | v_103 | v_108 | ~v_9;
assign x_249 = v_9 | ~v_107;
assign x_250 = ~v_107 | ~v_108;
assign x_251 = v_64 | ~v_107 | ~v_103;
assign x_252 = v_108 | ~v_68 | ~v_109;
assign x_253 = v_108 | ~v_68 | ~v_112;
assign x_254 = v_108 | ~v_68 | ~v_111;
assign x_255 = v_68 | ~v_108;
assign x_256 = v_109 | v_111 | v_112 | ~v_108;
assign x_257 = v_109 | v_355 | ~v_354 | ~v_110;
assign x_258 = v_109 | ~v_354 | ~v_355 | ~v_103;
assign x_259 = v_354 | ~v_109;
assign x_260 = v_103 | ~v_109 | ~v_355;
assign x_261 = v_355 | v_110 | ~v_109;
assign x_262 = v_112 | v_354 | ~v_113;
assign x_263 = v_112 | v_354 | v_72 | ~v_103;
assign x_264 = ~v_112 | ~v_354;
assign x_265 = v_113 | ~v_112 | ~v_72;
assign x_266 = v_103 | v_113 | ~v_112;
assign x_267 = v_114 | v_9 | v_103 | v_116;
assign x_268 = v_114 | v_9 | v_116 | ~v_115;
assign x_269 = ~v_114 | ~v_9;
assign x_270 = ~v_114 | ~v_116;
assign x_271 = v_115 | ~v_114 | ~v_103;
assign x_272 = v_116 | ~v_117 | ~v_118;
assign x_273 = v_116 | v_326 | ~v_50 | ~v_117;
assign x_274 = v_117 | ~v_116;
assign x_275 = v_118 | ~v_116 | ~v_326;
assign x_276 = v_50 | v_118 | ~v_116;
assign x_277 = v_119 | v_120 | ~v_313;
assign x_278 = v_119 | v_90 | ~v_93;
assign x_279 = v_119 | v_90 | v_120;
assign x_280 = v_119 | ~v_313 | ~v_93;
assign x_281 = v_313 | ~v_119 | ~v_90;
assign x_282 = v_93 | ~v_119 | ~v_120;
assign x_283 = v_121 | ~v_19 | ~v_122;
assign x_284 = v_121 | v_19 | ~v_128;
assign x_285 = v_121 | v_19 | ~v_123;
assign x_286 = v_122 | ~v_121 | ~v_19;
assign x_287 = v_19 | v_123 | v_128 | ~v_121;
assign x_288 = v_122 | v_313 | ~v_60;
assign x_289 = v_122 | v_61 | v_120;
assign x_290 = v_122 | v_61 | ~v_60;
assign x_291 = v_122 | v_313 | v_120;
assign x_292 = v_60 | ~v_122 | ~v_120;
assign x_293 = ~v_122 | ~v_313 | ~v_61;
assign x_294 = v_123 | v_28 | v_124 | ~v_115;
assign x_295 = v_123 | v_28 | v_120 | v_124;
assign x_296 = ~v_123 | ~v_28;
assign x_297 = ~v_123 | ~v_124;
assign x_298 = v_115 | ~v_123 | ~v_120;
assign x_299 = v_124 | ~v_117 | ~v_125;
assign x_300 = v_124 | ~v_117 | ~v_126;
assign x_301 = v_117 | ~v_124;
assign x_302 = v_125 | v_126 | ~v_124;
assign x_303 = v_126 | v_313 | v_127 | ~v_50;
assign x_304 = v_126 | ~v_313 | ~v_50 | ~v_127;
assign x_305 = v_50 | ~v_126;
assign x_306 = v_127 | ~v_126 | ~v_313;
assign x_307 = v_313 | ~v_126 | ~v_127;
assign x_308 = v_128 | v_313 | v_129 | ~v_28;
assign x_309 = v_128 | v_54 | v_129 | ~v_28;
assign x_310 = v_28 | ~v_128;
assign x_311 = ~v_128 | ~v_129;
assign x_312 = ~v_128 | ~v_313 | ~v_54;
assign x_313 = v_130 | ~v_62 | ~v_146;
assign x_314 = v_130 | ~v_131 | ~v_146;
assign x_315 = v_130 | ~v_140 | ~v_146;
assign x_316 = v_146 | ~v_130;
assign x_317 = v_62 | v_131 | v_140 | ~v_130;
assign x_318 = v_131 | v_9 | v_132 | v_139;
assign x_319 = v_131 | v_9 | v_132 | ~v_138;
assign x_320 = ~v_131 | ~v_9;
assign x_321 = ~v_131 | ~v_132;
assign x_322 = v_138 | ~v_131 | ~v_139;
assign x_323 = v_132 | v_38 | v_136 | ~v_34;
assign x_324 = v_132 | v_34 | v_38 | ~v_133;
assign x_325 = ~v_132 | ~v_38;
assign x_326 = ~v_132 | ~v_34 | ~v_136;
assign x_327 = v_34 | v_133 | ~v_132;
assign x_328 = v_133 | v_134 | v_135;
assign x_329 = v_133 | v_338 | v_134;
assign x_330 = v_133 | ~v_324 | ~v_338 | ~v_135;
assign x_331 = v_338 | ~v_133 | ~v_134;
assign x_332 = v_135 | ~v_133 | ~v_134;
assign x_333 = v_324 | ~v_133 | ~v_338 | ~v_135;
assign x_334 = v_136 | v_137 | ~v_134;
assign x_335 = v_361 | v_134 | ~v_136;
assign x_336 = v_137 | v_324 | ~v_351 | ~v_361;
assign x_337 = v_137 | v_324 | ~v_361 | ~v_363;
assign x_338 = v_137 | v_351 | v_363 | ~v_324 | ~v_361;
assign x_339 = ~v_137 | ~v_324 | ~v_351;
assign x_340 = ~v_137 | ~v_324 | ~v_363;
assign x_341 = v_324 | v_351 | v_363 | ~v_137;
assign x_342 = v_138 | v_50 | ~v_134;
assign x_343 = v_138 | v_338 | ~v_134;
assign x_344 = v_134 | ~v_138;
assign x_345 = ~v_138 | ~v_338 | ~v_50;
assign x_346 = v_139 | ~v_324 | ~v_38;
assign x_347 = v_139 | v_338 | ~v_38;
assign x_348 = v_139 | v_50 | ~v_38;
assign x_349 = v_38 | ~v_139;
assign x_350 = v_324 | ~v_139 | ~v_338 | ~v_50;
assign x_351 = v_140 | ~v_9 | ~v_141;
assign x_352 = v_140 | v_93 | ~v_9 | ~v_134;
assign x_353 = v_9 | ~v_140;
assign x_354 = v_141 | ~v_140 | ~v_93;
assign x_355 = v_134 | v_141 | ~v_140;
assign x_356 = v_141 | v_324 | ~v_145;
assign x_357 = v_141 | ~v_142 | ~v_143 | ~v_145;
assign x_358 = v_145 | ~v_141;
assign x_359 = v_142 | ~v_141 | ~v_324;
assign x_360 = v_143 | ~v_141 | ~v_324;
assign x_361 = v_143 | v_338 | v_359 | ~v_144;
assign x_362 = v_143 | v_338 | v_359 | ~v_357;
assign x_363 = ~v_143 | ~v_338;
assign x_364 = ~v_143 | ~v_359;
assign x_365 = v_357 | v_144 | ~v_143;
assign x_366 = v_145 | ~v_324 | ~v_90;
assign x_367 = v_145 | v_72 | ~v_90;
assign x_368 = v_145 | v_143 | ~v_90;
assign x_369 = v_90 | ~v_145;
assign x_370 = v_324 | ~v_145 | ~v_72 | ~v_143;
assign x_371 = v_146 | v_147 | ~v_166;
assign x_372 = v_146 | v_147 | v_161 | ~v_62;
assign x_373 = ~v_146 | ~v_147;
assign x_374 = v_166 | ~v_146 | ~v_161;
assign x_375 = v_62 | v_166 | ~v_146;
assign x_376 = v_147 | ~v_62 | ~v_148;
assign x_377 = v_147 | v_62 | ~v_159;
assign x_378 = v_147 | v_62 | ~v_154;
assign x_379 = v_148 | ~v_147 | ~v_62;
assign x_380 = v_62 | v_154 | v_159 | ~v_147;
assign x_381 = v_148 | v_151 | ~v_150;
assign x_382 = v_148 | v_149 | v_151;
assign x_383 = ~v_148 | ~v_151;
assign x_384 = v_150 | ~v_148 | ~v_149;
assign x_385 = v_151 | ~v_321 | ~v_152 | ~v_153;
assign x_386 = v_151 | v_153 | ~v_149 | ~v_152;
assign x_387 = v_152 | ~v_151;
assign x_388 = v_321 | ~v_151 | ~v_153;
assign x_389 = v_149 | v_153 | ~v_151;
assign x_390 = v_154 | v_9 | v_155 | v_157;
assign x_391 = v_154 | v_34 | v_9 | v_155;
assign x_392 = ~v_154 | ~v_155;
assign x_393 = ~v_154 | ~v_9;
assign x_394 = ~v_154 | ~v_34 | ~v_157;
assign x_395 = v_155 | v_34 | v_156 | ~v_149;
assign x_396 = v_155 | v_321 | v_34 | ~v_156;
assign x_397 = ~v_155 | ~v_34;
assign x_398 = v_156 | v_149 | ~v_155;
assign x_399 = ~v_155 | ~v_321 | ~v_156;
assign x_400 = v_157 | v_158 | ~v_149;
assign x_401 = v_157 | ~v_321 | ~v_158;
assign x_402 = v_149 | v_158 | ~v_157;
assign x_403 = v_321 | ~v_157 | ~v_158;
assign x_404 = v_159 | v_160 | ~v_321 | ~v_9;
assign x_405 = v_159 | v_90 | v_160 | ~v_9;
assign x_406 = v_9 | ~v_159;
assign x_407 = ~v_159 | ~v_160;
assign x_408 = v_321 | ~v_159 | ~v_90;
assign x_409 = v_161 | v_163 | ~v_150;
assign x_410 = v_161 | v_162 | v_163;
assign x_411 = ~v_161 | ~v_163;
assign x_412 = v_150 | ~v_161 | ~v_162;
assign x_413 = v_163 | ~v_323 | ~v_152 | ~v_164;
assign x_414 = v_163 | v_164 | ~v_152 | ~v_162;
assign x_415 = v_152 | ~v_163;
assign x_416 = v_323 | ~v_163 | ~v_164;
assign x_417 = v_162 | v_164 | ~v_163;
assign x_418 = v_166 | ~v_9 | ~v_172;
assign x_419 = v_166 | ~v_167 | ~v_172;
assign x_420 = v_166 | ~v_169 | ~v_172;
assign x_421 = v_172 | ~v_166;
assign x_422 = v_9 | v_167 | v_169 | ~v_166;
assign x_423 = v_167 | v_323 | v_34 | ~v_168;
assign x_424 = v_167 | v_34 | v_168 | ~v_162;
assign x_425 = ~v_167 | ~v_34;
assign x_426 = ~v_167 | ~v_323 | ~v_168;
assign x_427 = v_162 | v_168 | ~v_167;
assign x_428 = v_169 | ~v_323 | ~v_34 | ~v_170;
assign x_429 = v_169 | v_170 | ~v_34 | ~v_162;
assign x_430 = v_34 | ~v_169;
assign x_431 = v_323 | ~v_169 | ~v_170;
assign x_432 = v_162 | v_170 | ~v_169;
assign x_433 = v_172 | v_62 | v_173;
assign x_434 = v_172 | v_323 | v_62 | ~v_90;
assign x_435 = ~v_172 | ~v_62;
assign x_436 = ~v_172 | ~v_323 | ~v_173;
assign x_437 = v_90 | ~v_172 | ~v_173;
assign x_438 = v_173 | ~v_9 | ~v_93;
assign x_439 = v_173 | v_162 | ~v_9;
assign x_440 = v_9 | ~v_173;
assign x_441 = v_93 | ~v_173 | ~v_162;
assign x_442 = v_175 | v_62 | ~v_190;
assign x_443 = v_175 | ~v_176 | ~v_184 | ~v_190;
assign x_444 = v_190 | ~v_175;
assign x_445 = v_176 | ~v_175 | ~v_62;
assign x_446 = v_184 | ~v_175 | ~v_62;
assign x_447 = v_176 | v_177 | ~v_182;
assign x_448 = v_176 | v_150 | v_177 | ~v_181;
assign x_449 = ~v_176 | ~v_177;
assign x_450 = v_182 | ~v_176 | ~v_150;
assign x_451 = v_181 | v_182 | ~v_176;
assign x_452 = v_177 | v_179 | ~v_150;
assign x_453 = v_177 | v_178 | v_179;
assign x_454 = ~v_177 | ~v_179;
assign x_455 = v_150 | ~v_177 | ~v_178;
assign x_456 = v_178 | ~v_315 | ~v_357;
assign x_457 = v_178 | v_315 | v_357 | ~v_316 | ~v_358;
assign x_458 = v_178 | v_315 | v_316 | v_357 | v_358;
assign x_459 = v_357 | ~v_178 | ~v_315;
assign x_460 = v_315 | v_358 | ~v_178 | ~v_316;
assign x_461 = v_315 | ~v_178 | ~v_357;
assign x_462 = v_316 | v_357 | ~v_178 | ~v_358;
assign x_463 = v_179 | v_73 | v_180 | ~v_152;
assign x_464 = v_179 | ~v_73 | ~v_152 | ~v_178;
assign x_465 = v_152 | ~v_179;
assign x_466 = v_73 | ~v_179 | ~v_180;
assign x_467 = v_178 | ~v_179 | ~v_73;
assign x_468 = v_180 | v_338 | ~v_315;
assign x_469 = v_180 | v_315 | v_339 | ~v_316;
assign x_470 = v_180 | v_315 | ~v_338;
assign x_471 = v_180 | v_316 | v_338 | ~v_339;
assign x_472 = ~v_180 | ~v_315 | ~v_338;
assign x_473 = v_315 | v_338 | ~v_180 | ~v_316 | ~v_339;
assign x_474 = v_315 | v_316 | v_338 | v_339 | ~v_180;
assign x_475 = v_182 | ~v_73 | ~v_152 | ~v_183;
assign x_476 = v_182 | v_73 | ~v_152 | ~v_181;
assign x_477 = v_152 | ~v_182;
assign x_478 = v_183 | ~v_182 | ~v_73;
assign x_479 = v_73 | v_181 | ~v_182;
assign x_480 = v_183 | ~v_325 | ~v_365;
assign x_481 = v_183 | ~v_325 | ~v_165;
assign x_482 = v_183 | v_325 | v_365 | v_165;
assign x_483 = v_325 | ~v_183 | ~v_165;
assign x_484 = v_365 | v_165 | ~v_183 | ~v_325;
assign x_485 = v_325 | ~v_183 | ~v_365;
assign x_486 = v_184 | v_187 | ~v_185;
assign x_487 = v_184 | v_150 | v_187 | ~v_134;
assign x_488 = ~v_184 | ~v_187;
assign x_489 = v_185 | ~v_184 | ~v_150;
assign x_490 = v_134 | v_185 | ~v_184;
assign x_491 = v_185 | v_73 | ~v_134 | ~v_152;
assign x_492 = v_185 | ~v_73 | ~v_152 | ~v_186;
assign x_493 = v_152 | ~v_185;
assign x_494 = v_186 | ~v_185 | ~v_73;
assign x_495 = v_73 | v_134 | ~v_185;
assign x_496 = v_186 | ~v_324 | ~v_338;
assign x_497 = v_186 | ~v_324 | ~v_363;
assign x_498 = v_186 | v_324 | v_338 | v_363;
assign x_499 = v_324 | ~v_186 | ~v_363;
assign x_500 = v_338 | v_363 | ~v_186 | ~v_324;
assign x_501 = v_324 | ~v_186 | ~v_338;
assign x_502 = v_187 | v_189 | ~v_150;
assign x_503 = v_187 | v_188 | v_189;
assign x_504 = ~v_187 | ~v_189;
assign x_505 = v_150 | ~v_187 | ~v_188;
assign x_506 = v_189 | v_73 | ~v_152 | ~v_188;
assign x_507 = v_189 | ~v_322 | ~v_73 | ~v_152;
assign x_508 = v_152 | ~v_189;
assign x_509 = v_73 | v_188 | ~v_189;
assign x_510 = v_322 | ~v_189 | ~v_73;
assign x_511 = v_190 | v_9 | v_201 | ~v_204;
assign x_512 = v_190 | v_201 | ~v_191 | ~v_204;
assign x_513 = v_204 | ~v_190;
assign x_514 = ~v_190 | ~v_201;
assign x_515 = v_191 | ~v_190 | ~v_9;
assign x_516 = v_191 | v_192 | v_200;
assign x_517 = v_191 | v_322 | v_192 | ~v_90;
assign x_518 = ~v_191 | ~v_192;
assign x_519 = ~v_191 | ~v_322 | ~v_200;
assign x_520 = v_90 | ~v_191 | ~v_200;
assign x_521 = v_192 | v_193 | ~v_195;
assign x_522 = v_192 | v_90 | v_193;
assign x_523 = v_192 | v_142 | v_193;
assign x_524 = ~v_192 | ~v_193;
assign x_525 = v_195 | ~v_192 | ~v_90 | ~v_142;
assign x_526 = v_193 | v_93 | v_194;
assign x_527 = v_193 | v_72 | v_194 | ~v_68;
assign x_528 = ~v_193 | ~v_194;
assign x_529 = ~v_193 | ~v_72 | ~v_93;
assign x_530 = v_68 | ~v_193 | ~v_93;
assign x_531 = v_194 | v_374 | ~v_332;
assign x_532 = v_194 | v_332 | v_375 | ~v_333;
assign x_533 = v_194 | v_332 | ~v_374;
assign x_534 = v_194 | v_333 | v_374 | ~v_375;
assign x_535 = ~v_194 | ~v_332 | ~v_374;
assign x_536 = v_332 | v_374 | ~v_194 | ~v_333 | ~v_375;
assign x_537 = v_332 | v_333 | v_374 | v_375 | ~v_194;
assign x_538 = v_195 | ~v_74 | ~v_196;
assign x_539 = v_195 | ~v_77 | ~v_197;
assign x_540 = v_195 | ~v_77 | ~v_74;
assign x_541 = v_195 | ~v_196 | ~v_197;
assign x_542 = v_74 | v_197 | ~v_195;
assign x_543 = v_77 | v_196 | ~v_195;
assign x_544 = v_196 | v_357 | ~v_332;
assign x_545 = v_196 | v_332 | v_358 | ~v_333;
assign x_546 = v_196 | v_332 | ~v_357;
assign x_547 = v_196 | v_333 | v_357 | ~v_358;
assign x_548 = ~v_196 | ~v_332 | ~v_357;
assign x_549 = v_332 | v_357 | ~v_196 | ~v_333 | ~v_358;
assign x_550 = v_332 | v_333 | v_357 | v_358 | ~v_196;
assign x_551 = v_197 | v_332 | ~v_342 | ~v_198;
assign x_552 = v_197 | v_199 | ~v_332 | ~v_342;
assign x_553 = v_342 | ~v_197;
assign x_554 = ~v_197 | ~v_332 | ~v_199;
assign x_555 = v_332 | v_198 | ~v_197;
assign x_556 = v_198 | v_333 | v_365;
assign x_557 = v_198 | v_333 | ~v_165;
assign x_558 = ~v_198 | ~v_333;
assign x_559 = v_165 | ~v_198 | ~v_365;
assign x_560 = v_200 | v_62 | ~v_93;
assign x_561 = v_200 | v_62 | v_188;
assign x_562 = ~v_200 | ~v_62;
assign x_563 = v_93 | ~v_200 | ~v_188;
assign x_564 = v_201 | v_33 | v_37 | ~v_203;
assign x_565 = v_201 | v_37 | v_202 | ~v_33;
assign x_566 = ~v_201 | ~v_37;
assign x_567 = ~v_201 | ~v_33 | ~v_202;
assign x_568 = v_33 | v_203 | ~v_201;
assign x_569 = v_203 | v_361 | ~v_319;
assign x_570 = v_203 | v_319 | v_362 | ~v_320;
assign x_571 = v_203 | v_319 | ~v_361;
assign x_572 = v_203 | v_320 | v_361 | ~v_362;
assign x_573 = ~v_203 | ~v_319 | ~v_361;
assign x_574 = v_319 | v_361 | ~v_203 | ~v_320 | ~v_362;
assign x_575 = v_319 | v_320 | v_361 | v_362 | ~v_203;
assign x_576 = v_205 | v_319 | ~v_320 | ~v_37;
assign x_577 = v_205 | v_361 | ~v_319 | ~v_37;
assign x_578 = v_205 | v_319 | ~v_361 | ~v_37;
assign x_579 = v_37 | ~v_205;
assign x_580 = ~v_205 | ~v_319 | ~v_361;
assign x_581 = v_319 | v_320 | v_361 | ~v_205;
assign x_582 = v_206 | ~v_48 | ~v_207 | ~v_209;
assign x_583 = v_206 | v_48 | v_207 | ~v_208 | ~v_209;
assign x_584 = v_48 | ~v_206 | ~v_207;
assign x_585 = v_207 | ~v_206 | ~v_48;
assign x_586 = v_209 | ~v_206;
assign x_587 = v_48 | v_208 | ~v_206;
assign x_588 = v_209 | ~v_309 | ~v_380;
assign x_589 = v_209 | v_310 | ~v_380;
assign x_590 = v_209 | ~v_380 | ~v_210;
assign x_591 = v_380 | ~v_209;
assign x_592 = v_309 | v_210 | ~v_209 | ~v_310;
assign x_593 = v_211 | v_351 | ~v_309;
assign x_594 = v_211 | v_309 | v_310 | ~v_351;
assign x_595 = v_211 | v_310 | v_351 | ~v_352;
assign x_596 = v_309 | ~v_211 | ~v_310;
assign x_597 = ~v_211 | ~v_309 | ~v_351;
assign x_598 = v_309 | v_351 | v_352 | ~v_211;
assign x_599 = v_212 | v_214 | ~v_342;
assign x_600 = v_212 | v_213 | v_199 | v_214;
assign x_601 = ~v_212 | ~v_214;
assign x_602 = v_342 | ~v_212 | ~v_213;
assign x_603 = v_342 | ~v_212 | ~v_199;
assign x_604 = v_214 | v_344 | ~v_215;
assign x_605 = v_214 | v_338 | v_344 | ~v_366;
assign x_606 = ~v_214 | ~v_344;
assign x_607 = v_215 | ~v_214 | ~v_338;
assign x_608 = v_366 | v_215 | ~v_214;
assign x_609 = v_216 | v_217 | ~v_9;
assign x_610 = v_216 | v_217 | v_222 | v_226;
assign x_611 = ~v_216 | ~v_217;
assign x_612 = v_9 | ~v_216 | ~v_226;
assign x_613 = v_9 | ~v_216 | ~v_222;
assign x_614 = v_217 | v_62 | v_218 | ~v_221;
assign x_615 = v_217 | v_9 | v_62 | v_218;
assign x_616 = ~v_217 | ~v_218;
assign x_617 = ~v_217 | ~v_62;
assign x_618 = v_221 | ~v_217 | ~v_9;
assign x_619 = v_218 | v_9 | v_219 | ~v_178;
assign x_620 = v_218 | v_9 | v_220 | ~v_219;
assign x_621 = ~v_218 | ~v_9;
assign x_622 = v_178 | v_219 | ~v_218;
assign x_623 = ~v_218 | ~v_219 | ~v_220;
assign x_624 = v_220 | v_351 | ~v_315;
assign x_625 = v_220 | v_315 | v_352 | ~v_316;
assign x_626 = v_220 | v_315 | ~v_351;
assign x_627 = v_220 | v_316 | v_351 | ~v_352;
assign x_628 = ~v_220 | ~v_315 | ~v_351;
assign x_629 = v_315 | v_351 | ~v_220 | ~v_316 | ~v_352;
assign x_630 = v_315 | v_316 | v_351 | v_352 | ~v_220;
assign x_631 = v_221 | v_90 | v_178;
assign x_632 = v_221 | ~v_93 | ~v_180;
assign x_633 = v_221 | v_90 | ~v_93;
assign x_634 = v_221 | v_178 | ~v_180;
assign x_635 = v_180 | ~v_221 | ~v_90;
assign x_636 = v_93 | ~v_221 | ~v_178;
assign x_637 = v_222 | v_38 | ~v_194;
assign x_638 = v_222 | v_223 | ~v_38 | ~v_46;
assign x_639 = v_222 | v_223 | ~v_194;
assign x_640 = ~v_222 | ~v_38 | ~v_223;
assign x_641 = v_38 | v_194 | ~v_222;
assign x_642 = v_46 | v_194 | ~v_222;
assign x_643 = v_224 | v_332 | ~v_333;
assign x_644 = v_224 | ~v_332 | ~v_225;
assign x_645 = v_224 | v_332 | ~v_215;
assign x_646 = v_225 | ~v_224 | ~v_332;
assign x_647 = v_332 | v_333 | v_215 | ~v_224;
assign x_648 = v_226 | v_322 | v_62 | ~v_33;
assign x_649 = v_226 | v_33 | v_62 | v_188;
assign x_650 = ~v_226 | ~v_62;
assign x_651 = v_33 | ~v_226 | ~v_188;
assign x_652 = ~v_226 | ~v_322 | ~v_33;
assign x_653 = v_227 | ~v_62 | ~v_228;
assign x_654 = v_227 | v_62 | ~v_234;
assign x_655 = v_227 | v_62 | ~v_230;
assign x_656 = v_228 | ~v_227 | ~v_62;
assign x_657 = v_62 | v_230 | v_234 | ~v_227;
assign x_658 = v_228 | v_314 | ~v_150;
assign x_659 = v_228 | v_152 | v_229;
assign x_660 = v_228 | v_152 | ~v_150;
assign x_661 = v_228 | v_314 | v_229;
assign x_662 = v_150 | ~v_228 | ~v_229;
assign x_663 = ~v_228 | ~v_314 | ~v_152;
assign x_664 = v_230 | v_9 | v_231 | ~v_233;
assign x_665 = v_230 | v_28 | v_9 | v_231;
assign x_666 = ~v_230 | ~v_231;
assign x_667 = ~v_230 | ~v_9;
assign x_668 = v_233 | ~v_230 | ~v_28;
assign x_669 = v_231 | v_314 | v_28 | ~v_232;
assign x_670 = v_231 | v_28 | v_232 | ~v_229;
assign x_671 = ~v_231 | ~v_28;
assign x_672 = ~v_231 | ~v_314 | ~v_232;
assign x_673 = v_229 | v_232 | ~v_231;
assign x_674 = v_233 | v_229 | ~v_314;
assign x_675 = v_233 | v_54 | ~v_56;
assign x_676 = v_233 | v_54 | v_229;
assign x_677 = v_233 | ~v_314 | ~v_56;
assign x_678 = v_314 | ~v_233 | ~v_54;
assign x_679 = v_56 | ~v_233 | ~v_229;
assign x_680 = v_234 | v_314 | v_235 | ~v_9;
assign x_681 = v_234 | v_90 | v_235 | ~v_9;
assign x_682 = v_9 | ~v_234;
assign x_683 = ~v_234 | ~v_235;
assign x_684 = ~v_234 | ~v_314 | ~v_90;
assign x_685 = v_236 | v_62 | v_237 | ~v_245;
assign x_686 = v_236 | v_9 | v_62 | v_237;
assign x_687 = ~v_236 | ~v_237;
assign x_688 = ~v_236 | ~v_62;
assign x_689 = v_245 | ~v_236 | ~v_9;
assign x_690 = v_237 | v_9 | v_238 | v_243;
assign x_691 = v_237 | v_9 | v_238 | ~v_242;
assign x_692 = ~v_237 | ~v_9;
assign x_693 = ~v_237 | ~v_238;
assign x_694 = v_242 | ~v_237 | ~v_243;
assign x_695 = v_238 | v_38 | v_240 | ~v_34;
assign x_696 = v_238 | v_34 | v_38 | ~v_239;
assign x_697 = ~v_238 | ~v_38;
assign x_698 = ~v_238 | ~v_34 | ~v_240;
assign x_699 = v_34 | v_239 | ~v_238;
assign x_700 = v_239 | v_165 | v_181;
assign x_701 = v_239 | v_135 | v_181;
assign x_702 = v_239 | ~v_325 | ~v_165 | ~v_135;
assign x_703 = v_165 | ~v_239 | ~v_181;
assign x_704 = v_135 | ~v_239 | ~v_181;
assign x_705 = v_325 | ~v_239 | ~v_165 | ~v_135;
assign x_706 = v_240 | v_241 | ~v_181;
assign x_707 = v_361 | v_181 | ~v_240;
assign x_708 = v_241 | v_325 | ~v_361 | ~v_365;
assign x_709 = v_241 | v_325 | ~v_361 | ~v_171;
assign x_710 = v_241 | v_365 | v_171 | ~v_325 | ~v_361;
assign x_711 = ~v_241 | ~v_325 | ~v_365;
assign x_712 = v_325 | v_365 | v_171 | ~v_241;
assign x_713 = ~v_241 | ~v_325 | ~v_171;
assign x_714 = v_242 | v_50 | ~v_181;
assign x_715 = v_242 | v_165 | ~v_181;
assign x_716 = v_181 | ~v_242;
assign x_717 = ~v_242 | ~v_165 | ~v_50;
assign x_718 = v_243 | v_244 | ~v_38;
assign x_719 = v_243 | v_50 | ~v_38;
assign x_720 = v_38 | ~v_243;
assign x_721 = ~v_243 | ~v_50 | ~v_244;
assign x_722 = v_245 | v_246 | ~v_93;
assign x_723 = v_245 | v_181 | v_246;
assign x_724 = ~v_245 | ~v_246;
assign x_725 = v_93 | ~v_245 | ~v_181;
assign x_726 = v_246 | v_325 | ~v_250;
assign x_727 = v_246 | ~v_142 | ~v_247 | ~v_250;
assign x_728 = v_250 | ~v_246;
assign x_729 = v_142 | ~v_246 | ~v_325;
assign x_730 = v_247 | ~v_246 | ~v_325;
assign x_731 = v_247 | v_58 | v_165 | ~v_249;
assign x_732 = v_247 | v_58 | v_165 | ~v_248;
assign x_733 = ~v_247 | ~v_58;
assign x_734 = ~v_247 | ~v_165;
assign x_735 = v_248 | v_249 | ~v_247;
assign x_736 = v_250 | ~v_325 | ~v_90;
assign x_737 = v_250 | v_72 | ~v_90;
assign x_738 = v_250 | v_247 | ~v_90;
assign x_739 = v_90 | ~v_250;
assign x_740 = v_325 | ~v_250 | ~v_72 | ~v_247;
assign x_741 = v_251 | v_252 | ~v_253 | ~v_254;
assign x_742 = v_251 | ~v_207 | ~v_253 | ~v_254;
assign x_743 = v_254 | ~v_251;
assign x_744 = v_253 | ~v_251;
assign x_745 = v_207 | ~v_251 | ~v_252;
assign x_746 = v_255 | v_315 | v_256 | ~v_257;
assign x_747 = v_255 | v_256 | ~v_317 | ~v_257;
assign x_748 = v_257 | ~v_255;
assign x_749 = ~v_255 | ~v_256;
assign x_750 = v_317 | ~v_255 | ~v_315;
assign x_751 = v_256 | v_316 | v_317 | ~v_318;
assign x_752 = v_256 | v_315 | v_316 | ~v_317;
assign x_753 = ~v_256 | ~v_316;
assign x_754 = v_317 | v_318 | ~v_256;
assign x_755 = ~v_256 | ~v_315 | ~v_317;
assign x_756 = v_259 | v_337 | v_379 | ~v_120 | ~v_162;
assign x_757 = v_259 | ~v_337 | ~v_379 | ~v_120 | ~v_162;
assign x_758 = v_162 | ~v_259;
assign x_759 = v_379 | ~v_259 | ~v_337;
assign x_760 = v_120 | ~v_259;
assign x_761 = v_337 | ~v_259 | ~v_379;
assign x_762 = v_260 | ~v_330 | ~v_372 | ~v_103;
assign x_763 = v_260 | v_330 | v_372 | ~v_103;
assign x_764 = v_103 | ~v_260;
assign x_765 = v_372 | ~v_260 | ~v_330;
assign x_766 = v_330 | ~v_260 | ~v_372;
assign x_767 = v_261 | v_318 | v_360 | ~v_306 | ~v_348;
assign x_768 = v_261 | v_306 | v_348 | ~v_318 | ~v_360;
assign x_769 = v_261 | v_306 | v_318 | v_348 | v_360;
assign x_770 = v_261 | ~v_306 | ~v_318 | ~v_348 | ~v_360;
assign x_771 = v_348 | ~v_261 | ~v_306;
assign x_772 = v_306 | ~v_261 | ~v_348;
assign x_773 = v_318 | ~v_261 | ~v_360;
assign x_774 = v_360 | ~v_261 | ~v_318;
assign x_775 = v_267 | v_331 | v_373 | v_268 | ~v_269;
assign x_776 = v_267 | v_268 | ~v_331 | ~v_373 | ~v_269;
assign x_777 = ~v_267 | ~v_268;
assign x_778 = v_331 | ~v_267 | ~v_373;
assign x_779 = v_269 | ~v_267;
assign x_780 = v_373 | ~v_267 | ~v_331;
assign x_781 = v_269 | v_298 | v_340 | ~v_297 | ~v_339;
assign x_782 = v_269 | v_297 | v_339 | ~v_298 | ~v_340;
assign x_783 = v_269 | v_297 | v_298 | v_339 | v_340;
assign x_784 = v_269 | ~v_297 | ~v_298 | ~v_339 | ~v_340;
assign x_785 = v_339 | ~v_269 | ~v_297;
assign x_786 = v_297 | ~v_269 | ~v_339;
assign x_787 = v_298 | ~v_269 | ~v_340;
assign x_788 = v_340 | ~v_269 | ~v_298;
assign x_789 = v_270 | v_296 | v_338 | ~v_271 | ~v_273;
assign x_790 = v_270 | ~v_296 | ~v_338 | ~v_271 | ~v_273;
assign x_791 = v_273 | ~v_270;
assign x_792 = v_338 | ~v_270 | ~v_296;
assign x_793 = v_271 | ~v_270;
assign x_794 = v_296 | ~v_270 | ~v_338;
assign x_795 = v_271 | ~v_310 | ~v_352 | ~v_272;
assign x_796 = v_271 | v_310 | v_352 | ~v_272;
assign x_797 = v_272 | ~v_271;
assign x_798 = v_352 | ~v_271 | ~v_310;
assign x_799 = v_310 | ~v_271 | ~v_352;
assign x_800 = v_272 | v_308 | v_335;
assign x_801 = v_272 | ~v_350 | ~v_377;
assign x_802 = v_272 | v_308 | ~v_377;
assign x_803 = v_272 | v_335 | ~v_350;
assign x_804 = v_350 | ~v_272 | ~v_308;
assign x_805 = v_377 | ~v_272 | ~v_335;
assign x_806 = v_273 | ~v_308 | ~v_381;
assign x_807 = v_273 | v_350 | ~v_381;
assign x_808 = v_381 | ~v_273;
assign x_809 = v_308 | ~v_273 | ~v_350;
assign x_810 = v_275 | v_317 | v_359 | ~v_276 | ~v_277;
assign x_811 = v_275 | ~v_317 | ~v_359 | ~v_276 | ~v_277;
assign x_812 = v_277 | ~v_275;
assign x_813 = v_359 | ~v_275 | ~v_317;
assign x_814 = v_276 | ~v_275;
assign x_815 = v_317 | ~v_275 | ~v_359;
assign x_816 = v_277 | ~v_304 | ~v_346 | ~v_134;
assign x_817 = v_277 | v_304 | v_346 | ~v_134;
assign x_818 = v_134 | ~v_277;
assign x_819 = v_346 | ~v_277 | ~v_304;
assign x_820 = v_304 | ~v_277 | ~v_346;
assign x_821 = v_279 | v_333 | v_375 | ~v_332 | ~v_374;
assign x_822 = v_279 | v_332 | v_374 | ~v_333 | ~v_375;
assign x_823 = v_279 | v_332 | v_333 | v_374 | v_375;
assign x_824 = v_279 | ~v_332 | ~v_333 | ~v_374 | ~v_375;
assign x_825 = v_374 | ~v_279 | ~v_332;
assign x_826 = v_332 | ~v_279 | ~v_374;
assign x_827 = v_333 | ~v_279 | ~v_375;
assign x_828 = v_375 | ~v_279 | ~v_333;
assign x_829 = v_280 | v_320 | v_362 | ~v_319 | ~v_361;
assign x_830 = v_280 | v_319 | v_361 | ~v_320 | ~v_362;
assign x_831 = v_280 | v_319 | v_320 | v_361 | v_362;
assign x_832 = v_280 | ~v_319 | ~v_320 | ~v_361 | ~v_362;
assign x_833 = v_361 | ~v_280 | ~v_319;
assign x_834 = v_319 | ~v_280 | ~v_361;
assign x_835 = v_320 | ~v_280 | ~v_362;
assign x_836 = v_362 | ~v_280 | ~v_320;
assign x_837 = v_281 | v_300 | v_342 | ~v_299;
assign x_838 = v_281 | v_341 | ~v_300 | ~v_342;
assign x_839 = v_281 | ~v_299 | ~v_300 | ~v_342;
assign x_840 = v_281 | v_300 | v_341 | v_342;
assign x_841 = v_300 | ~v_281 | ~v_342;
assign x_842 = v_342 | ~v_281 | ~v_300;
assign x_843 = v_299 | ~v_281 | ~v_341;
assign x_844 = v_282 | v_336 | v_283 | ~v_284;
assign x_845 = v_282 | v_283 | ~v_378 | ~v_284;
assign x_846 = v_284 | ~v_282;
assign x_847 = ~v_282 | ~v_283;
assign x_848 = v_378 | ~v_282 | ~v_336;
assign x_849 = v_284 | ~v_301 | ~v_341;
assign x_850 = v_284 | v_299 | v_343;
assign x_851 = v_284 | v_299 | ~v_301;
assign x_852 = v_284 | v_343 | ~v_341;
assign x_853 = v_341 | ~v_284 | ~v_299;
assign x_854 = v_301 | ~v_284 | ~v_343;
assign x_855 = v_285 | v_334 | v_376 | ~v_286 | ~v_289;
assign x_856 = v_285 | ~v_334 | ~v_376 | ~v_286 | ~v_289;
assign x_857 = v_289 | ~v_285;
assign x_858 = v_376 | ~v_285 | ~v_334;
assign x_859 = v_286 | ~v_285;
assign x_860 = v_334 | ~v_285 | ~v_376;
assign x_861 = v_286 | v_327 | v_369 | v_287 | v_288;
assign x_862 = v_286 | v_287 | v_288 | ~v_327 | ~v_369;
assign x_863 = ~v_286 | ~v_287;
assign x_864 = v_369 | ~v_286 | ~v_327;
assign x_865 = ~v_286 | ~v_288;
assign x_866 = v_327 | ~v_286 | ~v_369;
assign x_867 = v_291 | ~v_302 | ~v_343;
assign x_868 = v_291 | v_301 | v_344;
assign x_869 = v_291 | v_301 | ~v_302;
assign x_870 = v_291 | v_344 | ~v_343;
assign x_871 = v_343 | ~v_291 | ~v_301;
assign x_872 = v_302 | ~v_291 | ~v_344;
assign x_873 = v_292 | ~v_336 | ~v_345;
assign x_874 = v_292 | v_303 | v_378;
assign x_875 = v_292 | v_303 | ~v_336;
assign x_876 = v_292 | v_378 | ~v_345;
assign x_877 = v_345 | ~v_292 | ~v_303;
assign x_878 = v_336 | ~v_292 | ~v_378;
assign x_879 = v_293 | v_329 | v_371 | v_294 | v_295;
assign x_880 = v_293 | v_294 | v_295 | ~v_329 | ~v_371;
assign x_881 = ~v_293 | ~v_294;
assign x_882 = v_371 | ~v_293 | ~v_329;
assign x_883 = ~v_293 | ~v_295;
assign x_884 = v_329 | ~v_293 | ~v_371;
assign x_885 = x_2 & x_3;
assign x_886 = x_1 & x_885;
assign x_887 = x_5 & x_6;
assign x_888 = x_4 & x_887;
assign x_889 = x_886 & x_888;
assign x_890 = x_8 & x_9;
assign x_891 = x_7 & x_890;
assign x_892 = x_10 & x_11;
assign x_893 = x_12 & x_13;
assign x_894 = x_892 & x_893;
assign x_895 = x_891 & x_894;
assign x_896 = x_889 & x_895;
assign x_897 = x_15 & x_16;
assign x_898 = x_14 & x_897;
assign x_899 = x_17 & x_18;
assign x_900 = x_19 & x_20;
assign x_901 = x_899 & x_900;
assign x_902 = x_898 & x_901;
assign x_903 = x_22 & x_23;
assign x_904 = x_21 & x_903;
assign x_905 = x_24 & x_25;
assign x_906 = x_26 & x_27;
assign x_907 = x_905 & x_906;
assign x_908 = x_904 & x_907;
assign x_909 = x_902 & x_908;
assign x_910 = x_896 & x_909;
assign x_911 = x_29 & x_30;
assign x_912 = x_28 & x_911;
assign x_913 = x_31 & x_32;
assign x_914 = x_33 & x_34;
assign x_915 = x_913 & x_914;
assign x_916 = x_912 & x_915;
assign x_917 = x_36 & x_37;
assign x_918 = x_35 & x_917;
assign x_919 = x_38 & x_39;
assign x_920 = x_40 & x_41;
assign x_921 = x_919 & x_920;
assign x_922 = x_918 & x_921;
assign x_923 = x_916 & x_922;
assign x_924 = x_43 & x_44;
assign x_925 = x_42 & x_924;
assign x_926 = x_45 & x_46;
assign x_927 = x_47 & x_48;
assign x_928 = x_926 & x_927;
assign x_929 = x_925 & x_928;
assign x_930 = x_50 & x_51;
assign x_931 = x_49 & x_930;
assign x_932 = x_52 & x_53;
assign x_933 = x_54 & x_55;
assign x_934 = x_932 & x_933;
assign x_935 = x_931 & x_934;
assign x_936 = x_929 & x_935;
assign x_937 = x_923 & x_936;
assign x_938 = x_910 & x_937;
assign x_939 = x_57 & x_58;
assign x_940 = x_56 & x_939;
assign x_941 = x_60 & x_61;
assign x_942 = x_59 & x_941;
assign x_943 = x_940 & x_942;
assign x_944 = x_63 & x_64;
assign x_945 = x_62 & x_944;
assign x_946 = x_65 & x_66;
assign x_947 = x_67 & x_68;
assign x_948 = x_946 & x_947;
assign x_949 = x_945 & x_948;
assign x_950 = x_943 & x_949;
assign x_951 = x_70 & x_71;
assign x_952 = x_69 & x_951;
assign x_953 = x_72 & x_73;
assign x_954 = x_74 & x_75;
assign x_955 = x_953 & x_954;
assign x_956 = x_952 & x_955;
assign x_957 = x_77 & x_78;
assign x_958 = x_76 & x_957;
assign x_959 = x_79 & x_80;
assign x_960 = x_81 & x_82;
assign x_961 = x_959 & x_960;
assign x_962 = x_958 & x_961;
assign x_963 = x_956 & x_962;
assign x_964 = x_950 & x_963;
assign x_965 = x_84 & x_85;
assign x_966 = x_83 & x_965;
assign x_967 = x_86 & x_87;
assign x_968 = x_88 & x_89;
assign x_969 = x_967 & x_968;
assign x_970 = x_966 & x_969;
assign x_971 = x_91 & x_92;
assign x_972 = x_90 & x_971;
assign x_973 = x_93 & x_94;
assign x_974 = x_95 & x_96;
assign x_975 = x_973 & x_974;
assign x_976 = x_972 & x_975;
assign x_977 = x_970 & x_976;
assign x_978 = x_98 & x_99;
assign x_979 = x_97 & x_978;
assign x_980 = x_100 & x_101;
assign x_981 = x_102 & x_103;
assign x_982 = x_980 & x_981;
assign x_983 = x_979 & x_982;
assign x_984 = x_105 & x_106;
assign x_985 = x_104 & x_984;
assign x_986 = x_107 & x_108;
assign x_987 = x_109 & x_110;
assign x_988 = x_986 & x_987;
assign x_989 = x_985 & x_988;
assign x_990 = x_983 & x_989;
assign x_991 = x_977 & x_990;
assign x_992 = x_964 & x_991;
assign x_993 = x_938 & x_992;
assign x_994 = x_112 & x_113;
assign x_995 = x_111 & x_994;
assign x_996 = x_115 & x_116;
assign x_997 = x_114 & x_996;
assign x_998 = x_995 & x_997;
assign x_999 = x_118 & x_119;
assign x_1000 = x_117 & x_999;
assign x_1001 = x_120 & x_121;
assign x_1002 = x_122 & x_123;
assign x_1003 = x_1001 & x_1002;
assign x_1004 = x_1000 & x_1003;
assign x_1005 = x_998 & x_1004;
assign x_1006 = x_125 & x_126;
assign x_1007 = x_124 & x_1006;
assign x_1008 = x_127 & x_128;
assign x_1009 = x_129 & x_130;
assign x_1010 = x_1008 & x_1009;
assign x_1011 = x_1007 & x_1010;
assign x_1012 = x_132 & x_133;
assign x_1013 = x_131 & x_1012;
assign x_1014 = x_134 & x_135;
assign x_1015 = x_136 & x_137;
assign x_1016 = x_1014 & x_1015;
assign x_1017 = x_1013 & x_1016;
assign x_1018 = x_1011 & x_1017;
assign x_1019 = x_1005 & x_1018;
assign x_1020 = x_139 & x_140;
assign x_1021 = x_138 & x_1020;
assign x_1022 = x_141 & x_142;
assign x_1023 = x_143 & x_144;
assign x_1024 = x_1022 & x_1023;
assign x_1025 = x_1021 & x_1024;
assign x_1026 = x_146 & x_147;
assign x_1027 = x_145 & x_1026;
assign x_1028 = x_148 & x_149;
assign x_1029 = x_150 & x_151;
assign x_1030 = x_1028 & x_1029;
assign x_1031 = x_1027 & x_1030;
assign x_1032 = x_1025 & x_1031;
assign x_1033 = x_153 & x_154;
assign x_1034 = x_152 & x_1033;
assign x_1035 = x_155 & x_156;
assign x_1036 = x_157 & x_158;
assign x_1037 = x_1035 & x_1036;
assign x_1038 = x_1034 & x_1037;
assign x_1039 = x_160 & x_161;
assign x_1040 = x_159 & x_1039;
assign x_1041 = x_162 & x_163;
assign x_1042 = x_164 & x_165;
assign x_1043 = x_1041 & x_1042;
assign x_1044 = x_1040 & x_1043;
assign x_1045 = x_1038 & x_1044;
assign x_1046 = x_1032 & x_1045;
assign x_1047 = x_1019 & x_1046;
assign x_1048 = x_167 & x_168;
assign x_1049 = x_166 & x_1048;
assign x_1050 = x_169 & x_170;
assign x_1051 = x_171 & x_172;
assign x_1052 = x_1050 & x_1051;
assign x_1053 = x_1049 & x_1052;
assign x_1054 = x_174 & x_175;
assign x_1055 = x_173 & x_1054;
assign x_1056 = x_176 & x_177;
assign x_1057 = x_178 & x_179;
assign x_1058 = x_1056 & x_1057;
assign x_1059 = x_1055 & x_1058;
assign x_1060 = x_1053 & x_1059;
assign x_1061 = x_181 & x_182;
assign x_1062 = x_180 & x_1061;
assign x_1063 = x_183 & x_184;
assign x_1064 = x_185 & x_186;
assign x_1065 = x_1063 & x_1064;
assign x_1066 = x_1062 & x_1065;
assign x_1067 = x_188 & x_189;
assign x_1068 = x_187 & x_1067;
assign x_1069 = x_190 & x_191;
assign x_1070 = x_192 & x_193;
assign x_1071 = x_1069 & x_1070;
assign x_1072 = x_1068 & x_1071;
assign x_1073 = x_1066 & x_1072;
assign x_1074 = x_1060 & x_1073;
assign x_1075 = x_195 & x_196;
assign x_1076 = x_194 & x_1075;
assign x_1077 = x_197 & x_198;
assign x_1078 = x_199 & x_200;
assign x_1079 = x_1077 & x_1078;
assign x_1080 = x_1076 & x_1079;
assign x_1081 = x_202 & x_203;
assign x_1082 = x_201 & x_1081;
assign x_1083 = x_204 & x_205;
assign x_1084 = x_206 & x_207;
assign x_1085 = x_1083 & x_1084;
assign x_1086 = x_1082 & x_1085;
assign x_1087 = x_1080 & x_1086;
assign x_1088 = x_209 & x_210;
assign x_1089 = x_208 & x_1088;
assign x_1090 = x_211 & x_212;
assign x_1091 = x_213 & x_214;
assign x_1092 = x_1090 & x_1091;
assign x_1093 = x_1089 & x_1092;
assign x_1094 = x_216 & x_217;
assign x_1095 = x_215 & x_1094;
assign x_1096 = x_218 & x_219;
assign x_1097 = x_220 & x_221;
assign x_1098 = x_1096 & x_1097;
assign x_1099 = x_1095 & x_1098;
assign x_1100 = x_1093 & x_1099;
assign x_1101 = x_1087 & x_1100;
assign x_1102 = x_1074 & x_1101;
assign x_1103 = x_1047 & x_1102;
assign x_1104 = x_993 & x_1103;
assign x_1105 = x_223 & x_224;
assign x_1106 = x_222 & x_1105;
assign x_1107 = x_226 & x_227;
assign x_1108 = x_225 & x_1107;
assign x_1109 = x_1106 & x_1108;
assign x_1110 = x_229 & x_230;
assign x_1111 = x_228 & x_1110;
assign x_1112 = x_231 & x_232;
assign x_1113 = x_233 & x_234;
assign x_1114 = x_1112 & x_1113;
assign x_1115 = x_1111 & x_1114;
assign x_1116 = x_1109 & x_1115;
assign x_1117 = x_236 & x_237;
assign x_1118 = x_235 & x_1117;
assign x_1119 = x_238 & x_239;
assign x_1120 = x_240 & x_241;
assign x_1121 = x_1119 & x_1120;
assign x_1122 = x_1118 & x_1121;
assign x_1123 = x_243 & x_244;
assign x_1124 = x_242 & x_1123;
assign x_1125 = x_245 & x_246;
assign x_1126 = x_247 & x_248;
assign x_1127 = x_1125 & x_1126;
assign x_1128 = x_1124 & x_1127;
assign x_1129 = x_1122 & x_1128;
assign x_1130 = x_1116 & x_1129;
assign x_1131 = x_250 & x_251;
assign x_1132 = x_249 & x_1131;
assign x_1133 = x_252 & x_253;
assign x_1134 = x_254 & x_255;
assign x_1135 = x_1133 & x_1134;
assign x_1136 = x_1132 & x_1135;
assign x_1137 = x_257 & x_258;
assign x_1138 = x_256 & x_1137;
assign x_1139 = x_259 & x_260;
assign x_1140 = x_261 & x_262;
assign x_1141 = x_1139 & x_1140;
assign x_1142 = x_1138 & x_1141;
assign x_1143 = x_1136 & x_1142;
assign x_1144 = x_264 & x_265;
assign x_1145 = x_263 & x_1144;
assign x_1146 = x_266 & x_267;
assign x_1147 = x_268 & x_269;
assign x_1148 = x_1146 & x_1147;
assign x_1149 = x_1145 & x_1148;
assign x_1150 = x_271 & x_272;
assign x_1151 = x_270 & x_1150;
assign x_1152 = x_273 & x_274;
assign x_1153 = x_275 & x_276;
assign x_1154 = x_1152 & x_1153;
assign x_1155 = x_1151 & x_1154;
assign x_1156 = x_1149 & x_1155;
assign x_1157 = x_1143 & x_1156;
assign x_1158 = x_1130 & x_1157;
assign x_1159 = x_278 & x_279;
assign x_1160 = x_277 & x_1159;
assign x_1161 = x_281 & x_282;
assign x_1162 = x_280 & x_1161;
assign x_1163 = x_1160 & x_1162;
assign x_1164 = x_284 & x_285;
assign x_1165 = x_283 & x_1164;
assign x_1166 = x_286 & x_287;
assign x_1167 = x_288 & x_289;
assign x_1168 = x_1166 & x_1167;
assign x_1169 = x_1165 & x_1168;
assign x_1170 = x_1163 & x_1169;
assign x_1171 = x_291 & x_292;
assign x_1172 = x_290 & x_1171;
assign x_1173 = x_293 & x_294;
assign x_1174 = x_295 & x_296;
assign x_1175 = x_1173 & x_1174;
assign x_1176 = x_1172 & x_1175;
assign x_1177 = x_298 & x_299;
assign x_1178 = x_297 & x_1177;
assign x_1179 = x_300 & x_301;
assign x_1180 = x_302 & x_303;
assign x_1181 = x_1179 & x_1180;
assign x_1182 = x_1178 & x_1181;
assign x_1183 = x_1176 & x_1182;
assign x_1184 = x_1170 & x_1183;
assign x_1185 = x_305 & x_306;
assign x_1186 = x_304 & x_1185;
assign x_1187 = x_307 & x_308;
assign x_1188 = x_309 & x_310;
assign x_1189 = x_1187 & x_1188;
assign x_1190 = x_1186 & x_1189;
assign x_1191 = x_312 & x_313;
assign x_1192 = x_311 & x_1191;
assign x_1193 = x_314 & x_315;
assign x_1194 = x_316 & x_317;
assign x_1195 = x_1193 & x_1194;
assign x_1196 = x_1192 & x_1195;
assign x_1197 = x_1190 & x_1196;
assign x_1198 = x_319 & x_320;
assign x_1199 = x_318 & x_1198;
assign x_1200 = x_321 & x_322;
assign x_1201 = x_323 & x_324;
assign x_1202 = x_1200 & x_1201;
assign x_1203 = x_1199 & x_1202;
assign x_1204 = x_326 & x_327;
assign x_1205 = x_325 & x_1204;
assign x_1206 = x_328 & x_329;
assign x_1207 = x_330 & x_331;
assign x_1208 = x_1206 & x_1207;
assign x_1209 = x_1205 & x_1208;
assign x_1210 = x_1203 & x_1209;
assign x_1211 = x_1197 & x_1210;
assign x_1212 = x_1184 & x_1211;
assign x_1213 = x_1158 & x_1212;
assign x_1214 = x_333 & x_334;
assign x_1215 = x_332 & x_1214;
assign x_1216 = x_336 & x_337;
assign x_1217 = x_335 & x_1216;
assign x_1218 = x_1215 & x_1217;
assign x_1219 = x_339 & x_340;
assign x_1220 = x_338 & x_1219;
assign x_1221 = x_341 & x_342;
assign x_1222 = x_343 & x_344;
assign x_1223 = x_1221 & x_1222;
assign x_1224 = x_1220 & x_1223;
assign x_1225 = x_1218 & x_1224;
assign x_1226 = x_346 & x_347;
assign x_1227 = x_345 & x_1226;
assign x_1228 = x_348 & x_349;
assign x_1229 = x_350 & x_351;
assign x_1230 = x_1228 & x_1229;
assign x_1231 = x_1227 & x_1230;
assign x_1232 = x_353 & x_354;
assign x_1233 = x_352 & x_1232;
assign x_1234 = x_355 & x_356;
assign x_1235 = x_357 & x_358;
assign x_1236 = x_1234 & x_1235;
assign x_1237 = x_1233 & x_1236;
assign x_1238 = x_1231 & x_1237;
assign x_1239 = x_1225 & x_1238;
assign x_1240 = x_360 & x_361;
assign x_1241 = x_359 & x_1240;
assign x_1242 = x_362 & x_363;
assign x_1243 = x_364 & x_365;
assign x_1244 = x_1242 & x_1243;
assign x_1245 = x_1241 & x_1244;
assign x_1246 = x_367 & x_368;
assign x_1247 = x_366 & x_1246;
assign x_1248 = x_369 & x_370;
assign x_1249 = x_371 & x_372;
assign x_1250 = x_1248 & x_1249;
assign x_1251 = x_1247 & x_1250;
assign x_1252 = x_1245 & x_1251;
assign x_1253 = x_374 & x_375;
assign x_1254 = x_373 & x_1253;
assign x_1255 = x_376 & x_377;
assign x_1256 = x_378 & x_379;
assign x_1257 = x_1255 & x_1256;
assign x_1258 = x_1254 & x_1257;
assign x_1259 = x_381 & x_382;
assign x_1260 = x_380 & x_1259;
assign x_1261 = x_383 & x_384;
assign x_1262 = x_385 & x_386;
assign x_1263 = x_1261 & x_1262;
assign x_1264 = x_1260 & x_1263;
assign x_1265 = x_1258 & x_1264;
assign x_1266 = x_1252 & x_1265;
assign x_1267 = x_1239 & x_1266;
assign x_1268 = x_388 & x_389;
assign x_1269 = x_387 & x_1268;
assign x_1270 = x_390 & x_391;
assign x_1271 = x_392 & x_393;
assign x_1272 = x_1270 & x_1271;
assign x_1273 = x_1269 & x_1272;
assign x_1274 = x_395 & x_396;
assign x_1275 = x_394 & x_1274;
assign x_1276 = x_397 & x_398;
assign x_1277 = x_399 & x_400;
assign x_1278 = x_1276 & x_1277;
assign x_1279 = x_1275 & x_1278;
assign x_1280 = x_1273 & x_1279;
assign x_1281 = x_402 & x_403;
assign x_1282 = x_401 & x_1281;
assign x_1283 = x_404 & x_405;
assign x_1284 = x_406 & x_407;
assign x_1285 = x_1283 & x_1284;
assign x_1286 = x_1282 & x_1285;
assign x_1287 = x_409 & x_410;
assign x_1288 = x_408 & x_1287;
assign x_1289 = x_411 & x_412;
assign x_1290 = x_413 & x_414;
assign x_1291 = x_1289 & x_1290;
assign x_1292 = x_1288 & x_1291;
assign x_1293 = x_1286 & x_1292;
assign x_1294 = x_1280 & x_1293;
assign x_1295 = x_416 & x_417;
assign x_1296 = x_415 & x_1295;
assign x_1297 = x_418 & x_419;
assign x_1298 = x_420 & x_421;
assign x_1299 = x_1297 & x_1298;
assign x_1300 = x_1296 & x_1299;
assign x_1301 = x_423 & x_424;
assign x_1302 = x_422 & x_1301;
assign x_1303 = x_425 & x_426;
assign x_1304 = x_427 & x_428;
assign x_1305 = x_1303 & x_1304;
assign x_1306 = x_1302 & x_1305;
assign x_1307 = x_1300 & x_1306;
assign x_1308 = x_430 & x_431;
assign x_1309 = x_429 & x_1308;
assign x_1310 = x_432 & x_433;
assign x_1311 = x_434 & x_435;
assign x_1312 = x_1310 & x_1311;
assign x_1313 = x_1309 & x_1312;
assign x_1314 = x_437 & x_438;
assign x_1315 = x_436 & x_1314;
assign x_1316 = x_439 & x_440;
assign x_1317 = x_441 & x_442;
assign x_1318 = x_1316 & x_1317;
assign x_1319 = x_1315 & x_1318;
assign x_1320 = x_1313 & x_1319;
assign x_1321 = x_1307 & x_1320;
assign x_1322 = x_1294 & x_1321;
assign x_1323 = x_1267 & x_1322;
assign x_1324 = x_1213 & x_1323;
assign x_1325 = x_1104 & x_1324;
assign x_1326 = x_444 & x_445;
assign x_1327 = x_443 & x_1326;
assign x_1328 = x_447 & x_448;
assign x_1329 = x_446 & x_1328;
assign x_1330 = x_1327 & x_1329;
assign x_1331 = x_450 & x_451;
assign x_1332 = x_449 & x_1331;
assign x_1333 = x_452 & x_453;
assign x_1334 = x_454 & x_455;
assign x_1335 = x_1333 & x_1334;
assign x_1336 = x_1332 & x_1335;
assign x_1337 = x_1330 & x_1336;
assign x_1338 = x_457 & x_458;
assign x_1339 = x_456 & x_1338;
assign x_1340 = x_459 & x_460;
assign x_1341 = x_461 & x_462;
assign x_1342 = x_1340 & x_1341;
assign x_1343 = x_1339 & x_1342;
assign x_1344 = x_464 & x_465;
assign x_1345 = x_463 & x_1344;
assign x_1346 = x_466 & x_467;
assign x_1347 = x_468 & x_469;
assign x_1348 = x_1346 & x_1347;
assign x_1349 = x_1345 & x_1348;
assign x_1350 = x_1343 & x_1349;
assign x_1351 = x_1337 & x_1350;
assign x_1352 = x_471 & x_472;
assign x_1353 = x_470 & x_1352;
assign x_1354 = x_473 & x_474;
assign x_1355 = x_475 & x_476;
assign x_1356 = x_1354 & x_1355;
assign x_1357 = x_1353 & x_1356;
assign x_1358 = x_478 & x_479;
assign x_1359 = x_477 & x_1358;
assign x_1360 = x_480 & x_481;
assign x_1361 = x_482 & x_483;
assign x_1362 = x_1360 & x_1361;
assign x_1363 = x_1359 & x_1362;
assign x_1364 = x_1357 & x_1363;
assign x_1365 = x_485 & x_486;
assign x_1366 = x_484 & x_1365;
assign x_1367 = x_487 & x_488;
assign x_1368 = x_489 & x_490;
assign x_1369 = x_1367 & x_1368;
assign x_1370 = x_1366 & x_1369;
assign x_1371 = x_492 & x_493;
assign x_1372 = x_491 & x_1371;
assign x_1373 = x_494 & x_495;
assign x_1374 = x_496 & x_497;
assign x_1375 = x_1373 & x_1374;
assign x_1376 = x_1372 & x_1375;
assign x_1377 = x_1370 & x_1376;
assign x_1378 = x_1364 & x_1377;
assign x_1379 = x_1351 & x_1378;
assign x_1380 = x_499 & x_500;
assign x_1381 = x_498 & x_1380;
assign x_1382 = x_502 & x_503;
assign x_1383 = x_501 & x_1382;
assign x_1384 = x_1381 & x_1383;
assign x_1385 = x_505 & x_506;
assign x_1386 = x_504 & x_1385;
assign x_1387 = x_507 & x_508;
assign x_1388 = x_509 & x_510;
assign x_1389 = x_1387 & x_1388;
assign x_1390 = x_1386 & x_1389;
assign x_1391 = x_1384 & x_1390;
assign x_1392 = x_512 & x_513;
assign x_1393 = x_511 & x_1392;
assign x_1394 = x_514 & x_515;
assign x_1395 = x_516 & x_517;
assign x_1396 = x_1394 & x_1395;
assign x_1397 = x_1393 & x_1396;
assign x_1398 = x_519 & x_520;
assign x_1399 = x_518 & x_1398;
assign x_1400 = x_521 & x_522;
assign x_1401 = x_523 & x_524;
assign x_1402 = x_1400 & x_1401;
assign x_1403 = x_1399 & x_1402;
assign x_1404 = x_1397 & x_1403;
assign x_1405 = x_1391 & x_1404;
assign x_1406 = x_526 & x_527;
assign x_1407 = x_525 & x_1406;
assign x_1408 = x_528 & x_529;
assign x_1409 = x_530 & x_531;
assign x_1410 = x_1408 & x_1409;
assign x_1411 = x_1407 & x_1410;
assign x_1412 = x_533 & x_534;
assign x_1413 = x_532 & x_1412;
assign x_1414 = x_535 & x_536;
assign x_1415 = x_537 & x_538;
assign x_1416 = x_1414 & x_1415;
assign x_1417 = x_1413 & x_1416;
assign x_1418 = x_1411 & x_1417;
assign x_1419 = x_540 & x_541;
assign x_1420 = x_539 & x_1419;
assign x_1421 = x_542 & x_543;
assign x_1422 = x_544 & x_545;
assign x_1423 = x_1421 & x_1422;
assign x_1424 = x_1420 & x_1423;
assign x_1425 = x_547 & x_548;
assign x_1426 = x_546 & x_1425;
assign x_1427 = x_549 & x_550;
assign x_1428 = x_551 & x_552;
assign x_1429 = x_1427 & x_1428;
assign x_1430 = x_1426 & x_1429;
assign x_1431 = x_1424 & x_1430;
assign x_1432 = x_1418 & x_1431;
assign x_1433 = x_1405 & x_1432;
assign x_1434 = x_1379 & x_1433;
assign x_1435 = x_554 & x_555;
assign x_1436 = x_553 & x_1435;
assign x_1437 = x_557 & x_558;
assign x_1438 = x_556 & x_1437;
assign x_1439 = x_1436 & x_1438;
assign x_1440 = x_560 & x_561;
assign x_1441 = x_559 & x_1440;
assign x_1442 = x_562 & x_563;
assign x_1443 = x_564 & x_565;
assign x_1444 = x_1442 & x_1443;
assign x_1445 = x_1441 & x_1444;
assign x_1446 = x_1439 & x_1445;
assign x_1447 = x_567 & x_568;
assign x_1448 = x_566 & x_1447;
assign x_1449 = x_569 & x_570;
assign x_1450 = x_571 & x_572;
assign x_1451 = x_1449 & x_1450;
assign x_1452 = x_1448 & x_1451;
assign x_1453 = x_574 & x_575;
assign x_1454 = x_573 & x_1453;
assign x_1455 = x_576 & x_577;
assign x_1456 = x_578 & x_579;
assign x_1457 = x_1455 & x_1456;
assign x_1458 = x_1454 & x_1457;
assign x_1459 = x_1452 & x_1458;
assign x_1460 = x_1446 & x_1459;
assign x_1461 = x_581 & x_582;
assign x_1462 = x_580 & x_1461;
assign x_1463 = x_583 & x_584;
assign x_1464 = x_585 & x_586;
assign x_1465 = x_1463 & x_1464;
assign x_1466 = x_1462 & x_1465;
assign x_1467 = x_588 & x_589;
assign x_1468 = x_587 & x_1467;
assign x_1469 = x_590 & x_591;
assign x_1470 = x_592 & x_593;
assign x_1471 = x_1469 & x_1470;
assign x_1472 = x_1468 & x_1471;
assign x_1473 = x_1466 & x_1472;
assign x_1474 = x_595 & x_596;
assign x_1475 = x_594 & x_1474;
assign x_1476 = x_597 & x_598;
assign x_1477 = x_599 & x_600;
assign x_1478 = x_1476 & x_1477;
assign x_1479 = x_1475 & x_1478;
assign x_1480 = x_602 & x_603;
assign x_1481 = x_601 & x_1480;
assign x_1482 = x_604 & x_605;
assign x_1483 = x_606 & x_607;
assign x_1484 = x_1482 & x_1483;
assign x_1485 = x_1481 & x_1484;
assign x_1486 = x_1479 & x_1485;
assign x_1487 = x_1473 & x_1486;
assign x_1488 = x_1460 & x_1487;
assign x_1489 = x_609 & x_610;
assign x_1490 = x_608 & x_1489;
assign x_1491 = x_611 & x_612;
assign x_1492 = x_613 & x_614;
assign x_1493 = x_1491 & x_1492;
assign x_1494 = x_1490 & x_1493;
assign x_1495 = x_616 & x_617;
assign x_1496 = x_615 & x_1495;
assign x_1497 = x_618 & x_619;
assign x_1498 = x_620 & x_621;
assign x_1499 = x_1497 & x_1498;
assign x_1500 = x_1496 & x_1499;
assign x_1501 = x_1494 & x_1500;
assign x_1502 = x_623 & x_624;
assign x_1503 = x_622 & x_1502;
assign x_1504 = x_625 & x_626;
assign x_1505 = x_627 & x_628;
assign x_1506 = x_1504 & x_1505;
assign x_1507 = x_1503 & x_1506;
assign x_1508 = x_630 & x_631;
assign x_1509 = x_629 & x_1508;
assign x_1510 = x_632 & x_633;
assign x_1511 = x_634 & x_635;
assign x_1512 = x_1510 & x_1511;
assign x_1513 = x_1509 & x_1512;
assign x_1514 = x_1507 & x_1513;
assign x_1515 = x_1501 & x_1514;
assign x_1516 = x_637 & x_638;
assign x_1517 = x_636 & x_1516;
assign x_1518 = x_639 & x_640;
assign x_1519 = x_641 & x_642;
assign x_1520 = x_1518 & x_1519;
assign x_1521 = x_1517 & x_1520;
assign x_1522 = x_644 & x_645;
assign x_1523 = x_643 & x_1522;
assign x_1524 = x_646 & x_647;
assign x_1525 = x_648 & x_649;
assign x_1526 = x_1524 & x_1525;
assign x_1527 = x_1523 & x_1526;
assign x_1528 = x_1521 & x_1527;
assign x_1529 = x_651 & x_652;
assign x_1530 = x_650 & x_1529;
assign x_1531 = x_653 & x_654;
assign x_1532 = x_655 & x_656;
assign x_1533 = x_1531 & x_1532;
assign x_1534 = x_1530 & x_1533;
assign x_1535 = x_658 & x_659;
assign x_1536 = x_657 & x_1535;
assign x_1537 = x_660 & x_661;
assign x_1538 = x_662 & x_663;
assign x_1539 = x_1537 & x_1538;
assign x_1540 = x_1536 & x_1539;
assign x_1541 = x_1534 & x_1540;
assign x_1542 = x_1528 & x_1541;
assign x_1543 = x_1515 & x_1542;
assign x_1544 = x_1488 & x_1543;
assign x_1545 = x_1434 & x_1544;
assign x_1546 = x_665 & x_666;
assign x_1547 = x_664 & x_1546;
assign x_1548 = x_668 & x_669;
assign x_1549 = x_667 & x_1548;
assign x_1550 = x_1547 & x_1549;
assign x_1551 = x_671 & x_672;
assign x_1552 = x_670 & x_1551;
assign x_1553 = x_673 & x_674;
assign x_1554 = x_675 & x_676;
assign x_1555 = x_1553 & x_1554;
assign x_1556 = x_1552 & x_1555;
assign x_1557 = x_1550 & x_1556;
assign x_1558 = x_678 & x_679;
assign x_1559 = x_677 & x_1558;
assign x_1560 = x_680 & x_681;
assign x_1561 = x_682 & x_683;
assign x_1562 = x_1560 & x_1561;
assign x_1563 = x_1559 & x_1562;
assign x_1564 = x_685 & x_686;
assign x_1565 = x_684 & x_1564;
assign x_1566 = x_687 & x_688;
assign x_1567 = x_689 & x_690;
assign x_1568 = x_1566 & x_1567;
assign x_1569 = x_1565 & x_1568;
assign x_1570 = x_1563 & x_1569;
assign x_1571 = x_1557 & x_1570;
assign x_1572 = x_692 & x_693;
assign x_1573 = x_691 & x_1572;
assign x_1574 = x_694 & x_695;
assign x_1575 = x_696 & x_697;
assign x_1576 = x_1574 & x_1575;
assign x_1577 = x_1573 & x_1576;
assign x_1578 = x_699 & x_700;
assign x_1579 = x_698 & x_1578;
assign x_1580 = x_701 & x_702;
assign x_1581 = x_703 & x_704;
assign x_1582 = x_1580 & x_1581;
assign x_1583 = x_1579 & x_1582;
assign x_1584 = x_1577 & x_1583;
assign x_1585 = x_706 & x_707;
assign x_1586 = x_705 & x_1585;
assign x_1587 = x_708 & x_709;
assign x_1588 = x_710 & x_711;
assign x_1589 = x_1587 & x_1588;
assign x_1590 = x_1586 & x_1589;
assign x_1591 = x_713 & x_714;
assign x_1592 = x_712 & x_1591;
assign x_1593 = x_715 & x_716;
assign x_1594 = x_717 & x_718;
assign x_1595 = x_1593 & x_1594;
assign x_1596 = x_1592 & x_1595;
assign x_1597 = x_1590 & x_1596;
assign x_1598 = x_1584 & x_1597;
assign x_1599 = x_1571 & x_1598;
assign x_1600 = x_720 & x_721;
assign x_1601 = x_719 & x_1600;
assign x_1602 = x_723 & x_724;
assign x_1603 = x_722 & x_1602;
assign x_1604 = x_1601 & x_1603;
assign x_1605 = x_726 & x_727;
assign x_1606 = x_725 & x_1605;
assign x_1607 = x_728 & x_729;
assign x_1608 = x_730 & x_731;
assign x_1609 = x_1607 & x_1608;
assign x_1610 = x_1606 & x_1609;
assign x_1611 = x_1604 & x_1610;
assign x_1612 = x_733 & x_734;
assign x_1613 = x_732 & x_1612;
assign x_1614 = x_735 & x_736;
assign x_1615 = x_737 & x_738;
assign x_1616 = x_1614 & x_1615;
assign x_1617 = x_1613 & x_1616;
assign x_1618 = x_740 & x_741;
assign x_1619 = x_739 & x_1618;
assign x_1620 = x_742 & x_743;
assign x_1621 = x_744 & x_745;
assign x_1622 = x_1620 & x_1621;
assign x_1623 = x_1619 & x_1622;
assign x_1624 = x_1617 & x_1623;
assign x_1625 = x_1611 & x_1624;
assign x_1626 = x_747 & x_748;
assign x_1627 = x_746 & x_1626;
assign x_1628 = x_749 & x_750;
assign x_1629 = x_751 & x_752;
assign x_1630 = x_1628 & x_1629;
assign x_1631 = x_1627 & x_1630;
assign x_1632 = x_754 & x_755;
assign x_1633 = x_753 & x_1632;
assign x_1634 = x_756 & x_757;
assign x_1635 = x_758 & x_759;
assign x_1636 = x_1634 & x_1635;
assign x_1637 = x_1633 & x_1636;
assign x_1638 = x_1631 & x_1637;
assign x_1639 = x_761 & x_762;
assign x_1640 = x_760 & x_1639;
assign x_1641 = x_763 & x_764;
assign x_1642 = x_765 & x_766;
assign x_1643 = x_1641 & x_1642;
assign x_1644 = x_1640 & x_1643;
assign x_1645 = x_768 & x_769;
assign x_1646 = x_767 & x_1645;
assign x_1647 = x_770 & x_771;
assign x_1648 = x_772 & x_773;
assign x_1649 = x_1647 & x_1648;
assign x_1650 = x_1646 & x_1649;
assign x_1651 = x_1644 & x_1650;
assign x_1652 = x_1638 & x_1651;
assign x_1653 = x_1625 & x_1652;
assign x_1654 = x_1599 & x_1653;
assign x_1655 = x_775 & x_776;
assign x_1656 = x_774 & x_1655;
assign x_1657 = x_778 & x_779;
assign x_1658 = x_777 & x_1657;
assign x_1659 = x_1656 & x_1658;
assign x_1660 = x_781 & x_782;
assign x_1661 = x_780 & x_1660;
assign x_1662 = x_783 & x_784;
assign x_1663 = x_785 & x_786;
assign x_1664 = x_1662 & x_1663;
assign x_1665 = x_1661 & x_1664;
assign x_1666 = x_1659 & x_1665;
assign x_1667 = x_788 & x_789;
assign x_1668 = x_787 & x_1667;
assign x_1669 = x_790 & x_791;
assign x_1670 = x_792 & x_793;
assign x_1671 = x_1669 & x_1670;
assign x_1672 = x_1668 & x_1671;
assign x_1673 = x_795 & x_796;
assign x_1674 = x_794 & x_1673;
assign x_1675 = x_797 & x_798;
assign x_1676 = x_799 & x_800;
assign x_1677 = x_1675 & x_1676;
assign x_1678 = x_1674 & x_1677;
assign x_1679 = x_1672 & x_1678;
assign x_1680 = x_1666 & x_1679;
assign x_1681 = x_802 & x_803;
assign x_1682 = x_801 & x_1681;
assign x_1683 = x_804 & x_805;
assign x_1684 = x_806 & x_807;
assign x_1685 = x_1683 & x_1684;
assign x_1686 = x_1682 & x_1685;
assign x_1687 = x_809 & x_810;
assign x_1688 = x_808 & x_1687;
assign x_1689 = x_811 & x_812;
assign x_1690 = x_813 & x_814;
assign x_1691 = x_1689 & x_1690;
assign x_1692 = x_1688 & x_1691;
assign x_1693 = x_1686 & x_1692;
assign x_1694 = x_816 & x_817;
assign x_1695 = x_815 & x_1694;
assign x_1696 = x_818 & x_819;
assign x_1697 = x_820 & x_821;
assign x_1698 = x_1696 & x_1697;
assign x_1699 = x_1695 & x_1698;
assign x_1700 = x_823 & x_824;
assign x_1701 = x_822 & x_1700;
assign x_1702 = x_825 & x_826;
assign x_1703 = x_827 & x_828;
assign x_1704 = x_1702 & x_1703;
assign x_1705 = x_1701 & x_1704;
assign x_1706 = x_1699 & x_1705;
assign x_1707 = x_1693 & x_1706;
assign x_1708 = x_1680 & x_1707;
assign x_1709 = x_830 & x_831;
assign x_1710 = x_829 & x_1709;
assign x_1711 = x_832 & x_833;
assign x_1712 = x_834 & x_835;
assign x_1713 = x_1711 & x_1712;
assign x_1714 = x_1710 & x_1713;
assign x_1715 = x_837 & x_838;
assign x_1716 = x_836 & x_1715;
assign x_1717 = x_839 & x_840;
assign x_1718 = x_841 & x_842;
assign x_1719 = x_1717 & x_1718;
assign x_1720 = x_1716 & x_1719;
assign x_1721 = x_1714 & x_1720;
assign x_1722 = x_844 & x_845;
assign x_1723 = x_843 & x_1722;
assign x_1724 = x_846 & x_847;
assign x_1725 = x_848 & x_849;
assign x_1726 = x_1724 & x_1725;
assign x_1727 = x_1723 & x_1726;
assign x_1728 = x_851 & x_852;
assign x_1729 = x_850 & x_1728;
assign x_1730 = x_853 & x_854;
assign x_1731 = x_855 & x_856;
assign x_1732 = x_1730 & x_1731;
assign x_1733 = x_1729 & x_1732;
assign x_1734 = x_1727 & x_1733;
assign x_1735 = x_1721 & x_1734;
assign x_1736 = x_858 & x_859;
assign x_1737 = x_857 & x_1736;
assign x_1738 = x_860 & x_861;
assign x_1739 = x_862 & x_863;
assign x_1740 = x_1738 & x_1739;
assign x_1741 = x_1737 & x_1740;
assign x_1742 = x_865 & x_866;
assign x_1743 = x_864 & x_1742;
assign x_1744 = x_867 & x_868;
assign x_1745 = x_869 & x_870;
assign x_1746 = x_1744 & x_1745;
assign x_1747 = x_1743 & x_1746;
assign x_1748 = x_1741 & x_1747;
assign x_1749 = x_872 & x_873;
assign x_1750 = x_871 & x_1749;
assign x_1751 = x_874 & x_875;
assign x_1752 = x_876 & x_877;
assign x_1753 = x_1751 & x_1752;
assign x_1754 = x_1750 & x_1753;
assign x_1755 = x_879 & x_880;
assign x_1756 = x_878 & x_1755;
assign x_1757 = x_881 & x_882;
assign x_1758 = x_883 & x_884;
assign x_1759 = x_1757 & x_1758;
assign x_1760 = x_1756 & x_1759;
assign x_1761 = x_1754 & x_1760;
assign x_1762 = x_1748 & x_1761;
assign x_1763 = x_1735 & x_1762;
assign x_1764 = x_1708 & x_1763;
assign x_1765 = x_1654 & x_1764;
assign x_1766 = x_1545 & x_1765;
assign x_1767 = x_1325 & x_1766;
assign o_1 = x_1767;
endmodule
