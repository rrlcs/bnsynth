module formula(v_1,v_2,v_3,v_4,v_5,v_6,v_7,v_8,v_9,v_10,v_11,v_12,v_13,v_14,v_15,v_16,v_17,v_18,v_19,v_20,v_21,v_22,v_23,v_24,v_25,o_1);
	input v_1;
	input v_2;
	input v_3;
	input v_4;
	input v_5;
	input v_6;
	input v_7;
	input v_8;
	input v_9;
	input v_10;
	input v_11;
	input v_12;
	input v_13;
	input v_14;
	input v_15;
	input v_16;
	input v_17;
	input v_18;
	input v_19;
	input v_20;
	input v_21;
	input v_22;
	input v_23;
	input v_24;
	input v_25;
	wire v_26;
	wire v_27;
	wire v_28;
	wire v_29;
	wire v_30;
	wire v_31;
	wire v_32;
	wire v_33;
	wire v_34;
	wire v_35;
	wire v_36;
	wire v_37;
	wire v_38;
	wire v_39;
	wire v_40;
	wire v_41;
	wire v_42;
	wire v_43;
	wire v_44;
	wire v_45;
	wire v_46;
	wire v_47;
	wire v_48;
	wire v_49;
	wire v_50;
	wire v_51;
	wire v_52;
	wire v_53;
	wire v_54;
	wire v_55;
	wire v_56;
	wire v_57;
	wire v_58;
	wire v_59;
	wire v_60;
	wire v_61;
	wire v_62;
	wire v_63;
	wire v_64;
	wire v_65;
	wire v_66;
	wire v_67;
	wire v_68;
	wire v_69;
	wire v_70;
	wire v_71;
	wire v_72;
	wire v_73;
	wire x_1;
	output o_1;
	assign v_51 = (~v_17 & v_22) ;
	assign v_47 = (~v_16 & v_19) ;
	assign v_43 = (~v_15 & v_21) ;
	assign v_38 = (~v_4 & v_11) ;
	assign v_34 = (~v_3 & v_9) ;
	assign v_30 = (~v_2 & v_6) ;
	assign v_26 = (~v_1 & v_8) ;
	assign v_52 = (~v_25 & v_51) ;
	assign v_48 = (~v_23 & v_47) ;
	assign v_44 = (~v_20 & v_43) ;
	assign v_39 = (~v_14 & v_38) ;
	assign v_35 = (~v_12 & v_34) ;
	assign v_31 = (~v_10 & v_30) ;
	assign v_27 = (~v_7 & v_26) ;
	assign v_53 = (v_25 | v_52) ;
	assign v_49 = (v_23 | v_48) ;
	assign v_45 = (v_20 | v_44) ;
	assign v_40 = (v_14 | v_39) ;
	assign v_36 = (v_12 | v_35) ;
	assign v_32 = (v_10 | v_31) ;
	assign v_28 = (v_7 | v_27) ;
	assign v_66 = (v_24 ^ v_13) ;
	assign v_65 = (v_18 ^ v_5) ;
	assign v_63 = (v_22 ^ v_13) ;
	assign v_62 = (v_17 ^ v_5) ;
	assign v_60 = (v_19 ^ v_13) ;
	assign v_59 = (v_16 ^ v_5) ;
	assign v_57 = (v_21 ^ v_13) ;
	assign v_56 = (v_15 ^ v_5) ;
	assign v_54 = (v_53 ^ v_24) ;
	assign v_50 = (v_49 ^ v_22) ;
	assign v_46 = (v_45 ^ v_19) ;
	assign v_41 = (v_40 ^ v_13) ;
	assign v_37 = (v_36 ^ v_11) ;
	assign v_33 = (v_32 ^ v_9) ;
	assign v_29 = (v_28 ^ v_6) ;
	assign v_67 = (~v_65 & ~v_66) ;
	assign v_64 = (~v_62 & ~v_63) ;
	assign v_61 = (~v_59 & ~v_60) ;
	assign v_58 = (~v_56 & ~v_57) ;
	assign v_73 = (~v_50 & ~v_54) ;
	assign v_72 = ((((~v_15 & ~v_16) & ~v_17) & ~v_18) & ~v_46) ;
	assign v_71 = (((~v_29 & ~v_33) & ~v_37) & ~v_41) ;
	assign v_70 = ((((~v_1 & ~v_2) & ~v_3) & ~v_4) & ~v_5) ;
	assign v_68 = (((v_58 | v_61) | v_64) | v_67) ;
	assign v_55 = (v_72 & v_73) ;
	assign v_42 = (v_70 & v_71) ;
	assign v_69 = (v_55 & v_68) ;
	assign x_1 = (v_69 | ~v_42) ;
	assign o_1 = x_1 ;
endmodule
