module formula(v_1,v_2,v_3,v_4,v_5,v_6,v_7,v_8,v_9,v_10,v_11,v_12,v_13,v_15,v_16,v_17,v_18,v_19,v_20,v_21,v_22,v_23,v_24,v_25,v_26,v_27,v_28,v_29,v_30,v_31,v_32,v_33,v_34,v_35,v_36,v_37,v_38,v_39,v_40,v_41,v_42,v_43,v_44,v_45,v_46,v_47,v_48,v_49,v_53,v_54,v_55,v_56,v_57,v_58,v_62,v_66,v_67,v_68,v_69,v_70,v_71,v_72,v_73,v_80,v_81,v_82,v_14,v_50,v_51,v_52,v_59,v_60,v_61,v_63,v_64,v_65,v_74,v_75,v_76,v_77,v_78,v_79,v_83,v_84,v_85,v_86,v_87,v_88,v_89,v_90,v_91,v_92,v_93,v_94,v_95,v_96,v_97,v_98,v_99,v_100,v_101,v_102,v_103,v_104,v_105,v_106,v_107,v_108,v_109,v_110,v_111,v_112,v_113,v_114,v_115,v_116,v_117,v_118,v_119,v_120,v_121,v_122,v_123,v_124,v_125,v_126,v_127,v_128,v_129,v_130,v_131,v_132,v_133,v_134,v_135,v_136,v_137,v_138,v_139,v_140,v_141,v_142,v_143,v_144,v_145,v_146,v_147,v_148,v_149,v_150,v_151,v_152,v_153,v_154,v_155,v_156,v_157,v_158,v_159,v_160,v_161,v_162,v_163,v_164,v_165,v_166,v_167,v_168,v_169,v_170,v_171,v_172,v_173,v_174,v_175,v_176,v_177,v_178,v_179,v_180,v_181,v_182,v_183,v_184,v_185,v_186,v_187,v_188,v_189,v_190,v_191,v_192,v_193,v_194,v_195,v_196,v_197,v_198,v_199,v_200,v_201,v_202,v_203,v_204,v_205,v_206,v_207,v_208,v_209,v_210,v_211,v_212,v_213,v_214,v_215,v_216,v_217,v_218,v_219,v_220,v_221,v_222,v_223,v_224,v_225,v_226,v_227,v_228,v_229,v_230,v_231,v_232,v_233,v_234,v_235,v_236,v_237,v_238,v_239,v_240,v_241,v_242,v_243,v_244,v_245,v_246,v_247,v_248,v_249,v_250,v_251,v_252,v_253,v_254,v_255,v_256,v_257,v_258,v_259,v_260,v_261,v_262,v_263,v_264,v_265,v_266,v_267,v_268,v_269,v_270,v_271,v_272,v_273,v_274,v_275,v_276,v_277,v_278,v_279,v_280,v_281,v_282,v_283,v_284,v_285,v_286,v_287,v_288,v_289,v_290,v_291,v_292,v_293,v_294,v_295,v_296,v_297,v_298,v_299,v_300,v_301,v_302,v_303,v_304,v_305,v_306,v_307,v_308,v_309,v_310,v_311,v_312,v_313,v_314,v_315,v_316,v_317,v_318,v_319,v_320,v_321,v_322,v_323,v_324,v_325,v_326,v_327,v_328,v_329,v_330,v_331,v_332,v_333,v_334,v_335,v_336,v_337,v_338,v_339,v_340,v_341,v_342,v_343,v_344,v_345,v_346,v_347,v_348,v_349,v_350,v_351,v_352,v_353,v_354,v_355,v_356,v_357,v_358,v_359,v_360,v_361,v_362,v_363,v_364,v_365,v_366,v_367,v_368,v_369,v_370,v_371,v_372,v_373,v_374,v_375,v_376,v_377,v_378,v_379,v_380,v_381,v_382,v_383,v_384,v_385,v_386,v_387,v_388,v_389,v_390,v_391,v_392,v_393,v_394,v_395,v_396,v_397,v_398,v_399,v_400,v_401,v_402,v_403,v_404,v_405,v_406,v_407,v_408,v_409,v_410,v_411,v_412,v_413,v_414,v_415,v_416,v_417,v_418,v_419,v_420,v_421,v_422,v_423,v_424,v_425,v_426,v_427,v_428,v_429,v_430,v_431,v_432,v_433,v_434,v_435,v_436,v_437,v_438,v_439,v_440,v_441,v_442,v_443,v_444,v_445,v_446,v_447,v_448,v_449,v_450,v_451,v_452,v_453,v_454,v_455,v_456,v_457,v_458,v_459,v_460,v_461,v_462,v_463,v_464,v_465,v_466,v_467,v_468,v_469,v_470,v_471,v_472,v_473,v_475,v_476,v_477,v_478,v_479,v_480,v_481,v_482,v_483,v_484,v_485,v_486,v_487,v_488,v_489,v_490,v_491,v_492,v_493,v_494,v_495,v_496,v_497,v_498,v_499,v_500,v_501,v_502,v_503,v_504,v_505,v_506,v_507,v_508,v_509,v_510,v_511,v_512,v_513,v_514,v_515,v_516,v_517,v_518,v_519,v_520,v_521,v_522,v_523,v_524,v_525,v_526,v_527,v_528,v_529,v_530,v_531,v_532,v_533,v_534,v_535,v_536,v_537,v_538,v_539,v_540,v_541,v_542,v_543,v_544,v_545,v_546,v_547,v_548,v_549,v_550,v_551,v_552,v_553,v_554,v_555,v_556,v_557,v_558,v_559,v_560,v_561,v_562,v_563,v_564,v_565,v_566,v_567,v_568,v_569,v_570,v_571,v_572,v_573,v_574,v_575,v_576,v_577,v_578,v_579,v_580,v_581,v_582,v_583,v_584,v_585,v_586,v_587,v_588,v_589,v_590,v_591,v_592,v_593,v_594,v_595,v_596,v_597,v_598,v_599,v_600,v_601,v_602,v_603,v_604,v_605,v_606,v_607,v_608,v_609,v_610,v_611,v_612,v_613,v_614,v_615,v_616,v_617,v_618,v_619,v_620,v_621,v_622,v_623,v_624,v_625,v_626,v_627,v_628,v_629,v_630,v_631,v_632,v_633,v_634,v_635,v_636,v_637,v_638,v_639,v_640,v_641,v_642,v_643,v_644,v_645,v_646,v_647,v_648,v_649,v_650,v_651,v_652,v_653,v_654,v_655,v_656,v_657,v_658,v_659,v_660,v_661,v_662,v_663,v_664,v_665,v_666,v_667,v_668,v_669,v_670,v_671,v_672,v_673,v_674,v_675,v_676,v_677,v_678,v_679,v_680,v_681,v_682,v_683,v_684,v_685,v_686,v_687,v_688,v_689,v_690,v_691,v_692,v_693,v_694,v_695,v_696,v_697,v_698,v_699,v_700,v_701,v_702,v_703,v_704,v_705,v_706,v_707,v_708,v_709,v_710,v_711,v_712,v_713,v_714,v_715,v_716,v_717,v_718,v_719,v_720,v_721,v_722,v_723,v_724,v_725,v_726,v_727,v_728,v_729,v_730,v_731,v_732,v_733,v_734,v_735,v_736,v_737,v_738,v_739,v_740,v_741,v_742,v_743,v_744,v_745,v_746,v_747,v_748,v_749,v_750,v_751,v_752,v_753,v_754,v_755,v_756,v_757,v_758,v_759,v_760,v_761,v_762,v_763,v_764,v_765,v_766,v_767,v_768,v_769,v_770,v_771,v_772,v_773,v_774,v_775,v_776,v_777,v_778,v_779,v_780,v_781,v_782,v_783,v_784,v_785,v_786,v_787,v_788,v_789,v_790,v_791,v_792,v_793,v_794,v_795,v_796,v_797,v_798,v_799,v_800,v_801,v_802,v_803,v_804,v_805,v_806,v_807,v_808,v_809,v_810,v_811,v_812,v_813,v_814,v_815,v_816,v_817,v_818,v_819,v_820,v_821,v_822,v_823,v_824,v_825,v_826,v_827,v_828,v_829,v_830,v_831,v_832,v_833,v_834,v_835,v_836,v_837,v_838,v_839,v_840,v_841,v_842,v_843,v_844,v_845,v_846,v_847,v_848,v_849,v_850,v_851,v_852,v_853,v_854,v_855,v_856,v_857,v_858,v_859,v_860,v_861,v_862,v_863,v_864,v_865,o_1);
	input v_1;
	input v_2;
	input v_3;
	input v_4;
	input v_5;
	input v_6;
	input v_7;
	input v_8;
	input v_9;
	input v_10;
	input v_11;
	input v_12;
	input v_13;
	input v_15;
	input v_16;
	input v_17;
	input v_18;
	input v_19;
	input v_20;
	input v_21;
	input v_22;
	input v_23;
	input v_24;
	input v_25;
	input v_26;
	input v_27;
	input v_28;
	input v_29;
	input v_30;
	input v_31;
	input v_32;
	input v_33;
	input v_34;
	input v_35;
	input v_36;
	input v_37;
	input v_38;
	input v_39;
	input v_40;
	input v_41;
	input v_42;
	input v_43;
	input v_44;
	input v_45;
	input v_46;
	input v_47;
	input v_48;
	input v_49;
	input v_53;
	input v_54;
	input v_55;
	input v_56;
	input v_57;
	input v_58;
	input v_62;
	input v_66;
	input v_67;
	input v_68;
	input v_69;
	input v_70;
	input v_71;
	input v_72;
	input v_73;
	input v_80;
	input v_81;
	input v_82;
	input v_14;
	input v_50;
	input v_51;
	input v_52;
	input v_59;
	input v_60;
	input v_61;
	input v_63;
	input v_64;
	input v_65;
	input v_74;
	input v_75;
	input v_76;
	input v_77;
	input v_78;
	input v_79;
	input v_83;
	input v_84;
	input v_85;
	input v_86;
	input v_87;
	input v_88;
	input v_89;
	input v_90;
	input v_91;
	input v_92;
	input v_93;
	input v_94;
	input v_95;
	input v_96;
	input v_97;
	input v_98;
	input v_99;
	input v_100;
	input v_101;
	input v_102;
	input v_103;
	input v_104;
	input v_105;
	input v_106;
	input v_107;
	input v_108;
	input v_109;
	input v_110;
	input v_111;
	input v_112;
	input v_113;
	input v_114;
	input v_115;
	input v_116;
	input v_117;
	input v_118;
	input v_119;
	input v_120;
	input v_121;
	input v_122;
	input v_123;
	input v_124;
	input v_125;
	input v_126;
	input v_127;
	input v_128;
	input v_129;
	input v_130;
	input v_131;
	input v_132;
	input v_133;
	input v_134;
	input v_135;
	input v_136;
	input v_137;
	input v_138;
	input v_139;
	input v_140;
	input v_141;
	input v_142;
	input v_143;
	input v_144;
	input v_145;
	input v_146;
	input v_147;
	input v_148;
	input v_149;
	input v_150;
	input v_151;
	input v_152;
	input v_153;
	input v_154;
	input v_155;
	input v_156;
	input v_157;
	input v_158;
	input v_159;
	input v_160;
	input v_161;
	input v_162;
	input v_163;
	input v_164;
	input v_165;
	input v_166;
	input v_167;
	input v_168;
	input v_169;
	input v_170;
	input v_171;
	input v_172;
	input v_173;
	input v_174;
	input v_175;
	input v_176;
	input v_177;
	input v_178;
	input v_179;
	input v_180;
	input v_181;
	input v_182;
	input v_183;
	input v_184;
	input v_185;
	input v_186;
	input v_187;
	input v_188;
	input v_189;
	input v_190;
	input v_191;
	input v_192;
	input v_193;
	input v_194;
	input v_195;
	input v_196;
	input v_197;
	input v_198;
	input v_199;
	input v_200;
	input v_201;
	input v_202;
	input v_203;
	input v_204;
	input v_205;
	input v_206;
	input v_207;
	input v_208;
	input v_209;
	input v_210;
	input v_211;
	input v_212;
	input v_213;
	input v_214;
	input v_215;
	input v_216;
	input v_217;
	input v_218;
	input v_219;
	input v_220;
	input v_221;
	input v_222;
	input v_223;
	input v_224;
	input v_225;
	input v_226;
	input v_227;
	input v_228;
	input v_229;
	input v_230;
	input v_231;
	input v_232;
	input v_233;
	input v_234;
	input v_235;
	input v_236;
	input v_237;
	input v_238;
	input v_239;
	input v_240;
	input v_241;
	input v_242;
	input v_243;
	input v_244;
	input v_245;
	input v_246;
	input v_247;
	input v_248;
	input v_249;
	input v_250;
	input v_251;
	input v_252;
	input v_253;
	input v_254;
	input v_255;
	input v_256;
	input v_257;
	input v_258;
	input v_259;
	input v_260;
	input v_261;
	input v_262;
	input v_263;
	input v_264;
	input v_265;
	input v_266;
	input v_267;
	input v_268;
	input v_269;
	input v_270;
	input v_271;
	input v_272;
	input v_273;
	input v_274;
	input v_275;
	input v_276;
	input v_277;
	input v_278;
	input v_279;
	input v_280;
	input v_281;
	input v_282;
	input v_283;
	input v_284;
	input v_285;
	input v_286;
	input v_287;
	input v_288;
	input v_289;
	input v_290;
	input v_291;
	input v_292;
	input v_293;
	input v_294;
	input v_295;
	input v_296;
	input v_297;
	input v_298;
	input v_299;
	input v_300;
	input v_301;
	input v_302;
	input v_303;
	input v_304;
	input v_305;
	input v_306;
	input v_307;
	input v_308;
	input v_309;
	input v_310;
	input v_311;
	input v_312;
	input v_313;
	input v_314;
	input v_315;
	input v_316;
	input v_317;
	input v_318;
	input v_319;
	input v_320;
	input v_321;
	input v_322;
	input v_323;
	input v_324;
	input v_325;
	input v_326;
	input v_327;
	input v_328;
	input v_329;
	input v_330;
	input v_331;
	input v_332;
	input v_333;
	input v_334;
	input v_335;
	input v_336;
	input v_337;
	input v_338;
	input v_339;
	input v_340;
	input v_341;
	input v_342;
	input v_343;
	input v_344;
	input v_345;
	input v_346;
	input v_347;
	input v_348;
	input v_349;
	input v_350;
	input v_351;
	input v_352;
	input v_353;
	input v_354;
	input v_355;
	input v_356;
	input v_357;
	input v_358;
	input v_359;
	input v_360;
	input v_361;
	input v_362;
	input v_363;
	input v_364;
	input v_365;
	input v_366;
	input v_367;
	input v_368;
	input v_369;
	input v_370;
	input v_371;
	input v_372;
	input v_373;
	input v_374;
	input v_375;
	input v_376;
	input v_377;
	input v_378;
	input v_379;
	input v_380;
	input v_381;
	input v_382;
	input v_383;
	input v_384;
	input v_385;
	input v_386;
	input v_387;
	input v_388;
	input v_389;
	input v_390;
	input v_391;
	input v_392;
	input v_393;
	input v_394;
	input v_395;
	input v_396;
	input v_397;
	input v_398;
	input v_399;
	input v_400;
	input v_401;
	input v_402;
	input v_403;
	input v_404;
	input v_405;
	input v_406;
	input v_407;
	input v_408;
	input v_409;
	input v_410;
	input v_411;
	input v_412;
	input v_413;
	input v_414;
	input v_415;
	input v_416;
	input v_417;
	input v_418;
	input v_419;
	input v_420;
	input v_421;
	input v_422;
	input v_423;
	input v_424;
	input v_425;
	input v_426;
	input v_427;
	input v_428;
	input v_429;
	input v_430;
	input v_431;
	input v_432;
	input v_433;
	input v_434;
	input v_435;
	input v_436;
	input v_437;
	input v_438;
	input v_439;
	input v_440;
	input v_441;
	input v_442;
	input v_443;
	input v_444;
	input v_445;
	input v_446;
	input v_447;
	input v_448;
	input v_449;
	input v_450;
	input v_451;
	input v_452;
	input v_453;
	input v_454;
	input v_455;
	input v_456;
	input v_457;
	input v_458;
	input v_459;
	input v_460;
	input v_461;
	input v_462;
	input v_463;
	input v_464;
	input v_465;
	input v_466;
	input v_467;
	input v_468;
	input v_469;
	input v_470;
	input v_471;
	input v_472;
	input v_473;
	input v_475;
	input v_476;
	input v_477;
	input v_478;
	input v_479;
	input v_480;
	input v_481;
	input v_482;
	input v_483;
	input v_484;
	input v_485;
	input v_486;
	input v_487;
	input v_488;
	input v_489;
	input v_490;
	input v_491;
	input v_492;
	input v_493;
	input v_494;
	input v_495;
	input v_496;
	input v_497;
	input v_498;
	input v_499;
	input v_500;
	input v_501;
	input v_502;
	input v_503;
	input v_504;
	input v_505;
	input v_506;
	input v_507;
	input v_508;
	input v_509;
	input v_510;
	input v_511;
	input v_512;
	input v_513;
	input v_514;
	input v_515;
	input v_516;
	input v_517;
	input v_518;
	input v_519;
	input v_520;
	input v_521;
	input v_522;
	input v_523;
	input v_524;
	input v_525;
	input v_526;
	input v_527;
	input v_528;
	input v_529;
	input v_530;
	input v_531;
	input v_532;
	input v_533;
	input v_534;
	input v_535;
	input v_536;
	input v_537;
	input v_538;
	input v_539;
	input v_540;
	input v_541;
	input v_542;
	input v_543;
	input v_544;
	input v_545;
	input v_546;
	input v_547;
	input v_548;
	input v_549;
	input v_550;
	input v_551;
	input v_552;
	input v_553;
	input v_554;
	input v_555;
	input v_556;
	input v_557;
	input v_558;
	input v_559;
	input v_560;
	input v_561;
	input v_562;
	input v_563;
	input v_564;
	input v_565;
	input v_566;
	input v_567;
	input v_568;
	input v_569;
	input v_570;
	input v_571;
	input v_572;
	input v_573;
	input v_574;
	input v_575;
	input v_576;
	input v_577;
	input v_578;
	input v_579;
	input v_580;
	input v_581;
	input v_582;
	input v_583;
	input v_584;
	input v_585;
	input v_586;
	input v_587;
	input v_588;
	input v_589;
	input v_590;
	input v_591;
	input v_592;
	input v_593;
	input v_594;
	input v_595;
	input v_596;
	input v_597;
	input v_598;
	input v_599;
	input v_600;
	input v_601;
	input v_602;
	input v_603;
	input v_604;
	input v_605;
	input v_606;
	input v_607;
	input v_608;
	input v_609;
	input v_610;
	input v_611;
	input v_612;
	input v_613;
	input v_614;
	input v_615;
	input v_616;
	input v_617;
	input v_618;
	input v_619;
	input v_620;
	input v_621;
	input v_622;
	input v_623;
	input v_624;
	input v_625;
	input v_626;
	input v_627;
	input v_628;
	input v_629;
	input v_630;
	input v_631;
	input v_632;
	input v_633;
	input v_634;
	input v_635;
	input v_636;
	input v_637;
	input v_638;
	input v_639;
	input v_640;
	input v_641;
	input v_642;
	input v_643;
	input v_644;
	input v_645;
	input v_646;
	input v_647;
	input v_648;
	input v_649;
	input v_650;
	input v_651;
	input v_652;
	input v_653;
	input v_654;
	input v_655;
	input v_656;
	input v_657;
	input v_658;
	input v_659;
	input v_660;
	input v_661;
	input v_662;
	input v_663;
	input v_664;
	input v_665;
	input v_666;
	input v_667;
	input v_668;
	input v_669;
	input v_670;
	input v_671;
	input v_672;
	input v_673;
	input v_674;
	input v_675;
	input v_676;
	input v_677;
	input v_678;
	input v_679;
	input v_680;
	input v_681;
	input v_682;
	input v_683;
	input v_684;
	input v_685;
	input v_686;
	input v_687;
	input v_688;
	input v_689;
	input v_690;
	input v_691;
	input v_692;
	input v_693;
	input v_694;
	input v_695;
	input v_696;
	input v_697;
	input v_698;
	input v_699;
	input v_700;
	input v_701;
	input v_702;
	input v_703;
	input v_704;
	input v_705;
	input v_706;
	input v_707;
	input v_708;
	input v_709;
	input v_710;
	input v_711;
	input v_712;
	input v_713;
	input v_714;
	input v_715;
	input v_716;
	input v_717;
	input v_718;
	input v_719;
	input v_720;
	input v_721;
	input v_722;
	input v_723;
	input v_724;
	input v_725;
	input v_726;
	input v_727;
	input v_728;
	input v_729;
	input v_730;
	input v_731;
	input v_732;
	input v_733;
	input v_734;
	input v_735;
	input v_736;
	input v_737;
	input v_738;
	input v_739;
	input v_740;
	input v_741;
	input v_742;
	input v_743;
	input v_744;
	input v_745;
	input v_746;
	input v_747;
	input v_748;
	input v_749;
	input v_750;
	input v_751;
	input v_752;
	input v_753;
	input v_754;
	input v_755;
	input v_756;
	input v_757;
	input v_758;
	input v_759;
	input v_760;
	input v_761;
	input v_762;
	input v_763;
	input v_764;
	input v_765;
	input v_766;
	input v_767;
	input v_768;
	input v_769;
	input v_770;
	input v_771;
	input v_772;
	input v_773;
	input v_774;
	input v_775;
	input v_776;
	input v_777;
	input v_778;
	input v_779;
	input v_780;
	input v_781;
	input v_782;
	input v_783;
	input v_784;
	input v_785;
	input v_786;
	input v_787;
	input v_788;
	input v_789;
	input v_790;
	input v_791;
	input v_792;
	input v_793;
	input v_794;
	input v_795;
	input v_796;
	input v_797;
	input v_798;
	input v_799;
	input v_800;
	input v_801;
	input v_802;
	input v_803;
	input v_804;
	input v_805;
	input v_806;
	input v_807;
	input v_808;
	input v_809;
	input v_810;
	input v_811;
	input v_812;
	input v_813;
	input v_814;
	input v_815;
	input v_816;
	input v_817;
	input v_818;
	input v_819;
	input v_820;
	input v_821;
	input v_822;
	input v_823;
	input v_824;
	input v_825;
	input v_826;
	input v_827;
	input v_828;
	input v_829;
	input v_830;
	input v_831;
	input v_832;
	input v_833;
	input v_834;
	input v_835;
	input v_836;
	input v_837;
	input v_838;
	input v_839;
	input v_840;
	input v_841;
	input v_842;
	input v_843;
	input v_844;
	input v_845;
	input v_846;
	input v_847;
	input v_848;
	input v_849;
	input v_850;
	input v_851;
	input v_852;
	input v_853;
	input v_854;
	input v_855;
	input v_856;
	input v_857;
	input v_858;
	input v_859;
	input v_860;
	input v_861;
	input v_862;
	input v_863;
	input v_864;
	input v_865;
	wire v_474;
	wire v_866;
	wire v_867;
	wire x_1;
	wire x_2;
	wire x_3;
	wire x_4;
	wire x_5;
	wire x_6;
	wire x_7;
	wire x_8;
	wire x_9;
	wire x_10;
	wire x_11;
	wire x_12;
	wire x_13;
	wire x_14;
	wire x_15;
	wire x_16;
	wire x_17;
	wire x_18;
	wire x_19;
	wire x_20;
	wire x_21;
	wire x_22;
	wire x_23;
	wire x_24;
	wire x_25;
	wire x_26;
	wire x_27;
	wire x_28;
	wire x_29;
	wire x_30;
	wire x_31;
	wire x_32;
	wire x_33;
	wire x_34;
	wire x_35;
	wire x_36;
	wire x_37;
	wire x_38;
	wire x_39;
	wire x_40;
	wire x_41;
	wire x_42;
	wire x_43;
	wire x_44;
	wire x_45;
	wire x_46;
	wire x_47;
	wire x_48;
	wire x_49;
	wire x_50;
	wire x_51;
	wire x_52;
	wire x_53;
	wire x_54;
	wire x_55;
	wire x_56;
	wire x_57;
	wire x_58;
	wire x_59;
	wire x_60;
	wire x_61;
	wire x_62;
	wire x_63;
	wire x_64;
	wire x_65;
	wire x_66;
	wire x_67;
	wire x_68;
	wire x_69;
	wire x_70;
	wire x_71;
	wire x_72;
	wire x_73;
	wire x_74;
	wire x_75;
	wire x_76;
	wire x_77;
	wire x_78;
	wire x_79;
	wire x_80;
	wire x_81;
	wire x_82;
	wire x_83;
	wire x_84;
	wire x_85;
	wire x_86;
	wire x_87;
	wire x_88;
	wire x_89;
	wire x_90;
	wire x_91;
	wire x_92;
	wire x_93;
	wire x_94;
	wire x_95;
	wire x_96;
	wire x_97;
	wire x_98;
	wire x_99;
	wire x_100;
	wire x_101;
	wire x_102;
	wire x_103;
	wire x_104;
	wire x_105;
	wire x_106;
	wire x_107;
	wire x_108;
	wire x_109;
	wire x_110;
	wire x_111;
	wire x_112;
	wire x_113;
	wire x_114;
	wire x_115;
	wire x_116;
	wire x_117;
	wire x_118;
	wire x_119;
	wire x_120;
	wire x_121;
	wire x_122;
	wire x_123;
	wire x_124;
	wire x_125;
	wire x_126;
	wire x_127;
	wire x_128;
	wire x_129;
	wire x_130;
	wire x_131;
	wire x_132;
	wire x_133;
	wire x_134;
	wire x_135;
	wire x_136;
	wire x_137;
	wire x_138;
	wire x_139;
	wire x_140;
	wire x_141;
	wire x_142;
	wire x_143;
	wire x_144;
	wire x_145;
	wire x_146;
	wire x_147;
	wire x_148;
	wire x_149;
	wire x_150;
	wire x_151;
	wire x_152;
	wire x_153;
	wire x_154;
	wire x_155;
	wire x_156;
	wire x_157;
	wire x_158;
	wire x_159;
	wire x_160;
	wire x_161;
	wire x_162;
	wire x_163;
	wire x_164;
	wire x_165;
	wire x_166;
	wire x_167;
	wire x_168;
	wire x_169;
	wire x_170;
	wire x_171;
	wire x_172;
	wire x_173;
	wire x_174;
	wire x_175;
	wire x_176;
	wire x_177;
	wire x_178;
	wire x_179;
	wire x_180;
	wire x_181;
	wire x_182;
	wire x_183;
	wire x_184;
	wire x_185;
	wire x_186;
	wire x_187;
	wire x_188;
	wire x_189;
	wire x_190;
	wire x_191;
	wire x_192;
	wire x_193;
	wire x_194;
	wire x_195;
	wire x_196;
	wire x_197;
	wire x_198;
	wire x_199;
	wire x_200;
	wire x_201;
	wire x_202;
	wire x_203;
	wire x_204;
	wire x_205;
	wire x_206;
	wire x_207;
	wire x_208;
	wire x_209;
	wire x_210;
	wire x_211;
	wire x_212;
	wire x_213;
	wire x_214;
	wire x_215;
	wire x_216;
	wire x_217;
	wire x_218;
	wire x_219;
	wire x_220;
	wire x_221;
	wire x_222;
	wire x_223;
	wire x_224;
	wire x_225;
	wire x_226;
	wire x_227;
	wire x_228;
	wire x_229;
	wire x_230;
	wire x_231;
	wire x_232;
	wire x_233;
	wire x_234;
	wire x_235;
	wire x_236;
	wire x_237;
	wire x_238;
	wire x_239;
	wire x_240;
	wire x_241;
	wire x_242;
	wire x_243;
	wire x_244;
	wire x_245;
	wire x_246;
	wire x_247;
	wire x_248;
	wire x_249;
	wire x_250;
	wire x_251;
	wire x_252;
	wire x_253;
	wire x_254;
	wire x_255;
	wire x_256;
	wire x_257;
	wire x_258;
	wire x_259;
	wire x_260;
	wire x_261;
	wire x_262;
	wire x_263;
	wire x_264;
	wire x_265;
	wire x_266;
	wire x_267;
	wire x_268;
	wire x_269;
	wire x_270;
	wire x_271;
	wire x_272;
	wire x_273;
	wire x_274;
	wire x_275;
	wire x_276;
	wire x_277;
	wire x_278;
	wire x_279;
	wire x_280;
	wire x_281;
	wire x_282;
	wire x_283;
	wire x_284;
	wire x_285;
	wire x_286;
	wire x_287;
	wire x_288;
	wire x_289;
	wire x_290;
	wire x_291;
	wire x_292;
	wire x_293;
	wire x_294;
	wire x_295;
	wire x_296;
	wire x_297;
	wire x_298;
	wire x_299;
	wire x_300;
	wire x_301;
	wire x_302;
	wire x_303;
	wire x_304;
	wire x_305;
	wire x_306;
	wire x_307;
	wire x_308;
	wire x_309;
	wire x_310;
	wire x_311;
	wire x_312;
	wire x_313;
	wire x_314;
	wire x_315;
	wire x_316;
	wire x_317;
	wire x_318;
	wire x_319;
	wire x_320;
	wire x_321;
	wire x_322;
	wire x_323;
	wire x_324;
	wire x_325;
	wire x_326;
	wire x_327;
	wire x_328;
	wire x_329;
	wire x_330;
	wire x_331;
	wire x_332;
	wire x_333;
	wire x_334;
	wire x_335;
	wire x_336;
	wire x_337;
	wire x_338;
	wire x_339;
	wire x_340;
	wire x_341;
	wire x_342;
	wire x_343;
	wire x_344;
	wire x_345;
	wire x_346;
	wire x_347;
	wire x_348;
	wire x_349;
	wire x_350;
	wire x_351;
	wire x_352;
	wire x_353;
	wire x_354;
	wire x_355;
	wire x_356;
	wire x_357;
	wire x_358;
	wire x_359;
	wire x_360;
	wire x_361;
	wire x_362;
	wire x_363;
	wire x_364;
	wire x_365;
	wire x_366;
	wire x_367;
	wire x_368;
	wire x_369;
	wire x_370;
	wire x_371;
	wire x_372;
	wire x_373;
	wire x_374;
	wire x_375;
	wire x_376;
	wire x_377;
	wire x_378;
	wire x_379;
	wire x_380;
	wire x_381;
	wire x_382;
	wire x_383;
	wire x_384;
	wire x_385;
	wire x_386;
	wire x_387;
	wire x_388;
	wire x_389;
	wire x_390;
	wire x_391;
	wire x_392;
	wire x_393;
	wire x_394;
	wire x_395;
	wire x_396;
	wire x_397;
	wire x_398;
	wire x_399;
	wire x_400;
	wire x_401;
	wire x_402;
	wire x_403;
	wire x_404;
	wire x_405;
	wire x_406;
	wire x_407;
	wire x_408;
	wire x_409;
	wire x_410;
	wire x_411;
	wire x_412;
	wire x_413;
	wire x_414;
	wire x_415;
	wire x_416;
	wire x_417;
	wire x_418;
	wire x_419;
	wire x_420;
	wire x_421;
	wire x_422;
	wire x_423;
	wire x_424;
	wire x_425;
	wire x_426;
	wire x_427;
	wire x_428;
	wire x_429;
	wire x_430;
	wire x_431;
	wire x_432;
	wire x_433;
	wire x_434;
	wire x_435;
	wire x_436;
	wire x_437;
	wire x_438;
	wire x_439;
	wire x_440;
	wire x_441;
	wire x_442;
	wire x_443;
	wire x_444;
	wire x_445;
	wire x_446;
	wire x_447;
	wire x_448;
	wire x_449;
	wire x_450;
	wire x_451;
	wire x_452;
	wire x_453;
	wire x_454;
	wire x_455;
	wire x_456;
	wire x_457;
	wire x_458;
	wire x_459;
	wire x_460;
	wire x_461;
	wire x_462;
	wire x_463;
	wire x_464;
	wire x_465;
	wire x_466;
	wire x_467;
	wire x_468;
	wire x_469;
	wire x_470;
	wire x_471;
	wire x_472;
	wire x_473;
	wire x_474;
	wire x_475;
	wire x_476;
	wire x_477;
	wire x_478;
	wire x_479;
	wire x_480;
	wire x_481;
	wire x_482;
	wire x_483;
	wire x_484;
	wire x_485;
	wire x_486;
	wire x_487;
	wire x_488;
	wire x_489;
	wire x_490;
	wire x_491;
	wire x_492;
	wire x_493;
	wire x_494;
	wire x_495;
	wire x_496;
	wire x_497;
	wire x_498;
	wire x_499;
	wire x_500;
	wire x_501;
	wire x_502;
	wire x_503;
	wire x_504;
	wire x_505;
	wire x_506;
	wire x_507;
	wire x_508;
	wire x_509;
	wire x_510;
	wire x_511;
	wire x_512;
	wire x_513;
	wire x_514;
	wire x_515;
	wire x_516;
	wire x_517;
	wire x_518;
	wire x_519;
	wire x_520;
	wire x_521;
	wire x_522;
	wire x_523;
	wire x_524;
	wire x_525;
	wire x_526;
	wire x_527;
	wire x_528;
	wire x_529;
	wire x_530;
	wire x_531;
	wire x_532;
	wire x_533;
	wire x_534;
	wire x_535;
	wire x_536;
	wire x_537;
	wire x_538;
	wire x_539;
	wire x_540;
	wire x_541;
	wire x_542;
	wire x_543;
	wire x_544;
	wire x_545;
	wire x_546;
	wire x_547;
	wire x_548;
	wire x_549;
	wire x_550;
	wire x_551;
	wire x_552;
	wire x_553;
	wire x_554;
	wire x_555;
	wire x_556;
	wire x_557;
	wire x_558;
	wire x_559;
	wire x_560;
	wire x_561;
	wire x_562;
	wire x_563;
	wire x_564;
	wire x_565;
	wire x_566;
	wire x_567;
	wire x_568;
	wire x_569;
	wire x_570;
	wire x_571;
	wire x_572;
	wire x_573;
	wire x_574;
	wire x_575;
	wire x_576;
	wire x_577;
	wire x_578;
	wire x_579;
	wire x_580;
	wire x_581;
	wire x_582;
	wire x_583;
	wire x_584;
	wire x_585;
	wire x_586;
	wire x_587;
	wire x_588;
	wire x_589;
	wire x_590;
	wire x_591;
	wire x_592;
	wire x_593;
	wire x_594;
	wire x_595;
	wire x_596;
	wire x_597;
	wire x_598;
	wire x_599;
	wire x_600;
	wire x_601;
	wire x_602;
	wire x_603;
	wire x_604;
	wire x_605;
	wire x_606;
	wire x_607;
	wire x_608;
	wire x_609;
	wire x_610;
	wire x_611;
	wire x_612;
	wire x_613;
	wire x_614;
	wire x_615;
	wire x_616;
	wire x_617;
	wire x_618;
	wire x_619;
	wire x_620;
	wire x_621;
	wire x_622;
	wire x_623;
	wire x_624;
	wire x_625;
	wire x_626;
	wire x_627;
	wire x_628;
	wire x_629;
	wire x_630;
	wire x_631;
	wire x_632;
	wire x_633;
	wire x_634;
	wire x_635;
	wire x_636;
	wire x_637;
	wire x_638;
	wire x_639;
	wire x_640;
	wire x_641;
	wire x_642;
	wire x_643;
	wire x_644;
	wire x_645;
	wire x_646;
	wire x_647;
	wire x_648;
	wire x_649;
	wire x_650;
	wire x_651;
	wire x_652;
	wire x_653;
	wire x_654;
	wire x_655;
	wire x_656;
	wire x_657;
	wire x_658;
	wire x_659;
	wire x_660;
	wire x_661;
	wire x_662;
	wire x_663;
	wire x_664;
	wire x_665;
	wire x_666;
	wire x_667;
	wire x_668;
	wire x_669;
	wire x_670;
	wire x_671;
	wire x_672;
	wire x_673;
	wire x_674;
	wire x_675;
	wire x_676;
	wire x_677;
	wire x_678;
	wire x_679;
	wire x_680;
	wire x_681;
	wire x_682;
	wire x_683;
	wire x_684;
	wire x_685;
	wire x_686;
	wire x_687;
	wire x_688;
	wire x_689;
	wire x_690;
	wire x_691;
	wire x_692;
	wire x_693;
	wire x_694;
	wire x_695;
	wire x_696;
	wire x_697;
	wire x_698;
	wire x_699;
	wire x_700;
	wire x_701;
	wire x_702;
	wire x_703;
	wire x_704;
	wire x_705;
	wire x_706;
	wire x_707;
	wire x_708;
	wire x_709;
	wire x_710;
	wire x_711;
	wire x_712;
	wire x_713;
	wire x_714;
	wire x_715;
	wire x_716;
	wire x_717;
	wire x_718;
	wire x_719;
	wire x_720;
	wire x_721;
	wire x_722;
	wire x_723;
	wire x_724;
	wire x_725;
	wire x_726;
	wire x_727;
	wire x_728;
	wire x_729;
	wire x_730;
	wire x_731;
	wire x_732;
	wire x_733;
	wire x_734;
	wire x_735;
	wire x_736;
	wire x_737;
	wire x_738;
	wire x_739;
	wire x_740;
	wire x_741;
	wire x_742;
	wire x_743;
	wire x_744;
	wire x_745;
	wire x_746;
	wire x_747;
	wire x_748;
	wire x_749;
	wire x_750;
	wire x_751;
	wire x_752;
	wire x_753;
	wire x_754;
	wire x_755;
	wire x_756;
	wire x_757;
	wire x_758;
	wire x_759;
	wire x_760;
	wire x_761;
	wire x_762;
	wire x_763;
	wire x_764;
	wire x_765;
	wire x_766;
	wire x_767;
	wire x_768;
	wire x_769;
	wire x_770;
	wire x_771;
	wire x_772;
	wire x_773;
	wire x_774;
	wire x_775;
	wire x_776;
	wire x_777;
	wire x_778;
	wire x_779;
	wire x_780;
	wire x_781;
	wire x_782;
	wire x_783;
	wire x_784;
	wire x_785;
	wire x_786;
	wire x_787;
	wire x_788;
	wire x_789;
	wire x_790;
	wire x_791;
	wire x_792;
	wire x_793;
	wire x_794;
	wire x_795;
	wire x_796;
	wire x_797;
	wire x_798;
	wire x_799;
	wire x_800;
	wire x_801;
	wire x_802;
	wire x_803;
	wire x_804;
	wire x_805;
	wire x_806;
	wire x_807;
	wire x_808;
	wire x_809;
	wire x_810;
	wire x_811;
	wire x_812;
	wire x_813;
	wire x_814;
	wire x_815;
	wire x_816;
	wire x_817;
	wire x_818;
	wire x_819;
	wire x_820;
	wire x_821;
	wire x_822;
	wire x_823;
	wire x_824;
	wire x_825;
	wire x_826;
	wire x_827;
	wire x_828;
	wire x_829;
	wire x_830;
	wire x_831;
	wire x_832;
	wire x_833;
	wire x_834;
	wire x_835;
	wire x_836;
	wire x_837;
	wire x_838;
	wire x_839;
	wire x_840;
	wire x_841;
	wire x_842;
	wire x_843;
	wire x_844;
	wire x_845;
	wire x_846;
	wire x_847;
	wire x_848;
	wire x_849;
	wire x_850;
	wire x_851;
	wire x_852;
	wire x_853;
	wire x_854;
	wire x_855;
	wire x_856;
	wire x_857;
	wire x_858;
	wire x_859;
	wire x_860;
	wire x_861;
	wire x_862;
	wire x_863;
	wire x_864;
	wire x_865;
	wire x_866;
	wire x_867;
	wire x_868;
	wire x_869;
	wire x_870;
	wire x_871;
	wire x_872;
	wire x_873;
	wire x_874;
	wire x_875;
	wire x_876;
	wire x_877;
	wire x_878;
	wire x_879;
	wire x_880;
	wire x_881;
	wire x_882;
	wire x_883;
	wire x_884;
	wire x_885;
	wire x_886;
	wire x_887;
	wire x_888;
	wire x_889;
	wire x_890;
	wire x_891;
	wire x_892;
	wire x_893;
	wire x_894;
	wire x_895;
	wire x_896;
	wire x_897;
	wire x_898;
	wire x_899;
	wire x_900;
	wire x_901;
	wire x_902;
	wire x_903;
	wire x_904;
	wire x_905;
	wire x_906;
	wire x_907;
	wire x_908;
	wire x_909;
	wire x_910;
	wire x_911;
	wire x_912;
	wire x_913;
	wire x_914;
	wire x_915;
	wire x_916;
	wire x_917;
	wire x_918;
	wire x_919;
	wire x_920;
	wire x_921;
	wire x_922;
	wire x_923;
	wire x_924;
	wire x_925;
	wire x_926;
	wire x_927;
	wire x_928;
	wire x_929;
	wire x_930;
	wire x_931;
	wire x_932;
	wire x_933;
	wire x_934;
	wire x_935;
	wire x_936;
	wire x_937;
	wire x_938;
	wire x_939;
	wire x_940;
	wire x_941;
	wire x_942;
	wire x_943;
	wire x_944;
	wire x_945;
	wire x_946;
	wire x_947;
	wire x_948;
	wire x_949;
	wire x_950;
	wire x_951;
	wire x_952;
	wire x_953;
	wire x_954;
	wire x_955;
	wire x_956;
	wire x_957;
	wire x_958;
	wire x_959;
	wire x_960;
	wire x_961;
	wire x_962;
	wire x_963;
	wire x_964;
	wire x_965;
	wire x_966;
	wire x_967;
	wire x_968;
	wire x_969;
	wire x_970;
	wire x_971;
	wire x_972;
	wire x_973;
	wire x_974;
	wire x_975;
	wire x_976;
	wire x_977;
	wire x_978;
	wire x_979;
	wire x_980;
	wire x_981;
	wire x_982;
	wire x_983;
	wire x_984;
	wire x_985;
	wire x_986;
	wire x_987;
	wire x_988;
	wire x_989;
	wire x_990;
	wire x_991;
	wire x_992;
	wire x_993;
	wire x_994;
	wire x_995;
	wire x_996;
	wire x_997;
	wire x_998;
	wire x_999;
	wire x_1000;
	wire x_1001;
	wire x_1002;
	wire x_1003;
	wire x_1004;
	wire x_1005;
	wire x_1006;
	wire x_1007;
	wire x_1008;
	wire x_1009;
	wire x_1010;
	wire x_1011;
	wire x_1012;
	wire x_1013;
	wire x_1014;
	wire x_1015;
	wire x_1016;
	wire x_1017;
	wire x_1018;
	wire x_1019;
	wire x_1020;
	wire x_1021;
	wire x_1022;
	wire x_1023;
	wire x_1024;
	wire x_1025;
	wire x_1026;
	wire x_1027;
	wire x_1028;
	wire x_1029;
	wire x_1030;
	wire x_1031;
	wire x_1032;
	wire x_1033;
	wire x_1034;
	wire x_1035;
	wire x_1036;
	wire x_1037;
	wire x_1038;
	wire x_1039;
	wire x_1040;
	wire x_1041;
	wire x_1042;
	wire x_1043;
	wire x_1044;
	wire x_1045;
	wire x_1046;
	wire x_1047;
	wire x_1048;
	wire x_1049;
	wire x_1050;
	wire x_1051;
	wire x_1052;
	wire x_1053;
	wire x_1054;
	wire x_1055;
	wire x_1056;
	wire x_1057;
	wire x_1058;
	wire x_1059;
	wire x_1060;
	wire x_1061;
	wire x_1062;
	wire x_1063;
	wire x_1064;
	wire x_1065;
	wire x_1066;
	wire x_1067;
	wire x_1068;
	wire x_1069;
	wire x_1070;
	wire x_1071;
	wire x_1072;
	wire x_1073;
	wire x_1074;
	wire x_1075;
	wire x_1076;
	wire x_1077;
	wire x_1078;
	wire x_1079;
	wire x_1080;
	wire x_1081;
	wire x_1082;
	wire x_1083;
	wire x_1084;
	wire x_1085;
	wire x_1086;
	wire x_1087;
	wire x_1088;
	wire x_1089;
	wire x_1090;
	wire x_1091;
	wire x_1092;
	wire x_1093;
	wire x_1094;
	wire x_1095;
	wire x_1096;
	wire x_1097;
	wire x_1098;
	wire x_1099;
	wire x_1100;
	wire x_1101;
	wire x_1102;
	wire x_1103;
	wire x_1104;
	wire x_1105;
	wire x_1106;
	wire x_1107;
	wire x_1108;
	wire x_1109;
	wire x_1110;
	wire x_1111;
	wire x_1112;
	wire x_1113;
	wire x_1114;
	wire x_1115;
	wire x_1116;
	wire x_1117;
	wire x_1118;
	wire x_1119;
	wire x_1120;
	wire x_1121;
	wire x_1122;
	wire x_1123;
	wire x_1124;
	wire x_1125;
	wire x_1126;
	wire x_1127;
	wire x_1128;
	wire x_1129;
	wire x_1130;
	wire x_1131;
	wire x_1132;
	wire x_1133;
	wire x_1134;
	wire x_1135;
	wire x_1136;
	wire x_1137;
	wire x_1138;
	wire x_1139;
	wire x_1140;
	wire x_1141;
	wire x_1142;
	wire x_1143;
	wire x_1144;
	wire x_1145;
	wire x_1146;
	wire x_1147;
	wire x_1148;
	wire x_1149;
	wire x_1150;
	wire x_1151;
	wire x_1152;
	wire x_1153;
	wire x_1154;
	wire x_1155;
	wire x_1156;
	wire x_1157;
	wire x_1158;
	wire x_1159;
	wire x_1160;
	wire x_1161;
	wire x_1162;
	wire x_1163;
	wire x_1164;
	wire x_1165;
	wire x_1166;
	wire x_1167;
	wire x_1168;
	wire x_1169;
	wire x_1170;
	wire x_1171;
	wire x_1172;
	wire x_1173;
	wire x_1174;
	wire x_1175;
	wire x_1176;
	wire x_1177;
	wire x_1178;
	wire x_1179;
	wire x_1180;
	wire x_1181;
	wire x_1182;
	wire x_1183;
	wire x_1184;
	wire x_1185;
	wire x_1186;
	wire x_1187;
	wire x_1188;
	wire x_1189;
	wire x_1190;
	wire x_1191;
	wire x_1192;
	wire x_1193;
	wire x_1194;
	wire x_1195;
	wire x_1196;
	wire x_1197;
	wire x_1198;
	wire x_1199;
	wire x_1200;
	wire x_1201;
	wire x_1202;
	wire x_1203;
	wire x_1204;
	wire x_1205;
	wire x_1206;
	wire x_1207;
	wire x_1208;
	wire x_1209;
	wire x_1210;
	wire x_1211;
	wire x_1212;
	wire x_1213;
	wire x_1214;
	wire x_1215;
	wire x_1216;
	wire x_1217;
	wire x_1218;
	wire x_1219;
	wire x_1220;
	wire x_1221;
	wire x_1222;
	wire x_1223;
	wire x_1224;
	wire x_1225;
	wire x_1226;
	wire x_1227;
	wire x_1228;
	wire x_1229;
	wire x_1230;
	wire x_1231;
	wire x_1232;
	wire x_1233;
	wire x_1234;
	wire x_1235;
	wire x_1236;
	wire x_1237;
	wire x_1238;
	wire x_1239;
	wire x_1240;
	wire x_1241;
	wire x_1242;
	wire x_1243;
	wire x_1244;
	wire x_1245;
	wire x_1246;
	wire x_1247;
	wire x_1248;
	wire x_1249;
	wire x_1250;
	wire x_1251;
	wire x_1252;
	wire x_1253;
	wire x_1254;
	wire x_1255;
	wire x_1256;
	wire x_1257;
	wire x_1258;
	wire x_1259;
	wire x_1260;
	wire x_1261;
	wire x_1262;
	wire x_1263;
	wire x_1264;
	wire x_1265;
	wire x_1266;
	wire x_1267;
	wire x_1268;
	wire x_1269;
	wire x_1270;
	wire x_1271;
	wire x_1272;
	wire x_1273;
	wire x_1274;
	wire x_1275;
	wire x_1276;
	wire x_1277;
	wire x_1278;
	wire x_1279;
	wire x_1280;
	wire x_1281;
	wire x_1282;
	wire x_1283;
	wire x_1284;
	wire x_1285;
	wire x_1286;
	wire x_1287;
	wire x_1288;
	wire x_1289;
	wire x_1290;
	wire x_1291;
	wire x_1292;
	wire x_1293;
	wire x_1294;
	wire x_1295;
	wire x_1296;
	wire x_1297;
	wire x_1298;
	wire x_1299;
	wire x_1300;
	wire x_1301;
	wire x_1302;
	wire x_1303;
	wire x_1304;
	wire x_1305;
	wire x_1306;
	wire x_1307;
	wire x_1308;
	wire x_1309;
	wire x_1310;
	wire x_1311;
	wire x_1312;
	wire x_1313;
	wire x_1314;
	wire x_1315;
	wire x_1316;
	wire x_1317;
	wire x_1318;
	wire x_1319;
	wire x_1320;
	wire x_1321;
	wire x_1322;
	wire x_1323;
	wire x_1324;
	wire x_1325;
	wire x_1326;
	wire x_1327;
	wire x_1328;
	wire x_1329;
	wire x_1330;
	wire x_1331;
	wire x_1332;
	wire x_1333;
	wire x_1334;
	wire x_1335;
	wire x_1336;
	wire x_1337;
	wire x_1338;
	wire x_1339;
	wire x_1340;
	wire x_1341;
	wire x_1342;
	wire x_1343;
	wire x_1344;
	wire x_1345;
	wire x_1346;
	wire x_1347;
	wire x_1348;
	wire x_1349;
	wire x_1350;
	wire x_1351;
	wire x_1352;
	wire x_1353;
	wire x_1354;
	wire x_1355;
	wire x_1356;
	wire x_1357;
	wire x_1358;
	wire x_1359;
	wire x_1360;
	wire x_1361;
	wire x_1362;
	wire x_1363;
	wire x_1364;
	wire x_1365;
	wire x_1366;
	wire x_1367;
	wire x_1368;
	wire x_1369;
	wire x_1370;
	wire x_1371;
	wire x_1372;
	wire x_1373;
	wire x_1374;
	wire x_1375;
	wire x_1376;
	wire x_1377;
	wire x_1378;
	wire x_1379;
	wire x_1380;
	wire x_1381;
	wire x_1382;
	wire x_1383;
	wire x_1384;
	wire x_1385;
	wire x_1386;
	wire x_1387;
	wire x_1388;
	wire x_1389;
	wire x_1390;
	wire x_1391;
	wire x_1392;
	wire x_1393;
	wire x_1394;
	wire x_1395;
	wire x_1396;
	wire x_1397;
	wire x_1398;
	wire x_1399;
	wire x_1400;
	wire x_1401;
	wire x_1402;
	wire x_1403;
	wire x_1404;
	wire x_1405;
	wire x_1406;
	wire x_1407;
	wire x_1408;
	wire x_1409;
	wire x_1410;
	wire x_1411;
	wire x_1412;
	wire x_1413;
	wire x_1414;
	wire x_1415;
	wire x_1416;
	wire x_1417;
	wire x_1418;
	wire x_1419;
	wire x_1420;
	wire x_1421;
	wire x_1422;
	wire x_1423;
	wire x_1424;
	wire x_1425;
	wire x_1426;
	wire x_1427;
	wire x_1428;
	wire x_1429;
	wire x_1430;
	wire x_1431;
	wire x_1432;
	wire x_1433;
	wire x_1434;
	wire x_1435;
	wire x_1436;
	wire x_1437;
	wire x_1438;
	wire x_1439;
	wire x_1440;
	wire x_1441;
	wire x_1442;
	wire x_1443;
	wire x_1444;
	wire x_1445;
	wire x_1446;
	wire x_1447;
	wire x_1448;
	wire x_1449;
	wire x_1450;
	wire x_1451;
	wire x_1452;
	wire x_1453;
	wire x_1454;
	wire x_1455;
	wire x_1456;
	wire x_1457;
	wire x_1458;
	wire x_1459;
	wire x_1460;
	wire x_1461;
	wire x_1462;
	wire x_1463;
	wire x_1464;
	wire x_1465;
	wire x_1466;
	wire x_1467;
	wire x_1468;
	wire x_1469;
	wire x_1470;
	wire x_1471;
	wire x_1472;
	wire x_1473;
	wire x_1474;
	wire x_1475;
	wire x_1476;
	wire x_1477;
	wire x_1478;
	wire x_1479;
	wire x_1480;
	wire x_1481;
	wire x_1482;
	wire x_1483;
	wire x_1484;
	wire x_1485;
	wire x_1486;
	wire x_1487;
	wire x_1488;
	wire x_1489;
	wire x_1490;
	wire x_1491;
	wire x_1492;
	wire x_1493;
	wire x_1494;
	wire x_1495;
	wire x_1496;
	wire x_1497;
	wire x_1498;
	wire x_1499;
	wire x_1500;
	wire x_1501;
	wire x_1502;
	wire x_1503;
	wire x_1504;
	wire x_1505;
	wire x_1506;
	wire x_1507;
	wire x_1508;
	wire x_1509;
	wire x_1510;
	wire x_1511;
	wire x_1512;
	wire x_1513;
	wire x_1514;
	wire x_1515;
	wire x_1516;
	wire x_1517;
	wire x_1518;
	wire x_1519;
	wire x_1520;
	wire x_1521;
	wire x_1522;
	wire x_1523;
	wire x_1524;
	wire x_1525;
	wire x_1526;
	wire x_1527;
	wire x_1528;
	wire x_1529;
	wire x_1530;
	wire x_1531;
	wire x_1532;
	wire x_1533;
	wire x_1534;
	wire x_1535;
	wire x_1536;
	wire x_1537;
	wire x_1538;
	wire x_1539;
	wire x_1540;
	wire x_1541;
	wire x_1542;
	wire x_1543;
	wire x_1544;
	wire x_1545;
	wire x_1546;
	wire x_1547;
	wire x_1548;
	wire x_1549;
	wire x_1550;
	wire x_1551;
	wire x_1552;
	wire x_1553;
	wire x_1554;
	wire x_1555;
	wire x_1556;
	wire x_1557;
	wire x_1558;
	wire x_1559;
	wire x_1560;
	wire x_1561;
	wire x_1562;
	wire x_1563;
	wire x_1564;
	wire x_1565;
	wire x_1566;
	wire x_1567;
	wire x_1568;
	wire x_1569;
	wire x_1570;
	wire x_1571;
	wire x_1572;
	wire x_1573;
	wire x_1574;
	wire x_1575;
	wire x_1576;
	wire x_1577;
	wire x_1578;
	wire x_1579;
	wire x_1580;
	wire x_1581;
	wire x_1582;
	wire x_1583;
	wire x_1584;
	wire x_1585;
	wire x_1586;
	wire x_1587;
	wire x_1588;
	wire x_1589;
	wire x_1590;
	wire x_1591;
	wire x_1592;
	wire x_1593;
	wire x_1594;
	wire x_1595;
	wire x_1596;
	wire x_1597;
	wire x_1598;
	wire x_1599;
	wire x_1600;
	wire x_1601;
	wire x_1602;
	wire x_1603;
	wire x_1604;
	wire x_1605;
	wire x_1606;
	wire x_1607;
	wire x_1608;
	wire x_1609;
	wire x_1610;
	wire x_1611;
	wire x_1612;
	wire x_1613;
	wire x_1614;
	wire x_1615;
	wire x_1616;
	wire x_1617;
	wire x_1618;
	wire x_1619;
	wire x_1620;
	wire x_1621;
	wire x_1622;
	wire x_1623;
	wire x_1624;
	wire x_1625;
	wire x_1626;
	wire x_1627;
	wire x_1628;
	wire x_1629;
	wire x_1630;
	wire x_1631;
	wire x_1632;
	wire x_1633;
	wire x_1634;
	wire x_1635;
	wire x_1636;
	wire x_1637;
	wire x_1638;
	wire x_1639;
	wire x_1640;
	wire x_1641;
	wire x_1642;
	wire x_1643;
	wire x_1644;
	wire x_1645;
	wire x_1646;
	wire x_1647;
	wire x_1648;
	wire x_1649;
	wire x_1650;
	wire x_1651;
	wire x_1652;
	wire x_1653;
	wire x_1654;
	wire x_1655;
	wire x_1656;
	wire x_1657;
	wire x_1658;
	wire x_1659;
	wire x_1660;
	wire x_1661;
	wire x_1662;
	wire x_1663;
	wire x_1664;
	wire x_1665;
	wire x_1666;
	wire x_1667;
	wire x_1668;
	wire x_1669;
	wire x_1670;
	wire x_1671;
	wire x_1672;
	wire x_1673;
	wire x_1674;
	wire x_1675;
	wire x_1676;
	wire x_1677;
	wire x_1678;
	wire x_1679;
	wire x_1680;
	wire x_1681;
	wire x_1682;
	wire x_1683;
	wire x_1684;
	wire x_1685;
	wire x_1686;
	wire x_1687;
	wire x_1688;
	wire x_1689;
	wire x_1690;
	wire x_1691;
	wire x_1692;
	wire x_1693;
	wire x_1694;
	wire x_1695;
	wire x_1696;
	wire x_1697;
	wire x_1698;
	wire x_1699;
	wire x_1700;
	wire x_1701;
	wire x_1702;
	wire x_1703;
	wire x_1704;
	wire x_1705;
	wire x_1706;
	wire x_1707;
	wire x_1708;
	wire x_1709;
	wire x_1710;
	wire x_1711;
	wire x_1712;
	wire x_1713;
	wire x_1714;
	wire x_1715;
	wire x_1716;
	wire x_1717;
	wire x_1718;
	wire x_1719;
	wire x_1720;
	wire x_1721;
	wire x_1722;
	wire x_1723;
	wire x_1724;
	wire x_1725;
	wire x_1726;
	wire x_1727;
	wire x_1728;
	wire x_1729;
	wire x_1730;
	wire x_1731;
	wire x_1732;
	wire x_1733;
	wire x_1734;
	wire x_1735;
	wire x_1736;
	wire x_1737;
	wire x_1738;
	wire x_1739;
	wire x_1740;
	wire x_1741;
	wire x_1742;
	wire x_1743;
	wire x_1744;
	wire x_1745;
	wire x_1746;
	wire x_1747;
	wire x_1748;
	wire x_1749;
	wire x_1750;
	wire x_1751;
	wire x_1752;
	wire x_1753;
	wire x_1754;
	wire x_1755;
	wire x_1756;
	wire x_1757;
	wire x_1758;
	wire x_1759;
	wire x_1760;
	wire x_1761;
	wire x_1762;
	wire x_1763;
	wire x_1764;
	wire x_1765;
	wire x_1766;
	wire x_1767;
	wire x_1768;
	wire x_1769;
	wire x_1770;
	wire x_1771;
	wire x_1772;
	wire x_1773;
	wire x_1774;
	wire x_1775;
	wire x_1776;
	wire x_1777;
	wire x_1778;
	wire x_1779;
	wire x_1780;
	wire x_1781;
	wire x_1782;
	wire x_1783;
	wire x_1784;
	wire x_1785;
	wire x_1786;
	wire x_1787;
	wire x_1788;
	wire x_1789;
	wire x_1790;
	wire x_1791;
	wire x_1792;
	wire x_1793;
	wire x_1794;
	wire x_1795;
	wire x_1796;
	wire x_1797;
	wire x_1798;
	wire x_1799;
	wire x_1800;
	wire x_1801;
	wire x_1802;
	wire x_1803;
	wire x_1804;
	wire x_1805;
	wire x_1806;
	wire x_1807;
	wire x_1808;
	wire x_1809;
	wire x_1810;
	wire x_1811;
	wire x_1812;
	wire x_1813;
	wire x_1814;
	wire x_1815;
	wire x_1816;
	wire x_1817;
	wire x_1818;
	wire x_1819;
	wire x_1820;
	wire x_1821;
	wire x_1822;
	wire x_1823;
	wire x_1824;
	wire x_1825;
	wire x_1826;
	wire x_1827;
	wire x_1828;
	wire x_1829;
	wire x_1830;
	wire x_1831;
	wire x_1832;
	wire x_1833;
	wire x_1834;
	wire x_1835;
	wire x_1836;
	wire x_1837;
	wire x_1838;
	wire x_1839;
	wire x_1840;
	wire x_1841;
	wire x_1842;
	wire x_1843;
	wire x_1844;
	wire x_1845;
	wire x_1846;
	wire x_1847;
	wire x_1848;
	wire x_1849;
	wire x_1850;
	wire x_1851;
	wire x_1852;
	wire x_1853;
	wire x_1854;
	wire x_1855;
	wire x_1856;
	wire x_1857;
	wire x_1858;
	wire x_1859;
	wire x_1860;
	wire x_1861;
	wire x_1862;
	wire x_1863;
	wire x_1864;
	wire x_1865;
	wire x_1866;
	wire x_1867;
	wire x_1868;
	wire x_1869;
	wire x_1870;
	wire x_1871;
	wire x_1872;
	wire x_1873;
	wire x_1874;
	wire x_1875;
	wire x_1876;
	wire x_1877;
	wire x_1878;
	wire x_1879;
	wire x_1880;
	wire x_1881;
	wire x_1882;
	wire x_1883;
	wire x_1884;
	wire x_1885;
	wire x_1886;
	wire x_1887;
	wire x_1888;
	wire x_1889;
	wire x_1890;
	wire x_1891;
	wire x_1892;
	wire x_1893;
	wire x_1894;
	wire x_1895;
	wire x_1896;
	wire x_1897;
	wire x_1898;
	wire x_1899;
	wire x_1900;
	wire x_1901;
	wire x_1902;
	wire x_1903;
	wire x_1904;
	wire x_1905;
	wire x_1906;
	wire x_1907;
	wire x_1908;
	wire x_1909;
	wire x_1910;
	wire x_1911;
	wire x_1912;
	wire x_1913;
	wire x_1914;
	wire x_1915;
	wire x_1916;
	wire x_1917;
	wire x_1918;
	wire x_1919;
	wire x_1920;
	wire x_1921;
	wire x_1922;
	wire x_1923;
	wire x_1924;
	wire x_1925;
	wire x_1926;
	wire x_1927;
	wire x_1928;
	wire x_1929;
	wire x_1930;
	wire x_1931;
	wire x_1932;
	wire x_1933;
	wire x_1934;
	wire x_1935;
	wire x_1936;
	wire x_1937;
	wire x_1938;
	wire x_1939;
	wire x_1940;
	wire x_1941;
	wire x_1942;
	wire x_1943;
	wire x_1944;
	wire x_1945;
	wire x_1946;
	wire x_1947;
	wire x_1948;
	wire x_1949;
	wire x_1950;
	wire x_1951;
	wire x_1952;
	wire x_1953;
	wire x_1954;
	wire x_1955;
	wire x_1956;
	wire x_1957;
	wire x_1958;
	wire x_1959;
	wire x_1960;
	wire x_1961;
	wire x_1962;
	wire x_1963;
	wire x_1964;
	wire x_1965;
	wire x_1966;
	wire x_1967;
	wire x_1968;
	wire x_1969;
	wire x_1970;
	wire x_1971;
	wire x_1972;
	wire x_1973;
	wire x_1974;
	wire x_1975;
	wire x_1976;
	wire x_1977;
	wire x_1978;
	wire x_1979;
	wire x_1980;
	wire x_1981;
	wire x_1982;
	wire x_1983;
	wire x_1984;
	wire x_1985;
	wire x_1986;
	wire x_1987;
	wire x_1988;
	wire x_1989;
	wire x_1990;
	wire x_1991;
	wire x_1992;
	wire x_1993;
	wire x_1994;
	wire x_1995;
	wire x_1996;
	wire x_1997;
	wire x_1998;
	wire x_1999;
	wire x_2000;
	wire x_2001;
	wire x_2002;
	wire x_2003;
	wire x_2004;
	wire x_2005;
	wire x_2006;
	wire x_2007;
	wire x_2008;
	wire x_2009;
	wire x_2010;
	wire x_2011;
	wire x_2012;
	wire x_2013;
	wire x_2014;
	wire x_2015;
	wire x_2016;
	wire x_2017;
	wire x_2018;
	wire x_2019;
	wire x_2020;
	wire x_2021;
	wire x_2022;
	wire x_2023;
	wire x_2024;
	wire x_2025;
	wire x_2026;
	wire x_2027;
	wire x_2028;
	wire x_2029;
	wire x_2030;
	wire x_2031;
	wire x_2032;
	wire x_2033;
	wire x_2034;
	wire x_2035;
	wire x_2036;
	wire x_2037;
	wire x_2038;
	wire x_2039;
	wire x_2040;
	wire x_2041;
	wire x_2042;
	wire x_2043;
	wire x_2044;
	wire x_2045;
	wire x_2046;
	wire x_2047;
	wire x_2048;
	wire x_2049;
	wire x_2050;
	wire x_2051;
	wire x_2052;
	wire x_2053;
	wire x_2054;
	wire x_2055;
	wire x_2056;
	wire x_2057;
	wire x_2058;
	wire x_2059;
	wire x_2060;
	wire x_2061;
	wire x_2062;
	wire x_2063;
	wire x_2064;
	wire x_2065;
	wire x_2066;
	wire x_2067;
	wire x_2068;
	wire x_2069;
	wire x_2070;
	wire x_2071;
	wire x_2072;
	wire x_2073;
	wire x_2074;
	wire x_2075;
	wire x_2076;
	wire x_2077;
	wire x_2078;
	wire x_2079;
	wire x_2080;
	wire x_2081;
	wire x_2082;
	wire x_2083;
	wire x_2084;
	wire x_2085;
	wire x_2086;
	wire x_2087;
	wire x_2088;
	wire x_2089;
	wire x_2090;
	wire x_2091;
	wire x_2092;
	wire x_2093;
	wire x_2094;
	wire x_2095;
	wire x_2096;
	wire x_2097;
	wire x_2098;
	wire x_2099;
	wire x_2100;
	wire x_2101;
	wire x_2102;
	wire x_2103;
	wire x_2104;
	wire x_2105;
	wire x_2106;
	wire x_2107;
	wire x_2108;
	wire x_2109;
	wire x_2110;
	wire x_2111;
	wire x_2112;
	wire x_2113;
	wire x_2114;
	wire x_2115;
	wire x_2116;
	wire x_2117;
	wire x_2118;
	wire x_2119;
	wire x_2120;
	wire x_2121;
	wire x_2122;
	wire x_2123;
	wire x_2124;
	wire x_2125;
	wire x_2126;
	wire x_2127;
	wire x_2128;
	wire x_2129;
	wire x_2130;
	wire x_2131;
	wire x_2132;
	wire x_2133;
	wire x_2134;
	wire x_2135;
	wire x_2136;
	wire x_2137;
	wire x_2138;
	wire x_2139;
	wire x_2140;
	wire x_2141;
	wire x_2142;
	wire x_2143;
	wire x_2144;
	wire x_2145;
	wire x_2146;
	wire x_2147;
	wire x_2148;
	wire x_2149;
	wire x_2150;
	wire x_2151;
	wire x_2152;
	wire x_2153;
	wire x_2154;
	wire x_2155;
	wire x_2156;
	wire x_2157;
	wire x_2158;
	wire x_2159;
	wire x_2160;
	wire x_2161;
	wire x_2162;
	wire x_2163;
	wire x_2164;
	wire x_2165;
	wire x_2166;
	wire x_2167;
	wire x_2168;
	wire x_2169;
	wire x_2170;
	wire x_2171;
	wire x_2172;
	wire x_2173;
	wire x_2174;
	wire x_2175;
	wire x_2176;
	wire x_2177;
	wire x_2178;
	wire x_2179;
	wire x_2180;
	wire x_2181;
	wire x_2182;
	wire x_2183;
	wire x_2184;
	wire x_2185;
	wire x_2186;
	wire x_2187;
	wire x_2188;
	wire x_2189;
	wire x_2190;
	wire x_2191;
	wire x_2192;
	wire x_2193;
	wire x_2194;
	wire x_2195;
	wire x_2196;
	wire x_2197;
	wire x_2198;
	wire x_2199;
	wire x_2200;
	wire x_2201;
	wire x_2202;
	wire x_2203;
	wire x_2204;
	wire x_2205;
	wire x_2206;
	wire x_2207;
	wire x_2208;
	wire x_2209;
	wire x_2210;
	wire x_2211;
	wire x_2212;
	wire x_2213;
	wire x_2214;
	wire x_2215;
	wire x_2216;
	wire x_2217;
	wire x_2218;
	wire x_2219;
	wire x_2220;
	wire x_2221;
	wire x_2222;
	wire x_2223;
	wire x_2224;
	wire x_2225;
	wire x_2226;
	wire x_2227;
	wire x_2228;
	wire x_2229;
	wire x_2230;
	wire x_2231;
	wire x_2232;
	wire x_2233;
	wire x_2234;
	wire x_2235;
	wire x_2236;
	wire x_2237;
	wire x_2238;
	wire x_2239;
	wire x_2240;
	wire x_2241;
	wire x_2242;
	wire x_2243;
	wire x_2244;
	wire x_2245;
	wire x_2246;
	wire x_2247;
	wire x_2248;
	wire x_2249;
	wire x_2250;
	wire x_2251;
	wire x_2252;
	wire x_2253;
	wire x_2254;
	wire x_2255;
	wire x_2256;
	wire x_2257;
	wire x_2258;
	wire x_2259;
	wire x_2260;
	wire x_2261;
	wire x_2262;
	wire x_2263;
	wire x_2264;
	wire x_2265;
	wire x_2266;
	wire x_2267;
	wire x_2268;
	wire x_2269;
	wire x_2270;
	wire x_2271;
	wire x_2272;
	wire x_2273;
	wire x_2274;
	wire x_2275;
	wire x_2276;
	wire x_2277;
	wire x_2278;
	wire x_2279;
	wire x_2280;
	wire x_2281;
	wire x_2282;
	wire x_2283;
	wire x_2284;
	wire x_2285;
	wire x_2286;
	wire x_2287;
	wire x_2288;
	wire x_2289;
	wire x_2290;
	wire x_2291;
	wire x_2292;
	wire x_2293;
	wire x_2294;
	wire x_2295;
	wire x_2296;
	wire x_2297;
	wire x_2298;
	wire x_2299;
	wire x_2300;
	wire x_2301;
	wire x_2302;
	wire x_2303;
	wire x_2304;
	wire x_2305;
	wire x_2306;
	wire x_2307;
	wire x_2308;
	wire x_2309;
	wire x_2310;
	wire x_2311;
	wire x_2312;
	wire x_2313;
	wire x_2314;
	wire x_2315;
	wire x_2316;
	wire x_2317;
	wire x_2318;
	wire x_2319;
	wire x_2320;
	wire x_2321;
	wire x_2322;
	wire x_2323;
	wire x_2324;
	wire x_2325;
	wire x_2326;
	wire x_2327;
	wire x_2328;
	wire x_2329;
	wire x_2330;
	wire x_2331;
	wire x_2332;
	wire x_2333;
	wire x_2334;
	wire x_2335;
	wire x_2336;
	wire x_2337;
	wire x_2338;
	wire x_2339;
	wire x_2340;
	wire x_2341;
	wire x_2342;
	wire x_2343;
	wire x_2344;
	wire x_2345;
	wire x_2346;
	wire x_2347;
	wire x_2348;
	wire x_2349;
	wire x_2350;
	wire x_2351;
	wire x_2352;
	wire x_2353;
	wire x_2354;
	wire x_2355;
	wire x_2356;
	wire x_2357;
	wire x_2358;
	wire x_2359;
	wire x_2360;
	wire x_2361;
	wire x_2362;
	wire x_2363;
	wire x_2364;
	wire x_2365;
	wire x_2366;
	wire x_2367;
	wire x_2368;
	wire x_2369;
	wire x_2370;
	wire x_2371;
	wire x_2372;
	wire x_2373;
	wire x_2374;
	wire x_2375;
	wire x_2376;
	wire x_2377;
	wire x_2378;
	wire x_2379;
	wire x_2380;
	wire x_2381;
	wire x_2382;
	wire x_2383;
	wire x_2384;
	wire x_2385;
	wire x_2386;
	wire x_2387;
	wire x_2388;
	wire x_2389;
	wire x_2390;
	wire x_2391;
	wire x_2392;
	wire x_2393;
	wire x_2394;
	wire x_2395;
	wire x_2396;
	wire x_2397;
	wire x_2398;
	wire x_2399;
	wire x_2400;
	wire x_2401;
	wire x_2402;
	wire x_2403;
	wire x_2404;
	wire x_2405;
	wire x_2406;
	wire x_2407;
	wire x_2408;
	wire x_2409;
	wire x_2410;
	wire x_2411;
	wire x_2412;
	wire x_2413;
	wire x_2414;
	wire x_2415;
	wire x_2416;
	wire x_2417;
	wire x_2418;
	wire x_2419;
	wire x_2420;
	wire x_2421;
	wire x_2422;
	wire x_2423;
	wire x_2424;
	wire x_2425;
	wire x_2426;
	wire x_2427;
	wire x_2428;
	wire x_2429;
	wire x_2430;
	wire x_2431;
	wire x_2432;
	wire x_2433;
	wire x_2434;
	wire x_2435;
	wire x_2436;
	wire x_2437;
	wire x_2438;
	wire x_2439;
	wire x_2440;
	wire x_2441;
	wire x_2442;
	wire x_2443;
	wire x_2444;
	wire x_2445;
	wire x_2446;
	wire x_2447;
	wire x_2448;
	wire x_2449;
	wire x_2450;
	wire x_2451;
	wire x_2452;
	wire x_2453;
	wire x_2454;
	wire x_2455;
	wire x_2456;
	wire x_2457;
	wire x_2458;
	wire x_2459;
	wire x_2460;
	wire x_2461;
	wire x_2462;
	wire x_2463;
	wire x_2464;
	wire x_2465;
	wire x_2466;
	wire x_2467;
	wire x_2468;
	wire x_2469;
	wire x_2470;
	wire x_2471;
	wire x_2472;
	wire x_2473;
	wire x_2474;
	wire x_2475;
	wire x_2476;
	wire x_2477;
	wire x_2478;
	wire x_2479;
	wire x_2480;
	wire x_2481;
	wire x_2482;
	wire x_2483;
	wire x_2484;
	wire x_2485;
	wire x_2486;
	wire x_2487;
	wire x_2488;
	wire x_2489;
	wire x_2490;
	wire x_2491;
	wire x_2492;
	wire x_2493;
	wire x_2494;
	wire x_2495;
	wire x_2496;
	wire x_2497;
	wire x_2498;
	wire x_2499;
	wire x_2500;
	wire x_2501;
	wire x_2502;
	wire x_2503;
	wire x_2504;
	wire x_2505;
	wire x_2506;
	wire x_2507;
	wire x_2508;
	wire x_2509;
	wire x_2510;
	wire x_2511;
	wire x_2512;
	wire x_2513;
	wire x_2514;
	wire x_2515;
	wire x_2516;
	wire x_2517;
	wire x_2518;
	wire x_2519;
	wire x_2520;
	wire x_2521;
	wire x_2522;
	wire x_2523;
	wire x_2524;
	wire x_2525;
	wire x_2526;
	wire x_2527;
	wire x_2528;
	wire x_2529;
	wire x_2530;
	wire x_2531;
	wire x_2532;
	wire x_2533;
	wire x_2534;
	wire x_2535;
	wire x_2536;
	wire x_2537;
	wire x_2538;
	wire x_2539;
	wire x_2540;
	wire x_2541;
	wire x_2542;
	wire x_2543;
	wire x_2544;
	wire x_2545;
	wire x_2546;
	wire x_2547;
	wire x_2548;
	wire x_2549;
	wire x_2550;
	wire x_2551;
	wire x_2552;
	wire x_2553;
	wire x_2554;
	wire x_2555;
	wire x_2556;
	wire x_2557;
	wire x_2558;
	wire x_2559;
	wire x_2560;
	wire x_2561;
	wire x_2562;
	wire x_2563;
	wire x_2564;
	wire x_2565;
	wire x_2566;
	wire x_2567;
	wire x_2568;
	wire x_2569;
	wire x_2570;
	wire x_2571;
	wire x_2572;
	wire x_2573;
	wire x_2574;
	wire x_2575;
	wire x_2576;
	wire x_2577;
	wire x_2578;
	wire x_2579;
	wire x_2580;
	wire x_2581;
	wire x_2582;
	wire x_2583;
	wire x_2584;
	wire x_2585;
	wire x_2586;
	wire x_2587;
	wire x_2588;
	wire x_2589;
	wire x_2590;
	wire x_2591;
	wire x_2592;
	wire x_2593;
	wire x_2594;
	wire x_2595;
	wire x_2596;
	wire x_2597;
	wire x_2598;
	wire x_2599;
	wire x_2600;
	wire x_2601;
	wire x_2602;
	wire x_2603;
	wire x_2604;
	wire x_2605;
	wire x_2606;
	wire x_2607;
	wire x_2608;
	wire x_2609;
	wire x_2610;
	wire x_2611;
	wire x_2612;
	wire x_2613;
	wire x_2614;
	wire x_2615;
	wire x_2616;
	wire x_2617;
	wire x_2618;
	wire x_2619;
	wire x_2620;
	wire x_2621;
	wire x_2622;
	wire x_2623;
	wire x_2624;
	wire x_2625;
	wire x_2626;
	wire x_2627;
	wire x_2628;
	wire x_2629;
	wire x_2630;
	wire x_2631;
	wire x_2632;
	wire x_2633;
	wire x_2634;
	wire x_2635;
	wire x_2636;
	wire x_2637;
	wire x_2638;
	wire x_2639;
	wire x_2640;
	wire x_2641;
	wire x_2642;
	wire x_2643;
	wire x_2644;
	wire x_2645;
	wire x_2646;
	wire x_2647;
	wire x_2648;
	wire x_2649;
	wire x_2650;
	wire x_2651;
	wire x_2652;
	wire x_2653;
	wire x_2654;
	wire x_2655;
	wire x_2656;
	wire x_2657;
	wire x_2658;
	wire x_2659;
	wire x_2660;
	wire x_2661;
	wire x_2662;
	wire x_2663;
	wire x_2664;
	wire x_2665;
	wire x_2666;
	wire x_2667;
	wire x_2668;
	wire x_2669;
	wire x_2670;
	wire x_2671;
	wire x_2672;
	wire x_2673;
	wire x_2674;
	wire x_2675;
	wire x_2676;
	wire x_2677;
	wire x_2678;
	wire x_2679;
	wire x_2680;
	wire x_2681;
	wire x_2682;
	wire x_2683;
	wire x_2684;
	wire x_2685;
	wire x_2686;
	wire x_2687;
	wire x_2688;
	wire x_2689;
	wire x_2690;
	wire x_2691;
	wire x_2692;
	wire x_2693;
	wire x_2694;
	wire x_2695;
	wire x_2696;
	wire x_2697;
	wire x_2698;
	wire x_2699;
	wire x_2700;
	wire x_2701;
	wire x_2702;
	wire x_2703;
	wire x_2704;
	wire x_2705;
	wire x_2706;
	wire x_2707;
	wire x_2708;
	wire x_2709;
	wire x_2710;
	wire x_2711;
	wire x_2712;
	wire x_2713;
	wire x_2714;
	wire x_2715;
	wire x_2716;
	wire x_2717;
	wire x_2718;
	wire x_2719;
	wire x_2720;
	wire x_2721;
	wire x_2722;
	wire x_2723;
	wire x_2724;
	wire x_2725;
	wire x_2726;
	wire x_2727;
	wire x_2728;
	wire x_2729;
	wire x_2730;
	wire x_2731;
	wire x_2732;
	wire x_2733;
	wire x_2734;
	wire x_2735;
	wire x_2736;
	wire x_2737;
	wire x_2738;
	wire x_2739;
	wire x_2740;
	wire x_2741;
	wire x_2742;
	wire x_2743;
	wire x_2744;
	wire x_2745;
	wire x_2746;
	wire x_2747;
	wire x_2748;
	wire x_2749;
	wire x_2750;
	wire x_2751;
	wire x_2752;
	wire x_2753;
	wire x_2754;
	wire x_2755;
	wire x_2756;
	wire x_2757;
	wire x_2758;
	wire x_2759;
	wire x_2760;
	wire x_2761;
	wire x_2762;
	wire x_2763;
	wire x_2764;
	wire x_2765;
	wire x_2766;
	wire x_2767;
	wire x_2768;
	wire x_2769;
	wire x_2770;
	wire x_2771;
	wire x_2772;
	wire x_2773;
	wire x_2774;
	wire x_2775;
	wire x_2776;
	wire x_2777;
	wire x_2778;
	wire x_2779;
	wire x_2780;
	wire x_2781;
	wire x_2782;
	wire x_2783;
	wire x_2784;
	wire x_2785;
	wire x_2786;
	wire x_2787;
	wire x_2788;
	wire x_2789;
	wire x_2790;
	wire x_2791;
	wire x_2792;
	wire x_2793;
	wire x_2794;
	wire x_2795;
	wire x_2796;
	wire x_2797;
	wire x_2798;
	wire x_2799;
	wire x_2800;
	wire x_2801;
	wire x_2802;
	wire x_2803;
	wire x_2804;
	wire x_2805;
	wire x_2806;
	wire x_2807;
	wire x_2808;
	wire x_2809;
	wire x_2810;
	wire x_2811;
	wire x_2812;
	wire x_2813;
	wire x_2814;
	wire x_2815;
	wire x_2816;
	wire x_2817;
	wire x_2818;
	wire x_2819;
	wire x_2820;
	wire x_2821;
	wire x_2822;
	wire x_2823;
	wire x_2824;
	wire x_2825;
	wire x_2826;
	wire x_2827;
	wire x_2828;
	wire x_2829;
	wire x_2830;
	wire x_2831;
	wire x_2832;
	wire x_2833;
	wire x_2834;
	wire x_2835;
	wire x_2836;
	wire x_2837;
	wire x_2838;
	wire x_2839;
	wire x_2840;
	wire x_2841;
	wire x_2842;
	wire x_2843;
	wire x_2844;
	wire x_2845;
	wire x_2846;
	wire x_2847;
	wire x_2848;
	wire x_2849;
	wire x_2850;
	wire x_2851;
	wire x_2852;
	wire x_2853;
	wire x_2854;
	wire x_2855;
	wire x_2856;
	wire x_2857;
	wire x_2858;
	wire x_2859;
	wire x_2860;
	wire x_2861;
	wire x_2862;
	wire x_2863;
	wire x_2864;
	wire x_2865;
	wire x_2866;
	wire x_2867;
	wire x_2868;
	wire x_2869;
	wire x_2870;
	wire x_2871;
	wire x_2872;
	wire x_2873;
	wire x_2874;
	wire x_2875;
	wire x_2876;
	wire x_2877;
	wire x_2878;
	wire x_2879;
	wire x_2880;
	wire x_2881;
	wire x_2882;
	wire x_2883;
	wire x_2884;
	wire x_2885;
	wire x_2886;
	wire x_2887;
	wire x_2888;
	wire x_2889;
	wire x_2890;
	wire x_2891;
	wire x_2892;
	wire x_2893;
	wire x_2894;
	wire x_2895;
	wire x_2896;
	wire x_2897;
	wire x_2898;
	wire x_2899;
	wire x_2900;
	wire x_2901;
	wire x_2902;
	wire x_2903;
	wire x_2904;
	wire x_2905;
	wire x_2906;
	wire x_2907;
	wire x_2908;
	wire x_2909;
	wire x_2910;
	wire x_2911;
	wire x_2912;
	wire x_2913;
	wire x_2914;
	wire x_2915;
	wire x_2916;
	wire x_2917;
	wire x_2918;
	wire x_2919;
	wire x_2920;
	wire x_2921;
	wire x_2922;
	wire x_2923;
	wire x_2924;
	wire x_2925;
	wire x_2926;
	wire x_2927;
	wire x_2928;
	wire x_2929;
	wire x_2930;
	wire x_2931;
	wire x_2932;
	wire x_2933;
	wire x_2934;
	wire x_2935;
	wire x_2936;
	wire x_2937;
	wire x_2938;
	wire x_2939;
	wire x_2940;
	wire x_2941;
	wire x_2942;
	wire x_2943;
	wire x_2944;
	wire x_2945;
	wire x_2946;
	wire x_2947;
	wire x_2948;
	wire x_2949;
	wire x_2950;
	wire x_2951;
	wire x_2952;
	wire x_2953;
	wire x_2954;
	wire x_2955;
	wire x_2956;
	wire x_2957;
	wire x_2958;
	wire x_2959;
	wire x_2960;
	wire x_2961;
	wire x_2962;
	wire x_2963;
	wire x_2964;
	wire x_2965;
	wire x_2966;
	wire x_2967;
	wire x_2968;
	wire x_2969;
	wire x_2970;
	wire x_2971;
	wire x_2972;
	wire x_2973;
	wire x_2974;
	wire x_2975;
	wire x_2976;
	wire x_2977;
	wire x_2978;
	wire x_2979;
	wire x_2980;
	wire x_2981;
	wire x_2982;
	wire x_2983;
	wire x_2984;
	wire x_2985;
	wire x_2986;
	wire x_2987;
	wire x_2988;
	wire x_2989;
	wire x_2990;
	wire x_2991;
	wire x_2992;
	wire x_2993;
	wire x_2994;
	wire x_2995;
	wire x_2996;
	wire x_2997;
	wire x_2998;
	wire x_2999;
	wire x_3000;
	wire x_3001;
	wire x_3002;
	wire x_3003;
	wire x_3004;
	wire x_3005;
	wire x_3006;
	wire x_3007;
	wire x_3008;
	wire x_3009;
	wire x_3010;
	wire x_3011;
	wire x_3012;
	wire x_3013;
	wire x_3014;
	wire x_3015;
	wire x_3016;
	wire x_3017;
	wire x_3018;
	wire x_3019;
	wire x_3020;
	wire x_3021;
	wire x_3022;
	wire x_3023;
	wire x_3024;
	wire x_3025;
	wire x_3026;
	wire x_3027;
	wire x_3028;
	wire x_3029;
	wire x_3030;
	wire x_3031;
	wire x_3032;
	wire x_3033;
	wire x_3034;
	wire x_3035;
	wire x_3036;
	wire x_3037;
	wire x_3038;
	wire x_3039;
	wire x_3040;
	wire x_3041;
	wire x_3042;
	wire x_3043;
	wire x_3044;
	wire x_3045;
	wire x_3046;
	wire x_3047;
	wire x_3048;
	wire x_3049;
	wire x_3050;
	wire x_3051;
	wire x_3052;
	wire x_3053;
	wire x_3054;
	wire x_3055;
	wire x_3056;
	wire x_3057;
	wire x_3058;
	wire x_3059;
	wire x_3060;
	wire x_3061;
	wire x_3062;
	wire x_3063;
	wire x_3064;
	wire x_3065;
	wire x_3066;
	wire x_3067;
	wire x_3068;
	wire x_3069;
	wire x_3070;
	wire x_3071;
	wire x_3072;
	wire x_3073;
	wire x_3074;
	wire x_3075;
	wire x_3076;
	wire x_3077;
	wire x_3078;
	wire x_3079;
	wire x_3080;
	wire x_3081;
	wire x_3082;
	wire x_3083;
	wire x_3084;
	wire x_3085;
	wire x_3086;
	wire x_3087;
	wire x_3088;
	wire x_3089;
	wire x_3090;
	wire x_3091;
	wire x_3092;
	wire x_3093;
	wire x_3094;
	wire x_3095;
	wire x_3096;
	wire x_3097;
	wire x_3098;
	wire x_3099;
	wire x_3100;
	wire x_3101;
	wire x_3102;
	wire x_3103;
	wire x_3104;
	wire x_3105;
	wire x_3106;
	wire x_3107;
	wire x_3108;
	wire x_3109;
	wire x_3110;
	wire x_3111;
	wire x_3112;
	wire x_3113;
	wire x_3114;
	wire x_3115;
	wire x_3116;
	wire x_3117;
	wire x_3118;
	wire x_3119;
	wire x_3120;
	wire x_3121;
	wire x_3122;
	wire x_3123;
	wire x_3124;
	wire x_3125;
	wire x_3126;
	wire x_3127;
	wire x_3128;
	wire x_3129;
	wire x_3130;
	wire x_3131;
	wire x_3132;
	wire x_3133;
	wire x_3134;
	wire x_3135;
	wire x_3136;
	wire x_3137;
	wire x_3138;
	wire x_3139;
	wire x_3140;
	wire x_3141;
	wire x_3142;
	wire x_3143;
	wire x_3144;
	wire x_3145;
	wire x_3146;
	wire x_3147;
	wire x_3148;
	wire x_3149;
	wire x_3150;
	wire x_3151;
	wire x_3152;
	wire x_3153;
	wire x_3154;
	wire x_3155;
	wire x_3156;
	wire x_3157;
	wire x_3158;
	wire x_3159;
	wire x_3160;
	wire x_3161;
	wire x_3162;
	wire x_3163;
	wire x_3164;
	wire x_3165;
	wire x_3166;
	wire x_3167;
	wire x_3168;
	wire x_3169;
	wire x_3170;
	wire x_3171;
	wire x_3172;
	wire x_3173;
	wire x_3174;
	wire x_3175;
	wire x_3176;
	wire x_3177;
	wire x_3178;
	wire x_3179;
	wire x_3180;
	wire x_3181;
	wire x_3182;
	wire x_3183;
	wire x_3184;
	wire x_3185;
	wire x_3186;
	wire x_3187;
	wire x_3188;
	wire x_3189;
	wire x_3190;
	wire x_3191;
	wire x_3192;
	wire x_3193;
	wire x_3194;
	wire x_3195;
	wire x_3196;
	wire x_3197;
	wire x_3198;
	wire x_3199;
	wire x_3200;
	wire x_3201;
	wire x_3202;
	wire x_3203;
	wire x_3204;
	wire x_3205;
	wire x_3206;
	wire x_3207;
	wire x_3208;
	wire x_3209;
	wire x_3210;
	wire x_3211;
	wire x_3212;
	wire x_3213;
	wire x_3214;
	wire x_3215;
	wire x_3216;
	wire x_3217;
	wire x_3218;
	wire x_3219;
	wire x_3220;
	wire x_3221;
	wire x_3222;
	wire x_3223;
	wire x_3224;
	wire x_3225;
	wire x_3226;
	wire x_3227;
	wire x_3228;
	wire x_3229;
	wire x_3230;
	wire x_3231;
	wire x_3232;
	wire x_3233;
	wire x_3234;
	wire x_3235;
	wire x_3236;
	wire x_3237;
	wire x_3238;
	wire x_3239;
	wire x_3240;
	wire x_3241;
	wire x_3242;
	wire x_3243;
	wire x_3244;
	wire x_3245;
	wire x_3246;
	wire x_3247;
	wire x_3248;
	wire x_3249;
	wire x_3250;
	wire x_3251;
	wire x_3252;
	wire x_3253;
	wire x_3254;
	wire x_3255;
	wire x_3256;
	wire x_3257;
	wire x_3258;
	wire x_3259;
	wire x_3260;
	wire x_3261;
	wire x_3262;
	wire x_3263;
	wire x_3264;
	wire x_3265;
	wire x_3266;
	wire x_3267;
	wire x_3268;
	wire x_3269;
	wire x_3270;
	wire x_3271;
	wire x_3272;
	wire x_3273;
	wire x_3274;
	wire x_3275;
	wire x_3276;
	wire x_3277;
	wire x_3278;
	wire x_3279;
	wire x_3280;
	wire x_3281;
	wire x_3282;
	wire x_3283;
	wire x_3284;
	wire x_3285;
	wire x_3286;
	wire x_3287;
	wire x_3288;
	wire x_3289;
	wire x_3290;
	wire x_3291;
	wire x_3292;
	wire x_3293;
	wire x_3294;
	wire x_3295;
	wire x_3296;
	wire x_3297;
	wire x_3298;
	wire x_3299;
	wire x_3300;
	wire x_3301;
	wire x_3302;
	wire x_3303;
	wire x_3304;
	wire x_3305;
	wire x_3306;
	wire x_3307;
	wire x_3308;
	wire x_3309;
	wire x_3310;
	wire x_3311;
	wire x_3312;
	wire x_3313;
	wire x_3314;
	wire x_3315;
	wire x_3316;
	wire x_3317;
	wire x_3318;
	wire x_3319;
	wire x_3320;
	wire x_3321;
	wire x_3322;
	wire x_3323;
	wire x_3324;
	wire x_3325;
	wire x_3326;
	wire x_3327;
	wire x_3328;
	wire x_3329;
	wire x_3330;
	wire x_3331;
	wire x_3332;
	wire x_3333;
	wire x_3334;
	wire x_3335;
	wire x_3336;
	wire x_3337;
	wire x_3338;
	wire x_3339;
	wire x_3340;
	wire x_3341;
	wire x_3342;
	wire x_3343;
	wire x_3344;
	wire x_3345;
	wire x_3346;
	wire x_3347;
	wire x_3348;
	wire x_3349;
	wire x_3350;
	wire x_3351;
	wire x_3352;
	wire x_3353;
	wire x_3354;
	wire x_3355;
	wire x_3356;
	wire x_3357;
	wire x_3358;
	wire x_3359;
	wire x_3360;
	wire x_3361;
	wire x_3362;
	wire x_3363;
	wire x_3364;
	wire x_3365;
	wire x_3366;
	wire x_3367;
	wire x_3368;
	wire x_3369;
	wire x_3370;
	wire x_3371;
	wire x_3372;
	wire x_3373;
	wire x_3374;
	wire x_3375;
	wire x_3376;
	wire x_3377;
	wire x_3378;
	wire x_3379;
	wire x_3380;
	wire x_3381;
	wire x_3382;
	wire x_3383;
	wire x_3384;
	wire x_3385;
	wire x_3386;
	wire x_3387;
	wire x_3388;
	wire x_3389;
	wire x_3390;
	wire x_3391;
	wire x_3392;
	wire x_3393;
	wire x_3394;
	wire x_3395;
	wire x_3396;
	wire x_3397;
	wire x_3398;
	wire x_3399;
	wire x_3400;
	wire x_3401;
	wire x_3402;
	wire x_3403;
	wire x_3404;
	wire x_3405;
	wire x_3406;
	wire x_3407;
	wire x_3408;
	wire x_3409;
	wire x_3410;
	wire x_3411;
	wire x_3412;
	wire x_3413;
	wire x_3414;
	wire x_3415;
	wire x_3416;
	wire x_3417;
	wire x_3418;
	wire x_3419;
	wire x_3420;
	wire x_3421;
	wire x_3422;
	wire x_3423;
	wire x_3424;
	wire x_3425;
	wire x_3426;
	wire x_3427;
	wire x_3428;
	wire x_3429;
	wire x_3430;
	wire x_3431;
	wire x_3432;
	wire x_3433;
	wire x_3434;
	wire x_3435;
	wire x_3436;
	wire x_3437;
	wire x_3438;
	wire x_3439;
	wire x_3440;
	wire x_3441;
	wire x_3442;
	wire x_3443;
	wire x_3444;
	wire x_3445;
	wire x_3446;
	wire x_3447;
	wire x_3448;
	wire x_3449;
	wire x_3450;
	wire x_3451;
	wire x_3452;
	wire x_3453;
	wire x_3454;
	wire x_3455;
	wire x_3456;
	wire x_3457;
	wire x_3458;
	wire x_3459;
	wire x_3460;
	wire x_3461;
	wire x_3462;
	wire x_3463;
	wire x_3464;
	wire x_3465;
	wire x_3466;
	wire x_3467;
	wire x_3468;
	wire x_3469;
	wire x_3470;
	wire x_3471;
	wire x_3472;
	wire x_3473;
	wire x_3474;
	wire x_3475;
	wire x_3476;
	wire x_3477;
	wire x_3478;
	wire x_3479;
	wire x_3480;
	wire x_3481;
	wire x_3482;
	wire x_3483;
	wire x_3484;
	wire x_3485;
	wire x_3486;
	wire x_3487;
	wire x_3488;
	wire x_3489;
	wire x_3490;
	wire x_3491;
	wire x_3492;
	wire x_3493;
	wire x_3494;
	wire x_3495;
	wire x_3496;
	wire x_3497;
	wire x_3498;
	wire x_3499;
	wire x_3500;
	wire x_3501;
	wire x_3502;
	wire x_3503;
	wire x_3504;
	wire x_3505;
	wire x_3506;
	wire x_3507;
	wire x_3508;
	wire x_3509;
	wire x_3510;
	wire x_3511;
	wire x_3512;
	wire x_3513;
	wire x_3514;
	wire x_3515;
	wire x_3516;
	wire x_3517;
	wire x_3518;
	wire x_3519;
	wire x_3520;
	wire x_3521;
	wire x_3522;
	wire x_3523;
	wire x_3524;
	wire x_3525;
	wire x_3526;
	wire x_3527;
	wire x_3528;
	wire x_3529;
	wire x_3530;
	wire x_3531;
	wire x_3532;
	wire x_3533;
	wire x_3534;
	wire x_3535;
	wire x_3536;
	wire x_3537;
	wire x_3538;
	wire x_3539;
	wire x_3540;
	wire x_3541;
	wire x_3542;
	wire x_3543;
	wire x_3544;
	wire x_3545;
	wire x_3546;
	wire x_3547;
	wire x_3548;
	wire x_3549;
	wire x_3550;
	wire x_3551;
	wire x_3552;
	wire x_3553;
	wire x_3554;
	wire x_3555;
	wire x_3556;
	wire x_3557;
	wire x_3558;
	wire x_3559;
	wire x_3560;
	wire x_3561;
	wire x_3562;
	wire x_3563;
	wire x_3564;
	wire x_3565;
	wire x_3566;
	wire x_3567;
	wire x_3568;
	wire x_3569;
	wire x_3570;
	wire x_3571;
	wire x_3572;
	wire x_3573;
	wire x_3574;
	wire x_3575;
	wire x_3576;
	wire x_3577;
	wire x_3578;
	wire x_3579;
	wire x_3580;
	wire x_3581;
	wire x_3582;
	wire x_3583;
	wire x_3584;
	wire x_3585;
	wire x_3586;
	wire x_3587;
	wire x_3588;
	wire x_3589;
	wire x_3590;
	wire x_3591;
	wire x_3592;
	wire x_3593;
	wire x_3594;
	wire x_3595;
	wire x_3596;
	wire x_3597;
	wire x_3598;
	wire x_3599;
	wire x_3600;
	wire x_3601;
	wire x_3602;
	wire x_3603;
	wire x_3604;
	wire x_3605;
	wire x_3606;
	wire x_3607;
	wire x_3608;
	wire x_3609;
	wire x_3610;
	wire x_3611;
	wire x_3612;
	wire x_3613;
	wire x_3614;
	wire x_3615;
	wire x_3616;
	wire x_3617;
	wire x_3618;
	wire x_3619;
	wire x_3620;
	wire x_3621;
	wire x_3622;
	wire x_3623;
	wire x_3624;
	wire x_3625;
	wire x_3626;
	wire x_3627;
	wire x_3628;
	wire x_3629;
	wire x_3630;
	wire x_3631;
	wire x_3632;
	wire x_3633;
	wire x_3634;
	wire x_3635;
	wire x_3636;
	wire x_3637;
	wire x_3638;
	wire x_3639;
	wire x_3640;
	wire x_3641;
	wire x_3642;
	wire x_3643;
	wire x_3644;
	wire x_3645;
	wire x_3646;
	wire x_3647;
	wire x_3648;
	wire x_3649;
	wire x_3650;
	wire x_3651;
	wire x_3652;
	wire x_3653;
	wire x_3654;
	wire x_3655;
	wire x_3656;
	wire x_3657;
	wire x_3658;
	wire x_3659;
	wire x_3660;
	wire x_3661;
	wire x_3662;
	wire x_3663;
	wire x_3664;
	wire x_3665;
	wire x_3666;
	wire x_3667;
	wire x_3668;
	wire x_3669;
	wire x_3670;
	wire x_3671;
	wire x_3672;
	wire x_3673;
	wire x_3674;
	wire x_3675;
	wire x_3676;
	wire x_3677;
	wire x_3678;
	wire x_3679;
	wire x_3680;
	wire x_3681;
	wire x_3682;
	wire x_3683;
	wire x_3684;
	wire x_3685;
	wire x_3686;
	wire x_3687;
	wire x_3688;
	wire x_3689;
	wire x_3690;
	wire x_3691;
	wire x_3692;
	wire x_3693;
	wire x_3694;
	wire x_3695;
	wire x_3696;
	wire x_3697;
	wire x_3698;
	wire x_3699;
	wire x_3700;
	wire x_3701;
	wire x_3702;
	wire x_3703;
	wire x_3704;
	wire x_3705;
	wire x_3706;
	wire x_3707;
	wire x_3708;
	wire x_3709;
	wire x_3710;
	wire x_3711;
	wire x_3712;
	wire x_3713;
	wire x_3714;
	wire x_3715;
	wire x_3716;
	wire x_3717;
	wire x_3718;
	wire x_3719;
	wire x_3720;
	wire x_3721;
	wire x_3722;
	wire x_3723;
	wire x_3724;
	wire x_3725;
	wire x_3726;
	wire x_3727;
	wire x_3728;
	wire x_3729;
	wire x_3730;
	wire x_3731;
	wire x_3732;
	wire x_3733;
	wire x_3734;
	wire x_3735;
	wire x_3736;
	wire x_3737;
	wire x_3738;
	wire x_3739;
	wire x_3740;
	wire x_3741;
	wire x_3742;
	wire x_3743;
	wire x_3744;
	wire x_3745;
	wire x_3746;
	wire x_3747;
	wire x_3748;
	wire x_3749;
	wire x_3750;
	wire x_3751;
	wire x_3752;
	wire x_3753;
	wire x_3754;
	wire x_3755;
	wire x_3756;
	wire x_3757;
	wire x_3758;
	wire x_3759;
	wire x_3760;
	wire x_3761;
	wire x_3762;
	wire x_3763;
	wire x_3764;
	wire x_3765;
	wire x_3766;
	wire x_3767;
	wire x_3768;
	wire x_3769;
	wire x_3770;
	wire x_3771;
	wire x_3772;
	wire x_3773;
	wire x_3774;
	wire x_3775;
	wire x_3776;
	wire x_3777;
	wire x_3778;
	wire x_3779;
	wire x_3780;
	wire x_3781;
	wire x_3782;
	wire x_3783;
	output o_1;
	assign x_1892 = (v_83 | v_59) ;
	assign x_1891 = (v_83 | v_78) ;
	assign x_1890 = (v_84 | v_76) ;
	assign x_1889 = (v_84 | v_50) ;
	assign x_1888 = (((v_63 | ~v_84) | ~v_83) | v_85) ;
	assign x_1887 = (v_86 | v_60) ;
	assign x_1886 = (v_86 | ~v_85) ;
	assign x_1885 = (v_87 | v_74) ;
	assign x_1884 = (v_87 | v_78) ;
	assign x_1883 = (v_88 | v_51) ;
	assign x_1882 = (v_88 | v_63) ;
	assign x_1881 = (((v_76 | ~v_88) | ~v_87) | v_89) ;
	assign x_1880 = (v_90 | v_75) ;
	assign x_1879 = (v_90 | ~v_89) ;
	assign x_1877 = (v_91 | v_75) ;
	assign x_1876 = (v_92 | v_63) ;
	assign x_1875 = (v_92 | v_60) ;
	assign x_1874 = (((((v_78 | ~v_92) | ~v_91) | ~v_90) | ~v_86) | v_93) ;
	assign x_1873 = (v_94 | v_76) ;
	assign x_1872 = (v_94 | v_79) ;
	assign x_1871 = (v_95 | v_51) ;
	assign x_1870 = (v_95 | v_59) ;
	assign x_1869 = (((v_74 | ~v_95) | ~v_94) | v_96) ;
	assign x_1868 = (v_97 | v_77) ;
	assign x_1867 = (v_97 | ~v_96) ;
	assign x_1866 = (v_98 | v_63) ;
	assign x_1865 = (v_98 | v_79) ;
	assign x_1864 = (v_99 | v_50) ;
	assign x_1862 = (((v_59 | ~v_99) | ~v_98) | v_100) ;
	assign x_1861 = (v_101 | v_64) ;
	assign x_1860 = (v_101 | ~v_100) ;
	assign x_1859 = (v_102 | v_74) ;
	assign x_1858 = (v_102 | v_77) ;
	assign x_1857 = (v_103 | v_64) ;
	assign x_1856 = (v_103 | v_59) ;
	assign x_1855 = (((((v_79 | ~v_103) | ~v_102) | ~v_101) | ~v_97) | v_104) ;
	assign x_1854 = (v_105 | ~v_104) ;
	assign x_1853 = (v_105 | ~v_93) ;
	assign x_1852 = (((v_78 | ~v_92) | ~v_91) | v_106) ;
	assign x_1851 = (v_107 | v_74) ;
	assign x_1850 = (v_107 | ~v_106) ;
	assign x_1849 = (v_108 | v_51) ;
	assign x_1847 = (((((v_76 | ~v_88) | ~v_87) | ~v_108) | ~v_107) | v_109) ;
	assign x_1846 = (v_110 | v_78) ;
	assign x_1845 = (v_110 | v_77) ;
	assign x_1844 = (v_111 | v_50) ;
	assign x_1843 = (v_111 | v_60) ;
	assign x_1842 = (((v_75 | ~v_111) | ~v_110) | v_112) ;
	assign x_1841 = (v_113 | v_79) ;
	assign x_1840 = (v_113 | ~v_112) ;
	assign x_1839 = (v_114 | v_63) ;
	assign x_1838 = (v_114 | v_77) ;
	assign x_1837 = (v_115 | v_59) ;
	assign x_1836 = (v_115 | v_75) ;
	assign x_1835 = (((v_50 | ~v_115) | ~v_114) | v_116) ;
	assign x_1834 = (v_117 | v_64) ;
	assign x_1832 = (v_118 | v_79) ;
	assign x_1831 = (v_118 | v_75) ;
	assign x_1830 = (v_119 | v_50) ;
	assign x_1829 = (v_119 | v_64) ;
	assign x_1828 = (((((v_77 | ~v_119) | ~v_118) | ~v_117) | ~v_113) | v_120) ;
	assign x_1827 = (v_121 | ~v_120) ;
	assign x_1826 = (v_121 | ~v_109) ;
	assign x_1825 = (v_122 | v_59) ;
	assign x_1824 = (v_122 | ~v_106) ;
	assign x_1823 = (v_123 | v_50) ;
	assign x_1822 = (v_123 | ~v_89) ;
	assign x_1821 = (((((v_63 | ~v_84) | ~v_123) | ~v_83) | ~v_122) | v_124) ;
	assign x_1820 = (v_125 | v_64) ;
	assign x_1819 = (v_125 | v_78) ;
	assign x_1817 = (v_126 | v_75) ;
	assign x_1816 = (((v_60 | ~v_126) | ~v_125) | v_127) ;
	assign x_1815 = (v_128 | v_79) ;
	assign x_1814 = (v_128 | ~v_127) ;
	assign x_1813 = (v_129 | v_60) ;
	assign x_1812 = (v_129 | v_74) ;
	assign x_1811 = (v_130 | v_76) ;
	assign x_1810 = (v_130 | v_64) ;
	assign x_1809 = (((v_51 | ~v_130) | ~v_129) | v_131) ;
	assign x_1808 = (v_132 | v_77) ;
	assign x_1807 = (v_132 | ~v_131) ;
	assign x_1806 = (v_133 | v_60) ;
	assign x_1805 = (v_133 | v_79) ;
	assign x_1804 = (v_134 | v_51) ;
	assign x_1802 = (((((v_64 | ~v_134) | ~v_133) | ~v_132) | ~v_128) | v_135) ;
	assign x_1801 = (v_136 | ~v_135) ;
	assign x_1800 = (v_136 | ~v_124) ;
	assign x_1799 = ((((v_65 | ~v_136) | ~v_121) | ~v_105) | v_137) ;
	assign x_1798 = (((v_79 | ~v_103) | ~v_102) | v_138) ;
	assign x_1797 = (v_139 | v_76) ;
	assign x_1796 = (v_139 | ~v_138) ;
	assign x_1795 = (v_140 | v_51) ;
	assign x_1794 = (v_140 | ~v_100) ;
	assign x_1793 = (((((v_74 | ~v_95) | ~v_94) | ~v_140) | ~v_139) | v_141) ;
	assign x_1792 = (((v_77 | ~v_119) | ~v_118) | v_142) ;
	assign x_1791 = (v_143 | v_78) ;
	assign x_1790 = (v_143 | ~v_142) ;
	assign x_1789 = (v_144 | v_60) ;
	assign x_1787 = (((((v_75 | ~v_111) | ~v_110) | ~v_144) | ~v_143) | v_145) ;
	assign x_1786 = (v_146 | ~v_145) ;
	assign x_1785 = (v_146 | ~v_141) ;
	assign x_1784 = (v_147 | v_63) ;
	assign x_1783 = (v_147 | ~v_138) ;
	assign x_1782 = (v_148 | v_50) ;
	assign x_1780 = (((((v_59 | ~v_99) | ~v_98) | ~v_148) | ~v_147) | v_149) ;
	assign x_1779 = (((v_64 | ~v_134) | ~v_133) | v_150) ;
	assign x_1778 = (v_151 | v_78) ;
	assign x_1777 = (v_151 | ~v_150) ;
	assign x_1776 = (v_152 | v_75) ;
	assign x_1775 = (v_152 | ~v_131) ;
	assign x_1773 = (v_154 | ~v_153) ;
	assign x_1772 = (v_154 | ~v_149) ;
	assign x_1771 = ((((v_61 | ~v_154) | ~v_146) | ~v_105) | v_155) ;
	assign x_1770 = (v_156 | v_63) ;
	assign x_1769 = (v_156 | ~v_142) ;
	assign x_1768 = (v_157 | v_59) ;
	assign x_1767 = (v_157 | ~v_112) ;
	assign x_1766 = (((((v_50 | ~v_115) | ~v_114) | ~v_157) | ~v_156) | v_158) ;
	assign x_1765 = (v_159 | v_76) ;
	assign x_1764 = (v_159 | ~v_150) ;
	assign x_1763 = (v_160 | v_74) ;
	assign x_1762 = (v_160 | ~v_127) ;
	assign x_1761 = (((((v_51 | ~v_130) | ~v_129) | ~v_160) | ~v_159) | v_161) ;
	assign x_1760 = (v_162 | ~v_161) ;
	assign x_1758 = ((((v_52 | ~v_162) | ~v_146) | ~v_121) | v_163) ;
	assign x_1757 = ((((v_14 | ~v_162) | ~v_154) | ~v_136) | v_164) ;
	assign x_1756 = (v_165 | ~v_164) ;
	assign x_1755 = (v_165 | ~v_163) ;
	assign x_1754 = (v_165 | ~v_155) ;
	assign x_1753 = (v_165 | ~v_137) ;
	assign x_1752 = (v_166 | v_1) ;
	assign x_1751 = (v_166 | ~v_78) ;
	assign x_1750 = (v_167 | v_16) ;
	assign x_1749 = (v_167 | ~v_79) ;
	assign x_1748 = (v_168 | v_5) ;
	assign x_1747 = (v_168 | v_78) ;
	assign x_1746 = (v_169 | v_17) ;
	assign x_1745 = (v_169 | ~v_65) ;
	assign x_1743 = (v_170 | v_65) ;
	assign x_1742 = (v_171 | v_18) ;
	assign x_1741 = (v_171 | v_61) ;
	assign x_1740 = (v_172 | v_19) ;
	assign x_1739 = (v_172 | v_79) ;
	assign x_1738 = (v_173 | v_15) ;
	assign x_1737 = (v_173 | ~v_61) ;
	assign x_1736 = (((((((((((((((v_13 | v_10) | v_68) | v_49) | v_48) | v_62) | v_47) | ~v_173) | ~v_172) | ~v_171) | ~v_170) | ~v_169) | ~v_168) | ~v_167) | ~v_166) | v_174) ;
	assign x_1735 = (v_175 | v_2) ;
	assign x_1734 = (v_175 | ~v_78) ;
	assign x_1733 = (v_176 | v_29) ;
	assign x_1732 = (v_176 | ~v_79) ;
	assign x_1731 = (v_177 | v_4) ;
	assign x_1730 = (v_177 | v_78) ;
	assign x_1728 = (v_178 | v_79) ;
	assign x_1727 = (v_179 | v_30) ;
	assign x_1726 = (v_179 | ~v_65) ;
	assign x_1725 = (v_180 | v_33) ;
	assign x_1724 = (v_180 | v_65) ;
	assign x_1723 = (v_181 | v_31) ;
	assign x_1721 = (v_182 | v_28) ;
	assign x_1720 = (v_182 | ~v_61) ;
	assign x_1719 = (((((((((((((((v_24 | v_27) | v_54) | v_53) | v_55) | v_66) | v_70) | ~v_182) | ~v_181) | ~v_180) | ~v_179) | ~v_178) | ~v_177) | ~v_176) | ~v_175) | v_183) ;
	assign x_1718 = (v_184 | v_3) ;
	assign x_1717 = (v_184 | ~v_78) ;
	assign x_1716 = (v_185 | ~v_79) ;
	assign x_1714 = (v_186 | v_6) ;
	assign x_1713 = (v_186 | v_78) ;
	assign x_1712 = (v_187 | v_45) ;
	assign x_1711 = (v_187 | v_79) ;
	assign x_1710 = (v_188 | ~v_65) ;
	assign x_1709 = (v_188 | v_43) ;
	assign x_1708 = (v_189 | v_46) ;
	assign x_1707 = (v_189 | v_65) ;
	assign x_1706 = (v_190 | v_61) ;
	assign x_1705 = (v_190 | v_44) ;
	assign x_1704 = (v_191 | ~v_61) ;
	assign x_1703 = (v_191 | v_41) ;
	assign x_1702 = (((((((((((((((v_37 | v_56) | v_67) | v_40) | v_58) | v_57) | v_72) | ~v_191) | ~v_190) | ~v_189) | ~v_188) | ~v_187) | ~v_186) | ~v_185) | ~v_184) | v_192) ;
	assign x_1701 = (v_193 | ~v_192) ;
	assign x_1699 = (v_193 | ~v_174) ;
	assign x_1698 = (v_194 | v_1) ;
	assign x_1697 = (v_194 | ~v_79) ;
	assign x_1696 = (v_195 | v_16) ;
	assign x_1695 = (v_195 | ~v_78) ;
	assign x_1694 = (v_196 | v_5) ;
	assign x_1693 = (v_196 | v_79) ;
	assign x_1692 = (v_197 | v_15) ;
	assign x_1691 = (v_197 | ~v_65) ;
	assign x_1690 = (v_198 | v_18) ;
	assign x_1689 = (v_198 | v_65) ;
	assign x_1688 = (v_199 | v_17) ;
	assign x_1687 = (v_199 | ~v_61) ;
	assign x_1686 = (v_200 | v_20) ;
	assign x_1684 = (v_201 | v_19) ;
	assign x_1683 = (v_201 | v_78) ;
	assign x_1682 = (((((((((((((((v_12 | v_11) | v_69) | v_68) | v_48) | v_47) | v_80) | ~v_201) | ~v_200) | ~v_199) | ~v_198) | ~v_197) | ~v_196) | ~v_195) | ~v_194) | v_202) ;
	assign x_1681 = (v_203 | v_2) ;
	assign x_1680 = (v_203 | ~v_79) ;
	assign x_1679 = (v_204 | v_29) ;
	assign x_1678 = (v_204 | ~v_78) ;
	assign x_1677 = (v_205 | v_4) ;
	assign x_1676 = (v_205 | v_79) ;
	assign x_1675 = (v_206 | v_32) ;
	assign x_1674 = (v_206 | v_78) ;
	assign x_1673 = (v_207 | v_28) ;
	assign x_1672 = (v_207 | ~v_65) ;
	assign x_1671 = (v_208 | v_31) ;
	assign x_1669 = (v_209 | v_30) ;
	assign x_1668 = (v_209 | ~v_61) ;
	assign x_1667 = (v_210 | v_33) ;
	assign x_1666 = (v_210 | v_61) ;
	assign x_1665 = (((((((((((((((v_25 | v_26) | v_54) | v_53) | v_81) | v_71) | v_70) | ~v_210) | ~v_209) | ~v_208) | ~v_207) | ~v_206) | ~v_205) | ~v_204) | ~v_203) | v_211) ;
	assign x_1664 = (v_212 | v_3) ;
	assign x_1662 = (v_213 | ~v_78) ;
	assign x_1661 = (v_213 | v_42) ;
	assign x_1660 = (v_214 | v_6) ;
	assign x_1659 = (v_214 | v_79) ;
	assign x_1658 = (v_215 | v_45) ;
	assign x_1657 = (v_215 | v_78) ;
	assign x_1655 = (v_216 | v_41) ;
	assign x_1654 = (v_217 | v_65) ;
	assign x_1653 = (v_217 | v_44) ;
	assign x_1652 = (v_218 | ~v_61) ;
	assign x_1651 = (v_218 | v_43) ;
	assign x_1650 = (v_219 | v_61) ;
	assign x_1649 = (v_219 | v_46) ;
	assign x_1648 = (((((((((((((((v_39 | v_38) | v_56) | v_57) | v_73) | v_72) | v_82) | ~v_219) | ~v_218) | ~v_217) | ~v_216) | ~v_215) | ~v_214) | ~v_213) | ~v_212) | v_220) ;
	assign x_1647 = (v_221 | ~v_220) ;
	assign x_1646 = (v_221 | ~v_211) ;
	assign x_1645 = (v_221 | ~v_202) ;
	assign x_1644 = (v_222 | v_1) ;
	assign x_1643 = (v_222 | ~v_76) ;
	assign x_1642 = (v_223 | v_16) ;
	assign x_1640 = (v_224 | v_5) ;
	assign x_1639 = (v_224 | v_76) ;
	assign x_1638 = (v_225 | v_18) ;
	assign x_1637 = (v_225 | v_52) ;
	assign x_1636 = (v_226 | v_19) ;
	assign x_1635 = (v_226 | v_77) ;
	assign x_1634 = (v_227 | v_15) ;
	assign x_1633 = (v_227 | ~v_52) ;
	assign x_1632 = (((((((((((((((v_13 | v_12) | v_10) | v_68) | v_48) | v_62) | v_47) | ~v_227) | ~v_226) | ~v_225) | ~v_170) | ~v_169) | ~v_224) | ~v_223) | ~v_222) | v_228) ;
	assign x_1631 = (v_229 | v_2) ;
	assign x_1630 = (v_229 | ~v_76) ;
	assign x_1629 = (v_230 | v_29) ;
	assign x_1628 = (v_230 | ~v_77) ;
	assign x_1627 = (v_231 | v_4) ;
	assign x_1625 = (v_232 | v_32) ;
	assign x_1624 = (v_232 | v_77) ;
	assign x_1623 = (v_233 | v_28) ;
	assign x_1622 = (v_233 | ~v_52) ;
	assign x_1621 = (v_234 | v_31) ;
	assign x_1620 = (v_234 | v_52) ;
	assign x_1619 = (((((((((((((((v_24 | v_27) | v_26) | v_54) | v_53) | v_66) | v_70) | ~v_234) | ~v_233) | ~v_180) | ~v_179) | ~v_232) | ~v_231) | ~v_230) | ~v_229) | v_235) ;
	assign x_1618 = (v_236 | v_3) ;
	assign x_1617 = (v_236 | ~v_76) ;
	assign x_1616 = (v_237 | ~v_77) ;
	assign x_1615 = (v_237 | v_42) ;
	assign x_1614 = (v_238 | v_6) ;
	assign x_1613 = (v_238 | v_76) ;
	assign x_1612 = (v_239 | v_45) ;
	assign x_1610 = (v_240 | ~v_52) ;
	assign x_1609 = (v_240 | v_41) ;
	assign x_1608 = (v_241 | v_52) ;
	assign x_1607 = (v_241 | v_44) ;
	assign x_1606 = (((((((((((((((v_39 | v_37) | v_56) | v_67) | v_40) | v_57) | v_72) | ~v_241) | ~v_240) | ~v_189) | ~v_188) | ~v_239) | ~v_238) | ~v_237) | ~v_236) | v_242) ;
	assign x_1605 = (v_243 | ~v_242) ;
	assign x_1603 = (v_243 | ~v_228) ;
	assign x_1602 = (v_244 | v_1) ;
	assign x_1601 = (v_244 | ~v_77) ;
	assign x_1600 = (v_245 | v_16) ;
	assign x_1599 = (v_245 | ~v_76) ;
	assign x_1598 = (v_246 | v_5) ;
	assign x_1596 = (v_247 | v_17) ;
	assign x_1595 = (v_247 | ~v_52) ;
	assign x_1594 = (v_248 | v_20) ;
	assign x_1593 = (v_248 | v_52) ;
	assign x_1592 = (v_249 | v_19) ;
	assign x_1591 = (v_249 | v_76) ;
	assign x_1590 = (((((((((((((((v_13 | v_12) | v_11) | v_68) | v_48) | v_47) | v_80) | ~v_249) | ~v_248) | ~v_247) | ~v_198) | ~v_197) | ~v_246) | ~v_245) | ~v_244) | v_250) ;
	assign x_1589 = (v_251 | v_2) ;
	assign x_1588 = (v_251 | ~v_77) ;
	assign x_1587 = (v_252 | v_29) ;
	assign x_1586 = (v_252 | ~v_76) ;
	assign x_1585 = (v_253 | v_4) ;
	assign x_1584 = (v_253 | v_77) ;
	assign x_1583 = (v_254 | v_32) ;
	assign x_1581 = (v_255 | v_30) ;
	assign x_1580 = (v_255 | ~v_52) ;
	assign x_1579 = (v_256 | v_33) ;
	assign x_1578 = (v_256 | v_52) ;
	assign x_1577 = (((((((((((((((v_25 | v_27) | v_26) | v_54) | v_53) | v_81) | v_70) | ~v_256) | ~v_255) | ~v_208) | ~v_207) | ~v_254) | ~v_253) | ~v_252) | ~v_251) | v_257) ;
	assign x_1576 = (v_258 | v_3) ;
	assign x_1575 = (v_258 | ~v_77) ;
	assign x_1574 = (v_259 | ~v_76) ;
	assign x_1573 = (v_259 | v_42) ;
	assign x_1572 = (v_260 | v_6) ;
	assign x_1571 = (v_260 | v_77) ;
	assign x_1570 = (v_261 | ~v_52) ;
	assign x_1569 = (v_261 | v_43) ;
	assign x_1568 = (v_262 | v_52) ;
	assign x_1566 = (v_263 | v_76) ;
	assign x_1565 = (v_263 | v_45) ;
	assign x_1564 = (((((((((((((((v_39 | v_38) | v_56) | v_40) | v_57) | v_72) | v_82) | ~v_263) | ~v_262) | ~v_261) | ~v_217) | ~v_216) | ~v_260) | ~v_259) | ~v_258) | v_264) ;
	assign x_1563 = (v_265 | ~v_264) ;
	assign x_1562 = (v_265 | ~v_257) ;
	assign x_1561 = (v_265 | ~v_250) ;
	assign x_1560 = (v_266 | v_1) ;
	assign x_1559 = (v_266 | ~v_74) ;
	assign x_1558 = (v_267 | v_5) ;
	assign x_1557 = (v_267 | v_74) ;
	assign x_1556 = (v_268 | v_19) ;
	assign x_1555 = (v_268 | v_75) ;
	assign x_1554 = (v_269 | v_16) ;
	assign x_1553 = (v_269 | ~v_75) ;
	assign x_1551 = (v_271 | v_2) ;
	assign x_1550 = (v_271 | ~v_74) ;
	assign x_1549 = (v_272 | v_4) ;
	assign x_1548 = (v_272 | v_74) ;
	assign x_1547 = (v_273 | v_32) ;
	assign x_1546 = (v_273 | v_75) ;
	assign x_1544 = (v_274 | ~v_75) ;
	assign x_1543 = (((((((((((((((v_25 | v_24) | v_27) | v_54) | v_53) | v_55) | v_70) | ~v_274) | ~v_273) | ~v_234) | ~v_233) | ~v_210) | ~v_209) | ~v_272) | ~v_271) | v_275) ;
	assign x_1542 = (v_276 | v_3) ;
	assign x_1541 = (v_276 | ~v_74) ;
	assign x_1540 = (v_277 | ~v_75) ;
	assign x_1539 = (v_277 | v_42) ;
	assign x_1537 = (v_278 | v_74) ;
	assign x_1536 = (v_279 | v_45) ;
	assign x_1535 = (v_279 | v_75) ;
	assign x_1534 = (((((((((((((((v_38 | v_37) | v_56) | v_40) | v_58) | v_57) | v_72) | ~v_279) | ~v_241) | ~v_240) | ~v_219) | ~v_218) | ~v_278) | ~v_277) | ~v_276) | v_280) ;
	assign x_1533 = (v_281 | ~v_280) ;
	assign x_1532 = (v_281 | ~v_275) ;
	assign x_1531 = (v_281 | ~v_270) ;
	assign x_1530 = (v_282 | v_1) ;
	assign x_1529 = (v_282 | ~v_63) ;
	assign x_1528 = (v_283 | v_16) ;
	assign x_1527 = (v_283 | ~v_64) ;
	assign x_1526 = (v_284 | v_5) ;
	assign x_1525 = (v_284 | v_63) ;
	assign x_1524 = (v_285 | v_19) ;
	assign x_1522 = (v_286 | v_18) ;
	assign x_1521 = (v_286 | v_14) ;
	assign x_1520 = (v_287 | ~v_14) ;
	assign x_1519 = (v_287 | v_15) ;
	assign x_1518 = (((((((((((((((v_13 | v_8) | v_12) | v_10) | v_48) | v_62) | v_47) | ~v_287) | ~v_286) | ~v_170) | ~v_169) | ~v_285) | ~v_284) | ~v_283) | ~v_282) | v_288) ;
	assign x_1517 = (v_289 | v_2) ;
	assign x_1516 = (v_289 | ~v_63) ;
	assign x_1515 = (v_290 | v_29) ;
	assign x_1514 = (v_290 | ~v_64) ;
	assign x_1513 = (v_291 | v_4) ;
	assign x_1512 = (v_291 | v_63) ;
	assign x_1511 = (v_292 | v_32) ;
	assign x_1510 = (v_292 | v_64) ;
	assign x_1509 = (v_293 | ~v_14) ;
	assign x_1507 = (v_294 | v_14) ;
	assign x_1506 = (v_294 | v_31) ;
	assign x_1505 = (((((((((((((((v_24 | v_22) | v_27) | v_26) | v_54) | v_53) | v_66) | ~v_294) | ~v_293) | ~v_180) | ~v_179) | ~v_292) | ~v_291) | ~v_290) | ~v_289) | v_295) ;
	assign x_1504 = (v_296 | v_3) ;
	assign x_1503 = (v_296 | ~v_63) ;
	assign x_1502 = (v_297 | ~v_64) ;
	assign x_1501 = (v_297 | v_42) ;
	assign x_1500 = (v_298 | v_45) ;
	assign x_1499 = (v_298 | v_64) ;
	assign x_1498 = (v_299 | ~v_14) ;
	assign x_1497 = (v_299 | v_41) ;
	assign x_1496 = (v_300 | v_14) ;
	assign x_1495 = (v_300 | v_44) ;
	assign x_1494 = (v_301 | v_6) ;
	assign x_1492 = (((((((((((((((v_39 | v_35) | v_37) | v_56) | v_67) | v_40) | v_57) | ~v_301) | ~v_300) | ~v_299) | ~v_189) | ~v_188) | ~v_298) | ~v_297) | ~v_296) | v_302) ;
	assign x_1491 = (v_303 | ~v_302) ;
	assign x_1490 = (v_303 | ~v_295) ;
	assign x_1489 = (v_303 | ~v_288) ;
	assign x_1488 = (v_304 | v_1) ;
	assign x_1487 = (v_304 | ~v_65) ;
	assign x_1485 = (v_305 | ~v_65) ;
	assign x_1484 = (v_306 | v_5) ;
	assign x_1483 = (v_306 | v_65) ;
	assign x_1482 = (v_307 | v_19) ;
	assign x_1481 = (v_307 | v_65) ;
	assign x_1480 = (((((((((((((((v_13 | v_7) | v_12) | v_68) | v_48) | v_62) | v_80) | ~v_198) | ~v_197) | ~v_307) | ~v_306) | ~v_305) | ~v_304) | ~v_170) | ~v_169) | v_308) ;
	assign x_1478 = (v_309 | ~v_65) ;
	assign x_1477 = (v_310 | v_29) ;
	assign x_1476 = (v_310 | ~v_65) ;
	assign x_1475 = (v_311 | v_4) ;
	assign x_1474 = (v_311 | v_65) ;
	assign x_1473 = (v_312 | v_32) ;
	assign x_1472 = (v_312 | v_65) ;
	assign x_1471 = (((((((((((((((v_21 | v_27) | v_26) | v_54) | v_81) | v_66) | v_70) | ~v_208) | ~v_207) | ~v_312) | ~v_311) | ~v_310) | ~v_309) | ~v_180) | ~v_179) | v_313) ;
	assign x_1470 = (v_314 | v_3) ;
	assign x_1469 = (v_314 | ~v_65) ;
	assign x_1468 = (v_315 | ~v_65) ;
	assign x_1467 = (v_315 | v_42) ;
	assign x_1466 = (v_316 | v_45) ;
	assign x_1465 = (v_316 | v_65) ;
	assign x_1463 = (v_317 | v_65) ;
	assign x_1462 = (((((((((((((((v_39 | v_34) | v_67) | v_40) | v_57) | v_72) | v_82) | ~v_317) | ~v_217) | ~v_216) | ~v_316) | ~v_315) | ~v_314) | ~v_189) | ~v_188) | v_318) ;
	assign x_1461 = (v_319 | ~v_318) ;
	assign x_1460 = (v_319 | ~v_313) ;
	assign x_1459 = (v_319 | ~v_308) ;
	assign x_1458 = (v_320 | v_1) ;
	assign x_1457 = (v_320 | ~v_64) ;
	assign x_1456 = (v_321 | v_16) ;
	assign x_1455 = (v_321 | ~v_63) ;
	assign x_1454 = (v_322 | v_5) ;
	assign x_1453 = (v_322 | v_64) ;
	assign x_1452 = (v_323 | v_19) ;
	assign x_1451 = (v_323 | v_63) ;
	assign x_1450 = (v_324 | ~v_14) ;
	assign x_1448 = (v_325 | v_20) ;
	assign x_1447 = (v_325 | v_14) ;
	assign x_1446 = (((((((((((((((v_13 | v_9) | v_12) | v_11) | v_68) | v_47) | v_80) | ~v_325) | ~v_324) | ~v_323) | ~v_322) | ~v_198) | ~v_321) | ~v_320) | ~v_197) | v_326) ;
	assign x_1445 = (v_327 | v_2) ;
	assign x_1444 = (v_327 | ~v_64) ;
	assign x_1443 = (v_328 | v_29) ;
	assign x_1442 = (v_328 | ~v_63) ;
	assign x_1441 = (v_329 | v_4) ;
	assign x_1440 = (v_329 | v_64) ;
	assign x_1439 = (v_330 | v_32) ;
	assign x_1438 = (v_330 | v_63) ;
	assign x_1437 = (v_331 | ~v_14) ;
	assign x_1436 = (v_331 | v_30) ;
	assign x_1435 = (v_332 | v_14) ;
	assign x_1433 = (((((((((((((((v_25 | v_23) | v_27) | v_26) | v_53) | v_81) | v_70) | ~v_332) | ~v_331) | ~v_330) | ~v_329) | ~v_208) | ~v_328) | ~v_327) | ~v_207) | v_333) ;
	assign x_1432 = (v_334 | v_3) ;
	assign x_1431 = (v_334 | ~v_64) ;
	assign x_1430 = (v_335 | ~v_63) ;
	assign x_1429 = (v_335 | v_42) ;
	assign x_1428 = (v_336 | v_45) ;
	assign x_1426 = (v_337 | ~v_14) ;
	assign x_1425 = (v_337 | v_43) ;
	assign x_1424 = (v_338 | v_14) ;
	assign x_1423 = (v_338 | v_46) ;
	assign x_1422 = (v_339 | v_6) ;
	assign x_1421 = (v_339 | v_64) ;
	assign x_1419 = (v_341 | ~v_340) ;
	assign x_1418 = (v_341 | ~v_333) ;
	assign x_1417 = (v_341 | ~v_326) ;
	assign x_1416 = (v_342 | v_16) ;
	assign x_1415 = (v_342 | ~v_60) ;
	assign x_1414 = (v_343 | v_1) ;
	assign x_1413 = (v_343 | ~v_59) ;
	assign x_1412 = (v_344 | v_5) ;
	assign x_1411 = (v_344 | v_59) ;
	assign x_1410 = (v_345 | v_19) ;
	assign x_1409 = (v_345 | v_60) ;
	assign x_1408 = (((((((((((((((v_13 | v_8) | v_12) | v_11) | v_10) | v_48) | v_47) | ~v_345) | ~v_344) | ~v_287) | ~v_343) | ~v_342) | ~v_286) | ~v_200) | ~v_199) | v_346) ;
	assign x_1407 = (v_347 | v_29) ;
	assign x_1406 = (v_347 | ~v_60) ;
	assign x_1404 = (v_348 | v_59) ;
	assign x_1403 = (v_349 | v_2) ;
	assign x_1402 = (v_349 | ~v_59) ;
	assign x_1401 = (v_350 | v_32) ;
	assign x_1400 = (v_350 | v_60) ;
	assign x_1399 = (((((((((((((((v_25 | v_24) | v_22) | v_27) | v_26) | v_54) | v_53) | ~v_350) | ~v_349) | ~v_348) | ~v_294) | ~v_293) | ~v_210) | ~v_209) | ~v_347) | v_351) ;
	assign x_1398 = (v_352 | ~v_60) ;
	assign x_1397 = (v_352 | v_42) ;
	assign x_1396 = (v_353 | v_6) ;
	assign x_1395 = (v_353 | v_59) ;
	assign x_1394 = (v_354 | v_3) ;
	assign x_1393 = (v_354 | ~v_59) ;
	assign x_1392 = (v_355 | v_45) ;
	assign x_1391 = (v_355 | v_60) ;
	assign x_1389 = (v_357 | ~v_356) ;
	assign x_1388 = (v_357 | ~v_351) ;
	assign x_1387 = (v_357 | ~v_346) ;
	assign x_1386 = (v_358 | v_16) ;
	assign x_1385 = (v_358 | ~v_61) ;
	assign x_1384 = (v_359 | v_19) ;
	assign x_1383 = (v_359 | v_61) ;
	assign x_1382 = (v_360 | v_1) ;
	assign x_1381 = (v_360 | ~v_61) ;
	assign x_1380 = (v_361 | v_5) ;
	assign x_1379 = (v_361 | v_61) ;
	assign x_1378 = (((((((((((((((v_13 | v_7) | v_12) | v_11) | v_10) | v_68) | v_48) | ~v_173) | ~v_361) | ~v_360) | ~v_171) | ~v_359) | ~v_358) | ~v_200) | ~v_199) | v_362) ;
	assign x_1377 = (v_363 | v_29) ;
	assign x_1376 = (v_363 | ~v_61) ;
	assign x_1374 = (v_364 | v_61) ;
	assign x_1373 = (v_365 | v_2) ;
	assign x_1372 = (v_365 | ~v_61) ;
	assign x_1371 = (v_366 | v_4) ;
	assign x_1370 = (v_366 | v_61) ;
	assign x_1369 = (((((((((((((((v_25 | v_24) | v_21) | v_27) | v_26) | v_54) | v_70) | ~v_182) | ~v_366) | ~v_365) | ~v_181) | ~v_364) | ~v_363) | ~v_210) | ~v_209) | v_367) ;
	assign x_1368 = (v_368 | ~v_61) ;
	assign x_1367 = (v_368 | v_42) ;
	assign x_1366 = (v_369 | v_61) ;
	assign x_1365 = (v_369 | v_45) ;
	assign x_1364 = (v_370 | v_3) ;
	assign x_1363 = (v_370 | ~v_61) ;
	assign x_1362 = (v_371 | v_6) ;
	assign x_1361 = (v_371 | v_61) ;
	assign x_1359 = (v_373 | ~v_372) ;
	assign x_1358 = (v_373 | ~v_367) ;
	assign x_1357 = (v_373 | ~v_362) ;
	assign x_1356 = (v_374 | v_19) ;
	assign x_1355 = (v_374 | v_59) ;
	assign x_1354 = (v_375 | v_16) ;
	assign x_1353 = (v_375 | ~v_59) ;
	assign x_1352 = (v_376 | v_1) ;
	assign x_1351 = (v_376 | ~v_60) ;
	assign x_1350 = (v_377 | v_5) ;
	assign x_1349 = (v_377 | v_60) ;
	assign x_1348 = (((((((((((((((v_13 | v_9) | v_12) | v_11) | v_10) | v_68) | v_47) | ~v_377) | ~v_376) | ~v_375) | ~v_173) | ~v_325) | ~v_171) | ~v_324) | ~v_374) | v_378) ;
	assign x_1347 = (v_379 | v_29) ;
	assign x_1346 = (v_379 | ~v_59) ;
	assign x_1344 = (v_380 | v_59) ;
	assign x_1343 = (v_381 | v_2) ;
	assign x_1342 = (v_381 | ~v_60) ;
	assign x_1341 = (v_382 | v_4) ;
	assign x_1340 = (v_382 | v_60) ;
	assign x_1339 = (((((((((((((((v_25 | v_24) | v_23) | v_27) | v_26) | v_53) | v_70) | ~v_382) | ~v_381) | ~v_182) | ~v_181) | ~v_332) | ~v_331) | ~v_380) | ~v_379) | v_383) ;
	assign x_1338 = (v_384 | v_45) ;
	assign x_1337 = (v_384 | v_59) ;
	assign x_1336 = (v_385 | ~v_59) ;
	assign x_1335 = (v_385 | v_42) ;
	assign x_1334 = (v_386 | v_3) ;
	assign x_1333 = (v_386 | ~v_60) ;
	assign x_1332 = (v_387 | v_6) ;
	assign x_1331 = (v_387 | v_60) ;
	assign x_1329 = (v_389 | ~v_388) ;
	assign x_1328 = (v_389 | ~v_383) ;
	assign x_1327 = (v_389 | ~v_378) ;
	assign x_1326 = (v_390 | v_1) ;
	assign x_1325 = (v_390 | ~v_50) ;
	assign x_1324 = (v_391 | v_16) ;
	assign x_1323 = (v_391 | ~v_51) ;
	assign x_1322 = (v_392 | v_5) ;
	assign x_1321 = (v_392 | v_50) ;
	assign x_1320 = (v_393 | v_19) ;
	assign x_1319 = (v_393 | v_51) ;
	assign x_1318 = (((((((((((((((v_13 | v_8) | v_11) | v_10) | v_49) | v_48) | v_47) | ~v_393) | ~v_287) | ~v_286) | ~v_248) | ~v_247) | ~v_392) | ~v_391) | ~v_390) | v_394) ;
	assign x_1317 = (v_395 | v_2) ;
	assign x_1316 = (v_395 | ~v_50) ;
	assign x_1314 = (v_396 | ~v_51) ;
	assign x_1313 = (v_397 | v_4) ;
	assign x_1312 = (v_397 | v_50) ;
	assign x_1311 = (v_398 | v_32) ;
	assign x_1310 = (v_398 | v_51) ;
	assign x_1309 = (((((((((((((((v_25 | v_24) | v_22) | v_27) | v_54) | v_53) | v_55) | ~v_398) | ~v_256) | ~v_255) | ~v_294) | ~v_293) | ~v_397) | ~v_396) | ~v_395) | v_399) ;
	assign x_1307 = (v_400 | ~v_50) ;
	assign x_1306 = (v_401 | ~v_51) ;
	assign x_1305 = (v_401 | v_42) ;
	assign x_1304 = (v_402 | v_6) ;
	assign x_1303 = (v_402 | v_50) ;
	assign x_1302 = (v_403 | v_51) ;
	assign x_1300 = (((((((((((((((v_38 | v_35) | v_37) | v_56) | v_40) | v_58) | v_57) | ~v_403) | ~v_402) | ~v_300) | ~v_262) | ~v_261) | ~v_299) | ~v_401) | ~v_400) | v_404) ;
	assign x_1299 = (v_405 | ~v_404) ;
	assign x_1298 = (v_405 | ~v_399) ;
	assign x_1297 = (v_405 | ~v_394) ;
	assign x_1296 = (v_406 | v_16) ;
	assign x_1295 = (v_406 | ~v_52) ;
	assign x_1294 = (v_407 | v_19) ;
	assign x_1293 = (v_407 | v_52) ;
	assign x_1292 = (v_408 | v_5) ;
	assign x_1291 = (v_408 | v_52) ;
	assign x_1290 = (v_409 | v_1) ;
	assign x_1289 = (v_409 | ~v_52) ;
	assign x_1288 = (((((((((((((((v_13 | v_7) | v_12) | v_11) | v_10) | v_68) | v_48) | ~v_409) | ~v_408) | ~v_227) | ~v_248) | ~v_247) | ~v_225) | ~v_407) | ~v_406) | v_410) ;
	assign x_1287 = (v_411 | v_29) ;
	assign x_1285 = (v_412 | v_4) ;
	assign x_1284 = (v_412 | v_52) ;
	assign x_1283 = (v_413 | v_2) ;
	assign x_1282 = (v_413 | ~v_52) ;
	assign x_1281 = (v_414 | v_32) ;
	assign x_1280 = (v_414 | v_52) ;
	assign x_1279 = (((((((((((((((v_25 | v_24) | v_21) | v_27) | v_26) | v_54) | v_70) | ~v_414) | ~v_413) | ~v_412) | ~v_234) | ~v_256) | ~v_255) | ~v_233) | ~v_411) | v_415) ;
	assign x_1278 = (v_416 | ~v_52) ;
	assign x_1277 = (v_416 | v_42) ;
	assign x_1276 = (v_417 | v_52) ;
	assign x_1275 = (v_417 | v_45) ;
	assign x_1274 = (v_418 | v_6) ;
	assign x_1273 = (v_418 | v_52) ;
	assign x_1272 = (v_419 | v_3) ;
	assign x_1270 = (((((((((((((((v_39 | v_38) | v_37) | v_34) | v_40) | v_57) | v_72) | ~v_419) | ~v_418) | ~v_262) | ~v_261) | ~v_241) | ~v_240) | ~v_417) | ~v_416) | v_420) ;
	assign x_1269 = (v_421 | ~v_420) ;
	assign x_1268 = (v_421 | ~v_415) ;
	assign x_1267 = (v_421 | ~v_410) ;
	assign x_1266 = (v_422 | v_16) ;
	assign x_1265 = (v_422 | ~v_50) ;
	assign x_1264 = (v_423 | v_19) ;
	assign x_1263 = (v_423 | v_50) ;
	assign x_1262 = (v_424 | v_1) ;
	assign x_1261 = (v_424 | ~v_51) ;
	assign x_1260 = (v_425 | v_5) ;
	assign x_1259 = (v_425 | v_51) ;
	assign x_1258 = (((((((((((((((v_9 | v_12) | v_11) | v_10) | v_69) | v_68) | v_47) | ~v_425) | ~v_424) | ~v_423) | ~v_227) | ~v_325) | ~v_324) | ~v_225) | ~v_422) | v_426) ;
	assign x_1257 = (v_427 | v_29) ;
	assign x_1255 = (v_428 | v_32) ;
	assign x_1254 = (v_428 | v_50) ;
	assign x_1253 = (v_429 | v_2) ;
	assign x_1252 = (v_429 | ~v_51) ;
	assign x_1251 = (v_430 | v_4) ;
	assign x_1250 = (v_430 | v_51) ;
	assign x_1248 = (v_432 | ~v_50) ;
	assign x_1247 = (v_432 | v_42) ;
	assign x_1246 = (v_433 | v_50) ;
	assign x_1245 = (v_433 | v_45) ;
	assign x_1244 = (v_434 | v_3) ;
	assign x_1243 = (v_434 | ~v_51) ;
	assign x_1241 = (v_435 | v_51) ;
	assign x_1240 = (((((((((((((((v_39 | v_38) | v_37) | v_36) | v_56) | v_73) | v_72) | ~v_435) | ~v_434) | ~v_338) | ~v_337) | ~v_433) | ~v_241) | ~v_432) | ~v_240) | v_436) ;
	assign x_1239 = (v_437 | ~v_436) ;
	assign x_1238 = (v_437 | ~v_431) ;
	assign x_1237 = (v_437 | ~v_426) ;
	assign x_1236 = (v_438 | ~v_14) ;
	assign x_1235 = (v_438 | v_16) ;
	assign x_1234 = (v_439 | v_19) ;
	assign x_1233 = (v_439 | v_14) ;
	assign x_1232 = (v_440 | ~v_14) ;
	assign x_1231 = (v_440 | v_1) ;
	assign x_1230 = (v_441 | v_5) ;
	assign x_1229 = (v_441 | v_14) ;
	assign x_1228 = (((((((((((((((v_13 | v_9) | v_7) | v_8) | v_12) | v_11) | v_10) | ~v_287) | ~v_441) | ~v_440) | ~v_286) | ~v_325) | ~v_439) | ~v_324) | ~v_438) | v_442) ;
	assign x_1226 = (v_443 | v_29) ;
	assign x_1225 = (v_444 | v_14) ;
	assign x_1224 = (v_444 | v_32) ;
	assign x_1223 = (v_445 | ~v_14) ;
	assign x_1222 = (v_445 | v_2) ;
	assign x_1221 = (v_446 | v_4) ;
	assign x_1220 = (v_446 | v_14) ;
	assign x_1219 = (((((((((((((((v_25 | v_24) | v_23) | v_22) | v_21) | v_27) | v_26) | ~v_446) | ~v_445) | ~v_332) | ~v_444) | ~v_294) | ~v_331) | ~v_443) | ~v_293) | v_447) ;
	assign x_1218 = (v_448 | ~v_14) ;
	assign x_1217 = (v_448 | v_42) ;
	assign x_1216 = (v_449 | v_14) ;
	assign x_1215 = (v_449 | v_45) ;
	assign x_1214 = (v_450 | ~v_14) ;
	assign x_1213 = (v_450 | v_3) ;
	assign x_1211 = (v_451 | v_14) ;
	assign x_1210 = (((((((((((((((v_39 | v_38) | v_35) | v_37) | v_36) | v_34) | v_40) | ~v_451) | ~v_450) | ~v_300) | ~v_449) | ~v_338) | ~v_337) | ~v_448) | ~v_299) | v_452) ;
	assign x_1209 = (v_453 | ~v_452) ;
	assign x_1208 = (v_453 | ~v_447) ;
	assign x_1207 = (v_453 | ~v_442) ;
	assign x_1206 = (v_454 | v_16) ;
	assign x_1205 = (v_454 | ~v_74) ;
	assign x_1204 = (v_455 | v_19) ;
	assign x_1203 = (v_455 | v_74) ;
	assign x_1202 = (v_456 | v_1) ;
	assign x_1201 = (v_456 | ~v_75) ;
	assign x_1200 = (v_457 | v_5) ;
	assign x_1199 = (v_457 | v_75) ;
	assign x_1198 = (((((((((((((((v_12 | v_11) | v_10) | v_69) | v_68) | v_48) | v_47) | ~v_173) | ~v_457) | ~v_456) | ~v_455) | ~v_454) | ~v_171) | ~v_248) | ~v_247) | v_458) ;
	assign x_1196 = (v_459 | ~v_74) ;
	assign x_1195 = (v_460 | v_32) ;
	assign x_1194 = (v_460 | v_74) ;
	assign x_1193 = (v_461 | v_2) ;
	assign x_1192 = (v_461 | ~v_75) ;
	assign x_1191 = (v_462 | v_4) ;
	assign x_1189 = (((((((((((((((v_25 | v_24) | v_26) | v_54) | v_53) | v_71) | v_70) | ~v_182) | ~v_462) | ~v_461) | ~v_181) | ~v_460) | ~v_459) | ~v_256) | ~v_255) | v_463) ;
	assign x_1188 = (v_464 | ~v_74) ;
	assign x_1187 = (v_464 | v_42) ;
	assign x_1186 = (v_465 | v_45) ;
	assign x_1185 = (v_465 | v_74) ;
	assign x_1184 = (v_466 | v_3) ;
	assign x_1182 = (v_467 | v_6) ;
	assign x_1181 = (v_467 | v_75) ;
	assign x_1180 = (((((((((((((((v_39 | v_38) | v_37) | v_56) | v_57) | v_73) | v_72) | ~v_191) | ~v_467) | ~v_466) | ~v_465) | ~v_464) | ~v_190) | ~v_262) | ~v_261) | v_468) ;
	assign x_1179 = (v_469 | ~v_468) ;
	assign x_1178 = (v_469 | ~v_463) ;
	assign x_1177 = (v_469 | ~v_458) ;
	assign x_1176 = (v_470 | ~v_1) ;
	assign x_1175 = (v_470 | v_2) ;
	assign x_1174 = (v_471 | ~v_2) ;
	assign x_1173 = (v_471 | v_3) ;
	assign x_1172 = (v_472 | ~v_6) ;
	assign x_1171 = (v_472 | v_4) ;
	assign x_1170 = (v_473 | ~v_4) ;
	assign x_1169 = (v_473 | v_5) ;
	assign x_1167 = ((~v_59 | ~v_78) | v_475) ;
	assign x_1166 = ((~v_50 | ~v_76) | v_476) ;
	assign x_1165 = (v_477 | ~v_63) ;
	assign x_1164 = (v_477 | ~v_476) ;
	assign x_1163 = (v_477 | ~v_475) ;
	assign x_1162 = ((~v_60 | ~v_477) | v_478) ;
	assign x_1161 = ((~v_74 | ~v_78) | v_479) ;
	assign x_1160 = ((~v_51 | ~v_63) | v_480) ;
	assign x_1159 = (v_481 | ~v_76) ;
	assign x_1158 = (v_481 | ~v_480) ;
	assign x_1157 = (v_481 | ~v_479) ;
	assign x_1156 = ((~v_75 | ~v_481) | v_482) ;
	assign x_1155 = ((~v_75 | ~v_76) | v_483) ;
	assign x_1154 = ((~v_60 | ~v_63) | v_484) ;
	assign x_1152 = (v_485 | ~v_484) ;
	assign x_1151 = (v_485 | ~v_483) ;
	assign x_1150 = (v_485 | ~v_482) ;
	assign x_1149 = (v_485 | ~v_478) ;
	assign x_1148 = ((~v_76 | ~v_79) | v_486) ;
	assign x_1147 = ((~v_51 | ~v_59) | v_487) ;
	assign x_1146 = (v_488 | ~v_74) ;
	assign x_1145 = (v_488 | ~v_487) ;
	assign x_1144 = (v_488 | ~v_486) ;
	assign x_1143 = ((~v_77 | ~v_488) | v_489) ;
	assign x_1142 = ((~v_63 | ~v_79) | v_490) ;
	assign x_1141 = ((~v_50 | ~v_74) | v_491) ;
	assign x_1140 = (v_492 | ~v_59) ;
	assign x_1139 = (v_492 | ~v_491) ;
	assign x_1137 = ((~v_64 | ~v_492) | v_493) ;
	assign x_1136 = ((~v_74 | ~v_77) | v_494) ;
	assign x_1135 = ((~v_59 | ~v_64) | v_495) ;
	assign x_1134 = (v_496 | ~v_79) ;
	assign x_1133 = (v_496 | ~v_495) ;
	assign x_1132 = (v_496 | ~v_494) ;
	assign x_1130 = (v_496 | ~v_489) ;
	assign x_1129 = ((~v_496 | ~v_485) | v_497) ;
	assign x_1128 = (v_498 | ~v_78) ;
	assign x_1127 = (v_498 | ~v_484) ;
	assign x_1126 = (v_498 | ~v_483) ;
	assign x_1125 = ((~v_74 | ~v_498) | v_499) ;
	assign x_1123 = (v_501 | ~v_76) ;
	assign x_1122 = (v_501 | ~v_480) ;
	assign x_1121 = (v_501 | ~v_479) ;
	assign x_1120 = (v_501 | ~v_500) ;
	assign x_1119 = (v_501 | ~v_499) ;
	assign x_1118 = ((~v_77 | ~v_78) | v_502) ;
	assign x_1117 = ((~v_50 | ~v_60) | v_503) ;
	assign x_1116 = (v_504 | ~v_75) ;
	assign x_1115 = (v_504 | ~v_503) ;
	assign x_1114 = (v_504 | ~v_502) ;
	assign x_1113 = ((~v_79 | ~v_504) | v_505) ;
	assign x_1112 = ((~v_63 | ~v_77) | v_506) ;
	assign x_1111 = ((~v_59 | ~v_75) | v_507) ;
	assign x_1110 = (v_508 | ~v_50) ;
	assign x_1108 = (v_508 | ~v_506) ;
	assign x_1107 = ((~v_64 | ~v_508) | v_509) ;
	assign x_1106 = ((~v_75 | ~v_79) | v_510) ;
	assign x_1105 = ((~v_50 | ~v_64) | v_511) ;
	assign x_1104 = (v_512 | ~v_77) ;
	assign x_1103 = (v_512 | ~v_511) ;
	assign x_1102 = (v_512 | ~v_510) ;
	assign x_1101 = (v_512 | ~v_509) ;
	assign x_1100 = (v_512 | ~v_505) ;
	assign x_1099 = ((~v_512 | ~v_501) | v_513) ;
	assign x_1098 = ((~v_59 | ~v_498) | v_514) ;
	assign x_1097 = ((~v_50 | ~v_481) | v_515) ;
	assign x_1096 = (v_516 | ~v_63) ;
	assign x_1095 = (v_516 | ~v_476) ;
	assign x_1093 = (v_516 | ~v_475) ;
	assign x_1092 = (v_516 | ~v_514) ;
	assign x_1091 = ((~v_64 | ~v_78) | v_517) ;
	assign x_1090 = ((~v_51 | ~v_75) | v_518) ;
	assign x_1089 = (v_519 | ~v_60) ;
	assign x_1088 = (v_519 | ~v_518) ;
	assign x_1087 = (v_519 | ~v_517) ;
	assign x_1086 = ((~v_79 | ~v_519) | v_520) ;
	assign x_1085 = ((~v_60 | ~v_74) | v_521) ;
	assign x_1084 = ((~v_64 | ~v_76) | v_522) ;
	assign x_1083 = (v_523 | ~v_51) ;
	assign x_1082 = (v_523 | ~v_522) ;
	assign x_1081 = (v_523 | ~v_521) ;
	assign x_1080 = ((~v_77 | ~v_523) | v_524) ;
	assign x_1078 = ((~v_51 | ~v_77) | v_526) ;
	assign x_1077 = (v_527 | ~v_64) ;
	assign x_1076 = (v_527 | ~v_526) ;
	assign x_1075 = (v_527 | ~v_525) ;
	assign x_1074 = (v_527 | ~v_524) ;
	assign x_1073 = (v_527 | ~v_520) ;
	assign x_1071 = (v_529 | ~v_65) ;
	assign x_1070 = (v_529 | ~v_528) ;
	assign x_1069 = (v_529 | ~v_513) ;
	assign x_1068 = (v_529 | ~v_497) ;
	assign x_1067 = (v_530 | ~v_79) ;
	assign x_1066 = (v_530 | ~v_495) ;
	assign x_1064 = ((~v_76 | ~v_530) | v_531) ;
	assign x_1063 = ((~v_51 | ~v_492) | v_532) ;
	assign x_1062 = (v_533 | ~v_74) ;
	assign x_1061 = (v_533 | ~v_487) ;
	assign x_1060 = (v_533 | ~v_486) ;
	assign x_1059 = (v_533 | ~v_532) ;
	assign x_1058 = (v_533 | ~v_531) ;
	assign x_1057 = (v_534 | ~v_77) ;
	assign x_1056 = (v_534 | ~v_511) ;
	assign x_1055 = (v_534 | ~v_510) ;
	assign x_1054 = ((~v_78 | ~v_534) | v_535) ;
	assign x_1053 = ((~v_60 | ~v_508) | v_536) ;
	assign x_1052 = (v_537 | ~v_75) ;
	assign x_1051 = (v_537 | ~v_503) ;
	assign x_1049 = (v_537 | ~v_536) ;
	assign x_1048 = (v_537 | ~v_535) ;
	assign x_1047 = ((~v_537 | ~v_533) | v_538) ;
	assign x_1046 = ((~v_63 | ~v_530) | v_539) ;
	assign x_1045 = ((~v_50 | ~v_488) | v_540) ;
	assign x_1044 = (v_541 | ~v_59) ;
	assign x_1043 = (v_541 | ~v_491) ;
	assign x_1042 = (v_541 | ~v_490) ;
	assign x_1041 = (v_541 | ~v_540) ;
	assign x_1040 = (v_541 | ~v_539) ;
	assign x_1039 = (v_542 | ~v_64) ;
	assign x_1038 = (v_542 | ~v_526) ;
	assign x_1037 = (v_542 | ~v_525) ;
	assign x_1036 = ((~v_78 | ~v_542) | v_543) ;
	assign x_1034 = (v_545 | ~v_60) ;
	assign x_1033 = (v_545 | ~v_518) ;
	assign x_1032 = (v_545 | ~v_517) ;
	assign x_1031 = (v_545 | ~v_544) ;
	assign x_1030 = (v_545 | ~v_543) ;
	assign x_1029 = ((~v_545 | ~v_541) | v_546) ;
	assign x_1028 = (v_547 | ~v_61) ;
	assign x_1027 = (v_547 | ~v_546) ;
	assign x_1026 = (v_547 | ~v_538) ;
	assign x_1025 = (v_547 | ~v_497) ;
	assign x_1024 = ((~v_63 | ~v_534) | v_548) ;
	assign x_1023 = ((~v_59 | ~v_504) | v_549) ;
	assign x_1022 = (v_550 | ~v_50) ;
	assign x_1021 = (v_550 | ~v_507) ;
	assign x_1019 = (v_550 | ~v_549) ;
	assign x_1018 = (v_550 | ~v_548) ;
	assign x_1017 = ((~v_76 | ~v_542) | v_551) ;
	assign x_1016 = ((~v_74 | ~v_519) | v_552) ;
	assign x_1015 = (v_553 | ~v_51) ;
	assign x_1014 = (v_553 | ~v_522) ;
	assign x_1012 = (v_553 | ~v_552) ;
	assign x_1011 = (v_553 | ~v_551) ;
	assign x_1010 = ((~v_553 | ~v_550) | v_554) ;
	assign x_1009 = (v_555 | ~v_52) ;
	assign x_1008 = (v_555 | ~v_554) ;
	assign x_1007 = (v_555 | ~v_538) ;
	assign x_1005 = (v_556 | ~v_14) ;
	assign x_1004 = (v_556 | ~v_554) ;
	assign x_1003 = (v_556 | ~v_546) ;
	assign x_1002 = (v_556 | ~v_528) ;
	assign x_1001 = ((~v_1 | v_78) | v_557) ;
	assign x_1000 = ((~v_16 | v_79) | v_558) ;
	assign x_999 = ((~v_5 | ~v_78) | v_559) ;
	assign x_998 = ((~v_17 | v_65) | v_560) ;
	assign x_997 = ((~v_20 | ~v_65) | v_561) ;
	assign x_996 = ((~v_18 | ~v_61) | v_562) ;
	assign x_995 = ((~v_19 | ~v_79) | v_563) ;
	assign x_994 = ((~v_15 | v_61) | v_564) ;
	assign x_993 = (v_565 | ~v_10) ;
	assign x_992 = (v_565 | ~v_13) ;
	assign x_990 = (v_565 | ~v_48) ;
	assign x_989 = (v_565 | ~v_49) ;
	assign x_988 = (v_565 | ~v_62) ;
	assign x_987 = (v_565 | ~v_68) ;
	assign x_986 = (v_565 | ~v_564) ;
	assign x_985 = (v_565 | ~v_563) ;
	assign x_984 = (v_565 | ~v_562) ;
	assign x_983 = (v_565 | ~v_561) ;
	assign x_982 = (v_565 | ~v_560) ;
	assign x_981 = (v_565 | ~v_559) ;
	assign x_980 = (v_565 | ~v_558) ;
	assign x_979 = (v_565 | ~v_557) ;
	assign x_978 = ((~v_2 | v_78) | v_566) ;
	assign x_977 = ((~v_29 | v_79) | v_567) ;
	assign x_975 = ((~v_32 | ~v_79) | v_569) ;
	assign x_974 = ((~v_30 | v_65) | v_570) ;
	assign x_973 = ((~v_33 | ~v_65) | v_571) ;
	assign x_972 = ((~v_31 | ~v_61) | v_572) ;
	assign x_971 = ((~v_28 | v_61) | v_573) ;
	assign x_970 = (v_574 | ~v_24) ;
	assign x_969 = (v_574 | ~v_27) ;
	assign x_968 = (v_574 | ~v_53) ;
	assign x_967 = (v_574 | ~v_54) ;
	assign x_966 = (v_574 | ~v_55) ;
	assign x_965 = (v_574 | ~v_66) ;
	assign x_964 = (v_574 | ~v_70) ;
	assign x_963 = (v_574 | ~v_573) ;
	assign x_962 = (v_574 | ~v_572) ;
	assign x_960 = (v_574 | ~v_570) ;
	assign x_959 = (v_574 | ~v_569) ;
	assign x_958 = (v_574 | ~v_568) ;
	assign x_957 = (v_574 | ~v_567) ;
	assign x_956 = (v_574 | ~v_566) ;
	assign x_955 = ((~v_3 | v_78) | v_575) ;
	assign x_953 = ((~v_6 | ~v_78) | v_577) ;
	assign x_952 = ((~v_45 | ~v_79) | v_578) ;
	assign x_951 = ((~v_43 | v_65) | v_579) ;
	assign x_950 = ((~v_46 | ~v_65) | v_580) ;
	assign x_949 = ((~v_44 | ~v_61) | v_581) ;
	assign x_948 = ((~v_41 | v_61) | v_582) ;
	assign x_946 = (v_583 | ~v_40) ;
	assign x_945 = (v_583 | ~v_56) ;
	assign x_944 = (v_583 | ~v_57) ;
	assign x_943 = (v_583 | ~v_58) ;
	assign x_942 = (v_583 | ~v_67) ;
	assign x_941 = (v_583 | ~v_72) ;
	assign x_940 = (v_583 | ~v_582) ;
	assign x_939 = (v_583 | ~v_581) ;
	assign x_938 = (v_583 | ~v_580) ;
	assign x_937 = (v_583 | ~v_579) ;
	assign x_936 = (v_583 | ~v_578) ;
	assign x_935 = (v_583 | ~v_577) ;
	assign x_934 = (v_583 | ~v_576) ;
	assign x_933 = (v_583 | ~v_575) ;
	assign x_931 = ((~v_1 | v_79) | v_585) ;
	assign x_930 = ((~v_16 | v_78) | v_586) ;
	assign x_929 = ((~v_5 | ~v_79) | v_587) ;
	assign x_928 = ((~v_15 | v_65) | v_588) ;
	assign x_927 = ((~v_18 | ~v_65) | v_589) ;
	assign x_926 = ((~v_17 | v_61) | v_590) ;
	assign x_925 = ((~v_20 | ~v_61) | v_591) ;
	assign x_924 = ((~v_19 | ~v_78) | v_592) ;
	assign x_923 = (v_593 | ~v_11) ;
	assign x_922 = (v_593 | ~v_12) ;
	assign x_921 = (v_593 | ~v_47) ;
	assign x_920 = (v_593 | ~v_48) ;
	assign x_919 = (v_593 | ~v_68) ;
	assign x_918 = (v_593 | ~v_69) ;
	assign x_916 = (v_593 | ~v_592) ;
	assign x_915 = (v_593 | ~v_591) ;
	assign x_914 = (v_593 | ~v_590) ;
	assign x_913 = (v_593 | ~v_589) ;
	assign x_912 = (v_593 | ~v_588) ;
	assign x_911 = (v_593 | ~v_587) ;
	assign x_910 = (v_593 | ~v_586) ;
	assign x_909 = (v_593 | ~v_585) ;
	assign x_908 = ((~v_2 | v_79) | v_594) ;
	assign x_907 = ((~v_29 | v_78) | v_595) ;
	assign x_906 = ((~v_4 | ~v_79) | v_596) ;
	assign x_905 = ((~v_32 | ~v_78) | v_597) ;
	assign x_904 = ((~v_28 | v_65) | v_598) ;
	assign x_903 = ((~v_31 | ~v_65) | v_599) ;
	assign x_901 = ((~v_33 | ~v_61) | v_601) ;
	assign x_900 = (v_602 | ~v_25) ;
	assign x_899 = (v_602 | ~v_26) ;
	assign x_898 = (v_602 | ~v_53) ;
	assign x_897 = (v_602 | ~v_54) ;
	assign x_896 = (v_602 | ~v_70) ;
	assign x_895 = (v_602 | ~v_71) ;
	assign x_894 = (v_602 | ~v_81) ;
	assign x_893 = (v_602 | ~v_601) ;
	assign x_892 = (v_602 | ~v_600) ;
	assign x_891 = (v_602 | ~v_599) ;
	assign x_890 = (v_602 | ~v_598) ;
	assign x_889 = (v_602 | ~v_597) ;
	assign x_888 = (v_602 | ~v_596) ;
	assign x_886 = (v_602 | ~v_594) ;
	assign x_885 = ((~v_3 | v_79) | v_603) ;
	assign x_884 = ((~v_42 | v_78) | v_604) ;
	assign x_883 = ((~v_6 | ~v_79) | v_605) ;
	assign x_882 = ((~v_45 | ~v_78) | v_606) ;
	assign x_881 = ((~v_41 | v_65) | v_607) ;
	assign x_880 = ((~v_44 | ~v_65) | v_608) ;
	assign x_879 = ((~v_43 | v_61) | v_609) ;
	assign x_878 = ((~v_46 | ~v_61) | v_610) ;
	assign x_877 = (v_611 | ~v_38) ;
	assign x_876 = (v_611 | ~v_39) ;
	assign x_875 = (v_611 | ~v_56) ;
	assign x_874 = (v_611 | ~v_57) ;
	assign x_873 = (v_611 | ~v_72) ;
	assign x_871 = (v_611 | ~v_82) ;
	assign x_870 = (v_611 | ~v_610) ;
	assign x_869 = (v_611 | ~v_609) ;
	assign x_868 = (v_611 | ~v_608) ;
	assign x_867 = (v_611 | ~v_607) ;
	assign x_866 = (v_611 | ~v_606) ;
	assign x_865 = (v_611 | ~v_605) ;
	assign x_864 = (v_611 | ~v_604) ;
	assign x_863 = (v_611 | ~v_603) ;
	assign x_862 = (((~v_611 | ~v_602) | ~v_593) | v_612) ;
	assign x_861 = ((~v_1 | v_76) | v_613) ;
	assign x_860 = ((~v_16 | v_77) | v_614) ;
	assign x_859 = ((~v_5 | ~v_76) | v_615) ;
	assign x_858 = ((~v_18 | ~v_52) | v_616) ;
	assign x_856 = ((~v_15 | v_52) | v_618) ;
	assign x_855 = (v_619 | ~v_10) ;
	assign x_854 = (v_619 | ~v_12) ;
	assign x_853 = (v_619 | ~v_13) ;
	assign x_852 = (v_619 | ~v_47) ;
	assign x_851 = (v_619 | ~v_48) ;
	assign x_850 = (v_619 | ~v_62) ;
	assign x_849 = (v_619 | ~v_68) ;
	assign x_848 = (v_619 | ~v_618) ;
	assign x_847 = (v_619 | ~v_617) ;
	assign x_846 = (v_619 | ~v_616) ;
	assign x_845 = (v_619 | ~v_561) ;
	assign x_844 = (v_619 | ~v_560) ;
	assign x_843 = (v_619 | ~v_615) ;
	assign x_841 = (v_619 | ~v_613) ;
	assign x_840 = ((~v_2 | v_76) | v_620) ;
	assign x_839 = ((~v_29 | v_77) | v_621) ;
	assign x_838 = ((~v_4 | ~v_76) | v_622) ;
	assign x_837 = ((~v_32 | ~v_77) | v_623) ;
	assign x_836 = ((~v_28 | v_52) | v_624) ;
	assign x_834 = (v_626 | ~v_24) ;
	assign x_833 = (v_626 | ~v_26) ;
	assign x_832 = (v_626 | ~v_27) ;
	assign x_831 = (v_626 | ~v_53) ;
	assign x_830 = (v_626 | ~v_54) ;
	assign x_829 = (v_626 | ~v_66) ;
	assign x_827 = (v_626 | ~v_625) ;
	assign x_826 = (v_626 | ~v_624) ;
	assign x_825 = (v_626 | ~v_571) ;
	assign x_824 = (v_626 | ~v_570) ;
	assign x_823 = (v_626 | ~v_623) ;
	assign x_822 = (v_626 | ~v_622) ;
	assign x_821 = (v_626 | ~v_621) ;
	assign x_820 = (v_626 | ~v_620) ;
	assign x_819 = ((~v_3 | v_76) | v_627) ;
	assign x_818 = ((~v_42 | v_77) | v_628) ;
	assign x_817 = ((~v_6 | ~v_76) | v_629) ;
	assign x_816 = ((~v_45 | ~v_77) | v_630) ;
	assign x_815 = ((~v_41 | v_52) | v_631) ;
	assign x_814 = ((~v_44 | ~v_52) | v_632) ;
	assign x_812 = (v_633 | ~v_39) ;
	assign x_811 = (v_633 | ~v_40) ;
	assign x_810 = (v_633 | ~v_56) ;
	assign x_809 = (v_633 | ~v_57) ;
	assign x_808 = (v_633 | ~v_67) ;
	assign x_807 = (v_633 | ~v_72) ;
	assign x_806 = (v_633 | ~v_632) ;
	assign x_805 = (v_633 | ~v_631) ;
	assign x_804 = (v_633 | ~v_580) ;
	assign x_803 = (v_633 | ~v_579) ;
	assign x_802 = (v_633 | ~v_630) ;
	assign x_801 = (v_633 | ~v_629) ;
	assign x_800 = (v_633 | ~v_628) ;
	assign x_799 = (v_633 | ~v_627) ;
	assign x_797 = ((~v_1 | v_77) | v_635) ;
	assign x_796 = ((~v_16 | v_76) | v_636) ;
	assign x_795 = ((~v_5 | ~v_77) | v_637) ;
	assign x_794 = ((~v_17 | v_52) | v_638) ;
	assign x_793 = ((~v_20 | ~v_52) | v_639) ;
	assign x_792 = ((~v_19 | ~v_76) | v_640) ;
	assign x_791 = (v_641 | ~v_11) ;
	assign x_790 = (v_641 | ~v_12) ;
	assign x_789 = (v_641 | ~v_13) ;
	assign x_788 = (v_641 | ~v_47) ;
	assign x_787 = (v_641 | ~v_48) ;
	assign x_786 = (v_641 | ~v_68) ;
	assign x_785 = (v_641 | ~v_80) ;
	assign x_784 = (v_641 | ~v_640) ;
	assign x_782 = (v_641 | ~v_638) ;
	assign x_781 = (v_641 | ~v_589) ;
	assign x_780 = (v_641 | ~v_588) ;
	assign x_779 = (v_641 | ~v_637) ;
	assign x_778 = (v_641 | ~v_636) ;
	assign x_777 = (v_641 | ~v_635) ;
	assign x_775 = ((~v_29 | v_76) | v_643) ;
	assign x_774 = ((~v_4 | ~v_77) | v_644) ;
	assign x_773 = ((~v_32 | ~v_76) | v_645) ;
	assign x_772 = ((~v_30 | v_52) | v_646) ;
	assign x_771 = ((~v_33 | ~v_52) | v_647) ;
	assign x_770 = (v_648 | ~v_25) ;
	assign x_768 = (v_648 | ~v_27) ;
	assign x_767 = (v_648 | ~v_53) ;
	assign x_766 = (v_648 | ~v_54) ;
	assign x_765 = (v_648 | ~v_70) ;
	assign x_764 = (v_648 | ~v_81) ;
	assign x_763 = (v_648 | ~v_647) ;
	assign x_762 = (v_648 | ~v_646) ;
	assign x_761 = (v_648 | ~v_599) ;
	assign x_760 = (v_648 | ~v_598) ;
	assign x_759 = (v_648 | ~v_645) ;
	assign x_758 = (v_648 | ~v_644) ;
	assign x_757 = (v_648 | ~v_643) ;
	assign x_756 = (v_648 | ~v_642) ;
	assign x_755 = ((~v_3 | v_77) | v_649) ;
	assign x_753 = ((~v_6 | ~v_77) | v_651) ;
	assign x_752 = ((~v_43 | v_52) | v_652) ;
	assign x_751 = ((~v_46 | ~v_52) | v_653) ;
	assign x_750 = ((~v_45 | ~v_76) | v_654) ;
	assign x_749 = (v_655 | ~v_38) ;
	assign x_748 = (v_655 | ~v_39) ;
	assign x_747 = (v_655 | ~v_40) ;
	assign x_746 = (v_655 | ~v_56) ;
	assign x_745 = (v_655 | ~v_57) ;
	assign x_744 = (v_655 | ~v_72) ;
	assign x_743 = (v_655 | ~v_82) ;
	assign x_742 = (v_655 | ~v_654) ;
	assign x_741 = (v_655 | ~v_653) ;
	assign x_740 = (v_655 | ~v_652) ;
	assign x_738 = (v_655 | ~v_607) ;
	assign x_737 = (v_655 | ~v_651) ;
	assign x_736 = (v_655 | ~v_650) ;
	assign x_735 = (v_655 | ~v_649) ;
	assign x_734 = (((~v_655 | ~v_648) | ~v_641) | v_656) ;
	assign x_733 = ((~v_1 | v_74) | v_657) ;
	assign x_732 = ((~v_5 | ~v_74) | v_658) ;
	assign x_731 = ((~v_19 | ~v_75) | v_659) ;
	assign x_730 = ((~v_16 | v_75) | v_660) ;
	assign x_729 = (v_661 | ~v_10) ;
	assign x_728 = (v_661 | ~v_11) ;
	assign x_727 = (v_661 | ~v_13) ;
	assign x_726 = (v_661 | ~v_47) ;
	assign x_725 = (v_661 | ~v_48) ;
	assign x_723 = (v_661 | ~v_68) ;
	assign x_722 = (v_661 | ~v_660) ;
	assign x_721 = (v_661 | ~v_659) ;
	assign x_720 = (v_661 | ~v_618) ;
	assign x_719 = (v_661 | ~v_616) ;
	assign x_718 = (v_661 | ~v_591) ;
	assign x_716 = (v_661 | ~v_658) ;
	assign x_715 = (v_661 | ~v_657) ;
	assign x_714 = ((~v_2 | v_74) | v_662) ;
	assign x_713 = ((~v_4 | ~v_74) | v_663) ;
	assign x_712 = ((~v_32 | ~v_75) | v_664) ;
	assign x_711 = ((~v_29 | v_75) | v_665) ;
	assign x_709 = (v_666 | ~v_25) ;
	assign x_708 = (v_666 | ~v_27) ;
	assign x_707 = (v_666 | ~v_53) ;
	assign x_706 = (v_666 | ~v_54) ;
	assign x_705 = (v_666 | ~v_55) ;
	assign x_704 = (v_666 | ~v_70) ;
	assign x_703 = (v_666 | ~v_665) ;
	assign x_702 = (v_666 | ~v_664) ;
	assign x_701 = (v_666 | ~v_625) ;
	assign x_700 = (v_666 | ~v_624) ;
	assign x_699 = (v_666 | ~v_601) ;
	assign x_698 = (v_666 | ~v_600) ;
	assign x_697 = (v_666 | ~v_663) ;
	assign x_696 = (v_666 | ~v_662) ;
	assign x_694 = ((~v_42 | v_75) | v_668) ;
	assign x_693 = ((~v_6 | ~v_74) | v_669) ;
	assign x_692 = ((~v_45 | ~v_75) | v_670) ;
	assign x_691 = (v_671 | ~v_37) ;
	assign x_690 = (v_671 | ~v_38) ;
	assign x_689 = (v_671 | ~v_40) ;
	assign x_688 = (v_671 | ~v_56) ;
	assign x_687 = (v_671 | ~v_57) ;
	assign x_686 = (v_671 | ~v_58) ;
	assign x_685 = (v_671 | ~v_72) ;
	assign x_684 = (v_671 | ~v_670) ;
	assign x_683 = (v_671 | ~v_632) ;
	assign x_682 = (v_671 | ~v_631) ;
	assign x_681 = (v_671 | ~v_610) ;
	assign x_679 = (v_671 | ~v_669) ;
	assign x_678 = (v_671 | ~v_668) ;
	assign x_677 = (v_671 | ~v_667) ;
	assign x_676 = (((~v_671 | ~v_666) | ~v_661) | v_672) ;
	assign x_675 = ((~v_1 | v_63) | v_673) ;
	assign x_674 = ((~v_16 | v_64) | v_674) ;
	assign x_673 = ((~v_5 | ~v_63) | v_675) ;
	assign x_672 = ((~v_19 | ~v_64) | v_676) ;
	assign x_671 = ((~v_14 | ~v_18) | v_677) ;
	assign x_670 = ((~v_15 | v_14) | v_678) ;
	assign x_669 = (v_679 | ~v_8) ;
	assign x_668 = (v_679 | ~v_10) ;
	assign x_667 = (v_679 | ~v_12) ;
	assign x_666 = (v_679 | ~v_13) ;
	assign x_664 = (v_679 | ~v_48) ;
	assign x_663 = (v_679 | ~v_62) ;
	assign x_662 = (v_679 | ~v_678) ;
	assign x_661 = (v_679 | ~v_677) ;
	assign x_660 = (v_679 | ~v_561) ;
	assign x_659 = (v_679 | ~v_560) ;
	assign x_657 = (v_679 | ~v_675) ;
	assign x_656 = (v_679 | ~v_674) ;
	assign x_655 = (v_679 | ~v_673) ;
	assign x_654 = ((~v_2 | v_63) | v_680) ;
	assign x_653 = ((~v_29 | v_64) | v_681) ;
	assign x_652 = ((~v_4 | ~v_63) | v_682) ;
	assign x_650 = ((~v_28 | v_14) | v_684) ;
	assign x_649 = ((~v_14 | ~v_31) | v_685) ;
	assign x_648 = (v_686 | ~v_22) ;
	assign x_647 = (v_686 | ~v_24) ;
	assign x_646 = (v_686 | ~v_26) ;
	assign x_645 = (v_686 | ~v_27) ;
	assign x_644 = (v_686 | ~v_53) ;
	assign x_643 = (v_686 | ~v_54) ;
	assign x_642 = (v_686 | ~v_66) ;
	assign x_641 = (v_686 | ~v_685) ;
	assign x_640 = (v_686 | ~v_684) ;
	assign x_639 = (v_686 | ~v_571) ;
	assign x_638 = (v_686 | ~v_570) ;
	assign x_637 = (v_686 | ~v_683) ;
	assign x_635 = (v_686 | ~v_681) ;
	assign x_634 = (v_686 | ~v_680) ;
	assign x_633 = ((~v_3 | v_63) | v_687) ;
	assign x_632 = ((~v_42 | v_64) | v_688) ;
	assign x_631 = ((~v_45 | ~v_64) | v_689) ;
	assign x_630 = ((v_14 | ~v_41) | v_690) ;
	assign x_629 = ((~v_14 | ~v_44) | v_691) ;
	assign x_628 = ((~v_6 | ~v_63) | v_692) ;
	assign x_627 = (v_693 | ~v_35) ;
	assign x_626 = (v_693 | ~v_37) ;
	assign x_625 = (v_693 | ~v_39) ;
	assign x_624 = (v_693 | ~v_40) ;
	assign x_623 = (v_693 | ~v_56) ;
	assign x_622 = (v_693 | ~v_57) ;
	assign x_620 = (v_693 | ~v_692) ;
	assign x_619 = (v_693 | ~v_691) ;
	assign x_618 = (v_693 | ~v_690) ;
	assign x_617 = (v_693 | ~v_580) ;
	assign x_616 = (v_693 | ~v_579) ;
	assign x_615 = (v_693 | ~v_689) ;
	assign x_614 = (v_693 | ~v_688) ;
	assign x_613 = (v_693 | ~v_687) ;
	assign x_612 = (((~v_693 | ~v_686) | ~v_679) | v_694) ;
	assign x_611 = ((~v_1 | v_65) | v_695) ;
	assign x_610 = ((~v_16 | v_65) | v_696) ;
	assign x_609 = ((~v_5 | ~v_65) | v_697) ;
	assign x_608 = ((~v_19 | ~v_65) | v_698) ;
	assign x_607 = (v_699 | ~v_7) ;
	assign x_605 = (v_699 | ~v_13) ;
	assign x_604 = (v_699 | ~v_48) ;
	assign x_603 = (v_699 | ~v_62) ;
	assign x_602 = (v_699 | ~v_68) ;
	assign x_601 = (v_699 | ~v_80) ;
	assign x_600 = (v_699 | ~v_589) ;
	assign x_598 = (v_699 | ~v_698) ;
	assign x_597 = (v_699 | ~v_697) ;
	assign x_596 = (v_699 | ~v_696) ;
	assign x_595 = (v_699 | ~v_695) ;
	assign x_594 = (v_699 | ~v_561) ;
	assign x_593 = (v_699 | ~v_560) ;
	assign x_591 = ((~v_29 | v_65) | v_701) ;
	assign x_590 = ((~v_4 | ~v_65) | v_702) ;
	assign x_589 = ((~v_32 | ~v_65) | v_703) ;
	assign x_588 = (v_704 | ~v_21) ;
	assign x_587 = (v_704 | ~v_26) ;
	assign x_586 = (v_704 | ~v_27) ;
	assign x_585 = (v_704 | ~v_54) ;
	assign x_584 = (v_704 | ~v_66) ;
	assign x_583 = (v_704 | ~v_70) ;
	assign x_582 = (v_704 | ~v_81) ;
	assign x_581 = (v_704 | ~v_599) ;
	assign x_580 = (v_704 | ~v_598) ;
	assign x_579 = (v_704 | ~v_703) ;
	assign x_578 = (v_704 | ~v_702) ;
	assign x_576 = (v_704 | ~v_700) ;
	assign x_575 = (v_704 | ~v_571) ;
	assign x_574 = (v_704 | ~v_570) ;
	assign x_573 = ((~v_3 | v_65) | v_705) ;
	assign x_572 = ((~v_42 | v_65) | v_706) ;
	assign x_571 = ((~v_45 | ~v_65) | v_707) ;
	assign x_570 = ((~v_6 | ~v_65) | v_708) ;
	assign x_569 = (v_709 | ~v_34) ;
	assign x_568 = (v_709 | ~v_39) ;
	assign x_567 = (v_709 | ~v_40) ;
	assign x_566 = (v_709 | ~v_57) ;
	assign x_565 = (v_709 | ~v_67) ;
	assign x_564 = (v_709 | ~v_72) ;
	assign x_563 = (v_709 | ~v_82) ;
	assign x_561 = (v_709 | ~v_608) ;
	assign x_560 = (v_709 | ~v_607) ;
	assign x_559 = (v_709 | ~v_707) ;
	assign x_558 = (v_709 | ~v_706) ;
	assign x_557 = (v_709 | ~v_705) ;
	assign x_556 = (v_709 | ~v_580) ;
	assign x_555 = (v_709 | ~v_579) ;
	assign x_554 = (((~v_709 | ~v_704) | ~v_699) | v_710) ;
	assign x_553 = ((~v_1 | v_64) | v_711) ;
	assign x_552 = ((~v_16 | v_63) | v_712) ;
	assign x_551 = ((~v_5 | ~v_64) | v_713) ;
	assign x_550 = ((~v_19 | ~v_63) | v_714) ;
	assign x_549 = ((~v_17 | v_14) | v_715) ;
	assign x_548 = ((~v_14 | ~v_20) | v_716) ;
	assign x_546 = (v_717 | ~v_11) ;
	assign x_545 = (v_717 | ~v_12) ;
	assign x_544 = (v_717 | ~v_13) ;
	assign x_543 = (v_717 | ~v_47) ;
	assign x_542 = (v_717 | ~v_68) ;
	assign x_541 = (v_717 | ~v_80) ;
	assign x_539 = (v_717 | ~v_715) ;
	assign x_538 = (v_717 | ~v_714) ;
	assign x_537 = (v_717 | ~v_713) ;
	assign x_536 = (v_717 | ~v_589) ;
	assign x_535 = (v_717 | ~v_712) ;
	assign x_534 = (v_717 | ~v_711) ;
	assign x_532 = ((~v_2 | v_64) | v_718) ;
	assign x_531 = ((~v_29 | v_63) | v_719) ;
	assign x_530 = ((~v_4 | ~v_64) | v_720) ;
	assign x_529 = ((~v_32 | ~v_63) | v_721) ;
	assign x_528 = ((~v_30 | v_14) | v_722) ;
	assign x_527 = ((~v_14 | ~v_33) | v_723) ;
	assign x_526 = (v_724 | ~v_23) ;
	assign x_525 = (v_724 | ~v_25) ;
	assign x_524 = (v_724 | ~v_26) ;
	assign x_523 = (v_724 | ~v_27) ;
	assign x_522 = (v_724 | ~v_53) ;
	assign x_521 = (v_724 | ~v_70) ;
	assign x_520 = (v_724 | ~v_81) ;
	assign x_519 = (v_724 | ~v_723) ;
	assign x_517 = (v_724 | ~v_721) ;
	assign x_516 = (v_724 | ~v_720) ;
	assign x_515 = (v_724 | ~v_599) ;
	assign x_514 = (v_724 | ~v_719) ;
	assign x_513 = (v_724 | ~v_718) ;
	assign x_512 = (v_724 | ~v_598) ;
	assign x_511 = ((~v_3 | v_64) | v_725) ;
	assign x_510 = ((~v_42 | v_63) | v_726) ;
	assign x_509 = ((~v_45 | ~v_63) | v_727) ;
	assign x_508 = ((v_14 | ~v_43) | v_728) ;
	assign x_507 = ((~v_14 | ~v_46) | v_729) ;
	assign x_506 = ((~v_6 | ~v_64) | v_730) ;
	assign x_505 = (v_731 | ~v_36) ;
	assign x_504 = (v_731 | ~v_38) ;
	assign x_502 = (v_731 | ~v_40) ;
	assign x_501 = (v_731 | ~v_56) ;
	assign x_500 = (v_731 | ~v_72) ;
	assign x_499 = (v_731 | ~v_82) ;
	assign x_498 = (v_731 | ~v_730) ;
	assign x_497 = (v_731 | ~v_729) ;
	assign x_496 = (v_731 | ~v_728) ;
	assign x_495 = (v_731 | ~v_727) ;
	assign x_494 = (v_731 | ~v_608) ;
	assign x_493 = (v_731 | ~v_726) ;
	assign x_492 = (v_731 | ~v_725) ;
	assign x_491 = (v_731 | ~v_607) ;
	assign x_490 = (((~v_731 | ~v_724) | ~v_717) | v_732) ;
	assign x_489 = ((~v_16 | v_60) | v_733) ;
	assign x_487 = ((~v_5 | ~v_59) | v_735) ;
	assign x_486 = ((~v_19 | ~v_60) | v_736) ;
	assign x_485 = (v_737 | ~v_8) ;
	assign x_484 = (v_737 | ~v_10) ;
	assign x_483 = (v_737 | ~v_11) ;
	assign x_482 = (v_737 | ~v_12) ;
	assign x_480 = (v_737 | ~v_47) ;
	assign x_479 = (v_737 | ~v_48) ;
	assign x_478 = (v_737 | ~v_736) ;
	assign x_477 = (v_737 | ~v_735) ;
	assign x_476 = (v_737 | ~v_678) ;
	assign x_475 = (v_737 | ~v_734) ;
	assign x_473 = (v_737 | ~v_677) ;
	assign x_472 = (v_737 | ~v_591) ;
	assign x_471 = (v_737 | ~v_590) ;
	assign x_470 = ((~v_29 | v_60) | v_738) ;
	assign x_469 = ((~v_4 | ~v_59) | v_739) ;
	assign x_468 = ((~v_2 | v_59) | v_740) ;
	assign x_467 = ((~v_32 | ~v_60) | v_741) ;
	assign x_466 = (v_742 | ~v_22) ;
	assign x_465 = (v_742 | ~v_24) ;
	assign x_464 = (v_742 | ~v_25) ;
	assign x_463 = (v_742 | ~v_26) ;
	assign x_462 = (v_742 | ~v_27) ;
	assign x_461 = (v_742 | ~v_53) ;
	assign x_460 = (v_742 | ~v_54) ;
	assign x_458 = (v_742 | ~v_740) ;
	assign x_457 = (v_742 | ~v_739) ;
	assign x_456 = (v_742 | ~v_685) ;
	assign x_455 = (v_742 | ~v_684) ;
	assign x_454 = (v_742 | ~v_601) ;
	assign x_453 = (v_742 | ~v_600) ;
	assign x_452 = (v_742 | ~v_738) ;
	assign x_451 = ((~v_42 | v_60) | v_743) ;
	assign x_450 = ((~v_6 | ~v_59) | v_744) ;
	assign x_449 = ((~v_3 | v_59) | v_745) ;
	assign x_448 = ((~v_45 | ~v_60) | v_746) ;
	assign x_447 = (v_747 | ~v_35) ;
	assign x_446 = (v_747 | ~v_37) ;
	assign x_445 = (v_747 | ~v_38) ;
	assign x_443 = (v_747 | ~v_40) ;
	assign x_442 = (v_747 | ~v_56) ;
	assign x_441 = (v_747 | ~v_57) ;
	assign x_440 = (v_747 | ~v_746) ;
	assign x_439 = (v_747 | ~v_745) ;
	assign x_438 = (v_747 | ~v_744) ;
	assign x_437 = (v_747 | ~v_691) ;
	assign x_436 = (v_747 | ~v_690) ;
	assign x_435 = (v_747 | ~v_610) ;
	assign x_434 = (v_747 | ~v_609) ;
	assign x_433 = (v_747 | ~v_743) ;
	assign x_432 = (((~v_747 | ~v_742) | ~v_737) | v_748) ;
	assign x_431 = ((~v_16 | v_61) | v_749) ;
	assign x_430 = ((~v_19 | ~v_61) | v_750) ;
	assign x_428 = ((~v_1 | v_61) | v_752) ;
	assign x_427 = (v_753 | ~v_7) ;
	assign x_426 = (v_753 | ~v_10) ;
	assign x_425 = (v_753 | ~v_11) ;
	assign x_424 = (v_753 | ~v_12) ;
	assign x_423 = (v_753 | ~v_13) ;
	assign x_422 = (v_753 | ~v_48) ;
	assign x_421 = (v_753 | ~v_68) ;
	assign x_420 = (v_753 | ~v_564) ;
	assign x_419 = (v_753 | ~v_752) ;
	assign x_418 = (v_753 | ~v_751) ;
	assign x_417 = (v_753 | ~v_562) ;
	assign x_416 = (v_753 | ~v_750) ;
	assign x_415 = (v_753 | ~v_749) ;
	assign x_413 = (v_753 | ~v_590) ;
	assign x_412 = ((~v_29 | v_61) | v_754) ;
	assign x_411 = ((~v_32 | ~v_61) | v_755) ;
	assign x_410 = ((~v_4 | ~v_61) | v_756) ;
	assign x_409 = ((~v_2 | v_61) | v_757) ;
	assign x_408 = (v_758 | ~v_21) ;
	assign x_407 = (v_758 | ~v_24) ;
	assign x_406 = (v_758 | ~v_25) ;
	assign x_405 = (v_758 | ~v_26) ;
	assign x_404 = (v_758 | ~v_27) ;
	assign x_403 = (v_758 | ~v_54) ;
	assign x_402 = (v_758 | ~v_70) ;
	assign x_401 = (v_758 | ~v_573) ;
	assign x_400 = (v_758 | ~v_757) ;
	assign x_398 = (v_758 | ~v_572) ;
	assign x_397 = (v_758 | ~v_755) ;
	assign x_396 = (v_758 | ~v_754) ;
	assign x_395 = (v_758 | ~v_601) ;
	assign x_394 = (v_758 | ~v_600) ;
	assign x_393 = ((~v_42 | v_61) | v_759) ;
	assign x_392 = ((~v_45 | ~v_61) | v_760) ;
	assign x_391 = ((~v_6 | ~v_61) | v_761) ;
	assign x_390 = ((~v_3 | v_61) | v_762) ;
	assign x_389 = (v_763 | ~v_34) ;
	assign x_388 = (v_763 | ~v_37) ;
	assign x_387 = (v_763 | ~v_38) ;
	assign x_386 = (v_763 | ~v_39) ;
	assign x_385 = (v_763 | ~v_40) ;
	assign x_383 = (v_763 | ~v_72) ;
	assign x_382 = (v_763 | ~v_582) ;
	assign x_381 = (v_763 | ~v_762) ;
	assign x_380 = (v_763 | ~v_761) ;
	assign x_379 = (v_763 | ~v_581) ;
	assign x_378 = (v_763 | ~v_760) ;
	assign x_377 = (v_763 | ~v_759) ;
	assign x_376 = (v_763 | ~v_610) ;
	assign x_375 = (v_763 | ~v_609) ;
	assign x_374 = (((~v_763 | ~v_758) | ~v_753) | v_764) ;
	assign x_373 = ((~v_19 | ~v_59) | v_765) ;
	assign x_372 = ((~v_16 | v_59) | v_766) ;
	assign x_371 = ((~v_1 | v_60) | v_767) ;
	assign x_370 = ((~v_5 | ~v_60) | v_768) ;
	assign x_368 = (v_769 | ~v_10) ;
	assign x_367 = (v_769 | ~v_11) ;
	assign x_366 = (v_769 | ~v_12) ;
	assign x_365 = (v_769 | ~v_13) ;
	assign x_364 = (v_769 | ~v_47) ;
	assign x_363 = (v_769 | ~v_68) ;
	assign x_361 = (v_769 | ~v_767) ;
	assign x_360 = (v_769 | ~v_766) ;
	assign x_359 = (v_769 | ~v_564) ;
	assign x_358 = (v_769 | ~v_716) ;
	assign x_357 = (v_769 | ~v_562) ;
	assign x_356 = (v_769 | ~v_715) ;
	assign x_354 = ((~v_29 | v_59) | v_770) ;
	assign x_353 = ((~v_32 | ~v_59) | v_771) ;
	assign x_352 = ((~v_2 | v_60) | v_772) ;
	assign x_351 = ((~v_4 | ~v_60) | v_773) ;
	assign x_350 = (v_774 | ~v_23) ;
	assign x_349 = (v_774 | ~v_24) ;
	assign x_348 = (v_774 | ~v_25) ;
	assign x_347 = (v_774 | ~v_26) ;
	assign x_346 = (v_774 | ~v_27) ;
	assign x_345 = (v_774 | ~v_53) ;
	assign x_344 = (v_774 | ~v_70) ;
	assign x_343 = (v_774 | ~v_773) ;
	assign x_342 = (v_774 | ~v_772) ;
	assign x_341 = (v_774 | ~v_573) ;
	assign x_339 = (v_774 | ~v_723) ;
	assign x_338 = (v_774 | ~v_722) ;
	assign x_337 = (v_774 | ~v_771) ;
	assign x_336 = (v_774 | ~v_770) ;
	assign x_335 = ((~v_45 | ~v_59) | v_775) ;
	assign x_334 = ((~v_42 | v_59) | v_776) ;
	assign x_333 = ((~v_3 | v_60) | v_777) ;
	assign x_332 = ((~v_6 | ~v_60) | v_778) ;
	assign x_331 = (v_779 | ~v_36) ;
	assign x_330 = (v_779 | ~v_37) ;
	assign x_329 = (v_779 | ~v_38) ;
	assign x_328 = (v_779 | ~v_39) ;
	assign x_327 = (v_779 | ~v_40) ;
	assign x_326 = (v_779 | ~v_56) ;
	assign x_324 = (v_779 | ~v_778) ;
	assign x_323 = (v_779 | ~v_777) ;
	assign x_322 = (v_779 | ~v_776) ;
	assign x_321 = (v_779 | ~v_582) ;
	assign x_320 = (v_779 | ~v_581) ;
	assign x_319 = (v_779 | ~v_729) ;
	assign x_318 = (v_779 | ~v_728) ;
	assign x_317 = (v_779 | ~v_775) ;
	assign x_316 = (((~v_779 | ~v_774) | ~v_769) | v_780) ;
	assign x_315 = ((~v_1 | v_50) | v_781) ;
	assign x_314 = ((~v_16 | v_51) | v_782) ;
	assign x_313 = ((~v_5 | ~v_50) | v_783) ;
	assign x_312 = ((~v_19 | ~v_51) | v_784) ;
	assign x_311 = (v_785 | ~v_8) ;
	assign x_309 = (v_785 | ~v_11) ;
	assign x_308 = (v_785 | ~v_13) ;
	assign x_307 = (v_785 | ~v_47) ;
	assign x_306 = (v_785 | ~v_48) ;
	assign x_305 = (v_785 | ~v_49) ;
	assign x_304 = (v_785 | ~v_784) ;
	assign x_302 = (v_785 | ~v_677) ;
	assign x_301 = (v_785 | ~v_639) ;
	assign x_300 = (v_785 | ~v_638) ;
	assign x_299 = (v_785 | ~v_783) ;
	assign x_298 = (v_785 | ~v_782) ;
	assign x_297 = (v_785 | ~v_781) ;
	assign x_295 = ((~v_29 | v_51) | v_787) ;
	assign x_294 = ((~v_4 | ~v_50) | v_788) ;
	assign x_293 = ((~v_32 | ~v_51) | v_789) ;
	assign x_292 = (v_790 | ~v_22) ;
	assign x_291 = (v_790 | ~v_24) ;
	assign x_290 = (v_790 | ~v_25) ;
	assign x_289 = (v_790 | ~v_27) ;
	assign x_288 = (v_790 | ~v_53) ;
	assign x_287 = (v_790 | ~v_54) ;
	assign x_286 = (v_790 | ~v_55) ;
	assign x_285 = (v_790 | ~v_789) ;
	assign x_284 = (v_790 | ~v_647) ;
	assign x_283 = (v_790 | ~v_646) ;
	assign x_282 = (v_790 | ~v_685) ;
	assign x_280 = (v_790 | ~v_788) ;
	assign x_279 = (v_790 | ~v_787) ;
	assign x_278 = (v_790 | ~v_786) ;
	assign x_277 = ((~v_3 | v_50) | v_791) ;
	assign x_276 = ((~v_42 | v_51) | v_792) ;
	assign x_275 = ((~v_6 | ~v_50) | v_793) ;
	assign x_274 = ((~v_45 | ~v_51) | v_794) ;
	assign x_273 = (v_795 | ~v_35) ;
	assign x_272 = (v_795 | ~v_37) ;
	assign x_271 = (v_795 | ~v_38) ;
	assign x_270 = (v_795 | ~v_40) ;
	assign x_269 = (v_795 | ~v_56) ;
	assign x_268 = (v_795 | ~v_57) ;
	assign x_267 = (v_795 | ~v_58) ;
	assign x_265 = (v_795 | ~v_793) ;
	assign x_264 = (v_795 | ~v_691) ;
	assign x_263 = (v_795 | ~v_653) ;
	assign x_262 = (v_795 | ~v_652) ;
	assign x_261 = (v_795 | ~v_690) ;
	assign x_260 = (v_795 | ~v_792) ;
	assign x_259 = (v_795 | ~v_791) ;
	assign x_258 = (((~v_795 | ~v_790) | ~v_785) | v_796) ;
	assign x_257 = ((~v_16 | v_52) | v_797) ;
	assign x_256 = ((~v_19 | ~v_52) | v_798) ;
	assign x_255 = ((~v_1 | v_52) | v_799) ;
	assign x_254 = ((~v_5 | ~v_52) | v_800) ;
	assign x_253 = (v_801 | ~v_7) ;
	assign x_252 = (v_801 | ~v_10) ;
	assign x_250 = (v_801 | ~v_12) ;
	assign x_249 = (v_801 | ~v_13) ;
	assign x_248 = (v_801 | ~v_48) ;
	assign x_247 = (v_801 | ~v_68) ;
	assign x_246 = (v_801 | ~v_800) ;
	assign x_245 = (v_801 | ~v_799) ;
	assign x_243 = (v_801 | ~v_639) ;
	assign x_242 = (v_801 | ~v_638) ;
	assign x_241 = (v_801 | ~v_616) ;
	assign x_240 = (v_801 | ~v_798) ;
	assign x_239 = (v_801 | ~v_797) ;
	assign x_238 = ((~v_29 | v_52) | v_802) ;
	assign x_236 = ((~v_4 | ~v_52) | v_804) ;
	assign x_235 = ((~v_32 | ~v_52) | v_805) ;
	assign x_234 = (v_806 | ~v_21) ;
	assign x_233 = (v_806 | ~v_24) ;
	assign x_232 = (v_806 | ~v_25) ;
	assign x_231 = (v_806 | ~v_26) ;
	assign x_230 = (v_806 | ~v_27) ;
	assign x_229 = (v_806 | ~v_54) ;
	assign x_228 = (v_806 | ~v_70) ;
	assign x_227 = (v_806 | ~v_805) ;
	assign x_226 = (v_806 | ~v_804) ;
	assign x_225 = (v_806 | ~v_803) ;
	assign x_224 = (v_806 | ~v_625) ;
	assign x_223 = (v_806 | ~v_647) ;
	assign x_221 = (v_806 | ~v_624) ;
	assign x_220 = (v_806 | ~v_802) ;
	assign x_219 = ((~v_42 | v_52) | v_807) ;
	assign x_218 = ((~v_45 | ~v_52) | v_808) ;
	assign x_217 = ((~v_3 | v_52) | v_809) ;
	assign x_216 = ((~v_6 | ~v_52) | v_810) ;
	assign x_215 = (v_811 | ~v_34) ;
	assign x_214 = (v_811 | ~v_37) ;
	assign x_213 = (v_811 | ~v_38) ;
	assign x_212 = (v_811 | ~v_39) ;
	assign x_211 = (v_811 | ~v_40) ;
	assign x_210 = (v_811 | ~v_57) ;
	assign x_209 = (v_811 | ~v_72) ;
	assign x_208 = (v_811 | ~v_810) ;
	assign x_206 = (v_811 | ~v_653) ;
	assign x_205 = (v_811 | ~v_652) ;
	assign x_204 = (v_811 | ~v_632) ;
	assign x_203 = (v_811 | ~v_631) ;
	assign x_202 = (v_811 | ~v_808) ;
	assign x_201 = (v_811 | ~v_807) ;
	assign x_200 = (((~v_811 | ~v_806) | ~v_801) | v_812) ;
	assign x_199 = ((~v_16 | v_50) | v_813) ;
	assign x_198 = ((~v_19 | ~v_50) | v_814) ;
	assign x_197 = ((~v_1 | v_51) | v_815) ;
	assign x_196 = ((~v_5 | ~v_51) | v_816) ;
	assign x_195 = (v_817 | ~v_9) ;
	assign x_194 = (v_817 | ~v_10) ;
	assign x_193 = (v_817 | ~v_11) ;
	assign x_191 = (v_817 | ~v_47) ;
	assign x_190 = (v_817 | ~v_68) ;
	assign x_189 = (v_817 | ~v_69) ;
	assign x_188 = (v_817 | ~v_816) ;
	assign x_187 = (v_817 | ~v_815) ;
	assign x_186 = (v_817 | ~v_814) ;
	assign x_184 = (v_817 | ~v_716) ;
	assign x_183 = (v_817 | ~v_715) ;
	assign x_182 = (v_817 | ~v_616) ;
	assign x_181 = (v_817 | ~v_813) ;
	assign x_180 = ((~v_29 | v_50) | v_818) ;
	assign x_179 = ((~v_32 | ~v_50) | v_819) ;
	assign x_177 = ((~v_4 | ~v_51) | v_821) ;
	assign x_176 = (v_822 | ~v_23) ;
	assign x_175 = (v_822 | ~v_24) ;
	assign x_174 = (v_822 | ~v_25) ;
	assign x_173 = (v_822 | ~v_26) ;
	assign x_172 = (v_822 | ~v_53) ;
	assign x_171 = (v_822 | ~v_70) ;
	assign x_170 = (v_822 | ~v_71) ;
	assign x_169 = (v_822 | ~v_821) ;
	assign x_168 = (v_822 | ~v_820) ;
	assign x_167 = (v_822 | ~v_819) ;
	assign x_166 = (v_822 | ~v_625) ;
	assign x_165 = (v_822 | ~v_723) ;
	assign x_164 = (v_822 | ~v_722) ;
	assign x_162 = (v_822 | ~v_624) ;
	assign x_161 = ((~v_42 | v_50) | v_823) ;
	assign x_160 = ((~v_45 | ~v_50) | v_824) ;
	assign x_159 = ((~v_3 | v_51) | v_825) ;
	assign x_158 = ((~v_6 | ~v_51) | v_826) ;
	assign x_157 = (v_827 | ~v_36) ;
	assign x_156 = (v_827 | ~v_37) ;
	assign x_155 = (v_827 | ~v_38) ;
	assign x_154 = (v_827 | ~v_39) ;
	assign x_153 = (v_827 | ~v_56) ;
	assign x_152 = (v_827 | ~v_72) ;
	assign x_151 = (v_827 | ~v_73) ;
	assign x_150 = (v_827 | ~v_826) ;
	assign x_149 = (v_827 | ~v_825) ;
	assign x_147 = (v_827 | ~v_728) ;
	assign x_146 = (v_827 | ~v_824) ;
	assign x_145 = (v_827 | ~v_632) ;
	assign x_144 = (v_827 | ~v_823) ;
	assign x_143 = (v_827 | ~v_631) ;
	assign x_142 = (((~v_827 | ~v_822) | ~v_817) | v_828) ;
	assign x_141 = ((~v_16 | v_14) | v_829) ;
	assign x_140 = ((~v_14 | ~v_19) | v_830) ;
	assign x_139 = ((~v_5 | ~v_14) | v_831) ;
	assign x_138 = ((~v_1 | v_14) | v_832) ;
	assign x_137 = (v_833 | ~v_7) ;
	assign x_136 = (v_833 | ~v_8) ;
	assign x_135 = (v_833 | ~v_9) ;
	assign x_134 = (v_833 | ~v_10) ;
	assign x_132 = (v_833 | ~v_12) ;
	assign x_131 = (v_833 | ~v_13) ;
	assign x_130 = (v_833 | ~v_832) ;
	assign x_129 = (v_833 | ~v_831) ;
	assign x_128 = (v_833 | ~v_678) ;
	assign x_127 = (v_833 | ~v_677) ;
	assign x_125 = (v_833 | ~v_830) ;
	assign x_124 = (v_833 | ~v_715) ;
	assign x_123 = (v_833 | ~v_829) ;
	assign x_122 = ((~v_29 | v_14) | v_834) ;
	assign x_121 = ((~v_14 | ~v_32) | v_835) ;
	assign x_120 = ((~v_4 | ~v_14) | v_836) ;
	assign x_118 = (v_838 | ~v_21) ;
	assign x_117 = (v_838 | ~v_22) ;
	assign x_116 = (v_838 | ~v_23) ;
	assign x_115 = (v_838 | ~v_24) ;
	assign x_114 = (v_838 | ~v_25) ;
	assign x_113 = (v_838 | ~v_26) ;
	assign x_112 = (v_838 | ~v_27) ;
	assign x_111 = (v_838 | ~v_837) ;
	assign x_110 = (v_838 | ~v_836) ;
	assign x_109 = (v_838 | ~v_723) ;
	assign x_108 = (v_838 | ~v_835) ;
	assign x_107 = (v_838 | ~v_685) ;
	assign x_106 = (v_838 | ~v_722) ;
	assign x_105 = (v_838 | ~v_834) ;
	assign x_103 = ((v_14 | ~v_42) | v_839) ;
	assign x_102 = ((~v_14 | ~v_45) | v_840) ;
	assign x_101 = ((~v_6 | ~v_14) | v_841) ;
	assign x_100 = ((~v_3 | v_14) | v_842) ;
	assign x_99 = (v_843 | ~v_34) ;
	assign x_98 = (v_843 | ~v_35) ;
	assign x_97 = (v_843 | ~v_36) ;
	assign x_96 = (v_843 | ~v_37) ;
	assign x_95 = (v_843 | ~v_38) ;
	assign x_94 = (v_843 | ~v_39) ;
	assign x_93 = (v_843 | ~v_40) ;
	assign x_92 = (v_843 | ~v_842) ;
	assign x_91 = (v_843 | ~v_841) ;
	assign x_90 = (v_843 | ~v_691) ;
	assign x_88 = (v_843 | ~v_729) ;
	assign x_87 = (v_843 | ~v_728) ;
	assign x_86 = (v_843 | ~v_839) ;
	assign x_85 = (v_843 | ~v_690) ;
	assign x_84 = (((~v_843 | ~v_838) | ~v_833) | v_844) ;
	assign x_83 = ((~v_16 | v_74) | v_845) ;
	assign x_82 = ((~v_19 | ~v_74) | v_846) ;
	assign x_81 = ((~v_5 | ~v_75) | v_847) ;
	assign x_80 = ((~v_1 | v_75) | v_848) ;
	assign x_79 = (v_849 | ~v_10) ;
	assign x_78 = (v_849 | ~v_11) ;
	assign x_77 = (v_849 | ~v_12) ;
	assign x_76 = (v_849 | ~v_47) ;
	assign x_75 = (v_849 | ~v_48) ;
	assign x_73 = (v_849 | ~v_69) ;
	assign x_72 = (v_849 | ~v_564) ;
	assign x_71 = (v_849 | ~v_848) ;
	assign x_70 = (v_849 | ~v_847) ;
	assign x_69 = (v_849 | ~v_846) ;
	assign x_68 = (v_849 | ~v_845) ;
	assign x_66 = (v_849 | ~v_639) ;
	assign x_65 = (v_849 | ~v_638) ;
	assign x_64 = ((~v_29 | v_74) | v_850) ;
	assign x_63 = ((~v_32 | ~v_74) | v_851) ;
	assign x_62 = ((~v_4 | ~v_75) | v_852) ;
	assign x_61 = ((~v_2 | v_75) | v_853) ;
	assign x_59 = (v_854 | ~v_25) ;
	assign x_58 = (v_854 | ~v_26) ;
	assign x_57 = (v_854 | ~v_53) ;
	assign x_56 = (v_854 | ~v_54) ;
	assign x_55 = (v_854 | ~v_70) ;
	assign x_54 = (v_854 | ~v_71) ;
	assign x_53 = (v_854 | ~v_573) ;
	assign x_52 = (v_854 | ~v_853) ;
	assign x_51 = (v_854 | ~v_852) ;
	assign x_50 = (v_854 | ~v_572) ;
	assign x_49 = (v_854 | ~v_851) ;
	assign x_48 = (v_854 | ~v_850) ;
	assign x_47 = (v_854 | ~v_647) ;
	assign x_46 = (v_854 | ~v_646) ;
	assign x_44 = ((~v_45 | ~v_74) | v_856) ;
	assign x_43 = ((~v_6 | ~v_75) | v_857) ;
	assign x_42 = ((~v_3 | v_75) | v_858) ;
	assign x_41 = (v_859 | ~v_37) ;
	assign x_40 = (v_859 | ~v_38) ;
	assign x_39 = (v_859 | ~v_39) ;
	assign x_38 = (v_859 | ~v_56) ;
	assign x_37 = (v_859 | ~v_57) ;
	assign x_36 = (v_859 | ~v_72) ;
	assign x_35 = (v_859 | ~v_73) ;
	assign x_34 = (v_859 | ~v_582) ;
	assign x_33 = (v_859 | ~v_858) ;
	assign x_32 = (v_859 | ~v_857) ;
	assign x_31 = (v_859 | ~v_856) ;
	assign x_29 = (v_859 | ~v_581) ;
	assign x_28 = (v_859 | ~v_653) ;
	assign x_27 = (v_859 | ~v_652) ;
	assign x_26 = (((~v_859 | ~v_854) | ~v_849) | v_860) ;
	assign x_25 = ((~v_2 | v_1) | v_861) ;
	assign x_24 = ((~v_3 | v_2) | v_862) ;
	assign x_23 = ((~v_4 | v_6) | v_863) ;
	assign x_22 = ((~v_5 | v_4) | v_864) ;
	assign x_21 = (v_865 | ~v_864) ;
	assign x_20 = (v_865 | ~v_863) ;
	assign x_19 = (v_865 | ~v_862) ;
	assign x_18 = (v_865 | ~v_861) ;
	assign x_17 = (v_865 | ~v_860) ;
	assign x_16 = (v_865 | ~v_844) ;
	assign x_14 = (v_865 | ~v_812) ;
	assign x_13 = (v_865 | ~v_796) ;
	assign x_12 = (v_865 | ~v_780) ;
	assign x_11 = (v_865 | ~v_764) ;
	assign x_10 = (v_865 | ~v_748) ;
	assign x_9 = (v_865 | ~v_732) ;
	assign x_7 = (v_865 | ~v_694) ;
	assign x_6 = (v_865 | ~v_672) ;
	assign x_5 = (v_865 | ~v_656) ;
	assign x_4 = (v_865 | ~v_634) ;
	assign x_3 = (v_865 | ~v_612) ;
	assign x_2 = (v_865 | ~v_584) ;
	assign x_3773 = (x_1891 & x_1892) ;
	assign x_3772 = (x_1889 & x_1890) ;
	assign x_3770 = (x_1887 & x_1888) ;
	assign x_3769 = (x_1885 & x_1886) ;
	assign x_3766 = (x_1883 & x_1884) ;
	assign x_3765 = (x_1881 & x_1882) ;
	assign x_3763 = (x_1879 & x_1880) ;
	assign x_1878 = (v_91 | v_76) ;
	assign x_3759 = (x_1876 & x_1877) ;
	assign x_3758 = (x_1874 & x_1875) ;
	assign x_3756 = (x_1872 & x_1873) ;
	assign x_3755 = (x_1870 & x_1871) ;
	assign x_3752 = (x_1868 & x_1869) ;
	assign x_3751 = (x_1866 & x_1867) ;
	assign x_3749 = (x_1864 & x_1865) ;
	assign x_1863 = (v_99 | v_74) ;
	assign x_3744 = (x_1861 & x_1862) ;
	assign x_3743 = (x_1859 & x_1860) ;
	assign x_3741 = (x_1857 & x_1858) ;
	assign x_3740 = (x_1855 & x_1856) ;
	assign x_3737 = (x_1853 & x_1854) ;
	assign x_3736 = (x_1851 & x_1852) ;
	assign x_3734 = (x_1849 & x_1850) ;
	assign x_1848 = (v_108 | ~v_85) ;
	assign x_3730 = (x_1846 & x_1847) ;
	assign x_3729 = (x_1844 & x_1845) ;
	assign x_3727 = (x_1842 & x_1843) ;
	assign x_3726 = (x_1840 & x_1841) ;
	assign x_3723 = (x_1838 & x_1839) ;
	assign x_3722 = (x_1836 & x_1837) ;
	assign x_3720 = (x_1834 & x_1835) ;
	assign x_1833 = (v_117 | ~v_116) ;
	assign x_3714 = (x_1831 & x_1832) ;
	assign x_3713 = (x_1829 & x_1830) ;
	assign x_3711 = (x_1827 & x_1828) ;
	assign x_3710 = (x_1825 & x_1826) ;
	assign x_3707 = (x_1823 & x_1824) ;
	assign x_3706 = (x_1821 & x_1822) ;
	assign x_3704 = (x_1819 & x_1820) ;
	assign x_1818 = (v_126 | v_51) ;
	assign x_3700 = (x_1816 & x_1817) ;
	assign x_3699 = (x_1814 & x_1815) ;
	assign x_3697 = (x_1812 & x_1813) ;
	assign x_3696 = (x_1810 & x_1811) ;
	assign x_3693 = (x_1808 & x_1809) ;
	assign x_3692 = (x_1806 & x_1807) ;
	assign x_3690 = (x_1804 & x_1805) ;
	assign x_1803 = (v_134 | v_77) ;
	assign x_3685 = (x_1801 & x_1802) ;
	assign x_3684 = (x_1799 & x_1800) ;
	assign x_3682 = (x_1797 & x_1798) ;
	assign x_3681 = (x_1795 & x_1796) ;
	assign x_3678 = (x_1793 & x_1794) ;
	assign x_3677 = (x_1791 & x_1792) ;
	assign x_3675 = (x_1789 & x_1790) ;
	assign x_1788 = (v_144 | ~v_116) ;
	assign x_3671 = (x_1786 & x_1787) ;
	assign x_3670 = (x_1784 & x_1785) ;
	assign x_3668 = (x_1782 & x_1783) ;
	assign x_1781 = (v_148 | ~v_96) ;
	assign x_3665 = (x_1779 & x_1780) ;
	assign x_3664 = (x_1777 & x_1778) ;
	assign x_3662 = (x_1775 & x_1776) ;
	assign x_1774 = (((((v_60 | ~v_126) | ~v_125) | ~v_152) | ~v_151) | v_153) ;
	assign x_3655 = (x_1772 & x_1773) ;
	assign x_3654 = (x_1770 & x_1771) ;
	assign x_3652 = (x_1768 & x_1769) ;
	assign x_3651 = (x_1766 & x_1767) ;
	assign x_3648 = (x_1764 & x_1765) ;
	assign x_3647 = (x_1762 & x_1763) ;
	assign x_3645 = (x_1760 & x_1761) ;
	assign x_1759 = (v_162 | ~v_158) ;
	assign x_3641 = (x_1757 & x_1758) ;
	assign x_3640 = (x_1755 & x_1756) ;
	assign x_3638 = (x_1753 & x_1754) ;
	assign x_3637 = (x_1751 & x_1752) ;
	assign x_3634 = (x_1749 & x_1750) ;
	assign x_3633 = (x_1747 & x_1748) ;
	assign x_3631 = (x_1745 & x_1746) ;
	assign x_1744 = (v_170 | v_20) ;
	assign x_3626 = (x_1742 & x_1743) ;
	assign x_3625 = (x_1740 & x_1741) ;
	assign x_3623 = (x_1738 & x_1739) ;
	assign x_3622 = (x_1736 & x_1737) ;
	assign x_3619 = (x_1734 & x_1735) ;
	assign x_3618 = (x_1732 & x_1733) ;
	assign x_3616 = (x_1730 & x_1731) ;
	assign x_1729 = (v_178 | v_32) ;
	assign x_3612 = (x_1727 & x_1728) ;
	assign x_3611 = (x_1725 & x_1726) ;
	assign x_3609 = (x_1723 & x_1724) ;
	assign x_1722 = (v_181 | v_61) ;
	assign x_3606 = (x_1720 & x_1721) ;
	assign x_3605 = (x_1718 & x_1719) ;
	assign x_3603 = (x_1716 & x_1717) ;
	assign x_1715 = (v_185 | v_42) ;
	assign x_3597 = (x_1713 & x_1714) ;
	assign x_3596 = (x_1711 & x_1712) ;
	assign x_3594 = (x_1709 & x_1710) ;
	assign x_3593 = (x_1707 & x_1708) ;
	assign x_3590 = (x_1705 & x_1706) ;
	assign x_3589 = (x_1703 & x_1704) ;
	assign x_3587 = (x_1701 & x_1702) ;
	assign x_1700 = (v_193 | ~v_183) ;
	assign x_3583 = (x_1698 & x_1699) ;
	assign x_3582 = (x_1696 & x_1697) ;
	assign x_3580 = (x_1694 & x_1695) ;
	assign x_3579 = (x_1692 & x_1693) ;
	assign x_3576 = (x_1690 & x_1691) ;
	assign x_3575 = (x_1688 & x_1689) ;
	assign x_3573 = (x_1686 & x_1687) ;
	assign x_1685 = (v_200 | v_61) ;
	assign x_3568 = (x_1683 & x_1684) ;
	assign x_3567 = (x_1681 & x_1682) ;
	assign x_3565 = (x_1679 & x_1680) ;
	assign x_3564 = (x_1677 & x_1678) ;
	assign x_3561 = (x_1675 & x_1676) ;
	assign x_3560 = (x_1673 & x_1674) ;
	assign x_3558 = (x_1671 & x_1672) ;
	assign x_1670 = (v_208 | v_65) ;
	assign x_3554 = (x_1668 & x_1669) ;
	assign x_3553 = (x_1666 & x_1667) ;
	assign x_3551 = (x_1664 & x_1665) ;
	assign x_1663 = (v_212 | ~v_79) ;
	assign x_3548 = (x_1661 & x_1662) ;
	assign x_3547 = (x_1659 & x_1660) ;
	assign x_3545 = (x_1657 & x_1658) ;
	assign x_1656 = (v_216 | ~v_65) ;
	assign x_3537 = (x_1654 & x_1655) ;
	assign x_3536 = (x_1652 & x_1653) ;
	assign x_3534 = (x_1650 & x_1651) ;
	assign x_3533 = (x_1648 & x_1649) ;
	assign x_3530 = (x_1646 & x_1647) ;
	assign x_3529 = (x_1644 & x_1645) ;
	assign x_3527 = (x_1642 & x_1643) ;
	assign x_1641 = (v_223 | ~v_77) ;
	assign x_3523 = (x_1639 & x_1640) ;
	assign x_3522 = (x_1637 & x_1638) ;
	assign x_3520 = (x_1635 & x_1636) ;
	assign x_3519 = (x_1633 & x_1634) ;
	assign x_3516 = (x_1631 & x_1632) ;
	assign x_3515 = (x_1629 & x_1630) ;
	assign x_3513 = (x_1627 & x_1628) ;
	assign x_1626 = (v_231 | v_76) ;
	assign x_3508 = (x_1624 & x_1625) ;
	assign x_3507 = (x_1622 & x_1623) ;
	assign x_3505 = (x_1620 & x_1621) ;
	assign x_3504 = (x_1618 & x_1619) ;
	assign x_3501 = (x_1616 & x_1617) ;
	assign x_3500 = (x_1614 & x_1615) ;
	assign x_3498 = (x_1612 & x_1613) ;
	assign x_1611 = (v_239 | v_77) ;
	assign x_3494 = (x_1609 & x_1610) ;
	assign x_3493 = (x_1607 & x_1608) ;
	assign x_3491 = (x_1605 & x_1606) ;
	assign x_1604 = (v_243 | ~v_235) ;
	assign x_3488 = (x_1602 & x_1603) ;
	assign x_3487 = (x_1600 & x_1601) ;
	assign x_3485 = (x_1598 & x_1599) ;
	assign x_1597 = (v_246 | v_77) ;
	assign x_3479 = (x_1595 & x_1596) ;
	assign x_3478 = (x_1593 & x_1594) ;
	assign x_3476 = (x_1591 & x_1592) ;
	assign x_3475 = (x_1589 & x_1590) ;
	assign x_3472 = (x_1587 & x_1588) ;
	assign x_3471 = (x_1585 & x_1586) ;
	assign x_3469 = (x_1583 & x_1584) ;
	assign x_1582 = (v_254 | v_76) ;
	assign x_3465 = (x_1580 & x_1581) ;
	assign x_3464 = (x_1578 & x_1579) ;
	assign x_3462 = (x_1576 & x_1577) ;
	assign x_3461 = (x_1574 & x_1575) ;
	assign x_3458 = (x_1572 & x_1573) ;
	assign x_3457 = (x_1570 & x_1571) ;
	assign x_3455 = (x_1568 & x_1569) ;
	assign x_1567 = (v_262 | v_46) ;
	assign x_3450 = (x_1565 & x_1566) ;
	assign x_3449 = (x_1563 & x_1564) ;
	assign x_3447 = (x_1561 & x_1562) ;
	assign x_3446 = (x_1559 & x_1560) ;
	assign x_3443 = (x_1557 & x_1558) ;
	assign x_3442 = (x_1555 & x_1556) ;
	assign x_3440 = (x_1553 & x_1554) ;
	assign x_1552 = (((((((((((((((v_13 | v_11) | v_10) | v_68) | v_49) | v_48) | v_47) | ~v_269) | ~v_268) | ~v_227) | ~v_225) | ~v_200) | ~v_199) | ~v_267) | ~v_266) | v_270) ;
	assign x_3436 = (x_1550 & x_1551) ;
	assign x_3435 = (x_1548 & x_1549) ;
	assign x_3433 = (x_1546 & x_1547) ;
	assign x_1545 = (v_274 | v_29) ;
	assign x_3430 = (x_1543 & x_1544) ;
	assign x_3429 = (x_1541 & x_1542) ;
	assign x_3427 = (x_1539 & x_1540) ;
	assign x_1538 = (v_278 | v_6) ;
	assign x_3420 = (x_1536 & x_1537) ;
	assign x_3419 = (x_1534 & x_1535) ;
	assign x_3417 = (x_1532 & x_1533) ;
	assign x_3416 = (x_1530 & x_1531) ;
	assign x_3413 = (x_1528 & x_1529) ;
	assign x_3412 = (x_1526 & x_1527) ;
	assign x_3410 = (x_1524 & x_1525) ;
	assign x_1523 = (v_285 | v_64) ;
	assign x_3406 = (x_1521 & x_1522) ;
	assign x_3405 = (x_1519 & x_1520) ;
	assign x_3403 = (x_1517 & x_1518) ;
	assign x_3402 = (x_1515 & x_1516) ;
	assign x_3399 = (x_1513 & x_1514) ;
	assign x_3398 = (x_1511 & x_1512) ;
	assign x_3396 = (x_1509 & x_1510) ;
	assign x_1508 = (v_293 | v_28) ;
	assign x_3391 = (x_1506 & x_1507) ;
	assign x_3390 = (x_1504 & x_1505) ;
	assign x_3388 = (x_1502 & x_1503) ;
	assign x_3387 = (x_1500 & x_1501) ;
	assign x_3384 = (x_1498 & x_1499) ;
	assign x_3383 = (x_1496 & x_1497) ;
	assign x_3381 = (x_1494 & x_1495) ;
	assign x_1493 = (v_301 | v_63) ;
	assign x_3377 = (x_1491 & x_1492) ;
	assign x_3376 = (x_1489 & x_1490) ;
	assign x_3374 = (x_1487 & x_1488) ;
	assign x_1486 = (v_305 | v_16) ;
	assign x_3371 = (x_1484 & x_1485) ;
	assign x_3370 = (x_1482 & x_1483) ;
	assign x_3368 = (x_1480 & x_1481) ;
	assign x_1479 = (v_309 | v_2) ;
	assign x_3362 = (x_1477 & x_1478) ;
	assign x_3361 = (x_1475 & x_1476) ;
	assign x_3359 = (x_1473 & x_1474) ;
	assign x_3358 = (x_1471 & x_1472) ;
	assign x_3355 = (x_1469 & x_1470) ;
	assign x_3354 = (x_1467 & x_1468) ;
	assign x_3352 = (x_1465 & x_1466) ;
	assign x_1464 = (v_317 | v_6) ;
	assign x_3348 = (x_1462 & x_1463) ;
	assign x_3347 = (x_1460 & x_1461) ;
	assign x_3345 = (x_1458 & x_1459) ;
	assign x_3344 = (x_1456 & x_1457) ;
	assign x_3341 = (x_1454 & x_1455) ;
	assign x_3340 = (x_1452 & x_1453) ;
	assign x_3338 = (x_1450 & x_1451) ;
	assign x_1449 = (v_324 | v_17) ;
	assign x_3333 = (x_1447 & x_1448) ;
	assign x_3332 = (x_1445 & x_1446) ;
	assign x_3330 = (x_1443 & x_1444) ;
	assign x_3329 = (x_1441 & x_1442) ;
	assign x_3326 = (x_1439 & x_1440) ;
	assign x_3325 = (x_1437 & x_1438) ;
	assign x_3323 = (x_1435 & x_1436) ;
	assign x_1434 = (v_332 | v_33) ;
	assign x_3319 = (x_1432 & x_1433) ;
	assign x_3318 = (x_1430 & x_1431) ;
	assign x_3316 = (x_1428 & x_1429) ;
	assign x_1427 = (v_336 | v_63) ;
	assign x_3313 = (x_1425 & x_1426) ;
	assign x_3312 = (x_1423 & x_1424) ;
	assign x_3310 = (x_1421 & x_1422) ;
	assign x_1420 = (((((((((((((((v_39 | v_38) | v_36) | v_56) | v_40) | v_72) | v_82) | ~v_339) | ~v_338) | ~v_337) | ~v_336) | ~v_217) | ~v_335) | ~v_334) | ~v_216) | v_340) ;
	assign x_3301 = (x_1418 & x_1419) ;
	assign x_3300 = (x_1416 & x_1417) ;
	assign x_3298 = (x_1414 & x_1415) ;
	assign x_3297 = (x_1412 & x_1413) ;
	assign x_3294 = (x_1410 & x_1411) ;
	assign x_3293 = (x_1408 & x_1409) ;
	assign x_3291 = (x_1406 & x_1407) ;
	assign x_1405 = (v_348 | v_4) ;
	assign x_3287 = (x_1403 & x_1404) ;
	assign x_3286 = (x_1401 & x_1402) ;
	assign x_3284 = (x_1399 & x_1400) ;
	assign x_3283 = (x_1397 & x_1398) ;
	assign x_3280 = (x_1395 & x_1396) ;
	assign x_3279 = (x_1393 & x_1394) ;
	assign x_3277 = (x_1391 & x_1392) ;
	assign x_1390 = (((((((((((((((v_39 | v_38) | v_35) | v_37) | v_56) | v_40) | v_57) | ~v_355) | ~v_354) | ~v_353) | ~v_300) | ~v_299) | ~v_219) | ~v_218) | ~v_352) | v_356) ;
	assign x_3272 = (x_1388 & x_1389) ;
	assign x_3271 = (x_1386 & x_1387) ;
	assign x_3269 = (x_1384 & x_1385) ;
	assign x_3268 = (x_1382 & x_1383) ;
	assign x_3265 = (x_1380 & x_1381) ;
	assign x_3264 = (x_1378 & x_1379) ;
	assign x_3262 = (x_1376 & x_1377) ;
	assign x_1375 = (v_364 | v_32) ;
	assign x_3258 = (x_1373 & x_1374) ;
	assign x_3257 = (x_1371 & x_1372) ;
	assign x_3255 = (x_1369 & x_1370) ;
	assign x_3254 = (x_1367 & x_1368) ;
	assign x_3251 = (x_1365 & x_1366) ;
	assign x_3250 = (x_1363 & x_1364) ;
	assign x_3248 = (x_1361 & x_1362) ;
	assign x_1360 = (((((((((((((((v_39 | v_38) | v_37) | v_34) | v_40) | v_57) | v_72) | ~v_191) | ~v_371) | ~v_370) | ~v_190) | ~v_369) | ~v_368) | ~v_219) | ~v_218) | v_372) ;
	assign x_3242 = (x_1358 & x_1359) ;
	assign x_3241 = (x_1356 & x_1357) ;
	assign x_3239 = (x_1354 & x_1355) ;
	assign x_3238 = (x_1352 & x_1353) ;
	assign x_3235 = (x_1350 & x_1351) ;
	assign x_3234 = (x_1348 & x_1349) ;
	assign x_3232 = (x_1346 & x_1347) ;
	assign x_1345 = (v_380 | v_32) ;
	assign x_3228 = (x_1343 & x_1344) ;
	assign x_3227 = (x_1341 & x_1342) ;
	assign x_3225 = (x_1339 & x_1340) ;
	assign x_3224 = (x_1337 & x_1338) ;
	assign x_3221 = (x_1335 & x_1336) ;
	assign x_3220 = (x_1333 & x_1334) ;
	assign x_3218 = (x_1331 & x_1332) ;
	assign x_1330 = (((((((((((((((v_39 | v_38) | v_37) | v_36) | v_56) | v_40) | v_72) | ~v_387) | ~v_386) | ~v_385) | ~v_191) | ~v_190) | ~v_338) | ~v_337) | ~v_384) | v_388) ;
	assign x_3213 = (x_1328 & x_1329) ;
	assign x_3212 = (x_1326 & x_1327) ;
	assign x_3210 = (x_1324 & x_1325) ;
	assign x_3209 = (x_1322 & x_1323) ;
	assign x_3206 = (x_1320 & x_1321) ;
	assign x_3205 = (x_1318 & x_1319) ;
	assign x_3203 = (x_1316 & x_1317) ;
	assign x_1315 = (v_396 | v_29) ;
	assign x_3199 = (x_1313 & x_1314) ;
	assign x_3198 = (x_1311 & x_1312) ;
	assign x_3196 = (x_1309 & x_1310) ;
	assign x_1308 = (v_400 | v_3) ;
	assign x_3193 = (x_1306 & x_1307) ;
	assign x_3192 = (x_1304 & x_1305) ;
	assign x_3190 = (x_1302 & x_1303) ;
	assign x_1301 = (v_403 | v_45) ;
	assign x_3183 = (x_1299 & x_1300) ;
	assign x_3182 = (x_1297 & x_1298) ;
	assign x_3180 = (x_1295 & x_1296) ;
	assign x_3179 = (x_1293 & x_1294) ;
	assign x_3176 = (x_1291 & x_1292) ;
	assign x_3175 = (x_1289 & x_1290) ;
	assign x_3173 = (x_1287 & x_1288) ;
	assign x_1286 = (v_411 | ~v_52) ;
	assign x_3169 = (x_1284 & x_1285) ;
	assign x_3168 = (x_1282 & x_1283) ;
	assign x_3166 = (x_1280 & x_1281) ;
	assign x_3165 = (x_1278 & x_1279) ;
	assign x_3162 = (x_1276 & x_1277) ;
	assign x_3161 = (x_1274 & x_1275) ;
	assign x_3159 = (x_1272 & x_1273) ;
	assign x_1271 = (v_419 | ~v_52) ;
	assign x_3154 = (x_1269 & x_1270) ;
	assign x_3153 = (x_1267 & x_1268) ;
	assign x_3151 = (x_1265 & x_1266) ;
	assign x_3150 = (x_1263 & x_1264) ;
	assign x_3147 = (x_1261 & x_1262) ;
	assign x_3146 = (x_1259 & x_1260) ;
	assign x_3144 = (x_1257 & x_1258) ;
	assign x_1256 = (v_427 | ~v_50) ;
	assign x_3140 = (x_1254 & x_1255) ;
	assign x_3139 = (x_1252 & x_1253) ;
	assign x_3137 = (x_1250 & x_1251) ;
	assign x_1249 = (((((((((((((((v_25 | v_24) | v_23) | v_26) | v_53) | v_71) | v_70) | ~v_430) | ~v_429) | ~v_428) | ~v_234) | ~v_332) | ~v_331) | ~v_427) | ~v_233) | v_431) ;
	assign x_3134 = (x_1247 & x_1248) ;
	assign x_3133 = (x_1245 & x_1246) ;
	assign x_3131 = (x_1243 & x_1244) ;
	assign x_1242 = (v_435 | v_6) ;
	assign x_3125 = (x_1240 & x_1241) ;
	assign x_3124 = (x_1238 & x_1239) ;
	assign x_3122 = (x_1236 & x_1237) ;
	assign x_3121 = (x_1234 & x_1235) ;
	assign x_3118 = (x_1232 & x_1233) ;
	assign x_3117 = (x_1230 & x_1231) ;
	assign x_3115 = (x_1228 & x_1229) ;
	assign x_1227 = (v_443 | ~v_14) ;
	assign x_3111 = (x_1225 & x_1226) ;
	assign x_3110 = (x_1223 & x_1224) ;
	assign x_3108 = (x_1221 & x_1222) ;
	assign x_3107 = (x_1219 & x_1220) ;
	assign x_3104 = (x_1217 & x_1218) ;
	assign x_3103 = (x_1215 & x_1216) ;
	assign x_3101 = (x_1213 & x_1214) ;
	assign x_1212 = (v_451 | v_6) ;
	assign x_3096 = (x_1210 & x_1211) ;
	assign x_3095 = (x_1208 & x_1209) ;
	assign x_3093 = (x_1206 & x_1207) ;
	assign x_3092 = (x_1204 & x_1205) ;
	assign x_3089 = (x_1202 & x_1203) ;
	assign x_3088 = (x_1200 & x_1201) ;
	assign x_3086 = (x_1198 & x_1199) ;
	assign x_1197 = (v_459 | v_29) ;
	assign x_3082 = (x_1195 & x_1196) ;
	assign x_3081 = (x_1193 & x_1194) ;
	assign x_3079 = (x_1191 & x_1192) ;
	assign x_1190 = (v_462 | v_75) ;
	assign x_3076 = (x_1188 & x_1189) ;
	assign x_3075 = (x_1186 & x_1187) ;
	assign x_3073 = (x_1184 & x_1185) ;
	assign x_1183 = (v_466 | ~v_75) ;
	assign x_3065 = (x_1181 & x_1182) ;
	assign x_3064 = (x_1179 & x_1180) ;
	assign x_3062 = (x_1177 & x_1178) ;
	assign x_3061 = (x_1175 & x_1176) ;
	assign x_3058 = (x_1173 & x_1174) ;
	assign x_3057 = (x_1171 & x_1172) ;
	assign x_3055 = (x_1169 & x_1170) ;
	assign x_1168 = ((((((((((((((((((((~v_473 | ~v_472) | ~v_471) | ~v_470) | ~v_469) | ~v_453) | ~v_437) | ~v_421) | ~v_405) | ~v_389) | ~v_373) | ~v_357) | ~v_341) | ~v_319) | ~v_303) | ~v_281) | ~v_265) | ~v_243) | ~v_221) | ~v_193) | ~v_165) ;
	assign x_3051 = (x_1166 & x_1167) ;
	assign x_3050 = (x_1164 & x_1165) ;
	assign x_3048 = (x_1162 & x_1163) ;
	assign x_3047 = (x_1160 & x_1161) ;
	assign x_3044 = (x_1158 & x_1159) ;
	assign x_3043 = (x_1156 & x_1157) ;
	assign x_3041 = (x_1154 & x_1155) ;
	assign x_1153 = (v_485 | ~v_78) ;
	assign x_3036 = (x_1151 & x_1152) ;
	assign x_3035 = (x_1149 & x_1150) ;
	assign x_3033 = (x_1147 & x_1148) ;
	assign x_3032 = (x_1145 & x_1146) ;
	assign x_3029 = (x_1143 & x_1144) ;
	assign x_3028 = (x_1141 & x_1142) ;
	assign x_3026 = (x_1139 & x_1140) ;
	assign x_1138 = (v_492 | ~v_490) ;
	assign x_3022 = (x_1136 & x_1137) ;
	assign x_3021 = (x_1134 & x_1135) ;
	assign x_3019 = (x_1132 & x_1133) ;
	assign x_1131 = (v_496 | ~v_493) ;
	assign x_3016 = (x_1129 & x_1130) ;
	assign x_3015 = (x_1127 & x_1128) ;
	assign x_3013 = (x_1125 & x_1126) ;
	assign x_1124 = ((~v_51 | ~v_477) | v_500) ;
	assign x_3007 = (x_1122 & x_1123) ;
	assign x_3006 = (x_1120 & x_1121) ;
	assign x_3004 = (x_1118 & x_1119) ;
	assign x_3003 = (x_1116 & x_1117) ;
	assign x_3000 = (x_1114 & x_1115) ;
	assign x_2999 = (x_1112 & x_1113) ;
	assign x_2997 = (x_1110 & x_1111) ;
	assign x_1109 = (v_508 | ~v_507) ;
	assign x_2993 = (x_1107 & x_1108) ;
	assign x_2992 = (x_1105 & x_1106) ;
	assign x_2990 = (x_1103 & x_1104) ;
	assign x_2989 = (x_1101 & x_1102) ;
	assign x_2986 = (x_1099 & x_1100) ;
	assign x_2985 = (x_1097 & x_1098) ;
	assign x_2983 = (x_1095 & x_1096) ;
	assign x_1094 = (v_516 | ~v_515) ;
	assign x_2978 = (x_1092 & x_1093) ;
	assign x_2977 = (x_1090 & x_1091) ;
	assign x_2975 = (x_1088 & x_1089) ;
	assign x_2974 = (x_1086 & x_1087) ;
	assign x_2971 = (x_1084 & x_1085) ;
	assign x_2970 = (x_1082 & x_1083) ;
	assign x_2968 = (x_1080 & x_1081) ;
	assign x_1079 = ((~v_60 | ~v_79) | v_525) ;
	assign x_2964 = (x_1077 & x_1078) ;
	assign x_2963 = (x_1075 & x_1076) ;
	assign x_2961 = (x_1073 & x_1074) ;
	assign x_1072 = ((~v_527 | ~v_516) | v_528) ;
	assign x_2958 = (x_1070 & x_1071) ;
	assign x_2957 = (x_1068 & x_1069) ;
	assign x_2955 = (x_1066 & x_1067) ;
	assign x_1065 = (v_530 | ~v_494) ;
	assign x_2948 = (x_1063 & x_1064) ;
	assign x_2947 = (x_1061 & x_1062) ;
	assign x_2945 = (x_1059 & x_1060) ;
	assign x_2944 = (x_1057 & x_1058) ;
	assign x_2941 = (x_1055 & x_1056) ;
	assign x_2940 = (x_1053 & x_1054) ;
	assign x_2938 = (x_1051 & x_1052) ;
	assign x_1050 = (v_537 | ~v_502) ;
	assign x_2934 = (x_1048 & x_1049) ;
	assign x_2933 = (x_1046 & x_1047) ;
	assign x_2931 = (x_1044 & x_1045) ;
	assign x_2930 = (x_1042 & x_1043) ;
	assign x_2927 = (x_1040 & x_1041) ;
	assign x_2926 = (x_1038 & x_1039) ;
	assign x_2924 = (x_1036 & x_1037) ;
	assign x_1035 = ((~v_75 | ~v_523) | v_544) ;
	assign x_2919 = (x_1033 & x_1034) ;
	assign x_2918 = (x_1031 & x_1032) ;
	assign x_2916 = (x_1029 & x_1030) ;
	assign x_2915 = (x_1027 & x_1028) ;
	assign x_2912 = (x_1025 & x_1026) ;
	assign x_2911 = (x_1023 & x_1024) ;
	assign x_2909 = (x_1021 & x_1022) ;
	assign x_1020 = (v_550 | ~v_506) ;
	assign x_2905 = (x_1018 & x_1019) ;
	assign x_2904 = (x_1016 & x_1017) ;
	assign x_2902 = (x_1014 & x_1015) ;
	assign x_1013 = (v_553 | ~v_521) ;
	assign x_2899 = (x_1011 & x_1012) ;
	assign x_2898 = (x_1009 & x_1010) ;
	assign x_2896 = (x_1007 & x_1008) ;
	assign x_1006 = (v_555 | ~v_513) ;
	assign x_2890 = (x_1004 & x_1005) ;
	assign x_2889 = (x_1002 & x_1003) ;
	assign x_2887 = (x_1000 & x_1001) ;
	assign x_2886 = (x_998 & x_999) ;
	assign x_2883 = (x_996 & x_997) ;
	assign x_2882 = (x_994 & x_995) ;
	assign x_2880 = (x_992 & x_993) ;
	assign x_991 = (v_565 | ~v_47) ;
	assign x_2876 = (x_989 & x_990) ;
	assign x_2875 = (x_987 & x_988) ;
	assign x_2873 = (x_985 & x_986) ;
	assign x_2872 = (x_983 & x_984) ;
	assign x_2869 = (x_981 & x_982) ;
	assign x_2868 = (x_979 & x_980) ;
	assign x_2866 = (x_977 & x_978) ;
	assign x_976 = ((~v_4 | ~v_78) | v_568) ;
	assign x_2861 = (x_974 & x_975) ;
	assign x_2860 = (x_972 & x_973) ;
	assign x_2858 = (x_970 & x_971) ;
	assign x_2857 = (x_968 & x_969) ;
	assign x_2854 = (x_966 & x_967) ;
	assign x_2853 = (x_964 & x_965) ;
	assign x_2851 = (x_962 & x_963) ;
	assign x_961 = (v_574 | ~v_571) ;
	assign x_2847 = (x_959 & x_960) ;
	assign x_2846 = (x_957 & x_958) ;
	assign x_2844 = (x_955 & x_956) ;
	assign x_954 = ((~v_42 | v_79) | v_576) ;
	assign x_2841 = (x_952 & x_953) ;
	assign x_2840 = (x_950 & x_951) ;
	assign x_2838 = (x_948 & x_949) ;
	assign x_947 = (v_583 | ~v_37) ;
	assign x_2828 = (x_945 & x_946) ;
	assign x_2827 = (x_943 & x_944) ;
	assign x_2825 = (x_941 & x_942) ;
	assign x_2824 = (x_939 & x_940) ;
	assign x_2821 = (x_937 & x_938) ;
	assign x_2820 = (x_935 & x_936) ;
	assign x_2818 = (x_933 & x_934) ;
	assign x_932 = (((~v_583 | ~v_574) | ~v_565) | v_584) ;
	assign x_2814 = (x_930 & x_931) ;
	assign x_2813 = (x_928 & x_929) ;
	assign x_2811 = (x_926 & x_927) ;
	assign x_2810 = (x_924 & x_925) ;
	assign x_2807 = (x_922 & x_923) ;
	assign x_2806 = (x_920 & x_921) ;
	assign x_2804 = (x_918 & x_919) ;
	assign x_917 = (v_593 | ~v_80) ;
	assign x_2799 = (x_915 & x_916) ;
	assign x_2798 = (x_913 & x_914) ;
	assign x_2796 = (x_911 & x_912) ;
	assign x_2795 = (x_909 & x_910) ;
	assign x_2792 = (x_907 & x_908) ;
	assign x_2791 = (x_905 & x_906) ;
	assign x_2789 = (x_903 & x_904) ;
	assign x_902 = ((~v_30 | v_61) | v_600) ;
	assign x_2785 = (x_900 & x_901) ;
	assign x_2784 = (x_898 & x_899) ;
	assign x_2782 = (x_896 & x_897) ;
	assign x_2781 = (x_894 & x_895) ;
	assign x_2778 = (x_892 & x_893) ;
	assign x_2777 = (x_890 & x_891) ;
	assign x_2775 = (x_888 & x_889) ;
	assign x_887 = (v_602 | ~v_595) ;
	assign x_2769 = (x_885 & x_886) ;
	assign x_2768 = (x_883 & x_884) ;
	assign x_2766 = (x_881 & x_882) ;
	assign x_2765 = (x_879 & x_880) ;
	assign x_2762 = (x_877 & x_878) ;
	assign x_2761 = (x_875 & x_876) ;
	assign x_2759 = (x_873 & x_874) ;
	assign x_872 = (v_611 | ~v_73) ;
	assign x_2755 = (x_870 & x_871) ;
	assign x_2754 = (x_868 & x_869) ;
	assign x_2752 = (x_866 & x_867) ;
	assign x_2751 = (x_864 & x_865) ;
	assign x_2748 = (x_862 & x_863) ;
	assign x_2747 = (x_860 & x_861) ;
	assign x_2745 = (x_858 & x_859) ;
	assign x_857 = ((~v_19 | ~v_77) | v_617) ;
	assign x_2740 = (x_855 & x_856) ;
	assign x_2739 = (x_853 & x_854) ;
	assign x_2737 = (x_851 & x_852) ;
	assign x_2736 = (x_849 & x_850) ;
	assign x_2733 = (x_847 & x_848) ;
	assign x_2732 = (x_845 & x_846) ;
	assign x_2730 = (x_843 & x_844) ;
	assign x_842 = (v_619 | ~v_614) ;
	assign x_2726 = (x_840 & x_841) ;
	assign x_2725 = (x_838 & x_839) ;
	assign x_2723 = (x_836 & x_837) ;
	assign x_835 = ((~v_31 | ~v_52) | v_625) ;
	assign x_2720 = (x_833 & x_834) ;
	assign x_2719 = (x_831 & x_832) ;
	assign x_2717 = (x_829 & x_830) ;
	assign x_828 = (v_626 | ~v_70) ;
	assign x_2710 = (x_826 & x_827) ;
	assign x_2709 = (x_824 & x_825) ;
	assign x_2707 = (x_822 & x_823) ;
	assign x_2706 = (x_820 & x_821) ;
	assign x_2703 = (x_818 & x_819) ;
	assign x_2702 = (x_816 & x_817) ;
	assign x_2700 = (x_814 & x_815) ;
	assign x_813 = (v_633 | ~v_37) ;
	assign x_2696 = (x_811 & x_812) ;
	assign x_2695 = (x_809 & x_810) ;
	assign x_2693 = (x_807 & x_808) ;
	assign x_2692 = (x_805 & x_806) ;
	assign x_2689 = (x_803 & x_804) ;
	assign x_2688 = (x_801 & x_802) ;
	assign x_2686 = (x_799 & x_800) ;
	assign x_798 = (((~v_633 | ~v_626) | ~v_619) | v_634) ;
	assign x_2681 = (x_796 & x_797) ;
	assign x_2680 = (x_794 & x_795) ;
	assign x_2678 = (x_792 & x_793) ;
	assign x_2677 = (x_790 & x_791) ;
	assign x_2674 = (x_788 & x_789) ;
	assign x_2673 = (x_786 & x_787) ;
	assign x_2671 = (x_784 & x_785) ;
	assign x_783 = (v_641 | ~v_639) ;
	assign x_2667 = (x_781 & x_782) ;
	assign x_2666 = (x_779 & x_780) ;
	assign x_2664 = (x_777 & x_778) ;
	assign x_776 = ((~v_2 | v_77) | v_642) ;
	assign x_2661 = (x_774 & x_775) ;
	assign x_2660 = (x_772 & x_773) ;
	assign x_2658 = (x_770 & x_771) ;
	assign x_769 = (v_648 | ~v_26) ;
	assign x_2652 = (x_767 & x_768) ;
	assign x_2651 = (x_765 & x_766) ;
	assign x_2649 = (x_763 & x_764) ;
	assign x_2648 = (x_761 & x_762) ;
	assign x_2645 = (x_759 & x_760) ;
	assign x_2644 = (x_757 & x_758) ;
	assign x_2642 = (x_755 & x_756) ;
	assign x_754 = ((~v_42 | v_76) | v_650) ;
	assign x_2638 = (x_752 & x_753) ;
	assign x_2637 = (x_750 & x_751) ;
	assign x_2635 = (x_748 & x_749) ;
	assign x_2634 = (x_746 & x_747) ;
	assign x_2631 = (x_744 & x_745) ;
	assign x_2630 = (x_742 & x_743) ;
	assign x_2628 = (x_740 & x_741) ;
	assign x_739 = (v_655 | ~v_608) ;
	assign x_2623 = (x_737 & x_738) ;
	assign x_2622 = (x_735 & x_736) ;
	assign x_2620 = (x_733 & x_734) ;
	assign x_2619 = (x_731 & x_732) ;
	assign x_2616 = (x_729 & x_730) ;
	assign x_2615 = (x_727 & x_728) ;
	assign x_2613 = (x_725 & x_726) ;
	assign x_724 = (v_661 | ~v_49) ;
	assign x_2609 = (x_722 & x_723) ;
	assign x_2608 = (x_720 & x_721) ;
	assign x_2606 = (x_718 & x_719) ;
	assign x_717 = (v_661 | ~v_590) ;
	assign x_2603 = (x_715 & x_716) ;
	assign x_2602 = (x_713 & x_714) ;
	assign x_2600 = (x_711 & x_712) ;
	assign x_710 = (v_666 | ~v_24) ;
	assign x_2592 = (x_708 & x_709) ;
	assign x_2591 = (x_706 & x_707) ;
	assign x_2589 = (x_704 & x_705) ;
	assign x_2588 = (x_702 & x_703) ;
	assign x_2585 = (x_700 & x_701) ;
	assign x_2584 = (x_698 & x_699) ;
	assign x_2582 = (x_696 & x_697) ;
	assign x_695 = ((~v_3 | v_74) | v_667) ;
	assign x_2578 = (x_693 & x_694) ;
	assign x_2577 = (x_691 & x_692) ;
	assign x_2575 = (x_689 & x_690) ;
	assign x_2574 = (x_687 & x_688) ;
	assign x_2571 = (x_685 & x_686) ;
	assign x_2570 = (x_683 & x_684) ;
	assign x_2568 = (x_681 & x_682) ;
	assign x_680 = (v_671 | ~v_609) ;
	assign x_2563 = (x_678 & x_679) ;
	assign x_2562 = (x_676 & x_677) ;
	assign x_2560 = (x_674 & x_675) ;
	assign x_2559 = (x_672 & x_673) ;
	assign x_2556 = (x_670 & x_671) ;
	assign x_2555 = (x_668 & x_669) ;
	assign x_2553 = (x_666 & x_667) ;
	assign x_665 = (v_679 | ~v_47) ;
	assign x_2549 = (x_663 & x_664) ;
	assign x_2548 = (x_661 & x_662) ;
	assign x_2546 = (x_659 & x_660) ;
	assign x_658 = (v_679 | ~v_676) ;
	assign x_2543 = (x_656 & x_657) ;
	assign x_2542 = (x_654 & x_655) ;
	assign x_2540 = (x_652 & x_653) ;
	assign x_651 = ((~v_32 | ~v_64) | v_683) ;
	assign x_2534 = (x_649 & x_650) ;
	assign x_2533 = (x_647 & x_648) ;
	assign x_2531 = (x_645 & x_646) ;
	assign x_2530 = (x_643 & x_644) ;
	assign x_2527 = (x_641 & x_642) ;
	assign x_2526 = (x_639 & x_640) ;
	assign x_2524 = (x_637 & x_638) ;
	assign x_636 = (v_686 | ~v_682) ;
	assign x_2520 = (x_634 & x_635) ;
	assign x_2519 = (x_632 & x_633) ;
	assign x_2517 = (x_630 & x_631) ;
	assign x_2516 = (x_628 & x_629) ;
	assign x_2513 = (x_626 & x_627) ;
	assign x_2512 = (x_624 & x_625) ;
	assign x_2510 = (x_622 & x_623) ;
	assign x_621 = (v_693 | ~v_67) ;
	assign x_2505 = (x_619 & x_620) ;
	assign x_2504 = (x_617 & x_618) ;
	assign x_2502 = (x_615 & x_616) ;
	assign x_2501 = (x_613 & x_614) ;
	assign x_2498 = (x_611 & x_612) ;
	assign x_2497 = (x_609 & x_610) ;
	assign x_2495 = (x_607 & x_608) ;
	assign x_606 = (v_699 | ~v_12) ;
	assign x_2491 = (x_604 & x_605) ;
	assign x_2490 = (x_602 & x_603) ;
	assign x_2488 = (x_600 & x_601) ;
	assign x_599 = (v_699 | ~v_588) ;
	assign x_2485 = (x_597 & x_598) ;
	assign x_2484 = (x_595 & x_596) ;
	assign x_2482 = (x_593 & x_594) ;
	assign x_592 = ((~v_2 | v_65) | v_700) ;
	assign x_2475 = (x_590 & x_591) ;
	assign x_2474 = (x_588 & x_589) ;
	assign x_2472 = (x_586 & x_587) ;
	assign x_2471 = (x_584 & x_585) ;
	assign x_2468 = (x_582 & x_583) ;
	assign x_2467 = (x_580 & x_581) ;
	assign x_2465 = (x_578 & x_579) ;
	assign x_577 = (v_704 | ~v_701) ;
	assign x_2461 = (x_575 & x_576) ;
	assign x_2460 = (x_573 & x_574) ;
	assign x_2458 = (x_571 & x_572) ;
	assign x_2457 = (x_569 & x_570) ;
	assign x_2454 = (x_567 & x_568) ;
	assign x_2453 = (x_565 & x_566) ;
	assign x_2451 = (x_563 & x_564) ;
	assign x_562 = (v_709 | ~v_708) ;
	assign x_2446 = (x_560 & x_561) ;
	assign x_2445 = (x_558 & x_559) ;
	assign x_2443 = (x_556 & x_557) ;
	assign x_2442 = (x_554 & x_555) ;
	assign x_2439 = (x_552 & x_553) ;
	assign x_2438 = (x_550 & x_551) ;
	assign x_2436 = (x_548 & x_549) ;
	assign x_547 = (v_717 | ~v_9) ;
	assign x_2432 = (x_545 & x_546) ;
	assign x_2431 = (x_543 & x_544) ;
	assign x_2429 = (x_541 & x_542) ;
	assign x_540 = (v_717 | ~v_716) ;
	assign x_2426 = (x_538 & x_539) ;
	assign x_2425 = (x_536 & x_537) ;
	assign x_2423 = (x_534 & x_535) ;
	assign x_533 = (v_717 | ~v_588) ;
	assign x_2417 = (x_531 & x_532) ;
	assign x_2416 = (x_529 & x_530) ;
	assign x_2414 = (x_527 & x_528) ;
	assign x_2413 = (x_525 & x_526) ;
	assign x_2410 = (x_523 & x_524) ;
	assign x_2409 = (x_521 & x_522) ;
	assign x_2407 = (x_519 & x_520) ;
	assign x_518 = (v_724 | ~v_722) ;
	assign x_2403 = (x_516 & x_517) ;
	assign x_2402 = (x_514 & x_515) ;
	assign x_2400 = (x_512 & x_513) ;
	assign x_2399 = (x_510 & x_511) ;
	assign x_2396 = (x_508 & x_509) ;
	assign x_2395 = (x_506 & x_507) ;
	assign x_2393 = (x_504 & x_505) ;
	assign x_503 = (v_731 | ~v_39) ;
	assign x_2388 = (x_501 & x_502) ;
	assign x_2387 = (x_499 & x_500) ;
	assign x_2385 = (x_497 & x_498) ;
	assign x_2384 = (x_495 & x_496) ;
	assign x_2381 = (x_493 & x_494) ;
	assign x_2380 = (x_491 & x_492) ;
	assign x_2378 = (x_489 & x_490) ;
	assign x_488 = ((~v_1 | v_59) | v_734) ;
	assign x_2374 = (x_486 & x_487) ;
	assign x_2373 = (x_484 & x_485) ;
	assign x_2371 = (x_482 & x_483) ;
	assign x_481 = (v_737 | ~v_13) ;
	assign x_2368 = (x_479 & x_480) ;
	assign x_2367 = (x_477 & x_478) ;
	assign x_2365 = (x_475 & x_476) ;
	assign x_474 = (v_737 | ~v_733) ;
	assign x_2356 = (x_472 & x_473) ;
	assign x_2355 = (x_470 & x_471) ;
	assign x_2353 = (x_468 & x_469) ;
	assign x_2352 = (x_466 & x_467) ;
	assign x_2349 = (x_464 & x_465) ;
	assign x_2348 = (x_462 & x_463) ;
	assign x_2346 = (x_460 & x_461) ;
	assign x_459 = (v_742 | ~v_741) ;
	assign x_2342 = (x_457 & x_458) ;
	assign x_2341 = (x_455 & x_456) ;
	assign x_2339 = (x_453 & x_454) ;
	assign x_2338 = (x_451 & x_452) ;
	assign x_2335 = (x_449 & x_450) ;
	assign x_2334 = (x_447 & x_448) ;
	assign x_2332 = (x_445 & x_446) ;
	assign x_444 = (v_747 | ~v_39) ;
	assign x_2327 = (x_442 & x_443) ;
	assign x_2326 = (x_440 & x_441) ;
	assign x_2324 = (x_438 & x_439) ;
	assign x_2323 = (x_436 & x_437) ;
	assign x_2320 = (x_434 & x_435) ;
	assign x_2319 = (x_432 & x_433) ;
	assign x_2317 = (x_430 & x_431) ;
	assign x_429 = ((~v_5 | ~v_61) | v_751) ;
	assign x_2313 = (x_427 & x_428) ;
	assign x_2312 = (x_425 & x_426) ;
	assign x_2310 = (x_423 & x_424) ;
	assign x_2309 = (x_421 & x_422) ;
	assign x_2306 = (x_419 & x_420) ;
	assign x_2305 = (x_417 & x_418) ;
	assign x_2303 = (x_415 & x_416) ;
	assign x_414 = (v_753 | ~v_591) ;
	assign x_2297 = (x_412 & x_413) ;
	assign x_2296 = (x_410 & x_411) ;
	assign x_2294 = (x_408 & x_409) ;
	assign x_2293 = (x_406 & x_407) ;
	assign x_2290 = (x_404 & x_405) ;
	assign x_2289 = (x_402 & x_403) ;
	assign x_2287 = (x_400 & x_401) ;
	assign x_399 = (v_758 | ~v_756) ;
	assign x_2283 = (x_397 & x_398) ;
	assign x_2282 = (x_395 & x_396) ;
	assign x_2280 = (x_393 & x_394) ;
	assign x_2279 = (x_391 & x_392) ;
	assign x_2276 = (x_389 & x_390) ;
	assign x_2275 = (x_387 & x_388) ;
	assign x_2273 = (x_385 & x_386) ;
	assign x_384 = (v_763 | ~v_57) ;
	assign x_2268 = (x_382 & x_383) ;
	assign x_2267 = (x_380 & x_381) ;
	assign x_2265 = (x_378 & x_379) ;
	assign x_2264 = (x_376 & x_377) ;
	assign x_2261 = (x_374 & x_375) ;
	assign x_2260 = (x_372 & x_373) ;
	assign x_2258 = (x_370 & x_371) ;
	assign x_369 = (v_769 | ~v_9) ;
	assign x_2254 = (x_367 & x_368) ;
	assign x_2253 = (x_365 & x_366) ;
	assign x_2251 = (x_363 & x_364) ;
	assign x_362 = (v_769 | ~v_768) ;
	assign x_2248 = (x_360 & x_361) ;
	assign x_2247 = (x_358 & x_359) ;
	assign x_2245 = (x_356 & x_357) ;
	assign x_355 = (v_769 | ~v_765) ;
	assign x_2238 = (x_353 & x_354) ;
	assign x_2237 = (x_351 & x_352) ;
	assign x_2235 = (x_349 & x_350) ;
	assign x_2234 = (x_347 & x_348) ;
	assign x_2231 = (x_345 & x_346) ;
	assign x_2230 = (x_343 & x_344) ;
	assign x_2228 = (x_341 & x_342) ;
	assign x_340 = (v_774 | ~v_572) ;
	assign x_2224 = (x_338 & x_339) ;
	assign x_2223 = (x_336 & x_337) ;
	assign x_2221 = (x_334 & x_335) ;
	assign x_2220 = (x_332 & x_333) ;
	assign x_2217 = (x_330 & x_331) ;
	assign x_2216 = (x_328 & x_329) ;
	assign x_2214 = (x_326 & x_327) ;
	assign x_325 = (v_779 | ~v_72) ;
	assign x_2209 = (x_323 & x_324) ;
	assign x_2208 = (x_321 & x_322) ;
	assign x_2206 = (x_319 & x_320) ;
	assign x_2205 = (x_317 & x_318) ;
	assign x_2202 = (x_315 & x_316) ;
	assign x_2201 = (x_313 & x_314) ;
	assign x_2199 = (x_311 & x_312) ;
	assign x_310 = (v_785 | ~v_10) ;
	assign x_2195 = (x_308 & x_309) ;
	assign x_2194 = (x_306 & x_307) ;
	assign x_2192 = (x_304 & x_305) ;
	assign x_303 = (v_785 | ~v_678) ;
	assign x_2189 = (x_301 & x_302) ;
	assign x_2188 = (x_299 & x_300) ;
	assign x_2186 = (x_297 & x_298) ;
	assign x_296 = ((~v_2 | v_50) | v_786) ;
	assign x_2180 = (x_294 & x_295) ;
	assign x_2179 = (x_292 & x_293) ;
	assign x_2177 = (x_290 & x_291) ;
	assign x_2176 = (x_288 & x_289) ;
	assign x_2173 = (x_286 & x_287) ;
	assign x_2172 = (x_284 & x_285) ;
	assign x_2170 = (x_282 & x_283) ;
	assign x_281 = (v_790 | ~v_684) ;
	assign x_2166 = (x_279 & x_280) ;
	assign x_2165 = (x_277 & x_278) ;
	assign x_2163 = (x_275 & x_276) ;
	assign x_2162 = (x_273 & x_274) ;
	assign x_2159 = (x_271 & x_272) ;
	assign x_2158 = (x_269 & x_270) ;
	assign x_2156 = (x_267 & x_268) ;
	assign x_266 = (v_795 | ~v_794) ;
	assign x_2151 = (x_264 & x_265) ;
	assign x_2150 = (x_262 & x_263) ;
	assign x_2148 = (x_260 & x_261) ;
	assign x_2147 = (x_258 & x_259) ;
	assign x_2144 = (x_256 & x_257) ;
	assign x_2143 = (x_254 & x_255) ;
	assign x_2141 = (x_252 & x_253) ;
	assign x_251 = (v_801 | ~v_11) ;
	assign x_2137 = (x_249 & x_250) ;
	assign x_2136 = (x_247 & x_248) ;
	assign x_2134 = (x_245 & x_246) ;
	assign x_244 = (v_801 | ~v_618) ;
	assign x_2131 = (x_242 & x_243) ;
	assign x_2130 = (x_240 & x_241) ;
	assign x_2128 = (x_238 & x_239) ;
	assign x_237 = ((~v_2 | v_52) | v_803) ;
	assign x_2120 = (x_235 & x_236) ;
	assign x_2119 = (x_233 & x_234) ;
	assign x_2117 = (x_231 & x_232) ;
	assign x_2116 = (x_229 & x_230) ;
	assign x_2113 = (x_227 & x_228) ;
	assign x_2112 = (x_225 & x_226) ;
	assign x_2110 = (x_223 & x_224) ;
	assign x_222 = (v_806 | ~v_646) ;
	assign x_2106 = (x_220 & x_221) ;
	assign x_2105 = (x_218 & x_219) ;
	assign x_2103 = (x_216 & x_217) ;
	assign x_2102 = (x_214 & x_215) ;
	assign x_2099 = (x_212 & x_213) ;
	assign x_2098 = (x_210 & x_211) ;
	assign x_2096 = (x_208 & x_209) ;
	assign x_207 = (v_811 | ~v_809) ;
	assign x_2091 = (x_205 & x_206) ;
	assign x_2090 = (x_203 & x_204) ;
	assign x_2088 = (x_201 & x_202) ;
	assign x_2087 = (x_199 & x_200) ;
	assign x_2084 = (x_197 & x_198) ;
	assign x_2083 = (x_195 & x_196) ;
	assign x_2081 = (x_193 & x_194) ;
	assign x_192 = (v_817 | ~v_12) ;
	assign x_2077 = (x_190 & x_191) ;
	assign x_2076 = (x_188 & x_189) ;
	assign x_2074 = (x_186 & x_187) ;
	assign x_185 = (v_817 | ~v_618) ;
	assign x_2071 = (x_183 & x_184) ;
	assign x_2070 = (x_181 & x_182) ;
	assign x_2068 = (x_179 & x_180) ;
	assign x_178 = ((~v_2 | v_51) | v_820) ;
	assign x_2062 = (x_176 & x_177) ;
	assign x_2061 = (x_174 & x_175) ;
	assign x_2059 = (x_172 & x_173) ;
	assign x_2058 = (x_170 & x_171) ;
	assign x_2055 = (x_168 & x_169) ;
	assign x_2054 = (x_166 & x_167) ;
	assign x_2052 = (x_164 & x_165) ;
	assign x_163 = (v_822 | ~v_818) ;
	assign x_2048 = (x_161 & x_162) ;
	assign x_2047 = (x_159 & x_160) ;
	assign x_2045 = (x_157 & x_158) ;
	assign x_2044 = (x_155 & x_156) ;
	assign x_2041 = (x_153 & x_154) ;
	assign x_2040 = (x_151 & x_152) ;
	assign x_2038 = (x_149 & x_150) ;
	assign x_148 = (v_827 | ~v_729) ;
	assign x_2033 = (x_146 & x_147) ;
	assign x_2032 = (x_144 & x_145) ;
	assign x_2030 = (x_142 & x_143) ;
	assign x_2029 = (x_140 & x_141) ;
	assign x_2026 = (x_138 & x_139) ;
	assign x_2025 = (x_136 & x_137) ;
	assign x_2023 = (x_134 & x_135) ;
	assign x_133 = (v_833 | ~v_11) ;
	assign x_2019 = (x_131 & x_132) ;
	assign x_2018 = (x_129 & x_130) ;
	assign x_2016 = (x_127 & x_128) ;
	assign x_126 = (v_833 | ~v_716) ;
	assign x_2013 = (x_124 & x_125) ;
	assign x_2012 = (x_122 & x_123) ;
	assign x_2010 = (x_120 & x_121) ;
	assign x_119 = ((~v_2 | v_14) | v_837) ;
	assign x_2003 = (x_117 & x_118) ;
	assign x_2002 = (x_115 & x_116) ;
	assign x_2000 = (x_113 & x_114) ;
	assign x_1999 = (x_111 & x_112) ;
	assign x_1996 = (x_109 & x_110) ;
	assign x_1995 = (x_107 & x_108) ;
	assign x_1993 = (x_105 & x_106) ;
	assign x_104 = (v_838 | ~v_684) ;
	assign x_1989 = (x_102 & x_103) ;
	assign x_1988 = (x_100 & x_101) ;
	assign x_1986 = (x_98 & x_99) ;
	assign x_1985 = (x_96 & x_97) ;
	assign x_1982 = (x_94 & x_95) ;
	assign x_1981 = (x_92 & x_93) ;
	assign x_1979 = (x_90 & x_91) ;
	assign x_89 = (v_843 | ~v_840) ;
	assign x_1974 = (x_87 & x_88) ;
	assign x_1973 = (x_85 & x_86) ;
	assign x_1971 = (x_83 & x_84) ;
	assign x_1970 = (x_81 & x_82) ;
	assign x_1967 = (x_79 & x_80) ;
	assign x_1966 = (x_77 & x_78) ;
	assign x_1964 = (x_75 & x_76) ;
	assign x_74 = (v_849 | ~v_68) ;
	assign x_1960 = (x_72 & x_73) ;
	assign x_1959 = (x_70 & x_71) ;
	assign x_1957 = (x_68 & x_69) ;
	assign x_67 = (v_849 | ~v_562) ;
	assign x_1954 = (x_65 & x_66) ;
	assign x_1953 = (x_63 & x_64) ;
	assign x_1951 = (x_61 & x_62) ;
	assign x_60 = (v_854 | ~v_24) ;
	assign x_1945 = (x_58 & x_59) ;
	assign x_1944 = (x_56 & x_57) ;
	assign x_1942 = (x_54 & x_55) ;
	assign x_1941 = (x_52 & x_53) ;
	assign x_1938 = (x_50 & x_51) ;
	assign x_1937 = (x_48 & x_49) ;
	assign x_1935 = (x_46 & x_47) ;
	assign x_45 = ((~v_42 | v_74) | v_855) ;
	assign x_1931 = (x_43 & x_44) ;
	assign x_1930 = (x_41 & x_42) ;
	assign x_1928 = (x_39 & x_40) ;
	assign x_1927 = (x_37 & x_38) ;
	assign x_1924 = (x_35 & x_36) ;
	assign x_1923 = (x_33 & x_34) ;
	assign x_1921 = (x_31 & x_32) ;
	assign x_30 = (v_859 | ~v_855) ;
	assign x_1916 = (x_28 & x_29) ;
	assign x_1915 = (x_26 & x_27) ;
	assign x_1913 = (x_24 & x_25) ;
	assign x_1912 = (x_22 & x_23) ;
	assign x_1909 = (x_20 & x_21) ;
	assign x_1908 = (x_18 & x_19) ;
	assign x_1906 = (x_16 & x_17) ;
	assign x_15 = (v_865 | ~v_828) ;
	assign x_1902 = (x_13 & x_14) ;
	assign x_1901 = (x_11 & x_12) ;
	assign x_1899 = (x_9 & x_10) ;
	assign x_8 = (v_865 | ~v_710) ;
	assign x_1896 = (x_6 & x_7) ;
	assign x_1895 = (x_4 & x_5) ;
	assign x_1893 = (x_2 & x_3) ;
	assign x_1 = ((((~v_865 | ~v_556) | ~v_555) | ~v_547) | ~v_529) ;
	assign x_3774 = (x_3772 & x_3773) ;
	assign x_3771 = (x_3769 & x_3770) ;
	assign x_3767 = (x_3765 & x_3766) ;
	assign x_3764 = (x_1878 & x_3763) ;
	assign x_3760 = (x_3758 & x_3759) ;
	assign x_3757 = (x_3755 & x_3756) ;
	assign x_3753 = (x_3751 & x_3752) ;
	assign x_3750 = (x_1863 & x_3749) ;
	assign x_3745 = (x_3743 & x_3744) ;
	assign x_3742 = (x_3740 & x_3741) ;
	assign x_3738 = (x_3736 & x_3737) ;
	assign x_3735 = (x_1848 & x_3734) ;
	assign x_3731 = (x_3729 & x_3730) ;
	assign x_3728 = (x_3726 & x_3727) ;
	assign x_3724 = (x_3722 & x_3723) ;
	assign x_3721 = (x_1833 & x_3720) ;
	assign x_3715 = (x_3713 & x_3714) ;
	assign x_3712 = (x_3710 & x_3711) ;
	assign x_3708 = (x_3706 & x_3707) ;
	assign x_3705 = (x_1818 & x_3704) ;
	assign x_3701 = (x_3699 & x_3700) ;
	assign x_3698 = (x_3696 & x_3697) ;
	assign x_3694 = (x_3692 & x_3693) ;
	assign x_3691 = (x_1803 & x_3690) ;
	assign x_3686 = (x_3684 & x_3685) ;
	assign x_3683 = (x_3681 & x_3682) ;
	assign x_3679 = (x_3677 & x_3678) ;
	assign x_3676 = (x_1788 & x_3675) ;
	assign x_3672 = (x_3670 & x_3671) ;
	assign x_3669 = (x_1781 & x_3668) ;
	assign x_3666 = (x_3664 & x_3665) ;
	assign x_3663 = (x_1774 & x_3662) ;
	assign x_3656 = (x_3654 & x_3655) ;
	assign x_3653 = (x_3651 & x_3652) ;
	assign x_3649 = (x_3647 & x_3648) ;
	assign x_3646 = (x_1759 & x_3645) ;
	assign x_3642 = (x_3640 & x_3641) ;
	assign x_3639 = (x_3637 & x_3638) ;
	assign x_3635 = (x_3633 & x_3634) ;
	assign x_3632 = (x_1744 & x_3631) ;
	assign x_3627 = (x_3625 & x_3626) ;
	assign x_3624 = (x_3622 & x_3623) ;
	assign x_3620 = (x_3618 & x_3619) ;
	assign x_3617 = (x_1729 & x_3616) ;
	assign x_3613 = (x_3611 & x_3612) ;
	assign x_3610 = (x_1722 & x_3609) ;
	assign x_3607 = (x_3605 & x_3606) ;
	assign x_3604 = (x_1715 & x_3603) ;
	assign x_3598 = (x_3596 & x_3597) ;
	assign x_3595 = (x_3593 & x_3594) ;
	assign x_3591 = (x_3589 & x_3590) ;
	assign x_3588 = (x_1700 & x_3587) ;
	assign x_3584 = (x_3582 & x_3583) ;
	assign x_3581 = (x_3579 & x_3580) ;
	assign x_3577 = (x_3575 & x_3576) ;
	assign x_3574 = (x_1685 & x_3573) ;
	assign x_3569 = (x_3567 & x_3568) ;
	assign x_3566 = (x_3564 & x_3565) ;
	assign x_3562 = (x_3560 & x_3561) ;
	assign x_3559 = (x_1670 & x_3558) ;
	assign x_3555 = (x_3553 & x_3554) ;
	assign x_3552 = (x_1663 & x_3551) ;
	assign x_3549 = (x_3547 & x_3548) ;
	assign x_3546 = (x_1656 & x_3545) ;
	assign x_3538 = (x_3536 & x_3537) ;
	assign x_3535 = (x_3533 & x_3534) ;
	assign x_3531 = (x_3529 & x_3530) ;
	assign x_3528 = (x_1641 & x_3527) ;
	assign x_3524 = (x_3522 & x_3523) ;
	assign x_3521 = (x_3519 & x_3520) ;
	assign x_3517 = (x_3515 & x_3516) ;
	assign x_3514 = (x_1626 & x_3513) ;
	assign x_3509 = (x_3507 & x_3508) ;
	assign x_3506 = (x_3504 & x_3505) ;
	assign x_3502 = (x_3500 & x_3501) ;
	assign x_3499 = (x_1611 & x_3498) ;
	assign x_3495 = (x_3493 & x_3494) ;
	assign x_3492 = (x_1604 & x_3491) ;
	assign x_3489 = (x_3487 & x_3488) ;
	assign x_3486 = (x_1597 & x_3485) ;
	assign x_3480 = (x_3478 & x_3479) ;
	assign x_3477 = (x_3475 & x_3476) ;
	assign x_3473 = (x_3471 & x_3472) ;
	assign x_3470 = (x_1582 & x_3469) ;
	assign x_3466 = (x_3464 & x_3465) ;
	assign x_3463 = (x_3461 & x_3462) ;
	assign x_3459 = (x_3457 & x_3458) ;
	assign x_3456 = (x_1567 & x_3455) ;
	assign x_3451 = (x_3449 & x_3450) ;
	assign x_3448 = (x_3446 & x_3447) ;
	assign x_3444 = (x_3442 & x_3443) ;
	assign x_3441 = (x_1552 & x_3440) ;
	assign x_3437 = (x_3435 & x_3436) ;
	assign x_3434 = (x_1545 & x_3433) ;
	assign x_3431 = (x_3429 & x_3430) ;
	assign x_3428 = (x_1538 & x_3427) ;
	assign x_3421 = (x_3419 & x_3420) ;
	assign x_3418 = (x_3416 & x_3417) ;
	assign x_3414 = (x_3412 & x_3413) ;
	assign x_3411 = (x_1523 & x_3410) ;
	assign x_3407 = (x_3405 & x_3406) ;
	assign x_3404 = (x_3402 & x_3403) ;
	assign x_3400 = (x_3398 & x_3399) ;
	assign x_3397 = (x_1508 & x_3396) ;
	assign x_3392 = (x_3390 & x_3391) ;
	assign x_3389 = (x_3387 & x_3388) ;
	assign x_3385 = (x_3383 & x_3384) ;
	assign x_3382 = (x_1493 & x_3381) ;
	assign x_3378 = (x_3376 & x_3377) ;
	assign x_3375 = (x_1486 & x_3374) ;
	assign x_3372 = (x_3370 & x_3371) ;
	assign x_3369 = (x_1479 & x_3368) ;
	assign x_3363 = (x_3361 & x_3362) ;
	assign x_3360 = (x_3358 & x_3359) ;
	assign x_3356 = (x_3354 & x_3355) ;
	assign x_3353 = (x_1464 & x_3352) ;
	assign x_3349 = (x_3347 & x_3348) ;
	assign x_3346 = (x_3344 & x_3345) ;
	assign x_3342 = (x_3340 & x_3341) ;
	assign x_3339 = (x_1449 & x_3338) ;
	assign x_3334 = (x_3332 & x_3333) ;
	assign x_3331 = (x_3329 & x_3330) ;
	assign x_3327 = (x_3325 & x_3326) ;
	assign x_3324 = (x_1434 & x_3323) ;
	assign x_3320 = (x_3318 & x_3319) ;
	assign x_3317 = (x_1427 & x_3316) ;
	assign x_3314 = (x_3312 & x_3313) ;
	assign x_3311 = (x_1420 & x_3310) ;
	assign x_3302 = (x_3300 & x_3301) ;
	assign x_3299 = (x_3297 & x_3298) ;
	assign x_3295 = (x_3293 & x_3294) ;
	assign x_3292 = (x_1405 & x_3291) ;
	assign x_3288 = (x_3286 & x_3287) ;
	assign x_3285 = (x_3283 & x_3284) ;
	assign x_3281 = (x_3279 & x_3280) ;
	assign x_3278 = (x_1390 & x_3277) ;
	assign x_3273 = (x_3271 & x_3272) ;
	assign x_3270 = (x_3268 & x_3269) ;
	assign x_3266 = (x_3264 & x_3265) ;
	assign x_3263 = (x_1375 & x_3262) ;
	assign x_3259 = (x_3257 & x_3258) ;
	assign x_3256 = (x_3254 & x_3255) ;
	assign x_3252 = (x_3250 & x_3251) ;
	assign x_3249 = (x_1360 & x_3248) ;
	assign x_3243 = (x_3241 & x_3242) ;
	assign x_3240 = (x_3238 & x_3239) ;
	assign x_3236 = (x_3234 & x_3235) ;
	assign x_3233 = (x_1345 & x_3232) ;
	assign x_3229 = (x_3227 & x_3228) ;
	assign x_3226 = (x_3224 & x_3225) ;
	assign x_3222 = (x_3220 & x_3221) ;
	assign x_3219 = (x_1330 & x_3218) ;
	assign x_3214 = (x_3212 & x_3213) ;
	assign x_3211 = (x_3209 & x_3210) ;
	assign x_3207 = (x_3205 & x_3206) ;
	assign x_3204 = (x_1315 & x_3203) ;
	assign x_3200 = (x_3198 & x_3199) ;
	assign x_3197 = (x_1308 & x_3196) ;
	assign x_3194 = (x_3192 & x_3193) ;
	assign x_3191 = (x_1301 & x_3190) ;
	assign x_3184 = (x_3182 & x_3183) ;
	assign x_3181 = (x_3179 & x_3180) ;
	assign x_3177 = (x_3175 & x_3176) ;
	assign x_3174 = (x_1286 & x_3173) ;
	assign x_3170 = (x_3168 & x_3169) ;
	assign x_3167 = (x_3165 & x_3166) ;
	assign x_3163 = (x_3161 & x_3162) ;
	assign x_3160 = (x_1271 & x_3159) ;
	assign x_3155 = (x_3153 & x_3154) ;
	assign x_3152 = (x_3150 & x_3151) ;
	assign x_3148 = (x_3146 & x_3147) ;
	assign x_3145 = (x_1256 & x_3144) ;
	assign x_3141 = (x_3139 & x_3140) ;
	assign x_3138 = (x_1249 & x_3137) ;
	assign x_3135 = (x_3133 & x_3134) ;
	assign x_3132 = (x_1242 & x_3131) ;
	assign x_3126 = (x_3124 & x_3125) ;
	assign x_3123 = (x_3121 & x_3122) ;
	assign x_3119 = (x_3117 & x_3118) ;
	assign x_3116 = (x_1227 & x_3115) ;
	assign x_3112 = (x_3110 & x_3111) ;
	assign x_3109 = (x_3107 & x_3108) ;
	assign x_3105 = (x_3103 & x_3104) ;
	assign x_3102 = (x_1212 & x_3101) ;
	assign x_3097 = (x_3095 & x_3096) ;
	assign x_3094 = (x_3092 & x_3093) ;
	assign x_3090 = (x_3088 & x_3089) ;
	assign x_3087 = (x_1197 & x_3086) ;
	assign x_3083 = (x_3081 & x_3082) ;
	assign x_3080 = (x_1190 & x_3079) ;
	assign x_3077 = (x_3075 & x_3076) ;
	assign x_3074 = (x_1183 & x_3073) ;
	assign x_3066 = (x_3064 & x_3065) ;
	assign x_3063 = (x_3061 & x_3062) ;
	assign x_3059 = (x_3057 & x_3058) ;
	assign x_3056 = (x_1168 & x_3055) ;
	assign x_3052 = (x_3050 & x_3051) ;
	assign x_3049 = (x_3047 & x_3048) ;
	assign x_3045 = (x_3043 & x_3044) ;
	assign x_3042 = (x_1153 & x_3041) ;
	assign x_3037 = (x_3035 & x_3036) ;
	assign x_3034 = (x_3032 & x_3033) ;
	assign x_3030 = (x_3028 & x_3029) ;
	assign x_3027 = (x_1138 & x_3026) ;
	assign x_3023 = (x_3021 & x_3022) ;
	assign x_3020 = (x_1131 & x_3019) ;
	assign x_3017 = (x_3015 & x_3016) ;
	assign x_3014 = (x_1124 & x_3013) ;
	assign x_3008 = (x_3006 & x_3007) ;
	assign x_3005 = (x_3003 & x_3004) ;
	assign x_3001 = (x_2999 & x_3000) ;
	assign x_2998 = (x_1109 & x_2997) ;
	assign x_2994 = (x_2992 & x_2993) ;
	assign x_2991 = (x_2989 & x_2990) ;
	assign x_2987 = (x_2985 & x_2986) ;
	assign x_2984 = (x_1094 & x_2983) ;
	assign x_2979 = (x_2977 & x_2978) ;
	assign x_2976 = (x_2974 & x_2975) ;
	assign x_2972 = (x_2970 & x_2971) ;
	assign x_2969 = (x_1079 & x_2968) ;
	assign x_2965 = (x_2963 & x_2964) ;
	assign x_2962 = (x_1072 & x_2961) ;
	assign x_2959 = (x_2957 & x_2958) ;
	assign x_2956 = (x_1065 & x_2955) ;
	assign x_2949 = (x_2947 & x_2948) ;
	assign x_2946 = (x_2944 & x_2945) ;
	assign x_2942 = (x_2940 & x_2941) ;
	assign x_2939 = (x_1050 & x_2938) ;
	assign x_2935 = (x_2933 & x_2934) ;
	assign x_2932 = (x_2930 & x_2931) ;
	assign x_2928 = (x_2926 & x_2927) ;
	assign x_2925 = (x_1035 & x_2924) ;
	assign x_2920 = (x_2918 & x_2919) ;
	assign x_2917 = (x_2915 & x_2916) ;
	assign x_2913 = (x_2911 & x_2912) ;
	assign x_2910 = (x_1020 & x_2909) ;
	assign x_2906 = (x_2904 & x_2905) ;
	assign x_2903 = (x_1013 & x_2902) ;
	assign x_2900 = (x_2898 & x_2899) ;
	assign x_2897 = (x_1006 & x_2896) ;
	assign x_2891 = (x_2889 & x_2890) ;
	assign x_2888 = (x_2886 & x_2887) ;
	assign x_2884 = (x_2882 & x_2883) ;
	assign x_2881 = (x_991 & x_2880) ;
	assign x_2877 = (x_2875 & x_2876) ;
	assign x_2874 = (x_2872 & x_2873) ;
	assign x_2870 = (x_2868 & x_2869) ;
	assign x_2867 = (x_976 & x_2866) ;
	assign x_2862 = (x_2860 & x_2861) ;
	assign x_2859 = (x_2857 & x_2858) ;
	assign x_2855 = (x_2853 & x_2854) ;
	assign x_2852 = (x_961 & x_2851) ;
	assign x_2848 = (x_2846 & x_2847) ;
	assign x_2845 = (x_954 & x_2844) ;
	assign x_2842 = (x_2840 & x_2841) ;
	assign x_2839 = (x_947 & x_2838) ;
	assign x_2829 = (x_2827 & x_2828) ;
	assign x_2826 = (x_2824 & x_2825) ;
	assign x_2822 = (x_2820 & x_2821) ;
	assign x_2819 = (x_932 & x_2818) ;
	assign x_2815 = (x_2813 & x_2814) ;
	assign x_2812 = (x_2810 & x_2811) ;
	assign x_2808 = (x_2806 & x_2807) ;
	assign x_2805 = (x_917 & x_2804) ;
	assign x_2800 = (x_2798 & x_2799) ;
	assign x_2797 = (x_2795 & x_2796) ;
	assign x_2793 = (x_2791 & x_2792) ;
	assign x_2790 = (x_902 & x_2789) ;
	assign x_2786 = (x_2784 & x_2785) ;
	assign x_2783 = (x_2781 & x_2782) ;
	assign x_2779 = (x_2777 & x_2778) ;
	assign x_2776 = (x_887 & x_2775) ;
	assign x_2770 = (x_2768 & x_2769) ;
	assign x_2767 = (x_2765 & x_2766) ;
	assign x_2763 = (x_2761 & x_2762) ;
	assign x_2760 = (x_872 & x_2759) ;
	assign x_2756 = (x_2754 & x_2755) ;
	assign x_2753 = (x_2751 & x_2752) ;
	assign x_2749 = (x_2747 & x_2748) ;
	assign x_2746 = (x_857 & x_2745) ;
	assign x_2741 = (x_2739 & x_2740) ;
	assign x_2738 = (x_2736 & x_2737) ;
	assign x_2734 = (x_2732 & x_2733) ;
	assign x_2731 = (x_842 & x_2730) ;
	assign x_2727 = (x_2725 & x_2726) ;
	assign x_2724 = (x_835 & x_2723) ;
	assign x_2721 = (x_2719 & x_2720) ;
	assign x_2718 = (x_828 & x_2717) ;
	assign x_2711 = (x_2709 & x_2710) ;
	assign x_2708 = (x_2706 & x_2707) ;
	assign x_2704 = (x_2702 & x_2703) ;
	assign x_2701 = (x_813 & x_2700) ;
	assign x_2697 = (x_2695 & x_2696) ;
	assign x_2694 = (x_2692 & x_2693) ;
	assign x_2690 = (x_2688 & x_2689) ;
	assign x_2687 = (x_798 & x_2686) ;
	assign x_2682 = (x_2680 & x_2681) ;
	assign x_2679 = (x_2677 & x_2678) ;
	assign x_2675 = (x_2673 & x_2674) ;
	assign x_2672 = (x_783 & x_2671) ;
	assign x_2668 = (x_2666 & x_2667) ;
	assign x_2665 = (x_776 & x_2664) ;
	assign x_2662 = (x_2660 & x_2661) ;
	assign x_2659 = (x_769 & x_2658) ;
	assign x_2653 = (x_2651 & x_2652) ;
	assign x_2650 = (x_2648 & x_2649) ;
	assign x_2646 = (x_2644 & x_2645) ;
	assign x_2643 = (x_754 & x_2642) ;
	assign x_2639 = (x_2637 & x_2638) ;
	assign x_2636 = (x_2634 & x_2635) ;
	assign x_2632 = (x_2630 & x_2631) ;
	assign x_2629 = (x_739 & x_2628) ;
	assign x_2624 = (x_2622 & x_2623) ;
	assign x_2621 = (x_2619 & x_2620) ;
	assign x_2617 = (x_2615 & x_2616) ;
	assign x_2614 = (x_724 & x_2613) ;
	assign x_2610 = (x_2608 & x_2609) ;
	assign x_2607 = (x_717 & x_2606) ;
	assign x_2604 = (x_2602 & x_2603) ;
	assign x_2601 = (x_710 & x_2600) ;
	assign x_2593 = (x_2591 & x_2592) ;
	assign x_2590 = (x_2588 & x_2589) ;
	assign x_2586 = (x_2584 & x_2585) ;
	assign x_2583 = (x_695 & x_2582) ;
	assign x_2579 = (x_2577 & x_2578) ;
	assign x_2576 = (x_2574 & x_2575) ;
	assign x_2572 = (x_2570 & x_2571) ;
	assign x_2569 = (x_680 & x_2568) ;
	assign x_2564 = (x_2562 & x_2563) ;
	assign x_2561 = (x_2559 & x_2560) ;
	assign x_2557 = (x_2555 & x_2556) ;
	assign x_2554 = (x_665 & x_2553) ;
	assign x_2550 = (x_2548 & x_2549) ;
	assign x_2547 = (x_658 & x_2546) ;
	assign x_2544 = (x_2542 & x_2543) ;
	assign x_2541 = (x_651 & x_2540) ;
	assign x_2535 = (x_2533 & x_2534) ;
	assign x_2532 = (x_2530 & x_2531) ;
	assign x_2528 = (x_2526 & x_2527) ;
	assign x_2525 = (x_636 & x_2524) ;
	assign x_2521 = (x_2519 & x_2520) ;
	assign x_2518 = (x_2516 & x_2517) ;
	assign x_2514 = (x_2512 & x_2513) ;
	assign x_2511 = (x_621 & x_2510) ;
	assign x_2506 = (x_2504 & x_2505) ;
	assign x_2503 = (x_2501 & x_2502) ;
	assign x_2499 = (x_2497 & x_2498) ;
	assign x_2496 = (x_606 & x_2495) ;
	assign x_2492 = (x_2490 & x_2491) ;
	assign x_2489 = (x_599 & x_2488) ;
	assign x_2486 = (x_2484 & x_2485) ;
	assign x_2483 = (x_592 & x_2482) ;
	assign x_2476 = (x_2474 & x_2475) ;
	assign x_2473 = (x_2471 & x_2472) ;
	assign x_2469 = (x_2467 & x_2468) ;
	assign x_2466 = (x_577 & x_2465) ;
	assign x_2462 = (x_2460 & x_2461) ;
	assign x_2459 = (x_2457 & x_2458) ;
	assign x_2455 = (x_2453 & x_2454) ;
	assign x_2452 = (x_562 & x_2451) ;
	assign x_2447 = (x_2445 & x_2446) ;
	assign x_2444 = (x_2442 & x_2443) ;
	assign x_2440 = (x_2438 & x_2439) ;
	assign x_2437 = (x_547 & x_2436) ;
	assign x_2433 = (x_2431 & x_2432) ;
	assign x_2430 = (x_540 & x_2429) ;
	assign x_2427 = (x_2425 & x_2426) ;
	assign x_2424 = (x_533 & x_2423) ;
	assign x_2418 = (x_2416 & x_2417) ;
	assign x_2415 = (x_2413 & x_2414) ;
	assign x_2411 = (x_2409 & x_2410) ;
	assign x_2408 = (x_518 & x_2407) ;
	assign x_2404 = (x_2402 & x_2403) ;
	assign x_2401 = (x_2399 & x_2400) ;
	assign x_2397 = (x_2395 & x_2396) ;
	assign x_2394 = (x_503 & x_2393) ;
	assign x_2389 = (x_2387 & x_2388) ;
	assign x_2386 = (x_2384 & x_2385) ;
	assign x_2382 = (x_2380 & x_2381) ;
	assign x_2379 = (x_488 & x_2378) ;
	assign x_2375 = (x_2373 & x_2374) ;
	assign x_2372 = (x_481 & x_2371) ;
	assign x_2369 = (x_2367 & x_2368) ;
	assign x_2366 = (x_474 & x_2365) ;
	assign x_2357 = (x_2355 & x_2356) ;
	assign x_2354 = (x_2352 & x_2353) ;
	assign x_2350 = (x_2348 & x_2349) ;
	assign x_2347 = (x_459 & x_2346) ;
	assign x_2343 = (x_2341 & x_2342) ;
	assign x_2340 = (x_2338 & x_2339) ;
	assign x_2336 = (x_2334 & x_2335) ;
	assign x_2333 = (x_444 & x_2332) ;
	assign x_2328 = (x_2326 & x_2327) ;
	assign x_2325 = (x_2323 & x_2324) ;
	assign x_2321 = (x_2319 & x_2320) ;
	assign x_2318 = (x_429 & x_2317) ;
	assign x_2314 = (x_2312 & x_2313) ;
	assign x_2311 = (x_2309 & x_2310) ;
	assign x_2307 = (x_2305 & x_2306) ;
	assign x_2304 = (x_414 & x_2303) ;
	assign x_2298 = (x_2296 & x_2297) ;
	assign x_2295 = (x_2293 & x_2294) ;
	assign x_2291 = (x_2289 & x_2290) ;
	assign x_2288 = (x_399 & x_2287) ;
	assign x_2284 = (x_2282 & x_2283) ;
	assign x_2281 = (x_2279 & x_2280) ;
	assign x_2277 = (x_2275 & x_2276) ;
	assign x_2274 = (x_384 & x_2273) ;
	assign x_2269 = (x_2267 & x_2268) ;
	assign x_2266 = (x_2264 & x_2265) ;
	assign x_2262 = (x_2260 & x_2261) ;
	assign x_2259 = (x_369 & x_2258) ;
	assign x_2255 = (x_2253 & x_2254) ;
	assign x_2252 = (x_362 & x_2251) ;
	assign x_2249 = (x_2247 & x_2248) ;
	assign x_2246 = (x_355 & x_2245) ;
	assign x_2239 = (x_2237 & x_2238) ;
	assign x_2236 = (x_2234 & x_2235) ;
	assign x_2232 = (x_2230 & x_2231) ;
	assign x_2229 = (x_340 & x_2228) ;
	assign x_2225 = (x_2223 & x_2224) ;
	assign x_2222 = (x_2220 & x_2221) ;
	assign x_2218 = (x_2216 & x_2217) ;
	assign x_2215 = (x_325 & x_2214) ;
	assign x_2210 = (x_2208 & x_2209) ;
	assign x_2207 = (x_2205 & x_2206) ;
	assign x_2203 = (x_2201 & x_2202) ;
	assign x_2200 = (x_310 & x_2199) ;
	assign x_2196 = (x_2194 & x_2195) ;
	assign x_2193 = (x_303 & x_2192) ;
	assign x_2190 = (x_2188 & x_2189) ;
	assign x_2187 = (x_296 & x_2186) ;
	assign x_2181 = (x_2179 & x_2180) ;
	assign x_2178 = (x_2176 & x_2177) ;
	assign x_2174 = (x_2172 & x_2173) ;
	assign x_2171 = (x_281 & x_2170) ;
	assign x_2167 = (x_2165 & x_2166) ;
	assign x_2164 = (x_2162 & x_2163) ;
	assign x_2160 = (x_2158 & x_2159) ;
	assign x_2157 = (x_266 & x_2156) ;
	assign x_2152 = (x_2150 & x_2151) ;
	assign x_2149 = (x_2147 & x_2148) ;
	assign x_2145 = (x_2143 & x_2144) ;
	assign x_2142 = (x_251 & x_2141) ;
	assign x_2138 = (x_2136 & x_2137) ;
	assign x_2135 = (x_244 & x_2134) ;
	assign x_2132 = (x_2130 & x_2131) ;
	assign x_2129 = (x_237 & x_2128) ;
	assign x_2121 = (x_2119 & x_2120) ;
	assign x_2118 = (x_2116 & x_2117) ;
	assign x_2114 = (x_2112 & x_2113) ;
	assign x_2111 = (x_222 & x_2110) ;
	assign x_2107 = (x_2105 & x_2106) ;
	assign x_2104 = (x_2102 & x_2103) ;
	assign x_2100 = (x_2098 & x_2099) ;
	assign x_2097 = (x_207 & x_2096) ;
	assign x_2092 = (x_2090 & x_2091) ;
	assign x_2089 = (x_2087 & x_2088) ;
	assign x_2085 = (x_2083 & x_2084) ;
	assign x_2082 = (x_192 & x_2081) ;
	assign x_2078 = (x_2076 & x_2077) ;
	assign x_2075 = (x_185 & x_2074) ;
	assign x_2072 = (x_2070 & x_2071) ;
	assign x_2069 = (x_178 & x_2068) ;
	assign x_2063 = (x_2061 & x_2062) ;
	assign x_2060 = (x_2058 & x_2059) ;
	assign x_2056 = (x_2054 & x_2055) ;
	assign x_2053 = (x_163 & x_2052) ;
	assign x_2049 = (x_2047 & x_2048) ;
	assign x_2046 = (x_2044 & x_2045) ;
	assign x_2042 = (x_2040 & x_2041) ;
	assign x_2039 = (x_148 & x_2038) ;
	assign x_2034 = (x_2032 & x_2033) ;
	assign x_2031 = (x_2029 & x_2030) ;
	assign x_2027 = (x_2025 & x_2026) ;
	assign x_2024 = (x_133 & x_2023) ;
	assign x_2020 = (x_2018 & x_2019) ;
	assign x_2017 = (x_126 & x_2016) ;
	assign x_2014 = (x_2012 & x_2013) ;
	assign x_2011 = (x_119 & x_2010) ;
	assign x_2004 = (x_2002 & x_2003) ;
	assign x_2001 = (x_1999 & x_2000) ;
	assign x_1997 = (x_1995 & x_1996) ;
	assign x_1994 = (x_104 & x_1993) ;
	assign x_1990 = (x_1988 & x_1989) ;
	assign x_1987 = (x_1985 & x_1986) ;
	assign x_1983 = (x_1981 & x_1982) ;
	assign x_1980 = (x_89 & x_1979) ;
	assign x_1975 = (x_1973 & x_1974) ;
	assign x_1972 = (x_1970 & x_1971) ;
	assign x_1968 = (x_1966 & x_1967) ;
	assign x_1965 = (x_74 & x_1964) ;
	assign x_1961 = (x_1959 & x_1960) ;
	assign x_1958 = (x_67 & x_1957) ;
	assign x_1955 = (x_1953 & x_1954) ;
	assign x_1952 = (x_60 & x_1951) ;
	assign x_1946 = (x_1944 & x_1945) ;
	assign x_1943 = (x_1941 & x_1942) ;
	assign x_1939 = (x_1937 & x_1938) ;
	assign x_1936 = (x_45 & x_1935) ;
	assign x_1932 = (x_1930 & x_1931) ;
	assign x_1929 = (x_1927 & x_1928) ;
	assign x_1925 = (x_1923 & x_1924) ;
	assign x_1922 = (x_30 & x_1921) ;
	assign x_1917 = (x_1915 & x_1916) ;
	assign x_1914 = (x_1912 & x_1913) ;
	assign x_1910 = (x_1908 & x_1909) ;
	assign x_1907 = (x_15 & x_1906) ;
	assign x_1903 = (x_1901 & x_1902) ;
	assign x_1900 = (x_8 & x_1899) ;
	assign x_1897 = (x_1895 & x_1896) ;
	assign x_1894 = (x_1 & x_1893) ;
	assign x_3775 = (x_3771 & x_3774) ;
	assign x_3768 = (x_3764 & x_3767) ;
	assign x_3761 = (x_3757 & x_3760) ;
	assign x_3754 = (x_3750 & x_3753) ;
	assign x_3746 = (x_3742 & x_3745) ;
	assign x_3739 = (x_3735 & x_3738) ;
	assign x_3732 = (x_3728 & x_3731) ;
	assign x_3725 = (x_3721 & x_3724) ;
	assign x_3716 = (x_3712 & x_3715) ;
	assign x_3709 = (x_3705 & x_3708) ;
	assign x_3702 = (x_3698 & x_3701) ;
	assign x_3695 = (x_3691 & x_3694) ;
	assign x_3687 = (x_3683 & x_3686) ;
	assign x_3680 = (x_3676 & x_3679) ;
	assign x_3673 = (x_3669 & x_3672) ;
	assign x_3667 = (x_3663 & x_3666) ;
	assign x_3657 = (x_3653 & x_3656) ;
	assign x_3650 = (x_3646 & x_3649) ;
	assign x_3643 = (x_3639 & x_3642) ;
	assign x_3636 = (x_3632 & x_3635) ;
	assign x_3628 = (x_3624 & x_3627) ;
	assign x_3621 = (x_3617 & x_3620) ;
	assign x_3614 = (x_3610 & x_3613) ;
	assign x_3608 = (x_3604 & x_3607) ;
	assign x_3599 = (x_3595 & x_3598) ;
	assign x_3592 = (x_3588 & x_3591) ;
	assign x_3585 = (x_3581 & x_3584) ;
	assign x_3578 = (x_3574 & x_3577) ;
	assign x_3570 = (x_3566 & x_3569) ;
	assign x_3563 = (x_3559 & x_3562) ;
	assign x_3556 = (x_3552 & x_3555) ;
	assign x_3550 = (x_3546 & x_3549) ;
	assign x_3539 = (x_3535 & x_3538) ;
	assign x_3532 = (x_3528 & x_3531) ;
	assign x_3525 = (x_3521 & x_3524) ;
	assign x_3518 = (x_3514 & x_3517) ;
	assign x_3510 = (x_3506 & x_3509) ;
	assign x_3503 = (x_3499 & x_3502) ;
	assign x_3496 = (x_3492 & x_3495) ;
	assign x_3490 = (x_3486 & x_3489) ;
	assign x_3481 = (x_3477 & x_3480) ;
	assign x_3474 = (x_3470 & x_3473) ;
	assign x_3467 = (x_3463 & x_3466) ;
	assign x_3460 = (x_3456 & x_3459) ;
	assign x_3452 = (x_3448 & x_3451) ;
	assign x_3445 = (x_3441 & x_3444) ;
	assign x_3438 = (x_3434 & x_3437) ;
	assign x_3432 = (x_3428 & x_3431) ;
	assign x_3422 = (x_3418 & x_3421) ;
	assign x_3415 = (x_3411 & x_3414) ;
	assign x_3408 = (x_3404 & x_3407) ;
	assign x_3401 = (x_3397 & x_3400) ;
	assign x_3393 = (x_3389 & x_3392) ;
	assign x_3386 = (x_3382 & x_3385) ;
	assign x_3379 = (x_3375 & x_3378) ;
	assign x_3373 = (x_3369 & x_3372) ;
	assign x_3364 = (x_3360 & x_3363) ;
	assign x_3357 = (x_3353 & x_3356) ;
	assign x_3350 = (x_3346 & x_3349) ;
	assign x_3343 = (x_3339 & x_3342) ;
	assign x_3335 = (x_3331 & x_3334) ;
	assign x_3328 = (x_3324 & x_3327) ;
	assign x_3321 = (x_3317 & x_3320) ;
	assign x_3315 = (x_3311 & x_3314) ;
	assign x_3303 = (x_3299 & x_3302) ;
	assign x_3296 = (x_3292 & x_3295) ;
	assign x_3289 = (x_3285 & x_3288) ;
	assign x_3282 = (x_3278 & x_3281) ;
	assign x_3274 = (x_3270 & x_3273) ;
	assign x_3267 = (x_3263 & x_3266) ;
	assign x_3260 = (x_3256 & x_3259) ;
	assign x_3253 = (x_3249 & x_3252) ;
	assign x_3244 = (x_3240 & x_3243) ;
	assign x_3237 = (x_3233 & x_3236) ;
	assign x_3230 = (x_3226 & x_3229) ;
	assign x_3223 = (x_3219 & x_3222) ;
	assign x_3215 = (x_3211 & x_3214) ;
	assign x_3208 = (x_3204 & x_3207) ;
	assign x_3201 = (x_3197 & x_3200) ;
	assign x_3195 = (x_3191 & x_3194) ;
	assign x_3185 = (x_3181 & x_3184) ;
	assign x_3178 = (x_3174 & x_3177) ;
	assign x_3171 = (x_3167 & x_3170) ;
	assign x_3164 = (x_3160 & x_3163) ;
	assign x_3156 = (x_3152 & x_3155) ;
	assign x_3149 = (x_3145 & x_3148) ;
	assign x_3142 = (x_3138 & x_3141) ;
	assign x_3136 = (x_3132 & x_3135) ;
	assign x_3127 = (x_3123 & x_3126) ;
	assign x_3120 = (x_3116 & x_3119) ;
	assign x_3113 = (x_3109 & x_3112) ;
	assign x_3106 = (x_3102 & x_3105) ;
	assign x_3098 = (x_3094 & x_3097) ;
	assign x_3091 = (x_3087 & x_3090) ;
	assign x_3084 = (x_3080 & x_3083) ;
	assign x_3078 = (x_3074 & x_3077) ;
	assign x_3067 = (x_3063 & x_3066) ;
	assign x_3060 = (x_3056 & x_3059) ;
	assign x_3053 = (x_3049 & x_3052) ;
	assign x_3046 = (x_3042 & x_3045) ;
	assign x_3038 = (x_3034 & x_3037) ;
	assign x_3031 = (x_3027 & x_3030) ;
	assign x_3024 = (x_3020 & x_3023) ;
	assign x_3018 = (x_3014 & x_3017) ;
	assign x_3009 = (x_3005 & x_3008) ;
	assign x_3002 = (x_2998 & x_3001) ;
	assign x_2995 = (x_2991 & x_2994) ;
	assign x_2988 = (x_2984 & x_2987) ;
	assign x_2980 = (x_2976 & x_2979) ;
	assign x_2973 = (x_2969 & x_2972) ;
	assign x_2966 = (x_2962 & x_2965) ;
	assign x_2960 = (x_2956 & x_2959) ;
	assign x_2950 = (x_2946 & x_2949) ;
	assign x_2943 = (x_2939 & x_2942) ;
	assign x_2936 = (x_2932 & x_2935) ;
	assign x_2929 = (x_2925 & x_2928) ;
	assign x_2921 = (x_2917 & x_2920) ;
	assign x_2914 = (x_2910 & x_2913) ;
	assign x_2907 = (x_2903 & x_2906) ;
	assign x_2901 = (x_2897 & x_2900) ;
	assign x_2892 = (x_2888 & x_2891) ;
	assign x_2885 = (x_2881 & x_2884) ;
	assign x_2878 = (x_2874 & x_2877) ;
	assign x_2871 = (x_2867 & x_2870) ;
	assign x_2863 = (x_2859 & x_2862) ;
	assign x_2856 = (x_2852 & x_2855) ;
	assign x_2849 = (x_2845 & x_2848) ;
	assign x_2843 = (x_2839 & x_2842) ;
	assign x_2830 = (x_2826 & x_2829) ;
	assign x_2823 = (x_2819 & x_2822) ;
	assign x_2816 = (x_2812 & x_2815) ;
	assign x_2809 = (x_2805 & x_2808) ;
	assign x_2801 = (x_2797 & x_2800) ;
	assign x_2794 = (x_2790 & x_2793) ;
	assign x_2787 = (x_2783 & x_2786) ;
	assign x_2780 = (x_2776 & x_2779) ;
	assign x_2771 = (x_2767 & x_2770) ;
	assign x_2764 = (x_2760 & x_2763) ;
	assign x_2757 = (x_2753 & x_2756) ;
	assign x_2750 = (x_2746 & x_2749) ;
	assign x_2742 = (x_2738 & x_2741) ;
	assign x_2735 = (x_2731 & x_2734) ;
	assign x_2728 = (x_2724 & x_2727) ;
	assign x_2722 = (x_2718 & x_2721) ;
	assign x_2712 = (x_2708 & x_2711) ;
	assign x_2705 = (x_2701 & x_2704) ;
	assign x_2698 = (x_2694 & x_2697) ;
	assign x_2691 = (x_2687 & x_2690) ;
	assign x_2683 = (x_2679 & x_2682) ;
	assign x_2676 = (x_2672 & x_2675) ;
	assign x_2669 = (x_2665 & x_2668) ;
	assign x_2663 = (x_2659 & x_2662) ;
	assign x_2654 = (x_2650 & x_2653) ;
	assign x_2647 = (x_2643 & x_2646) ;
	assign x_2640 = (x_2636 & x_2639) ;
	assign x_2633 = (x_2629 & x_2632) ;
	assign x_2625 = (x_2621 & x_2624) ;
	assign x_2618 = (x_2614 & x_2617) ;
	assign x_2611 = (x_2607 & x_2610) ;
	assign x_2605 = (x_2601 & x_2604) ;
	assign x_2594 = (x_2590 & x_2593) ;
	assign x_2587 = (x_2583 & x_2586) ;
	assign x_2580 = (x_2576 & x_2579) ;
	assign x_2573 = (x_2569 & x_2572) ;
	assign x_2565 = (x_2561 & x_2564) ;
	assign x_2558 = (x_2554 & x_2557) ;
	assign x_2551 = (x_2547 & x_2550) ;
	assign x_2545 = (x_2541 & x_2544) ;
	assign x_2536 = (x_2532 & x_2535) ;
	assign x_2529 = (x_2525 & x_2528) ;
	assign x_2522 = (x_2518 & x_2521) ;
	assign x_2515 = (x_2511 & x_2514) ;
	assign x_2507 = (x_2503 & x_2506) ;
	assign x_2500 = (x_2496 & x_2499) ;
	assign x_2493 = (x_2489 & x_2492) ;
	assign x_2487 = (x_2483 & x_2486) ;
	assign x_2477 = (x_2473 & x_2476) ;
	assign x_2470 = (x_2466 & x_2469) ;
	assign x_2463 = (x_2459 & x_2462) ;
	assign x_2456 = (x_2452 & x_2455) ;
	assign x_2448 = (x_2444 & x_2447) ;
	assign x_2441 = (x_2437 & x_2440) ;
	assign x_2434 = (x_2430 & x_2433) ;
	assign x_2428 = (x_2424 & x_2427) ;
	assign x_2419 = (x_2415 & x_2418) ;
	assign x_2412 = (x_2408 & x_2411) ;
	assign x_2405 = (x_2401 & x_2404) ;
	assign x_2398 = (x_2394 & x_2397) ;
	assign x_2390 = (x_2386 & x_2389) ;
	assign x_2383 = (x_2379 & x_2382) ;
	assign x_2376 = (x_2372 & x_2375) ;
	assign x_2370 = (x_2366 & x_2369) ;
	assign x_2358 = (x_2354 & x_2357) ;
	assign x_2351 = (x_2347 & x_2350) ;
	assign x_2344 = (x_2340 & x_2343) ;
	assign x_2337 = (x_2333 & x_2336) ;
	assign x_2329 = (x_2325 & x_2328) ;
	assign x_2322 = (x_2318 & x_2321) ;
	assign x_2315 = (x_2311 & x_2314) ;
	assign x_2308 = (x_2304 & x_2307) ;
	assign x_2299 = (x_2295 & x_2298) ;
	assign x_2292 = (x_2288 & x_2291) ;
	assign x_2285 = (x_2281 & x_2284) ;
	assign x_2278 = (x_2274 & x_2277) ;
	assign x_2270 = (x_2266 & x_2269) ;
	assign x_2263 = (x_2259 & x_2262) ;
	assign x_2256 = (x_2252 & x_2255) ;
	assign x_2250 = (x_2246 & x_2249) ;
	assign x_2240 = (x_2236 & x_2239) ;
	assign x_2233 = (x_2229 & x_2232) ;
	assign x_2226 = (x_2222 & x_2225) ;
	assign x_2219 = (x_2215 & x_2218) ;
	assign x_2211 = (x_2207 & x_2210) ;
	assign x_2204 = (x_2200 & x_2203) ;
	assign x_2197 = (x_2193 & x_2196) ;
	assign x_2191 = (x_2187 & x_2190) ;
	assign x_2182 = (x_2178 & x_2181) ;
	assign x_2175 = (x_2171 & x_2174) ;
	assign x_2168 = (x_2164 & x_2167) ;
	assign x_2161 = (x_2157 & x_2160) ;
	assign x_2153 = (x_2149 & x_2152) ;
	assign x_2146 = (x_2142 & x_2145) ;
	assign x_2139 = (x_2135 & x_2138) ;
	assign x_2133 = (x_2129 & x_2132) ;
	assign x_2122 = (x_2118 & x_2121) ;
	assign x_2115 = (x_2111 & x_2114) ;
	assign x_2108 = (x_2104 & x_2107) ;
	assign x_2101 = (x_2097 & x_2100) ;
	assign x_2093 = (x_2089 & x_2092) ;
	assign x_2086 = (x_2082 & x_2085) ;
	assign x_2079 = (x_2075 & x_2078) ;
	assign x_2073 = (x_2069 & x_2072) ;
	assign x_2064 = (x_2060 & x_2063) ;
	assign x_2057 = (x_2053 & x_2056) ;
	assign x_2050 = (x_2046 & x_2049) ;
	assign x_2043 = (x_2039 & x_2042) ;
	assign x_2035 = (x_2031 & x_2034) ;
	assign x_2028 = (x_2024 & x_2027) ;
	assign x_2021 = (x_2017 & x_2020) ;
	assign x_2015 = (x_2011 & x_2014) ;
	assign x_2005 = (x_2001 & x_2004) ;
	assign x_1998 = (x_1994 & x_1997) ;
	assign x_1991 = (x_1987 & x_1990) ;
	assign x_1984 = (x_1980 & x_1983) ;
	assign x_1976 = (x_1972 & x_1975) ;
	assign x_1969 = (x_1965 & x_1968) ;
	assign x_1962 = (x_1958 & x_1961) ;
	assign x_1956 = (x_1952 & x_1955) ;
	assign x_1947 = (x_1943 & x_1946) ;
	assign x_1940 = (x_1936 & x_1939) ;
	assign x_1933 = (x_1929 & x_1932) ;
	assign x_1926 = (x_1922 & x_1925) ;
	assign x_1918 = (x_1914 & x_1917) ;
	assign x_1911 = (x_1907 & x_1910) ;
	assign x_1904 = (x_1900 & x_1903) ;
	assign x_1898 = (x_1894 & x_1897) ;
	assign x_3776 = (x_3768 & x_3775) ;
	assign x_3762 = (x_3754 & x_3761) ;
	assign x_3747 = (x_3739 & x_3746) ;
	assign x_3733 = (x_3725 & x_3732) ;
	assign x_3717 = (x_3709 & x_3716) ;
	assign x_3703 = (x_3695 & x_3702) ;
	assign x_3688 = (x_3680 & x_3687) ;
	assign x_3674 = (x_3667 & x_3673) ;
	assign x_3658 = (x_3650 & x_3657) ;
	assign x_3644 = (x_3636 & x_3643) ;
	assign x_3629 = (x_3621 & x_3628) ;
	assign x_3615 = (x_3608 & x_3614) ;
	assign x_3600 = (x_3592 & x_3599) ;
	assign x_3586 = (x_3578 & x_3585) ;
	assign x_3571 = (x_3563 & x_3570) ;
	assign x_3557 = (x_3550 & x_3556) ;
	assign x_3540 = (x_3532 & x_3539) ;
	assign x_3526 = (x_3518 & x_3525) ;
	assign x_3511 = (x_3503 & x_3510) ;
	assign x_3497 = (x_3490 & x_3496) ;
	assign x_3482 = (x_3474 & x_3481) ;
	assign x_3468 = (x_3460 & x_3467) ;
	assign x_3453 = (x_3445 & x_3452) ;
	assign x_3439 = (x_3432 & x_3438) ;
	assign x_3423 = (x_3415 & x_3422) ;
	assign x_3409 = (x_3401 & x_3408) ;
	assign x_3394 = (x_3386 & x_3393) ;
	assign x_3380 = (x_3373 & x_3379) ;
	assign x_3365 = (x_3357 & x_3364) ;
	assign x_3351 = (x_3343 & x_3350) ;
	assign x_3336 = (x_3328 & x_3335) ;
	assign x_3322 = (x_3315 & x_3321) ;
	assign x_3304 = (x_3296 & x_3303) ;
	assign x_3290 = (x_3282 & x_3289) ;
	assign x_3275 = (x_3267 & x_3274) ;
	assign x_3261 = (x_3253 & x_3260) ;
	assign x_3245 = (x_3237 & x_3244) ;
	assign x_3231 = (x_3223 & x_3230) ;
	assign x_3216 = (x_3208 & x_3215) ;
	assign x_3202 = (x_3195 & x_3201) ;
	assign x_3186 = (x_3178 & x_3185) ;
	assign x_3172 = (x_3164 & x_3171) ;
	assign x_3157 = (x_3149 & x_3156) ;
	assign x_3143 = (x_3136 & x_3142) ;
	assign x_3128 = (x_3120 & x_3127) ;
	assign x_3114 = (x_3106 & x_3113) ;
	assign x_3099 = (x_3091 & x_3098) ;
	assign x_3085 = (x_3078 & x_3084) ;
	assign x_3068 = (x_3060 & x_3067) ;
	assign x_3054 = (x_3046 & x_3053) ;
	assign x_3039 = (x_3031 & x_3038) ;
	assign x_3025 = (x_3018 & x_3024) ;
	assign x_3010 = (x_3002 & x_3009) ;
	assign x_2996 = (x_2988 & x_2995) ;
	assign x_2981 = (x_2973 & x_2980) ;
	assign x_2967 = (x_2960 & x_2966) ;
	assign x_2951 = (x_2943 & x_2950) ;
	assign x_2937 = (x_2929 & x_2936) ;
	assign x_2922 = (x_2914 & x_2921) ;
	assign x_2908 = (x_2901 & x_2907) ;
	assign x_2893 = (x_2885 & x_2892) ;
	assign x_2879 = (x_2871 & x_2878) ;
	assign x_2864 = (x_2856 & x_2863) ;
	assign x_2850 = (x_2843 & x_2849) ;
	assign x_2831 = (x_2823 & x_2830) ;
	assign x_2817 = (x_2809 & x_2816) ;
	assign x_2802 = (x_2794 & x_2801) ;
	assign x_2788 = (x_2780 & x_2787) ;
	assign x_2772 = (x_2764 & x_2771) ;
	assign x_2758 = (x_2750 & x_2757) ;
	assign x_2743 = (x_2735 & x_2742) ;
	assign x_2729 = (x_2722 & x_2728) ;
	assign x_2713 = (x_2705 & x_2712) ;
	assign x_2699 = (x_2691 & x_2698) ;
	assign x_2684 = (x_2676 & x_2683) ;
	assign x_2670 = (x_2663 & x_2669) ;
	assign x_2655 = (x_2647 & x_2654) ;
	assign x_2641 = (x_2633 & x_2640) ;
	assign x_2626 = (x_2618 & x_2625) ;
	assign x_2612 = (x_2605 & x_2611) ;
	assign x_2595 = (x_2587 & x_2594) ;
	assign x_2581 = (x_2573 & x_2580) ;
	assign x_2566 = (x_2558 & x_2565) ;
	assign x_2552 = (x_2545 & x_2551) ;
	assign x_2537 = (x_2529 & x_2536) ;
	assign x_2523 = (x_2515 & x_2522) ;
	assign x_2508 = (x_2500 & x_2507) ;
	assign x_2494 = (x_2487 & x_2493) ;
	assign x_2478 = (x_2470 & x_2477) ;
	assign x_2464 = (x_2456 & x_2463) ;
	assign x_2449 = (x_2441 & x_2448) ;
	assign x_2435 = (x_2428 & x_2434) ;
	assign x_2420 = (x_2412 & x_2419) ;
	assign x_2406 = (x_2398 & x_2405) ;
	assign x_2391 = (x_2383 & x_2390) ;
	assign x_2377 = (x_2370 & x_2376) ;
	assign x_2359 = (x_2351 & x_2358) ;
	assign x_2345 = (x_2337 & x_2344) ;
	assign x_2330 = (x_2322 & x_2329) ;
	assign x_2316 = (x_2308 & x_2315) ;
	assign x_2300 = (x_2292 & x_2299) ;
	assign x_2286 = (x_2278 & x_2285) ;
	assign x_2271 = (x_2263 & x_2270) ;
	assign x_2257 = (x_2250 & x_2256) ;
	assign x_2241 = (x_2233 & x_2240) ;
	assign x_2227 = (x_2219 & x_2226) ;
	assign x_2212 = (x_2204 & x_2211) ;
	assign x_2198 = (x_2191 & x_2197) ;
	assign x_2183 = (x_2175 & x_2182) ;
	assign x_2169 = (x_2161 & x_2168) ;
	assign x_2154 = (x_2146 & x_2153) ;
	assign x_2140 = (x_2133 & x_2139) ;
	assign x_2123 = (x_2115 & x_2122) ;
	assign x_2109 = (x_2101 & x_2108) ;
	assign x_2094 = (x_2086 & x_2093) ;
	assign x_2080 = (x_2073 & x_2079) ;
	assign x_2065 = (x_2057 & x_2064) ;
	assign x_2051 = (x_2043 & x_2050) ;
	assign x_2036 = (x_2028 & x_2035) ;
	assign x_2022 = (x_2015 & x_2021) ;
	assign x_2006 = (x_1998 & x_2005) ;
	assign x_1992 = (x_1984 & x_1991) ;
	assign x_1977 = (x_1969 & x_1976) ;
	assign x_1963 = (x_1956 & x_1962) ;
	assign x_1948 = (x_1940 & x_1947) ;
	assign x_1934 = (x_1926 & x_1933) ;
	assign x_1919 = (x_1911 & x_1918) ;
	assign x_1905 = (x_1898 & x_1904) ;
	assign x_3777 = (x_3762 & x_3776) ;
	assign x_3748 = (x_3733 & x_3747) ;
	assign x_3718 = (x_3703 & x_3717) ;
	assign x_3689 = (x_3674 & x_3688) ;
	assign x_3659 = (x_3644 & x_3658) ;
	assign x_3630 = (x_3615 & x_3629) ;
	assign x_3601 = (x_3586 & x_3600) ;
	assign x_3572 = (x_3557 & x_3571) ;
	assign x_3541 = (x_3526 & x_3540) ;
	assign x_3512 = (x_3497 & x_3511) ;
	assign x_3483 = (x_3468 & x_3482) ;
	assign x_3454 = (x_3439 & x_3453) ;
	assign x_3424 = (x_3409 & x_3423) ;
	assign x_3395 = (x_3380 & x_3394) ;
	assign x_3366 = (x_3351 & x_3365) ;
	assign x_3337 = (x_3322 & x_3336) ;
	assign x_3305 = (x_3290 & x_3304) ;
	assign x_3276 = (x_3261 & x_3275) ;
	assign x_3246 = (x_3231 & x_3245) ;
	assign x_3217 = (x_3202 & x_3216) ;
	assign x_3187 = (x_3172 & x_3186) ;
	assign x_3158 = (x_3143 & x_3157) ;
	assign x_3129 = (x_3114 & x_3128) ;
	assign x_3100 = (x_3085 & x_3099) ;
	assign x_3069 = (x_3054 & x_3068) ;
	assign x_3040 = (x_3025 & x_3039) ;
	assign x_3011 = (x_2996 & x_3010) ;
	assign x_2982 = (x_2967 & x_2981) ;
	assign x_2952 = (x_2937 & x_2951) ;
	assign x_2923 = (x_2908 & x_2922) ;
	assign x_2894 = (x_2879 & x_2893) ;
	assign x_2865 = (x_2850 & x_2864) ;
	assign x_2832 = (x_2817 & x_2831) ;
	assign x_2803 = (x_2788 & x_2802) ;
	assign x_2773 = (x_2758 & x_2772) ;
	assign x_2744 = (x_2729 & x_2743) ;
	assign x_2714 = (x_2699 & x_2713) ;
	assign x_2685 = (x_2670 & x_2684) ;
	assign x_2656 = (x_2641 & x_2655) ;
	assign x_2627 = (x_2612 & x_2626) ;
	assign x_2596 = (x_2581 & x_2595) ;
	assign x_2567 = (x_2552 & x_2566) ;
	assign x_2538 = (x_2523 & x_2537) ;
	assign x_2509 = (x_2494 & x_2508) ;
	assign x_2479 = (x_2464 & x_2478) ;
	assign x_2450 = (x_2435 & x_2449) ;
	assign x_2421 = (x_2406 & x_2420) ;
	assign x_2392 = (x_2377 & x_2391) ;
	assign x_2360 = (x_2345 & x_2359) ;
	assign x_2331 = (x_2316 & x_2330) ;
	assign x_2301 = (x_2286 & x_2300) ;
	assign x_2272 = (x_2257 & x_2271) ;
	assign x_2242 = (x_2227 & x_2241) ;
	assign x_2213 = (x_2198 & x_2212) ;
	assign x_2184 = (x_2169 & x_2183) ;
	assign x_2155 = (x_2140 & x_2154) ;
	assign x_2124 = (x_2109 & x_2123) ;
	assign x_2095 = (x_2080 & x_2094) ;
	assign x_2066 = (x_2051 & x_2065) ;
	assign x_2037 = (x_2022 & x_2036) ;
	assign x_2007 = (x_1992 & x_2006) ;
	assign x_1978 = (x_1963 & x_1977) ;
	assign x_1949 = (x_1934 & x_1948) ;
	assign x_1920 = (x_1905 & x_1919) ;
	assign x_3778 = (x_3748 & x_3777) ;
	assign x_3719 = (x_3689 & x_3718) ;
	assign x_3660 = (x_3630 & x_3659) ;
	assign x_3602 = (x_3572 & x_3601) ;
	assign x_3542 = (x_3512 & x_3541) ;
	assign x_3484 = (x_3454 & x_3483) ;
	assign x_3425 = (x_3395 & x_3424) ;
	assign x_3367 = (x_3337 & x_3366) ;
	assign x_3306 = (x_3276 & x_3305) ;
	assign x_3247 = (x_3217 & x_3246) ;
	assign x_3188 = (x_3158 & x_3187) ;
	assign x_3130 = (x_3100 & x_3129) ;
	assign x_3070 = (x_3040 & x_3069) ;
	assign x_3012 = (x_2982 & x_3011) ;
	assign x_2953 = (x_2923 & x_2952) ;
	assign x_2895 = (x_2865 & x_2894) ;
	assign x_2833 = (x_2803 & x_2832) ;
	assign x_2774 = (x_2744 & x_2773) ;
	assign x_2715 = (x_2685 & x_2714) ;
	assign x_2657 = (x_2627 & x_2656) ;
	assign x_2597 = (x_2567 & x_2596) ;
	assign x_2539 = (x_2509 & x_2538) ;
	assign x_2480 = (x_2450 & x_2479) ;
	assign x_2422 = (x_2392 & x_2421) ;
	assign x_2361 = (x_2331 & x_2360) ;
	assign x_2302 = (x_2272 & x_2301) ;
	assign x_2243 = (x_2213 & x_2242) ;
	assign x_2185 = (x_2155 & x_2184) ;
	assign x_2125 = (x_2095 & x_2124) ;
	assign x_2067 = (x_2037 & x_2066) ;
	assign x_2008 = (x_1978 & x_2007) ;
	assign x_1950 = (x_1920 & x_1949) ;
	assign x_3779 = (x_3719 & x_3778) ;
	assign x_3661 = (x_3602 & x_3660) ;
	assign x_3543 = (x_3484 & x_3542) ;
	assign x_3426 = (x_3367 & x_3425) ;
	assign x_3307 = (x_3247 & x_3306) ;
	assign x_3189 = (x_3130 & x_3188) ;
	assign x_3071 = (x_3012 & x_3070) ;
	assign x_2954 = (x_2895 & x_2953) ;
	assign x_2834 = (x_2774 & x_2833) ;
	assign x_2716 = (x_2657 & x_2715) ;
	assign x_2598 = (x_2539 & x_2597) ;
	assign x_2481 = (x_2422 & x_2480) ;
	assign x_2362 = (x_2302 & x_2361) ;
	assign x_2244 = (x_2185 & x_2243) ;
	assign x_2126 = (x_2067 & x_2125) ;
	assign x_2009 = (x_1950 & x_2008) ;
	assign x_3780 = (x_3661 & x_3779) ;
	assign x_3544 = (x_3426 & x_3543) ;
	assign x_3308 = (x_3189 & x_3307) ;
	assign x_3072 = (x_2954 & x_3071) ;
	assign x_2835 = (x_2716 & x_2834) ;
	assign x_2599 = (x_2481 & x_2598) ;
	assign x_2363 = (x_2244 & x_2362) ;
	assign x_2127 = (x_2009 & x_2126) ;
	assign x_3781 = (x_3544 & x_3780) ;
	assign x_3309 = (x_3072 & x_3308) ;
	assign x_2836 = (x_2599 & x_2835) ;
	assign x_2364 = (x_2127 & x_2363) ;
	assign x_3782 = (x_3309 & x_3781) ;
	assign x_2837 = (x_2364 & x_2836) ;
	assign x_3783 = (x_2837 & x_3782) ;
	assign v_867 = 0 ;
	assign v_866 = 0 ;
	assign v_474 = 0 ;
	assign o_1 = x_3783 ;
endmodule
