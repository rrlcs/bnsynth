// Benchmark "SKOLEMFORMULA" written by ABC on Wed May 18 01:40:47 2022

module SKOLEMFORMULA ( 
    i0,
    i1, i2  );
  input  i0;
  output i1, i2;
  assign i2 = 1'b1;
  assign i1 = i0;
endmodule


