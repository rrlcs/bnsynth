module formula(v_380,v_509,v_510,v_511,v_512,v_513,v_514,v_515,v_516,v_517,v_518,v_519,v_520,v_521,v_522,v_523,v_524,v_525,v_526,v_527,v_528,v_529,v_530,v_531,v_532,v_533,v_534,v_535,v_536,v_537,v_538,v_539,v_540,v_541,v_542,v_543,v_544,v_545,v_546,v_547,v_548,v_549,v_550,v_551,v_552,v_553,v_554,v_555,v_556,v_557,v_558,v_559,v_560,v_561,v_562,v_563,v_564,v_565,v_566,v_567,v_568,v_569,v_570,v_571,v_381,v_383,v_385,v_387,v_389,v_391,v_393,v_395,v_396,v_397,v_399,v_401,v_403,v_405,v_407,v_409,v_411,v_413,v_415,v_417,v_419,v_421,v_423,v_425,v_427,v_428,v_429,v_431,v_433,v_435,v_437,v_439,v_441,v_443,v_445,v_447,v_449,v_451,v_453,v_455,v_457,v_459,v_460,v_461,v_463,v_465,v_467,v_469,v_471,v_473,v_475,v_477,v_479,v_481,v_482,v_483,v_485,v_487,v_489,v_491,v_493,v_495,v_497,v_499,v_501,v_502,v_503,v_505,v_507,v_7,v_8,v_9,v_10,v_11,v_12,v_13,v_14,v_15,v_16,v_17,v_18,v_19,v_22,v_23,v_24,v_25,v_26,v_27,v_28,v_29,v_30,v_31,v_32,v_33,v_34,v_35,v_36,v_37,v_38,v_39,v_40,v_41,v_42,v_43,v_44,v_45,v_46,v_47,v_48,v_49,v_50,v_51,v_54,v_55,v_56,v_57,v_58,v_59,v_60,v_61,v_62,v_63,v_64,v_65,v_66,v_67,v_68,v_69,v_70,v_71,v_72,v_73,v_74,v_75,v_76,v_77,v_78,v_79,v_80,v_81,v_82,v_83,v_86,v_87,v_88,v_89,v_90,v_91,v_92,v_93,v_94,v_95,v_96,v_97,v_98,v_99,v_100,v_101,v_102,v_103,v_104,v_105,v_108,v_109,v_110,v_111,v_112,v_113,v_114,v_115,v_116,v_117,v_118,v_119,v_120,v_121,v_122,v_123,v_124,v_125,v_136,v_137,o_1);
	input v_380;
	v_509;
	v_510;
	v_511;
	v_512;
	v_513;
	v_514;
	v_515;
	v_516;
	v_517;
	v_518;
	v_519;
	v_520;
	v_521;
	v_522;
	v_523;
	v_524;
	v_525;
	v_526;
	v_527;
	v_528;
	v_529;
	v_530;
	v_531;
	v_532;
	v_533;
	v_534;
	v_535;
	v_536;
	v_537;
	v_538;
	v_539;
	v_540;
	v_541;
	v_542;
	v_543;
	v_544;
	v_545;
	v_546;
	v_547;
	v_548;
	v_549;
	v_550;
	v_551;
	v_552;
	v_553;
	v_554;
	v_555;
	v_556;
	v_557;
	v_558;
	v_559;
	v_560;
	v_561;
	v_562;
	v_563;
	v_564;
	v_565;
	v_566;
	v_567;
	v_568;
	v_569;
	v_570;
	v_571;
	v_381;
	v_383;
	v_385;
	v_387;
	v_389;
	v_391;
	v_393;
	v_395;
	v_396;
	v_397;
	v_399;
	v_401;
	v_403;
	v_405;
	v_407;
	v_409;
	v_411;
	v_413;
	v_415;
	v_417;
	v_419;
	v_421;
	v_423;
	v_425;
	v_427;
	v_428;
	v_429;
	v_431;
	v_433;
	v_435;
	v_437;
	v_439;
	v_441;
	v_443;
	v_445;
	v_447;
	v_449;
	v_451;
	v_453;
	v_455;
	v_457;
	v_459;
	v_460;
	v_461;
	v_463;
	v_465;
	v_467;
	v_469;
	v_471;
	v_473;
	v_475;
	v_477;
	v_479;
	v_481;
	v_482;
	v_483;
	v_485;
	v_487;
	v_489;
	v_491;
	v_493;
	v_495;
	v_497;
	v_499;
	v_501;
	v_502;
	v_503;
	v_505;
	v_507;
	v_7;
	v_8;
	v_9;
	v_10;
	v_11;
	v_12;
	v_13;
	v_14;
	v_15;
	v_16;
	v_17;
	v_18;
	v_19;
	v_22;
	v_23;
	v_24;
	v_25;
	v_26;
	v_27;
	v_28;
	v_29;
	v_30;
	v_31;
	v_32;
	v_33;
	v_34;
	v_35;
	v_36;
	v_37;
	v_38;
	v_39;
	v_40;
	v_41;
	v_42;
	v_43;
	v_44;
	v_45;
	v_46;
	v_47;
	v_48;
	v_49;
	v_50;
	v_51;
	v_54;
	v_55;
	v_56;
	v_57;
	v_58;
	v_59;
	v_60;
	v_61;
	v_62;
	v_63;
	v_64;
	v_65;
	v_66;
	v_67;
	v_68;
	v_69;
	v_70;
	v_71;
	v_72;
	v_73;
	v_74;
	v_75;
	v_76;
	v_77;
	v_78;
	v_79;
	v_80;
	v_81;
	v_82;
	v_83;
	v_86;
	v_87;
	v_88;
	v_89;
	v_90;
	v_91;
	v_92;
	v_93;
	v_94;
	v_95;
	v_96;
	v_97;
	v_98;
	v_99;
	v_100;
	v_101;
	v_102;
	v_103;
	v_104;
	v_105;
	v_108;
	v_109;
	v_110;
	v_111;
	v_112;
	v_113;
	v_114;
	v_115;
	v_116;
	v_117;
	v_118;
	v_119;
	v_120;
	v_121;
	v_122;
	v_123;
	v_124;
	v_125;
	v_136;
	v_137;
	wire v_382;
	wire v_384;
	wire v_386;
	wire v_388;
	wire v_390;
	wire v_392;
	wire v_394;
	wire v_398;
	wire v_400;
	wire v_402;
	wire v_404;
	wire v_406;
	wire v_408;
	wire v_410;
	wire v_412;
	wire v_414;
	wire v_416;
	wire v_418;
	wire v_420;
	wire v_422;
	wire v_424;
	wire v_426;
	wire v_430;
	wire v_432;
	wire v_434;
	wire v_436;
	wire v_438;
	wire v_440;
	wire v_442;
	wire v_444;
	wire v_446;
	wire v_448;
	wire v_450;
	wire v_452;
	wire v_454;
	wire v_456;
	wire v_458;
	wire v_462;
	wire v_464;
	wire v_466;
	wire v_468;
	wire v_470;
	wire v_472;
	wire v_474;
	wire v_476;
	wire v_478;
	wire v_480;
	wire v_484;
	wire v_486;
	wire v_488;
	wire v_490;
	wire v_492;
	wire v_494;
	wire v_496;
	wire v_498;
	wire v_500;
	wire v_504;
	wire v_506;
	wire v_508;
	wire v_1;
	wire v_2;
	wire v_3;
	wire v_4;
	wire v_5;
	wire v_6;
	wire v_20;
	wire v_21;
	wire v_52;
	wire v_53;
	wire v_84;
	wire v_85;
	wire v_106;
	wire v_107;
	wire v_126;
	wire v_127;
	wire v_128;
	wire v_129;
	wire v_130;
	wire v_131;
	wire v_132;
	wire v_133;
	wire v_134;
	wire v_135;
	wire v_138;
	wire v_139;
	wire v_140;
	wire v_141;
	wire v_142;
	wire v_143;
	wire v_144;
	wire v_145;
	wire v_146;
	wire v_147;
	wire v_148;
	wire v_149;
	wire v_150;
	wire v_151;
	wire v_152;
	wire v_153;
	wire v_154;
	wire v_155;
	wire v_156;
	wire v_157;
	wire v_158;
	wire v_159;
	wire v_160;
	wire v_161;
	wire v_162;
	wire v_163;
	wire v_164;
	wire v_165;
	wire v_166;
	wire v_167;
	wire v_168;
	wire v_169;
	wire v_170;
	wire v_171;
	wire v_172;
	wire v_173;
	wire v_174;
	wire v_175;
	wire v_176;
	wire v_177;
	wire v_178;
	wire v_179;
	wire v_180;
	wire v_181;
	wire v_182;
	wire v_183;
	wire v_184;
	wire v_185;
	wire v_186;
	wire v_187;
	wire v_188;
	wire v_189;
	wire v_190;
	wire v_191;
	wire v_192;
	wire v_193;
	wire v_194;
	wire v_195;
	wire v_196;
	wire v_197;
	wire v_198;
	wire v_199;
	wire v_200;
	wire v_201;
	wire v_202;
	wire v_203;
	wire v_204;
	wire v_205;
	wire v_206;
	wire v_207;
	wire v_208;
	wire v_209;
	wire v_210;
	wire v_211;
	wire v_212;
	wire v_213;
	wire v_214;
	wire v_215;
	wire v_216;
	wire v_217;
	wire v_218;
	wire v_219;
	wire v_220;
	wire v_221;
	wire v_222;
	wire v_223;
	wire v_224;
	wire v_225;
	wire v_226;
	wire v_227;
	wire v_228;
	wire v_229;
	wire v_230;
	wire v_231;
	wire v_232;
	wire v_233;
	wire v_234;
	wire v_235;
	wire v_236;
	wire v_237;
	wire v_238;
	wire v_239;
	wire v_240;
	wire v_241;
	wire v_242;
	wire v_243;
	wire v_244;
	wire v_245;
	wire v_246;
	wire v_247;
	wire v_248;
	wire v_249;
	wire v_250;
	wire v_251;
	wire v_252;
	wire v_253;
	wire v_254;
	wire v_255;
	wire v_256;
	wire v_257;
	wire v_258;
	wire v_259;
	wire v_260;
	wire v_261;
	wire v_262;
	wire v_263;
	wire v_264;
	wire v_265;
	wire v_266;
	wire v_267;
	wire v_268;
	wire v_269;
	wire v_270;
	wire v_271;
	wire v_272;
	wire v_273;
	wire v_274;
	wire v_275;
	wire v_276;
	wire v_277;
	wire v_278;
	wire v_279;
	wire v_280;
	wire v_281;
	wire v_282;
	wire v_283;
	wire v_284;
	wire v_285;
	wire v_286;
	wire v_287;
	wire v_288;
	wire v_289;
	wire v_290;
	wire v_291;
	wire v_292;
	wire v_293;
	wire v_294;
	wire v_295;
	wire v_296;
	wire v_297;
	wire v_298;
	wire v_299;
	wire v_300;
	wire v_301;
	wire v_302;
	wire v_303;
	wire v_304;
	wire v_305;
	wire v_306;
	wire v_307;
	wire v_308;
	wire v_309;
	wire v_310;
	wire v_311;
	wire v_312;
	wire v_313;
	wire v_314;
	wire v_315;
	wire v_316;
	wire v_317;
	wire v_318;
	wire v_319;
	wire v_320;
	wire v_321;
	wire v_322;
	wire v_323;
	wire v_324;
	wire v_325;
	wire v_326;
	wire v_327;
	wire v_328;
	wire v_329;
	wire v_330;
	wire v_331;
	wire v_332;
	wire v_333;
	wire v_334;
	wire v_335;
	wire v_336;
	wire v_337;
	wire v_338;
	wire v_339;
	wire v_340;
	wire v_341;
	wire v_342;
	wire v_343;
	wire v_344;
	wire v_345;
	wire v_346;
	wire v_347;
	wire v_348;
	wire v_349;
	wire v_350;
	wire v_351;
	wire v_352;
	wire v_353;
	wire v_354;
	wire v_355;
	wire v_356;
	wire v_357;
	wire v_358;
	wire v_359;
	wire v_360;
	wire v_361;
	wire v_362;
	wire v_363;
	wire v_364;
	wire v_365;
	wire v_366;
	wire v_367;
	wire v_368;
	wire v_369;
	wire v_370;
	wire v_371;
	wire v_372;
	wire v_373;
	wire v_374;
	wire v_375;
	wire v_376;
	wire v_377;
	wire v_378;
	wire v_379;
	wire v_572;
	wire x_1;
	wire x_2;
	wire x_3;
	wire x_4;
	wire x_5;
	wire x_6;
	wire x_7;
	wire x_8;
	wire x_9;
	wire x_10;
	wire x_11;
	wire x_12;
	wire x_13;
	wire x_14;
	wire x_15;
	wire x_16;
	wire x_17;
	wire x_18;
	wire x_19;
	wire x_20;
	wire x_21;
	wire x_22;
	wire x_23;
	wire x_24;
	wire x_25;
	wire x_26;
	wire x_27;
	wire x_28;
	wire x_29;
	wire x_30;
	wire x_31;
	wire x_32;
	wire x_33;
	wire x_34;
	wire x_35;
	wire x_36;
	wire x_37;
	wire x_38;
	wire x_39;
	wire x_40;
	wire x_41;
	wire x_42;
	wire x_43;
	wire x_44;
	wire x_45;
	wire x_46;
	wire x_47;
	wire x_48;
	wire x_49;
	wire x_50;
	wire x_51;
	wire x_52;
	wire x_53;
	wire x_54;
	wire x_55;
	wire x_56;
	wire x_57;
	wire x_58;
	wire x_59;
	wire x_60;
	wire x_61;
	wire x_62;
	wire x_63;
	wire x_64;
	wire x_65;
	wire x_66;
	wire x_67;
	wire x_68;
	wire x_69;
	wire x_70;
	wire x_71;
	wire x_72;
	wire x_73;
	wire x_74;
	wire x_75;
	wire x_76;
	wire x_77;
	wire x_78;
	wire x_79;
	wire x_80;
	wire x_81;
	wire x_82;
	wire x_83;
	wire x_84;
	wire x_85;
	wire x_86;
	wire x_87;
	wire x_88;
	wire x_89;
	wire x_90;
	wire x_91;
	wire x_92;
	wire x_93;
	wire x_94;
	wire x_95;
	wire x_96;
	wire x_97;
	wire x_98;
	wire x_99;
	wire x_100;
	wire x_101;
	wire x_102;
	wire x_103;
	wire x_104;
	wire x_105;
	wire x_106;
	wire x_107;
	wire x_108;
	wire x_109;
	wire x_110;
	wire x_111;
	wire x_112;
	wire x_113;
	wire x_114;
	wire x_115;
	wire x_116;
	wire x_117;
	wire x_118;
	wire x_119;
	wire x_120;
	wire x_121;
	wire x_122;
	wire x_123;
	wire x_124;
	wire x_125;
	wire x_126;
	wire x_127;
	wire x_128;
	wire x_129;
	wire x_130;
	wire x_131;
	wire x_132;
	wire x_133;
	wire x_134;
	wire x_135;
	wire x_136;
	wire x_137;
	wire x_138;
	wire x_139;
	wire x_140;
	wire x_141;
	wire x_142;
	wire x_143;
	wire x_144;
	wire x_145;
	wire x_146;
	wire x_147;
	wire x_148;
	wire x_149;
	wire x_150;
	wire x_151;
	wire x_152;
	wire x_153;
	wire x_154;
	wire x_155;
	wire x_156;
	wire x_157;
	wire x_158;
	wire x_159;
	wire x_160;
	wire x_161;
	wire x_162;
	wire x_163;
	wire x_164;
	wire x_165;
	wire x_166;
	wire x_167;
	wire x_168;
	wire x_169;
	wire x_170;
	wire x_171;
	wire x_172;
	wire x_173;
	wire x_174;
	wire x_175;
	wire x_176;
	wire x_177;
	wire x_178;
	wire x_179;
	wire x_180;
	wire x_181;
	wire x_182;
	wire x_183;
	wire x_184;
	wire x_185;
	wire x_186;
	wire x_187;
	wire x_188;
	wire x_189;
	wire x_190;
	wire x_191;
	wire x_192;
	wire x_193;
	wire x_194;
	wire x_195;
	wire x_196;
	wire x_197;
	wire x_198;
	wire x_199;
	wire x_200;
	wire x_201;
	wire x_202;
	wire x_203;
	wire x_204;
	wire x_205;
	wire x_206;
	wire x_207;
	wire x_208;
	wire x_209;
	wire x_210;
	wire x_211;
	wire x_212;
	wire x_213;
	wire x_214;
	wire x_215;
	wire x_216;
	wire x_217;
	wire x_218;
	wire x_219;
	wire x_220;
	wire x_221;
	wire x_222;
	wire x_223;
	wire x_224;
	wire x_225;
	wire x_226;
	wire x_227;
	wire x_228;
	wire x_229;
	wire x_230;
	wire x_231;
	wire x_232;
	wire x_233;
	wire x_234;
	wire x_235;
	wire x_236;
	wire x_237;
	wire x_238;
	wire x_239;
	wire x_240;
	wire x_241;
	wire x_242;
	wire x_243;
	wire x_244;
	wire x_245;
	wire x_246;
	wire x_247;
	wire x_248;
	wire x_249;
	wire x_250;
	wire x_251;
	wire x_252;
	wire x_253;
	wire x_254;
	wire x_255;
	wire x_256;
	wire x_257;
	wire x_258;
	wire x_259;
	wire x_260;
	wire x_261;
	wire x_262;
	wire x_263;
	wire x_264;
	wire x_265;
	wire x_266;
	wire x_267;
	wire x_268;
	wire x_269;
	wire x_270;
	wire x_271;
	wire x_272;
	wire x_273;
	wire x_274;
	wire x_275;
	wire x_276;
	wire x_277;
	wire x_278;
	wire x_279;
	wire x_280;
	wire x_281;
	wire x_282;
	wire x_283;
	wire x_284;
	wire x_285;
	wire x_286;
	wire x_287;
	wire x_288;
	wire x_289;
	wire x_290;
	wire x_291;
	wire x_292;
	wire x_293;
	wire x_294;
	wire x_295;
	wire x_296;
	wire x_297;
	wire x_298;
	wire x_299;
	wire x_300;
	wire x_301;
	wire x_302;
	wire x_303;
	wire x_304;
	wire x_305;
	wire x_306;
	wire x_307;
	wire x_308;
	wire x_309;
	wire x_310;
	wire x_311;
	wire x_312;
	wire x_313;
	wire x_314;
	wire x_315;
	wire x_316;
	wire x_317;
	wire x_318;
	wire x_319;
	wire x_320;
	wire x_321;
	wire x_322;
	wire x_323;
	wire x_324;
	wire x_325;
	wire x_326;
	wire x_327;
	wire x_328;
	wire x_329;
	wire x_330;
	wire x_331;
	wire x_332;
	wire x_333;
	wire x_334;
	wire x_335;
	wire x_336;
	wire x_337;
	wire x_338;
	wire x_339;
	wire x_340;
	wire x_341;
	wire x_342;
	wire x_343;
	wire x_344;
	wire x_345;
	wire x_346;
	wire x_347;
	wire x_348;
	wire x_349;
	wire x_350;
	wire x_351;
	wire x_352;
	wire x_353;
	wire x_354;
	wire x_355;
	wire x_356;
	wire x_357;
	wire x_358;
	wire x_359;
	wire x_360;
	wire x_361;
	wire x_362;
	wire x_363;
	wire x_364;
	wire x_365;
	wire x_366;
	wire x_367;
	wire x_368;
	wire x_369;
	wire x_370;
	wire x_371;
	wire x_372;
	wire x_373;
	wire x_374;
	wire x_375;
	wire x_376;
	wire x_377;
	wire x_378;
	wire x_379;
	wire x_380;
	wire x_381;
	wire x_382;
	wire x_383;
	wire x_384;
	wire x_385;
	wire x_386;
	wire x_387;
	wire x_388;
	wire x_389;
	wire x_390;
	wire x_391;
	wire x_392;
	wire x_393;
	wire x_394;
	wire x_395;
	wire x_396;
	wire x_397;
	wire x_398;
	wire x_399;
	wire x_400;
	wire x_401;
	wire x_402;
	wire x_403;
	wire x_404;
	wire x_405;
	wire x_406;
	wire x_407;
	wire x_408;
	wire x_409;
	wire x_410;
	wire x_411;
	wire x_412;
	wire x_413;
	wire x_414;
	wire x_415;
	wire x_416;
	wire x_417;
	wire x_418;
	wire x_419;
	wire x_420;
	wire x_421;
	wire x_422;
	wire x_423;
	wire x_424;
	wire x_425;
	wire x_426;
	wire x_427;
	wire x_428;
	wire x_429;
	wire x_430;
	wire x_431;
	wire x_432;
	wire x_433;
	wire x_434;
	wire x_435;
	wire x_436;
	wire x_437;
	wire x_438;
	wire x_439;
	wire x_440;
	wire x_441;
	wire x_442;
	wire x_443;
	wire x_444;
	wire x_445;
	wire x_446;
	wire x_447;
	wire x_448;
	wire x_449;
	wire x_450;
	wire x_451;
	wire x_452;
	wire x_453;
	wire x_454;
	wire x_455;
	wire x_456;
	wire x_457;
	wire x_458;
	wire x_459;
	wire x_460;
	wire x_461;
	wire x_462;
	wire x_463;
	wire x_464;
	wire x_465;
	wire x_466;
	wire x_467;
	wire x_468;
	wire x_469;
	wire x_470;
	wire x_471;
	wire x_472;
	wire x_473;
	wire x_474;
	wire x_475;
	wire x_476;
	wire x_477;
	wire x_478;
	wire x_479;
	wire x_480;
	wire x_481;
	wire x_482;
	wire x_483;
	wire x_484;
	wire x_485;
	wire x_486;
	wire x_487;
	wire x_488;
	wire x_489;
	wire x_490;
	wire x_491;
	wire x_492;
	wire x_493;
	wire x_494;
	wire x_495;
	wire x_496;
	wire x_497;
	wire x_498;
	wire x_499;
	wire x_500;
	wire x_501;
	wire x_502;
	wire x_503;
	wire x_504;
	wire x_505;
	wire x_506;
	wire x_507;
	wire x_508;
	wire x_509;
	wire x_510;
	wire x_511;
	wire x_512;
	wire x_513;
	wire x_514;
	wire x_515;
	wire x_516;
	wire x_517;
	wire x_518;
	wire x_519;
	wire x_520;
	wire x_521;
	wire x_522;
	wire x_523;
	wire x_524;
	wire x_525;
	wire x_526;
	wire x_527;
	wire x_528;
	wire x_529;
	wire x_530;
	wire x_531;
	wire x_532;
	wire x_533;
	wire x_534;
	wire x_535;
	wire x_536;
	wire x_537;
	wire x_538;
	wire x_539;
	wire x_540;
	wire x_541;
	wire x_542;
	wire x_543;
	wire x_544;
	wire x_545;
	wire x_546;
	wire x_547;
	wire x_548;
	wire x_549;
	wire x_550;
	wire x_551;
	wire x_552;
	wire x_553;
	wire x_554;
	wire x_555;
	wire x_556;
	wire x_557;
	wire x_558;
	wire x_559;
	wire x_560;
	wire x_561;
	wire x_562;
	wire x_563;
	wire x_564;
	wire x_565;
	wire x_566;
	wire x_567;
	wire x_568;
	wire x_569;
	wire x_570;
	wire x_571;
	wire x_572;
	wire x_573;
	wire x_574;
	wire x_575;
	wire x_576;
	wire x_577;
	wire x_578;
	wire x_579;
	wire x_580;
	wire x_581;
	wire x_582;
	wire x_583;
	wire x_584;
	wire x_585;
	wire x_586;
	wire x_587;
	wire x_588;
	wire x_589;
	wire x_590;
	wire x_591;
	wire x_592;
	wire x_593;
	wire x_594;
	wire x_595;
	wire x_596;
	wire x_597;
	wire x_598;
	wire x_599;
	wire x_600;
	wire x_601;
	wire x_602;
	wire x_603;
	wire x_604;
	wire x_605;
	wire x_606;
	wire x_607;
	wire x_608;
	wire x_609;
	wire x_610;
	wire x_611;
	wire x_612;
	wire x_613;
	wire x_614;
	wire x_615;
	wire x_616;
	wire x_617;
	wire x_618;
	wire x_619;
	wire x_620;
	wire x_621;
	wire x_622;
	wire x_623;
	wire x_624;
	wire x_625;
	wire x_626;
	wire x_627;
	wire x_628;
	wire x_629;
	wire x_630;
	wire x_631;
	wire x_632;
	wire x_633;
	wire x_634;
	wire x_635;
	wire x_636;
	wire x_637;
	wire x_638;
	wire x_639;
	wire x_640;
	wire x_641;
	wire x_642;
	wire x_643;
	wire x_644;
	wire x_645;
	wire x_646;
	wire x_647;
	wire x_648;
	wire x_649;
	wire x_650;
	wire x_651;
	wire x_652;
	wire x_653;
	wire x_654;
	wire x_655;
	wire x_656;
	wire x_657;
	wire x_658;
	wire x_659;
	wire x_660;
	wire x_661;
	wire x_662;
	wire x_663;
	wire x_664;
	wire x_665;
	wire x_666;
	wire x_667;
	wire x_668;
	wire x_669;
	wire x_670;
	wire x_671;
	wire x_672;
	wire x_673;
	wire x_674;
	wire x_675;
	wire x_676;
	wire x_677;
	wire x_678;
	wire x_679;
	wire x_680;
	wire x_681;
	wire x_682;
	wire x_683;
	wire x_684;
	wire x_685;
	wire x_686;
	wire x_687;
	wire x_688;
	wire x_689;
	wire x_690;
	wire x_691;
	wire x_692;
	wire x_693;
	wire x_694;
	wire x_695;
	wire x_696;
	wire x_697;
	wire x_698;
	wire x_699;
	wire x_700;
	wire x_701;
	wire x_702;
	wire x_703;
	wire x_704;
	wire x_705;
	wire x_706;
	wire x_707;
	wire x_708;
	wire x_709;
	wire x_710;
	wire x_711;
	wire x_712;
	wire x_713;
	wire x_714;
	wire x_715;
	wire x_716;
	wire x_717;
	wire x_718;
	wire x_719;
	wire x_720;
	wire x_721;
	wire x_722;
	wire x_723;
	wire x_724;
	wire x_725;
	wire x_726;
	wire x_727;
	wire x_728;
	wire x_729;
	wire x_730;
	wire x_731;
	wire x_732;
	wire x_733;
	wire x_734;
	wire x_735;
	wire x_736;
	wire x_737;
	wire x_738;
	wire x_739;
	wire x_740;
	wire x_741;
	wire x_742;
	wire x_743;
	wire x_744;
	wire x_745;
	wire x_746;
	wire x_747;
	wire x_748;
	wire x_749;
	wire x_750;
	wire x_751;
	wire x_752;
	wire x_753;
	wire x_754;
	wire x_755;
	wire x_756;
	wire x_757;
	wire x_758;
	wire x_759;
	wire x_760;
	wire x_761;
	wire x_762;
	wire x_763;
	wire x_764;
	wire x_765;
	wire x_766;
	wire x_767;
	wire x_768;
	wire x_769;
	wire x_770;
	wire x_771;
	wire x_772;
	wire x_773;
	wire x_774;
	wire x_775;
	wire x_776;
	wire x_777;
	wire x_778;
	wire x_779;
	wire x_780;
	wire x_781;
	wire x_782;
	wire x_783;
	wire x_784;
	wire x_785;
	wire x_786;
	wire x_787;
	wire x_788;
	wire x_789;
	wire x_790;
	wire x_791;
	wire x_792;
	wire x_793;
	wire x_794;
	wire x_795;
	wire x_796;
	wire x_797;
	wire x_798;
	wire x_799;
	wire x_800;
	wire x_801;
	wire x_802;
	wire x_803;
	wire x_804;
	wire x_805;
	wire x_806;
	wire x_807;
	wire x_808;
	wire x_809;
	wire x_810;
	wire x_811;
	wire x_812;
	wire x_813;
	wire x_814;
	wire x_815;
	wire x_816;
	wire x_817;
	wire x_818;
	wire x_819;
	wire x_820;
	wire x_821;
	wire x_822;
	wire x_823;
	wire x_824;
	wire x_825;
	wire x_826;
	wire x_827;
	wire x_828;
	wire x_829;
	wire x_830;
	wire x_831;
	wire x_832;
	wire x_833;
	wire x_834;
	wire x_835;
	wire x_836;
	wire x_837;
	wire x_838;
	wire x_839;
	wire x_840;
	wire x_841;
	wire x_842;
	wire x_843;
	wire x_844;
	wire x_845;
	wire x_846;
	wire x_847;
	wire x_848;
	wire x_849;
	wire x_850;
	wire x_851;
	wire x_852;
	wire x_853;
	wire x_854;
	wire x_855;
	wire x_856;
	wire x_857;
	wire x_858;
	wire x_859;
	wire x_860;
	wire x_861;
	wire x_862;
	wire x_863;
	wire x_864;
	wire x_865;
	wire x_866;
	wire x_867;
	wire x_868;
	wire x_869;
	wire x_870;
	wire x_871;
	wire x_872;
	wire x_873;
	wire x_874;
	wire x_875;
	wire x_876;
	wire x_877;
	wire x_878;
	wire x_879;
	wire x_880;
	wire x_881;
	wire x_882;
	wire x_883;
	wire x_884;
	wire x_885;
	wire x_886;
	wire x_887;
	wire x_888;
	wire x_889;
	wire x_890;
	wire x_891;
	wire x_892;
	wire x_893;
	wire x_894;
	wire x_895;
	wire x_896;
	wire x_897;
	wire x_898;
	wire x_899;
	wire x_900;
	wire x_901;
	wire x_902;
	wire x_903;
	wire x_904;
	wire x_905;
	wire x_906;
	wire x_907;
	wire x_908;
	wire x_909;
	wire x_910;
	wire x_911;
	wire x_912;
	wire x_913;
	wire x_914;
	wire x_915;
	wire x_916;
	wire x_917;
	wire x_918;
	wire x_919;
	wire x_920;
	wire x_921;
	wire x_922;
	wire x_923;
	wire x_924;
	wire x_925;
	wire x_926;
	wire x_927;
	wire x_928;
	wire x_929;
	wire x_930;
	wire x_931;
	wire x_932;
	wire x_933;
	wire x_934;
	wire x_935;
	wire x_936;
	wire x_937;
	wire x_938;
	wire x_939;
	wire x_940;
	wire x_941;
	wire x_942;
	wire x_943;
	wire x_944;
	wire x_945;
	wire x_946;
	wire x_947;
	wire x_948;
	wire x_949;
	wire x_950;
	wire x_951;
	wire x_952;
	wire x_953;
	wire x_954;
	wire x_955;
	wire x_956;
	wire x_957;
	wire x_958;
	wire x_959;
	wire x_960;
	wire x_961;
	wire x_962;
	wire x_963;
	wire x_964;
	wire x_965;
	wire x_966;
	wire x_967;
	wire x_968;
	wire x_969;
	wire x_970;
	wire x_971;
	wire x_972;
	wire x_973;
	wire x_974;
	wire x_975;
	wire x_976;
	wire x_977;
	wire x_978;
	wire x_979;
	wire x_980;
	wire x_981;
	wire x_982;
	wire x_983;
	wire x_984;
	wire x_985;
	wire x_986;
	wire x_987;
	wire x_988;
	wire x_989;
	wire x_990;
	wire x_991;
	wire x_992;
	wire x_993;
	wire x_994;
	wire x_995;
	wire x_996;
	wire x_997;
	wire x_998;
	wire x_999;
	wire x_1000;
	wire x_1001;
	wire x_1002;
	wire x_1003;
	wire x_1004;
	wire x_1005;
	wire x_1006;
	wire x_1007;
	wire x_1008;
	wire x_1009;
	wire x_1010;
	wire x_1011;
	wire x_1012;
	wire x_1013;
	wire x_1014;
	wire x_1015;
	wire x_1016;
	wire x_1017;
	wire x_1018;
	wire x_1019;
	wire x_1020;
	wire x_1021;
	wire x_1022;
	wire x_1023;
	wire x_1024;
	wire x_1025;
	wire x_1026;
	wire x_1027;
	wire x_1028;
	wire x_1029;
	wire x_1030;
	wire x_1031;
	wire x_1032;
	wire x_1033;
	wire x_1034;
	wire x_1035;
	wire x_1036;
	wire x_1037;
	wire x_1038;
	wire x_1039;
	wire x_1040;
	wire x_1041;
	wire x_1042;
	wire x_1043;
	wire x_1044;
	wire x_1045;
	wire x_1046;
	wire x_1047;
	wire x_1048;
	wire x_1049;
	wire x_1050;
	wire x_1051;
	wire x_1052;
	wire x_1053;
	wire x_1054;
	wire x_1055;
	wire x_1056;
	wire x_1057;
	wire x_1058;
	wire x_1059;
	output o_1;
	assign v_6 = v_50);
	assign v_142 = v_51);
	assign v_145 = v_51);
	assign v_149 = v_51);
	assign v_152 = v_51);
	assign v_156 = v_51);
	assign v_159 = v_51);
	assign v_163 = v_51);
	assign v_165 = v_51);
	assign v_169 = v_51);
	assign v_172 = v_51);
	assign v_176 = v_52);
	assign v_179 = v_52);
	assign v_183 = v_52);
	assign v_186 = v_52);
	assign v_190 = v_52);
	assign v_193 = v_52);
	assign v_197 = v_52);
	assign v_200 = v_52);
	assign v_204 = v_52);
	assign v_207 = v_52);
	assign v_211 = v_53);
	assign v_214 = v_53);
	assign v_218 = v_53);
	assign v_220 = v_53);
	assign v_224 = v_53);
	assign v_227 = v_53);
	assign v_231 = v_53);
	assign v_234 = v_53);
	assign v_238 = v_53);
	assign v_241 = v_53);
	assign v_245 = v_54);
	assign v_248 = v_54);
	assign v_252 = v_54);
	assign v_255 = v_54);
	assign v_259 = v_54);
	assign v_262 = v_54);
	assign v_266 = v_54);
	assign v_269 = v_54);
	assign v_273 = v_54);
	assign v_275 = v_54);
	assign v_279 = v_55);
	assign v_282 = v_55);
	assign v_286 = v_55);
	assign v_289 = v_55);
	assign v_293 = v_55);
	assign v_296 = v_55);
	assign v_300 = v_55);
	assign v_303 = v_55);
	assign v_307 = v_55);
	assign v_310 = v_55);
	assign v_313 = v_56);
	assign v_316 = v_56);
	assign v_320 = v_56);
	assign v_323 = v_56);
	assign v_327 = v_56);
	assign v_330 = v_56);
	assign v_334 = v_56);
	assign v_337 = v_56);
	assign v_340 = v_56);
	assign v_344 = v_56);
	assign v_346 = v_57);
	assign v_349 = v_57);
	assign v_133 = (v_395 ^ v_396);
	assign v_132 = (v_427 ^ v_428);
	assign v_131 = (v_459 ^ v_460);
	assign v_130 = (v_481 ^ v_482);
	assign v_129 = (v_501 ^ v_502);
	assign x_3 = (~v_7 | ~v_8);
	assign x_1 = (((v_7 | v_383)) | v_8);
	assign x_7 = (~v_8 | ~v_9);
	assign x_12 = (~v_9 | ~v_10);
	assign x_10 = (((v_9 | v_385)) | v_10);
	assign x_16 = (~v_10 | ~v_11);
	assign x_21 = (~v_11 | ~v_12);
	assign x_19 = (((v_11 | v_387)) | v_12);
	assign x_25 = (~v_12 | ~v_13);
	assign x_30 = (~v_13 | ~v_14);
	assign x_28 = (((v_13 | v_389)) | v_14);
	assign x_34 = (~v_14 | ~v_15);
	assign x_39 = (~v_15 | ~v_16);
	assign x_37 = (((v_15 | v_391)) | v_16);
	assign x_43 = (~v_16 | ~v_17);
	assign x_48 = (~v_17 | ~v_18);
	assign x_46 = (((v_17 | v_393)) | v_18);
	assign x_58 = (((~v_19 | ~v_395)) | ~v_396);
	assign x_52 = (~v_18 | ~v_19);
	assign x_65 = (~v_22 | ~v_23);
	assign x_70 = (~v_23 | ~v_24);
	assign x_68 = (((v_23 | v_399)) | v_24);
	assign x_74 = (~v_24 | ~v_25);
	assign x_79 = (~v_25 | ~v_26);
	assign x_77 = (((v_25 | v_401)) | v_26);
	assign x_83 = (~v_26 | ~v_27);
	assign x_88 = (~v_27 | ~v_28);
	assign x_86 = (((v_27 | v_403)) | v_28);
	assign x_92 = (~v_28 | ~v_29);
	assign x_97 = (~v_29 | ~v_30);
	assign x_95 = (((v_29 | v_405)) | v_30);
	assign x_101 = (~v_30 | ~v_31);
	assign x_106 = (~v_31 | ~v_32);
	assign x_104 = (((v_31 | v_407)) | v_32);
	assign x_110 = (~v_32 | ~v_33);
	assign x_115 = (~v_33 | ~v_34);
	assign x_113 = (((v_33 | v_409)) | v_34);
	assign x_119 = (~v_34 | ~v_35);
	assign x_124 = (~v_35 | ~v_36);
	assign x_122 = (((v_35 | v_411)) | v_36);
	assign x_128 = (~v_36 | ~v_37);
	assign x_131 = (((v_37 | v_413)) | v_38);
	assign x_133 = (~v_37 | ~v_38);
	assign x_137 = (~v_38 | ~v_39);
	assign x_142 = (~v_39 | ~v_40);
	assign x_140 = (((v_39 | v_415)) | v_40);
	assign x_146 = (~v_40 | ~v_41);
	assign x_151 = (~v_41 | ~v_42);
	assign x_149 = (((v_41 | v_417)) | v_42);
	assign x_155 = (~v_42 | ~v_43);
	assign x_160 = (~v_43 | ~v_44);
	assign x_158 = (((v_43 | v_419)) | v_44);
	assign x_164 = (~v_44 | ~v_45);
	assign x_169 = (~v_45 | ~v_46);
	assign x_167 = (((v_45 | v_421)) | v_46);
	assign x_173 = (~v_46 | ~v_47);
	assign x_178 = (~v_47 | ~v_48);
	assign x_176 = (((v_47 | v_423)) | v_48);
	assign x_182 = (~v_48 | ~v_49);
	assign x_187 = (~v_49 | ~v_50);
	assign x_185 = (((v_49 | v_425)) | v_50);
	assign x_197 = (((~v_51 | ~v_427)) | ~v_428);
	assign x_191 = (~v_50 | ~v_51);
	assign x_204 = (~v_54 | ~v_55);
	assign x_209 = (~v_55 | ~v_56);
	assign x_207 = (((v_55 | v_431)) | v_56);
	assign x_213 = (~v_56 | ~v_57);
	assign x_218 = (~v_57 | ~v_58);
	assign x_216 = (((v_57 | v_433)) | v_58);
	assign x_222 = (~v_58 | ~v_59);
	assign x_227 = (~v_59 | ~v_60);
	assign x_225 = (((v_59 | v_435)) | v_60);
	assign x_231 = (~v_60 | ~v_61);
	assign x_236 = (~v_61 | ~v_62);
	assign x_234 = (((v_61 | v_437)) | v_62);
	assign x_240 = (~v_62 | ~v_63);
	assign x_245 = (~v_63 | ~v_64);
	assign x_243 = (((v_63 | v_439)) | v_64);
	assign x_249 = (~v_64 | ~v_65);
	assign x_254 = (~v_65 | ~v_66);
	assign x_252 = (((v_65 | v_441)) | v_66);
	assign x_258 = (~v_66 | ~v_67);
	assign x_263 = (~v_67 | ~v_68);
	assign x_261 = (((v_67 | v_443)) | v_68);
	assign x_267 = (~v_68 | ~v_69);
	assign x_272 = (~v_69 | ~v_70);
	assign x_270 = (((v_69 | v_445)) | v_70);
	assign x_276 = (~v_70 | ~v_71);
	assign x_281 = (~v_71 | ~v_72);
	assign x_279 = (((v_71 | v_447)) | v_72);
	assign x_285 = (~v_72 | ~v_73);
	assign x_290 = (~v_73 | ~v_74);
	assign x_288 = (((v_73 | v_449)) | v_74);
	assign x_294 = (~v_74 | ~v_75);
	assign x_297 = (((v_75 | v_451)) | v_76);
	assign x_299 = (~v_75 | ~v_76);
	assign x_303 = (~v_76 | ~v_77);
	assign x_308 = (~v_77 | ~v_78);
	assign x_306 = (((v_77 | v_453)) | v_78);
	assign x_312 = (~v_78 | ~v_79);
	assign x_317 = (~v_79 | ~v_80);
	assign x_315 = (((v_79 | v_455)) | v_80);
	assign x_321 = (~v_80 | ~v_81);
	assign x_326 = (~v_81 | ~v_82);
	assign x_324 = (((v_81 | v_457)) | v_82);
	assign x_330 = (~v_82 | ~v_83);
	assign x_336 = (((~v_83 | ~v_459)) | ~v_460);
	assign x_343 = (~v_86 | ~v_87);
	assign x_348 = (~v_87 | ~v_88);
	assign x_346 = (((v_87 | v_463)) | v_88);
	assign x_352 = (~v_88 | ~v_89);
	assign x_357 = (~v_89 | ~v_90);
	assign x_355 = (((v_89 | v_465)) | v_90);
	assign x_361 = (~v_90 | ~v_91);
	assign x_364 = (((v_91 | v_467)) | v_92);
	assign x_366 = (~v_91 | ~v_92);
	assign x_370 = (~v_92 | ~v_93);
	assign x_375 = (~v_93 | ~v_94);
	assign x_373 = (((v_93 | v_469)) | v_94);
	assign x_379 = (~v_94 | ~v_95);
	assign x_384 = (~v_95 | ~v_96);
	assign x_382 = (((v_95 | v_471)) | v_96);
	assign x_388 = (~v_96 | ~v_97);
	assign x_393 = (~v_97 | ~v_98);
	assign x_391 = (((v_97 | v_473)) | v_98);
	assign x_397 = (~v_98 | ~v_99);
	assign x_402 = (~v_99 | ~v_100);
	assign x_400 = (((v_99 | v_475)) | v_100);
	assign x_406 = (~v_100 | ~v_101);
	assign x_411 = (~v_101 | ~v_102);
	assign x_409 = (((v_101 | v_477)) | v_102);
	assign x_415 = (~v_102 | ~v_103);
	assign x_420 = (~v_103 | ~v_104);
	assign x_418 = (((v_103 | v_479)) | v_104);
	assign x_430 = (((~v_105 | ~v_481)) | ~v_482);
	assign x_424 = (~v_104 | ~v_105);
	assign x_437 = (~v_108 | ~v_109);
	assign x_442 = (~v_109 | ~v_110);
	assign x_440 = (((v_109 | v_485)) | v_110);
	assign x_446 = (~v_110 | ~v_111);
	assign x_451 = (~v_111 | ~v_112);
	assign x_449 = (((v_111 | v_487)) | v_112);
	assign x_455 = (~v_112 | ~v_113);
	assign x_460 = (~v_113 | ~v_114);
	assign x_458 = (((v_113 | v_489)) | v_114);
	assign x_464 = (~v_114 | ~v_115);
	assign x_469 = (~v_115 | ~v_116);
	assign x_467 = (((v_115 | v_491)) | v_116);
	assign x_473 = (~v_116 | ~v_117);
	assign x_478 = (~v_117 | ~v_118);
	assign x_476 = (((v_117 | v_493)) | v_118);
	assign x_482 = (~v_118 | ~v_119);
	assign x_487 = (~v_119 | ~v_120);
	assign x_485 = (((v_119 | v_495)) | v_120);
	assign x_491 = (~v_120 | ~v_121);
	assign x_496 = (~v_121 | ~v_122);
	assign x_494 = (((v_121 | v_497)) | v_122);
	assign x_500 = (~v_122 | ~v_123);
	assign x_505 = (~v_123 | ~v_124);
	assign x_503 = (((v_123 | v_499)) | v_124);
	assign x_515 = (((~v_125 | ~v_501)) | ~v_502);
	assign x_509 = (~v_124 | ~v_125);
	assign v_138 = ~v_13);
	assign x_528 = (~v_137 | ~v_7);
	assign x_524 = (~v_136 | ~v_137);
	assign x_522 = (((v_136 | v_381)) | v_137);
	assign v_134 = (v_6 ^ ~v_7);
	assign v_143 = (v_142 ^ ~v_9);
	assign v_146 = (v_145 ^ ~v_11);
	assign v_150 = (v_149 ^ ~v_13);
	assign v_153 = (v_152 ^ ~v_15);
	assign v_157 = (v_156 ^ ~v_17);
	assign v_160 = (v_159 ^ ~v_19);
	assign v_166 = (v_165 ^ ~v_23);
	assign v_170 = (v_169 ^ ~v_25);
	assign v_173 = (v_172 ^ ~v_27);
	assign v_177 = (v_176 ^ ~v_29);
	assign v_180 = (v_179 ^ ~v_31);
	assign v_184 = (v_183 ^ ~v_33);
	assign v_187 = (v_186 ^ ~v_35);
	assign v_191 = (v_190 ^ ~v_37);
	assign v_194 = (v_193 ^ ~v_39);
	assign v_198 = (v_197 ^ ~v_41);
	assign v_201 = (v_200 ^ ~v_43);
	assign v_205 = (v_204 ^ ~v_45);
	assign v_208 = (v_207 ^ ~v_47);
	assign v_212 = (v_211 ^ ~v_49);
	assign v_215 = (v_214 ^ ~v_51);
	assign v_221 = (v_220 ^ ~v_55);
	assign v_225 = (v_224 ^ ~v_57);
	assign v_228 = (v_227 ^ ~v_59);
	assign v_232 = (v_231 ^ ~v_61);
	assign v_235 = (v_234 ^ ~v_63);
	assign v_239 = (v_238 ^ ~v_65);
	assign v_242 = (v_241 ^ ~v_67);
	assign v_246 = (v_245 ^ ~v_69);
	assign v_249 = (v_248 ^ ~v_71);
	assign v_253 = (v_252 ^ ~v_73);
	assign v_256 = (v_255 ^ ~v_75);
	assign v_260 = (v_259 ^ ~v_77);
	assign v_263 = (v_262 ^ ~v_79);
	assign v_267 = (v_266 ^ ~v_81);
	assign v_270 = (v_269 ^ ~v_83);
	assign v_276 = (v_275 ^ ~v_87);
	assign v_280 = (v_279 ^ ~v_89);
	assign v_283 = (v_282 ^ ~v_91);
	assign v_287 = (v_286 ^ ~v_93);
	assign v_290 = (v_289 ^ ~v_95);
	assign v_294 = (v_293 ^ ~v_97);
	assign v_297 = (v_296 ^ ~v_99);
	assign v_301 = (v_300 ^ ~v_101);
	assign v_304 = (v_303 ^ ~v_103);
	assign v_308 = (v_307 ^ ~v_105);
	assign v_314 = (v_313 ^ ~v_109);
	assign v_317 = (v_316 ^ ~v_111);
	assign v_321 = (v_320 ^ ~v_113);
	assign v_324 = (v_323 ^ ~v_115);
	assign v_328 = (v_327 ^ ~v_117);
	assign v_331 = (v_330 ^ ~v_119);
	assign v_335 = (v_334 ^ ~v_121);
	assign v_338 = (v_337 ^ ~v_123);
	assign v_341 = (v_340 ^ ~v_125);
	assign v_506 = (v_349 ^ v_505);
	assign v_21 = (v_163 ^ ~v_133);
	assign v_53 = (v_218 ^ ~v_132);
	assign v_85 = (v_273 ^ ~v_131);
	assign v_107 = (v_310 ^ ~v_130);
	assign v_127 = (v_344 ^ ~v_129);
	assign v_139 = (v_138 ^ v_380);
	assign v_382 = (v_134 ^ v_381);
	assign v_384 = (v_143 ^ v_383);
	assign v_386 = (v_146 ^ v_385);
	assign v_388 = (v_150 ^ v_387);
	assign v_390 = (v_153 ^ v_389);
	assign v_392 = (v_157 ^ v_391);
	assign v_394 = (v_160 ^ v_393);
	assign v_398 = (v_166 ^ v_397);
	assign v_400 = (v_170 ^ v_399);
	assign v_402 = (v_173 ^ v_401);
	assign v_404 = (v_177 ^ v_403);
	assign v_406 = (v_180 ^ v_405);
	assign v_408 = (v_184 ^ v_407);
	assign v_410 = (v_187 ^ v_409);
	assign v_412 = (v_191 ^ v_411);
	assign v_414 = (v_194 ^ v_413);
	assign v_416 = (v_198 ^ v_415);
	assign v_418 = (v_201 ^ v_417);
	assign v_420 = (v_205 ^ v_419);
	assign v_422 = (v_208 ^ v_421);
	assign v_424 = (v_212 ^ v_423);
	assign v_426 = (v_215 ^ v_425);
	assign v_430 = (v_221 ^ v_429);
	assign v_432 = (v_225 ^ v_431);
	assign v_434 = (v_228 ^ v_433);
	assign v_436 = (v_232 ^ v_435);
	assign v_438 = (v_235 ^ v_437);
	assign v_440 = (v_239 ^ v_439);
	assign v_442 = (v_242 ^ v_441);
	assign v_444 = (v_246 ^ v_443);
	assign v_446 = (v_249 ^ v_445);
	assign v_448 = (v_253 ^ v_447);
	assign v_450 = (v_256 ^ v_449);
	assign v_452 = (v_260 ^ v_451);
	assign v_454 = (v_263 ^ v_453);
	assign v_456 = (v_267 ^ v_455);
	assign v_458 = (v_270 ^ v_457);
	assign v_462 = (v_276 ^ v_461);
	assign v_464 = (v_280 ^ v_463);
	assign v_466 = (v_283 ^ v_465);
	assign v_468 = (v_287 ^ v_467);
	assign v_470 = (v_290 ^ v_469);
	assign v_472 = (v_294 ^ v_471);
	assign v_474 = (v_297 ^ v_473);
	assign v_476 = (v_301 ^ v_475);
	assign v_478 = (v_304 ^ v_477);
	assign v_480 = (v_308 ^ v_479);
	assign v_484 = (v_314 ^ v_483);
	assign v_486 = (v_317 ^ v_485);
	assign v_488 = (v_321 ^ v_487);
	assign v_490 = (v_324 ^ v_489);
	assign v_492 = (v_328 ^ v_491);
	assign v_494 = (v_331 ^ v_493);
	assign v_496 = (v_335 ^ v_495);
	assign v_498 = (v_338 ^ v_497);
	assign v_500 = (v_341 ^ v_499);
	assign v_128 = (v_505 & v_506);
	assign v_20 = (~v_21 & v_133);
	assign x_61 = (~v_21 | ~v_22);
	assign x_59 = (((v_21 | v_397)) | v_22);
	assign x_198 = (((v_53 | v_429)) | v_54);
	assign v_52 = (~v_53 & v_132);
	assign x_200 = (~v_53 | ~v_54);
	assign v_84 = (~v_85 & v_131);
	assign x_339 = (~v_85 | ~v_86);
	assign x_337 = (((v_85 | v_461)) | v_86);
	assign v_106 = (~v_107 & v_130);
	assign x_433 = (~v_107 | ~v_108);
	assign x_431 = (((v_107 | v_483)) | v_108);
	assign v_126 = (~v_127 & v_129);
	assign v_508 = (v_139 ^ v_507);
	assign x_530 = (((~v_137 | ~v_381)) | ~v_382);
	assign x_529 = (((~v_137 | v_381)) | v_382);
	assign x_527 = (((((v_137 | ~v_381)) | v_382)) | v_7);
	assign x_526 = (((((v_137 | v_381)) | ~v_382)) | v_7);
	assign x_525 = (((~v_136 | ~v_381)) | ~v_382);
	assign x_523 = (((v_136 | v_382)) | v_137);
	assign x_9 = (((~v_8 | ~v_383)) | ~v_384);
	assign x_8 = (((~v_8 | v_383)) | v_384);
	assign x_6 = (((((v_8 | ~v_383)) | v_384)) | v_9);
	assign x_5 = (((((v_8 | v_383)) | ~v_384)) | v_9);
	assign x_4 = (((~v_7 | ~v_383)) | ~v_384);
	assign x_2 = (((v_7 | v_384)) | v_8);
	assign x_18 = (((~v_10 | ~v_385)) | ~v_386);
	assign x_17 = (((~v_10 | v_385)) | v_386);
	assign x_15 = (((((v_10 | ~v_385)) | v_386)) | v_11);
	assign x_14 = (((((v_10 | v_385)) | ~v_386)) | v_11);
	assign x_13 = (((~v_9 | ~v_385)) | ~v_386);
	assign x_11 = (((v_9 | v_386)) | v_10);
	assign x_27 = (((~v_12 | ~v_387)) | ~v_388);
	assign x_26 = (((~v_12 | v_387)) | v_388);
	assign x_24 = (((((v_12 | ~v_387)) | v_388)) | v_13);
	assign x_23 = (((((v_12 | v_387)) | ~v_388)) | v_13);
	assign x_22 = (((~v_11 | ~v_387)) | ~v_388);
	assign x_20 = (((v_11 | v_388)) | v_12);
	assign x_33 = (((((v_14 | ~v_389)) | v_390)) | v_15);
	assign x_32 = (((((v_14 | v_389)) | ~v_390)) | v_15);
	assign x_36 = (((~v_14 | ~v_389)) | ~v_390);
	assign x_35 = (((~v_14 | v_389)) | v_390);
	assign x_31 = (((~v_13 | ~v_389)) | ~v_390);
	assign x_29 = (((v_13 | v_390)) | v_14);
	assign x_45 = (((~v_16 | ~v_391)) | ~v_392);
	assign x_44 = (((~v_16 | v_391)) | v_392);
	assign x_42 = (((((v_16 | ~v_391)) | v_392)) | v_17);
	assign x_41 = (((((v_16 | v_391)) | ~v_392)) | v_17);
	assign x_40 = (((~v_15 | ~v_391)) | ~v_392);
	assign x_38 = (((v_15 | v_392)) | v_16);
	assign x_54 = (((~v_18 | ~v_393)) | ~v_394);
	assign x_53 = (((~v_18 | v_393)) | v_394);
	assign x_51 = (((((v_18 | ~v_393)) | v_394)) | v_19);
	assign x_50 = (((((v_18 | v_393)) | ~v_394)) | v_19);
	assign x_49 = (((~v_17 | ~v_393)) | ~v_394);
	assign x_47 = (((v_17 | v_394)) | v_18);
	assign x_66 = (((~v_22 | v_397)) | v_398);
	assign x_67 = (((~v_22 | ~v_397)) | ~v_398);
	assign x_64 = (((((v_22 | ~v_397)) | v_398)) | v_23);
	assign x_63 = (((((v_22 | v_397)) | ~v_398)) | v_23);
	assign x_62 = (((~v_21 | ~v_397)) | ~v_398);
	assign x_60 = (((v_21 | v_398)) | v_22);
	assign x_76 = (((~v_24 | ~v_399)) | ~v_400);
	assign x_75 = (((~v_24 | v_399)) | v_400);
	assign x_73 = (((((v_24 | ~v_399)) | v_400)) | v_25);
	assign x_72 = (((((v_24 | v_399)) | ~v_400)) | v_25);
	assign x_71 = (((~v_23 | ~v_399)) | ~v_400);
	assign x_69 = (((v_23 | v_400)) | v_24);
	assign x_85 = (((~v_26 | ~v_401)) | ~v_402);
	assign x_84 = (((~v_26 | v_401)) | v_402);
	assign x_82 = (((((v_26 | ~v_401)) | v_402)) | v_27);
	assign x_81 = (((((v_26 | v_401)) | ~v_402)) | v_27);
	assign x_80 = (((~v_25 | ~v_401)) | ~v_402);
	assign x_78 = (((v_25 | v_402)) | v_26);
	assign x_94 = (((~v_28 | ~v_403)) | ~v_404);
	assign x_93 = (((~v_28 | v_403)) | v_404);
	assign x_91 = (((((v_28 | ~v_403)) | v_404)) | v_29);
	assign x_90 = (((((v_28 | v_403)) | ~v_404)) | v_29);
	assign x_89 = (((~v_27 | ~v_403)) | ~v_404);
	assign x_87 = (((v_27 | v_404)) | v_28);
	assign x_99 = (((((v_30 | v_405)) | ~v_406)) | v_31);
	assign x_98 = (((~v_29 | ~v_405)) | ~v_406);
	assign x_103 = (((~v_30 | ~v_405)) | ~v_406);
	assign x_102 = (((~v_30 | v_405)) | v_406);
	assign x_100 = (((((v_30 | ~v_405)) | v_406)) | v_31);
	assign x_96 = (((v_29 | v_406)) | v_30);
	assign x_112 = (((~v_32 | ~v_407)) | ~v_408);
	assign x_111 = (((~v_32 | v_407)) | v_408);
	assign x_109 = (((((v_32 | ~v_407)) | v_408)) | v_33);
	assign x_108 = (((((v_32 | v_407)) | ~v_408)) | v_33);
	assign x_107 = (((~v_31 | ~v_407)) | ~v_408);
	assign x_105 = (((v_31 | v_408)) | v_32);
	assign x_121 = (((~v_34 | ~v_409)) | ~v_410);
	assign x_120 = (((~v_34 | v_409)) | v_410);
	assign x_118 = (((((v_34 | ~v_409)) | v_410)) | v_35);
	assign x_117 = (((((v_34 | v_409)) | ~v_410)) | v_35);
	assign x_116 = (((~v_33 | ~v_409)) | ~v_410);
	assign x_114 = (((v_33 | v_410)) | v_34);
	assign x_130 = (((~v_36 | ~v_411)) | ~v_412);
	assign x_129 = (((~v_36 | v_411)) | v_412);
	assign x_127 = (((((v_36 | ~v_411)) | v_412)) | v_37);
	assign x_126 = (((((v_36 | v_411)) | ~v_412)) | v_37);
	assign x_125 = (((~v_35 | ~v_411)) | ~v_412);
	assign x_123 = (((v_35 | v_412)) | v_36);
	assign x_132 = (((v_37 | v_414)) | v_38);
	assign x_139 = (((~v_38 | ~v_413)) | ~v_414);
	assign x_138 = (((~v_38 | v_413)) | v_414);
	assign x_136 = (((((v_38 | ~v_413)) | v_414)) | v_39);
	assign x_135 = (((((v_38 | v_413)) | ~v_414)) | v_39);
	assign x_134 = (((~v_37 | ~v_413)) | ~v_414);
	assign x_148 = (((~v_40 | ~v_415)) | ~v_416);
	assign x_147 = (((~v_40 | v_415)) | v_416);
	assign x_145 = (((((v_40 | ~v_415)) | v_416)) | v_41);
	assign x_144 = (((((v_40 | v_415)) | ~v_416)) | v_41);
	assign x_143 = (((~v_39 | ~v_415)) | ~v_416);
	assign x_141 = (((v_39 | v_416)) | v_40);
	assign x_157 = (((~v_42 | ~v_417)) | ~v_418);
	assign x_156 = (((~v_42 | v_417)) | v_418);
	assign x_154 = (((((v_42 | ~v_417)) | v_418)) | v_43);
	assign x_153 = (((((v_42 | v_417)) | ~v_418)) | v_43);
	assign x_152 = (((~v_41 | ~v_417)) | ~v_418);
	assign x_150 = (((v_41 | v_418)) | v_42);
	assign x_165 = (((~v_44 | v_419)) | v_420);
	assign x_166 = (((~v_44 | ~v_419)) | ~v_420);
	assign x_163 = (((((v_44 | ~v_419)) | v_420)) | v_45);
	assign x_162 = (((((v_44 | v_419)) | ~v_420)) | v_45);
	assign x_161 = (((~v_43 | ~v_419)) | ~v_420);
	assign x_159 = (((v_43 | v_420)) | v_44);
	assign x_175 = (((~v_46 | ~v_421)) | ~v_422);
	assign x_174 = (((~v_46 | v_421)) | v_422);
	assign x_172 = (((((v_46 | ~v_421)) | v_422)) | v_47);
	assign x_171 = (((((v_46 | v_421)) | ~v_422)) | v_47);
	assign x_170 = (((~v_45 | ~v_421)) | ~v_422);
	assign x_168 = (((v_45 | v_422)) | v_46);
	assign x_184 = (((~v_48 | ~v_423)) | ~v_424);
	assign x_183 = (((~v_48 | v_423)) | v_424);
	assign x_181 = (((((v_48 | ~v_423)) | v_424)) | v_49);
	assign x_180 = (((((v_48 | v_423)) | ~v_424)) | v_49);
	assign x_179 = (((~v_47 | ~v_423)) | ~v_424);
	assign x_177 = (((v_47 | v_424)) | v_48);
	assign x_193 = (((~v_50 | ~v_425)) | ~v_426);
	assign x_192 = (((~v_50 | v_425)) | v_426);
	assign x_190 = (((((v_50 | ~v_425)) | v_426)) | v_51);
	assign x_189 = (((((v_50 | v_425)) | ~v_426)) | v_51);
	assign x_188 = (((~v_49 | ~v_425)) | ~v_426);
	assign x_186 = (((v_49 | v_426)) | v_50);
	assign x_206 = (((~v_54 | ~v_429)) | ~v_430);
	assign x_205 = (((~v_54 | v_429)) | v_430);
	assign x_203 = (((((v_54 | ~v_429)) | v_430)) | v_55);
	assign x_202 = (((((v_54 | v_429)) | ~v_430)) | v_55);
	assign x_201 = (((~v_53 | ~v_429)) | ~v_430);
	assign x_199 = (((v_53 | v_430)) | v_54);
	assign x_215 = (((~v_56 | ~v_431)) | ~v_432);
	assign x_214 = (((~v_56 | v_431)) | v_432);
	assign x_212 = (((((v_56 | ~v_431)) | v_432)) | v_57);
	assign x_211 = (((((v_56 | v_431)) | ~v_432)) | v_57);
	assign x_210 = (((~v_55 | ~v_431)) | ~v_432);
	assign x_208 = (((v_55 | v_432)) | v_56);
	assign x_224 = (((~v_58 | ~v_433)) | ~v_434);
	assign x_223 = (((~v_58 | v_433)) | v_434);
	assign x_221 = (((((v_58 | ~v_433)) | v_434)) | v_59);
	assign x_220 = (((((v_58 | v_433)) | ~v_434)) | v_59);
	assign x_219 = (((~v_57 | ~v_433)) | ~v_434);
	assign x_217 = (((v_57 | v_434)) | v_58);
	assign x_230 = (((((v_60 | ~v_435)) | v_436)) | v_61);
	assign x_233 = (((~v_60 | ~v_435)) | ~v_436);
	assign x_232 = (((~v_60 | v_435)) | v_436);
	assign x_229 = (((((v_60 | v_435)) | ~v_436)) | v_61);
	assign x_228 = (((~v_59 | ~v_435)) | ~v_436);
	assign x_226 = (((v_59 | v_436)) | v_60);
	assign x_242 = (((~v_62 | ~v_437)) | ~v_438);
	assign x_241 = (((~v_62 | v_437)) | v_438);
	assign x_239 = (((((v_62 | ~v_437)) | v_438)) | v_63);
	assign x_238 = (((((v_62 | v_437)) | ~v_438)) | v_63);
	assign x_237 = (((~v_61 | ~v_437)) | ~v_438);
	assign x_235 = (((v_61 | v_438)) | v_62);
	assign x_248 = (((((v_64 | ~v_439)) | v_440)) | v_65);
	assign x_247 = (((((v_64 | v_439)) | ~v_440)) | v_65);
	assign x_251 = (((~v_64 | ~v_439)) | ~v_440);
	assign x_250 = (((~v_64 | v_439)) | v_440);
	assign x_246 = (((~v_63 | ~v_439)) | ~v_440);
	assign x_244 = (((v_63 | v_440)) | v_64);
	assign x_260 = (((~v_66 | ~v_441)) | ~v_442);
	assign x_259 = (((~v_66 | v_441)) | v_442);
	assign x_257 = (((((v_66 | ~v_441)) | v_442)) | v_67);
	assign x_256 = (((((v_66 | v_441)) | ~v_442)) | v_67);
	assign x_255 = (((~v_65 | ~v_441)) | ~v_442);
	assign x_253 = (((v_65 | v_442)) | v_66);
	assign x_265 = (((((v_68 | v_443)) | ~v_444)) | v_69);
	assign x_264 = (((~v_67 | ~v_443)) | ~v_444);
	assign x_269 = (((~v_68 | ~v_443)) | ~v_444);
	assign x_268 = (((~v_68 | v_443)) | v_444);
	assign x_266 = (((((v_68 | ~v_443)) | v_444)) | v_69);
	assign x_262 = (((v_67 | v_444)) | v_68);
	assign x_278 = (((~v_70 | ~v_445)) | ~v_446);
	assign x_277 = (((~v_70 | v_445)) | v_446);
	assign x_275 = (((((v_70 | ~v_445)) | v_446)) | v_71);
	assign x_274 = (((((v_70 | v_445)) | ~v_446)) | v_71);
	assign x_273 = (((~v_69 | ~v_445)) | ~v_446);
	assign x_271 = (((v_69 | v_446)) | v_70);
	assign x_287 = (((~v_72 | ~v_447)) | ~v_448);
	assign x_286 = (((~v_72 | v_447)) | v_448);
	assign x_284 = (((((v_72 | ~v_447)) | v_448)) | v_73);
	assign x_283 = (((((v_72 | v_447)) | ~v_448)) | v_73);
	assign x_282 = (((~v_71 | ~v_447)) | ~v_448);
	assign x_280 = (((v_71 | v_448)) | v_72);
	assign x_296 = (((~v_74 | ~v_449)) | ~v_450);
	assign x_295 = (((~v_74 | v_449)) | v_450);
	assign x_293 = (((((v_74 | ~v_449)) | v_450)) | v_75);
	assign x_292 = (((((v_74 | v_449)) | ~v_450)) | v_75);
	assign x_291 = (((~v_73 | ~v_449)) | ~v_450);
	assign x_289 = (((v_73 | v_450)) | v_74);
	assign x_298 = (((v_75 | v_452)) | v_76);
	assign x_305 = (((~v_76 | ~v_451)) | ~v_452);
	assign x_304 = (((~v_76 | v_451)) | v_452);
	assign x_302 = (((((v_76 | ~v_451)) | v_452)) | v_77);
	assign x_301 = (((((v_76 | v_451)) | ~v_452)) | v_77);
	assign x_300 = (((~v_75 | ~v_451)) | ~v_452);
	assign x_314 = (((~v_78 | ~v_453)) | ~v_454);
	assign x_313 = (((~v_78 | v_453)) | v_454);
	assign x_311 = (((((v_78 | ~v_453)) | v_454)) | v_79);
	assign x_310 = (((((v_78 | v_453)) | ~v_454)) | v_79);
	assign x_309 = (((~v_77 | ~v_453)) | ~v_454);
	assign x_307 = (((v_77 | v_454)) | v_78);
	assign x_323 = (((~v_80 | ~v_455)) | ~v_456);
	assign x_322 = (((~v_80 | v_455)) | v_456);
	assign x_320 = (((((v_80 | ~v_455)) | v_456)) | v_81);
	assign x_319 = (((((v_80 | v_455)) | ~v_456)) | v_81);
	assign x_318 = (((~v_79 | ~v_455)) | ~v_456);
	assign x_316 = (((v_79 | v_456)) | v_80);
	assign x_331 = (((~v_82 | v_457)) | v_458);
	assign x_332 = (((~v_82 | ~v_457)) | ~v_458);
	assign x_329 = (((((v_82 | ~v_457)) | v_458)) | v_83);
	assign x_328 = (((((v_82 | v_457)) | ~v_458)) | v_83);
	assign x_327 = (((~v_81 | ~v_457)) | ~v_458);
	assign x_325 = (((v_81 | v_458)) | v_82);
	assign x_345 = (((~v_86 | ~v_461)) | ~v_462);
	assign x_344 = (((~v_86 | v_461)) | v_462);
	assign x_342 = (((((v_86 | ~v_461)) | v_462)) | v_87);
	assign x_341 = (((((v_86 | v_461)) | ~v_462)) | v_87);
	assign x_340 = (((~v_85 | ~v_461)) | ~v_462);
	assign x_338 = (((v_85 | v_462)) | v_86);
	assign x_354 = (((~v_88 | ~v_463)) | ~v_464);
	assign x_353 = (((~v_88 | v_463)) | v_464);
	assign x_351 = (((((v_88 | ~v_463)) | v_464)) | v_89);
	assign x_350 = (((((v_88 | v_463)) | ~v_464)) | v_89);
	assign x_349 = (((~v_87 | ~v_463)) | ~v_464);
	assign x_347 = (((v_87 | v_464)) | v_88);
	assign x_363 = (((~v_90 | ~v_465)) | ~v_466);
	assign x_362 = (((~v_90 | v_465)) | v_466);
	assign x_360 = (((((v_90 | ~v_465)) | v_466)) | v_91);
	assign x_359 = (((((v_90 | v_465)) | ~v_466)) | v_91);
	assign x_358 = (((~v_89 | ~v_465)) | ~v_466);
	assign x_356 = (((v_89 | v_466)) | v_90);
	assign x_372 = (((~v_92 | ~v_467)) | ~v_468);
	assign x_371 = (((~v_92 | v_467)) | v_468);
	assign x_369 = (((((v_92 | ~v_467)) | v_468)) | v_93);
	assign x_368 = (((((v_92 | v_467)) | ~v_468)) | v_93);
	assign x_367 = (((~v_91 | ~v_467)) | ~v_468);
	assign x_365 = (((v_91 | v_468)) | v_92);
	assign x_381 = (((~v_94 | ~v_469)) | ~v_470);
	assign x_380 = (((~v_94 | v_469)) | v_470);
	assign x_378 = (((((v_94 | ~v_469)) | v_470)) | v_95);
	assign x_377 = (((((v_94 | v_469)) | ~v_470)) | v_95);
	assign x_376 = (((~v_93 | ~v_469)) | ~v_470);
	assign x_374 = (((v_93 | v_470)) | v_94);
	assign x_390 = (((~v_96 | ~v_471)) | ~v_472);
	assign x_389 = (((~v_96 | v_471)) | v_472);
	assign x_387 = (((((v_96 | ~v_471)) | v_472)) | v_97);
	assign x_386 = (((((v_96 | v_471)) | ~v_472)) | v_97);
	assign x_385 = (((~v_95 | ~v_471)) | ~v_472);
	assign x_383 = (((v_95 | v_472)) | v_96);
	assign x_396 = (((((v_98 | ~v_473)) | v_474)) | v_99);
	assign x_399 = (((~v_98 | ~v_473)) | ~v_474);
	assign x_398 = (((~v_98 | v_473)) | v_474);
	assign x_395 = (((((v_98 | v_473)) | ~v_474)) | v_99);
	assign x_394 = (((~v_97 | ~v_473)) | ~v_474);
	assign x_392 = (((v_97 | v_474)) | v_98);
	assign x_408 = (((~v_100 | ~v_475)) | ~v_476);
	assign x_407 = (((~v_100 | v_475)) | v_476);
	assign x_405 = (((((v_100 | ~v_475)) | v_476)) | v_101);
	assign x_404 = (((((v_100 | v_475)) | ~v_476)) | v_101);
	assign x_403 = (((~v_99 | ~v_475)) | ~v_476);
	assign x_401 = (((v_99 | v_476)) | v_100);
	assign x_417 = (((~v_102 | ~v_477)) | ~v_478);
	assign x_416 = (((~v_102 | v_477)) | v_478);
	assign x_414 = (((((v_102 | ~v_477)) | v_478)) | v_103);
	assign x_413 = (((((v_102 | v_477)) | ~v_478)) | v_103);
	assign x_412 = (((~v_101 | ~v_477)) | ~v_478);
	assign x_410 = (((v_101 | v_478)) | v_102);
	assign x_426 = (((~v_104 | ~v_479)) | ~v_480);
	assign x_425 = (((~v_104 | v_479)) | v_480);
	assign x_423 = (((((v_104 | ~v_479)) | v_480)) | v_105);
	assign x_422 = (((((v_104 | v_479)) | ~v_480)) | v_105);
	assign x_421 = (((~v_103 | ~v_479)) | ~v_480);
	assign x_419 = (((v_103 | v_480)) | v_104);
	assign x_439 = (((~v_108 | ~v_483)) | ~v_484);
	assign x_438 = (((~v_108 | v_483)) | v_484);
	assign x_436 = (((((v_108 | ~v_483)) | v_484)) | v_109);
	assign x_435 = (((((v_108 | v_483)) | ~v_484)) | v_109);
	assign x_434 = (((~v_107 | ~v_483)) | ~v_484);
	assign x_432 = (((v_107 | v_484)) | v_108);
	assign x_448 = (((~v_110 | ~v_485)) | ~v_486);
	assign x_447 = (((~v_110 | v_485)) | v_486);
	assign x_445 = (((((v_110 | ~v_485)) | v_486)) | v_111);
	assign x_444 = (((((v_110 | v_485)) | ~v_486)) | v_111);
	assign x_443 = (((~v_109 | ~v_485)) | ~v_486);
	assign x_441 = (((v_109 | v_486)) | v_110);
	assign x_457 = (((~v_112 | ~v_487)) | ~v_488);
	assign x_456 = (((~v_112 | v_487)) | v_488);
	assign x_454 = (((((v_112 | ~v_487)) | v_488)) | v_113);
	assign x_453 = (((((v_112 | v_487)) | ~v_488)) | v_113);
	assign x_452 = (((~v_111 | ~v_487)) | ~v_488);
	assign x_450 = (((v_111 | v_488)) | v_112);
	assign x_463 = (((((v_114 | ~v_489)) | v_490)) | v_115);
	assign x_462 = (((((v_114 | v_489)) | ~v_490)) | v_115);
	assign x_466 = (((~v_114 | ~v_489)) | ~v_490);
	assign x_465 = (((~v_114 | v_489)) | v_490);
	assign x_461 = (((~v_113 | ~v_489)) | ~v_490);
	assign x_459 = (((v_113 | v_490)) | v_114);
	assign x_475 = (((~v_116 | ~v_491)) | ~v_492);
	assign x_474 = (((~v_116 | v_491)) | v_492);
	assign x_472 = (((((v_116 | ~v_491)) | v_492)) | v_117);
	assign x_471 = (((((v_116 | v_491)) | ~v_492)) | v_117);
	assign x_470 = (((~v_115 | ~v_491)) | ~v_492);
	assign x_468 = (((v_115 | v_492)) | v_116);
	assign x_484 = (((~v_118 | ~v_493)) | ~v_494);
	assign x_483 = (((~v_118 | v_493)) | v_494);
	assign x_481 = (((((v_118 | ~v_493)) | v_494)) | v_119);
	assign x_480 = (((((v_118 | v_493)) | ~v_494)) | v_119);
	assign x_479 = (((~v_117 | ~v_493)) | ~v_494);
	assign x_477 = (((v_117 | v_494)) | v_118);
	assign x_493 = (((~v_120 | ~v_495)) | ~v_496);
	assign x_492 = (((~v_120 | v_495)) | v_496);
	assign x_490 = (((((v_120 | ~v_495)) | v_496)) | v_121);
	assign x_489 = (((((v_120 | v_495)) | ~v_496)) | v_121);
	assign x_488 = (((~v_119 | ~v_495)) | ~v_496);
	assign x_486 = (((v_119 | v_496)) | v_120);
	assign x_495 = (((v_121 | v_498)) | v_122);
	assign x_502 = (((~v_122 | ~v_497)) | ~v_498);
	assign x_501 = (((~v_122 | v_497)) | v_498);
	assign x_499 = (((((v_122 | ~v_497)) | v_498)) | v_123);
	assign x_498 = (((((v_122 | v_497)) | ~v_498)) | v_123);
	assign x_497 = (((~v_121 | ~v_497)) | ~v_498);
	assign x_511 = (((~v_124 | ~v_499)) | ~v_500);
	assign x_510 = (((~v_124 | v_499)) | v_500);
	assign x_508 = (((((v_124 | ~v_499)) | v_500)) | v_125);
	assign x_507 = (((((v_124 | v_499)) | ~v_500)) | v_125);
	assign x_506 = (((~v_123 | ~v_499)) | ~v_500);
	assign x_504 = (((v_123 | v_500)) | v_124);
	assign v_347 = (v_346 ^ v_128);
	assign x_521 = (((~v_127 | ~v_503)) | ~v_128);
	assign x_516 = (((v_127 | v_503)) | v_128);
	assign x_57 = (~v_19 | ~v_20);
	assign x_56 = (((v_19 | v_396)) | v_20);
	assign x_55 = (((v_19 | v_395)) | v_20);
	assign x_585 = (x_58 & x_59);
	assign x_720 = (x_197 & x_198);
	assign x_196 = (~v_51 | ~v_52);
	assign x_195 = (((v_51 | v_428)) | v_52);
	assign x_194 = (((v_51 | v_427)) | v_52);
	assign x_335 = (~v_83 | ~v_84);
	assign x_334 = (((v_83 | v_460)) | v_84);
	assign x_333 = (((v_83 | v_459)) | v_84);
	assign x_863 = (x_336 & x_337);
	assign x_429 = (~v_105 | ~v_106);
	assign x_428 = (((v_105 | v_482)) | v_106);
	assign x_427 = (((v_105 | v_481)) | v_106);
	assign x_513 = (((v_125 | v_502)) | v_126);
	assign x_512 = (((v_125 | v_501)) | v_126);
	assign x_514 = (~v_125 | ~v_126);
	assign x_1050 = (x_529 & x_530);
	assign x_1049 = (x_526 & x_527);
	assign x_1047 = (x_524 & x_525);
	assign x_1046 = (x_522 & x_523);
	assign x_538 = (x_9 & x_10);
	assign x_535 = (x_7 & x_8);
	assign x_534 = (x_5 & x_6);
	assign x_532 = (x_3 & x_4);
	assign x_531 = (x_1 & x_2);
	assign x_546 = (x_17 & x_18);
	assign x_542 = (x_15 & x_16);
	assign x_541 = (x_13 & x_14);
	assign x_539 = (x_11 & x_12);
	assign x_554 = (x_27 & x_28);
	assign x_553 = (x_25 & x_26);
	assign x_550 = (x_23 & x_24);
	assign x_549 = (x_21 & x_22);
	assign x_547 = (x_19 & x_20);
	assign x_557 = (x_32 & x_33);
	assign x_564 = (x_36 & x_37);
	assign x_563 = (x_34 & x_35);
	assign x_556 = (x_29 & x_30);
	assign x_571 = (x_44 & x_45);
	assign x_570 = (x_42 & x_43);
	assign x_567 = (x_40 & x_41);
	assign x_566 = (x_38 & x_39);
	assign x_579 = (x_52 & x_53);
	assign x_578 = (x_50 & x_51);
	assign x_574 = (x_48 & x_49);
	assign x_573 = (x_46 & x_47);
	assign x_589 = (x_65 & x_66);
	assign x_596 = (x_67 & x_68);
	assign x_588 = (x_62 & x_63);
	assign x_586 = (x_60 & x_61);
	assign x_603 = (x_75 & x_76);
	assign x_600 = (x_73 & x_74);
	assign x_599 = (x_71 & x_72);
	assign x_597 = (x_69 & x_70);
	assign x_612 = (x_85 & x_86);
	assign x_611 = (x_83 & x_84);
	assign x_607 = (x_81 & x_82);
	assign x_606 = (x_79 & x_80);
	assign x_604 = (x_77 & x_78);
	assign x_619 = (x_93 & x_94);
	assign x_618 = (x_91 & x_92);
	assign x_615 = (x_89 & x_90);
	assign x_614 = (x_87 & x_88);
	assign x_622 = (x_98 & x_99);
	assign x_629 = (x_102 & x_103);
	assign x_628 = (x_100 & x_101);
	assign x_621 = (x_95 & x_96);
	assign x_638 = (x_112 & x_113);
	assign x_636 = (x_110 & x_111);
	assign x_635 = (x_108 & x_109);
	assign x_632 = (x_106 & x_107);
	assign x_631 = (x_104 & x_105);
	assign x_646 = (x_120 & x_121);
	assign x_644 = (x_118 & x_119);
	assign x_643 = (x_116 & x_117);
	assign x_639 = (x_114 & x_115);
	assign x_653 = (x_128 & x_129);
	assign x_651 = (x_126 & x_127);
	assign x_650 = (x_124 & x_125);
	assign x_647 = (x_122 & x_123);
	assign x_654 = (x_131 & x_132);
	assign x_666 = (x_139 & x_140);
	assign x_665 = (x_137 & x_138);
	assign x_663 = (x_135 & x_136);
	assign x_662 = (x_133 & x_134);
	assign x_673 = (x_147 & x_148);
	assign x_672 = (x_145 & x_146);
	assign x_670 = (x_143 & x_144);
	assign x_669 = (x_141 & x_142);
	assign x_684 = (x_157 & x_158);
	assign x_681 = (x_155 & x_156);
	assign x_680 = (x_153 & x_154);
	assign x_678 = (x_151 & x_152);
	assign x_677 = (x_149 & x_150);
	assign x_688 = (x_164 & x_165);
	assign x_694 = (x_166 & x_167);
	assign x_687 = (x_161 & x_162);
	assign x_685 = (x_159 & x_160);
	assign x_701 = (x_174 & x_175);
	assign x_698 = (x_172 & x_173);
	assign x_697 = (x_170 & x_171);
	assign x_695 = (x_168 & x_169);
	assign x_710 = (x_184 & x_185);
	assign x_709 = (x_182 & x_183);
	assign x_705 = (x_180 & x_181);
	assign x_704 = (x_178 & x_179);
	assign x_702 = (x_176 & x_177);
	assign x_717 = (x_192 & x_193);
	assign x_716 = (x_190 & x_191);
	assign x_713 = (x_188 & x_189);
	assign x_712 = (x_186 & x_187);
	assign x_731 = (x_205 & x_206);
	assign x_730 = (x_203 & x_204);
	assign x_728 = (x_201 & x_202);
	assign x_727 = (x_199 & x_200);
	assign x_742 = (x_215 & x_216);
	assign x_738 = (x_213 & x_214);
	assign x_737 = (x_211 & x_212);
	assign x_735 = (x_209 & x_210);
	assign x_734 = (x_207 & x_208);
	assign x_749 = (x_223 & x_224);
	assign x_746 = (x_221 & x_222);
	assign x_745 = (x_219 & x_220);
	assign x_743 = (x_217 & x_218);
	assign x_753 = (x_230 & x_231);
	assign x_759 = (x_232 & x_233);
	assign x_752 = (x_227 & x_228);
	assign x_750 = (x_225 & x_226);
	assign x_767 = (x_242 & x_243);
	assign x_766 = (x_240 & x_241);
	assign x_763 = (x_238 & x_239);
	assign x_762 = (x_236 & x_237);
	assign x_760 = (x_234 & x_235);
	assign x_770 = (x_247 & x_248);
	assign x_776 = (x_251 & x_252);
	assign x_775 = (x_249 & x_250);
	assign x_769 = (x_244 & x_245);
	assign x_783 = (x_259 & x_260);
	assign x_782 = (x_257 & x_258);
	assign x_779 = (x_255 & x_256);
	assign x_778 = (x_253 & x_254);
	assign x_786 = (x_264 & x_265);
	assign x_796 = (x_268 & x_269);
	assign x_795 = (x_266 & x_267);
	assign x_785 = (x_261 & x_262);
	assign x_805 = (x_278 & x_279);
	assign x_803 = (x_276 & x_277);
	assign x_802 = (x_274 & x_275);
	assign x_799 = (x_272 & x_273);
	assign x_798 = (x_270 & x_271);
	assign x_813 = (x_286 & x_287);
	assign x_811 = (x_284 & x_285);
	assign x_810 = (x_282 & x_283);
	assign x_806 = (x_280 & x_281);
	assign x_820 = (x_294 & x_295);
	assign x_818 = (x_292 & x_293);
	assign x_817 = (x_290 & x_291);
	assign x_814 = (x_288 & x_289);
	assign x_821 = (x_297 & x_298);
	assign x_831 = (x_305 & x_306);
	assign x_830 = (x_303 & x_304);
	assign x_828 = (x_301 & x_302);
	assign x_827 = (x_299 & x_300);
	assign x_838 = (x_313 & x_314);
	assign x_837 = (x_311 & x_312);
	assign x_835 = (x_309 & x_310);
	assign x_834 = (x_307 & x_308);
	assign x_849 = (x_323 & x_324);
	assign x_846 = (x_321 & x_322);
	assign x_845 = (x_319 & x_320);
	assign x_843 = (x_317 & x_318);
	assign x_842 = (x_315 & x_316);
	assign x_853 = (x_330 & x_331);
	assign x_852 = (x_327 & x_328);
	assign x_850 = (x_325 & x_326);
	assign x_870 = (x_344 & x_345);
	assign x_868 = (x_342 & x_343);
	assign x_867 = (x_340 & x_341);
	assign x_864 = (x_338 & x_339);
	assign x_879 = (x_354 & x_355);
	assign x_878 = (x_352 & x_353);
	assign x_876 = (x_350 & x_351);
	assign x_875 = (x_348 & x_349);
	assign x_871 = (x_346 & x_347);
	assign x_886 = (x_363 & x_364);
	assign x_885 = (x_360 & x_361);
	assign x_883 = (x_358 & x_359);
	assign x_882 = (x_356 & x_357);
	assign x_896 = (x_371 & x_372);
	assign x_895 = (x_369 & x_370);
	assign x_893 = (x_367 & x_368);
	assign x_892 = (x_365 & x_366);
	assign x_907 = (x_381 & x_382);
	assign x_903 = (x_379 & x_380);
	assign x_902 = (x_377 & x_378);
	assign x_900 = (x_375 & x_376);
	assign x_899 = (x_373 & x_374);
	assign x_914 = (x_389 & x_390);
	assign x_911 = (x_387 & x_388);
	assign x_910 = (x_385 & x_386);
	assign x_908 = (x_383 & x_384);
	assign x_918 = (x_396 & x_397);
	assign x_926 = (x_398 & x_399);
	assign x_917 = (x_393 & x_394);
	assign x_915 = (x_391 & x_392);
	assign x_934 = (x_408 & x_409);
	assign x_933 = (x_406 & x_407);
	assign x_930 = (x_404 & x_405);
	assign x_929 = (x_402 & x_403);
	assign x_927 = (x_400 & x_401);
	assign x_942 = (x_416 & x_417);
	assign x_941 = (x_414 & x_415);
	assign x_937 = (x_412 & x_413);
	assign x_936 = (x_410 & x_411);
	assign x_949 = (x_424 & x_425);
	assign x_948 = (x_422 & x_423);
	assign x_945 = (x_420 & x_421);
	assign x_944 = (x_418 & x_419);
	assign x_965 = (x_439 & x_440);
	assign x_962 = (x_437 & x_438);
	assign x_961 = (x_435 & x_436);
	assign x_959 = (x_433 & x_434);
	assign x_958 = (x_431 & x_432);
	assign x_973 = (x_447 & x_448);
	assign x_969 = (x_445 & x_446);
	assign x_968 = (x_443 & x_444);
	assign x_966 = (x_441 & x_442);
	assign x_981 = (x_457 & x_458);
	assign x_980 = (x_455 & x_456);
	assign x_977 = (x_453 & x_454);
	assign x_976 = (x_451 & x_452);
	assign x_974 = (x_449 & x_450);
	assign x_984 = (x_462 & x_463);
	assign x_992 = (x_466 & x_467);
	assign x_991 = (x_464 & x_465);
	assign x_983 = (x_459 & x_460);
	assign x_999 = (x_474 & x_475);
	assign x_998 = (x_472 & x_473);
	assign x_995 = (x_470 & x_471);
	assign x_994 = (x_468 & x_469);
	assign x_1009 = (x_484 & x_485);
	assign x_1007 = (x_482 & x_483);
	assign x_1006 = (x_480 & x_481);
	assign x_1002 = (x_478 & x_479);
	assign x_1001 = (x_476 & x_477);
	assign x_1016 = (x_492 & x_493);
	assign x_1014 = (x_490 & x_491);
	assign x_1013 = (x_488 & x_489);
	assign x_1010 = (x_486 & x_487);
	assign x_1017 = (x_495 & x_496);
	assign x_1026 = (x_501 & x_502);
	assign x_1024 = (x_499 & x_500);
	assign x_1023 = (x_497 & x_498);
	assign x_1033 = (x_509 & x_510);
	assign x_1031 = (x_507 & x_508);
	assign x_1030 = (x_505 & x_506);
	assign x_1027 = (x_503 & x_504);
	assign v_504 = (v_347 ^ v_503);
	assign x_582 = (x_56 & x_57);
	assign x_581 = (x_54 & x_55);
	assign x_721 = (x_196 & x_720);
	assign x_719 = (x_194 & x_195);
	assign x_861 = (x_334 & x_335);
	assign x_860 = (x_332 & x_333);
	assign x_952 = (x_429 & x_430);
	assign x_951 = (x_426 & x_427);
	assign x_1034 = (x_512 & x_513);
	assign x_1039 = (x_514 & x_515);
	assign x_1051 = (x_528 & x_1050);
	assign x_1048 = (x_1046 & x_1047);
	assign x_536 = (x_534 & x_535);
	assign x_533 = (x_531 & x_532);
	assign x_543 = (x_541 & x_542);
	assign x_540 = (x_538 & x_539);
	assign x_555 = (x_553 & x_554);
	assign x_551 = (x_549 & x_550);
	assign x_548 = (x_546 & x_547);
	assign x_558 = (x_31 & x_557);
	assign x_565 = (x_563 & x_564);
	assign x_572 = (x_570 & x_571);
	assign x_568 = (x_566 & x_567);
	assign x_580 = (x_578 & x_579);
	assign x_575 = (x_573 & x_574);
	assign x_590 = (x_64 & x_589);
	assign x_587 = (x_585 & x_586);
	assign x_601 = (x_599 & x_600);
	assign x_598 = (x_596 & x_597);
	assign x_613 = (x_611 & x_612);
	assign x_608 = (x_606 & x_607);
	assign x_605 = (x_603 & x_604);
	assign x_620 = (x_618 & x_619);
	assign x_616 = (x_614 & x_615);
	assign x_623 = (x_97 & x_622);
	assign x_630 = (x_628 & x_629);
	assign x_637 = (x_635 & x_636);
	assign x_633 = (x_631 & x_632);
	assign x_645 = (x_643 & x_644);
	assign x_640 = (x_638 & x_639);
	assign x_652 = (x_650 & x_651);
	assign x_648 = (x_646 & x_647);
	assign x_655 = (x_130 & x_654);
	assign x_667 = (x_665 & x_666);
	assign x_664 = (x_662 & x_663);
	assign x_674 = (x_672 & x_673);
	assign x_671 = (x_669 & x_670);
	assign x_682 = (x_680 & x_681);
	assign x_679 = (x_677 & x_678);
	assign x_689 = (x_163 & x_688);
	assign x_686 = (x_684 & x_685);
	assign x_699 = (x_697 & x_698);
	assign x_696 = (x_694 & x_695);
	assign x_711 = (x_709 & x_710);
	assign x_706 = (x_704 & x_705);
	assign x_703 = (x_701 & x_702);
	assign x_718 = (x_716 & x_717);
	assign x_714 = (x_712 & x_713);
	assign x_732 = (x_730 & x_731);
	assign x_729 = (x_727 & x_728);
	assign x_739 = (x_737 & x_738);
	assign x_736 = (x_734 & x_735);
	assign x_747 = (x_745 & x_746);
	assign x_744 = (x_742 & x_743);
	assign x_754 = (x_229 & x_753);
	assign x_751 = (x_749 & x_750);
	assign x_768 = (x_766 & x_767);
	assign x_764 = (x_762 & x_763);
	assign x_761 = (x_759 & x_760);
	assign x_771 = (x_246 & x_770);
	assign x_777 = (x_775 & x_776);
	assign x_784 = (x_782 & x_783);
	assign x_780 = (x_778 & x_779);
	assign x_787 = (x_263 & x_786);
	assign x_797 = (x_795 & x_796);
	assign x_804 = (x_802 & x_803);
	assign x_800 = (x_798 & x_799);
	assign x_812 = (x_810 & x_811);
	assign x_807 = (x_805 & x_806);
	assign x_819 = (x_817 & x_818);
	assign x_815 = (x_813 & x_814);
	assign x_822 = (x_296 & x_821);
	assign x_832 = (x_830 & x_831);
	assign x_829 = (x_827 & x_828);
	assign x_839 = (x_837 & x_838);
	assign x_836 = (x_834 & x_835);
	assign x_847 = (x_845 & x_846);
	assign x_844 = (x_842 & x_843);
	assign x_854 = (x_329 & x_853);
	assign x_851 = (x_849 & x_850);
	assign x_869 = (x_867 & x_868);
	assign x_865 = (x_863 & x_864);
	assign x_880 = (x_878 & x_879);
	assign x_877 = (x_875 & x_876);
	assign x_872 = (x_870 & x_871);
	assign x_887 = (x_362 & x_886);
	assign x_884 = (x_882 & x_883);
	assign x_897 = (x_895 & x_896);
	assign x_894 = (x_892 & x_893);
	assign x_904 = (x_902 & x_903);
	assign x_901 = (x_899 & x_900);
	assign x_912 = (x_910 & x_911);
	assign x_909 = (x_907 & x_908);
	assign x_919 = (x_395 & x_918);
	assign x_916 = (x_914 & x_915);
	assign x_935 = (x_933 & x_934);
	assign x_931 = (x_929 & x_930);
	assign x_928 = (x_926 & x_927);
	assign x_943 = (x_941 & x_942);
	assign x_938 = (x_936 & x_937);
	assign x_950 = (x_948 & x_949);
	assign x_946 = (x_944 & x_945);
	assign x_963 = (x_961 & x_962);
	assign x_960 = (x_958 & x_959);
	assign x_970 = (x_968 & x_969);
	assign x_967 = (x_965 & x_966);
	assign x_982 = (x_980 & x_981);
	assign x_978 = (x_976 & x_977);
	assign x_975 = (x_973 & x_974);
	assign x_985 = (x_461 & x_984);
	assign x_993 = (x_991 & x_992);
	assign x_1000 = (x_998 & x_999);
	assign x_996 = (x_994 & x_995);
	assign x_1008 = (x_1006 & x_1007);
	assign x_1003 = (x_1001 & x_1002);
	assign x_1015 = (x_1013 & x_1014);
	assign x_1011 = (x_1009 & x_1010);
	assign x_1018 = (x_494 & x_1017);
	assign x_1025 = (x_1023 & x_1024);
	assign x_1032 = (x_1030 & x_1031);
	assign x_1028 = (x_1026 & x_1027);
	assign x_520 = (((~v_127 | ~v_504)) | ~v_128);
	assign x_519 = (((~v_127 | ~v_503)) | ~v_504);
	assign x_518 = (((v_127 | v_503)) | v_504);
	assign x_517 = (((v_127 | v_504)) | v_128);
	assign x_583 = (x_581 & x_582);
	assign x_722 = (x_719 & x_721);
	assign x_862 = (x_860 & x_861);
	assign x_953 = (x_428 & x_952);
	assign x_1035 = (x_511 & x_1034);
	assign x_1052 = (x_1049 & x_1051);
	assign x_537 = (x_533 & x_536);
	assign x_544 = (x_540 & x_543);
	assign x_552 = (x_548 & x_551);
	assign x_559 = (x_556 & x_558);
	assign x_569 = (x_565 & x_568);
	assign x_576 = (x_572 & x_575);
	assign x_591 = (x_588 & x_590);
	assign x_602 = (x_598 & x_601);
	assign x_609 = (x_605 & x_608);
	assign x_617 = (x_613 & x_616);
	assign x_624 = (x_621 & x_623);
	assign x_634 = (x_630 & x_633);
	assign x_641 = (x_637 & x_640);
	assign x_649 = (x_645 & x_648);
	assign x_656 = (x_653 & x_655);
	assign x_668 = (x_664 & x_667);
	assign x_675 = (x_671 & x_674);
	assign x_683 = (x_679 & x_682);
	assign x_690 = (x_687 & x_689);
	assign x_700 = (x_696 & x_699);
	assign x_707 = (x_703 & x_706);
	assign x_715 = (x_711 & x_714);
	assign x_733 = (x_729 & x_732);
	assign x_740 = (x_736 & x_739);
	assign x_748 = (x_744 & x_747);
	assign x_755 = (x_752 & x_754);
	assign x_765 = (x_761 & x_764);
	assign x_772 = (x_769 & x_771);
	assign x_781 = (x_777 & x_780);
	assign x_788 = (x_785 & x_787);
	assign x_801 = (x_797 & x_800);
	assign x_808 = (x_804 & x_807);
	assign x_816 = (x_812 & x_815);
	assign x_823 = (x_820 & x_822);
	assign x_833 = (x_829 & x_832);
	assign x_840 = (x_836 & x_839);
	assign x_848 = (x_844 & x_847);
	assign x_855 = (x_852 & x_854);
	assign x_881 = (x_877 & x_880);
	assign x_873 = (x_869 & x_872);
	assign x_888 = (x_885 & x_887);
	assign x_898 = (x_894 & x_897);
	assign x_905 = (x_901 & x_904);
	assign x_913 = (x_909 & x_912);
	assign x_920 = (x_917 & x_919);
	assign x_932 = (x_928 & x_931);
	assign x_939 = (x_935 & x_938);
	assign x_947 = (x_943 & x_946);
	assign x_964 = (x_960 & x_963);
	assign x_971 = (x_967 & x_970);
	assign x_979 = (x_975 & x_978);
	assign x_986 = (x_983 & x_985);
	assign x_997 = (x_993 & x_996);
	assign x_1004 = (x_1000 & x_1003);
	assign x_1012 = (x_1008 & x_1011);
	assign x_1019 = (x_1016 & x_1018);
	assign x_1029 = (x_1025 & x_1028);
	assign x_1043 = (x_520 & x_521);
	assign x_1042 = (x_518 & x_519);
	assign x_1040 = (x_516 & x_517);
	assign x_584 = (x_580 & x_583);
	assign x_723 = (x_718 & x_722);
	assign x_866 = (x_862 & x_865);
	assign x_954 = (x_951 & x_953);
	assign x_1036 = (x_1033 & x_1035);
	assign x_1053 = (x_1048 & x_1052);
	assign x_545 = (x_537 & x_544);
	assign x_560 = (x_555 & x_559);
	assign x_577 = (x_569 & x_576);
	assign x_592 = (x_587 & x_591);
	assign x_610 = (x_602 & x_609);
	assign x_625 = (x_620 & x_624);
	assign x_642 = (x_634 & x_641);
	assign x_657 = (x_652 & x_656);
	assign x_676 = (x_668 & x_675);
	assign x_691 = (x_686 & x_690);
	assign x_708 = (x_700 & x_707);
	assign x_741 = (x_733 & x_740);
	assign x_756 = (x_751 & x_755);
	assign x_773 = (x_768 & x_772);
	assign x_789 = (x_784 & x_788);
	assign x_809 = (x_801 & x_808);
	assign x_824 = (x_819 & x_823);
	assign x_841 = (x_833 & x_840);
	assign x_856 = (x_851 & x_855);
	assign x_889 = (x_884 & x_888);
	assign x_906 = (x_898 & x_905);
	assign x_921 = (x_916 & x_920);
	assign x_940 = (x_932 & x_939);
	assign x_972 = (x_964 & x_971);
	assign x_987 = (x_982 & x_986);
	assign x_1005 = (x_997 & x_1004);
	assign x_1020 = (x_1015 & x_1019);
	assign x_1044 = (x_1042 & x_1043);
	assign x_1041 = (x_1039 & x_1040);
	assign x_724 = (x_715 & x_723);
	assign x_874 = (x_866 & x_873);
	assign x_955 = (x_950 & x_954);
	assign x_1037 = (x_1032 & x_1036);
	assign x_561 = (x_552 & x_560);
	assign x_593 = (x_584 & x_592);
	assign x_626 = (x_617 & x_625);
	assign x_658 = (x_649 & x_657);
	assign x_692 = (x_683 & x_691);
	assign x_757 = (x_748 & x_756);
	assign x_774 = (x_765 & x_773);
	assign x_790 = (x_781 & x_789);
	assign x_825 = (x_816 & x_824);
	assign x_857 = (x_848 & x_856);
	assign x_890 = (x_881 & x_889);
	assign x_922 = (x_913 & x_921);
	assign x_988 = (x_979 & x_987);
	assign x_1021 = (x_1012 & x_1020);
	assign x_1045 = (x_1041 & x_1044);
	assign x_725 = (x_708 & x_724);
	assign x_956 = (x_947 & x_955);
	assign x_1038 = (x_1029 & x_1037);
	assign x_562 = (x_545 & x_561);
	assign x_594 = (x_577 & x_593);
	assign x_627 = (x_610 & x_626);
	assign x_659 = (x_642 & x_658);
	assign x_693 = (x_676 & x_692);
	assign x_758 = (x_741 & x_757);
	assign x_791 = (x_774 & x_790);
	assign x_826 = (x_809 & x_825);
	assign x_858 = (x_841 & x_857);
	assign x_891 = (x_874 & x_890);
	assign x_923 = (x_906 & x_922);
	assign x_989 = (x_972 & x_988);
	assign x_1022 = (x_1005 & x_1021);
	assign x_1054 = (x_1045 & x_1053);
	assign x_957 = (x_940 & x_956);
	assign x_595 = (x_562 & x_594);
	assign x_660 = (x_627 & x_659);
	assign x_726 = (x_693 & x_725);
	assign x_792 = (x_758 & x_791);
	assign x_859 = (x_826 & x_858);
	assign x_924 = (x_891 & x_923);
	assign x_1055 = (x_1038 & x_1054);
	assign x_990 = (x_957 & x_989);
	assign x_661 = (x_595 & x_660);
	assign x_793 = (x_726 & x_792);
	assign x_925 = (x_859 & x_924);
	assign x_1056 = (x_1022 & x_1055);
	assign x_794 = (x_661 & x_793);
	assign x_1057 = (x_990 & x_1056);
	assign x_1058 = (x_925 & x_1057);
	assign x_1059 = (x_794 & x_1058);
	assign o_1 = x_105);
endmodule
