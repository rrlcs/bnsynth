module formula(v_1,v_2,v_3,v_4,v_5,v_6,v_7,v_8,v_13,v_14,v_15,v_16,v_17,v_18,v_19,v_20,v_21,v_22,v_23,v_24,v_25,v_26,v_27,v_28,v_29,v_30,v_31,v_32,v_33,v_34,v_35,v_36,v_37,v_38,v_39,v_40,v_41,v_42,v_43,v_44,v_45,v_46,v_47,v_48,v_49,v_50,v_51,v_52,v_53,v_54,v_55,v_56,v_57,v_58,v_59,v_60,v_61,v_62,v_63,v_64,v_65,v_66,v_9,v_10,v_11,v_12,v_67,v_68,v_69,v_70,v_71,v_72,v_73,v_74,v_75,v_76,v_77,v_78,v_79,v_80,v_81,v_82,v_83,v_84,v_85,v_86,v_87,v_88,v_89,v_90,v_91,v_92,v_93,v_94,v_95,v_96,v_97,v_98,v_99,v_100,v_101,v_102,v_103,v_104,v_105,v_106,v_107,v_108,v_109,v_110,v_111,v_112,v_113,v_114,v_115,v_116,v_117,v_118,v_119,v_120,v_121,v_122,v_123,v_124,v_125,v_126,v_127,v_128,v_129,v_130,v_131,v_132,v_133,v_134,v_135,v_136,v_137,v_138,v_139,v_140,v_141,v_142,v_143,v_144,v_145,v_146,v_147,v_148,v_149,v_150,v_151,v_152,v_153,v_154,v_155,v_156,v_157,v_158,v_159,v_160,v_161,v_162,v_163,v_164,v_165,v_166,v_167,v_168,v_169,v_170,v_171,v_172,v_173,v_174,v_175,v_176,v_177,v_178,v_179,v_180,v_181,v_182,v_183,v_184,v_185,v_186,v_187,v_188,v_189,v_190,v_191,v_192,v_193,v_194,v_195,v_196,v_197,v_198,v_199,v_200,v_201,v_202,v_203,v_204,v_205,v_206,v_207,v_208,v_209,v_210,v_211,v_212,v_213,v_214,v_215,v_216,v_217,v_218,v_219,v_220,v_221,v_222,v_223,v_224,v_225,v_226,v_227,v_228,v_229,v_230,v_231,v_232,v_233,v_234,v_235,v_236,v_237,v_238,v_239,v_240,v_241,v_242,v_243,v_244,v_245,v_246,v_247,v_248,v_249,v_250,v_251,v_252,v_253,v_254,v_255,v_256,v_257,v_258,v_259,v_260,v_261,v_262,v_263,v_264,v_265,v_266,v_267,v_268,v_269,v_270,v_271,v_272,v_273,v_274,v_275,v_276,v_277,v_278,v_279,v_280,v_281,v_282,v_283,v_284,v_285,v_286,v_287,v_288,v_289,v_290,v_291,v_292,v_293,v_294,v_295,v_296,v_297,v_298,v_299,v_300,v_301,v_302,v_303,v_304,v_305,v_306,v_307,v_308,v_309,v_310,v_311,v_312,v_313,v_314,v_315,v_316,v_317,v_318,v_319,v_320,v_321,v_322,v_323,v_324,v_325,v_326,v_327,v_328,v_329,v_330,v_331,v_332,v_333,v_334,v_335,v_336,v_337,v_338,v_339,v_340,v_341,v_342,v_343,v_344,v_345,v_346,v_347,v_348,v_349,v_350,v_351,v_352,v_353,v_354,v_355,v_356,v_357,v_358,v_359,v_360,v_361,v_362,v_363,v_364,v_365,v_366,v_367,v_368,v_369,v_370,v_371,v_372,v_373,v_375,v_376,v_377,v_378,v_379,v_380,v_381,v_382,v_383,v_384,v_385,v_386,v_387,v_388,v_389,v_390,v_391,v_392,v_393,v_394,v_395,v_396,v_397,v_398,v_400,v_401,v_402,v_403,v_404,v_405,v_406,v_407,v_408,v_409,v_410,v_411,v_412,v_413,v_414,v_415,v_416,v_417,v_418,v_419,v_420,v_421,v_422,v_423,v_424,v_425,v_426,v_427,v_428,v_429,v_430,v_431,v_432,v_433,v_434,v_435,v_436,v_437,v_438,v_439,v_440,v_441,v_442,v_443,v_444,v_445,v_446,v_447,v_449,v_450,v_451,v_452,v_453,v_454,v_455,v_456,v_457,v_458,v_459,v_460,v_461,v_462,v_463,v_464,v_465,v_466,v_467,v_468,v_469,v_470,v_471,v_472,v_474,v_475,v_476,v_477,v_478,v_479,v_480,v_481,v_483,v_484,v_485,v_486,v_487,v_488,v_489,v_490,v_492,v_493,v_494,v_495,v_496,v_497,v_498,v_499,v_500,v_501,v_502,v_503,v_504,v_505,v_506,v_507,v_508,v_509,v_510,v_511,v_513,v_514,v_515,v_516,v_517,v_518,v_519,v_520,v_521,v_522,v_523,v_524,v_525,v_526,v_527,v_528,v_529,v_530,v_532,v_533,v_534,v_535,v_536,v_537,v_538,v_539,v_540,v_541,v_542,v_543,v_544,v_545,v_546,v_547,v_549,v_550,v_551,v_552,v_553,v_554,v_555,v_556,v_558,v_559,v_560,v_561,v_562,v_563,v_564,v_565,v_567,v_568,v_569,v_570,v_571,v_572,v_573,v_574,v_576,v_577,v_578,v_579,v_580,v_581,v_582,v_583,v_585,v_586,v_587,v_588,v_589,v_590,v_591,v_592,v_593,v_594,v_595,v_596,v_597,v_598,v_600,v_601,v_602,v_603,v_604,v_605,v_606,v_607,v_609,v_610,v_611,v_612,v_613,v_614,v_615,v_616,o_1);
	input v_1;
	v_2;
	v_3;
	v_4;
	v_5;
	v_6;
	v_7;
	v_8;
	v_13;
	v_14;
	v_15;
	v_16;
	v_17;
	v_18;
	v_19;
	v_20;
	v_21;
	v_22;
	v_23;
	v_24;
	v_25;
	v_26;
	v_27;
	v_28;
	v_29;
	v_30;
	v_31;
	v_32;
	v_33;
	v_34;
	v_35;
	v_36;
	v_37;
	v_38;
	v_39;
	v_40;
	v_41;
	v_42;
	v_43;
	v_44;
	v_45;
	v_46;
	v_47;
	v_48;
	v_49;
	v_50;
	v_51;
	v_52;
	v_53;
	v_54;
	v_55;
	v_56;
	v_57;
	v_58;
	v_59;
	v_60;
	v_61;
	v_62;
	v_63;
	v_64;
	v_65;
	v_66;
	v_9;
	v_10;
	v_11;
	v_12;
	v_67;
	v_68;
	v_69;
	v_70;
	v_71;
	v_72;
	v_73;
	v_74;
	v_75;
	v_76;
	v_77;
	v_78;
	v_79;
	v_80;
	v_81;
	v_82;
	v_83;
	v_84;
	v_85;
	v_86;
	v_87;
	v_88;
	v_89;
	v_90;
	v_91;
	v_92;
	v_93;
	v_94;
	v_95;
	v_96;
	v_97;
	v_98;
	v_99;
	v_100;
	v_101;
	v_102;
	v_103;
	v_104;
	v_105;
	v_106;
	v_107;
	v_108;
	v_109;
	v_110;
	v_111;
	v_112;
	v_113;
	v_114;
	v_115;
	v_116;
	v_117;
	v_118;
	v_119;
	v_120;
	v_121;
	v_122;
	v_123;
	v_124;
	v_125;
	v_126;
	v_127;
	v_128;
	v_129;
	v_130;
	v_131;
	v_132;
	v_133;
	v_134;
	v_135;
	v_136;
	v_137;
	v_138;
	v_139;
	v_140;
	v_141;
	v_142;
	v_143;
	v_144;
	v_145;
	v_146;
	v_147;
	v_148;
	v_149;
	v_150;
	v_151;
	v_152;
	v_153;
	v_154;
	v_155;
	v_156;
	v_157;
	v_158;
	v_159;
	v_160;
	v_161;
	v_162;
	v_163;
	v_164;
	v_165;
	v_166;
	v_167;
	v_168;
	v_169;
	v_170;
	v_171;
	v_172;
	v_173;
	v_174;
	v_175;
	v_176;
	v_177;
	v_178;
	v_179;
	v_180;
	v_181;
	v_182;
	v_183;
	v_184;
	v_185;
	v_186;
	v_187;
	v_188;
	v_189;
	v_190;
	v_191;
	v_192;
	v_193;
	v_194;
	v_195;
	v_196;
	v_197;
	v_198;
	v_199;
	v_200;
	v_201;
	v_202;
	v_203;
	v_204;
	v_205;
	v_206;
	v_207;
	v_208;
	v_209;
	v_210;
	v_211;
	v_212;
	v_213;
	v_214;
	v_215;
	v_216;
	v_217;
	v_218;
	v_219;
	v_220;
	v_221;
	v_222;
	v_223;
	v_224;
	v_225;
	v_226;
	v_227;
	v_228;
	v_229;
	v_230;
	v_231;
	v_232;
	v_233;
	v_234;
	v_235;
	v_236;
	v_237;
	v_238;
	v_239;
	v_240;
	v_241;
	v_242;
	v_243;
	v_244;
	v_245;
	v_246;
	v_247;
	v_248;
	v_249;
	v_250;
	v_251;
	v_252;
	v_253;
	v_254;
	v_255;
	v_256;
	v_257;
	v_258;
	v_259;
	v_260;
	v_261;
	v_262;
	v_263;
	v_264;
	v_265;
	v_266;
	v_267;
	v_268;
	v_269;
	v_270;
	v_271;
	v_272;
	v_273;
	v_274;
	v_275;
	v_276;
	v_277;
	v_278;
	v_279;
	v_280;
	v_281;
	v_282;
	v_283;
	v_284;
	v_285;
	v_286;
	v_287;
	v_288;
	v_289;
	v_290;
	v_291;
	v_292;
	v_293;
	v_294;
	v_295;
	v_296;
	v_297;
	v_298;
	v_299;
	v_300;
	v_301;
	v_302;
	v_303;
	v_304;
	v_305;
	v_306;
	v_307;
	v_308;
	v_309;
	v_310;
	v_311;
	v_312;
	v_313;
	v_314;
	v_315;
	v_316;
	v_317;
	v_318;
	v_319;
	v_320;
	v_321;
	v_322;
	v_323;
	v_324;
	v_325;
	v_326;
	v_327;
	v_328;
	v_329;
	v_330;
	v_331;
	v_332;
	v_333;
	v_334;
	v_335;
	v_336;
	v_337;
	v_338;
	v_339;
	v_340;
	v_341;
	v_342;
	v_343;
	v_344;
	v_345;
	v_346;
	v_347;
	v_348;
	v_349;
	v_350;
	v_351;
	v_352;
	v_353;
	v_354;
	v_355;
	v_356;
	v_357;
	v_358;
	v_359;
	v_360;
	v_361;
	v_362;
	v_363;
	v_364;
	v_365;
	v_366;
	v_367;
	v_368;
	v_369;
	v_370;
	v_371;
	v_372;
	v_373;
	v_375;
	v_376;
	v_377;
	v_378;
	v_379;
	v_380;
	v_381;
	v_382;
	v_383;
	v_384;
	v_385;
	v_386;
	v_387;
	v_388;
	v_389;
	v_390;
	v_391;
	v_392;
	v_393;
	v_394;
	v_395;
	v_396;
	v_397;
	v_398;
	v_400;
	v_401;
	v_402;
	v_403;
	v_404;
	v_405;
	v_406;
	v_407;
	v_408;
	v_409;
	v_410;
	v_411;
	v_412;
	v_413;
	v_414;
	v_415;
	v_416;
	v_417;
	v_418;
	v_419;
	v_420;
	v_421;
	v_422;
	v_423;
	v_424;
	v_425;
	v_426;
	v_427;
	v_428;
	v_429;
	v_430;
	v_431;
	v_432;
	v_433;
	v_434;
	v_435;
	v_436;
	v_437;
	v_438;
	v_439;
	v_440;
	v_441;
	v_442;
	v_443;
	v_444;
	v_445;
	v_446;
	v_447;
	v_449;
	v_450;
	v_451;
	v_452;
	v_453;
	v_454;
	v_455;
	v_456;
	v_457;
	v_458;
	v_459;
	v_460;
	v_461;
	v_462;
	v_463;
	v_464;
	v_465;
	v_466;
	v_467;
	v_468;
	v_469;
	v_470;
	v_471;
	v_472;
	v_474;
	v_475;
	v_476;
	v_477;
	v_478;
	v_479;
	v_480;
	v_481;
	v_483;
	v_484;
	v_485;
	v_486;
	v_487;
	v_488;
	v_489;
	v_490;
	v_492;
	v_493;
	v_494;
	v_495;
	v_496;
	v_497;
	v_498;
	v_499;
	v_500;
	v_501;
	v_502;
	v_503;
	v_504;
	v_505;
	v_506;
	v_507;
	v_508;
	v_509;
	v_510;
	v_511;
	v_513;
	v_514;
	v_515;
	v_516;
	v_517;
	v_518;
	v_519;
	v_520;
	v_521;
	v_522;
	v_523;
	v_524;
	v_525;
	v_526;
	v_527;
	v_528;
	v_529;
	v_530;
	v_532;
	v_533;
	v_534;
	v_535;
	v_536;
	v_537;
	v_538;
	v_539;
	v_540;
	v_541;
	v_542;
	v_543;
	v_544;
	v_545;
	v_546;
	v_547;
	v_549;
	v_550;
	v_551;
	v_552;
	v_553;
	v_554;
	v_555;
	v_556;
	v_558;
	v_559;
	v_560;
	v_561;
	v_562;
	v_563;
	v_564;
	v_565;
	v_567;
	v_568;
	v_569;
	v_570;
	v_571;
	v_572;
	v_573;
	v_574;
	v_576;
	v_577;
	v_578;
	v_579;
	v_580;
	v_581;
	v_582;
	v_583;
	v_585;
	v_586;
	v_587;
	v_588;
	v_589;
	v_590;
	v_591;
	v_592;
	v_593;
	v_594;
	v_595;
	v_596;
	v_597;
	v_598;
	v_600;
	v_601;
	v_602;
	v_603;
	v_604;
	v_605;
	v_606;
	v_607;
	v_609;
	v_610;
	v_611;
	v_612;
	v_613;
	v_614;
	v_615;
	v_616;
	wire v_374;
	wire v_399;
	wire v_448;
	wire v_473;
	wire v_482;
	wire v_491;
	wire v_512;
	wire v_531;
	wire v_548;
	wire v_557;
	wire v_566;
	wire v_575;
	wire v_584;
	wire v_599;
	wire v_608;
	wire v_617;
	wire v_618;
	wire x_1;
	wire x_2;
	wire x_3;
	wire x_4;
	wire x_5;
	wire x_6;
	wire x_7;
	wire x_8;
	wire x_9;
	wire x_10;
	wire x_11;
	wire x_12;
	wire x_13;
	wire x_14;
	wire x_15;
	wire x_16;
	wire x_17;
	wire x_18;
	wire x_19;
	wire x_20;
	wire x_21;
	wire x_22;
	wire x_23;
	wire x_24;
	wire x_25;
	wire x_26;
	wire x_27;
	wire x_28;
	wire x_29;
	wire x_30;
	wire x_31;
	wire x_32;
	wire x_33;
	wire x_34;
	wire x_35;
	wire x_36;
	wire x_37;
	wire x_38;
	wire x_39;
	wire x_40;
	wire x_41;
	wire x_42;
	wire x_43;
	wire x_44;
	wire x_45;
	wire x_46;
	wire x_47;
	wire x_48;
	wire x_49;
	wire x_50;
	wire x_51;
	wire x_52;
	wire x_53;
	wire x_54;
	wire x_55;
	wire x_56;
	wire x_57;
	wire x_58;
	wire x_59;
	wire x_60;
	wire x_61;
	wire x_62;
	wire x_63;
	wire x_64;
	wire x_65;
	wire x_66;
	wire x_67;
	wire x_68;
	wire x_69;
	wire x_70;
	wire x_71;
	wire x_72;
	wire x_73;
	wire x_74;
	wire x_75;
	wire x_76;
	wire x_77;
	wire x_78;
	wire x_79;
	wire x_80;
	wire x_81;
	wire x_82;
	wire x_83;
	wire x_84;
	wire x_85;
	wire x_86;
	wire x_87;
	wire x_88;
	wire x_89;
	wire x_90;
	wire x_91;
	wire x_92;
	wire x_93;
	wire x_94;
	wire x_95;
	wire x_96;
	wire x_97;
	wire x_98;
	wire x_99;
	wire x_100;
	wire x_101;
	wire x_102;
	wire x_103;
	wire x_104;
	wire x_105;
	wire x_106;
	wire x_107;
	wire x_108;
	wire x_109;
	wire x_110;
	wire x_111;
	wire x_112;
	wire x_113;
	wire x_114;
	wire x_115;
	wire x_116;
	wire x_117;
	wire x_118;
	wire x_119;
	wire x_120;
	wire x_121;
	wire x_122;
	wire x_123;
	wire x_124;
	wire x_125;
	wire x_126;
	wire x_127;
	wire x_128;
	wire x_129;
	wire x_130;
	wire x_131;
	wire x_132;
	wire x_133;
	wire x_134;
	wire x_135;
	wire x_136;
	wire x_137;
	wire x_138;
	wire x_139;
	wire x_140;
	wire x_141;
	wire x_142;
	wire x_143;
	wire x_144;
	wire x_145;
	wire x_146;
	wire x_147;
	wire x_148;
	wire x_149;
	wire x_150;
	wire x_151;
	wire x_152;
	wire x_153;
	wire x_154;
	wire x_155;
	wire x_156;
	wire x_157;
	wire x_158;
	wire x_159;
	wire x_160;
	wire x_161;
	wire x_162;
	wire x_163;
	wire x_164;
	wire x_165;
	wire x_166;
	wire x_167;
	wire x_168;
	wire x_169;
	wire x_170;
	wire x_171;
	wire x_172;
	wire x_173;
	wire x_174;
	wire x_175;
	wire x_176;
	wire x_177;
	wire x_178;
	wire x_179;
	wire x_180;
	wire x_181;
	wire x_182;
	wire x_183;
	wire x_184;
	wire x_185;
	wire x_186;
	wire x_187;
	wire x_188;
	wire x_189;
	wire x_190;
	wire x_191;
	wire x_192;
	wire x_193;
	wire x_194;
	wire x_195;
	wire x_196;
	wire x_197;
	wire x_198;
	wire x_199;
	wire x_200;
	wire x_201;
	wire x_202;
	wire x_203;
	wire x_204;
	wire x_205;
	wire x_206;
	wire x_207;
	wire x_208;
	wire x_209;
	wire x_210;
	wire x_211;
	wire x_212;
	wire x_213;
	wire x_214;
	wire x_215;
	wire x_216;
	wire x_217;
	wire x_218;
	wire x_219;
	wire x_220;
	wire x_221;
	wire x_222;
	wire x_223;
	wire x_224;
	wire x_225;
	wire x_226;
	wire x_227;
	wire x_228;
	wire x_229;
	wire x_230;
	wire x_231;
	wire x_232;
	wire x_233;
	wire x_234;
	wire x_235;
	wire x_236;
	wire x_237;
	wire x_238;
	wire x_239;
	wire x_240;
	wire x_241;
	wire x_242;
	wire x_243;
	wire x_244;
	wire x_245;
	wire x_246;
	wire x_247;
	wire x_248;
	wire x_249;
	wire x_250;
	wire x_251;
	wire x_252;
	wire x_253;
	wire x_254;
	wire x_255;
	wire x_256;
	wire x_257;
	wire x_258;
	wire x_259;
	wire x_260;
	wire x_261;
	wire x_262;
	wire x_263;
	wire x_264;
	wire x_265;
	wire x_266;
	wire x_267;
	wire x_268;
	wire x_269;
	wire x_270;
	wire x_271;
	wire x_272;
	wire x_273;
	wire x_274;
	wire x_275;
	wire x_276;
	wire x_277;
	wire x_278;
	wire x_279;
	wire x_280;
	wire x_281;
	wire x_282;
	wire x_283;
	wire x_284;
	wire x_285;
	wire x_286;
	wire x_287;
	wire x_288;
	wire x_289;
	wire x_290;
	wire x_291;
	wire x_292;
	wire x_293;
	wire x_294;
	wire x_295;
	wire x_296;
	wire x_297;
	wire x_298;
	wire x_299;
	wire x_300;
	wire x_301;
	wire x_302;
	wire x_303;
	wire x_304;
	wire x_305;
	wire x_306;
	wire x_307;
	wire x_308;
	wire x_309;
	wire x_310;
	wire x_311;
	wire x_312;
	wire x_313;
	wire x_314;
	wire x_315;
	wire x_316;
	wire x_317;
	wire x_318;
	wire x_319;
	wire x_320;
	wire x_321;
	wire x_322;
	wire x_323;
	wire x_324;
	wire x_325;
	wire x_326;
	wire x_327;
	wire x_328;
	wire x_329;
	wire x_330;
	wire x_331;
	wire x_332;
	wire x_333;
	wire x_334;
	wire x_335;
	wire x_336;
	wire x_337;
	wire x_338;
	wire x_339;
	wire x_340;
	wire x_341;
	wire x_342;
	wire x_343;
	wire x_344;
	wire x_345;
	wire x_346;
	wire x_347;
	wire x_348;
	wire x_349;
	wire x_350;
	wire x_351;
	wire x_352;
	wire x_353;
	wire x_354;
	wire x_355;
	wire x_356;
	wire x_357;
	wire x_358;
	wire x_359;
	wire x_360;
	wire x_361;
	wire x_362;
	wire x_363;
	wire x_364;
	wire x_365;
	wire x_366;
	wire x_367;
	wire x_368;
	wire x_369;
	wire x_370;
	wire x_371;
	wire x_372;
	wire x_373;
	wire x_374;
	wire x_375;
	wire x_376;
	wire x_377;
	wire x_378;
	wire x_379;
	wire x_380;
	wire x_381;
	wire x_382;
	wire x_383;
	wire x_384;
	wire x_385;
	wire x_386;
	wire x_387;
	wire x_388;
	wire x_389;
	wire x_390;
	wire x_391;
	wire x_392;
	wire x_393;
	wire x_394;
	wire x_395;
	wire x_396;
	wire x_397;
	wire x_398;
	wire x_399;
	wire x_400;
	wire x_401;
	wire x_402;
	wire x_403;
	wire x_404;
	wire x_405;
	wire x_406;
	wire x_407;
	wire x_408;
	wire x_409;
	wire x_410;
	wire x_411;
	wire x_412;
	wire x_413;
	wire x_414;
	wire x_415;
	wire x_416;
	wire x_417;
	wire x_418;
	wire x_419;
	wire x_420;
	wire x_421;
	wire x_422;
	wire x_423;
	wire x_424;
	wire x_425;
	wire x_426;
	wire x_427;
	wire x_428;
	wire x_429;
	wire x_430;
	wire x_431;
	wire x_432;
	wire x_433;
	wire x_434;
	wire x_435;
	wire x_436;
	wire x_437;
	wire x_438;
	wire x_439;
	wire x_440;
	wire x_441;
	wire x_442;
	wire x_443;
	wire x_444;
	wire x_445;
	wire x_446;
	wire x_447;
	wire x_448;
	wire x_449;
	wire x_450;
	wire x_451;
	wire x_452;
	wire x_453;
	wire x_454;
	wire x_455;
	wire x_456;
	wire x_457;
	wire x_458;
	wire x_459;
	wire x_460;
	wire x_461;
	wire x_462;
	wire x_463;
	wire x_464;
	wire x_465;
	wire x_466;
	wire x_467;
	wire x_468;
	wire x_469;
	wire x_470;
	wire x_471;
	wire x_472;
	wire x_473;
	wire x_474;
	wire x_475;
	wire x_476;
	wire x_477;
	wire x_478;
	wire x_479;
	wire x_480;
	wire x_481;
	wire x_482;
	wire x_483;
	wire x_484;
	wire x_485;
	wire x_486;
	wire x_487;
	wire x_488;
	wire x_489;
	wire x_490;
	wire x_491;
	wire x_492;
	wire x_493;
	wire x_494;
	wire x_495;
	wire x_496;
	wire x_497;
	wire x_498;
	wire x_499;
	wire x_500;
	wire x_501;
	wire x_502;
	wire x_503;
	wire x_504;
	wire x_505;
	wire x_506;
	wire x_507;
	wire x_508;
	wire x_509;
	wire x_510;
	wire x_511;
	wire x_512;
	wire x_513;
	wire x_514;
	wire x_515;
	wire x_516;
	wire x_517;
	wire x_518;
	wire x_519;
	wire x_520;
	wire x_521;
	wire x_522;
	wire x_523;
	wire x_524;
	wire x_525;
	wire x_526;
	wire x_527;
	wire x_528;
	wire x_529;
	wire x_530;
	wire x_531;
	wire x_532;
	wire x_533;
	wire x_534;
	wire x_535;
	wire x_536;
	wire x_537;
	wire x_538;
	wire x_539;
	wire x_540;
	wire x_541;
	wire x_542;
	wire x_543;
	wire x_544;
	wire x_545;
	wire x_546;
	wire x_547;
	wire x_548;
	wire x_549;
	wire x_550;
	wire x_551;
	wire x_552;
	wire x_553;
	wire x_554;
	wire x_555;
	wire x_556;
	wire x_557;
	wire x_558;
	wire x_559;
	wire x_560;
	wire x_561;
	wire x_562;
	wire x_563;
	wire x_564;
	wire x_565;
	wire x_566;
	wire x_567;
	wire x_568;
	wire x_569;
	wire x_570;
	wire x_571;
	wire x_572;
	wire x_573;
	wire x_574;
	wire x_575;
	wire x_576;
	wire x_577;
	wire x_578;
	wire x_579;
	wire x_580;
	wire x_581;
	wire x_582;
	wire x_583;
	wire x_584;
	wire x_585;
	wire x_586;
	wire x_587;
	wire x_588;
	wire x_589;
	wire x_590;
	wire x_591;
	wire x_592;
	wire x_593;
	wire x_594;
	wire x_595;
	wire x_596;
	wire x_597;
	wire x_598;
	wire x_599;
	wire x_600;
	wire x_601;
	wire x_602;
	wire x_603;
	wire x_604;
	wire x_605;
	wire x_606;
	wire x_607;
	wire x_608;
	wire x_609;
	wire x_610;
	wire x_611;
	wire x_612;
	wire x_613;
	wire x_614;
	wire x_615;
	wire x_616;
	wire x_617;
	wire x_618;
	wire x_619;
	wire x_620;
	wire x_621;
	wire x_622;
	wire x_623;
	wire x_624;
	wire x_625;
	wire x_626;
	wire x_627;
	wire x_628;
	wire x_629;
	wire x_630;
	wire x_631;
	wire x_632;
	wire x_633;
	wire x_634;
	wire x_635;
	wire x_636;
	wire x_637;
	wire x_638;
	wire x_639;
	wire x_640;
	wire x_641;
	wire x_642;
	wire x_643;
	wire x_644;
	wire x_645;
	wire x_646;
	wire x_647;
	wire x_648;
	wire x_649;
	wire x_650;
	wire x_651;
	wire x_652;
	wire x_653;
	wire x_654;
	wire x_655;
	wire x_656;
	wire x_657;
	wire x_658;
	wire x_659;
	wire x_660;
	wire x_661;
	wire x_662;
	wire x_663;
	wire x_664;
	wire x_665;
	wire x_666;
	wire x_667;
	wire x_668;
	wire x_669;
	wire x_670;
	wire x_671;
	wire x_672;
	wire x_673;
	wire x_674;
	wire x_675;
	wire x_676;
	wire x_677;
	wire x_678;
	wire x_679;
	wire x_680;
	wire x_681;
	wire x_682;
	wire x_683;
	wire x_684;
	wire x_685;
	wire x_686;
	wire x_687;
	wire x_688;
	wire x_689;
	wire x_690;
	wire x_691;
	wire x_692;
	wire x_693;
	wire x_694;
	wire x_695;
	wire x_696;
	wire x_697;
	wire x_698;
	wire x_699;
	wire x_700;
	wire x_701;
	wire x_702;
	wire x_703;
	wire x_704;
	wire x_705;
	wire x_706;
	wire x_707;
	wire x_708;
	wire x_709;
	wire x_710;
	wire x_711;
	wire x_712;
	wire x_713;
	wire x_714;
	wire x_715;
	wire x_716;
	wire x_717;
	wire x_718;
	wire x_719;
	wire x_720;
	wire x_721;
	wire x_722;
	wire x_723;
	wire x_724;
	wire x_725;
	wire x_726;
	wire x_727;
	wire x_728;
	wire x_729;
	wire x_730;
	wire x_731;
	wire x_732;
	wire x_733;
	wire x_734;
	wire x_735;
	wire x_736;
	wire x_737;
	wire x_738;
	wire x_739;
	wire x_740;
	wire x_741;
	wire x_742;
	wire x_743;
	wire x_744;
	wire x_745;
	wire x_746;
	wire x_747;
	wire x_748;
	wire x_749;
	wire x_750;
	wire x_751;
	wire x_752;
	wire x_753;
	wire x_754;
	wire x_755;
	wire x_756;
	wire x_757;
	wire x_758;
	wire x_759;
	wire x_760;
	wire x_761;
	wire x_762;
	wire x_763;
	wire x_764;
	wire x_765;
	wire x_766;
	wire x_767;
	wire x_768;
	wire x_769;
	wire x_770;
	wire x_771;
	wire x_772;
	wire x_773;
	wire x_774;
	wire x_775;
	wire x_776;
	wire x_777;
	wire x_778;
	wire x_779;
	wire x_780;
	wire x_781;
	wire x_782;
	wire x_783;
	wire x_784;
	wire x_785;
	wire x_786;
	wire x_787;
	wire x_788;
	wire x_789;
	wire x_790;
	wire x_791;
	wire x_792;
	wire x_793;
	wire x_794;
	wire x_795;
	wire x_796;
	wire x_797;
	wire x_798;
	wire x_799;
	wire x_800;
	wire x_801;
	wire x_802;
	wire x_803;
	wire x_804;
	wire x_805;
	wire x_806;
	wire x_807;
	wire x_808;
	wire x_809;
	wire x_810;
	wire x_811;
	wire x_812;
	wire x_813;
	wire x_814;
	wire x_815;
	wire x_816;
	wire x_817;
	wire x_818;
	wire x_819;
	wire x_820;
	wire x_821;
	wire x_822;
	wire x_823;
	wire x_824;
	wire x_825;
	wire x_826;
	wire x_827;
	wire x_828;
	wire x_829;
	wire x_830;
	wire x_831;
	wire x_832;
	wire x_833;
	wire x_834;
	wire x_835;
	wire x_836;
	wire x_837;
	wire x_838;
	wire x_839;
	wire x_840;
	wire x_841;
	wire x_842;
	wire x_843;
	wire x_844;
	wire x_845;
	wire x_846;
	wire x_847;
	wire x_848;
	wire x_849;
	wire x_850;
	wire x_851;
	wire x_852;
	wire x_853;
	wire x_854;
	wire x_855;
	wire x_856;
	wire x_857;
	wire x_858;
	wire x_859;
	wire x_860;
	wire x_861;
	wire x_862;
	wire x_863;
	wire x_864;
	wire x_865;
	wire x_866;
	wire x_867;
	wire x_868;
	wire x_869;
	wire x_870;
	wire x_871;
	wire x_872;
	wire x_873;
	wire x_874;
	wire x_875;
	wire x_876;
	wire x_877;
	wire x_878;
	wire x_879;
	wire x_880;
	wire x_881;
	wire x_882;
	wire x_883;
	wire x_884;
	wire x_885;
	wire x_886;
	wire x_887;
	wire x_888;
	wire x_889;
	wire x_890;
	wire x_891;
	wire x_892;
	wire x_893;
	wire x_894;
	wire x_895;
	wire x_896;
	wire x_897;
	wire x_898;
	wire x_899;
	wire x_900;
	wire x_901;
	wire x_902;
	wire x_903;
	wire x_904;
	wire x_905;
	wire x_906;
	wire x_907;
	wire x_908;
	wire x_909;
	wire x_910;
	wire x_911;
	wire x_912;
	wire x_913;
	wire x_914;
	wire x_915;
	wire x_916;
	wire x_917;
	wire x_918;
	wire x_919;
	wire x_920;
	wire x_921;
	wire x_922;
	wire x_923;
	wire x_924;
	wire x_925;
	wire x_926;
	wire x_927;
	wire x_928;
	wire x_929;
	wire x_930;
	wire x_931;
	wire x_932;
	wire x_933;
	wire x_934;
	wire x_935;
	wire x_936;
	wire x_937;
	wire x_938;
	wire x_939;
	wire x_940;
	wire x_941;
	wire x_942;
	wire x_943;
	wire x_944;
	wire x_945;
	wire x_946;
	wire x_947;
	wire x_948;
	wire x_949;
	wire x_950;
	wire x_951;
	wire x_952;
	wire x_953;
	wire x_954;
	wire x_955;
	wire x_956;
	wire x_957;
	wire x_958;
	wire x_959;
	wire x_960;
	wire x_961;
	wire x_962;
	wire x_963;
	wire x_964;
	wire x_965;
	wire x_966;
	wire x_967;
	wire x_968;
	wire x_969;
	wire x_970;
	wire x_971;
	wire x_972;
	wire x_973;
	wire x_974;
	wire x_975;
	wire x_976;
	wire x_977;
	wire x_978;
	wire x_979;
	wire x_980;
	wire x_981;
	wire x_982;
	wire x_983;
	wire x_984;
	wire x_985;
	wire x_986;
	wire x_987;
	wire x_988;
	wire x_989;
	wire x_990;
	wire x_991;
	wire x_992;
	wire x_993;
	wire x_994;
	wire x_995;
	wire x_996;
	wire x_997;
	wire x_998;
	wire x_999;
	wire x_1000;
	wire x_1001;
	wire x_1002;
	wire x_1003;
	wire x_1004;
	wire x_1005;
	wire x_1006;
	wire x_1007;
	wire x_1008;
	wire x_1009;
	wire x_1010;
	wire x_1011;
	wire x_1012;
	wire x_1013;
	wire x_1014;
	wire x_1015;
	wire x_1016;
	wire x_1017;
	wire x_1018;
	wire x_1019;
	wire x_1020;
	wire x_1021;
	wire x_1022;
	wire x_1023;
	wire x_1024;
	wire x_1025;
	wire x_1026;
	wire x_1027;
	wire x_1028;
	wire x_1029;
	wire x_1030;
	wire x_1031;
	wire x_1032;
	wire x_1033;
	wire x_1034;
	wire x_1035;
	wire x_1036;
	wire x_1037;
	wire x_1038;
	wire x_1039;
	wire x_1040;
	wire x_1041;
	wire x_1042;
	wire x_1043;
	wire x_1044;
	wire x_1045;
	wire x_1046;
	wire x_1047;
	wire x_1048;
	wire x_1049;
	wire x_1050;
	wire x_1051;
	wire x_1052;
	wire x_1053;
	wire x_1054;
	wire x_1055;
	wire x_1056;
	wire x_1057;
	wire x_1058;
	wire x_1059;
	wire x_1060;
	wire x_1061;
	wire x_1062;
	wire x_1063;
	wire x_1064;
	wire x_1065;
	wire x_1066;
	wire x_1067;
	wire x_1068;
	wire x_1069;
	wire x_1070;
	wire x_1071;
	wire x_1072;
	wire x_1073;
	wire x_1074;
	wire x_1075;
	wire x_1076;
	wire x_1077;
	wire x_1078;
	wire x_1079;
	wire x_1080;
	wire x_1081;
	wire x_1082;
	wire x_1083;
	wire x_1084;
	wire x_1085;
	wire x_1086;
	wire x_1087;
	wire x_1088;
	wire x_1089;
	wire x_1090;
	wire x_1091;
	wire x_1092;
	wire x_1093;
	wire x_1094;
	wire x_1095;
	wire x_1096;
	wire x_1097;
	wire x_1098;
	wire x_1099;
	wire x_1100;
	wire x_1101;
	wire x_1102;
	wire x_1103;
	wire x_1104;
	wire x_1105;
	wire x_1106;
	wire x_1107;
	wire x_1108;
	wire x_1109;
	wire x_1110;
	wire x_1111;
	wire x_1112;
	wire x_1113;
	wire x_1114;
	wire x_1115;
	wire x_1116;
	wire x_1117;
	wire x_1118;
	wire x_1119;
	wire x_1120;
	wire x_1121;
	wire x_1122;
	wire x_1123;
	wire x_1124;
	wire x_1125;
	wire x_1126;
	wire x_1127;
	wire x_1128;
	wire x_1129;
	wire x_1130;
	wire x_1131;
	wire x_1132;
	wire x_1133;
	wire x_1134;
	wire x_1135;
	wire x_1136;
	wire x_1137;
	wire x_1138;
	wire x_1139;
	wire x_1140;
	wire x_1141;
	wire x_1142;
	wire x_1143;
	wire x_1144;
	wire x_1145;
	wire x_1146;
	wire x_1147;
	wire x_1148;
	wire x_1149;
	wire x_1150;
	wire x_1151;
	wire x_1152;
	wire x_1153;
	wire x_1154;
	wire x_1155;
	wire x_1156;
	wire x_1157;
	wire x_1158;
	wire x_1159;
	wire x_1160;
	wire x_1161;
	wire x_1162;
	wire x_1163;
	wire x_1164;
	wire x_1165;
	wire x_1166;
	wire x_1167;
	wire x_1168;
	wire x_1169;
	wire x_1170;
	wire x_1171;
	wire x_1172;
	wire x_1173;
	wire x_1174;
	wire x_1175;
	wire x_1176;
	wire x_1177;
	wire x_1178;
	wire x_1179;
	wire x_1180;
	wire x_1181;
	wire x_1182;
	wire x_1183;
	wire x_1184;
	wire x_1185;
	wire x_1186;
	wire x_1187;
	wire x_1188;
	wire x_1189;
	wire x_1190;
	wire x_1191;
	wire x_1192;
	wire x_1193;
	wire x_1194;
	wire x_1195;
	wire x_1196;
	wire x_1197;
	wire x_1198;
	wire x_1199;
	wire x_1200;
	wire x_1201;
	wire x_1202;
	wire x_1203;
	wire x_1204;
	wire x_1205;
	wire x_1206;
	wire x_1207;
	wire x_1208;
	wire x_1209;
	wire x_1210;
	wire x_1211;
	wire x_1212;
	wire x_1213;
	wire x_1214;
	wire x_1215;
	wire x_1216;
	wire x_1217;
	wire x_1218;
	wire x_1219;
	wire x_1220;
	wire x_1221;
	wire x_1222;
	wire x_1223;
	wire x_1224;
	wire x_1225;
	wire x_1226;
	wire x_1227;
	wire x_1228;
	wire x_1229;
	wire x_1230;
	wire x_1231;
	wire x_1232;
	wire x_1233;
	wire x_1234;
	wire x_1235;
	wire x_1236;
	wire x_1237;
	wire x_1238;
	wire x_1239;
	wire x_1240;
	wire x_1241;
	wire x_1242;
	wire x_1243;
	wire x_1244;
	wire x_1245;
	wire x_1246;
	wire x_1247;
	wire x_1248;
	wire x_1249;
	wire x_1250;
	wire x_1251;
	wire x_1252;
	wire x_1253;
	wire x_1254;
	wire x_1255;
	wire x_1256;
	wire x_1257;
	wire x_1258;
	wire x_1259;
	wire x_1260;
	wire x_1261;
	wire x_1262;
	wire x_1263;
	wire x_1264;
	wire x_1265;
	wire x_1266;
	wire x_1267;
	wire x_1268;
	wire x_1269;
	wire x_1270;
	wire x_1271;
	wire x_1272;
	wire x_1273;
	wire x_1274;
	wire x_1275;
	wire x_1276;
	wire x_1277;
	wire x_1278;
	wire x_1279;
	wire x_1280;
	wire x_1281;
	wire x_1282;
	wire x_1283;
	wire x_1284;
	wire x_1285;
	wire x_1286;
	wire x_1287;
	wire x_1288;
	wire x_1289;
	wire x_1290;
	wire x_1291;
	wire x_1292;
	wire x_1293;
	wire x_1294;
	wire x_1295;
	wire x_1296;
	wire x_1297;
	wire x_1298;
	wire x_1299;
	wire x_1300;
	wire x_1301;
	wire x_1302;
	wire x_1303;
	wire x_1304;
	wire x_1305;
	wire x_1306;
	wire x_1307;
	wire x_1308;
	wire x_1309;
	wire x_1310;
	wire x_1311;
	wire x_1312;
	wire x_1313;
	wire x_1314;
	wire x_1315;
	wire x_1316;
	wire x_1317;
	wire x_1318;
	wire x_1319;
	wire x_1320;
	wire x_1321;
	wire x_1322;
	wire x_1323;
	wire x_1324;
	wire x_1325;
	wire x_1326;
	wire x_1327;
	wire x_1328;
	wire x_1329;
	wire x_1330;
	wire x_1331;
	wire x_1332;
	wire x_1333;
	wire x_1334;
	wire x_1335;
	wire x_1336;
	wire x_1337;
	wire x_1338;
	wire x_1339;
	wire x_1340;
	wire x_1341;
	wire x_1342;
	wire x_1343;
	wire x_1344;
	wire x_1345;
	wire x_1346;
	wire x_1347;
	wire x_1348;
	wire x_1349;
	wire x_1350;
	wire x_1351;
	wire x_1352;
	wire x_1353;
	wire x_1354;
	wire x_1355;
	wire x_1356;
	wire x_1357;
	wire x_1358;
	wire x_1359;
	wire x_1360;
	wire x_1361;
	wire x_1362;
	wire x_1363;
	wire x_1364;
	wire x_1365;
	wire x_1366;
	wire x_1367;
	wire x_1368;
	wire x_1369;
	wire x_1370;
	wire x_1371;
	wire x_1372;
	wire x_1373;
	wire x_1374;
	wire x_1375;
	wire x_1376;
	wire x_1377;
	wire x_1378;
	wire x_1379;
	wire x_1380;
	wire x_1381;
	wire x_1382;
	wire x_1383;
	wire x_1384;
	wire x_1385;
	wire x_1386;
	wire x_1387;
	wire x_1388;
	wire x_1389;
	wire x_1390;
	wire x_1391;
	wire x_1392;
	wire x_1393;
	wire x_1394;
	wire x_1395;
	wire x_1396;
	wire x_1397;
	wire x_1398;
	wire x_1399;
	wire x_1400;
	wire x_1401;
	wire x_1402;
	wire x_1403;
	wire x_1404;
	wire x_1405;
	wire x_1406;
	wire x_1407;
	wire x_1408;
	wire x_1409;
	wire x_1410;
	wire x_1411;
	wire x_1412;
	wire x_1413;
	wire x_1414;
	wire x_1415;
	wire x_1416;
	wire x_1417;
	wire x_1418;
	wire x_1419;
	wire x_1420;
	wire x_1421;
	wire x_1422;
	wire x_1423;
	wire x_1424;
	wire x_1425;
	wire x_1426;
	wire x_1427;
	wire x_1428;
	wire x_1429;
	wire x_1430;
	wire x_1431;
	wire x_1432;
	wire x_1433;
	wire x_1434;
	wire x_1435;
	wire x_1436;
	wire x_1437;
	wire x_1438;
	wire x_1439;
	wire x_1440;
	wire x_1441;
	wire x_1442;
	wire x_1443;
	wire x_1444;
	wire x_1445;
	wire x_1446;
	wire x_1447;
	wire x_1448;
	wire x_1449;
	wire x_1450;
	wire x_1451;
	wire x_1452;
	wire x_1453;
	wire x_1454;
	wire x_1455;
	wire x_1456;
	wire x_1457;
	wire x_1458;
	wire x_1459;
	wire x_1460;
	wire x_1461;
	wire x_1462;
	wire x_1463;
	wire x_1464;
	wire x_1465;
	wire x_1466;
	wire x_1467;
	wire x_1468;
	wire x_1469;
	wire x_1470;
	wire x_1471;
	wire x_1472;
	wire x_1473;
	wire x_1474;
	wire x_1475;
	wire x_1476;
	wire x_1477;
	wire x_1478;
	wire x_1479;
	wire x_1480;
	wire x_1481;
	wire x_1482;
	wire x_1483;
	wire x_1484;
	wire x_1485;
	wire x_1486;
	wire x_1487;
	wire x_1488;
	wire x_1489;
	wire x_1490;
	wire x_1491;
	wire x_1492;
	wire x_1493;
	wire x_1494;
	wire x_1495;
	wire x_1496;
	wire x_1497;
	wire x_1498;
	wire x_1499;
	wire x_1500;
	wire x_1501;
	wire x_1502;
	wire x_1503;
	wire x_1504;
	wire x_1505;
	wire x_1506;
	wire x_1507;
	wire x_1508;
	wire x_1509;
	wire x_1510;
	wire x_1511;
	wire x_1512;
	wire x_1513;
	wire x_1514;
	wire x_1515;
	wire x_1516;
	wire x_1517;
	wire x_1518;
	wire x_1519;
	wire x_1520;
	wire x_1521;
	wire x_1522;
	wire x_1523;
	wire x_1524;
	wire x_1525;
	wire x_1526;
	wire x_1527;
	wire x_1528;
	wire x_1529;
	wire x_1530;
	wire x_1531;
	wire x_1532;
	wire x_1533;
	wire x_1534;
	wire x_1535;
	wire x_1536;
	wire x_1537;
	wire x_1538;
	wire x_1539;
	wire x_1540;
	wire x_1541;
	wire x_1542;
	wire x_1543;
	wire x_1544;
	wire x_1545;
	wire x_1546;
	wire x_1547;
	wire x_1548;
	wire x_1549;
	wire x_1550;
	wire x_1551;
	wire x_1552;
	wire x_1553;
	wire x_1554;
	wire x_1555;
	wire x_1556;
	wire x_1557;
	wire x_1558;
	wire x_1559;
	wire x_1560;
	wire x_1561;
	wire x_1562;
	wire x_1563;
	wire x_1564;
	wire x_1565;
	wire x_1566;
	wire x_1567;
	wire x_1568;
	wire x_1569;
	wire x_1570;
	wire x_1571;
	wire x_1572;
	wire x_1573;
	wire x_1574;
	wire x_1575;
	wire x_1576;
	wire x_1577;
	wire x_1578;
	wire x_1579;
	wire x_1580;
	wire x_1581;
	wire x_1582;
	wire x_1583;
	wire x_1584;
	wire x_1585;
	wire x_1586;
	wire x_1587;
	wire x_1588;
	wire x_1589;
	wire x_1590;
	wire x_1591;
	wire x_1592;
	wire x_1593;
	wire x_1594;
	wire x_1595;
	wire x_1596;
	wire x_1597;
	wire x_1598;
	wire x_1599;
	wire x_1600;
	wire x_1601;
	wire x_1602;
	wire x_1603;
	wire x_1604;
	wire x_1605;
	wire x_1606;
	wire x_1607;
	wire x_1608;
	wire x_1609;
	wire x_1610;
	wire x_1611;
	wire x_1612;
	wire x_1613;
	wire x_1614;
	wire x_1615;
	wire x_1616;
	wire x_1617;
	wire x_1618;
	wire x_1619;
	wire x_1620;
	wire x_1621;
	wire x_1622;
	wire x_1623;
	wire x_1624;
	wire x_1625;
	wire x_1626;
	wire x_1627;
	wire x_1628;
	wire x_1629;
	wire x_1630;
	wire x_1631;
	wire x_1632;
	wire x_1633;
	wire x_1634;
	wire x_1635;
	wire x_1636;
	wire x_1637;
	wire x_1638;
	wire x_1639;
	wire x_1640;
	wire x_1641;
	wire x_1642;
	wire x_1643;
	wire x_1644;
	wire x_1645;
	wire x_1646;
	wire x_1647;
	wire x_1648;
	wire x_1649;
	wire x_1650;
	wire x_1651;
	wire x_1652;
	wire x_1653;
	wire x_1654;
	wire x_1655;
	wire x_1656;
	wire x_1657;
	wire x_1658;
	wire x_1659;
	wire x_1660;
	wire x_1661;
	wire x_1662;
	wire x_1663;
	wire x_1664;
	wire x_1665;
	wire x_1666;
	wire x_1667;
	wire x_1668;
	wire x_1669;
	wire x_1670;
	wire x_1671;
	wire x_1672;
	wire x_1673;
	wire x_1674;
	wire x_1675;
	wire x_1676;
	wire x_1677;
	wire x_1678;
	wire x_1679;
	wire x_1680;
	wire x_1681;
	wire x_1682;
	wire x_1683;
	wire x_1684;
	wire x_1685;
	wire x_1686;
	wire x_1687;
	wire x_1688;
	wire x_1689;
	wire x_1690;
	wire x_1691;
	wire x_1692;
	wire x_1693;
	wire x_1694;
	wire x_1695;
	wire x_1696;
	wire x_1697;
	wire x_1698;
	wire x_1699;
	wire x_1700;
	wire x_1701;
	wire x_1702;
	wire x_1703;
	wire x_1704;
	wire x_1705;
	wire x_1706;
	wire x_1707;
	wire x_1708;
	wire x_1709;
	wire x_1710;
	wire x_1711;
	wire x_1712;
	wire x_1713;
	wire x_1714;
	wire x_1715;
	wire x_1716;
	wire x_1717;
	wire x_1718;
	wire x_1719;
	wire x_1720;
	wire x_1721;
	wire x_1722;
	wire x_1723;
	wire x_1724;
	wire x_1725;
	wire x_1726;
	wire x_1727;
	wire x_1728;
	wire x_1729;
	wire x_1730;
	wire x_1731;
	wire x_1732;
	wire x_1733;
	wire x_1734;
	wire x_1735;
	wire x_1736;
	wire x_1737;
	wire x_1738;
	wire x_1739;
	wire x_1740;
	wire x_1741;
	wire x_1742;
	wire x_1743;
	wire x_1744;
	wire x_1745;
	wire x_1746;
	wire x_1747;
	wire x_1748;
	wire x_1749;
	wire x_1750;
	wire x_1751;
	wire x_1752;
	wire x_1753;
	wire x_1754;
	wire x_1755;
	wire x_1756;
	wire x_1757;
	wire x_1758;
	wire x_1759;
	wire x_1760;
	wire x_1761;
	wire x_1762;
	wire x_1763;
	wire x_1764;
	wire x_1765;
	wire x_1766;
	wire x_1767;
	wire x_1768;
	wire x_1769;
	wire x_1770;
	wire x_1771;
	wire x_1772;
	wire x_1773;
	wire x_1774;
	wire x_1775;
	wire x_1776;
	wire x_1777;
	wire x_1778;
	wire x_1779;
	wire x_1780;
	wire x_1781;
	wire x_1782;
	wire x_1783;
	wire x_1784;
	wire x_1785;
	wire x_1786;
	wire x_1787;
	wire x_1788;
	wire x_1789;
	wire x_1790;
	wire x_1791;
	wire x_1792;
	wire x_1793;
	wire x_1794;
	wire x_1795;
	wire x_1796;
	wire x_1797;
	wire x_1798;
	wire x_1799;
	wire x_1800;
	wire x_1801;
	wire x_1802;
	wire x_1803;
	wire x_1804;
	wire x_1805;
	wire x_1806;
	wire x_1807;
	wire x_1808;
	wire x_1809;
	wire x_1810;
	wire x_1811;
	wire x_1812;
	wire x_1813;
	wire x_1814;
	wire x_1815;
	wire x_1816;
	wire x_1817;
	wire x_1818;
	wire x_1819;
	wire x_1820;
	wire x_1821;
	wire x_1822;
	wire x_1823;
	wire x_1824;
	wire x_1825;
	wire x_1826;
	wire x_1827;
	wire x_1828;
	wire x_1829;
	wire x_1830;
	wire x_1831;
	wire x_1832;
	wire x_1833;
	wire x_1834;
	wire x_1835;
	wire x_1836;
	wire x_1837;
	wire x_1838;
	wire x_1839;
	wire x_1840;
	wire x_1841;
	wire x_1842;
	wire x_1843;
	wire x_1844;
	wire x_1845;
	wire x_1846;
	wire x_1847;
	wire x_1848;
	wire x_1849;
	wire x_1850;
	wire x_1851;
	wire x_1852;
	wire x_1853;
	wire x_1854;
	wire x_1855;
	wire x_1856;
	wire x_1857;
	wire x_1858;
	wire x_1859;
	wire x_1860;
	wire x_1861;
	wire x_1862;
	wire x_1863;
	wire x_1864;
	wire x_1865;
	wire x_1866;
	wire x_1867;
	wire x_1868;
	wire x_1869;
	wire x_1870;
	wire x_1871;
	wire x_1872;
	wire x_1873;
	wire x_1874;
	wire x_1875;
	wire x_1876;
	wire x_1877;
	wire x_1878;
	wire x_1879;
	wire x_1880;
	wire x_1881;
	wire x_1882;
	wire x_1883;
	wire x_1884;
	wire x_1885;
	wire x_1886;
	wire x_1887;
	wire x_1888;
	wire x_1889;
	wire x_1890;
	wire x_1891;
	wire x_1892;
	wire x_1893;
	wire x_1894;
	wire x_1895;
	wire x_1896;
	wire x_1897;
	wire x_1898;
	wire x_1899;
	wire x_1900;
	wire x_1901;
	wire x_1902;
	wire x_1903;
	wire x_1904;
	wire x_1905;
	wire x_1906;
	wire x_1907;
	wire x_1908;
	wire x_1909;
	wire x_1910;
	wire x_1911;
	wire x_1912;
	wire x_1913;
	wire x_1914;
	wire x_1915;
	wire x_1916;
	wire x_1917;
	wire x_1918;
	wire x_1919;
	wire x_1920;
	wire x_1921;
	wire x_1922;
	wire x_1923;
	wire x_1924;
	wire x_1925;
	wire x_1926;
	wire x_1927;
	wire x_1928;
	wire x_1929;
	wire x_1930;
	wire x_1931;
	wire x_1932;
	wire x_1933;
	wire x_1934;
	wire x_1935;
	wire x_1936;
	wire x_1937;
	wire x_1938;
	wire x_1939;
	wire x_1940;
	wire x_1941;
	wire x_1942;
	wire x_1943;
	wire x_1944;
	wire x_1945;
	wire x_1946;
	wire x_1947;
	wire x_1948;
	wire x_1949;
	wire x_1950;
	wire x_1951;
	wire x_1952;
	wire x_1953;
	wire x_1954;
	wire x_1955;
	wire x_1956;
	wire x_1957;
	wire x_1958;
	wire x_1959;
	wire x_1960;
	wire x_1961;
	wire x_1962;
	wire x_1963;
	wire x_1964;
	wire x_1965;
	wire x_1966;
	wire x_1967;
	wire x_1968;
	wire x_1969;
	wire x_1970;
	wire x_1971;
	wire x_1972;
	wire x_1973;
	wire x_1974;
	wire x_1975;
	wire x_1976;
	wire x_1977;
	wire x_1978;
	wire x_1979;
	wire x_1980;
	wire x_1981;
	wire x_1982;
	wire x_1983;
	wire x_1984;
	wire x_1985;
	wire x_1986;
	wire x_1987;
	wire x_1988;
	wire x_1989;
	wire x_1990;
	wire x_1991;
	wire x_1992;
	wire x_1993;
	wire x_1994;
	wire x_1995;
	wire x_1996;
	wire x_1997;
	wire x_1998;
	wire x_1999;
	wire x_2000;
	wire x_2001;
	wire x_2002;
	wire x_2003;
	wire x_2004;
	wire x_2005;
	wire x_2006;
	wire x_2007;
	wire x_2008;
	wire x_2009;
	wire x_2010;
	wire x_2011;
	wire x_2012;
	wire x_2013;
	wire x_2014;
	wire x_2015;
	wire x_2016;
	wire x_2017;
	wire x_2018;
	wire x_2019;
	wire x_2020;
	wire x_2021;
	wire x_2022;
	wire x_2023;
	wire x_2024;
	wire x_2025;
	wire x_2026;
	wire x_2027;
	wire x_2028;
	wire x_2029;
	wire x_2030;
	wire x_2031;
	wire x_2032;
	wire x_2033;
	wire x_2034;
	wire x_2035;
	wire x_2036;
	wire x_2037;
	wire x_2038;
	wire x_2039;
	wire x_2040;
	wire x_2041;
	wire x_2042;
	wire x_2043;
	wire x_2044;
	wire x_2045;
	wire x_2046;
	wire x_2047;
	wire x_2048;
	wire x_2049;
	wire x_2050;
	wire x_2051;
	wire x_2052;
	wire x_2053;
	wire x_2054;
	wire x_2055;
	wire x_2056;
	wire x_2057;
	wire x_2058;
	wire x_2059;
	wire x_2060;
	wire x_2061;
	wire x_2062;
	wire x_2063;
	wire x_2064;
	wire x_2065;
	wire x_2066;
	wire x_2067;
	wire x_2068;
	wire x_2069;
	wire x_2070;
	wire x_2071;
	wire x_2072;
	wire x_2073;
	wire x_2074;
	wire x_2075;
	wire x_2076;
	wire x_2077;
	wire x_2078;
	wire x_2079;
	wire x_2080;
	wire x_2081;
	wire x_2082;
	wire x_2083;
	wire x_2084;
	wire x_2085;
	wire x_2086;
	wire x_2087;
	wire x_2088;
	wire x_2089;
	wire x_2090;
	wire x_2091;
	wire x_2092;
	wire x_2093;
	wire x_2094;
	wire x_2095;
	wire x_2096;
	wire x_2097;
	wire x_2098;
	wire x_2099;
	wire x_2100;
	wire x_2101;
	wire x_2102;
	wire x_2103;
	wire x_2104;
	wire x_2105;
	wire x_2106;
	wire x_2107;
	wire x_2108;
	wire x_2109;
	wire x_2110;
	wire x_2111;
	wire x_2112;
	wire x_2113;
	wire x_2114;
	wire x_2115;
	wire x_2116;
	wire x_2117;
	wire x_2118;
	wire x_2119;
	wire x_2120;
	wire x_2121;
	wire x_2122;
	wire x_2123;
	wire x_2124;
	wire x_2125;
	wire x_2126;
	wire x_2127;
	wire x_2128;
	wire x_2129;
	wire x_2130;
	wire x_2131;
	wire x_2132;
	wire x_2133;
	wire x_2134;
	wire x_2135;
	wire x_2136;
	wire x_2137;
	wire x_2138;
	wire x_2139;
	wire x_2140;
	wire x_2141;
	wire x_2142;
	wire x_2143;
	wire x_2144;
	wire x_2145;
	wire x_2146;
	wire x_2147;
	wire x_2148;
	wire x_2149;
	wire x_2150;
	wire x_2151;
	wire x_2152;
	wire x_2153;
	wire x_2154;
	wire x_2155;
	wire x_2156;
	wire x_2157;
	wire x_2158;
	wire x_2159;
	wire x_2160;
	wire x_2161;
	wire x_2162;
	wire x_2163;
	wire x_2164;
	wire x_2165;
	wire x_2166;
	wire x_2167;
	wire x_2168;
	wire x_2169;
	wire x_2170;
	wire x_2171;
	wire x_2172;
	wire x_2173;
	wire x_2174;
	wire x_2175;
	wire x_2176;
	wire x_2177;
	wire x_2178;
	wire x_2179;
	wire x_2180;
	wire x_2181;
	wire x_2182;
	wire x_2183;
	wire x_2184;
	wire x_2185;
	wire x_2186;
	wire x_2187;
	wire x_2188;
	wire x_2189;
	wire x_2190;
	wire x_2191;
	wire x_2192;
	wire x_2193;
	wire x_2194;
	wire x_2195;
	wire x_2196;
	wire x_2197;
	wire x_2198;
	wire x_2199;
	wire x_2200;
	wire x_2201;
	wire x_2202;
	wire x_2203;
	wire x_2204;
	wire x_2205;
	wire x_2206;
	wire x_2207;
	wire x_2208;
	wire x_2209;
	wire x_2210;
	wire x_2211;
	wire x_2212;
	wire x_2213;
	wire x_2214;
	wire x_2215;
	wire x_2216;
	wire x_2217;
	wire x_2218;
	wire x_2219;
	wire x_2220;
	wire x_2221;
	wire x_2222;
	wire x_2223;
	wire x_2224;
	wire x_2225;
	wire x_2226;
	wire x_2227;
	wire x_2228;
	wire x_2229;
	wire x_2230;
	wire x_2231;
	wire x_2232;
	wire x_2233;
	wire x_2234;
	wire x_2235;
	wire x_2236;
	wire x_2237;
	wire x_2238;
	wire x_2239;
	wire x_2240;
	wire x_2241;
	wire x_2242;
	wire x_2243;
	wire x_2244;
	wire x_2245;
	wire x_2246;
	wire x_2247;
	wire x_2248;
	wire x_2249;
	wire x_2250;
	wire x_2251;
	wire x_2252;
	wire x_2253;
	wire x_2254;
	wire x_2255;
	wire x_2256;
	wire x_2257;
	wire x_2258;
	wire x_2259;
	wire x_2260;
	wire x_2261;
	wire x_2262;
	wire x_2263;
	wire x_2264;
	wire x_2265;
	wire x_2266;
	wire x_2267;
	wire x_2268;
	wire x_2269;
	wire x_2270;
	wire x_2271;
	wire x_2272;
	wire x_2273;
	wire x_2274;
	wire x_2275;
	wire x_2276;
	wire x_2277;
	wire x_2278;
	wire x_2279;
	wire x_2280;
	wire x_2281;
	wire x_2282;
	wire x_2283;
	wire x_2284;
	wire x_2285;
	wire x_2286;
	wire x_2287;
	wire x_2288;
	wire x_2289;
	wire x_2290;
	wire x_2291;
	wire x_2292;
	wire x_2293;
	wire x_2294;
	wire x_2295;
	wire x_2296;
	wire x_2297;
	wire x_2298;
	wire x_2299;
	wire x_2300;
	wire x_2301;
	wire x_2302;
	wire x_2303;
	wire x_2304;
	wire x_2305;
	wire x_2306;
	wire x_2307;
	wire x_2308;
	wire x_2309;
	wire x_2310;
	wire x_2311;
	wire x_2312;
	wire x_2313;
	wire x_2314;
	wire x_2315;
	wire x_2316;
	wire x_2317;
	wire x_2318;
	wire x_2319;
	wire x_2320;
	wire x_2321;
	wire x_2322;
	wire x_2323;
	wire x_2324;
	wire x_2325;
	wire x_2326;
	wire x_2327;
	wire x_2328;
	wire x_2329;
	wire x_2330;
	wire x_2331;
	wire x_2332;
	wire x_2333;
	wire x_2334;
	wire x_2335;
	wire x_2336;
	wire x_2337;
	wire x_2338;
	wire x_2339;
	wire x_2340;
	wire x_2341;
	wire x_2342;
	wire x_2343;
	wire x_2344;
	wire x_2345;
	wire x_2346;
	wire x_2347;
	wire x_2348;
	wire x_2349;
	wire x_2350;
	wire x_2351;
	wire x_2352;
	wire x_2353;
	wire x_2354;
	wire x_2355;
	wire x_2356;
	wire x_2357;
	wire x_2358;
	wire x_2359;
	wire x_2360;
	wire x_2361;
	wire x_2362;
	wire x_2363;
	wire x_2364;
	wire x_2365;
	wire x_2366;
	wire x_2367;
	wire x_2368;
	wire x_2369;
	wire x_2370;
	wire x_2371;
	wire x_2372;
	wire x_2373;
	wire x_2374;
	wire x_2375;
	wire x_2376;
	wire x_2377;
	wire x_2378;
	wire x_2379;
	wire x_2380;
	wire x_2381;
	wire x_2382;
	wire x_2383;
	wire x_2384;
	wire x_2385;
	wire x_2386;
	wire x_2387;
	wire x_2388;
	wire x_2389;
	wire x_2390;
	wire x_2391;
	wire x_2392;
	wire x_2393;
	wire x_2394;
	wire x_2395;
	wire x_2396;
	wire x_2397;
	wire x_2398;
	wire x_2399;
	wire x_2400;
	wire x_2401;
	wire x_2402;
	wire x_2403;
	wire x_2404;
	wire x_2405;
	wire x_2406;
	wire x_2407;
	wire x_2408;
	wire x_2409;
	wire x_2410;
	wire x_2411;
	wire x_2412;
	wire x_2413;
	wire x_2414;
	wire x_2415;
	wire x_2416;
	wire x_2417;
	wire x_2418;
	wire x_2419;
	wire x_2420;
	wire x_2421;
	wire x_2422;
	wire x_2423;
	wire x_2424;
	wire x_2425;
	wire x_2426;
	wire x_2427;
	wire x_2428;
	wire x_2429;
	wire x_2430;
	wire x_2431;
	wire x_2432;
	wire x_2433;
	wire x_2434;
	wire x_2435;
	wire x_2436;
	wire x_2437;
	wire x_2438;
	wire x_2439;
	wire x_2440;
	wire x_2441;
	wire x_2442;
	wire x_2443;
	wire x_2444;
	wire x_2445;
	wire x_2446;
	wire x_2447;
	wire x_2448;
	wire x_2449;
	wire x_2450;
	wire x_2451;
	wire x_2452;
	wire x_2453;
	wire x_2454;
	wire x_2455;
	wire x_2456;
	wire x_2457;
	wire x_2458;
	wire x_2459;
	wire x_2460;
	wire x_2461;
	wire x_2462;
	wire x_2463;
	wire x_2464;
	wire x_2465;
	wire x_2466;
	wire x_2467;
	wire x_2468;
	wire x_2469;
	wire x_2470;
	wire x_2471;
	wire x_2472;
	wire x_2473;
	wire x_2474;
	wire x_2475;
	wire x_2476;
	wire x_2477;
	wire x_2478;
	wire x_2479;
	wire x_2480;
	wire x_2481;
	wire x_2482;
	wire x_2483;
	wire x_2484;
	wire x_2485;
	wire x_2486;
	wire x_2487;
	wire x_2488;
	wire x_2489;
	wire x_2490;
	wire x_2491;
	wire x_2492;
	wire x_2493;
	wire x_2494;
	wire x_2495;
	wire x_2496;
	wire x_2497;
	wire x_2498;
	wire x_2499;
	wire x_2500;
	wire x_2501;
	wire x_2502;
	wire x_2503;
	wire x_2504;
	wire x_2505;
	wire x_2506;
	wire x_2507;
	wire x_2508;
	wire x_2509;
	wire x_2510;
	wire x_2511;
	wire x_2512;
	wire x_2513;
	wire x_2514;
	wire x_2515;
	wire x_2516;
	wire x_2517;
	wire x_2518;
	wire x_2519;
	wire x_2520;
	wire x_2521;
	wire x_2522;
	wire x_2523;
	wire x_2524;
	wire x_2525;
	wire x_2526;
	wire x_2527;
	wire x_2528;
	wire x_2529;
	wire x_2530;
	wire x_2531;
	wire x_2532;
	wire x_2533;
	wire x_2534;
	wire x_2535;
	wire x_2536;
	wire x_2537;
	wire x_2538;
	wire x_2539;
	wire x_2540;
	wire x_2541;
	wire x_2542;
	wire x_2543;
	wire x_2544;
	wire x_2545;
	wire x_2546;
	wire x_2547;
	wire x_2548;
	wire x_2549;
	wire x_2550;
	wire x_2551;
	wire x_2552;
	wire x_2553;
	wire x_2554;
	wire x_2555;
	wire x_2556;
	wire x_2557;
	wire x_2558;
	wire x_2559;
	wire x_2560;
	wire x_2561;
	wire x_2562;
	wire x_2563;
	wire x_2564;
	wire x_2565;
	wire x_2566;
	wire x_2567;
	wire x_2568;
	wire x_2569;
	wire x_2570;
	wire x_2571;
	wire x_2572;
	wire x_2573;
	wire x_2574;
	wire x_2575;
	wire x_2576;
	wire x_2577;
	wire x_2578;
	wire x_2579;
	wire x_2580;
	wire x_2581;
	wire x_2582;
	wire x_2583;
	wire x_2584;
	wire x_2585;
	wire x_2586;
	wire x_2587;
	wire x_2588;
	wire x_2589;
	wire x_2590;
	wire x_2591;
	wire x_2592;
	wire x_2593;
	wire x_2594;
	wire x_2595;
	wire x_2596;
	wire x_2597;
	wire x_2598;
	wire x_2599;
	wire x_2600;
	wire x_2601;
	wire x_2602;
	wire x_2603;
	wire x_2604;
	wire x_2605;
	wire x_2606;
	wire x_2607;
	wire x_2608;
	wire x_2609;
	wire x_2610;
	wire x_2611;
	wire x_2612;
	wire x_2613;
	wire x_2614;
	wire x_2615;
	wire x_2616;
	wire x_2617;
	wire x_2618;
	wire x_2619;
	wire x_2620;
	wire x_2621;
	wire x_2622;
	wire x_2623;
	wire x_2624;
	wire x_2625;
	wire x_2626;
	wire x_2627;
	wire x_2628;
	wire x_2629;
	wire x_2630;
	wire x_2631;
	wire x_2632;
	wire x_2633;
	wire x_2634;
	wire x_2635;
	wire x_2636;
	wire x_2637;
	wire x_2638;
	wire x_2639;
	wire x_2640;
	wire x_2641;
	wire x_2642;
	wire x_2643;
	wire x_2644;
	wire x_2645;
	wire x_2646;
	wire x_2647;
	wire x_2648;
	wire x_2649;
	wire x_2650;
	wire x_2651;
	wire x_2652;
	wire x_2653;
	wire x_2654;
	wire x_2655;
	wire x_2656;
	wire x_2657;
	wire x_2658;
	wire x_2659;
	wire x_2660;
	wire x_2661;
	wire x_2662;
	wire x_2663;
	wire x_2664;
	wire x_2665;
	wire x_2666;
	wire x_2667;
	wire x_2668;
	wire x_2669;
	wire x_2670;
	wire x_2671;
	wire x_2672;
	wire x_2673;
	wire x_2674;
	wire x_2675;
	wire x_2676;
	wire x_2677;
	wire x_2678;
	wire x_2679;
	wire x_2680;
	wire x_2681;
	wire x_2682;
	wire x_2683;
	wire x_2684;
	wire x_2685;
	wire x_2686;
	wire x_2687;
	wire x_2688;
	wire x_2689;
	wire x_2690;
	wire x_2691;
	wire x_2692;
	wire x_2693;
	wire x_2694;
	wire x_2695;
	wire x_2696;
	wire x_2697;
	wire x_2698;
	wire x_2699;
	wire x_2700;
	wire x_2701;
	wire x_2702;
	wire x_2703;
	wire x_2704;
	wire x_2705;
	wire x_2706;
	wire x_2707;
	wire x_2708;
	wire x_2709;
	wire x_2710;
	wire x_2711;
	wire x_2712;
	wire x_2713;
	wire x_2714;
	wire x_2715;
	wire x_2716;
	wire x_2717;
	wire x_2718;
	wire x_2719;
	wire x_2720;
	wire x_2721;
	wire x_2722;
	wire x_2723;
	wire x_2724;
	wire x_2725;
	wire x_2726;
	wire x_2727;
	wire x_2728;
	wire x_2729;
	wire x_2730;
	wire x_2731;
	wire x_2732;
	wire x_2733;
	wire x_2734;
	wire x_2735;
	wire x_2736;
	wire x_2737;
	wire x_2738;
	wire x_2739;
	wire x_2740;
	wire x_2741;
	wire x_2742;
	wire x_2743;
	wire x_2744;
	wire x_2745;
	wire x_2746;
	wire x_2747;
	wire x_2748;
	wire x_2749;
	wire x_2750;
	wire x_2751;
	wire x_2752;
	wire x_2753;
	wire x_2754;
	wire x_2755;
	wire x_2756;
	wire x_2757;
	wire x_2758;
	wire x_2759;
	wire x_2760;
	wire x_2761;
	wire x_2762;
	wire x_2763;
	wire x_2764;
	wire x_2765;
	wire x_2766;
	wire x_2767;
	wire x_2768;
	wire x_2769;
	wire x_2770;
	wire x_2771;
	wire x_2772;
	wire x_2773;
	wire x_2774;
	wire x_2775;
	wire x_2776;
	wire x_2777;
	wire x_2778;
	wire x_2779;
	wire x_2780;
	wire x_2781;
	wire x_2782;
	wire x_2783;
	wire x_2784;
	wire x_2785;
	wire x_2786;
	wire x_2787;
	wire x_2788;
	wire x_2789;
	wire x_2790;
	wire x_2791;
	wire x_2792;
	wire x_2793;
	wire x_2794;
	wire x_2795;
	wire x_2796;
	wire x_2797;
	wire x_2798;
	wire x_2799;
	wire x_2800;
	wire x_2801;
	wire x_2802;
	wire x_2803;
	wire x_2804;
	wire x_2805;
	wire x_2806;
	wire x_2807;
	wire x_2808;
	wire x_2809;
	wire x_2810;
	wire x_2811;
	wire x_2812;
	wire x_2813;
	wire x_2814;
	wire x_2815;
	wire x_2816;
	wire x_2817;
	wire x_2818;
	wire x_2819;
	wire x_2820;
	wire x_2821;
	wire x_2822;
	wire x_2823;
	wire x_2824;
	wire x_2825;
	wire x_2826;
	wire x_2827;
	wire x_2828;
	wire x_2829;
	wire x_2830;
	wire x_2831;
	wire x_2832;
	wire x_2833;
	wire x_2834;
	wire x_2835;
	wire x_2836;
	wire x_2837;
	wire x_2838;
	wire x_2839;
	wire x_2840;
	wire x_2841;
	wire x_2842;
	wire x_2843;
	wire x_2844;
	wire x_2845;
	wire x_2846;
	wire x_2847;
	wire x_2848;
	wire x_2849;
	wire x_2850;
	wire x_2851;
	wire x_2852;
	wire x_2853;
	wire x_2854;
	wire x_2855;
	wire x_2856;
	wire x_2857;
	wire x_2858;
	wire x_2859;
	wire x_2860;
	wire x_2861;
	wire x_2862;
	wire x_2863;
	wire x_2864;
	wire x_2865;
	wire x_2866;
	wire x_2867;
	wire x_2868;
	wire x_2869;
	wire x_2870;
	wire x_2871;
	wire x_2872;
	wire x_2873;
	wire x_2874;
	wire x_2875;
	wire x_2876;
	wire x_2877;
	wire x_2878;
	wire x_2879;
	wire x_2880;
	wire x_2881;
	wire x_2882;
	wire x_2883;
	wire x_2884;
	wire x_2885;
	wire x_2886;
	wire x_2887;
	wire x_2888;
	wire x_2889;
	wire x_2890;
	wire x_2891;
	wire x_2892;
	wire x_2893;
	wire x_2894;
	wire x_2895;
	wire x_2896;
	wire x_2897;
	wire x_2898;
	wire x_2899;
	wire x_2900;
	wire x_2901;
	wire x_2902;
	wire x_2903;
	wire x_2904;
	wire x_2905;
	wire x_2906;
	wire x_2907;
	wire x_2908;
	wire x_2909;
	wire x_2910;
	wire x_2911;
	wire x_2912;
	wire x_2913;
	wire x_2914;
	wire x_2915;
	wire x_2916;
	wire x_2917;
	wire x_2918;
	wire x_2919;
	wire x_2920;
	wire x_2921;
	wire x_2922;
	wire x_2923;
	wire x_2924;
	wire x_2925;
	wire x_2926;
	wire x_2927;
	wire x_2928;
	wire x_2929;
	wire x_2930;
	wire x_2931;
	wire x_2932;
	wire x_2933;
	wire x_2934;
	wire x_2935;
	wire x_2936;
	wire x_2937;
	wire x_2938;
	wire x_2939;
	wire x_2940;
	wire x_2941;
	wire x_2942;
	wire x_2943;
	wire x_2944;
	wire x_2945;
	wire x_2946;
	wire x_2947;
	wire x_2948;
	wire x_2949;
	wire x_2950;
	wire x_2951;
	wire x_2952;
	wire x_2953;
	wire x_2954;
	wire x_2955;
	wire x_2956;
	wire x_2957;
	wire x_2958;
	wire x_2959;
	wire x_2960;
	wire x_2961;
	wire x_2962;
	wire x_2963;
	wire x_2964;
	wire x_2965;
	wire x_2966;
	wire x_2967;
	wire x_2968;
	wire x_2969;
	wire x_2970;
	wire x_2971;
	wire x_2972;
	wire x_2973;
	wire x_2974;
	wire x_2975;
	wire x_2976;
	wire x_2977;
	wire x_2978;
	wire x_2979;
	wire x_2980;
	wire x_2981;
	wire x_2982;
	wire x_2983;
	wire x_2984;
	wire x_2985;
	wire x_2986;
	wire x_2987;
	wire x_2988;
	wire x_2989;
	wire x_2990;
	wire x_2991;
	wire x_2992;
	wire x_2993;
	wire x_2994;
	wire x_2995;
	wire x_2996;
	wire x_2997;
	wire x_2998;
	wire x_2999;
	wire x_3000;
	wire x_3001;
	wire x_3002;
	wire x_3003;
	wire x_3004;
	wire x_3005;
	wire x_3006;
	wire x_3007;
	wire x_3008;
	wire x_3009;
	wire x_3010;
	wire x_3011;
	wire x_3012;
	wire x_3013;
	wire x_3014;
	wire x_3015;
	wire x_3016;
	wire x_3017;
	wire x_3018;
	wire x_3019;
	wire x_3020;
	wire x_3021;
	wire x_3022;
	wire x_3023;
	wire x_3024;
	wire x_3025;
	wire x_3026;
	wire x_3027;
	wire x_3028;
	wire x_3029;
	wire x_3030;
	wire x_3031;
	wire x_3032;
	wire x_3033;
	wire x_3034;
	wire x_3035;
	wire x_3036;
	wire x_3037;
	wire x_3038;
	wire x_3039;
	wire x_3040;
	wire x_3041;
	wire x_3042;
	wire x_3043;
	wire x_3044;
	wire x_3045;
	wire x_3046;
	wire x_3047;
	wire x_3048;
	wire x_3049;
	wire x_3050;
	wire x_3051;
	wire x_3052;
	wire x_3053;
	wire x_3054;
	wire x_3055;
	wire x_3056;
	wire x_3057;
	wire x_3058;
	wire x_3059;
	wire x_3060;
	wire x_3061;
	wire x_3062;
	wire x_3063;
	wire x_3064;
	wire x_3065;
	wire x_3066;
	wire x_3067;
	wire x_3068;
	wire x_3069;
	wire x_3070;
	wire x_3071;
	wire x_3072;
	wire x_3073;
	wire x_3074;
	wire x_3075;
	wire x_3076;
	wire x_3077;
	wire x_3078;
	wire x_3079;
	wire x_3080;
	wire x_3081;
	wire x_3082;
	wire x_3083;
	wire x_3084;
	wire x_3085;
	wire x_3086;
	wire x_3087;
	wire x_3088;
	wire x_3089;
	wire x_3090;
	wire x_3091;
	wire x_3092;
	wire x_3093;
	wire x_3094;
	wire x_3095;
	wire x_3096;
	wire x_3097;
	wire x_3098;
	wire x_3099;
	wire x_3100;
	wire x_3101;
	wire x_3102;
	wire x_3103;
	wire x_3104;
	wire x_3105;
	wire x_3106;
	wire x_3107;
	wire x_3108;
	wire x_3109;
	wire x_3110;
	wire x_3111;
	wire x_3112;
	wire x_3113;
	wire x_3114;
	wire x_3115;
	wire x_3116;
	wire x_3117;
	wire x_3118;
	wire x_3119;
	wire x_3120;
	wire x_3121;
	wire x_3122;
	wire x_3123;
	wire x_3124;
	wire x_3125;
	wire x_3126;
	wire x_3127;
	wire x_3128;
	wire x_3129;
	wire x_3130;
	wire x_3131;
	wire x_3132;
	wire x_3133;
	wire x_3134;
	wire x_3135;
	wire x_3136;
	wire x_3137;
	wire x_3138;
	wire x_3139;
	wire x_3140;
	wire x_3141;
	wire x_3142;
	wire x_3143;
	wire x_3144;
	wire x_3145;
	wire x_3146;
	wire x_3147;
	wire x_3148;
	wire x_3149;
	wire x_3150;
	wire x_3151;
	wire x_3152;
	wire x_3153;
	wire x_3154;
	wire x_3155;
	wire x_3156;
	wire x_3157;
	wire x_3158;
	wire x_3159;
	wire x_3160;
	wire x_3161;
	wire x_3162;
	wire x_3163;
	wire x_3164;
	wire x_3165;
	wire x_3166;
	wire x_3167;
	wire x_3168;
	wire x_3169;
	wire x_3170;
	wire x_3171;
	wire x_3172;
	wire x_3173;
	wire x_3174;
	wire x_3175;
	wire x_3176;
	wire x_3177;
	wire x_3178;
	wire x_3179;
	wire x_3180;
	wire x_3181;
	wire x_3182;
	wire x_3183;
	wire x_3184;
	wire x_3185;
	wire x_3186;
	wire x_3187;
	wire x_3188;
	wire x_3189;
	wire x_3190;
	wire x_3191;
	wire x_3192;
	wire x_3193;
	wire x_3194;
	wire x_3195;
	wire x_3196;
	wire x_3197;
	wire x_3198;
	wire x_3199;
	wire x_3200;
	wire x_3201;
	wire x_3202;
	wire x_3203;
	wire x_3204;
	wire x_3205;
	wire x_3206;
	wire x_3207;
	wire x_3208;
	wire x_3209;
	wire x_3210;
	wire x_3211;
	wire x_3212;
	wire x_3213;
	wire x_3214;
	wire x_3215;
	wire x_3216;
	wire x_3217;
	wire x_3218;
	wire x_3219;
	wire x_3220;
	wire x_3221;
	wire x_3222;
	wire x_3223;
	wire x_3224;
	wire x_3225;
	wire x_3226;
	wire x_3227;
	wire x_3228;
	wire x_3229;
	wire x_3230;
	wire x_3231;
	wire x_3232;
	wire x_3233;
	wire x_3234;
	wire x_3235;
	wire x_3236;
	wire x_3237;
	wire x_3238;
	wire x_3239;
	wire x_3240;
	wire x_3241;
	wire x_3242;
	wire x_3243;
	wire x_3244;
	wire x_3245;
	wire x_3246;
	wire x_3247;
	wire x_3248;
	wire x_3249;
	wire x_3250;
	wire x_3251;
	wire x_3252;
	wire x_3253;
	wire x_3254;
	wire x_3255;
	wire x_3256;
	wire x_3257;
	wire x_3258;
	wire x_3259;
	output o_1;
	assign x_1630 = (v_67 | v_17);
	assign x_1629 = (v_67 | v_12);
	assign x_1628 = (v_68 | ~v_11);
	assign x_1627 = (v_68 | v_26);
	assign x_1626 = (v_69 | v_11);
	assign x_1625 = (v_69 | v_27);
	assign x_1623 = (v_70 | v_13);
	assign x_1624 = (v_70 | ~v_12);
	assign x_1622 = (((((((((((((((((((((v_24 | v_23)) | v_55)) | v_46)) | v_64)) | v_58)) | v_47)) | ~v_70)) | ~v_69)) | ~v_68)) | ~v_67)) | v_71);
	assign x_1620 = (v_72 | v_12);
	assign x_1621 = (v_72 | v_16);
	assign x_1619 = (v_73 | ~v_11);
	assign x_1618 = (v_73 | v_35);
	assign x_1617 = (v_74 | v_11);
	assign x_1616 = (v_74 | v_36);
	assign x_1615 = (v_75 | ~v_12);
	assign x_1614 = (v_75 | v_14);
	assign x_1613 = (((((((((((((((((((((v_32 | v_33)) | v_56)) | v_50)) | v_49)) | v_65)) | v_59)) | ~v_75)) | ~v_74)) | ~v_73)) | ~v_72)) | v_76);
	assign x_1612 = (v_77 | v_18);
	assign x_1611 = (v_77 | v_12);
	assign x_1610 = (v_78 | ~v_11);
	assign x_1609 = (v_78 | v_44);
	assign x_1607 = (v_79 | v_45);
	assign x_1608 = (v_79 | v_11);
	assign x_1606 = (v_80 | ~v_12);
	assign x_1605 = (v_80 | v_15);
	assign x_1604 = (((((((((((((((((((((v_53 | v_52)) | v_66)) | v_60)) | v_57)) | v_42)) | v_41)) | ~v_80)) | ~v_79)) | ~v_78)) | ~v_77)) | v_81);
	assign x_1603 = (v_82 | ~v_81);
	assign x_1602 = (v_82 | ~v_76);
	assign x_1601 = (v_82 | ~v_71);
	assign x_1600 = (v_83 | ~v_10);
	assign x_1599 = (v_83 | v_26);
	assign x_1597 = (v_84 | v_27);
	assign x_1598 = (v_84 | v_10);
	assign x_1596 = (v_85 | ~v_11);
	assign x_1595 = (v_85 | v_13);
	assign x_1594 = (v_86 | v_17);
	assign x_1593 = (v_86 | v_11);
	assign x_1592 = (((((((((((((((((((((v_24 | v_23)) | v_22)) | v_55)) | v_46)) | v_58)) | v_47)) | ~v_86)) | ~v_85)) | ~v_84)) | ~v_83)) | v_87);
	assign x_1591 = (v_88 | ~v_10);
	assign x_1590 = (v_88 | v_35);
	assign x_1588 = (v_89 | v_36);
	assign x_1589 = (v_89 | v_10);
	assign x_1587 = (v_90 | v_16);
	assign x_1586 = (v_90 | v_11);
	assign x_1585 = (v_91 | ~v_11);
	assign x_1584 = (v_91 | v_14);
	assign x_1583 = (((((((((((((((((((((v_32 | v_31)) | v_33)) | v_56)) | v_50)) | v_49)) | v_59)) | ~v_91)) | ~v_90)) | ~v_89)) | ~v_88)) | v_92);
	assign x_1582 = (v_93 | ~v_10);
	assign x_1581 = (v_93 | v_44);
	assign x_1579 = (v_94 | v_45);
	assign x_1580 = (v_94 | v_10);
	assign x_1578 = (v_95 | ~v_11);
	assign x_1577 = (v_95 | v_15);
	assign x_1576 = (v_96 | v_18);
	assign x_1575 = (v_96 | v_11);
	assign x_1574 = (((((((((((((((((((((v_53 | v_52)) | v_40)) | v_60)) | v_57)) | v_42)) | v_41)) | ~v_96)) | ~v_95)) | ~v_94)) | ~v_93)) | v_97);
	assign x_1572 = (v_98 | ~v_92);
	assign x_1571 = (v_98 | ~v_87);
	assign x_1573 = (v_98 | ~v_97);
	assign x_1569 = (v_99 | v_16);
	assign x_1570 = (v_99 | ~v_18);
	assign x_1568 = (v_100 | ~v_14);
	assign x_1567 = (v_100 | v_15);
	assign x_1566 = (v_101 | ~v_16);
	assign x_1565 = (v_101 | v_17);
	assign x_1564 = (v_102 | ~v_13);
	assign x_1563 = (v_102 | v_14);
	assign x_1562 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_98)) | ~v_82)) | v_103);
	assign x_1561 = (v_104 | ~v_9);
	assign x_1560 = (v_104 | v_26);
	assign x_1559 = (v_105 | v_9);
	assign x_1558 = (v_105 | v_27);
	assign x_1557 = (((((((((((((((((((((v_25 | v_24)) | v_23)) | v_21)) | v_55)) | v_46)) | v_64)) | ~v_70)) | ~v_105)) | ~v_104)) | ~v_67)) | v_106);
	assign x_1556 = (v_107 | ~v_9);
	assign x_1555 = (v_107 | v_35);
	assign x_1553 = (v_108 | v_36);
	assign x_1554 = (v_108 | v_9);
	assign x_1552 = (((((((((((((((((((((v_32 | v_30)) | v_33)) | v_34)) | v_56)) | v_49)) | v_65)) | ~v_75)) | ~v_108)) | ~v_107)) | ~v_72)) | v_109);
	assign x_1551 = (v_110 | ~v_9);
	assign x_1550 = (v_110 | v_44);
	assign x_1549 = (v_111 | v_9);
	assign x_1548 = (v_111 | v_45);
	assign x_1547 = (((((((((((((((((((((v_39 | v_52)) | v_66)) | v_43)) | v_57)) | v_42)) | v_41)) | ~v_80)) | ~v_111)) | ~v_110)) | ~v_77)) | v_112);
	assign x_1546 = (v_113 | ~v_112);
	assign x_1545 = (v_113 | ~v_109);
	assign x_1544 = (v_113 | ~v_106);
	assign x_1543 = (v_114 | ~v_9);
	assign x_1542 = (v_114 | v_13);
	assign x_1540 = (v_115 | v_17);
	assign x_1541 = (v_115 | v_9);
	assign x_1539 = (((((((((((((((((((((v_25 | v_23)) | v_22)) | v_20)) | v_48)) | v_46)) | v_47)) | ~v_115)) | ~v_114)) | ~v_84)) | ~v_83)) | v_116);
	assign x_1537 = (v_117 | v_16);
	assign x_1538 = (v_117 | v_9);
	assign x_1536 = (v_118 | ~v_9);
	assign x_1535 = (v_118 | v_14);
	assign x_1534 = (((((((((((((((((((((v_32 | v_31)) | v_29)) | v_34)) | v_50)) | v_51)) | v_49)) | ~v_118)) | ~v_117)) | ~v_89)) | ~v_88)) | v_119);
	assign x_1533 = (v_120 | v_9);
	assign x_1532 = (v_120 | v_18);
	assign x_1531 = (v_121 | ~v_9);
	assign x_1530 = (v_121 | v_15);
	assign x_1529 = (((((((((((((((((((((v_38 | v_54)) | v_53)) | v_52)) | v_43)) | v_40)) | v_41)) | ~v_121)) | ~v_120)) | ~v_94)) | ~v_93)) | v_122);
	assign x_1528 = (v_123 | ~v_122);
	assign x_1527 = (v_123 | ~v_119);
	assign x_1526 = (v_123 | ~v_116);
	assign x_1525 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_123)) | ~v_113)) | v_124);
	assign x_1524 = (((((((((((((((((((((v_32 | v_33)) | v_34)) | v_56)) | v_50)) | v_49)) | v_65)) | ~v_75)) | ~v_89)) | ~v_88)) | ~v_72)) | v_125);
	assign x_1523 = (((((((((((((((((((((v_53 | v_52)) | v_66)) | v_43)) | v_57)) | v_42)) | v_41)) | ~v_80)) | ~v_94)) | ~v_93)) | ~v_77)) | v_126);
	assign x_1522 = (((((((((((((((((((((v_25 | v_24)) | v_23)) | v_55)) | v_46)) | v_64)) | v_47)) | ~v_70)) | ~v_84)) | ~v_83)) | ~v_67)) | v_127);
	assign x_1521 = (v_128 | ~v_127);
	assign x_1520 = (v_128 | ~v_126);
	assign x_1519 = (v_128 | ~v_125);
	assign x_1518 = (((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_128)) | v_129);
	assign x_1517 = (v_130 | ~v_129);
	assign x_1515 = (v_130 | ~v_103);
	assign x_1516 = (v_130 | ~v_124);
	assign x_1514 = (v_131 | ~v_12);
	assign x_1513 = (v_131 | v_26);
	assign x_1512 = (v_132 | v_12);
	assign x_1511 = (v_132 | v_27);
	assign x_1510 = (((((((((((((((((((((v_25 | v_24)) | v_22)) | v_20)) | v_61)) | v_46)) | v_47)) | ~v_115)) | ~v_132)) | ~v_114)) | ~v_131)) | v_133);
	assign x_1508 = (v_134 | v_35);
	assign x_1509 = (v_134 | ~v_12);
	assign x_1507 = (v_135 | v_12);
	assign x_1506 = (v_135 | v_36);
	assign x_1505 = (((((((((((((((((((((v_31 | v_29)) | v_33)) | v_34)) | v_50)) | v_49)) | v_62)) | ~v_118)) | ~v_117)) | ~v_135)) | ~v_134)) | v_136);
	assign x_1504 = (v_137 | ~v_12);
	assign x_1503 = (v_137 | v_44);
	assign x_1502 = (v_138 | v_12);
	assign x_1501 = (v_138 | v_45);
	assign x_1500 = (((((((((((((((((((((v_38 | v_53)) | v_52)) | v_43)) | v_40)) | v_63)) | v_42)) | ~v_121)) | ~v_120)) | ~v_138)) | ~v_137)) | v_139);
	assign x_1499 = (v_140 | ~v_139);
	assign x_1498 = (v_140 | ~v_136);
	assign x_1497 = (v_140 | ~v_133);
	assign x_1496 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_140)) | ~v_130)) | v_141);
	assign x_1495 = (((((((((((((((((((((v_25 | v_22)) | v_55)) | v_61)) | v_48)) | v_46)) | v_47)) | ~v_86)) | ~v_85)) | ~v_132)) | ~v_131)) | v_142);
	assign x_1494 = (((((((((((((((((((((v_31 | v_34)) | v_56)) | v_50)) | v_51)) | v_49)) | v_62)) | ~v_91)) | ~v_90)) | ~v_135)) | ~v_134)) | v_143);
	assign x_1493 = (((((((((((((((((((((v_54 | v_53)) | v_52)) | v_43)) | v_40)) | v_63)) | v_57)) | ~v_138)) | ~v_137)) | ~v_96)) | ~v_95)) | v_144);
	assign x_1492 = (v_145 | ~v_144);
	assign x_1491 = (v_145 | ~v_143);
	assign x_1490 = (v_145 | ~v_142);
	assign x_1489 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_145)) | ~v_128)) | v_146);
	assign x_1488 = (((((((((((((((((((((v_25 | v_24)) | v_23)) | v_22)) | v_21)) | v_55)) | v_46)) | ~v_86)) | ~v_85)) | ~v_105)) | ~v_104)) | v_147);
	assign x_1487 = (((((((((((((((((((((v_32 | v_31)) | v_30)) | v_33)) | v_34)) | v_56)) | v_49)) | ~v_91)) | ~v_90)) | ~v_108)) | ~v_107)) | v_148);
	assign x_1486 = (((((((((((((((((((((v_39 | v_52)) | v_43)) | v_40)) | v_57)) | v_42)) | v_41)) | ~v_96)) | ~v_95)) | ~v_111)) | ~v_110)) | v_149);
	assign x_1485 = (v_150 | ~v_149);
	assign x_1483 = (v_150 | ~v_147);
	assign x_1484 = (v_150 | ~v_148);
	assign x_1482 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_150)) | ~v_123)) | v_151);
	assign x_1481 = (((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_98)) | v_152);
	assign x_1480 = (v_153 | ~v_152);
	assign x_1479 = (v_153 | ~v_151);
	assign x_1478 = (v_153 | ~v_146);
	assign x_1477 = (((((((((((((((((((((v_25 | v_24)) | v_23)) | v_22)) | v_20)) | v_46)) | v_47)) | ~v_115)) | ~v_69)) | ~v_68)) | ~v_114)) | v_154);
	assign x_1476 = (((((((((((((((((((((v_32 | v_31)) | v_29)) | v_33)) | v_34)) | v_50)) | v_49)) | ~v_118)) | ~v_117)) | ~v_74)) | ~v_73)) | v_155);
	assign x_1475 = (((((((((((((((((((((v_38 | v_53)) | v_52)) | v_43)) | v_40)) | v_42)) | v_41)) | ~v_121)) | ~v_120)) | ~v_79)) | ~v_78)) | v_156);
	assign x_1474 = (v_157 | ~v_156);
	assign x_1473 = (v_157 | ~v_155);
	assign x_1472 = (v_157 | ~v_154);
	assign x_1471 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_157)) | ~v_153)) | v_158);
	assign x_1470 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_140)) | ~v_128)) | v_159);
	assign x_1469 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_98)) | ~v_157)) | v_160);
	assign x_1468 = (((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_123)) | v_161);
	assign x_1467 = (v_162 | ~v_161);
	assign x_1466 = (v_162 | ~v_160);
	assign x_1464 = (v_162 | ~v_158);
	assign x_1463 = (v_162 | ~v_141);
	assign x_1465 = (v_162 | ~v_159);
	assign x_1462 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_145)) | ~v_157)) | v_163);
	assign x_1461 = (v_164 | ~v_10);
	assign x_1460 = (v_164 | v_14);
	assign x_1459 = (v_165 | v_16);
	assign x_1458 = (v_165 | v_10);
	assign x_1457 = (((((((((((((((((((((v_31 | v_33)) | v_34)) | v_56)) | v_50)) | v_49)) | v_62)) | ~v_165)) | ~v_164)) | ~v_135)) | ~v_134)) | v_166);
	assign x_1456 = (v_167 | ~v_10);
	assign x_1455 = (v_167 | v_15);
	assign x_1454 = (v_168 | v_18);
	assign x_1453 = (v_168 | v_10);
	assign x_1452 = (((((((((((((((((((((v_53 | v_52)) | v_43)) | v_40)) | v_63)) | v_57)) | v_42)) | ~v_138)) | ~v_137)) | ~v_168)) | ~v_167)) | v_169);
	assign x_1451 = (v_170 | ~v_10);
	assign x_1450 = (v_170 | v_13);
	assign x_1449 = (v_171 | v_17);
	assign x_1448 = (v_171 | v_10);
	assign x_1447 = (((((((((((((((((((((v_25 | v_24)) | v_22)) | v_55)) | v_61)) | v_46)) | v_47)) | ~v_171)) | ~v_132)) | ~v_170)) | ~v_131)) | v_172);
	assign x_1446 = (v_173 | ~v_172);
	assign x_1444 = (v_173 | ~v_166);
	assign x_1445 = (v_173 | ~v_169);
	assign x_1443 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_173)) | ~v_123)) | v_174);
	assign x_1442 = (((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_140)) | v_175);
	assign x_1441 = (v_176 | ~v_175);
	assign x_1440 = (v_176 | ~v_174);
	assign x_1439 = (v_176 | ~v_163);
	assign x_1438 = (((((((((((((((((((((v_24 | v_23)) | v_22)) | v_21)) | v_55)) | v_46)) | v_58)) | ~v_171)) | ~v_105)) | ~v_104)) | ~v_170)) | v_177);
	assign x_1437 = (((((((((((((((((((((v_32 | v_31)) | v_30)) | v_33)) | v_56)) | v_49)) | v_59)) | ~v_165)) | ~v_108)) | ~v_107)) | ~v_164)) | v_178);
	assign x_1436 = (((((((((((((((((((((v_39 | v_52)) | v_40)) | v_60)) | v_57)) | v_42)) | v_41)) | ~v_111)) | ~v_110)) | ~v_168)) | ~v_167)) | v_179);
	assign x_1435 = (v_180 | ~v_179);
	assign x_1434 = (v_180 | ~v_178);
	assign x_1433 = (v_180 | ~v_177);
	assign x_1432 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_180)) | ~v_176)) | v_181);
	assign x_1431 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_140)) | ~v_150)) | v_182);
	assign x_1430 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_173)) | ~v_98)) | v_183);
	assign x_1429 = (((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_145)) | v_184);
	assign x_1428 = (v_185 | ~v_184);
	assign x_1426 = (v_185 | ~v_182);
	assign x_1427 = (v_185 | ~v_183);
	assign x_1425 = (((((((((((((((((((((v_25 | v_23)) | v_22)) | v_55)) | v_48)) | v_46)) | v_47)) | ~v_171)) | ~v_69)) | ~v_68)) | ~v_170)) | v_186);
	assign x_1424 = (((((((((((((((((((((v_32 | v_31)) | v_34)) | v_56)) | v_50)) | v_51)) | v_49)) | ~v_165)) | ~v_74)) | ~v_73)) | ~v_164)) | v_187);
	assign x_1423 = (((((((((((((((((((((v_54 | v_53)) | v_52)) | v_43)) | v_40)) | v_57)) | v_41)) | ~v_79)) | ~v_78)) | ~v_168)) | ~v_167)) | v_188);
	assign x_1422 = (v_189 | ~v_188);
	assign x_1421 = (v_189 | ~v_187);
	assign x_1420 = (v_189 | ~v_186);
	assign x_1419 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_189)) | ~v_185)) | v_190);
	assign x_1418 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_189)) | ~v_145)) | v_191);
	assign x_1417 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_180)) | ~v_140)) | v_192);
	assign x_1416 = (((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_173)) | v_193);
	assign x_1415 = (v_194 | ~v_193);
	assign x_1413 = (v_194 | ~v_191);
	assign x_1412 = (v_194 | ~v_190);
	assign x_1411 = (v_194 | ~v_181);
	assign x_1414 = (v_194 | ~v_192);
	assign x_1410 = (((~v_194 | ~v_162)) | v_195);
	assign x_1409 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_189)) | ~v_128)) | v_196);
	assign x_1408 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_157)) | ~v_113)) | v_197);
	assign x_1407 = (((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_82)) | v_198);
	assign x_1406 = (v_199 | ~v_198);
	assign x_1405 = (v_199 | ~v_197);
	assign x_1404 = (v_199 | ~v_196);
	assign x_1403 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_140)) | ~v_199)) | v_200);
	assign x_1402 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_173)) | ~v_82)) | v_201);
	assign x_1401 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_180)) | ~v_157)) | v_202);
	assign x_1400 = (((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_189)) | v_203);
	assign x_1399 = (v_204 | ~v_203);
	assign x_1398 = (v_204 | ~v_202);
	assign x_1397 = (v_204 | ~v_201);
	assign x_1396 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_123)) | ~v_204)) | v_205);
	assign x_1395 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_189)) | ~v_123)) | v_206);
	assign x_1394 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_140)) | ~v_82)) | v_207);
	assign x_1393 = (((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_157)) | v_208);
	assign x_1392 = (v_209 | ~v_208);
	assign x_1390 = (v_209 | ~v_206);
	assign x_1389 = (v_209 | ~v_205);
	assign x_1391 = (v_209 | ~v_207);
	assign x_1388 = (v_209 | ~v_200);
	assign x_1387 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_150)) | ~v_176)) | v_210);
	assign x_1386 = (v_211 | ~v_193);
	assign x_1384 = (v_211 | ~v_191);
	assign x_1385 = (v_211 | ~v_192);
	assign x_1383 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_211)) | ~v_98)) | v_212);
	assign x_1381 = (v_213 | ~v_183);
	assign x_1380 = (v_213 | ~v_182);
	assign x_1378 = (v_213 | ~v_210);
	assign x_1382 = (v_213 | ~v_184);
	assign x_1379 = (v_213 | ~v_212);
	assign x_1377 = (((~v_213 | ~v_209)) | v_214);
	assign x_1376 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_185)) | ~v_157)) | v_215);
	assign x_1375 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_211)) | ~v_123)) | v_216);
	assign x_1374 = (v_217 | ~v_175);
	assign x_1373 = (v_217 | ~v_174);
	assign x_1372 = (v_217 | ~v_163);
	assign x_1371 = (v_217 | ~v_216);
	assign x_1370 = (v_217 | ~v_215);
	assign x_1368 = (v_217 | ~v_195);
	assign x_1369 = (v_217 | ~v_214);
	assign x_1367 = (((((((((~v_9 | ~v_10)) | ~v_11)) | ~v_12)) | ~v_217)) | v_218);
	assign x_1365 = (v_219 | v_12);
	assign x_1364 = (v_219 | v_11);
	assign x_1366 = (v_219 | v_9);
	assign x_1363 = (v_219 | v_10);
	assign x_1362 = (((~v_12 | ~v_17)) | v_220);
	assign x_1361 = (((~v_26 | v_11)) | v_221);
	assign x_1360 = (((~v_11 | ~v_27)) | v_222);
	assign x_1359 = (((~v_13 | v_12)) | v_223);
	assign x_1358 = (v_224 | ~v_23);
	assign x_1357 = (v_224 | ~v_24);
	assign x_1355 = (v_224 | ~v_47);
	assign x_1354 = (v_224 | ~v_55);
	assign x_1352 = (v_224 | ~v_64);
	assign x_1351 = (v_224 | ~v_223);
	assign x_1349 = (v_224 | ~v_221);
	assign x_1348 = (v_224 | ~v_220);
	assign x_1356 = (v_224 | ~v_46);
	assign x_1353 = (v_224 | ~v_58);
	assign x_1350 = (v_224 | ~v_222);
	assign x_1347 = (((~v_12 | ~v_16)) | v_225);
	assign x_1346 = (((~v_35 | v_11)) | v_226);
	assign x_1345 = (((~v_11 | ~v_36)) | v_227);
	assign x_1344 = (((~v_14 | v_12)) | v_228);
	assign x_1342 = (v_229 | ~v_33);
	assign x_1341 = (v_229 | ~v_49);
	assign x_1339 = (v_229 | ~v_56);
	assign x_1338 = (v_229 | ~v_59);
	assign x_1336 = (v_229 | ~v_228);
	assign x_1335 = (v_229 | ~v_227);
	assign x_1333 = (v_229 | ~v_225);
	assign x_1343 = (v_229 | ~v_32);
	assign x_1340 = (v_229 | ~v_50);
	assign x_1337 = (v_229 | ~v_65);
	assign x_1334 = (v_229 | ~v_226);
	assign x_1332 = (((~v_12 | ~v_18)) | v_230);
	assign x_1331 = (((v_11 | ~v_44)) | v_231);
	assign x_1330 = (((~v_11 | ~v_45)) | v_232);
	assign x_1329 = (((~v_15 | v_12)) | v_233);
	assign x_1327 = (v_234 | ~v_42);
	assign x_1326 = (v_234 | ~v_52);
	assign x_1324 = (v_234 | ~v_57);
	assign x_1323 = (v_234 | ~v_60);
	assign x_1322 = (v_234 | ~v_66);
	assign x_1321 = (v_234 | ~v_233);
	assign x_1320 = (v_234 | ~v_232);
	assign x_1319 = (v_234 | ~v_231);
	assign x_1328 = (v_234 | ~v_41);
	assign x_1325 = (v_234 | ~v_53);
	assign x_1318 = (v_234 | ~v_230);
	assign x_1317 = (((((~v_234 | ~v_229)) | ~v_224)) | v_235);
	assign x_1316 = (((~v_26 | v_10)) | v_236);
	assign x_1315 = (((~v_10 | ~v_27)) | v_237);
	assign x_1314 = (((~v_13 | v_11)) | v_238);
	assign x_1313 = (((~v_11 | ~v_17)) | v_239);
	assign x_1311 = (v_240 | ~v_23);
	assign x_1310 = (v_240 | ~v_24);
	assign x_1309 = (v_240 | ~v_46);
	assign x_1308 = (v_240 | ~v_47);
	assign x_1307 = (v_240 | ~v_55);
	assign x_1306 = (v_240 | ~v_58);
	assign x_1304 = (v_240 | ~v_238);
	assign x_1303 = (v_240 | ~v_237);
	assign x_1312 = (v_240 | ~v_22);
	assign x_1305 = (v_240 | ~v_239);
	assign x_1302 = (v_240 | ~v_236);
	assign x_1301 = (((~v_35 | v_10)) | v_241);
	assign x_1300 = (((~v_10 | ~v_36)) | v_242);
	assign x_1299 = (((~v_11 | ~v_16)) | v_243);
	assign x_1298 = (((~v_14 | v_11)) | v_244);
	assign x_1297 = (v_245 | ~v_31);
	assign x_1296 = (v_245 | ~v_32);
	assign x_1295 = (v_245 | ~v_33);
	assign x_1294 = (v_245 | ~v_49);
	assign x_1293 = (v_245 | ~v_50);
	assign x_1291 = (v_245 | ~v_59);
	assign x_1290 = (v_245 | ~v_244);
	assign x_1288 = (v_245 | ~v_242);
	assign x_1287 = (v_245 | ~v_241);
	assign x_1292 = (v_245 | ~v_56);
	assign x_1289 = (v_245 | ~v_243);
	assign x_1286 = (((v_10 | ~v_44)) | v_246);
	assign x_1285 = (((~v_10 | ~v_45)) | v_247);
	assign x_1284 = (((~v_15 | v_11)) | v_248);
	assign x_1283 = (((~v_11 | ~v_18)) | v_249);
	assign x_1282 = (v_250 | ~v_40);
	assign x_1281 = (v_250 | ~v_41);
	assign x_1279 = (v_250 | ~v_52);
	assign x_1278 = (v_250 | ~v_53);
	assign x_1276 = (v_250 | ~v_60);
	assign x_1275 = (v_250 | ~v_249);
	assign x_1273 = (v_250 | ~v_247);
	assign x_1272 = (v_250 | ~v_246);
	assign x_1280 = (v_250 | ~v_42);
	assign x_1277 = (v_250 | ~v_57);
	assign x_1274 = (v_250 | ~v_248);
	assign x_1271 = (((((~v_250 | ~v_245)) | ~v_240)) | v_251);
	assign x_1270 = (((~v_16 | v_18)) | v_252);
	assign x_1269 = (((~v_15 | v_14)) | v_253);
	assign x_1268 = (((~v_17 | v_16)) | v_254);
	assign x_1267 = (((~v_14 | v_13)) | v_255);
	assign x_1266 = (v_256 | ~v_255);
	assign x_1265 = (v_256 | ~v_254);
	assign x_1263 = (v_256 | ~v_252);
	assign x_1262 = (v_256 | ~v_251);
	assign x_1264 = (v_256 | ~v_253);
	assign x_1261 = (v_256 | ~v_235);
	assign x_1260 = (((~v_26 | v_9)) | v_257);
	assign x_1259 = (((~v_9 | ~v_27)) | v_258);
	assign x_1258 = (v_259 | ~v_21);
	assign x_1257 = (v_259 | ~v_23);
	assign x_1256 = (v_259 | ~v_24);
	assign x_1255 = (v_259 | ~v_25);
	assign x_1253 = (v_259 | ~v_55);
	assign x_1252 = (v_259 | ~v_64);
	assign x_1250 = (v_259 | ~v_258);
	assign x_1249 = (v_259 | ~v_257);
	assign x_1254 = (v_259 | ~v_46);
	assign x_1251 = (v_259 | ~v_223);
	assign x_1248 = (v_259 | ~v_220);
	assign x_1247 = (((~v_35 | v_9)) | v_260);
	assign x_1246 = (((~v_9 | ~v_36)) | v_261);
	assign x_1245 = (v_262 | ~v_30);
	assign x_1244 = (v_262 | ~v_32);
	assign x_1243 = (v_262 | ~v_33);
	assign x_1242 = (v_262 | ~v_34);
	assign x_1240 = (v_262 | ~v_56);
	assign x_1239 = (v_262 | ~v_65);
	assign x_1237 = (v_262 | ~v_261);
	assign x_1236 = (v_262 | ~v_260);
	assign x_1241 = (v_262 | ~v_49);
	assign x_1238 = (v_262 | ~v_228);
	assign x_1235 = (v_262 | ~v_225);
	assign x_1234 = (((v_9 | ~v_44)) | v_263);
	assign x_1233 = (((~v_9 | ~v_45)) | v_264);
	assign x_1231 = (v_265 | ~v_41);
	assign x_1230 = (v_265 | ~v_42);
	assign x_1228 = (v_265 | ~v_52);
	assign x_1227 = (v_265 | ~v_57);
	assign x_1225 = (v_265 | ~v_233);
	assign x_1224 = (v_265 | ~v_264);
	assign x_1222 = (v_265 | ~v_230);
	assign x_1232 = (v_265 | ~v_39);
	assign x_1229 = (v_265 | ~v_43);
	assign x_1226 = (v_265 | ~v_66);
	assign x_1223 = (v_265 | ~v_263);
	assign x_1221 = (((((~v_265 | ~v_262)) | ~v_259)) | v_266);
	assign x_1220 = (((~v_13 | v_9)) | v_267);
	assign x_1219 = (((~v_9 | ~v_17)) | v_268);
	assign x_1218 = (v_269 | ~v_20);
	assign x_1217 = (v_269 | ~v_22);
	assign x_1215 = (v_269 | ~v_25);
	assign x_1214 = (v_269 | ~v_46);
	assign x_1212 = (v_269 | ~v_48);
	assign x_1211 = (v_269 | ~v_268);
	assign x_1209 = (v_269 | ~v_237);
	assign x_1208 = (v_269 | ~v_236);
	assign x_1216 = (v_269 | ~v_23);
	assign x_1213 = (v_269 | ~v_47);
	assign x_1210 = (v_269 | ~v_267);
	assign x_1207 = (((~v_9 | ~v_16)) | v_270);
	assign x_1206 = (((~v_14 | v_9)) | v_271);
	assign x_1205 = (v_272 | ~v_29);
	assign x_1204 = (v_272 | ~v_31);
	assign x_1202 = (v_272 | ~v_34);
	assign x_1201 = (v_272 | ~v_49);
	assign x_1199 = (v_272 | ~v_51);
	assign x_1198 = (v_272 | ~v_271);
	assign x_1196 = (v_272 | ~v_242);
	assign x_1195 = (v_272 | ~v_241);
	assign x_1203 = (v_272 | ~v_32);
	assign x_1200 = (v_272 | ~v_50);
	assign x_1197 = (v_272 | ~v_270);
	assign x_1194 = (((~v_15 | v_9)) | v_273);
	assign x_1193 = (((~v_9 | ~v_18)) | v_274);
	assign x_1192 = (v_275 | ~v_38);
	assign x_1191 = (v_275 | ~v_40);
	assign x_1189 = (v_275 | ~v_43);
	assign x_1188 = (v_275 | ~v_52);
	assign x_1186 = (v_275 | ~v_54);
	assign x_1185 = (v_275 | ~v_274);
	assign x_1183 = (v_275 | ~v_247);
	assign x_1182 = (v_275 | ~v_246);
	assign x_1190 = (v_275 | ~v_41);
	assign x_1187 = (v_275 | ~v_53);
	assign x_1184 = (v_275 | ~v_273);
	assign x_1181 = (((((~v_275 | ~v_272)) | ~v_269)) | v_276);
	assign x_1180 = (v_277 | ~v_255);
	assign x_1179 = (v_277 | ~v_254);
	assign x_1177 = (v_277 | ~v_252);
	assign x_1176 = (v_277 | ~v_276);
	assign x_1178 = (v_277 | ~v_253);
	assign x_1175 = (v_277 | ~v_266);
	assign x_1174 = (v_278 | ~v_32);
	assign x_1173 = (v_278 | ~v_33);
	assign x_1171 = (v_278 | ~v_49);
	assign x_1170 = (v_278 | ~v_50);
	assign x_1169 = (v_278 | ~v_56);
	assign x_1168 = (v_278 | ~v_65);
	assign x_1167 = (v_278 | ~v_228);
	assign x_1166 = (v_278 | ~v_242);
	assign x_1164 = (v_278 | ~v_225);
	assign x_1172 = (v_278 | ~v_34);
	assign x_1165 = (v_278 | ~v_241);
	assign x_1163 = (v_279 | ~v_41);
	assign x_1161 = (v_279 | ~v_43);
	assign x_1160 = (v_279 | ~v_52);
	assign x_1158 = (v_279 | ~v_57);
	assign x_1157 = (v_279 | ~v_66);
	assign x_1156 = (v_279 | ~v_233);
	assign x_1155 = (v_279 | ~v_247);
	assign x_1154 = (v_279 | ~v_246);
	assign x_1153 = (v_279 | ~v_230);
	assign x_1162 = (v_279 | ~v_42);
	assign x_1159 = (v_279 | ~v_53);
	assign x_1151 = (v_280 | ~v_24);
	assign x_1150 = (v_280 | ~v_25);
	assign x_1148 = (v_280 | ~v_47);
	assign x_1147 = (v_280 | ~v_55);
	assign x_1145 = (v_280 | ~v_223);
	assign x_1144 = (v_280 | ~v_237);
	assign x_1143 = (v_280 | ~v_236);
	assign x_1142 = (v_280 | ~v_220);
	assign x_1152 = (v_280 | ~v_23);
	assign x_1149 = (v_280 | ~v_46);
	assign x_1146 = (v_280 | ~v_64);
	assign x_1141 = (((((~v_280 | ~v_279)) | ~v_278)) | v_281);
	assign x_1140 = (v_282 | ~v_255);
	assign x_1138 = (v_282 | ~v_253);
	assign x_1137 = (v_282 | ~v_252);
	assign x_1139 = (v_282 | ~v_254);
	assign x_1136 = (v_282 | ~v_281);
	assign x_1135 = (((((~v_282 | ~v_277)) | ~v_256)) | v_283);
	assign x_1134 = (((~v_26 | v_12)) | v_284);
	assign x_1133 = (((~v_12 | ~v_27)) | v_285);
	assign x_1132 = (v_286 | ~v_20);
	assign x_1131 = (v_286 | ~v_22);
	assign x_1129 = (v_286 | ~v_25);
	assign x_1128 = (v_286 | ~v_46);
	assign x_1126 = (v_286 | ~v_61);
	assign x_1125 = (v_286 | ~v_268);
	assign x_1123 = (v_286 | ~v_267);
	assign x_1122 = (v_286 | ~v_284);
	assign x_1130 = (v_286 | ~v_24);
	assign x_1127 = (v_286 | ~v_47);
	assign x_1124 = (v_286 | ~v_285);
	assign x_1121 = (((~v_35 | v_12)) | v_287);
	assign x_1120 = (((~v_12 | ~v_36)) | v_288);
	assign x_1119 = (v_289 | ~v_29);
	assign x_1118 = (v_289 | ~v_31);
	assign x_1117 = (v_289 | ~v_33);
	assign x_1116 = (v_289 | ~v_34);
	assign x_1115 = (v_289 | ~v_49);
	assign x_1113 = (v_289 | ~v_62);
	assign x_1112 = (v_289 | ~v_271);
	assign x_1110 = (v_289 | ~v_288);
	assign x_1109 = (v_289 | ~v_287);
	assign x_1114 = (v_289 | ~v_50);
	assign x_1111 = (v_289 | ~v_270);
	assign x_1108 = (((v_12 | ~v_44)) | v_290);
	assign x_1107 = (((~v_12 | ~v_45)) | v_291);
	assign x_1106 = (v_292 | ~v_38);
	assign x_1105 = (v_292 | ~v_40);
	assign x_1104 = (v_292 | ~v_42);
	assign x_1103 = (v_292 | ~v_43);
	assign x_1102 = (v_292 | ~v_52);
	assign x_1100 = (v_292 | ~v_63);
	assign x_1099 = (v_292 | ~v_274);
	assign x_1097 = (v_292 | ~v_291);
	assign x_1096 = (v_292 | ~v_290);
	assign x_1101 = (v_292 | ~v_53);
	assign x_1098 = (v_292 | ~v_273);
	assign x_1095 = (((((~v_292 | ~v_289)) | ~v_286)) | v_293);
	assign x_1094 = (v_294 | ~v_255);
	assign x_1093 = (v_294 | ~v_254);
	assign x_1092 = (v_294 | ~v_253);
	assign x_1091 = (v_294 | ~v_252);
	assign x_1090 = (v_294 | ~v_293);
	assign x_1089 = (v_294 | ~v_283);
	assign x_1087 = (v_295 | ~v_25);
	assign x_1086 = (v_295 | ~v_46);
	assign x_1084 = (v_295 | ~v_48);
	assign x_1083 = (v_295 | ~v_55);
	assign x_1081 = (v_295 | ~v_239);
	assign x_1080 = (v_295 | ~v_238);
	assign x_1078 = (v_295 | ~v_284);
	assign x_1088 = (v_295 | ~v_22);
	assign x_1085 = (v_295 | ~v_47);
	assign x_1082 = (v_295 | ~v_61);
	assign x_1079 = (v_295 | ~v_285);
	assign x_1077 = (v_296 | ~v_31);
	assign x_1075 = (v_296 | ~v_49);
	assign x_1074 = (v_296 | ~v_50);
	assign x_1072 = (v_296 | ~v_56);
	assign x_1071 = (v_296 | ~v_62);
	assign x_1069 = (v_296 | ~v_243);
	assign x_1068 = (v_296 | ~v_288);
	assign x_1067 = (v_296 | ~v_287);
	assign x_1076 = (v_296 | ~v_34);
	assign x_1073 = (v_296 | ~v_51);
	assign x_1070 = (v_296 | ~v_244);
	assign x_1066 = (v_297 | ~v_40);
	assign x_1065 = (v_297 | ~v_43);
	assign x_1064 = (v_297 | ~v_52);
	assign x_1062 = (v_297 | ~v_54);
	assign x_1061 = (v_297 | ~v_57);
	assign x_1059 = (v_297 | ~v_291);
	assign x_1058 = (v_297 | ~v_290);
	assign x_1056 = (v_297 | ~v_248);
	assign x_1063 = (v_297 | ~v_53);
	assign x_1060 = (v_297 | ~v_63);
	assign x_1057 = (v_297 | ~v_249);
	assign x_1055 = (((((~v_297 | ~v_296)) | ~v_295)) | v_298);
	assign x_1054 = (v_299 | ~v_255);
	assign x_1053 = (v_299 | ~v_254);
	assign x_1052 = (v_299 | ~v_253);
	assign x_1051 = (v_299 | ~v_252);
	assign x_1049 = (v_299 | ~v_281);
	assign x_1050 = (v_299 | ~v_298);
	assign x_1048 = (v_300 | ~v_21);
	assign x_1046 = (v_300 | ~v_23);
	assign x_1045 = (v_300 | ~v_24);
	assign x_1043 = (v_300 | ~v_46);
	assign x_1042 = (v_300 | ~v_55);
	assign x_1041 = (v_300 | ~v_239);
	assign x_1040 = (v_300 | ~v_238);
	assign x_1039 = (v_300 | ~v_258);
	assign x_1038 = (v_300 | ~v_257);
	assign x_1047 = (v_300 | ~v_22);
	assign x_1044 = (v_300 | ~v_25);
	assign x_1036 = (v_301 | ~v_31);
	assign x_1035 = (v_301 | ~v_32);
	assign x_1033 = (v_301 | ~v_34);
	assign x_1032 = (v_301 | ~v_49);
	assign x_1030 = (v_301 | ~v_244);
	assign x_1029 = (v_301 | ~v_243);
	assign x_1027 = (v_301 | ~v_260);
	assign x_1037 = (v_301 | ~v_30);
	assign x_1034 = (v_301 | ~v_33);
	assign x_1031 = (v_301 | ~v_56);
	assign x_1028 = (v_301 | ~v_261);
	assign x_1026 = (v_302 | ~v_39);
	assign x_1024 = (v_302 | ~v_41);
	assign x_1023 = (v_302 | ~v_42);
	assign x_1021 = (v_302 | ~v_52);
	assign x_1020 = (v_302 | ~v_57);
	assign x_1018 = (v_302 | ~v_248);
	assign x_1017 = (v_302 | ~v_264);
	assign x_1016 = (v_302 | ~v_263);
	assign x_1025 = (v_302 | ~v_40);
	assign x_1022 = (v_302 | ~v_43);
	assign x_1019 = (v_302 | ~v_249);
	assign x_1015 = (((((~v_302 | ~v_301)) | ~v_300)) | v_303);
	assign x_1014 = (v_304 | ~v_255);
	assign x_1013 = (v_304 | ~v_254);
	assign x_1011 = (v_304 | ~v_252);
	assign x_1010 = (v_304 | ~v_303);
	assign x_1012 = (v_304 | ~v_253);
	assign x_1009 = (v_304 | ~v_276);
	assign x_1008 = (v_305 | ~v_255);
	assign x_1007 = (v_305 | ~v_254);
	assign x_1005 = (v_305 | ~v_252);
	assign x_1004 = (v_305 | ~v_251);
	assign x_1006 = (v_305 | ~v_253);
	assign x_1003 = (((((~v_305 | ~v_304)) | ~v_299)) | v_306);
	assign x_1002 = (v_307 | ~v_20);
	assign x_1001 = (v_307 | ~v_22);
	assign x_1000 = (v_307 | ~v_23);
	assign x_998 = (v_307 | ~v_25);
	assign x_997 = (v_307 | ~v_46);
	assign x_995 = (v_307 | ~v_268);
	assign x_994 = (v_307 | ~v_222);
	assign x_992 = (v_307 | ~v_267);
	assign x_999 = (v_307 | ~v_24);
	assign x_996 = (v_307 | ~v_47);
	assign x_993 = (v_307 | ~v_221);
	assign x_991 = (v_308 | ~v_29);
	assign x_990 = (v_308 | ~v_31);
	assign x_989 = (v_308 | ~v_32);
	assign x_988 = (v_308 | ~v_33);
	assign x_987 = (v_308 | ~v_34);
	assign x_985 = (v_308 | ~v_50);
	assign x_984 = (v_308 | ~v_271);
	assign x_982 = (v_308 | ~v_227);
	assign x_981 = (v_308 | ~v_226);
	assign x_986 = (v_308 | ~v_49);
	assign x_983 = (v_308 | ~v_270);
	assign x_979 = (v_309 | ~v_40);
	assign x_978 = (v_309 | ~v_41);
	assign x_976 = (v_309 | ~v_43);
	assign x_975 = (v_309 | ~v_52);
	assign x_973 = (v_309 | ~v_274);
	assign x_972 = (v_309 | ~v_273);
	assign x_970 = (v_309 | ~v_231);
	assign x_980 = (v_309 | ~v_38);
	assign x_977 = (v_309 | ~v_42);
	assign x_974 = (v_309 | ~v_53);
	assign x_971 = (v_309 | ~v_232);
	assign x_969 = (((((~v_309 | ~v_308)) | ~v_307)) | v_310);
	assign x_967 = (v_311 | ~v_254);
	assign x_966 = (v_311 | ~v_253);
	assign x_965 = (v_311 | ~v_252);
	assign x_964 = (v_311 | ~v_310);
	assign x_963 = (v_311 | ~v_306);
	assign x_968 = (v_311 | ~v_255);
	assign x_962 = (v_312 | ~v_255);
	assign x_960 = (v_312 | ~v_253);
	assign x_959 = (v_312 | ~v_252);
	assign x_957 = (v_312 | ~v_281);
	assign x_961 = (v_312 | ~v_254);
	assign x_958 = (v_312 | ~v_293);
	assign x_956 = (v_313 | ~v_255);
	assign x_954 = (v_313 | ~v_253);
	assign x_953 = (v_313 | ~v_252);
	assign x_952 = (v_313 | ~v_251);
	assign x_951 = (v_313 | ~v_310);
	assign x_955 = (v_313 | ~v_254);
	assign x_950 = (v_314 | ~v_255);
	assign x_949 = (v_314 | ~v_254);
	assign x_947 = (v_314 | ~v_252);
	assign x_946 = (v_314 | ~v_276);
	assign x_948 = (v_314 | ~v_253);
	assign x_945 = (((((((((~v_314 | ~v_313)) | ~v_312)) | ~v_311)) | ~v_294)) | v_315);
	assign x_944 = (v_316 | ~v_255);
	assign x_943 = (v_316 | ~v_254);
	assign x_941 = (v_316 | ~v_252);
	assign x_940 = (v_316 | ~v_298);
	assign x_939 = (v_316 | ~v_310);
	assign x_942 = (v_316 | ~v_253);
	assign x_938 = (((~v_14 | v_10)) | v_317);
	assign x_937 = (((~v_10 | ~v_16)) | v_318);
	assign x_936 = (v_319 | ~v_31);
	assign x_934 = (v_319 | ~v_34);
	assign x_933 = (v_319 | ~v_49);
	assign x_931 = (v_319 | ~v_56);
	assign x_930 = (v_319 | ~v_62);
	assign x_928 = (v_319 | ~v_317);
	assign x_927 = (v_319 | ~v_288);
	assign x_935 = (v_319 | ~v_33);
	assign x_932 = (v_319 | ~v_50);
	assign x_929 = (v_319 | ~v_318);
	assign x_926 = (v_319 | ~v_287);
	assign x_925 = (((~v_15 | v_10)) | v_320);
	assign x_924 = (((~v_10 | ~v_18)) | v_321);
	assign x_922 = (v_322 | ~v_42);
	assign x_921 = (v_322 | ~v_43);
	assign x_919 = (v_322 | ~v_53);
	assign x_918 = (v_322 | ~v_57);
	assign x_916 = (v_322 | ~v_291);
	assign x_915 = (v_322 | ~v_290);
	assign x_914 = (v_322 | ~v_321);
	assign x_913 = (v_322 | ~v_320);
	assign x_923 = (v_322 | ~v_40);
	assign x_920 = (v_322 | ~v_52);
	assign x_917 = (v_322 | ~v_63);
	assign x_912 = (((~v_13 | v_10)) | v_323);
	assign x_911 = (((~v_10 | ~v_17)) | v_324);
	assign x_909 = (v_325 | ~v_24);
	assign x_908 = (v_325 | ~v_25);
	assign x_906 = (v_325 | ~v_47);
	assign x_905 = (v_325 | ~v_55);
	assign x_903 = (v_325 | ~v_324);
	assign x_902 = (v_325 | ~v_285);
	assign x_901 = (v_325 | ~v_323);
	assign x_900 = (v_325 | ~v_284);
	assign x_910 = (v_325 | ~v_22);
	assign x_907 = (v_325 | ~v_46);
	assign x_904 = (v_325 | ~v_61);
	assign x_899 = (((((~v_325 | ~v_322)) | ~v_319)) | v_326);
	assign x_898 = (v_327 | ~v_255);
	assign x_896 = (v_327 | ~v_253);
	assign x_895 = (v_327 | ~v_252);
	assign x_893 = (v_327 | ~v_276);
	assign x_897 = (v_327 | ~v_254);
	assign x_894 = (v_327 | ~v_326);
	assign x_892 = (v_328 | ~v_255);
	assign x_890 = (v_328 | ~v_253);
	assign x_889 = (v_328 | ~v_252);
	assign x_888 = (v_328 | ~v_293);
	assign x_891 = (v_328 | ~v_254);
	assign x_887 = (((((~v_328 | ~v_327)) | ~v_316)) | v_329);
	assign x_886 = (v_330 | ~v_21);
	assign x_885 = (v_330 | ~v_22);
	assign x_883 = (v_330 | ~v_24);
	assign x_882 = (v_330 | ~v_46);
	assign x_880 = (v_330 | ~v_58);
	assign x_879 = (v_330 | ~v_324);
	assign x_877 = (v_330 | ~v_257);
	assign x_876 = (v_330 | ~v_323);
	assign x_884 = (v_330 | ~v_23);
	assign x_881 = (v_330 | ~v_55);
	assign x_878 = (v_330 | ~v_258);
	assign x_874 = (v_331 | ~v_31);
	assign x_873 = (v_331 | ~v_32);
	assign x_871 = (v_331 | ~v_49);
	assign x_870 = (v_331 | ~v_56);
	assign x_868 = (v_331 | ~v_318);
	assign x_867 = (v_331 | ~v_261);
	assign x_865 = (v_331 | ~v_317);
	assign x_875 = (v_331 | ~v_30);
	assign x_872 = (v_331 | ~v_33);
	assign x_869 = (v_331 | ~v_59);
	assign x_866 = (v_331 | ~v_260);
	assign x_864 = (v_332 | ~v_39);
	assign x_863 = (v_332 | ~v_40);
	assign x_862 = (v_332 | ~v_41);
	assign x_861 = (v_332 | ~v_42);
	assign x_860 = (v_332 | ~v_52);
	assign x_858 = (v_332 | ~v_60);
	assign x_857 = (v_332 | ~v_264);
	assign x_855 = (v_332 | ~v_321);
	assign x_854 = (v_332 | ~v_320);
	assign x_859 = (v_332 | ~v_57);
	assign x_856 = (v_332 | ~v_263);
	assign x_853 = (((((~v_332 | ~v_331)) | ~v_330)) | v_333);
	assign x_852 = (v_334 | ~v_255);
	assign x_851 = (v_334 | ~v_254);
	assign x_849 = (v_334 | ~v_252);
	assign x_848 = (v_334 | ~v_333);
	assign x_850 = (v_334 | ~v_253);
	assign x_847 = (v_334 | ~v_329);
	assign x_846 = (v_335 | ~v_255);
	assign x_845 = (v_335 | ~v_254);
	assign x_843 = (v_335 | ~v_252);
	assign x_842 = (v_335 | ~v_293);
	assign x_844 = (v_335 | ~v_253);
	assign x_841 = (v_335 | ~v_303);
	assign x_840 = (v_336 | ~v_255);
	assign x_839 = (v_336 | ~v_254);
	assign x_838 = (v_336 | ~v_253);
	assign x_837 = (v_336 | ~v_252);
	assign x_836 = (v_336 | ~v_326);
	assign x_835 = (v_336 | ~v_251);
	assign x_833 = (v_337 | ~v_254);
	assign x_832 = (v_337 | ~v_253);
	assign x_830 = (v_337 | ~v_298);
	assign x_834 = (v_337 | ~v_255);
	assign x_831 = (v_337 | ~v_252);
	assign x_829 = (((((~v_337 | ~v_336)) | ~v_335)) | v_338);
	assign x_827 = (v_339 | ~v_23);
	assign x_826 = (v_339 | ~v_25);
	assign x_824 = (v_339 | ~v_47);
	assign x_823 = (v_339 | ~v_48);
	assign x_821 = (v_339 | ~v_324);
	assign x_820 = (v_339 | ~v_222);
	assign x_818 = (v_339 | ~v_323);
	assign x_828 = (v_339 | ~v_22);
	assign x_825 = (v_339 | ~v_46);
	assign x_822 = (v_339 | ~v_55);
	assign x_819 = (v_339 | ~v_221);
	assign x_817 = (v_340 | ~v_31);
	assign x_815 = (v_340 | ~v_34);
	assign x_814 = (v_340 | ~v_49);
	assign x_813 = (v_340 | ~v_50);
	assign x_812 = (v_340 | ~v_51);
	assign x_811 = (v_340 | ~v_56);
	assign x_810 = (v_340 | ~v_318);
	assign x_808 = (v_340 | ~v_226);
	assign x_807 = (v_340 | ~v_317);
	assign x_816 = (v_340 | ~v_32);
	assign x_809 = (v_340 | ~v_227);
	assign x_805 = (v_341 | ~v_41);
	assign x_804 = (v_341 | ~v_43);
	assign x_802 = (v_341 | ~v_53);
	assign x_801 = (v_341 | ~v_54);
	assign x_800 = (v_341 | ~v_57);
	assign x_799 = (v_341 | ~v_232);
	assign x_798 = (v_341 | ~v_231);
	assign x_797 = (v_341 | ~v_321);
	assign x_806 = (v_341 | ~v_40);
	assign x_803 = (v_341 | ~v_52);
	assign x_796 = (v_341 | ~v_320);
	assign x_795 = (((((~v_341 | ~v_340)) | ~v_339)) | v_342);
	assign x_794 = (v_343 | ~v_255);
	assign x_792 = (v_343 | ~v_253);
	assign x_791 = (v_343 | ~v_252);
	assign x_789 = (v_343 | ~v_338);
	assign x_793 = (v_343 | ~v_254);
	assign x_790 = (v_343 | ~v_342);
	assign x_788 = (v_344 | ~v_255);
	assign x_787 = (v_344 | ~v_254);
	assign x_786 = (v_344 | ~v_253);
	assign x_785 = (v_344 | ~v_252);
	assign x_784 = (v_344 | ~v_342);
	assign x_783 = (v_344 | ~v_298);
	assign x_782 = (v_345 | ~v_255);
	assign x_781 = (v_345 | ~v_254);
	assign x_779 = (v_345 | ~v_252);
	assign x_778 = (v_345 | ~v_333);
	assign x_780 = (v_345 | ~v_253);
	assign x_777 = (v_345 | ~v_293);
	assign x_776 = (v_346 | ~v_255);
	assign x_775 = (v_346 | ~v_254);
	assign x_773 = (v_346 | ~v_252);
	assign x_772 = (v_346 | ~v_326);
	assign x_774 = (v_346 | ~v_253);
	assign x_771 = (((((((((~v_346 | ~v_345)) | ~v_344)) | ~v_343)) | ~v_334)) | v_347);
	assign x_770 = (v_348 | ~v_347);
	assign x_769 = (v_348 | ~v_315);
	assign x_767 = (v_349 | ~v_254);
	assign x_766 = (v_349 | ~v_253);
	assign x_764 = (v_349 | ~v_342);
	assign x_763 = (v_349 | ~v_281);
	assign x_768 = (v_349 | ~v_255);
	assign x_765 = (v_349 | ~v_252);
	assign x_762 = (v_350 | ~v_255);
	assign x_761 = (v_350 | ~v_254);
	assign x_760 = (v_350 | ~v_253);
	assign x_759 = (v_350 | ~v_252);
	assign x_757 = (v_350 | ~v_266);
	assign x_758 = (v_350 | ~v_310);
	assign x_756 = (v_351 | ~v_255);
	assign x_754 = (v_351 | ~v_253);
	assign x_753 = (v_351 | ~v_252);
	assign x_755 = (v_351 | ~v_254);
	assign x_752 = (v_351 | ~v_235);
	assign x_751 = (((((~v_351 | ~v_350)) | ~v_349)) | v_352);
	assign x_750 = (v_353 | ~v_255);
	assign x_749 = (v_353 | ~v_254);
	assign x_748 = (v_353 | ~v_253);
	assign x_747 = (v_353 | ~v_252);
	assign x_746 = (v_353 | ~v_293);
	assign x_745 = (v_353 | ~v_352);
	assign x_744 = (v_354 | ~v_255);
	assign x_743 = (v_354 | ~v_254);
	assign x_741 = (v_354 | ~v_252);
	assign x_740 = (v_354 | ~v_326);
	assign x_742 = (v_354 | ~v_253);
	assign x_739 = (v_354 | ~v_235);
	assign x_738 = (v_355 | ~v_255);
	assign x_737 = (v_355 | ~v_254);
	assign x_736 = (v_355 | ~v_253);
	assign x_735 = (v_355 | ~v_252);
	assign x_734 = (v_355 | ~v_333);
	assign x_733 = (v_355 | ~v_310);
	assign x_731 = (v_356 | ~v_254);
	assign x_730 = (v_356 | ~v_253);
	assign x_728 = (v_356 | ~v_342);
	assign x_732 = (v_356 | ~v_255);
	assign x_729 = (v_356 | ~v_252);
	assign x_727 = (((((~v_356 | ~v_355)) | ~v_354)) | v_357);
	assign x_725 = (v_358 | ~v_254);
	assign x_724 = (v_358 | ~v_253);
	assign x_722 = (v_358 | ~v_276);
	assign x_721 = (v_358 | ~v_357);
	assign x_726 = (v_358 | ~v_255);
	assign x_723 = (v_358 | ~v_252);
	assign x_719 = (v_359 | ~v_254);
	assign x_718 = (v_359 | ~v_253);
	assign x_716 = (v_359 | ~v_342);
	assign x_715 = (v_359 | ~v_276);
	assign x_720 = (v_359 | ~v_255);
	assign x_717 = (v_359 | ~v_252);
	assign x_713 = (v_360 | ~v_254);
	assign x_712 = (v_360 | ~v_253);
	assign x_711 = (v_360 | ~v_252);
	assign x_710 = (v_360 | ~v_293);
	assign x_709 = (v_360 | ~v_235);
	assign x_714 = (v_360 | ~v_255);
	assign x_708 = (v_361 | ~v_255);
	assign x_706 = (v_361 | ~v_253);
	assign x_705 = (v_361 | ~v_252);
	assign x_707 = (v_361 | ~v_254);
	assign x_704 = (v_361 | ~v_310);
	assign x_703 = (((((((((~v_361 | ~v_360)) | ~v_359)) | ~v_358)) | ~v_353)) | v_362);
	assign x_702 = (v_363 | ~v_255);
	assign x_700 = (v_363 | ~v_253);
	assign x_699 = (v_363 | ~v_252);
	assign x_698 = (v_363 | ~v_303);
	assign x_697 = (v_363 | ~v_329);
	assign x_701 = (v_363 | ~v_254);
	assign x_696 = (((((~v_346 | ~v_345)) | ~v_344)) | v_364);
	assign x_695 = (v_365 | ~v_255);
	assign x_693 = (v_365 | ~v_253);
	assign x_692 = (v_365 | ~v_252);
	assign x_690 = (v_365 | ~v_251);
	assign x_694 = (v_365 | ~v_254);
	assign x_691 = (v_365 | ~v_364);
	assign x_689 = (((((((((~v_337 | ~v_336)) | ~v_335)) | ~v_365)) | ~v_363)) | v_366);
	assign x_687 = (v_367 | ~v_362);
	assign x_688 = (v_367 | ~v_366);
	assign x_686 = (v_368 | ~v_255);
	assign x_685 = (v_368 | ~v_254);
	assign x_684 = (v_368 | ~v_253);
	assign x_683 = (v_368 | ~v_252);
	assign x_682 = (v_368 | ~v_338);
	assign x_681 = (v_368 | ~v_310);
	assign x_680 = (v_369 | ~v_255);
	assign x_679 = (v_369 | ~v_254);
	assign x_677 = (v_369 | ~v_252);
	assign x_676 = (v_369 | ~v_364);
	assign x_678 = (v_369 | ~v_253);
	assign x_675 = (v_369 | ~v_276);
	assign x_674 = (((((((((((((((~v_328 | ~v_327)) | ~v_316)) | ~v_369)) | ~v_368)) | ~v_367)) | ~v_348)) | ~v_219)) | v_370);
	assign x_673 = (v_371 | ~v_370);
	assign x_672 = (v_371 | ~v_218);
	assign x_671 = (v_372 | ~v_4);
	assign x_670 = (v_372 | ~v_5);
	assign x_668 = (v_372 | ~v_8);
	assign x_669 = (v_372 | ~v_6);
	assign x_667 = (v_373 | ~v_1);
	assign x_665 = (v_373 | ~v_3);
	assign x_664 = (v_373 | ~v_7);
	assign x_666 = (v_373 | ~v_2);
	assign x_663 = (((((((((((((((v_5 | v_6)) | v_8)) | v_3)) | v_2)) | v_1)) | ~v_373)) | ~v_372)) | ~v_371);
	assign x_662 = (v_375 | ~v_208);
	assign x_661 = (v_375 | ~v_207);
	assign x_660 = (v_375 | ~v_206);
	assign x_659 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_180)) | ~v_375)) | v_376);
	assign x_658 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_173)) | ~v_199)) | v_377);
	assign x_657 = (v_378 | ~v_203);
	assign x_655 = (v_378 | ~v_201);
	assign x_654 = (v_378 | ~v_377);
	assign x_656 = (v_378 | ~v_202);
	assign x_653 = (v_378 | ~v_376);
	assign x_652 = (((~v_378 | ~v_162)) | v_379);
	assign x_651 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_113)) | ~v_375)) | v_380);
	assign x_650 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_204)) | ~v_128)) | v_381);
	assign x_649 = (v_382 | ~v_198);
	assign x_648 = (v_382 | ~v_197);
	assign x_647 = (v_382 | ~v_196);
	assign x_646 = (v_382 | ~v_381);
	assign x_645 = (v_382 | ~v_380);
	assign x_644 = (v_383 | ~v_175);
	assign x_642 = (v_383 | ~v_163);
	assign x_641 = (v_383 | ~v_216);
	assign x_643 = (v_383 | ~v_174);
	assign x_640 = (v_383 | ~v_215);
	assign x_639 = (((~v_383 | ~v_382)) | v_384);
	assign x_638 = (v_385 | ~v_208);
	assign x_636 = (v_385 | ~v_206);
	assign x_635 = (v_385 | ~v_205);
	assign x_634 = (v_385 | ~v_200);
	assign x_633 = (v_385 | ~v_384);
	assign x_632 = (v_385 | ~v_379);
	assign x_637 = (v_385 | ~v_207);
	assign x_631 = (((((((((~v_9 | ~v_10)) | ~v_11)) | ~v_12)) | ~v_385)) | v_386);
	assign x_630 = (((((~v_361 | ~v_360)) | ~v_359)) | v_387);
	assign x_629 = (v_388 | ~v_255);
	assign x_628 = (v_388 | ~v_254);
	assign x_626 = (v_388 | ~v_252);
	assign x_625 = (v_388 | ~v_333);
	assign x_627 = (v_388 | ~v_253);
	assign x_624 = (v_388 | ~v_387);
	assign x_623 = (v_389 | ~v_255);
	assign x_622 = (v_389 | ~v_254);
	assign x_620 = (v_389 | ~v_252);
	assign x_619 = (v_389 | ~v_326);
	assign x_621 = (v_389 | ~v_253);
	assign x_618 = (v_389 | ~v_352);
	assign x_617 = (((((((((~v_356 | ~v_355)) | ~v_354)) | ~v_389)) | ~v_388)) | v_390);
	assign x_616 = (v_391 | ~v_390);
	assign x_615 = (v_391 | ~v_315);
	assign x_614 = (v_392 | ~v_255);
	assign x_613 = (v_392 | ~v_254);
	assign x_611 = (v_392 | ~v_252);
	assign x_610 = (v_392 | ~v_266);
	assign x_609 = (v_392 | ~v_387);
	assign x_612 = (v_392 | ~v_253);
	assign x_608 = (v_393 | ~v_255);
	assign x_607 = (v_393 | ~v_254);
	assign x_606 = (v_393 | ~v_253);
	assign x_604 = (v_393 | ~v_357);
	assign x_603 = (v_393 | ~v_281);
	assign x_605 = (v_393 | ~v_252);
	assign x_602 = (((((((((~v_351 | ~v_350)) | ~v_349)) | ~v_393)) | ~v_392)) | v_394);
	assign x_601 = (((((((((~v_328 | ~v_327)) | ~v_316)) | ~v_369)) | ~v_368)) | v_395);
	assign x_600 = (v_396 | ~v_395);
	assign x_599 = (v_396 | ~v_394);
	assign x_598 = (((((((((((((((~v_361 | ~v_360)) | ~v_359)) | ~v_358)) | ~v_353)) | ~v_396)) | ~v_391)) | ~v_219)) | v_397);
	assign x_597 = (v_398 | ~v_397);
	assign x_596 = (v_398 | ~v_386);
	assign x_595 = (((((((((((((((v_4 | v_6)) | v_8)) | v_3)) | v_2)) | v_1)) | ~v_373)) | ~v_372)) | ~v_398);
	assign x_594 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_145)) | ~v_113)) | v_400);
	assign x_593 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_180)) | ~v_98)) | v_401);
	assign x_592 = (((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_150)) | v_402);
	assign x_591 = (v_403 | ~v_402);
	assign x_590 = (v_403 | ~v_401);
	assign x_589 = (v_403 | ~v_400);
	assign x_588 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_82)) | ~v_403)) | v_404);
	assign x_587 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_189)) | ~v_150)) | v_405);
	assign x_586 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_173)) | ~v_113)) | v_406);
	assign x_585 = (((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_180)) | v_407);
	assign x_584 = (v_408 | ~v_407);
	assign x_583 = (v_408 | ~v_406);
	assign x_582 = (v_408 | ~v_405);
	assign x_581 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_128)) | ~v_408)) | v_409);
	assign x_580 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_150)) | ~v_82)) | v_410);
	assign x_579 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_180)) | ~v_128)) | v_411);
	assign x_578 = (((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_113)) | v_412);
	assign x_577 = (v_413 | ~v_412);
	assign x_575 = (v_413 | ~v_410);
	assign x_574 = (v_413 | ~v_409);
	assign x_576 = (v_413 | ~v_411);
	assign x_573 = (v_413 | ~v_404);
	assign x_572 = (((~v_413 | ~v_162)) | v_414);
	assign x_571 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_145)) | ~v_130)) | v_415);
	assign x_569 = (v_416 | ~v_160);
	assign x_568 = (v_416 | ~v_159);
	assign x_570 = (v_416 | ~v_161);
	assign x_567 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_150)) | ~v_416)) | v_417);
	assign x_566 = (v_418 | ~v_152);
	assign x_565 = (v_418 | ~v_151);
	assign x_563 = (v_418 | ~v_417);
	assign x_562 = (v_418 | ~v_415);
	assign x_564 = (v_418 | ~v_146);
	assign x_561 = (((~v_418 | ~v_382)) | v_419);
	assign x_560 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_82)) | ~v_153)) | v_420);
	assign x_559 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_113)) | ~v_416)) | v_421);
	assign x_558 = (v_422 | ~v_129);
	assign x_557 = (v_422 | ~v_421);
	assign x_556 = (v_422 | ~v_420);
	assign x_555 = (v_422 | ~v_124);
	assign x_553 = (v_422 | ~v_419);
	assign x_552 = (v_422 | ~v_414);
	assign x_554 = (v_422 | ~v_103);
	assign x_551 = (((((((((~v_9 | ~v_10)) | ~v_11)) | ~v_12)) | ~v_422)) | v_423);
	assign x_550 = (v_424 | ~v_255);
	assign x_549 = (v_424 | ~v_254);
	assign x_547 = (v_424 | ~v_252);
	assign x_546 = (v_424 | ~v_298);
	assign x_545 = (v_424 | ~v_266);
	assign x_548 = (v_424 | ~v_253);
	assign x_544 = (v_425 | ~v_255);
	assign x_543 = (v_425 | ~v_254);
	assign x_542 = (v_425 | ~v_253);
	assign x_540 = (v_425 | ~v_333);
	assign x_539 = (v_425 | ~v_251);
	assign x_541 = (v_425 | ~v_252);
	assign x_537 = (v_426 | ~v_254);
	assign x_536 = (v_426 | ~v_253);
	assign x_534 = (v_426 | ~v_303);
	assign x_538 = (v_426 | ~v_255);
	assign x_535 = (v_426 | ~v_252);
	assign x_533 = (((((~v_426 | ~v_425)) | ~v_424)) | v_427);
	assign x_532 = (v_428 | ~v_255);
	assign x_531 = (v_428 | ~v_254);
	assign x_530 = (v_428 | ~v_253);
	assign x_529 = (v_428 | ~v_252);
	assign x_527 = (v_428 | ~v_427);
	assign x_528 = (v_428 | ~v_235);
	assign x_526 = (v_429 | ~v_255);
	assign x_524 = (v_429 | ~v_253);
	assign x_523 = (v_429 | ~v_252);
	assign x_521 = (v_429 | ~v_303);
	assign x_525 = (v_429 | ~v_254);
	assign x_522 = (v_429 | ~v_342);
	assign x_520 = (v_430 | ~v_255);
	assign x_518 = (v_430 | ~v_253);
	assign x_517 = (v_430 | ~v_252);
	assign x_515 = (v_430 | ~v_266);
	assign x_519 = (v_430 | ~v_254);
	assign x_516 = (v_430 | ~v_326);
	assign x_514 = (v_431 | ~v_255);
	assign x_512 = (v_431 | ~v_253);
	assign x_511 = (v_431 | ~v_252);
	assign x_513 = (v_431 | ~v_254);
	assign x_510 = (v_431 | ~v_333);
	assign x_509 = (((((~v_431 | ~v_430)) | ~v_429)) | v_432);
	assign x_508 = (v_433 | ~v_255);
	assign x_507 = (v_433 | ~v_254);
	assign x_506 = (v_433 | ~v_253);
	assign x_505 = (v_433 | ~v_252);
	assign x_504 = (v_433 | ~v_281);
	assign x_503 = (v_433 | ~v_432);
	assign x_502 = (v_434 | ~v_255);
	assign x_501 = (v_434 | ~v_254);
	assign x_499 = (v_434 | ~v_252);
	assign x_498 = (v_434 | ~v_303);
	assign x_500 = (v_434 | ~v_253);
	assign x_497 = (v_434 | ~v_235);
	assign x_496 = (v_435 | ~v_255);
	assign x_495 = (v_435 | ~v_254);
	assign x_494 = (v_435 | ~v_253);
	assign x_493 = (v_435 | ~v_252);
	assign x_492 = (v_435 | ~v_333);
	assign x_491 = (v_435 | ~v_281);
	assign x_489 = (v_436 | ~v_254);
	assign x_488 = (v_436 | ~v_253);
	assign x_486 = (v_436 | ~v_266);
	assign x_490 = (v_436 | ~v_255);
	assign x_487 = (v_436 | ~v_252);
	assign x_485 = (((((((((~v_436 | ~v_435)) | ~v_434)) | ~v_433)) | ~v_428)) | v_437);
	assign x_483 = (v_438 | ~v_315);
	assign x_484 = (v_438 | ~v_437);
	assign x_482 = (v_439 | ~v_255);
	assign x_481 = (v_439 | ~v_254);
	assign x_480 = (v_439 | ~v_253);
	assign x_479 = (v_439 | ~v_252);
	assign x_478 = (v_439 | ~v_298);
	assign x_477 = (v_439 | ~v_283);
	assign x_476 = (((((~v_314 | ~v_313)) | ~v_312)) | v_440);
	assign x_475 = (v_441 | ~v_255);
	assign x_473 = (v_441 | ~v_253);
	assign x_472 = (v_441 | ~v_252);
	assign x_470 = (v_441 | ~v_440);
	assign x_474 = (v_441 | ~v_254);
	assign x_471 = (v_441 | ~v_303);
	assign x_469 = (((((((((~v_305 | ~v_304)) | ~v_299)) | ~v_441)) | ~v_439)) | v_442);
	assign x_467 = (v_443 | ~v_394);
	assign x_468 = (v_443 | ~v_442);
	assign x_466 = (v_444 | ~v_255);
	assign x_464 = (v_444 | ~v_253);
	assign x_463 = (v_444 | ~v_252);
	assign x_461 = (v_444 | ~v_306);
	assign x_465 = (v_444 | ~v_254);
	assign x_462 = (v_444 | ~v_235);
	assign x_460 = (v_445 | ~v_255);
	assign x_458 = (v_445 | ~v_253);
	assign x_457 = (v_445 | ~v_252);
	assign x_456 = (v_445 | ~v_266);
	assign x_455 = (v_445 | ~v_440);
	assign x_459 = (v_445 | ~v_254);
	assign x_454 = (((((((((((((((~v_282 | ~v_445)) | ~v_444)) | ~v_277)) | ~v_256)) | ~v_443)) | ~v_438)) | ~v_219)) | v_446);
	assign x_453 = (v_447 | ~v_446);
	assign x_451 = (((((((((((((((v_7 | v_5)) | v_4)) | v_8)) | v_3)) | v_2)) | ~v_373)) | ~v_372)) | ~v_447);
	assign x_452 = (v_447 | ~v_423);
	assign x_450 = (v_449 | ~v_129);
	assign x_448 = (v_449 | ~v_420);
	assign x_447 = (v_449 | ~v_124);
	assign x_449 = (v_449 | ~v_421);
	assign x_446 = (v_449 | ~v_103);
	assign x_445 = (v_450 | ~v_412);
	assign x_444 = (v_450 | ~v_411);
	assign x_443 = (v_450 | ~v_410);
	assign x_442 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_173)) | ~v_450)) | v_451);
	assign x_441 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_189)) | ~v_403)) | v_452);
	assign x_440 = (v_453 | ~v_407);
	assign x_438 = (v_453 | ~v_405);
	assign x_437 = (v_453 | ~v_452);
	assign x_439 = (v_453 | ~v_406);
	assign x_436 = (v_453 | ~v_451);
	assign x_435 = (((~v_453 | ~v_449)) | v_454);
	assign x_434 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_145)) | ~v_450)) | v_455);
	assign x_433 = (((((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_98)) | ~v_408)) | v_456);
	assign x_432 = (v_457 | ~v_402);
	assign x_431 = (v_457 | ~v_401);
	assign x_430 = (v_457 | ~v_400);
	assign x_429 = (v_457 | ~v_456);
	assign x_428 = (v_457 | ~v_455);
	assign x_427 = (((~v_457 | ~v_382)) | v_458);
	assign x_425 = (v_459 | ~v_411);
	assign x_424 = (v_459 | ~v_410);
	assign x_422 = (v_459 | ~v_404);
	assign x_421 = (v_459 | ~v_458);
	assign x_426 = (v_459 | ~v_412);
	assign x_423 = (v_459 | ~v_409);
	assign x_420 = (v_459 | ~v_454);
	assign x_419 = (((((((((~v_9 | ~v_10)) | ~v_11)) | ~v_12)) | ~v_459)) | v_460);
	assign x_418 = (((((((((~v_282 | ~v_445)) | ~v_444)) | ~v_277)) | ~v_256)) | v_461);
	assign x_417 = (((((~v_436 | ~v_435)) | ~v_434)) | v_462);
	assign x_416 = (v_463 | ~v_255);
	assign x_415 = (v_463 | ~v_254);
	assign x_413 = (v_463 | ~v_252);
	assign x_412 = (v_463 | ~v_326);
	assign x_414 = (v_463 | ~v_253);
	assign x_411 = (v_463 | ~v_462);
	assign x_410 = (v_464 | ~v_255);
	assign x_409 = (v_464 | ~v_254);
	assign x_407 = (v_464 | ~v_252);
	assign x_406 = (v_464 | ~v_342);
	assign x_405 = (v_464 | ~v_427);
	assign x_408 = (v_464 | ~v_253);
	assign x_404 = (((((((((~v_431 | ~v_430)) | ~v_429)) | ~v_464)) | ~v_463)) | v_465);
	assign x_403 = (v_466 | ~v_465);
	assign x_402 = (v_466 | ~v_461);
	assign x_400 = (v_467 | ~v_254);
	assign x_399 = (v_467 | ~v_253);
	assign x_397 = (v_467 | ~v_298);
	assign x_396 = (v_467 | ~v_462);
	assign x_401 = (v_467 | ~v_255);
	assign x_398 = (v_467 | ~v_252);
	assign x_394 = (v_468 | ~v_254);
	assign x_393 = (v_468 | ~v_253);
	assign x_392 = (v_468 | ~v_252);
	assign x_391 = (v_468 | ~v_251);
	assign x_390 = (v_468 | ~v_432);
	assign x_395 = (v_468 | ~v_255);
	assign x_389 = (((((((((~v_426 | ~v_425)) | ~v_424)) | ~v_468)) | ~v_467)) | v_469);
	assign x_387 = (v_470 | ~v_394);
	assign x_388 = (v_470 | ~v_469);
	assign x_386 = (((((((((((((((~v_436 | ~v_435)) | ~v_434)) | ~v_433)) | ~v_428)) | ~v_470)) | ~v_466)) | ~v_219)) | v_471);
	assign x_384 = (v_472 | ~v_460);
	assign x_383 = (((((((((((((((v_7 | v_5)) | v_4)) | v_6)) | v_3)) | v_2)) | ~v_373)) | ~v_372)) | ~v_472);
	assign x_385 = (v_472 | ~v_471);
	assign x_382 = (((~v_413 | ~v_209)) | v_474);
	assign x_381 = (((~v_378 | ~v_449)) | v_475);
	assign x_380 = (v_476 | ~v_198);
	assign x_379 = (v_476 | ~v_197);
	assign x_378 = (v_476 | ~v_196);
	assign x_377 = (v_476 | ~v_381);
	assign x_376 = (v_476 | ~v_380);
	assign x_374 = (v_476 | ~v_474);
	assign x_375 = (v_476 | ~v_475);
	assign x_373 = (((((((((~v_9 | ~v_10)) | ~v_11)) | ~v_12)) | ~v_476)) | v_477);
	assign x_371 = (v_478 | ~v_362);
	assign x_372 = (v_478 | ~v_437);
	assign x_370 = (v_479 | ~v_390);
	assign x_369 = (v_479 | ~v_461);
	assign x_368 = (((((((((((((((~v_351 | ~v_350)) | ~v_349)) | ~v_393)) | ~v_392)) | ~v_479)) | ~v_478)) | ~v_219)) | v_480);
	assign x_367 = (v_481 | ~v_480);
	assign x_365 = (((((((((((((((v_7 | v_4)) | v_6)) | v_8)) | v_3)) | v_2)) | ~v_373)) | ~v_372)) | ~v_481);
	assign x_366 = (v_481 | ~v_477);
	assign x_364 = (((~v_418 | ~v_209)) | v_483);
	assign x_363 = (((~v_383 | ~v_449)) | v_484);
	assign x_362 = (v_485 | ~v_161);
	assign x_361 = (v_485 | ~v_160);
	assign x_359 = (v_485 | ~v_158);
	assign x_358 = (v_485 | ~v_141);
	assign x_356 = (v_485 | ~v_483);
	assign x_360 = (v_485 | ~v_159);
	assign x_357 = (v_485 | ~v_484);
	assign x_355 = (((((((((~v_9 | ~v_10)) | ~v_11)) | ~v_12)) | ~v_485)) | v_486);
	assign x_354 = (v_487 | ~v_442);
	assign x_353 = (v_487 | ~v_362);
	assign x_352 = (v_488 | ~v_395);
	assign x_351 = (v_488 | ~v_461);
	assign x_350 = (((((((((((((((~v_314 | ~v_313)) | ~v_312)) | ~v_311)) | ~v_294)) | ~v_488)) | ~v_487)) | ~v_219)) | v_489);
	assign x_349 = (v_490 | ~v_489);
	assign x_348 = (v_490 | ~v_486);
	assign x_347 = (((((((((((((((v_5 | v_4)) | v_8)) | v_3)) | v_2)) | v_1)) | ~v_373)) | ~v_372)) | ~v_490);
	assign x_346 = (((((((((((((((((((((v_25 | v_24)) | v_23)) | v_22)) | v_21)) | v_20)) | v_19)) | ~v_115)) | ~v_105)) | ~v_104)) | ~v_114)) | v_492);
	assign x_345 = (((((((((((((((((((((v_28 | v_32)) | v_31)) | v_30)) | v_29)) | v_33)) | v_34)) | ~v_118)) | ~v_117)) | ~v_108)) | ~v_107)) | v_493);
	assign x_344 = (((((((((((((((((((((v_39 | v_38)) | v_37)) | v_43)) | v_40)) | v_42)) | v_41)) | ~v_121)) | ~v_120)) | ~v_111)) | ~v_110)) | v_494);
	assign x_343 = (v_495 | ~v_494);
	assign x_342 = (v_495 | ~v_493);
	assign x_341 = (v_495 | ~v_492);
	assign x_340 = (((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_495)) | v_496);
	assign x_339 = (((~v_457 | ~v_209)) | v_497);
	assign x_338 = (((~v_383 | ~v_413)) | v_498);
	assign x_337 = (((~v_453 | ~v_162)) | v_499);
	assign x_336 = (v_500 | ~v_499);
	assign x_335 = (v_500 | ~v_498);
	assign x_333 = (v_500 | ~v_496);
	assign x_334 = (v_500 | ~v_497);
	assign x_332 = (((((((((~v_9 | ~v_10)) | ~v_11)) | ~v_12)) | ~v_500)) | v_501);
	assign x_330 = (v_502 | ~v_20);
	assign x_329 = (v_502 | ~v_21);
	assign x_328 = (v_502 | ~v_22);
	assign x_327 = (v_502 | ~v_23);
	assign x_326 = (v_502 | ~v_24);
	assign x_325 = (v_502 | ~v_25);
	assign x_323 = (v_502 | ~v_258);
	assign x_322 = (v_502 | ~v_257);
	assign x_331 = (v_502 | ~v_19);
	assign x_324 = (v_502 | ~v_268);
	assign x_321 = (v_502 | ~v_267);
	assign x_320 = (v_503 | ~v_28);
	assign x_319 = (v_503 | ~v_29);
	assign x_317 = (v_503 | ~v_31);
	assign x_316 = (v_503 | ~v_32);
	assign x_314 = (v_503 | ~v_34);
	assign x_313 = (v_503 | ~v_271);
	assign x_311 = (v_503 | ~v_261);
	assign x_310 = (v_503 | ~v_260);
	assign x_318 = (v_503 | ~v_30);
	assign x_315 = (v_503 | ~v_33);
	assign x_312 = (v_503 | ~v_270);
	assign x_308 = (v_504 | ~v_38);
	assign x_307 = (v_504 | ~v_39);
	assign x_305 = (v_504 | ~v_41);
	assign x_304 = (v_504 | ~v_42);
	assign x_303 = (v_504 | ~v_43);
	assign x_302 = (v_504 | ~v_274);
	assign x_301 = (v_504 | ~v_273);
	assign x_300 = (v_504 | ~v_264);
	assign x_309 = (v_504 | ~v_37);
	assign x_306 = (v_504 | ~v_40);
	assign x_299 = (v_504 | ~v_263);
	assign x_298 = (((((~v_504 | ~v_503)) | ~v_502)) | v_505);
	assign x_297 = (v_506 | ~v_255);
	assign x_295 = (v_506 | ~v_253);
	assign x_294 = (v_506 | ~v_252);
	assign x_296 = (v_506 | ~v_254);
	assign x_293 = (v_506 | ~v_505);
	assign x_292 = (v_507 | ~v_469);
	assign x_291 = (v_507 | ~v_362);
	assign x_290 = (v_508 | ~v_395);
	assign x_289 = (v_508 | ~v_437);
	assign x_288 = (v_509 | ~v_465);
	assign x_287 = (v_509 | ~v_315);
	assign x_286 = (((((((((~v_509 | ~v_508)) | ~v_507)) | ~v_506)) | ~v_219)) | v_510);
	assign x_285 = (v_511 | ~v_510);
	assign x_284 = (v_511 | ~v_501);
	assign x_283 = (((((((((((((((v_5 | v_4)) | v_6)) | v_3)) | v_2)) | v_1)) | ~v_373)) | ~v_372)) | ~v_511);
	assign x_282 = (((((((((((((((((((((v_25 | v_24)) | v_23)) | v_22)) | v_19)) | v_55)) | v_47)) | ~v_86)) | ~v_85)) | ~v_69)) | ~v_68)) | v_513);
	assign x_281 = (((((((((((((((((((((v_28 | v_32)) | v_31)) | v_33)) | v_34)) | v_56)) | v_50)) | ~v_91)) | ~v_90)) | ~v_74)) | ~v_73)) | v_514);
	assign x_280 = (((((((((((((((((((((v_37 | v_53)) | v_43)) | v_40)) | v_57)) | v_42)) | v_41)) | ~v_96)) | ~v_95)) | ~v_79)) | ~v_78)) | v_515);
	assign x_279 = (v_516 | ~v_515);
	assign x_278 = (v_516 | ~v_514);
	assign x_277 = (v_516 | ~v_513);
	assign x_276 = (((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_516)) | v_517);
	assign x_275 = (((~v_213 | ~v_382)) | v_518);
	assign x_274 = (((~v_378 | ~v_418)) | v_519);
	assign x_272 = (v_520 | ~v_518);
	assign x_271 = (v_520 | ~v_497);
	assign x_273 = (v_520 | ~v_519);
	assign x_270 = (v_520 | ~v_517);
	assign x_269 = (((((((((~v_9 | ~v_10)) | ~v_11)) | ~v_12)) | ~v_520)) | v_521);
	assign x_268 = (v_522 | ~v_19);
	assign x_266 = (v_522 | ~v_23);
	assign x_265 = (v_522 | ~v_24);
	assign x_263 = (v_522 | ~v_47);
	assign x_262 = (v_522 | ~v_55);
	assign x_260 = (v_522 | ~v_238);
	assign x_259 = (v_522 | ~v_222);
	assign x_267 = (v_522 | ~v_22);
	assign x_264 = (v_522 | ~v_25);
	assign x_261 = (v_522 | ~v_239);
	assign x_258 = (v_522 | ~v_221);
	assign x_257 = (v_523 | ~v_28);
	assign x_256 = (v_523 | ~v_31);
	assign x_254 = (v_523 | ~v_33);
	assign x_253 = (v_523 | ~v_34);
	assign x_252 = (v_523 | ~v_50);
	assign x_251 = (v_523 | ~v_56);
	assign x_250 = (v_523 | ~v_244);
	assign x_249 = (v_523 | ~v_243);
	assign x_247 = (v_523 | ~v_226);
	assign x_255 = (v_523 | ~v_32);
	assign x_248 = (v_523 | ~v_227);
	assign x_246 = (v_524 | ~v_37);
	assign x_244 = (v_524 | ~v_41);
	assign x_243 = (v_524 | ~v_42);
	assign x_241 = (v_524 | ~v_53);
	assign x_240 = (v_524 | ~v_57);
	assign x_239 = (v_524 | ~v_249);
	assign x_238 = (v_524 | ~v_248);
	assign x_237 = (v_524 | ~v_232);
	assign x_236 = (v_524 | ~v_231);
	assign x_245 = (v_524 | ~v_40);
	assign x_242 = (v_524 | ~v_43);
	assign x_235 = (((((~v_524 | ~v_523)) | ~v_522)) | v_525);
	assign x_234 = (v_526 | ~v_255);
	assign x_233 = (v_526 | ~v_254);
	assign x_231 = (v_526 | ~v_252);
	assign x_230 = (v_526 | ~v_525);
	assign x_232 = (v_526 | ~v_253);
	assign x_228 = (v_527 | ~v_394);
	assign x_229 = (v_527 | ~v_366);
	assign x_227 = (v_528 | ~v_390);
	assign x_226 = (v_528 | ~v_442);
	assign x_225 = (((((((((~v_528 | ~v_527)) | ~v_507)) | ~v_526)) | ~v_219)) | v_529);
	assign x_224 = (v_530 | ~v_529);
	assign x_223 = (v_530 | ~v_521);
	assign x_222 = (((((((((((((((v_7 | v_4)) | v_6)) | v_8)) | v_3)) | v_1)) | ~v_373)) | ~v_372)) | ~v_530);
	assign x_221 = (((((((((((((((((((((v_25 | v_24)) | v_19)) | v_55)) | v_61)) | v_64)) | v_47)) | ~v_70)) | ~v_132)) | ~v_67)) | ~v_131)) | v_532);
	assign x_220 = (((((((((((((((((((((v_28 | v_33)) | v_34)) | v_56)) | v_50)) | v_65)) | v_62)) | ~v_75)) | ~v_72)) | ~v_135)) | ~v_134)) | v_533);
	assign x_219 = (((((((((((((((((((((v_37 | v_53)) | v_66)) | v_43)) | v_63)) | v_57)) | v_42)) | ~v_138)) | ~v_137)) | ~v_80)) | ~v_77)) | v_534);
	assign x_218 = (v_535 | ~v_534);
	assign x_217 = (v_535 | ~v_533);
	assign x_216 = (v_535 | ~v_532);
	assign x_215 = (((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_535)) | v_536);
	assign x_214 = (((~v_194 | ~v_449)) | v_537);
	assign x_212 = (v_538 | ~v_518);
	assign x_211 = (v_538 | ~v_498);
	assign x_213 = (v_538 | ~v_537);
	assign x_210 = (v_538 | ~v_536);
	assign x_209 = (((((((((~v_9 | ~v_10)) | ~v_11)) | ~v_12)) | ~v_538)) | v_539);
	assign x_208 = (v_540 | ~v_19);
	assign x_206 = (v_540 | ~v_25);
	assign x_205 = (v_540 | ~v_47);
	assign x_203 = (v_540 | ~v_61);
	assign x_202 = (v_540 | ~v_64);
	assign x_201 = (v_540 | ~v_223);
	assign x_200 = (v_540 | ~v_285);
	assign x_199 = (v_540 | ~v_220);
	assign x_198 = (v_540 | ~v_284);
	assign x_207 = (v_540 | ~v_24);
	assign x_204 = (v_540 | ~v_55);
	assign x_196 = (v_541 | ~v_33);
	assign x_195 = (v_541 | ~v_34);
	assign x_193 = (v_541 | ~v_56);
	assign x_192 = (v_541 | ~v_62);
	assign x_190 = (v_541 | ~v_228);
	assign x_189 = (v_541 | ~v_225);
	assign x_188 = (v_541 | ~v_288);
	assign x_187 = (v_541 | ~v_287);
	assign x_197 = (v_541 | ~v_28);
	assign x_194 = (v_541 | ~v_50);
	assign x_191 = (v_541 | ~v_65);
	assign x_186 = (v_542 | ~v_37);
	assign x_185 = (v_542 | ~v_42);
	assign x_183 = (v_542 | ~v_53);
	assign x_182 = (v_542 | ~v_57);
	assign x_180 = (v_542 | ~v_66);
	assign x_179 = (v_542 | ~v_291);
	assign x_177 = (v_542 | ~v_233);
	assign x_176 = (v_542 | ~v_230);
	assign x_184 = (v_542 | ~v_43);
	assign x_181 = (v_542 | ~v_63);
	assign x_178 = (v_542 | ~v_290);
	assign x_175 = (((((~v_542 | ~v_541)) | ~v_540)) | v_543);
	assign x_174 = (v_544 | ~v_255);
	assign x_173 = (v_544 | ~v_254);
	assign x_172 = (v_544 | ~v_253);
	assign x_170 = (v_544 | ~v_543);
	assign x_171 = (v_544 | ~v_252);
	assign x_169 = (v_545 | ~v_347);
	assign x_168 = (v_545 | ~v_461);
	assign x_167 = (((((((((~v_545 | ~v_527)) | ~v_508)) | ~v_544)) | ~v_219)) | v_546);
	assign x_166 = (v_547 | ~v_546);
	assign x_164 = (((((((((((((((v_7 | v_5)) | v_6)) | v_8)) | v_3)) | v_2)) | ~v_373)) | ~v_372)) | ~v_547);
	assign x_165 = (v_547 | ~v_539);
	assign x_163 = (((~v_457 | ~v_162)) | v_549);
	assign x_162 = (((~v_213 | ~v_449)) | v_550);
	assign x_161 = (v_551 | ~v_152);
	assign x_160 = (v_551 | ~v_151);
	assign x_158 = (v_551 | ~v_417);
	assign x_157 = (v_551 | ~v_415);
	assign x_155 = (v_551 | ~v_549);
	assign x_159 = (v_551 | ~v_146);
	assign x_156 = (v_551 | ~v_550);
	assign x_154 = (((((((((~v_9 | ~v_10)) | ~v_11)) | ~v_12)) | ~v_551)) | v_552);
	assign x_152 = (v_553 | ~v_315);
	assign x_153 = (v_553 | ~v_469);
	assign x_151 = (v_554 | ~v_366);
	assign x_150 = (v_554 | ~v_461);
	assign x_149 = (((((((((((((((~v_305 | ~v_304)) | ~v_299)) | ~v_441)) | ~v_439)) | ~v_554)) | ~v_553)) | ~v_219)) | v_555);
	assign x_148 = (v_556 | ~v_555);
	assign x_147 = (v_556 | ~v_552);
	assign x_146 = (((((((((((((((v_7 | v_5)) | v_4)) | v_8)) | v_3)) | v_1)) | ~v_373)) | ~v_372)) | ~v_556);
	assign x_145 = (((~v_453 | ~v_418)) | v_558);
	assign x_144 = (((~v_213 | ~v_413)) | v_559);
	assign x_142 = (v_560 | ~v_401);
	assign x_141 = (v_560 | ~v_400);
	assign x_139 = (v_560 | ~v_455);
	assign x_138 = (v_560 | ~v_559);
	assign x_137 = (v_560 | ~v_558);
	assign x_143 = (v_560 | ~v_402);
	assign x_140 = (v_560 | ~v_456);
	assign x_136 = (((((((((~v_9 | ~v_10)) | ~v_11)) | ~v_12)) | ~v_560)) | v_561);
	assign x_135 = (v_562 | ~v_465);
	assign x_134 = (v_562 | ~v_442);
	assign x_132 = (v_563 | ~v_437);
	assign x_133 = (v_563 | ~v_366);
	assign x_131 = (((((((((((((((~v_426 | ~v_425)) | ~v_424)) | ~v_468)) | ~v_467)) | ~v_563)) | ~v_562)) | ~v_219)) | v_564);
	assign x_129 = (v_565 | ~v_561);
	assign x_128 = (((((((((((((((v_7 | v_5)) | v_4)) | v_6)) | v_3)) | v_1)) | ~v_373)) | ~v_372)) | ~v_565);
	assign x_130 = (v_565 | ~v_564);
	assign x_127 = (((~v_383 | ~v_457)) | v_567);
	assign x_126 = (((~v_194 | ~v_418)) | v_568);
	assign x_125 = (v_569 | ~v_184);
	assign x_124 = (v_569 | ~v_183);
	assign x_123 = (v_569 | ~v_182);
	assign x_122 = (v_569 | ~v_212);
	assign x_121 = (v_569 | ~v_210);
	assign x_119 = (v_569 | ~v_567);
	assign x_120 = (v_569 | ~v_568);
	assign x_118 = (((((((((~v_9 | ~v_10)) | ~v_11)) | ~v_12)) | ~v_569)) | v_570);
	assign x_116 = (v_571 | ~v_469);
	assign x_117 = (v_571 | ~v_395);
	assign x_115 = (v_572 | ~v_347);
	assign x_114 = (v_572 | ~v_442);
	assign x_113 = (((((((((((((((~v_337 | ~v_336)) | ~v_335)) | ~v_365)) | ~v_363)) | ~v_572)) | ~v_571)) | ~v_219)) | v_573);
	assign x_112 = (v_574 | ~v_573);
	assign x_110 = (((((((((((((((v_7 | v_5)) | v_6)) | v_8)) | v_3)) | v_1)) | ~v_373)) | ~v_372)) | ~v_574);
	assign x_111 = (v_574 | ~v_570);
	assign x_109 = (((~v_453 | ~v_209)) | v_576);
	assign x_108 = (((~v_194 | ~v_382)) | v_577);
	assign x_107 = (v_578 | ~v_203);
	assign x_106 = (v_578 | ~v_202);
	assign x_104 = (v_578 | ~v_377);
	assign x_103 = (v_578 | ~v_376);
	assign x_101 = (v_578 | ~v_576);
	assign x_105 = (v_578 | ~v_201);
	assign x_102 = (v_578 | ~v_577);
	assign x_100 = (((((((((~v_9 | ~v_10)) | ~v_11)) | ~v_12)) | ~v_578)) | v_579);
	assign x_99 = (v_580 | ~v_465);
	assign x_98 = (v_580 | ~v_362);
	assign x_97 = (v_581 | ~v_347);
	assign x_96 = (v_581 | ~v_394);
	assign x_95 = (((((((((((((((~v_356 | ~v_355)) | ~v_354)) | ~v_389)) | ~v_388)) | ~v_581)) | ~v_580)) | ~v_219)) | v_582);
	assign x_94 = (v_583 | ~v_582);
	assign x_93 = (v_583 | ~v_579);
	assign x_92 = (((((((((((((((v_7 | v_4)) | v_6)) | v_8)) | v_2)) | v_1)) | ~v_373)) | ~v_372)) | ~v_583);
	assign x_91 = (((((((((((((((((((((v_25 | v_24)) | v_23)) | v_22)) | v_19)) | v_55)) | v_47)) | ~v_171)) | ~v_84)) | ~v_83)) | ~v_170)) | v_585);
	assign x_90 = (((((((((((((((((((((v_28 | v_32)) | v_31)) | v_33)) | v_34)) | v_56)) | v_50)) | ~v_165)) | ~v_89)) | ~v_88)) | ~v_164)) | v_586);
	assign x_89 = (((((((((((((((((((((v_37 | v_53)) | v_43)) | v_40)) | v_57)) | v_42)) | v_41)) | ~v_94)) | ~v_93)) | ~v_168)) | ~v_167)) | v_587);
	assign x_88 = (v_588 | ~v_587);
	assign x_87 = (v_588 | ~v_586);
	assign x_86 = (v_588 | ~v_585);
	assign x_85 = (((((((((~v_102 | ~v_101)) | ~v_100)) | ~v_99)) | ~v_588)) | v_589);
	assign x_84 = (v_590 | ~v_537);
	assign x_83 = (v_590 | ~v_519);
	assign x_81 = (v_590 | ~v_589);
	assign x_82 = (v_590 | ~v_499);
	assign x_80 = (((((((((~v_9 | ~v_10)) | ~v_11)) | ~v_12)) | ~v_590)) | v_591);
	assign x_78 = (v_592 | ~v_22);
	assign x_77 = (v_592 | ~v_23);
	assign x_75 = (v_592 | ~v_25);
	assign x_74 = (v_592 | ~v_47);
	assign x_73 = (v_592 | ~v_55);
	assign x_72 = (v_592 | ~v_324);
	assign x_71 = (v_592 | ~v_237);
	assign x_70 = (v_592 | ~v_236);
	assign x_79 = (v_592 | ~v_19);
	assign x_76 = (v_592 | ~v_24);
	assign x_69 = (v_592 | ~v_323);
	assign x_68 = (v_593 | ~v_28);
	assign x_67 = (v_593 | ~v_31);
	assign x_65 = (v_593 | ~v_33);
	assign x_64 = (v_593 | ~v_34);
	assign x_62 = (v_593 | ~v_56);
	assign x_61 = (v_593 | ~v_318);
	assign x_59 = (v_593 | ~v_241);
	assign x_58 = (v_593 | ~v_317);
	assign x_66 = (v_593 | ~v_32);
	assign x_63 = (v_593 | ~v_50);
	assign x_60 = (v_593 | ~v_242);
	assign x_56 = (v_594 | ~v_40);
	assign x_55 = (v_594 | ~v_41);
	assign x_53 = (v_594 | ~v_43);
	assign x_52 = (v_594 | ~v_53);
	assign x_50 = (v_594 | ~v_247);
	assign x_49 = (v_594 | ~v_246);
	assign x_48 = (v_594 | ~v_321);
	assign x_47 = (v_594 | ~v_320);
	assign x_57 = (v_594 | ~v_37);
	assign x_54 = (v_594 | ~v_42);
	assign x_51 = (v_594 | ~v_57);
	assign x_46 = (((((~v_594 | ~v_593)) | ~v_592)) | v_595);
	assign x_45 = (v_596 | ~v_255);
	assign x_43 = (v_596 | ~v_253);
	assign x_42 = (v_596 | ~v_252);
	assign x_44 = (v_596 | ~v_254);
	assign x_41 = (v_596 | ~v_595);
	assign x_40 = (((((((((~v_545 | ~v_528)) | ~v_509)) | ~v_596)) | ~v_219)) | v_597);
	assign x_39 = (v_598 | ~v_597);
	assign x_37 = (((((((((((((((v_7 | v_5)) | v_4)) | v_8)) | v_2)) | v_1)) | ~v_373)) | ~v_372)) | ~v_598);
	assign x_38 = (v_598 | ~v_591);
	assign x_36 = (((~v_378 | ~v_457)) | v_600);
	assign x_35 = (((~v_194 | ~v_413)) | v_601);
	assign x_34 = (v_602 | ~v_407);
	assign x_33 = (v_602 | ~v_406);
	assign x_31 = (v_602 | ~v_452);
	assign x_30 = (v_602 | ~v_451);
	assign x_28 = (v_602 | ~v_600);
	assign x_32 = (v_602 | ~v_405);
	assign x_29 = (v_602 | ~v_601);
	assign x_27 = (((((((((~v_9 | ~v_10)) | ~v_11)) | ~v_12)) | ~v_602)) | v_603);
	assign x_25 = (v_604 | ~v_469);
	assign x_26 = (v_604 | ~v_390);
	assign x_24 = (v_605 | ~v_347);
	assign x_23 = (v_605 | ~v_437);
	assign x_22 = (((((((((((((((~v_431 | ~v_430)) | ~v_429)) | ~v_464)) | ~v_463)) | ~v_605)) | ~v_604)) | ~v_219)) | v_606);
	assign x_21 = (v_607 | ~v_606);
	assign x_20 = (v_607 | ~v_603);
	assign x_19 = (((((((((((((((v_7 | v_5)) | v_4)) | v_6)) | v_2)) | v_1)) | ~v_373)) | ~v_372)) | ~v_607);
	assign x_18 = (((~v_383 | ~v_453)) | v_609);
	assign x_17 = (((~v_213 | ~v_378)) | v_610);
	assign x_15 = (v_611 | ~v_192);
	assign x_14 = (v_611 | ~v_191);
	assign x_12 = (v_611 | ~v_181);
	assign x_11 = (v_611 | ~v_610);
	assign x_16 = (v_611 | ~v_193);
	assign x_13 = (v_611 | ~v_190);
	assign x_10 = (v_611 | ~v_609);
	assign x_9 = (((((((((~v_9 | ~v_10)) | ~v_11)) | ~v_12)) | ~v_611)) | v_612);
	assign x_8 = (v_613 | ~v_395);
	assign x_7 = (v_613 | ~v_465);
	assign x_6 = (v_614 | ~v_366);
	assign x_5 = (v_614 | ~v_390);
	assign x_4 = (((((((((((((((~v_346 | ~v_345)) | ~v_344)) | ~v_343)) | ~v_334)) | ~v_614)) | ~v_613)) | ~v_219)) | v_615);
	assign x_3 = (v_616 | ~v_615);
	assign x_2 = (v_616 | ~v_612);
	assign x_1 = (((((((((((((((v_7 | v_5)) | v_6)) | v_8)) | v_2)) | v_1)) | ~v_373)) | ~v_372)) | ~v_616);
	assign x_3249 = (x_1629 & x_1630);
	assign x_3248 = (x_1627 & x_1628);
	assign x_3246 = (x_1625 & x_1626);
	assign x_3243 = (x_1622 & x_1623);
	assign x_3241 = (x_1619 & x_1620);
	assign x_3237 = (x_1616 & x_1617);
	assign x_3236 = (x_1614 & x_1615);
	assign x_3234 = (x_1612 & x_1613);
	assign x_3231 = (x_1609 & x_1610);
	assign x_3229 = (x_1606 & x_1607);
	assign x_3224 = (x_1603 & x_1604);
	assign x_3223 = (x_1601 & x_1602);
	assign x_3221 = (x_1599 & x_1600);
	assign x_3218 = (x_1596 & x_1597);
	assign x_3216 = (x_1593 & x_1594);
	assign x_3212 = (x_1590 & x_1591);
	assign x_3210 = (x_1587 & x_1588);
	assign x_3207 = (x_1584 & x_1585);
	assign x_3205 = (x_1581 & x_1582);
	assign x_3199 = (x_1578 & x_1579);
	assign x_3198 = (x_1576 & x_1577);
	assign x_3196 = (x_1574 & x_1575);
	assign x_3193 = (x_1571 & x_1572);
	assign x_3191 = (x_1568 & x_1569);
	assign x_3187 = (x_1565 & x_1566);
	assign x_3186 = (x_1563 & x_1564);
	assign x_3184 = (x_1561 & x_1562);
	assign x_3181 = (x_1558 & x_1559);
	assign x_3179 = (x_1555 & x_1556);
	assign x_3174 = (x_1552 & x_1553);
	assign x_3173 = (x_1550 & x_1551);
	assign x_3171 = (x_1548 & x_1549);
	assign x_3168 = (x_1545 & x_1546);
	assign x_3166 = (x_1542 & x_1543);
	assign x_3162 = (x_1539 & x_1540);
	assign x_3160 = (x_1536 & x_1537);
	assign x_3157 = (x_1533 & x_1534);
	assign x_3155 = (x_1530 & x_1531);
	assign x_3148 = (x_1527 & x_1528);
	assign x_3147 = (x_1525 & x_1526);
	assign x_3145 = (x_1523 & x_1524);
	assign x_3142 = (x_1520 & x_1521);
	assign x_3140 = (x_1517 & x_1518);
	assign x_3136 = (x_1514 & x_1515);
	assign x_3135 = (x_1512 & x_1513);
	assign x_3133 = (x_1510 & x_1511);
	assign x_3130 = (x_1507 & x_1508);
	assign x_3128 = (x_1504 & x_1505);
	assign x_3123 = (x_1501 & x_1502);
	assign x_3122 = (x_1499 & x_1500);
	assign x_3120 = (x_1497 & x_1498);
	assign x_3117 = (x_1494 & x_1495);
	assign x_3115 = (x_1491 & x_1492);
	assign x_3111 = (x_1488 & x_1489);
	assign x_3109 = (x_1485 & x_1486);
	assign x_3106 = (x_1482 & x_1483);
	assign x_3104 = (x_1479 & x_1480);
	assign x_3098 = (x_1476 & x_1477);
	assign x_3097 = (x_1474 & x_1475);
	assign x_3095 = (x_1472 & x_1473);
	assign x_3092 = (x_1469 & x_1470);
	assign x_3090 = (x_1466 & x_1467);
	assign x_3086 = (x_1463 & x_1464);
	assign x_3085 = (x_1461 & x_1462);
	assign x_3083 = (x_1459 & x_1460);
	assign x_3080 = (x_1456 & x_1457);
	assign x_3078 = (x_1453 & x_1454);
	assign x_3073 = (x_1450 & x_1451);
	assign x_3072 = (x_1448 & x_1449);
	assign x_3070 = (x_1446 & x_1447);
	assign x_3067 = (x_1443 & x_1444);
	assign x_3065 = (x_1440 & x_1441);
	assign x_3061 = (x_1437 & x_1438);
	assign x_3059 = (x_1434 & x_1435);
	assign x_3056 = (x_1431 & x_1432);
	assign x_3054 = (x_1428 & x_1429);
	assign x_3046 = (x_1425 & x_1426);
	assign x_3045 = (x_1423 & x_1424);
	assign x_3043 = (x_1421 & x_1422);
	assign x_3040 = (x_1418 & x_1419);
	assign x_3038 = (x_1415 & x_1416);
	assign x_3034 = (x_1412 & x_1413);
	assign x_3033 = (x_1410 & x_1411);
	assign x_3031 = (x_1408 & x_1409);
	assign x_3028 = (x_1405 & x_1406);
	assign x_3026 = (x_1402 & x_1403);
	assign x_3021 = (x_1399 & x_1400);
	assign x_3020 = (x_1397 & x_1398);
	assign x_3018 = (x_1395 & x_1396);
	assign x_3015 = (x_1392 & x_1393);
	assign x_3013 = (x_1389 & x_1390);
	assign x_3009 = (x_1386 & x_1387);
	assign x_3007 = (x_1383 & x_1384);
	assign x_3004 = (x_1380 & x_1381);
	assign x_3002 = (x_1377 & x_1378);
	assign x_2996 = (x_1374 & x_1375);
	assign x_2995 = (x_1372 & x_1373);
	assign x_2993 = (x_1370 & x_1371);
	assign x_2990 = (x_1367 & x_1368);
	assign x_2988 = (x_1364 & x_1365);
	assign x_2984 = (x_1361 & x_1362);
	assign x_2983 = (x_1359 & x_1360);
	assign x_2981 = (x_1357 & x_1358);
	assign x_2978 = (x_1354 & x_1355);
	assign x_2976 = (x_1351 & x_1352);
	assign x_2971 = (x_1348 & x_1349);
	assign x_2970 = (x_1346 & x_1347);
	assign x_2968 = (x_1344 & x_1345);
	assign x_2965 = (x_1341 & x_1342);
	assign x_2963 = (x_1338 & x_1339);
	assign x_2959 = (x_1335 & x_1336);
	assign x_2957 = (x_1332 & x_1333);
	assign x_2954 = (x_1329 & x_1330);
	assign x_2952 = (x_1326 & x_1327);
	assign x_2945 = (x_1323 & x_1324);
	assign x_2944 = (x_1321 & x_1322);
	assign x_2942 = (x_1319 & x_1320);
	assign x_2939 = (x_1316 & x_1317);
	assign x_2937 = (x_1313 & x_1314);
	assign x_2933 = (x_1310 & x_1311);
	assign x_2932 = (x_1308 & x_1309);
	assign x_2930 = (x_1306 & x_1307);
	assign x_2927 = (x_1303 & x_1304);
	assign x_2925 = (x_1300 & x_1301);
	assign x_2920 = (x_1297 & x_1298);
	assign x_2919 = (x_1295 & x_1296);
	assign x_2917 = (x_1293 & x_1294);
	assign x_2914 = (x_1290 & x_1291);
	assign x_2912 = (x_1287 & x_1288);
	assign x_2908 = (x_1284 & x_1285);
	assign x_2906 = (x_1281 & x_1282);
	assign x_2903 = (x_1278 & x_1279);
	assign x_2901 = (x_1275 & x_1276);
	assign x_2895 = (x_1272 & x_1273);
	assign x_2894 = (x_1270 & x_1271);
	assign x_2892 = (x_1268 & x_1269);
	assign x_2889 = (x_1265 & x_1266);
	assign x_2887 = (x_1262 & x_1263);
	assign x_2883 = (x_1259 & x_1260);
	assign x_2882 = (x_1257 & x_1258);
	assign x_2880 = (x_1255 & x_1256);
	assign x_2877 = (x_1252 & x_1253);
	assign x_2875 = (x_1249 & x_1250);
	assign x_2870 = (x_1246 & x_1247);
	assign x_2869 = (x_1244 & x_1245);
	assign x_2867 = (x_1242 & x_1243);
	assign x_2864 = (x_1239 & x_1240);
	assign x_2862 = (x_1236 & x_1237);
	assign x_2858 = (x_1233 & x_1234);
	assign x_2856 = (x_1230 & x_1231);
	assign x_2853 = (x_1227 & x_1228);
	assign x_2851 = (x_1224 & x_1225);
	assign x_2842 = (x_1221 & x_1222);
	assign x_2841 = (x_1219 & x_1220);
	assign x_2839 = (x_1217 & x_1218);
	assign x_2836 = (x_1214 & x_1215);
	assign x_2834 = (x_1211 & x_1212);
	assign x_2830 = (x_1208 & x_1209);
	assign x_2829 = (x_1206 & x_1207);
	assign x_2827 = (x_1204 & x_1205);
	assign x_2824 = (x_1201 & x_1202);
	assign x_2822 = (x_1198 & x_1199);
	assign x_2817 = (x_1195 & x_1196);
	assign x_2816 = (x_1193 & x_1194);
	assign x_2814 = (x_1191 & x_1192);
	assign x_2811 = (x_1188 & x_1189);
	assign x_2809 = (x_1185 & x_1186);
	assign x_2805 = (x_1182 & x_1183);
	assign x_2803 = (x_1179 & x_1180);
	assign x_2800 = (x_1176 & x_1177);
	assign x_2798 = (x_1173 & x_1174);
	assign x_2792 = (x_1170 & x_1171);
	assign x_2791 = (x_1168 & x_1169);
	assign x_2789 = (x_1166 & x_1167);
	assign x_2786 = (x_1163 & x_1164);
	assign x_2784 = (x_1160 & x_1161);
	assign x_2780 = (x_1157 & x_1158);
	assign x_2779 = (x_1155 & x_1156);
	assign x_2777 = (x_1153 & x_1154);
	assign x_2774 = (x_1150 & x_1151);
	assign x_2772 = (x_1147 & x_1148);
	assign x_2767 = (x_1144 & x_1145);
	assign x_2766 = (x_1142 & x_1143);
	assign x_2764 = (x_1140 & x_1141);
	assign x_2761 = (x_1137 & x_1138);
	assign x_2759 = (x_1134 & x_1135);
	assign x_2755 = (x_1131 & x_1132);
	assign x_2753 = (x_1128 & x_1129);
	assign x_2750 = (x_1125 & x_1126);
	assign x_2748 = (x_1122 & x_1123);
	assign x_2741 = (x_1119 & x_1120);
	assign x_2740 = (x_1117 & x_1118);
	assign x_2738 = (x_1115 & x_1116);
	assign x_2735 = (x_1112 & x_1113);
	assign x_2733 = (x_1109 & x_1110);
	assign x_2729 = (x_1106 & x_1107);
	assign x_2728 = (x_1104 & x_1105);
	assign x_2726 = (x_1102 & x_1103);
	assign x_2723 = (x_1099 & x_1100);
	assign x_2721 = (x_1096 & x_1097);
	assign x_2716 = (x_1093 & x_1094);
	assign x_2715 = (x_1091 & x_1092);
	assign x_2713 = (x_1089 & x_1090);
	assign x_2710 = (x_1086 & x_1087);
	assign x_2708 = (x_1083 & x_1084);
	assign x_2704 = (x_1080 & x_1081);
	assign x_2702 = (x_1077 & x_1078);
	assign x_2699 = (x_1074 & x_1075);
	assign x_2697 = (x_1071 & x_1072);
	assign x_2691 = (x_1068 & x_1069);
	assign x_2690 = (x_1066 & x_1067);
	assign x_2688 = (x_1064 & x_1065);
	assign x_2685 = (x_1061 & x_1062);
	assign x_2683 = (x_1058 & x_1059);
	assign x_2679 = (x_1055 & x_1056);
	assign x_2678 = (x_1053 & x_1054);
	assign x_2676 = (x_1051 & x_1052);
	assign x_2673 = (x_1048 & x_1049);
	assign x_2671 = (x_1045 & x_1046);
	assign x_2666 = (x_1042 & x_1043);
	assign x_2665 = (x_1040 & x_1041);
	assign x_2663 = (x_1038 & x_1039);
	assign x_2660 = (x_1035 & x_1036);
	assign x_2658 = (x_1032 & x_1033);
	assign x_2654 = (x_1029 & x_1030);
	assign x_2652 = (x_1026 & x_1027);
	assign x_2649 = (x_1023 & x_1024);
	assign x_2647 = (x_1020 & x_1021);
	assign x_2639 = (x_1017 & x_1018);
	assign x_2638 = (x_1015 & x_1016);
	assign x_2636 = (x_1013 & x_1014);
	assign x_2633 = (x_1010 & x_1011);
	assign x_2631 = (x_1007 & x_1008);
	assign x_2627 = (x_1004 & x_1005);
	assign x_2626 = (x_1002 & x_1003);
	assign x_2624 = (x_1000 & x_1001);
	assign x_2621 = (x_997 & x_998);
	assign x_2619 = (x_994 & x_995);
	assign x_2614 = (x_991 & x_992);
	assign x_2613 = (x_989 & x_990);
	assign x_2611 = (x_987 & x_988);
	assign x_2608 = (x_984 & x_985);
	assign x_2606 = (x_981 & x_982);
	assign x_2602 = (x_978 & x_979);
	assign x_2600 = (x_975 & x_976);
	assign x_2597 = (x_972 & x_973);
	assign x_2595 = (x_969 & x_970);
	assign x_2589 = (x_966 & x_967);
	assign x_2588 = (x_964 & x_965);
	assign x_2586 = (x_962 & x_963);
	assign x_2583 = (x_959 & x_960);
	assign x_2581 = (x_956 & x_957);
	assign x_2577 = (x_953 & x_954);
	assign x_2576 = (x_951 & x_952);
	assign x_2574 = (x_949 & x_950);
	assign x_2571 = (x_946 & x_947);
	assign x_2569 = (x_943 & x_944);
	assign x_2564 = (x_940 & x_941);
	assign x_2563 = (x_938 & x_939);
	assign x_2561 = (x_936 & x_937);
	assign x_2558 = (x_933 & x_934);
	assign x_2556 = (x_930 & x_931);
	assign x_2552 = (x_927 & x_928);
	assign x_2550 = (x_924 & x_925);
	assign x_2547 = (x_921 & x_922);
	assign x_2545 = (x_918 & x_919);
	assign x_2538 = (x_915 & x_916);
	assign x_2537 = (x_913 & x_914);
	assign x_2535 = (x_911 & x_912);
	assign x_2532 = (x_908 & x_909);
	assign x_2530 = (x_905 & x_906);
	assign x_2526 = (x_902 & x_903);
	assign x_2525 = (x_900 & x_901);
	assign x_2523 = (x_898 & x_899);
	assign x_2520 = (x_895 & x_896);
	assign x_2518 = (x_892 & x_893);
	assign x_2513 = (x_889 & x_890);
	assign x_2512 = (x_887 & x_888);
	assign x_2510 = (x_885 & x_886);
	assign x_2507 = (x_882 & x_883);
	assign x_2505 = (x_879 & x_880);
	assign x_2501 = (x_876 & x_877);
	assign x_2499 = (x_873 & x_874);
	assign x_2496 = (x_870 & x_871);
	assign x_2494 = (x_867 & x_868);
	assign x_2488 = (x_864 & x_865);
	assign x_2487 = (x_862 & x_863);
	assign x_2485 = (x_860 & x_861);
	assign x_2482 = (x_857 & x_858);
	assign x_2480 = (x_854 & x_855);
	assign x_2476 = (x_851 & x_852);
	assign x_2474 = (x_848 & x_849);
	assign x_2471 = (x_845 & x_846);
	assign x_2469 = (x_842 & x_843);
	assign x_2464 = (x_839 & x_840);
	assign x_2463 = (x_837 & x_838);
	assign x_2461 = (x_835 & x_836);
	assign x_2458 = (x_832 & x_833);
	assign x_2456 = (x_829 & x_830);
	assign x_2452 = (x_826 & x_827);
	assign x_2450 = (x_823 & x_824);
	assign x_2447 = (x_820 & x_821);
	assign x_2445 = (x_817 & x_818);
	assign x_2435 = (x_814 & x_815);
	assign x_2434 = (x_812 & x_813);
	assign x_2432 = (x_810 & x_811);
	assign x_2429 = (x_807 & x_808);
	assign x_2427 = (x_804 & x_805);
	assign x_2423 = (x_801 & x_802);
	assign x_2422 = (x_799 & x_800);
	assign x_2420 = (x_797 & x_798);
	assign x_2417 = (x_794 & x_795);
	assign x_2415 = (x_791 & x_792);
	assign x_2410 = (x_788 & x_789);
	assign x_2409 = (x_786 & x_787);
	assign x_2407 = (x_784 & x_785);
	assign x_2404 = (x_781 & x_782);
	assign x_2402 = (x_778 & x_779);
	assign x_2398 = (x_775 & x_776);
	assign x_2396 = (x_772 & x_773);
	assign x_2393 = (x_769 & x_770);
	assign x_2391 = (x_766 & x_767);
	assign x_2385 = (x_763 & x_764);
	assign x_2384 = (x_761 & x_762);
	assign x_2382 = (x_759 & x_760);
	assign x_2379 = (x_756 & x_757);
	assign x_2377 = (x_753 & x_754);
	assign x_2373 = (x_750 & x_751);
	assign x_2372 = (x_748 & x_749);
	assign x_2370 = (x_746 & x_747);
	assign x_2367 = (x_743 & x_744);
	assign x_2365 = (x_740 & x_741);
	assign x_2360 = (x_737 & x_738);
	assign x_2359 = (x_735 & x_736);
	assign x_2357 = (x_733 & x_734);
	assign x_2354 = (x_730 & x_731);
	assign x_2352 = (x_727 & x_728);
	assign x_2348 = (x_724 & x_725);
	assign x_2346 = (x_721 & x_722);
	assign x_2343 = (x_718 & x_719);
	assign x_2341 = (x_715 & x_716);
	assign x_2334 = (x_712 & x_713);
	assign x_2333 = (x_710 & x_711);
	assign x_2331 = (x_708 & x_709);
	assign x_2328 = (x_705 & x_706);
	assign x_2326 = (x_702 & x_703);
	assign x_2322 = (x_699 & x_700);
	assign x_2321 = (x_697 & x_698);
	assign x_2319 = (x_695 & x_696);
	assign x_2316 = (x_692 & x_693);
	assign x_2314 = (x_689 & x_690);
	assign x_2309 = (x_686 & x_687);
	assign x_2308 = (x_684 & x_685);
	assign x_2306 = (x_682 & x_683);
	assign x_2303 = (x_679 & x_680);
	assign x_2301 = (x_676 & x_677);
	assign x_2297 = (x_673 & x_674);
	assign x_2295 = (x_670 & x_671);
	assign x_2292 = (x_667 & x_668);
	assign x_2290 = (x_664 & x_665);
	assign x_2284 = (x_661 & x_662);
	assign x_2283 = (x_659 & x_660);
	assign x_2281 = (x_657 & x_658);
	assign x_2278 = (x_654 & x_655);
	assign x_2276 = (x_651 & x_652);
	assign x_2272 = (x_648 & x_649);
	assign x_2271 = (x_646 & x_647);
	assign x_2269 = (x_644 & x_645);
	assign x_2266 = (x_641 & x_642);
	assign x_2264 = (x_638 & x_639);
	assign x_2259 = (x_635 & x_636);
	assign x_2258 = (x_633 & x_634);
	assign x_2256 = (x_631 & x_632);
	assign x_2253 = (x_628 & x_629);
	assign x_2251 = (x_625 & x_626);
	assign x_2247 = (x_622 & x_623);
	assign x_2245 = (x_619 & x_620);
	assign x_2242 = (x_616 & x_617);
	assign x_2240 = (x_613 & x_614);
	assign x_2232 = (x_610 & x_611);
	assign x_2231 = (x_608 & x_609);
	assign x_2229 = (x_606 & x_607);
	assign x_2226 = (x_603 & x_604);
	assign x_2224 = (x_600 & x_601);
	assign x_2220 = (x_597 & x_598);
	assign x_2219 = (x_595 & x_596);
	assign x_2217 = (x_593 & x_594);
	assign x_2214 = (x_590 & x_591);
	assign x_2212 = (x_587 & x_588);
	assign x_2207 = (x_584 & x_585);
	assign x_2206 = (x_582 & x_583);
	assign x_2204 = (x_580 & x_581);
	assign x_2201 = (x_577 & x_578);
	assign x_2199 = (x_574 & x_575);
	assign x_2195 = (x_571 & x_572);
	assign x_2193 = (x_568 & x_569);
	assign x_2190 = (x_565 & x_566);
	assign x_2188 = (x_562 & x_563);
	assign x_2182 = (x_559 & x_560);
	assign x_2181 = (x_557 & x_558);
	assign x_2179 = (x_555 & x_556);
	assign x_2176 = (x_552 & x_553);
	assign x_2174 = (x_549 & x_550);
	assign x_2170 = (x_546 & x_547);
	assign x_2169 = (x_544 & x_545);
	assign x_2167 = (x_542 & x_543);
	assign x_2164 = (x_539 & x_540);
	assign x_2162 = (x_536 & x_537);
	assign x_2157 = (x_533 & x_534);
	assign x_2156 = (x_531 & x_532);
	assign x_2154 = (x_529 & x_530);
	assign x_2151 = (x_526 & x_527);
	assign x_2149 = (x_523 & x_524);
	assign x_2145 = (x_520 & x_521);
	assign x_2143 = (x_517 & x_518);
	assign x_2140 = (x_514 & x_515);
	assign x_2138 = (x_511 & x_512);
	assign x_2131 = (x_508 & x_509);
	assign x_2130 = (x_506 & x_507);
	assign x_2128 = (x_504 & x_505);
	assign x_2125 = (x_501 & x_502);
	assign x_2123 = (x_498 & x_499);
	assign x_2119 = (x_495 & x_496);
	assign x_2118 = (x_493 & x_494);
	assign x_2116 = (x_491 & x_492);
	assign x_2113 = (x_488 & x_489);
	assign x_2111 = (x_485 & x_486);
	assign x_2106 = (x_482 & x_483);
	assign x_2105 = (x_480 & x_481);
	assign x_2103 = (x_478 & x_479);
	assign x_2100 = (x_475 & x_476);
	assign x_2098 = (x_472 & x_473);
	assign x_2094 = (x_469 & x_470);
	assign x_2092 = (x_466 & x_467);
	assign x_2089 = (x_463 & x_464);
	assign x_2087 = (x_460 & x_461);
	assign x_2081 = (x_457 & x_458);
	assign x_2080 = (x_455 & x_456);
	assign x_2078 = (x_453 & x_454);
	assign x_2075 = (x_450 & x_451);
	assign x_2073 = (x_447 & x_448);
	assign x_2069 = (x_444 & x_445);
	assign x_2068 = (x_442 & x_443);
	assign x_2066 = (x_440 & x_441);
	assign x_2063 = (x_437 & x_438);
	assign x_2061 = (x_434 & x_435);
	assign x_2056 = (x_431 & x_432);
	assign x_2055 = (x_429 & x_430);
	assign x_2053 = (x_427 & x_428);
	assign x_2050 = (x_424 & x_425);
	assign x_2048 = (x_421 & x_422);
	assign x_2044 = (x_418 & x_419);
	assign x_2042 = (x_415 & x_416);
	assign x_2039 = (x_412 & x_413);
	assign x_2037 = (x_409 & x_410);
	assign x_2028 = (x_406 & x_407);
	assign x_2027 = (x_404 & x_405);
	assign x_2025 = (x_402 & x_403);
	assign x_2022 = (x_399 & x_400);
	assign x_2020 = (x_396 & x_397);
	assign x_2016 = (x_393 & x_394);
	assign x_2015 = (x_391 & x_392);
	assign x_2013 = (x_389 & x_390);
	assign x_2010 = (x_386 & x_387);
	assign x_2008 = (x_383 & x_384);
	assign x_2003 = (x_380 & x_381);
	assign x_2002 = (x_378 & x_379);
	assign x_2000 = (x_376 & x_377);
	assign x_1997 = (x_373 & x_374);
	assign x_1995 = (x_370 & x_371);
	assign x_1991 = (x_367 & x_368);
	assign x_1989 = (x_364 & x_365);
	assign x_1986 = (x_361 & x_362);
	assign x_1984 = (x_358 & x_359);
	assign x_1978 = (x_355 & x_356);
	assign x_1977 = (x_353 & x_354);
	assign x_1975 = (x_351 & x_352);
	assign x_1972 = (x_348 & x_349);
	assign x_1970 = (x_345 & x_346);
	assign x_1966 = (x_342 & x_343);
	assign x_1965 = (x_340 & x_341);
	assign x_1963 = (x_338 & x_339);
	assign x_1960 = (x_335 & x_336);
	assign x_1958 = (x_332 & x_333);
	assign x_1953 = (x_329 & x_330);
	assign x_1952 = (x_327 & x_328);
	assign x_1950 = (x_325 & x_326);
	assign x_1947 = (x_322 & x_323);
	assign x_1945 = (x_319 & x_320);
	assign x_1941 = (x_316 & x_317);
	assign x_1939 = (x_313 & x_314);
	assign x_1936 = (x_310 & x_311);
	assign x_1934 = (x_307 & x_308);
	assign x_1927 = (x_304 & x_305);
	assign x_1926 = (x_302 & x_303);
	assign x_1924 = (x_300 & x_301);
	assign x_1921 = (x_297 & x_298);
	assign x_1919 = (x_294 & x_295);
	assign x_1915 = (x_291 & x_292);
	assign x_1914 = (x_289 & x_290);
	assign x_1912 = (x_287 & x_288);
	assign x_1909 = (x_284 & x_285);
	assign x_1907 = (x_281 & x_282);
	assign x_1902 = (x_278 & x_279);
	assign x_1901 = (x_276 & x_277);
	assign x_1899 = (x_274 & x_275);
	assign x_1896 = (x_271 & x_272);
	assign x_1894 = (x_268 & x_269);
	assign x_1890 = (x_265 & x_266);
	assign x_1888 = (x_262 & x_263);
	assign x_1885 = (x_259 & x_260);
	assign x_1883 = (x_256 & x_257);
	assign x_1877 = (x_253 & x_254);
	assign x_1876 = (x_251 & x_252);
	assign x_1874 = (x_249 & x_250);
	assign x_1871 = (x_246 & x_247);
	assign x_1869 = (x_243 & x_244);
	assign x_1865 = (x_240 & x_241);
	assign x_1864 = (x_238 & x_239);
	assign x_1862 = (x_236 & x_237);
	assign x_1859 = (x_233 & x_234);
	assign x_1857 = (x_230 & x_231);
	assign x_1852 = (x_227 & x_228);
	assign x_1851 = (x_225 & x_226);
	assign x_1849 = (x_223 & x_224);
	assign x_1846 = (x_220 & x_221);
	assign x_1844 = (x_217 & x_218);
	assign x_1840 = (x_214 & x_215);
	assign x_1838 = (x_211 & x_212);
	assign x_1835 = (x_208 & x_209);
	assign x_1833 = (x_205 & x_206);
	assign x_1825 = (x_202 & x_203);
	assign x_1824 = (x_200 & x_201);
	assign x_1822 = (x_198 & x_199);
	assign x_1819 = (x_195 & x_196);
	assign x_1817 = (x_192 & x_193);
	assign x_1813 = (x_189 & x_190);
	assign x_1812 = (x_187 & x_188);
	assign x_1810 = (x_185 & x_186);
	assign x_1807 = (x_182 & x_183);
	assign x_1805 = (x_179 & x_180);
	assign x_1800 = (x_176 & x_177);
	assign x_1799 = (x_174 & x_175);
	assign x_1797 = (x_172 & x_173);
	assign x_1794 = (x_169 & x_170);
	assign x_1792 = (x_166 & x_167);
	assign x_1788 = (x_163 & x_164);
	assign x_1786 = (x_160 & x_161);
	assign x_1783 = (x_157 & x_158);
	assign x_1781 = (x_154 & x_155);
	assign x_1775 = (x_151 & x_152);
	assign x_1774 = (x_149 & x_150);
	assign x_1772 = (x_147 & x_148);
	assign x_1769 = (x_144 & x_145);
	assign x_1767 = (x_141 & x_142);
	assign x_1763 = (x_138 & x_139);
	assign x_1762 = (x_136 & x_137);
	assign x_1760 = (x_134 & x_135);
	assign x_1757 = (x_131 & x_132);
	assign x_1755 = (x_128 & x_129);
	assign x_1750 = (x_125 & x_126);
	assign x_1749 = (x_123 & x_124);
	assign x_1747 = (x_121 & x_122);
	assign x_1744 = (x_118 & x_119);
	assign x_1742 = (x_115 & x_116);
	assign x_1738 = (x_112 & x_113);
	assign x_1736 = (x_109 & x_110);
	assign x_1733 = (x_106 & x_107);
	assign x_1731 = (x_103 & x_104);
	assign x_1724 = (x_100 & x_101);
	assign x_1723 = (x_98 & x_99);
	assign x_1721 = (x_96 & x_97);
	assign x_1718 = (x_93 & x_94);
	assign x_1716 = (x_90 & x_91);
	assign x_1712 = (x_87 & x_88);
	assign x_1711 = (x_85 & x_86);
	assign x_1709 = (x_83 & x_84);
	assign x_1706 = (x_80 & x_81);
	assign x_1704 = (x_77 & x_78);
	assign x_1699 = (x_74 & x_75);
	assign x_1698 = (x_72 & x_73);
	assign x_1696 = (x_70 & x_71);
	assign x_1693 = (x_67 & x_68);
	assign x_1691 = (x_64 & x_65);
	assign x_1687 = (x_61 & x_62);
	assign x_1685 = (x_58 & x_59);
	assign x_1682 = (x_55 & x_56);
	assign x_1680 = (x_52 & x_53);
	assign x_1674 = (x_49 & x_50);
	assign x_1673 = (x_47 & x_48);
	assign x_1671 = (x_45 & x_46);
	assign x_1668 = (x_42 & x_43);
	assign x_1666 = (x_39 & x_40);
	assign x_1662 = (x_36 & x_37);
	assign x_1660 = (x_33 & x_34);
	assign x_1657 = (x_30 & x_31);
	assign x_1655 = (x_27 & x_28);
	assign x_1650 = (x_24 & x_25);
	assign x_1649 = (x_22 & x_23);
	assign x_1647 = (x_20 & x_21);
	assign x_1644 = (x_17 & x_18);
	assign x_1642 = (x_14 & x_15);
	assign x_1638 = (x_11 & x_12);
	assign x_1636 = (x_8 & x_9);
	assign x_1633 = (x_5 & x_6);
	assign x_1631 = (x_2 & x_3);
	assign x_3250 = (x_3248 & x_3249);
	assign x_3247 = (x_1624 & x_3246);
	assign x_3244 = (x_1621 & x_3243);
	assign x_3242 = (x_1618 & x_3241);
	assign x_3238 = (x_3236 & x_3237);
	assign x_3235 = (x_1611 & x_3234);
	assign x_3232 = (x_1608 & x_3231);
	assign x_3230 = (x_1605 & x_3229);
	assign x_3225 = (x_3223 & x_3224);
	assign x_3222 = (x_1598 & x_3221);
	assign x_3219 = (x_1595 & x_3218);
	assign x_3217 = (x_1592 & x_3216);
	assign x_3213 = (x_1589 & x_3212);
	assign x_3211 = (x_1586 & x_3210);
	assign x_3208 = (x_1583 & x_3207);
	assign x_3206 = (x_1580 & x_3205);
	assign x_3200 = (x_3198 & x_3199);
	assign x_3197 = (x_1573 & x_3196);
	assign x_3194 = (x_1570 & x_3193);
	assign x_3192 = (x_1567 & x_3191);
	assign x_3188 = (x_3186 & x_3187);
	assign x_3185 = (x_1560 & x_3184);
	assign x_3182 = (x_1557 & x_3181);
	assign x_3180 = (x_1554 & x_3179);
	assign x_3175 = (x_3173 & x_3174);
	assign x_3172 = (x_1547 & x_3171);
	assign x_3169 = (x_1544 & x_3168);
	assign x_3167 = (x_1541 & x_3166);
	assign x_3163 = (x_1538 & x_3162);
	assign x_3161 = (x_1535 & x_3160);
	assign x_3158 = (x_1532 & x_3157);
	assign x_3156 = (x_1529 & x_3155);
	assign x_3149 = (x_3147 & x_3148);
	assign x_3146 = (x_1522 & x_3145);
	assign x_3143 = (x_1519 & x_3142);
	assign x_3141 = (x_1516 & x_3140);
	assign x_3137 = (x_3135 & x_3136);
	assign x_3134 = (x_1509 & x_3133);
	assign x_3131 = (x_1506 & x_3130);
	assign x_3129 = (x_1503 & x_3128);
	assign x_3124 = (x_3122 & x_3123);
	assign x_3121 = (x_1496 & x_3120);
	assign x_3118 = (x_1493 & x_3117);
	assign x_3116 = (x_1490 & x_3115);
	assign x_3112 = (x_1487 & x_3111);
	assign x_3110 = (x_1484 & x_3109);
	assign x_3107 = (x_1481 & x_3106);
	assign x_3105 = (x_1478 & x_3104);
	assign x_3099 = (x_3097 & x_3098);
	assign x_3096 = (x_1471 & x_3095);
	assign x_3093 = (x_1468 & x_3092);
	assign x_3091 = (x_1465 & x_3090);
	assign x_3087 = (x_3085 & x_3086);
	assign x_3084 = (x_1458 & x_3083);
	assign x_3081 = (x_1455 & x_3080);
	assign x_3079 = (x_1452 & x_3078);
	assign x_3074 = (x_3072 & x_3073);
	assign x_3071 = (x_1445 & x_3070);
	assign x_3068 = (x_1442 & x_3067);
	assign x_3066 = (x_1439 & x_3065);
	assign x_3062 = (x_1436 & x_3061);
	assign x_3060 = (x_1433 & x_3059);
	assign x_3057 = (x_1430 & x_3056);
	assign x_3055 = (x_1427 & x_3054);
	assign x_3047 = (x_3045 & x_3046);
	assign x_3044 = (x_1420 & x_3043);
	assign x_3041 = (x_1417 & x_3040);
	assign x_3039 = (x_1414 & x_3038);
	assign x_3035 = (x_3033 & x_3034);
	assign x_3032 = (x_1407 & x_3031);
	assign x_3029 = (x_1404 & x_3028);
	assign x_3027 = (x_1401 & x_3026);
	assign x_3022 = (x_3020 & x_3021);
	assign x_3019 = (x_1394 & x_3018);
	assign x_3016 = (x_1391 & x_3015);
	assign x_3014 = (x_1388 & x_3013);
	assign x_3010 = (x_1385 & x_3009);
	assign x_3008 = (x_1382 & x_3007);
	assign x_3005 = (x_1379 & x_3004);
	assign x_3003 = (x_1376 & x_3002);
	assign x_2997 = (x_2995 & x_2996);
	assign x_2994 = (x_1369 & x_2993);
	assign x_2991 = (x_1366 & x_2990);
	assign x_2989 = (x_1363 & x_2988);
	assign x_2985 = (x_2983 & x_2984);
	assign x_2982 = (x_1356 & x_2981);
	assign x_2979 = (x_1353 & x_2978);
	assign x_2977 = (x_1350 & x_2976);
	assign x_2972 = (x_2970 & x_2971);
	assign x_2969 = (x_1343 & x_2968);
	assign x_2966 = (x_1340 & x_2965);
	assign x_2964 = (x_1337 & x_2963);
	assign x_2960 = (x_1334 & x_2959);
	assign x_2958 = (x_1331 & x_2957);
	assign x_2955 = (x_1328 & x_2954);
	assign x_2953 = (x_1325 & x_2952);
	assign x_2946 = (x_2944 & x_2945);
	assign x_2943 = (x_1318 & x_2942);
	assign x_2940 = (x_1315 & x_2939);
	assign x_2938 = (x_1312 & x_2937);
	assign x_2934 = (x_2932 & x_2933);
	assign x_2931 = (x_1305 & x_2930);
	assign x_2928 = (x_1302 & x_2927);
	assign x_2926 = (x_1299 & x_2925);
	assign x_2921 = (x_2919 & x_2920);
	assign x_2918 = (x_1292 & x_2917);
	assign x_2915 = (x_1289 & x_2914);
	assign x_2913 = (x_1286 & x_2912);
	assign x_2909 = (x_1283 & x_2908);
	assign x_2907 = (x_1280 & x_2906);
	assign x_2904 = (x_1277 & x_2903);
	assign x_2902 = (x_1274 & x_2901);
	assign x_2896 = (x_2894 & x_2895);
	assign x_2893 = (x_1267 & x_2892);
	assign x_2890 = (x_1264 & x_2889);
	assign x_2888 = (x_1261 & x_2887);
	assign x_2884 = (x_2882 & x_2883);
	assign x_2881 = (x_1254 & x_2880);
	assign x_2878 = (x_1251 & x_2877);
	assign x_2876 = (x_1248 & x_2875);
	assign x_2871 = (x_2869 & x_2870);
	assign x_2868 = (x_1241 & x_2867);
	assign x_2865 = (x_1238 & x_2864);
	assign x_2863 = (x_1235 & x_2862);
	assign x_2859 = (x_1232 & x_2858);
	assign x_2857 = (x_1229 & x_2856);
	assign x_2854 = (x_1226 & x_2853);
	assign x_2852 = (x_1223 & x_2851);
	assign x_2843 = (x_2841 & x_2842);
	assign x_2840 = (x_1216 & x_2839);
	assign x_2837 = (x_1213 & x_2836);
	assign x_2835 = (x_1210 & x_2834);
	assign x_2831 = (x_2829 & x_2830);
	assign x_2828 = (x_1203 & x_2827);
	assign x_2825 = (x_1200 & x_2824);
	assign x_2823 = (x_1197 & x_2822);
	assign x_2818 = (x_2816 & x_2817);
	assign x_2815 = (x_1190 & x_2814);
	assign x_2812 = (x_1187 & x_2811);
	assign x_2810 = (x_1184 & x_2809);
	assign x_2806 = (x_1181 & x_2805);
	assign x_2804 = (x_1178 & x_2803);
	assign x_2801 = (x_1175 & x_2800);
	assign x_2799 = (x_1172 & x_2798);
	assign x_2793 = (x_2791 & x_2792);
	assign x_2790 = (x_1165 & x_2789);
	assign x_2787 = (x_1162 & x_2786);
	assign x_2785 = (x_1159 & x_2784);
	assign x_2781 = (x_2779 & x_2780);
	assign x_2778 = (x_1152 & x_2777);
	assign x_2775 = (x_1149 & x_2774);
	assign x_2773 = (x_1146 & x_2772);
	assign x_2768 = (x_2766 & x_2767);
	assign x_2765 = (x_1139 & x_2764);
	assign x_2762 = (x_1136 & x_2761);
	assign x_2760 = (x_1133 & x_2759);
	assign x_2756 = (x_1130 & x_2755);
	assign x_2754 = (x_1127 & x_2753);
	assign x_2751 = (x_1124 & x_2750);
	assign x_2749 = (x_1121 & x_2748);
	assign x_2742 = (x_2740 & x_2741);
	assign x_2739 = (x_1114 & x_2738);
	assign x_2736 = (x_1111 & x_2735);
	assign x_2734 = (x_1108 & x_2733);
	assign x_2730 = (x_2728 & x_2729);
	assign x_2727 = (x_1101 & x_2726);
	assign x_2724 = (x_1098 & x_2723);
	assign x_2722 = (x_1095 & x_2721);
	assign x_2717 = (x_2715 & x_2716);
	assign x_2714 = (x_1088 & x_2713);
	assign x_2711 = (x_1085 & x_2710);
	assign x_2709 = (x_1082 & x_2708);
	assign x_2705 = (x_1079 & x_2704);
	assign x_2703 = (x_1076 & x_2702);
	assign x_2700 = (x_1073 & x_2699);
	assign x_2698 = (x_1070 & x_2697);
	assign x_2692 = (x_2690 & x_2691);
	assign x_2689 = (x_1063 & x_2688);
	assign x_2686 = (x_1060 & x_2685);
	assign x_2684 = (x_1057 & x_2683);
	assign x_2680 = (x_2678 & x_2679);
	assign x_2677 = (x_1050 & x_2676);
	assign x_2674 = (x_1047 & x_2673);
	assign x_2672 = (x_1044 & x_2671);
	assign x_2667 = (x_2665 & x_2666);
	assign x_2664 = (x_1037 & x_2663);
	assign x_2661 = (x_1034 & x_2660);
	assign x_2659 = (x_1031 & x_2658);
	assign x_2655 = (x_1028 & x_2654);
	assign x_2653 = (x_1025 & x_2652);
	assign x_2650 = (x_1022 & x_2649);
	assign x_2648 = (x_1019 & x_2647);
	assign x_2640 = (x_2638 & x_2639);
	assign x_2637 = (x_1012 & x_2636);
	assign x_2634 = (x_1009 & x_2633);
	assign x_2632 = (x_1006 & x_2631);
	assign x_2628 = (x_2626 & x_2627);
	assign x_2625 = (x_999 & x_2624);
	assign x_2622 = (x_996 & x_2621);
	assign x_2620 = (x_993 & x_2619);
	assign x_2615 = (x_2613 & x_2614);
	assign x_2612 = (x_986 & x_2611);
	assign x_2609 = (x_983 & x_2608);
	assign x_2607 = (x_980 & x_2606);
	assign x_2603 = (x_977 & x_2602);
	assign x_2601 = (x_974 & x_2600);
	assign x_2598 = (x_971 & x_2597);
	assign x_2596 = (x_968 & x_2595);
	assign x_2590 = (x_2588 & x_2589);
	assign x_2587 = (x_961 & x_2586);
	assign x_2584 = (x_958 & x_2583);
	assign x_2582 = (x_955 & x_2581);
	assign x_2578 = (x_2576 & x_2577);
	assign x_2575 = (x_948 & x_2574);
	assign x_2572 = (x_945 & x_2571);
	assign x_2570 = (x_942 & x_2569);
	assign x_2565 = (x_2563 & x_2564);
	assign x_2562 = (x_935 & x_2561);
	assign x_2559 = (x_932 & x_2558);
	assign x_2557 = (x_929 & x_2556);
	assign x_2553 = (x_926 & x_2552);
	assign x_2551 = (x_923 & x_2550);
	assign x_2548 = (x_920 & x_2547);
	assign x_2546 = (x_917 & x_2545);
	assign x_2539 = (x_2537 & x_2538);
	assign x_2536 = (x_910 & x_2535);
	assign x_2533 = (x_907 & x_2532);
	assign x_2531 = (x_904 & x_2530);
	assign x_2527 = (x_2525 & x_2526);
	assign x_2524 = (x_897 & x_2523);
	assign x_2521 = (x_894 & x_2520);
	assign x_2519 = (x_891 & x_2518);
	assign x_2514 = (x_2512 & x_2513);
	assign x_2511 = (x_884 & x_2510);
	assign x_2508 = (x_881 & x_2507);
	assign x_2506 = (x_878 & x_2505);
	assign x_2502 = (x_875 & x_2501);
	assign x_2500 = (x_872 & x_2499);
	assign x_2497 = (x_869 & x_2496);
	assign x_2495 = (x_866 & x_2494);
	assign x_2489 = (x_2487 & x_2488);
	assign x_2486 = (x_859 & x_2485);
	assign x_2483 = (x_856 & x_2482);
	assign x_2481 = (x_853 & x_2480);
	assign x_2477 = (x_850 & x_2476);
	assign x_2475 = (x_847 & x_2474);
	assign x_2472 = (x_844 & x_2471);
	assign x_2470 = (x_841 & x_2469);
	assign x_2465 = (x_2463 & x_2464);
	assign x_2462 = (x_834 & x_2461);
	assign x_2459 = (x_831 & x_2458);
	assign x_2457 = (x_828 & x_2456);
	assign x_2453 = (x_825 & x_2452);
	assign x_2451 = (x_822 & x_2450);
	assign x_2448 = (x_819 & x_2447);
	assign x_2446 = (x_816 & x_2445);
	assign x_2436 = (x_2434 & x_2435);
	assign x_2433 = (x_809 & x_2432);
	assign x_2430 = (x_806 & x_2429);
	assign x_2428 = (x_803 & x_2427);
	assign x_2424 = (x_2422 & x_2423);
	assign x_2421 = (x_796 & x_2420);
	assign x_2418 = (x_793 & x_2417);
	assign x_2416 = (x_790 & x_2415);
	assign x_2411 = (x_2409 & x_2410);
	assign x_2408 = (x_783 & x_2407);
	assign x_2405 = (x_780 & x_2404);
	assign x_2403 = (x_777 & x_2402);
	assign x_2399 = (x_774 & x_2398);
	assign x_2397 = (x_771 & x_2396);
	assign x_2394 = (x_768 & x_2393);
	assign x_2392 = (x_765 & x_2391);
	assign x_2386 = (x_2384 & x_2385);
	assign x_2383 = (x_758 & x_2382);
	assign x_2380 = (x_755 & x_2379);
	assign x_2378 = (x_752 & x_2377);
	assign x_2374 = (x_2372 & x_2373);
	assign x_2371 = (x_745 & x_2370);
	assign x_2368 = (x_742 & x_2367);
	assign x_2366 = (x_739 & x_2365);
	assign x_2361 = (x_2359 & x_2360);
	assign x_2358 = (x_732 & x_2357);
	assign x_2355 = (x_729 & x_2354);
	assign x_2353 = (x_726 & x_2352);
	assign x_2349 = (x_723 & x_2348);
	assign x_2347 = (x_720 & x_2346);
	assign x_2344 = (x_717 & x_2343);
	assign x_2342 = (x_714 & x_2341);
	assign x_2335 = (x_2333 & x_2334);
	assign x_2332 = (x_707 & x_2331);
	assign x_2329 = (x_704 & x_2328);
	assign x_2327 = (x_701 & x_2326);
	assign x_2323 = (x_2321 & x_2322);
	assign x_2320 = (x_694 & x_2319);
	assign x_2317 = (x_691 & x_2316);
	assign x_2315 = (x_688 & x_2314);
	assign x_2310 = (x_2308 & x_2309);
	assign x_2307 = (x_681 & x_2306);
	assign x_2304 = (x_678 & x_2303);
	assign x_2302 = (x_675 & x_2301);
	assign x_2298 = (x_672 & x_2297);
	assign x_2296 = (x_669 & x_2295);
	assign x_2293 = (x_666 & x_2292);
	assign x_2291 = (x_663 & x_2290);
	assign x_2285 = (x_2283 & x_2284);
	assign x_2282 = (x_656 & x_2281);
	assign x_2279 = (x_653 & x_2278);
	assign x_2277 = (x_650 & x_2276);
	assign x_2273 = (x_2271 & x_2272);
	assign x_2270 = (x_643 & x_2269);
	assign x_2267 = (x_640 & x_2266);
	assign x_2265 = (x_637 & x_2264);
	assign x_2260 = (x_2258 & x_2259);
	assign x_2257 = (x_630 & x_2256);
	assign x_2254 = (x_627 & x_2253);
	assign x_2252 = (x_624 & x_2251);
	assign x_2248 = (x_621 & x_2247);
	assign x_2246 = (x_618 & x_2245);
	assign x_2243 = (x_615 & x_2242);
	assign x_2241 = (x_612 & x_2240);
	assign x_2233 = (x_2231 & x_2232);
	assign x_2230 = (x_605 & x_2229);
	assign x_2227 = (x_602 & x_2226);
	assign x_2225 = (x_599 & x_2224);
	assign x_2221 = (x_2219 & x_2220);
	assign x_2218 = (x_592 & x_2217);
	assign x_2215 = (x_589 & x_2214);
	assign x_2213 = (x_586 & x_2212);
	assign x_2208 = (x_2206 & x_2207);
	assign x_2205 = (x_579 & x_2204);
	assign x_2202 = (x_576 & x_2201);
	assign x_2200 = (x_573 & x_2199);
	assign x_2196 = (x_570 & x_2195);
	assign x_2194 = (x_567 & x_2193);
	assign x_2191 = (x_564 & x_2190);
	assign x_2189 = (x_561 & x_2188);
	assign x_2183 = (x_2181 & x_2182);
	assign x_2180 = (x_554 & x_2179);
	assign x_2177 = (x_551 & x_2176);
	assign x_2175 = (x_548 & x_2174);
	assign x_2171 = (x_2169 & x_2170);
	assign x_2168 = (x_541 & x_2167);
	assign x_2165 = (x_538 & x_2164);
	assign x_2163 = (x_535 & x_2162);
	assign x_2158 = (x_2156 & x_2157);
	assign x_2155 = (x_528 & x_2154);
	assign x_2152 = (x_525 & x_2151);
	assign x_2150 = (x_522 & x_2149);
	assign x_2146 = (x_519 & x_2145);
	assign x_2144 = (x_516 & x_2143);
	assign x_2141 = (x_513 & x_2140);
	assign x_2139 = (x_510 & x_2138);
	assign x_2132 = (x_2130 & x_2131);
	assign x_2129 = (x_503 & x_2128);
	assign x_2126 = (x_500 & x_2125);
	assign x_2124 = (x_497 & x_2123);
	assign x_2120 = (x_2118 & x_2119);
	assign x_2117 = (x_490 & x_2116);
	assign x_2114 = (x_487 & x_2113);
	assign x_2112 = (x_484 & x_2111);
	assign x_2107 = (x_2105 & x_2106);
	assign x_2104 = (x_477 & x_2103);
	assign x_2101 = (x_474 & x_2100);
	assign x_2099 = (x_471 & x_2098);
	assign x_2095 = (x_468 & x_2094);
	assign x_2093 = (x_465 & x_2092);
	assign x_2090 = (x_462 & x_2089);
	assign x_2088 = (x_459 & x_2087);
	assign x_2082 = (x_2080 & x_2081);
	assign x_2079 = (x_452 & x_2078);
	assign x_2076 = (x_449 & x_2075);
	assign x_2074 = (x_446 & x_2073);
	assign x_2070 = (x_2068 & x_2069);
	assign x_2067 = (x_439 & x_2066);
	assign x_2064 = (x_436 & x_2063);
	assign x_2062 = (x_433 & x_2061);
	assign x_2057 = (x_2055 & x_2056);
	assign x_2054 = (x_426 & x_2053);
	assign x_2051 = (x_423 & x_2050);
	assign x_2049 = (x_420 & x_2048);
	assign x_2045 = (x_417 & x_2044);
	assign x_2043 = (x_414 & x_2042);
	assign x_2040 = (x_411 & x_2039);
	assign x_2038 = (x_408 & x_2037);
	assign x_2029 = (x_2027 & x_2028);
	assign x_2026 = (x_401 & x_2025);
	assign x_2023 = (x_398 & x_2022);
	assign x_2021 = (x_395 & x_2020);
	assign x_2017 = (x_2015 & x_2016);
	assign x_2014 = (x_388 & x_2013);
	assign x_2011 = (x_385 & x_2010);
	assign x_2009 = (x_382 & x_2008);
	assign x_2004 = (x_2002 & x_2003);
	assign x_2001 = (x_375 & x_2000);
	assign x_1998 = (x_372 & x_1997);
	assign x_1996 = (x_369 & x_1995);
	assign x_1992 = (x_366 & x_1991);
	assign x_1990 = (x_363 & x_1989);
	assign x_1987 = (x_360 & x_1986);
	assign x_1985 = (x_357 & x_1984);
	assign x_1979 = (x_1977 & x_1978);
	assign x_1976 = (x_350 & x_1975);
	assign x_1973 = (x_347 & x_1972);
	assign x_1971 = (x_344 & x_1970);
	assign x_1967 = (x_1965 & x_1966);
	assign x_1964 = (x_337 & x_1963);
	assign x_1961 = (x_334 & x_1960);
	assign x_1959 = (x_331 & x_1958);
	assign x_1954 = (x_1952 & x_1953);
	assign x_1951 = (x_324 & x_1950);
	assign x_1948 = (x_321 & x_1947);
	assign x_1946 = (x_318 & x_1945);
	assign x_1942 = (x_315 & x_1941);
	assign x_1940 = (x_312 & x_1939);
	assign x_1937 = (x_309 & x_1936);
	assign x_1935 = (x_306 & x_1934);
	assign x_1928 = (x_1926 & x_1927);
	assign x_1925 = (x_299 & x_1924);
	assign x_1922 = (x_296 & x_1921);
	assign x_1920 = (x_293 & x_1919);
	assign x_1916 = (x_1914 & x_1915);
	assign x_1913 = (x_286 & x_1912);
	assign x_1910 = (x_283 & x_1909);
	assign x_1908 = (x_280 & x_1907);
	assign x_1903 = (x_1901 & x_1902);
	assign x_1900 = (x_273 & x_1899);
	assign x_1897 = (x_270 & x_1896);
	assign x_1895 = (x_267 & x_1894);
	assign x_1891 = (x_264 & x_1890);
	assign x_1889 = (x_261 & x_1888);
	assign x_1886 = (x_258 & x_1885);
	assign x_1884 = (x_255 & x_1883);
	assign x_1878 = (x_1876 & x_1877);
	assign x_1875 = (x_248 & x_1874);
	assign x_1872 = (x_245 & x_1871);
	assign x_1870 = (x_242 & x_1869);
	assign x_1866 = (x_1864 & x_1865);
	assign x_1863 = (x_235 & x_1862);
	assign x_1860 = (x_232 & x_1859);
	assign x_1858 = (x_229 & x_1857);
	assign x_1853 = (x_1851 & x_1852);
	assign x_1850 = (x_222 & x_1849);
	assign x_1847 = (x_219 & x_1846);
	assign x_1845 = (x_216 & x_1844);
	assign x_1841 = (x_213 & x_1840);
	assign x_1839 = (x_210 & x_1838);
	assign x_1836 = (x_207 & x_1835);
	assign x_1834 = (x_204 & x_1833);
	assign x_1826 = (x_1824 & x_1825);
	assign x_1823 = (x_197 & x_1822);
	assign x_1820 = (x_194 & x_1819);
	assign x_1818 = (x_191 & x_1817);
	assign x_1814 = (x_1812 & x_1813);
	assign x_1811 = (x_184 & x_1810);
	assign x_1808 = (x_181 & x_1807);
	assign x_1806 = (x_178 & x_1805);
	assign x_1801 = (x_1799 & x_1800);
	assign x_1798 = (x_171 & x_1797);
	assign x_1795 = (x_168 & x_1794);
	assign x_1793 = (x_165 & x_1792);
	assign x_1789 = (x_162 & x_1788);
	assign x_1787 = (x_159 & x_1786);
	assign x_1784 = (x_156 & x_1783);
	assign x_1782 = (x_153 & x_1781);
	assign x_1776 = (x_1774 & x_1775);
	assign x_1773 = (x_146 & x_1772);
	assign x_1770 = (x_143 & x_1769);
	assign x_1768 = (x_140 & x_1767);
	assign x_1764 = (x_1762 & x_1763);
	assign x_1761 = (x_133 & x_1760);
	assign x_1758 = (x_130 & x_1757);
	assign x_1756 = (x_127 & x_1755);
	assign x_1751 = (x_1749 & x_1750);
	assign x_1748 = (x_120 & x_1747);
	assign x_1745 = (x_117 & x_1744);
	assign x_1743 = (x_114 & x_1742);
	assign x_1739 = (x_111 & x_1738);
	assign x_1737 = (x_108 & x_1736);
	assign x_1734 = (x_105 & x_1733);
	assign x_1732 = (x_102 & x_1731);
	assign x_1725 = (x_1723 & x_1724);
	assign x_1722 = (x_95 & x_1721);
	assign x_1719 = (x_92 & x_1718);
	assign x_1717 = (x_89 & x_1716);
	assign x_1713 = (x_1711 & x_1712);
	assign x_1710 = (x_82 & x_1709);
	assign x_1707 = (x_79 & x_1706);
	assign x_1705 = (x_76 & x_1704);
	assign x_1700 = (x_1698 & x_1699);
	assign x_1697 = (x_69 & x_1696);
	assign x_1694 = (x_66 & x_1693);
	assign x_1692 = (x_63 & x_1691);
	assign x_1688 = (x_60 & x_1687);
	assign x_1686 = (x_57 & x_1685);
	assign x_1683 = (x_54 & x_1682);
	assign x_1681 = (x_51 & x_1680);
	assign x_1675 = (x_1673 & x_1674);
	assign x_1672 = (x_44 & x_1671);
	assign x_1669 = (x_41 & x_1668);
	assign x_1667 = (x_38 & x_1666);
	assign x_1663 = (x_35 & x_1662);
	assign x_1661 = (x_32 & x_1660);
	assign x_1658 = (x_29 & x_1657);
	assign x_1656 = (x_26 & x_1655);
	assign x_1651 = (x_1649 & x_1650);
	assign x_1648 = (x_19 & x_1647);
	assign x_1645 = (x_16 & x_1644);
	assign x_1643 = (x_13 & x_1642);
	assign x_1639 = (x_10 & x_1638);
	assign x_1637 = (x_7 & x_1636);
	assign x_1634 = (x_4 & x_1633);
	assign x_1632 = (x_1 & x_1631);
	assign x_3251 = (x_3247 & x_3250);
	assign x_3245 = (x_3242 & x_3244);
	assign x_3239 = (x_3235 & x_3238);
	assign x_3233 = (x_3230 & x_3232);
	assign x_3226 = (x_3222 & x_3225);
	assign x_3220 = (x_3217 & x_3219);
	assign x_3214 = (x_3211 & x_3213);
	assign x_3209 = (x_3206 & x_3208);
	assign x_3201 = (x_3197 & x_3200);
	assign x_3195 = (x_3192 & x_3194);
	assign x_3189 = (x_3185 & x_3188);
	assign x_3183 = (x_3180 & x_3182);
	assign x_3176 = (x_3172 & x_3175);
	assign x_3170 = (x_3167 & x_3169);
	assign x_3164 = (x_3161 & x_3163);
	assign x_3159 = (x_3156 & x_3158);
	assign x_3150 = (x_3146 & x_3149);
	assign x_3144 = (x_3141 & x_3143);
	assign x_3138 = (x_3134 & x_3137);
	assign x_3132 = (x_3129 & x_3131);
	assign x_3125 = (x_3121 & x_3124);
	assign x_3119 = (x_3116 & x_3118);
	assign x_3113 = (x_3110 & x_3112);
	assign x_3108 = (x_3105 & x_3107);
	assign x_3100 = (x_3096 & x_3099);
	assign x_3094 = (x_3091 & x_3093);
	assign x_3088 = (x_3084 & x_3087);
	assign x_3082 = (x_3079 & x_3081);
	assign x_3075 = (x_3071 & x_3074);
	assign x_3069 = (x_3066 & x_3068);
	assign x_3063 = (x_3060 & x_3062);
	assign x_3058 = (x_3055 & x_3057);
	assign x_3048 = (x_3044 & x_3047);
	assign x_3042 = (x_3039 & x_3041);
	assign x_3036 = (x_3032 & x_3035);
	assign x_3030 = (x_3027 & x_3029);
	assign x_3023 = (x_3019 & x_3022);
	assign x_3017 = (x_3014 & x_3016);
	assign x_3011 = (x_3008 & x_3010);
	assign x_3006 = (x_3003 & x_3005);
	assign x_2998 = (x_2994 & x_2997);
	assign x_2992 = (x_2989 & x_2991);
	assign x_2986 = (x_2982 & x_2985);
	assign x_2980 = (x_2977 & x_2979);
	assign x_2973 = (x_2969 & x_2972);
	assign x_2967 = (x_2964 & x_2966);
	assign x_2961 = (x_2958 & x_2960);
	assign x_2956 = (x_2953 & x_2955);
	assign x_2947 = (x_2943 & x_2946);
	assign x_2941 = (x_2938 & x_2940);
	assign x_2935 = (x_2931 & x_2934);
	assign x_2929 = (x_2926 & x_2928);
	assign x_2922 = (x_2918 & x_2921);
	assign x_2916 = (x_2913 & x_2915);
	assign x_2910 = (x_2907 & x_2909);
	assign x_2905 = (x_2902 & x_2904);
	assign x_2897 = (x_2893 & x_2896);
	assign x_2891 = (x_2888 & x_2890);
	assign x_2885 = (x_2881 & x_2884);
	assign x_2879 = (x_2876 & x_2878);
	assign x_2872 = (x_2868 & x_2871);
	assign x_2866 = (x_2863 & x_2865);
	assign x_2860 = (x_2857 & x_2859);
	assign x_2855 = (x_2852 & x_2854);
	assign x_2844 = (x_2840 & x_2843);
	assign x_2838 = (x_2835 & x_2837);
	assign x_2832 = (x_2828 & x_2831);
	assign x_2826 = (x_2823 & x_2825);
	assign x_2819 = (x_2815 & x_2818);
	assign x_2813 = (x_2810 & x_2812);
	assign x_2807 = (x_2804 & x_2806);
	assign x_2802 = (x_2799 & x_2801);
	assign x_2794 = (x_2790 & x_2793);
	assign x_2788 = (x_2785 & x_2787);
	assign x_2782 = (x_2778 & x_2781);
	assign x_2776 = (x_2773 & x_2775);
	assign x_2769 = (x_2765 & x_2768);
	assign x_2763 = (x_2760 & x_2762);
	assign x_2757 = (x_2754 & x_2756);
	assign x_2752 = (x_2749 & x_2751);
	assign x_2743 = (x_2739 & x_2742);
	assign x_2737 = (x_2734 & x_2736);
	assign x_2731 = (x_2727 & x_2730);
	assign x_2725 = (x_2722 & x_2724);
	assign x_2718 = (x_2714 & x_2717);
	assign x_2712 = (x_2709 & x_2711);
	assign x_2706 = (x_2703 & x_2705);
	assign x_2701 = (x_2698 & x_2700);
	assign x_2693 = (x_2689 & x_2692);
	assign x_2687 = (x_2684 & x_2686);
	assign x_2681 = (x_2677 & x_2680);
	assign x_2675 = (x_2672 & x_2674);
	assign x_2668 = (x_2664 & x_2667);
	assign x_2662 = (x_2659 & x_2661);
	assign x_2656 = (x_2653 & x_2655);
	assign x_2651 = (x_2648 & x_2650);
	assign x_2641 = (x_2637 & x_2640);
	assign x_2635 = (x_2632 & x_2634);
	assign x_2629 = (x_2625 & x_2628);
	assign x_2623 = (x_2620 & x_2622);
	assign x_2616 = (x_2612 & x_2615);
	assign x_2610 = (x_2607 & x_2609);
	assign x_2604 = (x_2601 & x_2603);
	assign x_2599 = (x_2596 & x_2598);
	assign x_2591 = (x_2587 & x_2590);
	assign x_2585 = (x_2582 & x_2584);
	assign x_2579 = (x_2575 & x_2578);
	assign x_2573 = (x_2570 & x_2572);
	assign x_2566 = (x_2562 & x_2565);
	assign x_2560 = (x_2557 & x_2559);
	assign x_2554 = (x_2551 & x_2553);
	assign x_2549 = (x_2546 & x_2548);
	assign x_2540 = (x_2536 & x_2539);
	assign x_2534 = (x_2531 & x_2533);
	assign x_2528 = (x_2524 & x_2527);
	assign x_2522 = (x_2519 & x_2521);
	assign x_2515 = (x_2511 & x_2514);
	assign x_2509 = (x_2506 & x_2508);
	assign x_2503 = (x_2500 & x_2502);
	assign x_2498 = (x_2495 & x_2497);
	assign x_2490 = (x_2486 & x_2489);
	assign x_2484 = (x_2481 & x_2483);
	assign x_2478 = (x_2475 & x_2477);
	assign x_2473 = (x_2470 & x_2472);
	assign x_2466 = (x_2462 & x_2465);
	assign x_2460 = (x_2457 & x_2459);
	assign x_2454 = (x_2451 & x_2453);
	assign x_2449 = (x_2446 & x_2448);
	assign x_2437 = (x_2433 & x_2436);
	assign x_2431 = (x_2428 & x_2430);
	assign x_2425 = (x_2421 & x_2424);
	assign x_2419 = (x_2416 & x_2418);
	assign x_2412 = (x_2408 & x_2411);
	assign x_2406 = (x_2403 & x_2405);
	assign x_2400 = (x_2397 & x_2399);
	assign x_2395 = (x_2392 & x_2394);
	assign x_2387 = (x_2383 & x_2386);
	assign x_2381 = (x_2378 & x_2380);
	assign x_2375 = (x_2371 & x_2374);
	assign x_2369 = (x_2366 & x_2368);
	assign x_2362 = (x_2358 & x_2361);
	assign x_2356 = (x_2353 & x_2355);
	assign x_2350 = (x_2347 & x_2349);
	assign x_2345 = (x_2342 & x_2344);
	assign x_2336 = (x_2332 & x_2335);
	assign x_2330 = (x_2327 & x_2329);
	assign x_2324 = (x_2320 & x_2323);
	assign x_2318 = (x_2315 & x_2317);
	assign x_2311 = (x_2307 & x_2310);
	assign x_2305 = (x_2302 & x_2304);
	assign x_2299 = (x_2296 & x_2298);
	assign x_2294 = (x_2291 & x_2293);
	assign x_2286 = (x_2282 & x_2285);
	assign x_2280 = (x_2277 & x_2279);
	assign x_2274 = (x_2270 & x_2273);
	assign x_2268 = (x_2265 & x_2267);
	assign x_2261 = (x_2257 & x_2260);
	assign x_2255 = (x_2252 & x_2254);
	assign x_2249 = (x_2246 & x_2248);
	assign x_2244 = (x_2241 & x_2243);
	assign x_2234 = (x_2230 & x_2233);
	assign x_2228 = (x_2225 & x_2227);
	assign x_2222 = (x_2218 & x_2221);
	assign x_2216 = (x_2213 & x_2215);
	assign x_2209 = (x_2205 & x_2208);
	assign x_2203 = (x_2200 & x_2202);
	assign x_2197 = (x_2194 & x_2196);
	assign x_2192 = (x_2189 & x_2191);
	assign x_2184 = (x_2180 & x_2183);
	assign x_2178 = (x_2175 & x_2177);
	assign x_2172 = (x_2168 & x_2171);
	assign x_2166 = (x_2163 & x_2165);
	assign x_2159 = (x_2155 & x_2158);
	assign x_2153 = (x_2150 & x_2152);
	assign x_2147 = (x_2144 & x_2146);
	assign x_2142 = (x_2139 & x_2141);
	assign x_2133 = (x_2129 & x_2132);
	assign x_2127 = (x_2124 & x_2126);
	assign x_2121 = (x_2117 & x_2120);
	assign x_2115 = (x_2112 & x_2114);
	assign x_2108 = (x_2104 & x_2107);
	assign x_2102 = (x_2099 & x_2101);
	assign x_2096 = (x_2093 & x_2095);
	assign x_2091 = (x_2088 & x_2090);
	assign x_2083 = (x_2079 & x_2082);
	assign x_2077 = (x_2074 & x_2076);
	assign x_2071 = (x_2067 & x_2070);
	assign x_2065 = (x_2062 & x_2064);
	assign x_2058 = (x_2054 & x_2057);
	assign x_2052 = (x_2049 & x_2051);
	assign x_2046 = (x_2043 & x_2045);
	assign x_2041 = (x_2038 & x_2040);
	assign x_2030 = (x_2026 & x_2029);
	assign x_2024 = (x_2021 & x_2023);
	assign x_2018 = (x_2014 & x_2017);
	assign x_2012 = (x_2009 & x_2011);
	assign x_2005 = (x_2001 & x_2004);
	assign x_1999 = (x_1996 & x_1998);
	assign x_1993 = (x_1990 & x_1992);
	assign x_1988 = (x_1985 & x_1987);
	assign x_1980 = (x_1976 & x_1979);
	assign x_1974 = (x_1971 & x_1973);
	assign x_1968 = (x_1964 & x_1967);
	assign x_1962 = (x_1959 & x_1961);
	assign x_1955 = (x_1951 & x_1954);
	assign x_1949 = (x_1946 & x_1948);
	assign x_1943 = (x_1940 & x_1942);
	assign x_1938 = (x_1935 & x_1937);
	assign x_1929 = (x_1925 & x_1928);
	assign x_1923 = (x_1920 & x_1922);
	assign x_1917 = (x_1913 & x_1916);
	assign x_1911 = (x_1908 & x_1910);
	assign x_1904 = (x_1900 & x_1903);
	assign x_1898 = (x_1895 & x_1897);
	assign x_1892 = (x_1889 & x_1891);
	assign x_1887 = (x_1884 & x_1886);
	assign x_1879 = (x_1875 & x_1878);
	assign x_1873 = (x_1870 & x_1872);
	assign x_1867 = (x_1863 & x_1866);
	assign x_1861 = (x_1858 & x_1860);
	assign x_1854 = (x_1850 & x_1853);
	assign x_1848 = (x_1845 & x_1847);
	assign x_1842 = (x_1839 & x_1841);
	assign x_1837 = (x_1834 & x_1836);
	assign x_1827 = (x_1823 & x_1826);
	assign x_1821 = (x_1818 & x_1820);
	assign x_1815 = (x_1811 & x_1814);
	assign x_1809 = (x_1806 & x_1808);
	assign x_1802 = (x_1798 & x_1801);
	assign x_1796 = (x_1793 & x_1795);
	assign x_1790 = (x_1787 & x_1789);
	assign x_1785 = (x_1782 & x_1784);
	assign x_1777 = (x_1773 & x_1776);
	assign x_1771 = (x_1768 & x_1770);
	assign x_1765 = (x_1761 & x_1764);
	assign x_1759 = (x_1756 & x_1758);
	assign x_1752 = (x_1748 & x_1751);
	assign x_1746 = (x_1743 & x_1745);
	assign x_1740 = (x_1737 & x_1739);
	assign x_1735 = (x_1732 & x_1734);
	assign x_1726 = (x_1722 & x_1725);
	assign x_1720 = (x_1717 & x_1719);
	assign x_1714 = (x_1710 & x_1713);
	assign x_1708 = (x_1705 & x_1707);
	assign x_1701 = (x_1697 & x_1700);
	assign x_1695 = (x_1692 & x_1694);
	assign x_1689 = (x_1686 & x_1688);
	assign x_1684 = (x_1681 & x_1683);
	assign x_1676 = (x_1672 & x_1675);
	assign x_1670 = (x_1667 & x_1669);
	assign x_1664 = (x_1661 & x_1663);
	assign x_1659 = (x_1656 & x_1658);
	assign x_1652 = (x_1648 & x_1651);
	assign x_1646 = (x_1643 & x_1645);
	assign x_1640 = (x_1637 & x_1639);
	assign x_1635 = (x_1632 & x_1634);
	assign x_3252 = (x_3245 & x_3251);
	assign x_3240 = (x_3233 & x_3239);
	assign x_3227 = (x_3220 & x_3226);
	assign x_3215 = (x_3209 & x_3214);
	assign x_3202 = (x_3195 & x_3201);
	assign x_3190 = (x_3183 & x_3189);
	assign x_3177 = (x_3170 & x_3176);
	assign x_3165 = (x_3159 & x_3164);
	assign x_3151 = (x_3144 & x_3150);
	assign x_3139 = (x_3132 & x_3138);
	assign x_3126 = (x_3119 & x_3125);
	assign x_3114 = (x_3108 & x_3113);
	assign x_3101 = (x_3094 & x_3100);
	assign x_3089 = (x_3082 & x_3088);
	assign x_3076 = (x_3069 & x_3075);
	assign x_3064 = (x_3058 & x_3063);
	assign x_3049 = (x_3042 & x_3048);
	assign x_3037 = (x_3030 & x_3036);
	assign x_3024 = (x_3017 & x_3023);
	assign x_3012 = (x_3006 & x_3011);
	assign x_2999 = (x_2992 & x_2998);
	assign x_2987 = (x_2980 & x_2986);
	assign x_2974 = (x_2967 & x_2973);
	assign x_2962 = (x_2956 & x_2961);
	assign x_2948 = (x_2941 & x_2947);
	assign x_2936 = (x_2929 & x_2935);
	assign x_2923 = (x_2916 & x_2922);
	assign x_2911 = (x_2905 & x_2910);
	assign x_2898 = (x_2891 & x_2897);
	assign x_2886 = (x_2879 & x_2885);
	assign x_2873 = (x_2866 & x_2872);
	assign x_2861 = (x_2855 & x_2860);
	assign x_2845 = (x_2838 & x_2844);
	assign x_2833 = (x_2826 & x_2832);
	assign x_2820 = (x_2813 & x_2819);
	assign x_2808 = (x_2802 & x_2807);
	assign x_2795 = (x_2788 & x_2794);
	assign x_2783 = (x_2776 & x_2782);
	assign x_2770 = (x_2763 & x_2769);
	assign x_2758 = (x_2752 & x_2757);
	assign x_2744 = (x_2737 & x_2743);
	assign x_2732 = (x_2725 & x_2731);
	assign x_2719 = (x_2712 & x_2718);
	assign x_2707 = (x_2701 & x_2706);
	assign x_2694 = (x_2687 & x_2693);
	assign x_2682 = (x_2675 & x_2681);
	assign x_2669 = (x_2662 & x_2668);
	assign x_2657 = (x_2651 & x_2656);
	assign x_2642 = (x_2635 & x_2641);
	assign x_2630 = (x_2623 & x_2629);
	assign x_2617 = (x_2610 & x_2616);
	assign x_2605 = (x_2599 & x_2604);
	assign x_2592 = (x_2585 & x_2591);
	assign x_2580 = (x_2573 & x_2579);
	assign x_2567 = (x_2560 & x_2566);
	assign x_2555 = (x_2549 & x_2554);
	assign x_2541 = (x_2534 & x_2540);
	assign x_2529 = (x_2522 & x_2528);
	assign x_2516 = (x_2509 & x_2515);
	assign x_2504 = (x_2498 & x_2503);
	assign x_2491 = (x_2484 & x_2490);
	assign x_2479 = (x_2473 & x_2478);
	assign x_2467 = (x_2460 & x_2466);
	assign x_2455 = (x_2449 & x_2454);
	assign x_2438 = (x_2431 & x_2437);
	assign x_2426 = (x_2419 & x_2425);
	assign x_2413 = (x_2406 & x_2412);
	assign x_2401 = (x_2395 & x_2400);
	assign x_2388 = (x_2381 & x_2387);
	assign x_2376 = (x_2369 & x_2375);
	assign x_2363 = (x_2356 & x_2362);
	assign x_2351 = (x_2345 & x_2350);
	assign x_2337 = (x_2330 & x_2336);
	assign x_2325 = (x_2318 & x_2324);
	assign x_2312 = (x_2305 & x_2311);
	assign x_2300 = (x_2294 & x_2299);
	assign x_2287 = (x_2280 & x_2286);
	assign x_2275 = (x_2268 & x_2274);
	assign x_2262 = (x_2255 & x_2261);
	assign x_2250 = (x_2244 & x_2249);
	assign x_2235 = (x_2228 & x_2234);
	assign x_2223 = (x_2216 & x_2222);
	assign x_2210 = (x_2203 & x_2209);
	assign x_2198 = (x_2192 & x_2197);
	assign x_2185 = (x_2178 & x_2184);
	assign x_2173 = (x_2166 & x_2172);
	assign x_2160 = (x_2153 & x_2159);
	assign x_2148 = (x_2142 & x_2147);
	assign x_2134 = (x_2127 & x_2133);
	assign x_2122 = (x_2115 & x_2121);
	assign x_2109 = (x_2102 & x_2108);
	assign x_2097 = (x_2091 & x_2096);
	assign x_2084 = (x_2077 & x_2083);
	assign x_2072 = (x_2065 & x_2071);
	assign x_2059 = (x_2052 & x_2058);
	assign x_2047 = (x_2041 & x_2046);
	assign x_2031 = (x_2024 & x_2030);
	assign x_2019 = (x_2012 & x_2018);
	assign x_2006 = (x_1999 & x_2005);
	assign x_1994 = (x_1988 & x_1993);
	assign x_1981 = (x_1974 & x_1980);
	assign x_1969 = (x_1962 & x_1968);
	assign x_1956 = (x_1949 & x_1955);
	assign x_1944 = (x_1938 & x_1943);
	assign x_1930 = (x_1923 & x_1929);
	assign x_1918 = (x_1911 & x_1917);
	assign x_1905 = (x_1898 & x_1904);
	assign x_1893 = (x_1887 & x_1892);
	assign x_1880 = (x_1873 & x_1879);
	assign x_1868 = (x_1861 & x_1867);
	assign x_1855 = (x_1848 & x_1854);
	assign x_1843 = (x_1837 & x_1842);
	assign x_1828 = (x_1821 & x_1827);
	assign x_1816 = (x_1809 & x_1815);
	assign x_1803 = (x_1796 & x_1802);
	assign x_1791 = (x_1785 & x_1790);
	assign x_1778 = (x_1771 & x_1777);
	assign x_1766 = (x_1759 & x_1765);
	assign x_1753 = (x_1746 & x_1752);
	assign x_1741 = (x_1735 & x_1740);
	assign x_1727 = (x_1720 & x_1726);
	assign x_1715 = (x_1708 & x_1714);
	assign x_1702 = (x_1695 & x_1701);
	assign x_1690 = (x_1684 & x_1689);
	assign x_1677 = (x_1670 & x_1676);
	assign x_1665 = (x_1659 & x_1664);
	assign x_1653 = (x_1646 & x_1652);
	assign x_1641 = (x_1635 & x_1640);
	assign x_3253 = (x_3240 & x_3252);
	assign x_3228 = (x_3215 & x_3227);
	assign x_3203 = (x_3190 & x_3202);
	assign x_3178 = (x_3165 & x_3177);
	assign x_3152 = (x_3139 & x_3151);
	assign x_3127 = (x_3114 & x_3126);
	assign x_3102 = (x_3089 & x_3101);
	assign x_3077 = (x_3064 & x_3076);
	assign x_3050 = (x_3037 & x_3049);
	assign x_3025 = (x_3012 & x_3024);
	assign x_3000 = (x_2987 & x_2999);
	assign x_2975 = (x_2962 & x_2974);
	assign x_2949 = (x_2936 & x_2948);
	assign x_2924 = (x_2911 & x_2923);
	assign x_2899 = (x_2886 & x_2898);
	assign x_2874 = (x_2861 & x_2873);
	assign x_2846 = (x_2833 & x_2845);
	assign x_2821 = (x_2808 & x_2820);
	assign x_2796 = (x_2783 & x_2795);
	assign x_2771 = (x_2758 & x_2770);
	assign x_2745 = (x_2732 & x_2744);
	assign x_2720 = (x_2707 & x_2719);
	assign x_2695 = (x_2682 & x_2694);
	assign x_2670 = (x_2657 & x_2669);
	assign x_2643 = (x_2630 & x_2642);
	assign x_2618 = (x_2605 & x_2617);
	assign x_2593 = (x_2580 & x_2592);
	assign x_2568 = (x_2555 & x_2567);
	assign x_2542 = (x_2529 & x_2541);
	assign x_2517 = (x_2504 & x_2516);
	assign x_2492 = (x_2479 & x_2491);
	assign x_2468 = (x_2455 & x_2467);
	assign x_2439 = (x_2426 & x_2438);
	assign x_2414 = (x_2401 & x_2413);
	assign x_2389 = (x_2376 & x_2388);
	assign x_2364 = (x_2351 & x_2363);
	assign x_2338 = (x_2325 & x_2337);
	assign x_2313 = (x_2300 & x_2312);
	assign x_2288 = (x_2275 & x_2287);
	assign x_2263 = (x_2250 & x_2262);
	assign x_2236 = (x_2223 & x_2235);
	assign x_2211 = (x_2198 & x_2210);
	assign x_2186 = (x_2173 & x_2185);
	assign x_2161 = (x_2148 & x_2160);
	assign x_2135 = (x_2122 & x_2134);
	assign x_2110 = (x_2097 & x_2109);
	assign x_2085 = (x_2072 & x_2084);
	assign x_2060 = (x_2047 & x_2059);
	assign x_2032 = (x_2019 & x_2031);
	assign x_2007 = (x_1994 & x_2006);
	assign x_1982 = (x_1969 & x_1981);
	assign x_1957 = (x_1944 & x_1956);
	assign x_1931 = (x_1918 & x_1930);
	assign x_1906 = (x_1893 & x_1905);
	assign x_1881 = (x_1868 & x_1880);
	assign x_1856 = (x_1843 & x_1855);
	assign x_1829 = (x_1816 & x_1828);
	assign x_1804 = (x_1791 & x_1803);
	assign x_1779 = (x_1766 & x_1778);
	assign x_1754 = (x_1741 & x_1753);
	assign x_1728 = (x_1715 & x_1727);
	assign x_1703 = (x_1690 & x_1702);
	assign x_1678 = (x_1665 & x_1677);
	assign x_1654 = (x_1641 & x_1653);
	assign x_3254 = (x_3228 & x_3253);
	assign x_3204 = (x_3178 & x_3203);
	assign x_3153 = (x_3127 & x_3152);
	assign x_3103 = (x_3077 & x_3102);
	assign x_3051 = (x_3025 & x_3050);
	assign x_3001 = (x_2975 & x_3000);
	assign x_2950 = (x_2924 & x_2949);
	assign x_2900 = (x_2874 & x_2899);
	assign x_2847 = (x_2821 & x_2846);
	assign x_2797 = (x_2771 & x_2796);
	assign x_2746 = (x_2720 & x_2745);
	assign x_2696 = (x_2670 & x_2695);
	assign x_2644 = (x_2618 & x_2643);
	assign x_2594 = (x_2568 & x_2593);
	assign x_2543 = (x_2517 & x_2542);
	assign x_2493 = (x_2468 & x_2492);
	assign x_2440 = (x_2414 & x_2439);
	assign x_2390 = (x_2364 & x_2389);
	assign x_2339 = (x_2313 & x_2338);
	assign x_2289 = (x_2263 & x_2288);
	assign x_2237 = (x_2211 & x_2236);
	assign x_2187 = (x_2161 & x_2186);
	assign x_2136 = (x_2110 & x_2135);
	assign x_2086 = (x_2060 & x_2085);
	assign x_2033 = (x_2007 & x_2032);
	assign x_1983 = (x_1957 & x_1982);
	assign x_1932 = (x_1906 & x_1931);
	assign x_1882 = (x_1856 & x_1881);
	assign x_1830 = (x_1804 & x_1829);
	assign x_1780 = (x_1754 & x_1779);
	assign x_1729 = (x_1703 & x_1728);
	assign x_1679 = (x_1654 & x_1678);
	assign x_3255 = (x_3204 & x_3254);
	assign x_3154 = (x_3103 & x_3153);
	assign x_3052 = (x_3001 & x_3051);
	assign x_2951 = (x_2900 & x_2950);
	assign x_2848 = (x_2797 & x_2847);
	assign x_2747 = (x_2696 & x_2746);
	assign x_2645 = (x_2594 & x_2644);
	assign x_2544 = (x_2493 & x_2543);
	assign x_2441 = (x_2390 & x_2440);
	assign x_2340 = (x_2289 & x_2339);
	assign x_2238 = (x_2187 & x_2237);
	assign x_2137 = (x_2086 & x_2136);
	assign x_2034 = (x_1983 & x_2033);
	assign x_1933 = (x_1882 & x_1932);
	assign x_1831 = (x_1780 & x_1830);
	assign x_1730 = (x_1679 & x_1729);
	assign x_3256 = (x_3154 & x_3255);
	assign x_3053 = (x_2951 & x_3052);
	assign x_2849 = (x_2747 & x_2848);
	assign x_2646 = (x_2544 & x_2645);
	assign x_2442 = (x_2340 & x_2441);
	assign x_2239 = (x_2137 & x_2238);
	assign x_2035 = (x_1933 & x_2034);
	assign x_1832 = (x_1730 & x_1831);
	assign x_3257 = (x_3053 & x_3256);
	assign x_2850 = (x_2646 & x_2849);
	assign x_2443 = (x_2239 & x_2442);
	assign x_2036 = (x_1832 & x_2035);
	assign x_3258 = (x_2850 & x_3257);
	assign x_2444 = (x_2036 & x_2443);
	assign x_3259 = (x_2444 & x_3258);
	assign o_1 = x_325);
endmodule
