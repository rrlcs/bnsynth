// Benchmark "SKOLEMFORMULA" written by ABC on Fri May 20 19:42:52 2022

module SKOLEMFORMULA ( 
    i0,
    i1  );
  input  i0;
  output i1;
  assign i1 = 1'b1;
endmodule


