// Benchmark "SKOLEMFORMULA" written by ABC on Wed May 18 00:57:13 2022

module SKOLEMFORMULA ( 
    i0,
    i1  );
  input  i0;
  output i1;
  assign i1 = 1'b1;
endmodule


