module add20ysat(v_14,v_9,v_40,v_67,v_94,v_121,v_148,v_175,v_202,v_229,v_256,v_283,v_310,v_337,v_364,v_391,v_418,v_445,v_472,v_510,v_13,v_8,v_39,v_66,v_93,v_120,v_147,v_174,v_201,v_228,v_255,v_282,v_309,v_336,v_363,v_390,v_417,v_444,v_471,v_502,v_607,v_1,v_3,v_32,v_23,v_58,v_85,v_112,v_139,v_166,v_193,v_220,v_247,v_274,v_301,v_328,v_355,v_382,v_409,v_436,v_463,v_490,v_517,v_6,v_7,v_606,o_1);
	input v_14;
	input v_9;
	input v_40;
	input v_67;
	input v_94;
	input v_121;
	input v_148;
	input v_175;
	input v_202;
	input v_229;
	input v_256;
	input v_283;
	input v_310;
	input v_337;
	input v_364;
	input v_391;
	input v_418;
	input v_445;
	input v_472;
	input v_510;
	input v_13;
	input v_8;
	input v_39;
	input v_66;
	input v_93;
	input v_120;
	input v_147;
	input v_174;
	input v_201;
	input v_228;
	input v_255;
	input v_282;
	input v_309;
	input v_336;
	input v_363;
	input v_390;
	input v_417;
	input v_444;
	input v_471;
	input v_502;
	input v_607;
	input v_1;
	input v_3;
	input v_32;
	input v_23;
	input v_58;
	input v_85;
	input v_112;
	input v_139;
	input v_166;
	input v_193;
	input v_220;
	input v_247;
	input v_274;
	input v_301;
	input v_328;
	input v_355;
	input v_382;
	input v_409;
	input v_436;
	input v_463;
	input v_490;
	input v_517;
	input v_6;
	input v_7;
	input v_606;
	wire v_2;
	wire v_4;
	wire v_5;
	wire v_10;
	wire v_11;
	wire v_12;
	wire v_15;
	wire v_16;
	wire v_17;
	wire v_18;
	wire v_19;
	wire v_20;
	wire v_21;
	wire v_22;
	wire v_24;
	wire v_25;
	wire v_26;
	wire v_27;
	wire v_28;
	wire v_29;
	wire v_30;
	wire v_31;
	wire v_33;
	wire v_34;
	wire v_35;
	wire v_36;
	wire v_37;
	wire v_38;
	wire v_41;
	wire v_42;
	wire v_43;
	wire v_44;
	wire v_45;
	wire v_46;
	wire v_47;
	wire v_48;
	wire v_49;
	wire v_50;
	wire v_51;
	wire v_52;
	wire v_53;
	wire v_54;
	wire v_55;
	wire v_56;
	wire v_57;
	wire v_59;
	wire v_60;
	wire v_61;
	wire v_62;
	wire v_63;
	wire v_64;
	wire v_65;
	wire v_68;
	wire v_69;
	wire v_70;
	wire v_71;
	wire v_72;
	wire v_73;
	wire v_74;
	wire v_75;
	wire v_76;
	wire v_77;
	wire v_78;
	wire v_79;
	wire v_80;
	wire v_81;
	wire v_82;
	wire v_83;
	wire v_84;
	wire v_86;
	wire v_87;
	wire v_88;
	wire v_89;
	wire v_90;
	wire v_91;
	wire v_92;
	wire v_95;
	wire v_96;
	wire v_97;
	wire v_98;
	wire v_99;
	wire v_100;
	wire v_101;
	wire v_102;
	wire v_103;
	wire v_104;
	wire v_105;
	wire v_106;
	wire v_107;
	wire v_108;
	wire v_109;
	wire v_110;
	wire v_111;
	wire v_113;
	wire v_114;
	wire v_115;
	wire v_116;
	wire v_117;
	wire v_118;
	wire v_119;
	wire v_122;
	wire v_123;
	wire v_124;
	wire v_125;
	wire v_126;
	wire v_127;
	wire v_128;
	wire v_129;
	wire v_130;
	wire v_131;
	wire v_132;
	wire v_133;
	wire v_134;
	wire v_135;
	wire v_136;
	wire v_137;
	wire v_138;
	wire v_140;
	wire v_141;
	wire v_142;
	wire v_143;
	wire v_144;
	wire v_145;
	wire v_146;
	wire v_149;
	wire v_150;
	wire v_151;
	wire v_152;
	wire v_153;
	wire v_154;
	wire v_155;
	wire v_156;
	wire v_157;
	wire v_158;
	wire v_159;
	wire v_160;
	wire v_161;
	wire v_162;
	wire v_163;
	wire v_164;
	wire v_165;
	wire v_167;
	wire v_168;
	wire v_169;
	wire v_170;
	wire v_171;
	wire v_172;
	wire v_173;
	wire v_176;
	wire v_177;
	wire v_178;
	wire v_179;
	wire v_180;
	wire v_181;
	wire v_182;
	wire v_183;
	wire v_184;
	wire v_185;
	wire v_186;
	wire v_187;
	wire v_188;
	wire v_189;
	wire v_190;
	wire v_191;
	wire v_192;
	wire v_194;
	wire v_195;
	wire v_196;
	wire v_197;
	wire v_198;
	wire v_199;
	wire v_200;
	wire v_203;
	wire v_204;
	wire v_205;
	wire v_206;
	wire v_207;
	wire v_208;
	wire v_209;
	wire v_210;
	wire v_211;
	wire v_212;
	wire v_213;
	wire v_214;
	wire v_215;
	wire v_216;
	wire v_217;
	wire v_218;
	wire v_219;
	wire v_221;
	wire v_222;
	wire v_223;
	wire v_224;
	wire v_225;
	wire v_226;
	wire v_227;
	wire v_230;
	wire v_231;
	wire v_232;
	wire v_233;
	wire v_234;
	wire v_235;
	wire v_236;
	wire v_237;
	wire v_238;
	wire v_239;
	wire v_240;
	wire v_241;
	wire v_242;
	wire v_243;
	wire v_244;
	wire v_245;
	wire v_246;
	wire v_248;
	wire v_249;
	wire v_250;
	wire v_251;
	wire v_252;
	wire v_253;
	wire v_254;
	wire v_257;
	wire v_258;
	wire v_259;
	wire v_260;
	wire v_261;
	wire v_262;
	wire v_263;
	wire v_264;
	wire v_265;
	wire v_266;
	wire v_267;
	wire v_268;
	wire v_269;
	wire v_270;
	wire v_271;
	wire v_272;
	wire v_273;
	wire v_275;
	wire v_276;
	wire v_277;
	wire v_278;
	wire v_279;
	wire v_280;
	wire v_281;
	wire v_284;
	wire v_285;
	wire v_286;
	wire v_287;
	wire v_288;
	wire v_289;
	wire v_290;
	wire v_291;
	wire v_292;
	wire v_293;
	wire v_294;
	wire v_295;
	wire v_296;
	wire v_297;
	wire v_298;
	wire v_299;
	wire v_300;
	wire v_302;
	wire v_303;
	wire v_304;
	wire v_305;
	wire v_306;
	wire v_307;
	wire v_308;
	wire v_311;
	wire v_312;
	wire v_313;
	wire v_314;
	wire v_315;
	wire v_316;
	wire v_317;
	wire v_318;
	wire v_319;
	wire v_320;
	wire v_321;
	wire v_322;
	wire v_323;
	wire v_324;
	wire v_325;
	wire v_326;
	wire v_327;
	wire v_329;
	wire v_330;
	wire v_331;
	wire v_332;
	wire v_333;
	wire v_334;
	wire v_335;
	wire v_338;
	wire v_339;
	wire v_340;
	wire v_341;
	wire v_342;
	wire v_343;
	wire v_344;
	wire v_345;
	wire v_346;
	wire v_347;
	wire v_348;
	wire v_349;
	wire v_350;
	wire v_351;
	wire v_352;
	wire v_353;
	wire v_354;
	wire v_356;
	wire v_357;
	wire v_358;
	wire v_359;
	wire v_360;
	wire v_361;
	wire v_362;
	wire v_365;
	wire v_366;
	wire v_367;
	wire v_368;
	wire v_369;
	wire v_370;
	wire v_371;
	wire v_372;
	wire v_373;
	wire v_374;
	wire v_375;
	wire v_376;
	wire v_377;
	wire v_378;
	wire v_379;
	wire v_380;
	wire v_381;
	wire v_383;
	wire v_384;
	wire v_385;
	wire v_386;
	wire v_387;
	wire v_388;
	wire v_389;
	wire v_392;
	wire v_393;
	wire v_394;
	wire v_395;
	wire v_396;
	wire v_397;
	wire v_398;
	wire v_399;
	wire v_400;
	wire v_401;
	wire v_402;
	wire v_403;
	wire v_404;
	wire v_405;
	wire v_406;
	wire v_407;
	wire v_408;
	wire v_410;
	wire v_411;
	wire v_412;
	wire v_413;
	wire v_414;
	wire v_415;
	wire v_416;
	wire v_419;
	wire v_420;
	wire v_421;
	wire v_422;
	wire v_423;
	wire v_424;
	wire v_425;
	wire v_426;
	wire v_427;
	wire v_428;
	wire v_429;
	wire v_430;
	wire v_431;
	wire v_432;
	wire v_433;
	wire v_434;
	wire v_435;
	wire v_437;
	wire v_438;
	wire v_439;
	wire v_440;
	wire v_441;
	wire v_442;
	wire v_443;
	wire v_446;
	wire v_447;
	wire v_448;
	wire v_449;
	wire v_450;
	wire v_451;
	wire v_452;
	wire v_453;
	wire v_454;
	wire v_455;
	wire v_456;
	wire v_457;
	wire v_458;
	wire v_459;
	wire v_460;
	wire v_461;
	wire v_462;
	wire v_464;
	wire v_465;
	wire v_466;
	wire v_467;
	wire v_468;
	wire v_469;
	wire v_470;
	wire v_473;
	wire v_474;
	wire v_475;
	wire v_476;
	wire v_477;
	wire v_478;
	wire v_479;
	wire v_480;
	wire v_481;
	wire v_482;
	wire v_483;
	wire v_484;
	wire v_485;
	wire v_486;
	wire v_487;
	wire v_488;
	wire v_489;
	wire v_491;
	wire v_492;
	wire v_493;
	wire v_494;
	wire v_495;
	wire v_496;
	wire v_497;
	wire v_498;
	wire v_499;
	wire v_500;
	wire v_501;
	wire v_503;
	wire v_504;
	wire v_505;
	wire v_506;
	wire v_507;
	wire v_508;
	wire v_509;
	wire v_511;
	wire v_512;
	wire v_513;
	wire v_514;
	wire v_515;
	wire v_516;
	wire v_518;
	wire v_519;
	wire v_520;
	wire v_521;
	wire v_522;
	wire v_523;
	wire v_524;
	wire v_525;
	wire v_526;
	wire v_527;
	wire v_528;
	wire v_529;
	wire v_530;
	wire v_531;
	wire v_532;
	wire v_533;
	wire v_534;
	wire v_535;
	wire v_536;
	wire v_537;
	wire v_538;
	wire v_539;
	wire v_540;
	wire v_541;
	wire v_542;
	wire v_543;
	wire v_544;
	wire v_545;
	wire v_546;
	wire v_547;
	wire v_548;
	wire v_549;
	wire v_550;
	wire v_551;
	wire v_552;
	wire v_553;
	wire v_554;
	wire v_555;
	wire v_556;
	wire v_557;
	wire v_558;
	wire v_559;
	wire v_560;
	wire v_561;
	wire v_562;
	wire v_563;
	wire v_564;
	wire v_565;
	wire v_566;
	wire v_567;
	wire v_568;
	wire v_569;
	wire v_570;
	wire v_571;
	wire v_572;
	wire v_573;
	wire v_574;
	wire v_575;
	wire v_576;
	wire v_577;
	wire v_578;
	wire v_579;
	wire v_580;
	wire v_581;
	wire v_582;
	wire v_583;
	wire v_584;
	wire v_585;
	wire v_586;
	wire v_587;
	wire v_588;
	wire v_589;
	wire v_590;
	wire v_591;
	wire v_592;
	wire v_593;
	wire v_594;
	wire v_595;
	wire v_596;
	wire v_597;
	wire v_598;
	wire v_599;
	wire v_600;
	wire v_601;
	wire v_602;
	wire v_603;
	wire v_604;
	wire v_605;
	wire v_608;
	wire v_609;
	wire v_610;
	wire v_611;
	wire v_612;
	wire v_613;
	wire v_614;
	wire v_615;
	wire v_616;
	wire v_617;
	wire v_618;
	wire x_1;
	output o_1;
	assign v_15 = (v_13 & v_14);
	assign v_30 = (~v_13 & ~v_14);
	assign v_20 = (~v_13 | ~v_14);
	assign v_34 = (v_13 | v_14);
	assign v_17 = (~v_8 & v_9);
	assign v_18 = (v_8 & ~v_9);
	assign v_44 = (~v_8 & ~v_9);
	assign v_54 = (v_8 & v_9);
	assign v_10 = (v_8 | ~v_9);
	assign v_11 = (~v_8 | v_9);
	assign v_46 = (~v_8 | ~v_9);
	assign v_52 = (v_8 | v_9);
	assign v_49 = (~v_39 & v_40);
	assign v_50 = (v_39 & ~v_40);
	assign v_71 = (~v_39 & ~v_40);
	assign v_81 = (v_39 & v_40);
	assign v_41 = (v_39 | ~v_40);
	assign v_42 = (~v_39 | v_40);
	assign v_73 = (~v_39 | ~v_40);
	assign v_79 = (v_39 | v_40);
	assign v_76 = (~v_66 & v_67);
	assign v_77 = (v_66 & ~v_67);
	assign v_98 = (~v_66 & ~v_67);
	assign v_108 = (v_66 & v_67);
	assign v_68 = (v_66 | ~v_67);
	assign v_69 = (~v_66 | v_67);
	assign v_100 = (~v_66 | ~v_67);
	assign v_106 = (v_66 | v_67);
	assign v_103 = (~v_93 & v_94);
	assign v_104 = (v_93 & ~v_94);
	assign v_125 = (~v_93 & ~v_94);
	assign v_135 = (v_93 & v_94);
	assign v_95 = (v_93 | ~v_94);
	assign v_96 = (~v_93 | v_94);
	assign v_127 = (~v_93 | ~v_94);
	assign v_133 = (v_93 | v_94);
	assign v_130 = (~v_120 & v_121);
	assign v_131 = (v_120 & ~v_121);
	assign v_152 = (~v_120 & ~v_121);
	assign v_162 = (v_120 & v_121);
	assign v_122 = (v_120 | ~v_121);
	assign v_123 = (~v_120 | v_121);
	assign v_154 = (~v_120 | ~v_121);
	assign v_160 = (v_120 | v_121);
	assign v_157 = (~v_147 & v_148);
	assign v_158 = (v_147 & ~v_148);
	assign v_179 = (~v_147 & ~v_148);
	assign v_189 = (v_147 & v_148);
	assign v_149 = (v_147 | ~v_148);
	assign v_150 = (~v_147 | v_148);
	assign v_181 = (~v_147 | ~v_148);
	assign v_187 = (v_147 | v_148);
	assign v_184 = (~v_174 & v_175);
	assign v_185 = (v_174 & ~v_175);
	assign v_206 = (~v_174 & ~v_175);
	assign v_216 = (v_174 & v_175);
	assign v_176 = (v_174 | ~v_175);
	assign v_177 = (~v_174 | v_175);
	assign v_208 = (~v_174 | ~v_175);
	assign v_214 = (v_174 | v_175);
	assign v_211 = (~v_201 & v_202);
	assign v_212 = (v_201 & ~v_202);
	assign v_233 = (~v_201 & ~v_202);
	assign v_243 = (v_201 & v_202);
	assign v_203 = (v_201 | ~v_202);
	assign v_204 = (~v_201 | v_202);
	assign v_235 = (~v_201 | ~v_202);
	assign v_241 = (v_201 | v_202);
	assign v_238 = (~v_228 & v_229);
	assign v_239 = (v_228 & ~v_229);
	assign v_260 = (~v_228 & ~v_229);
	assign v_270 = (v_228 & v_229);
	assign v_230 = (v_228 | ~v_229);
	assign v_231 = (~v_228 | v_229);
	assign v_262 = (~v_228 | ~v_229);
	assign v_268 = (v_228 | v_229);
	assign v_265 = (~v_255 & v_256);
	assign v_266 = (v_255 & ~v_256);
	assign v_287 = (~v_255 & ~v_256);
	assign v_297 = (v_255 & v_256);
	assign v_257 = (v_255 | ~v_256);
	assign v_258 = (~v_255 | v_256);
	assign v_289 = (~v_255 | ~v_256);
	assign v_295 = (v_255 | v_256);
	assign v_292 = (~v_282 & v_283);
	assign v_293 = (v_282 & ~v_283);
	assign v_314 = (~v_282 & ~v_283);
	assign v_324 = (v_282 & v_283);
	assign v_284 = (v_282 | ~v_283);
	assign v_285 = (~v_282 | v_283);
	assign v_316 = (~v_282 | ~v_283);
	assign v_322 = (v_282 | v_283);
	assign v_319 = (~v_309 & v_310);
	assign v_320 = (v_309 & ~v_310);
	assign v_341 = (~v_309 & ~v_310);
	assign v_351 = (v_309 & v_310);
	assign v_311 = (v_309 | ~v_310);
	assign v_312 = (~v_309 | v_310);
	assign v_343 = (~v_309 | ~v_310);
	assign v_349 = (v_309 | v_310);
	assign v_346 = (~v_336 & v_337);
	assign v_347 = (v_336 & ~v_337);
	assign v_368 = (~v_336 & ~v_337);
	assign v_378 = (v_336 & v_337);
	assign v_338 = (v_336 | ~v_337);
	assign v_339 = (~v_336 | v_337);
	assign v_370 = (~v_336 | ~v_337);
	assign v_376 = (v_336 | v_337);
	assign v_373 = (~v_363 & v_364);
	assign v_374 = (v_363 & ~v_364);
	assign v_395 = (~v_363 & ~v_364);
	assign v_405 = (v_363 & v_364);
	assign v_365 = (v_363 | ~v_364);
	assign v_366 = (~v_363 | v_364);
	assign v_397 = (~v_363 | ~v_364);
	assign v_403 = (v_363 | v_364);
	assign v_400 = (~v_390 & v_391);
	assign v_401 = (v_390 & ~v_391);
	assign v_422 = (~v_390 & ~v_391);
	assign v_432 = (v_390 & v_391);
	assign v_392 = (v_390 | ~v_391);
	assign v_393 = (~v_390 | v_391);
	assign v_424 = (~v_390 | ~v_391);
	assign v_430 = (v_390 | v_391);
	assign v_427 = (~v_417 & v_418);
	assign v_428 = (v_417 & ~v_418);
	assign v_449 = (~v_417 & ~v_418);
	assign v_459 = (v_417 & v_418);
	assign v_419 = (v_417 | ~v_418);
	assign v_420 = (~v_417 | v_418);
	assign v_451 = (~v_417 | ~v_418);
	assign v_457 = (v_417 | v_418);
	assign v_454 = (~v_444 & v_445);
	assign v_455 = (v_444 & ~v_445);
	assign v_476 = (~v_444 & ~v_445);
	assign v_486 = (v_444 & v_445);
	assign v_446 = (v_444 | ~v_445);
	assign v_447 = (~v_444 | v_445);
	assign v_478 = (~v_444 | ~v_445);
	assign v_484 = (v_444 | v_445);
	assign v_481 = (~v_471 & v_472);
	assign v_482 = (v_471 & ~v_472);
	assign v_500 = (v_471 & v_472);
	assign v_504 = (~v_471 & ~v_472);
	assign v_473 = (v_471 | ~v_472);
	assign v_474 = (~v_471 | v_472);
	assign v_498 = (v_471 | v_472);
	assign v_506 = (~v_471 | ~v_472);
	assign v_2 = v_1;
	assign v_608 = (v_1 & v_607);
	assign v_610 = (~v_1 | ~v_607);
	assign v_4 = v_3;
	assign v_612 = ~v_7;
	assign v_613 = ~v_606;
	assign v_31 = (v_15 | v_30);
	assign v_35 = (v_20 & v_34);
	assign v_19 = (v_17 | v_18);
	assign v_45 = (v_20 | v_44);
	assign v_12 = (v_10 & v_11);
	assign v_53 = (v_15 & v_52);
	assign v_51 = (v_49 | v_50);
	assign v_43 = (v_41 & v_42);
	assign v_78 = (v_76 | v_77);
	assign v_70 = (v_68 & v_69);
	assign v_105 = (v_103 | v_104);
	assign v_97 = (v_95 & v_96);
	assign v_132 = (v_130 | v_131);
	assign v_124 = (v_122 & v_123);
	assign v_159 = (v_157 | v_158);
	assign v_151 = (v_149 & v_150);
	assign v_186 = (v_184 | v_185);
	assign v_178 = (v_176 & v_177);
	assign v_213 = (v_211 | v_212);
	assign v_205 = (v_203 & v_204);
	assign v_240 = (v_238 | v_239);
	assign v_232 = (v_230 & v_231);
	assign v_267 = (v_265 | v_266);
	assign v_259 = (v_257 & v_258);
	assign v_294 = (v_292 | v_293);
	assign v_286 = (v_284 & v_285);
	assign v_321 = (v_319 | v_320);
	assign v_313 = (v_311 & v_312);
	assign v_348 = (v_346 | v_347);
	assign v_340 = (v_338 & v_339);
	assign v_375 = (v_373 | v_374);
	assign v_367 = (v_365 & v_366);
	assign v_402 = (v_400 | v_401);
	assign v_394 = (v_392 & v_393);
	assign v_429 = (v_427 | v_428);
	assign v_421 = (v_419 & v_420);
	assign v_456 = (v_454 | v_455);
	assign v_448 = (v_446 & v_447);
	assign v_483 = (v_481 | v_482);
	assign v_475 = (v_473 & v_474);
	assign v_609 = (~v_606 | v_608);
	assign v_611 = (v_606 | v_610);
	assign v_5 = (v_2 | v_4);
	assign v_614 = (v_612 & v_613);
	assign v_33 = (v_31 & v_32);
	assign v_530 = (v_31 | v_32);
	assign v_36 = (~v_32 & v_35);
	assign v_529 = (~v_32 | v_35);
	assign v_25 = (v_19 & v_20);
	assign v_21 = (v_19 | v_20);
	assign v_47 = (v_45 & v_46);
	assign v_26 = (v_12 & v_15);
	assign v_16 = (v_12 | v_15);
	assign v_55 = (v_53 | v_54);
	assign v_618 = v_614;
	assign v_37 = (v_33 | v_36);
	assign v_531 = (v_529 & v_530);
	assign v_48 = (v_43 & v_47);
	assign v_61 = (v_43 | v_47);
	assign v_72 = (v_47 | v_71);
	assign v_27 = (v_25 | v_26);
	assign v_22 = (v_16 & v_21);
	assign v_56 = (v_51 & v_55);
	assign v_80 = (v_55 & v_79);
	assign v_60 = (v_51 | v_55);
	assign v_74 = (v_72 & v_73);
	assign v_28 = (~v_23 & v_27);
	assign v_526 = (~v_23 | v_27);
	assign v_24 = (v_22 & v_23);
	assign v_527 = (v_22 | v_23);
	assign v_57 = (v_48 | v_56);
	assign v_82 = (v_80 | v_81);
	assign v_62 = (v_60 & v_61);
	assign v_75 = (v_70 & v_74);
	assign v_88 = (v_70 | v_74);
	assign v_99 = (v_74 | v_98);
	assign v_29 = (v_24 | v_28);
	assign v_528 = (v_526 & v_527);
	assign v_59 = (v_57 & v_58);
	assign v_534 = (v_57 | v_58);
	assign v_83 = (v_78 & v_82);
	assign v_107 = (v_82 & v_106);
	assign v_87 = (v_78 | v_82);
	assign v_63 = (~v_58 & v_62);
	assign v_533 = (~v_58 | v_62);
	assign v_101 = (v_99 & v_100);
	assign v_38 = (v_29 | v_37);
	assign v_532 = (v_528 & v_531);
	assign v_84 = (v_75 | v_83);
	assign v_109 = (v_107 | v_108);
	assign v_89 = (v_87 & v_88);
	assign v_64 = (v_59 | v_63);
	assign v_535 = (v_533 & v_534);
	assign v_102 = (v_97 & v_101);
	assign v_115 = (v_97 | v_101);
	assign v_126 = (v_101 | v_125);
	assign v_86 = (v_84 & v_85);
	assign v_538 = (v_84 | v_85);
	assign v_110 = (v_105 & v_109);
	assign v_134 = (v_109 & v_133);
	assign v_114 = (v_105 | v_109);
	assign v_90 = (~v_85 & v_89);
	assign v_537 = (~v_85 | v_89);
	assign v_65 = (v_38 | v_64);
	assign v_536 = (v_532 & v_535);
	assign v_128 = (v_126 & v_127);
	assign v_111 = (v_102 | v_110);
	assign v_136 = (v_134 | v_135);
	assign v_116 = (v_114 & v_115);
	assign v_91 = (v_86 | v_90);
	assign v_539 = (v_537 & v_538);
	assign v_129 = (v_124 & v_128);
	assign v_142 = (v_124 | v_128);
	assign v_153 = (v_128 | v_152);
	assign v_113 = (v_111 & v_112);
	assign v_542 = (v_111 | v_112);
	assign v_137 = (v_132 & v_136);
	assign v_161 = (v_136 & v_160);
	assign v_141 = (v_132 | v_136);
	assign v_117 = (~v_112 & v_116);
	assign v_541 = (~v_112 | v_116);
	assign v_92 = (v_65 | v_91);
	assign v_540 = (v_536 & v_539);
	assign v_155 = (v_153 & v_154);
	assign v_138 = (v_129 | v_137);
	assign v_163 = (v_161 | v_162);
	assign v_143 = (v_141 & v_142);
	assign v_118 = (v_113 | v_117);
	assign v_543 = (v_541 & v_542);
	assign v_156 = (v_151 & v_155);
	assign v_169 = (v_151 | v_155);
	assign v_180 = (v_155 | v_179);
	assign v_140 = (v_138 & v_139);
	assign v_546 = (v_138 | v_139);
	assign v_164 = (v_159 & v_163);
	assign v_188 = (v_163 & v_187);
	assign v_168 = (v_159 | v_163);
	assign v_144 = (~v_139 & v_143);
	assign v_545 = (~v_139 | v_143);
	assign v_119 = (v_92 | v_118);
	assign v_544 = (v_540 & v_543);
	assign v_182 = (v_180 & v_181);
	assign v_165 = (v_156 | v_164);
	assign v_190 = (v_188 | v_189);
	assign v_170 = (v_168 & v_169);
	assign v_145 = (v_140 | v_144);
	assign v_547 = (v_545 & v_546);
	assign v_183 = (v_178 & v_182);
	assign v_196 = (v_178 | v_182);
	assign v_207 = (v_182 | v_206);
	assign v_167 = (v_165 & v_166);
	assign v_550 = (v_165 | v_166);
	assign v_191 = (v_186 & v_190);
	assign v_215 = (v_190 & v_214);
	assign v_195 = (v_186 | v_190);
	assign v_171 = (~v_166 & v_170);
	assign v_549 = (~v_166 | v_170);
	assign v_146 = (v_119 | v_145);
	assign v_548 = (v_544 & v_547);
	assign v_209 = (v_207 & v_208);
	assign v_192 = (v_183 | v_191);
	assign v_217 = (v_215 | v_216);
	assign v_197 = (v_195 & v_196);
	assign v_172 = (v_167 | v_171);
	assign v_551 = (v_549 & v_550);
	assign v_210 = (v_205 & v_209);
	assign v_223 = (v_205 | v_209);
	assign v_234 = (v_209 | v_233);
	assign v_194 = (v_192 & v_193);
	assign v_554 = (v_192 | v_193);
	assign v_218 = (v_213 & v_217);
	assign v_242 = (v_217 & v_241);
	assign v_222 = (v_213 | v_217);
	assign v_198 = (~v_193 & v_197);
	assign v_553 = (~v_193 | v_197);
	assign v_173 = (v_146 | v_172);
	assign v_552 = (v_548 & v_551);
	assign v_236 = (v_234 & v_235);
	assign v_219 = (v_210 | v_218);
	assign v_244 = (v_242 | v_243);
	assign v_224 = (v_222 & v_223);
	assign v_199 = (v_194 | v_198);
	assign v_555 = (v_553 & v_554);
	assign v_237 = (v_232 & v_236);
	assign v_250 = (v_232 | v_236);
	assign v_261 = (v_236 | v_260);
	assign v_221 = (v_219 & v_220);
	assign v_558 = (v_219 | v_220);
	assign v_245 = (v_240 & v_244);
	assign v_269 = (v_244 & v_268);
	assign v_249 = (v_240 | v_244);
	assign v_225 = (~v_220 & v_224);
	assign v_557 = (~v_220 | v_224);
	assign v_200 = (v_173 | v_199);
	assign v_556 = (v_552 & v_555);
	assign v_263 = (v_261 & v_262);
	assign v_246 = (v_237 | v_245);
	assign v_271 = (v_269 | v_270);
	assign v_251 = (v_249 & v_250);
	assign v_226 = (v_221 | v_225);
	assign v_559 = (v_557 & v_558);
	assign v_264 = (v_259 & v_263);
	assign v_277 = (v_259 | v_263);
	assign v_288 = (v_263 | v_287);
	assign v_248 = (v_246 & v_247);
	assign v_562 = (v_246 | v_247);
	assign v_272 = (v_267 & v_271);
	assign v_296 = (v_271 & v_295);
	assign v_276 = (v_267 | v_271);
	assign v_252 = (~v_247 & v_251);
	assign v_561 = (~v_247 | v_251);
	assign v_227 = (v_200 | v_226);
	assign v_560 = (v_556 & v_559);
	assign v_290 = (v_288 & v_289);
	assign v_273 = (v_264 | v_272);
	assign v_298 = (v_296 | v_297);
	assign v_278 = (v_276 & v_277);
	assign v_253 = (v_248 | v_252);
	assign v_563 = (v_561 & v_562);
	assign v_291 = (v_286 & v_290);
	assign v_304 = (v_286 | v_290);
	assign v_315 = (v_290 | v_314);
	assign v_275 = (v_273 & v_274);
	assign v_566 = (v_273 | v_274);
	assign v_299 = (v_294 & v_298);
	assign v_323 = (v_298 & v_322);
	assign v_303 = (v_294 | v_298);
	assign v_279 = (~v_274 & v_278);
	assign v_565 = (~v_274 | v_278);
	assign v_254 = (v_227 | v_253);
	assign v_564 = (v_560 & v_563);
	assign v_317 = (v_315 & v_316);
	assign v_300 = (v_291 | v_299);
	assign v_325 = (v_323 | v_324);
	assign v_305 = (v_303 & v_304);
	assign v_280 = (v_275 | v_279);
	assign v_567 = (v_565 & v_566);
	assign v_318 = (v_313 & v_317);
	assign v_331 = (v_313 | v_317);
	assign v_342 = (v_317 | v_341);
	assign v_302 = (v_300 & v_301);
	assign v_570 = (v_300 | v_301);
	assign v_326 = (v_321 & v_325);
	assign v_350 = (v_325 & v_349);
	assign v_330 = (v_321 | v_325);
	assign v_306 = (~v_301 & v_305);
	assign v_569 = (~v_301 | v_305);
	assign v_281 = (v_254 | v_280);
	assign v_568 = (v_564 & v_567);
	assign v_344 = (v_342 & v_343);
	assign v_327 = (v_318 | v_326);
	assign v_352 = (v_350 | v_351);
	assign v_332 = (v_330 & v_331);
	assign v_307 = (v_302 | v_306);
	assign v_571 = (v_569 & v_570);
	assign v_345 = (v_340 & v_344);
	assign v_358 = (v_340 | v_344);
	assign v_369 = (v_344 | v_368);
	assign v_329 = (v_327 & v_328);
	assign v_574 = (v_327 | v_328);
	assign v_353 = (v_348 & v_352);
	assign v_377 = (v_352 & v_376);
	assign v_357 = (v_348 | v_352);
	assign v_333 = (~v_328 & v_332);
	assign v_573 = (~v_328 | v_332);
	assign v_308 = (v_281 | v_307);
	assign v_572 = (v_568 & v_571);
	assign v_371 = (v_369 & v_370);
	assign v_354 = (v_345 | v_353);
	assign v_379 = (v_377 | v_378);
	assign v_359 = (v_357 & v_358);
	assign v_334 = (v_329 | v_333);
	assign v_575 = (v_573 & v_574);
	assign v_372 = (v_367 & v_371);
	assign v_385 = (v_367 | v_371);
	assign v_396 = (v_371 | v_395);
	assign v_356 = (v_354 & v_355);
	assign v_578 = (v_354 | v_355);
	assign v_380 = (v_375 & v_379);
	assign v_404 = (v_379 & v_403);
	assign v_384 = (v_375 | v_379);
	assign v_360 = (~v_355 & v_359);
	assign v_577 = (~v_355 | v_359);
	assign v_335 = (v_308 | v_334);
	assign v_576 = (v_572 & v_575);
	assign v_398 = (v_396 & v_397);
	assign v_381 = (v_372 | v_380);
	assign v_406 = (v_404 | v_405);
	assign v_386 = (v_384 & v_385);
	assign v_361 = (v_356 | v_360);
	assign v_579 = (v_577 & v_578);
	assign v_399 = (v_394 & v_398);
	assign v_412 = (v_394 | v_398);
	assign v_423 = (v_398 | v_422);
	assign v_383 = (v_381 & v_382);
	assign v_582 = (v_381 | v_382);
	assign v_407 = (v_402 & v_406);
	assign v_431 = (v_406 & v_430);
	assign v_411 = (v_402 | v_406);
	assign v_387 = (~v_382 & v_386);
	assign v_581 = (~v_382 | v_386);
	assign v_362 = (v_335 | v_361);
	assign v_580 = (v_576 & v_579);
	assign v_425 = (v_423 & v_424);
	assign v_408 = (v_399 | v_407);
	assign v_433 = (v_431 | v_432);
	assign v_413 = (v_411 & v_412);
	assign v_388 = (v_383 | v_387);
	assign v_583 = (v_581 & v_582);
	assign v_426 = (v_421 & v_425);
	assign v_439 = (v_421 | v_425);
	assign v_450 = (v_425 | v_449);
	assign v_410 = (v_408 & v_409);
	assign v_586 = (v_408 | v_409);
	assign v_434 = (v_429 & v_433);
	assign v_458 = (v_433 & v_457);
	assign v_438 = (v_429 | v_433);
	assign v_414 = (~v_409 & v_413);
	assign v_585 = (~v_409 | v_413);
	assign v_389 = (v_362 | v_388);
	assign v_584 = (v_580 & v_583);
	assign v_452 = (v_450 & v_451);
	assign v_435 = (v_426 | v_434);
	assign v_460 = (v_458 | v_459);
	assign v_440 = (v_438 & v_439);
	assign v_415 = (v_410 | v_414);
	assign v_587 = (v_585 & v_586);
	assign v_453 = (v_448 & v_452);
	assign v_466 = (v_448 | v_452);
	assign v_477 = (v_452 | v_476);
	assign v_437 = (v_435 & v_436);
	assign v_590 = (v_435 | v_436);
	assign v_461 = (v_456 & v_460);
	assign v_485 = (v_460 & v_484);
	assign v_465 = (v_456 | v_460);
	assign v_441 = (~v_436 & v_440);
	assign v_589 = (~v_436 | v_440);
	assign v_416 = (v_389 | v_415);
	assign v_588 = (v_584 & v_587);
	assign v_479 = (v_477 & v_478);
	assign v_462 = (v_453 | v_461);
	assign v_487 = (v_485 | v_486);
	assign v_467 = (v_465 & v_466);
	assign v_442 = (v_437 | v_441);
	assign v_591 = (v_589 & v_590);
	assign v_480 = (v_475 & v_479);
	assign v_493 = (v_475 | v_479);
	assign v_505 = (v_479 | v_504);
	assign v_464 = (v_462 & v_463);
	assign v_594 = (v_462 | v_463);
	assign v_488 = (v_483 & v_487);
	assign v_499 = (v_487 & v_498);
	assign v_492 = (v_483 | v_487);
	assign v_468 = (~v_463 & v_467);
	assign v_593 = (~v_463 | v_467);
	assign v_443 = (v_416 | v_442);
	assign v_592 = (v_588 & v_591);
	assign v_507 = (v_505 & v_506);
	assign v_489 = (v_480 | v_488);
	assign v_501 = (v_499 | v_500);
	assign v_494 = (v_492 & v_493);
	assign v_469 = (v_464 | v_468);
	assign v_595 = (v_593 & v_594);
	assign v_512 = (~v_502 & v_507);
	assign v_508 = (~v_502 | v_507);
	assign v_491 = (v_489 & v_490);
	assign v_598 = (v_489 | v_490);
	assign v_513 = (v_501 & v_502);
	assign v_503 = (v_501 | v_502);
	assign v_495 = (~v_490 & v_494);
	assign v_597 = (~v_490 | v_494);
	assign v_470 = (v_443 | v_469);
	assign v_596 = (v_592 & v_595);
	assign v_514 = (v_512 | v_513);
	assign v_509 = (v_503 & v_508);
	assign v_496 = (v_491 | v_495);
	assign v_599 = (v_597 & v_598);
	assign v_515 = (~v_510 & v_514);
	assign v_519 = (~v_510 | v_514);
	assign v_511 = (v_509 & v_510);
	assign v_520 = (v_509 | v_510);
	assign v_497 = (v_470 | v_496);
	assign v_600 = (v_596 & v_599);
	assign v_516 = (v_511 | v_515);
	assign v_521 = (v_519 & v_520);
	assign v_518 = (v_516 & v_517);
	assign v_602 = (v_516 | v_517);
	assign v_522 = (~v_517 & v_521);
	assign v_601 = (~v_517 | v_521);
	assign v_523 = (v_518 | v_522);
	assign v_603 = (v_601 & v_602);
	assign v_524 = (v_497 | v_523);
	assign v_604 = (v_600 & v_603);
	assign v_525 = (~v_7 | v_524);
	assign v_605 = (v_7 | v_604);
	assign v_617 = (((((((v_6 & v_525)) & v_605)) & v_609)) & v_611);
	assign v_615 = (v_617 & v_618);
	assign x_1 = (v_5 | v_615);
	assign o_1 = x_1;
endmodule
