// skolem function for order file variables
// Generated using findDep.cpp 
module small-dyn-partition-fixpoint-1 (v_1, v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_12, v_13, v_14, v_15, v_16, v_17, v_18, v_19, v_20, v_21, v_22, v_23, v_24, o_1);
input v_1;
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_13;
input v_14;
input v_15;
input v_16;
input v_17;
input v_18;
input v_19;
input v_20;
input v_21;
input v_22;
input v_23;
input v_24;
output o_1;
wire v_25;
wire v_26;
wire v_27;
wire v_28;
wire v_29;
wire v_30;
wire v_31;
wire v_32;
wire v_33;
wire v_34;
wire v_35;
wire v_36;
wire v_37;
wire v_38;
wire v_39;
wire v_40;
wire v_41;
wire v_42;
wire v_43;
wire v_44;
wire v_45;
wire v_46;
wire v_47;
wire v_48;
wire v_49;
wire v_50;
wire v_51;
wire v_52;
wire v_53;
wire v_54;
wire v_55;
wire v_56;
wire v_57;
wire v_58;
wire v_59;
wire v_60;
wire v_61;
wire v_62;
wire v_63;
wire v_64;
wire v_65;
wire v_66;
wire v_67;
wire v_68;
wire v_69;
wire v_70;
wire v_71;
wire v_72;
wire v_73;
wire v_74;
wire v_75;
wire v_76;
wire v_77;
wire v_78;
wire v_79;
wire v_80;
wire v_81;
wire v_82;
wire v_83;
wire v_84;
wire v_85;
wire v_86;
wire v_87;
wire x_1;
assign v_25 = ~v_1 & ~v_2 & ~v_3;
assign v_26 = ~v_4 & ~v_5 & ~v_6;
assign v_27 = ~v_7 & ~v_8 & v_25 & v_26;
assign v_29 = v_1;
assign v_31 = v_2 & v_29;
assign v_32 = v_31;
assign v_34 = v_3 & v_32;
assign v_35 = v_34;
assign v_36 = ~v_28 & ~v_1;
assign v_37 = v_28 & v_1;
assign v_39 = ~v_28 & v_30;
assign v_40 = v_28 & v_2;
assign v_42 = ~v_28 & v_33;
assign v_43 = v_28 & v_3;
assign v_48 = ~v_45 & ~v_46 & ~v_47;
assign v_49 = v_4;
assign v_51 = v_5 & v_49;
assign v_52 = v_51;
assign v_54 = v_6 & v_52;
assign v_55 = v_54;
assign v_56 = ~v_28 & v_4;
assign v_57 = ~v_4 & v_28;
assign v_59 = ~v_28 & v_5;
assign v_60 = v_28 & v_50;
assign v_62 = ~v_28 & v_6;
assign v_63 = v_28 & v_53;
assign v_68 = ~v_65 & ~v_66 & ~v_67;
assign v_71 = ~v_69 & ~v_70 & v_48 & v_68;
assign v_72 = v_27 & v_71;
assign v_73 = ~v_17 & ~v_18 & ~v_19;
assign v_74 = ~v_20 & ~v_21 & ~v_22;
assign v_75 = ~v_23 & ~v_24 & v_73 & v_74;
assign v_79 = ~v_76 & ~v_77 & ~v_78;
assign v_83 = ~v_80 & ~v_81 & ~v_82;
assign v_86 = ~v_84 & ~v_85 & v_79 & v_83;
assign v_87 = v_75 & v_86;
assign v_38 = v_36 | v_37;
assign v_41 = v_39 | v_40;
assign v_44 = v_42 | v_43;
assign v_58 = v_56 | v_57;
assign v_61 = v_59 | v_60;
assign v_64 = v_62 | v_63;
assign v_28 = v_8 ^ v_7;
assign v_30 = v_29 ^ v_2;
assign v_33 = v_32 ^ v_3;
assign v_45 = v_38 ^ v_9;
assign v_46 = v_41 ^ v_10;
assign v_47 = v_44 ^ v_11;
assign v_50 = v_49 ^ v_5;
assign v_53 = v_52 ^ v_6;
assign v_65 = v_58 ^ v_12;
assign v_66 = v_61 ^ v_13;
assign v_67 = v_64 ^ v_14;
assign v_69 = ~v_15 ^ v_8;
assign v_70 = v_7 ^ v_16;
assign v_76 = v_17 ^ v_9;
assign v_77 = v_18 ^ v_10;
assign v_78 = v_19 ^ v_11;
assign v_80 = v_20 ^ v_12;
assign v_81 = v_21 ^ v_13;
assign v_82 = v_22 ^ v_14;
assign v_84 = v_23 ^ v_15;
assign v_85 = v_24 ^ v_16;
assign x_1 = v_87 | ~v_72;
assign o_1 = x_1;
endmodule
