// skolem function for order file variables
// Generated using findDep.cpp 
module small-dyn-partition-fixpoint-2 (v_1, v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_12, v_13, v_14, v_15, v_16, v_17, v_18, v_19, v_20, v_21, v_22, v_23, v_24, v_25, v_26, v_27, v_28, v_29, v_30, v_31, v_32, v_33, v_34, v_35, v_36, v_37, v_38, v_39, v_40, o_1);
input v_1;
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_13;
input v_14;
input v_15;
input v_16;
input v_17;
input v_18;
input v_19;
input v_20;
input v_21;
input v_22;
input v_23;
input v_24;
input v_25;
input v_26;
input v_27;
input v_28;
input v_29;
input v_30;
input v_31;
input v_32;
input v_33;
input v_34;
input v_35;
input v_36;
input v_37;
input v_38;
input v_39;
input v_40;
output o_1;
wire v_41;
wire v_42;
wire v_43;
wire v_44;
wire v_45;
wire v_46;
wire v_47;
wire v_48;
wire v_49;
wire v_50;
wire v_51;
wire v_52;
wire v_53;
wire v_54;
wire v_55;
wire v_56;
wire v_57;
wire v_58;
wire v_59;
wire v_60;
wire v_61;
wire v_62;
wire v_63;
wire v_64;
wire v_65;
wire v_66;
wire v_67;
wire v_68;
wire v_69;
wire v_70;
wire v_71;
wire v_72;
wire v_73;
wire v_74;
wire v_75;
wire v_76;
wire v_77;
wire v_78;
wire v_79;
wire v_80;
wire v_81;
wire v_82;
wire v_83;
wire v_84;
wire v_85;
wire v_86;
wire v_87;
wire v_88;
wire v_89;
wire v_90;
wire v_91;
wire v_92;
wire v_93;
wire v_94;
wire v_95;
wire v_96;
wire v_97;
wire v_98;
wire v_99;
wire v_100;
wire v_101;
wire v_102;
wire v_103;
wire v_104;
wire v_105;
wire v_106;
wire v_107;
wire v_108;
wire v_109;
wire v_110;
wire v_111;
wire v_112;
wire v_113;
wire v_114;
wire v_115;
wire v_116;
wire v_117;
wire v_118;
wire v_119;
wire v_120;
wire v_121;
wire v_122;
wire v_123;
wire v_124;
wire v_125;
wire v_126;
wire v_127;
wire v_128;
wire v_129;
wire v_130;
wire v_131;
wire v_132;
wire v_133;
wire v_134;
wire v_135;
wire v_136;
wire v_137;
wire v_138;
wire v_139;
wire v_140;
wire v_141;
wire v_142;
wire v_143;
wire v_144;
wire v_145;
wire v_146;
wire v_147;
wire v_148;
wire v_149;
wire v_150;
wire v_151;
wire v_152;
wire v_153;
wire v_154;
wire v_155;
wire v_156;
wire v_157;
wire v_158;
wire v_159;
wire v_160;
wire v_161;
wire v_162;
wire v_163;
wire v_164;
wire v_165;
wire v_166;
wire v_167;
wire v_168;
wire v_169;
wire v_170;
wire v_171;
wire v_172;
wire v_173;
wire v_174;
wire v_175;
wire v_176;
wire v_177;
wire v_178;
wire v_179;
wire v_180;
wire v_181;
wire v_182;
wire v_183;
wire v_184;
wire v_185;
wire v_186;
wire v_187;
wire v_188;
wire v_189;
wire v_190;
wire v_191;
wire v_192;
wire v_193;
wire v_194;
wire v_195;
wire v_196;
wire v_197;
wire v_198;
wire v_199;
wire v_200;
wire v_201;
wire v_202;
wire v_203;
wire v_204;
wire x_1;
assign v_41 = ~v_1 & ~v_2 & ~v_3;
assign v_42 = ~v_4 & ~v_5 & ~v_6;
assign v_43 = ~v_7 & ~v_8 & v_41 & v_42;
assign v_45 = v_1;
assign v_47 = v_2 & v_45;
assign v_48 = v_47;
assign v_50 = v_3 & v_48;
assign v_51 = v_50;
assign v_52 = ~v_44 & ~v_1;
assign v_53 = v_44 & v_1;
assign v_55 = ~v_44 & v_46;
assign v_56 = v_44 & v_2;
assign v_58 = ~v_44 & v_49;
assign v_59 = v_44 & v_3;
assign v_64 = ~v_61 & ~v_62 & ~v_63;
assign v_65 = v_4;
assign v_67 = v_5 & v_65;
assign v_68 = v_67;
assign v_70 = v_6 & v_68;
assign v_71 = v_70;
assign v_72 = ~v_44 & v_4;
assign v_73 = ~v_4 & v_44;
assign v_75 = ~v_44 & v_5;
assign v_76 = v_44 & v_66;
assign v_78 = ~v_44 & v_6;
assign v_79 = v_44 & v_69;
assign v_84 = ~v_81 & ~v_82 & ~v_83;
assign v_87 = ~v_85 & ~v_86 & v_64 & v_84;
assign v_89 = v_9;
assign v_91 = v_10 & v_89;
assign v_92 = v_91;
assign v_94 = v_11 & v_92;
assign v_95 = v_94;
assign v_96 = ~v_88 & ~v_9;
assign v_97 = v_88 & v_9;
assign v_99 = ~v_88 & v_90;
assign v_100 = v_88 & v_10;
assign v_102 = ~v_88 & v_93;
assign v_103 = v_88 & v_11;
assign v_108 = ~v_105 & ~v_106 & ~v_107;
assign v_109 = v_12;
assign v_111 = v_13 & v_109;
assign v_112 = v_111;
assign v_114 = v_14 & v_112;
assign v_115 = v_114;
assign v_116 = ~v_88 & v_12;
assign v_117 = ~v_12 & v_88;
assign v_119 = ~v_88 & v_13;
assign v_120 = v_88 & v_110;
assign v_122 = ~v_88 & v_14;
assign v_123 = v_88 & v_113;
assign v_128 = ~v_125 & ~v_126 & ~v_127;
assign v_131 = ~v_129 & ~v_130 & v_108 & v_128;
assign v_132 = v_43 & v_87 & v_131;
assign v_133 = ~v_25 & ~v_26 & ~v_27;
assign v_134 = ~v_28 & ~v_29 & ~v_30;
assign v_135 = ~v_31 & ~v_32 & v_133 & v_134;
assign v_137 = v_25;
assign v_139 = v_26 & v_137;
assign v_140 = v_139;
assign v_142 = v_27 & v_140;
assign v_143 = v_142;
assign v_144 = ~v_136 & ~v_25;
assign v_145 = v_136 & v_25;
assign v_147 = ~v_136 & v_138;
assign v_148 = v_136 & v_26;
assign v_150 = ~v_136 & v_141;
assign v_151 = v_136 & v_27;
assign v_156 = ~v_153 & ~v_154 & ~v_155;
assign v_157 = v_28;
assign v_159 = v_29 & v_157;
assign v_160 = v_159;
assign v_162 = v_30 & v_160;
assign v_163 = v_162;
assign v_164 = ~v_136 & v_28;
assign v_165 = ~v_28 & v_136;
assign v_167 = ~v_136 & v_29;
assign v_168 = v_136 & v_158;
assign v_170 = ~v_136 & v_30;
assign v_171 = v_136 & v_161;
assign v_176 = ~v_173 & ~v_174 & ~v_175;
assign v_179 = ~v_177 & ~v_178 & v_156 & v_176;
assign v_180 = v_135 & v_179;
assign v_184 = ~v_181 & ~v_182 & ~v_183;
assign v_188 = ~v_185 & ~v_186 & ~v_187;
assign v_191 = ~v_189 & ~v_190 & v_184 & v_188;
assign v_195 = ~v_192 & ~v_193 & ~v_194;
assign v_199 = ~v_196 & ~v_197 & ~v_198;
assign v_202 = ~v_200 & ~v_201 & v_195 & v_199;
assign v_204 = v_180 & v_203;
assign v_54 = v_52 | v_53;
assign v_57 = v_55 | v_56;
assign v_60 = v_58 | v_59;
assign v_74 = v_72 | v_73;
assign v_77 = v_75 | v_76;
assign v_80 = v_78 | v_79;
assign v_98 = v_96 | v_97;
assign v_101 = v_99 | v_100;
assign v_104 = v_102 | v_103;
assign v_118 = v_116 | v_117;
assign v_121 = v_119 | v_120;
assign v_124 = v_122 | v_123;
assign v_146 = v_144 | v_145;
assign v_149 = v_147 | v_148;
assign v_152 = v_150 | v_151;
assign v_166 = v_164 | v_165;
assign v_169 = v_167 | v_168;
assign v_172 = v_170 | v_171;
assign v_203 = v_191 | v_202;
assign v_44 = v_8 ^ v_7;
assign v_46 = v_45 ^ v_2;
assign v_49 = v_48 ^ v_3;
assign v_61 = v_54 ^ v_9;
assign v_62 = v_57 ^ v_10;
assign v_63 = v_60 ^ v_11;
assign v_66 = v_65 ^ v_5;
assign v_69 = v_68 ^ v_6;
assign v_81 = v_74 ^ v_12;
assign v_82 = v_77 ^ v_13;
assign v_83 = v_80 ^ v_14;
assign v_85 = ~v_15 ^ v_8;
assign v_86 = v_7 ^ v_16;
assign v_88 = v_16 ^ v_15;
assign v_90 = v_89 ^ v_10;
assign v_93 = v_92 ^ v_11;
assign v_105 = v_98 ^ v_17;
assign v_106 = v_101 ^ v_18;
assign v_107 = v_104 ^ v_19;
assign v_110 = v_109 ^ v_13;
assign v_113 = v_112 ^ v_14;
assign v_125 = v_118 ^ v_20;
assign v_126 = v_121 ^ v_21;
assign v_127 = v_124 ^ v_22;
assign v_129 = ~v_23 ^ v_16;
assign v_130 = v_15 ^ v_24;
assign v_136 = v_32 ^ v_31;
assign v_138 = v_137 ^ v_26;
assign v_141 = v_140 ^ v_27;
assign v_153 = v_146 ^ v_33;
assign v_154 = v_149 ^ v_34;
assign v_155 = v_152 ^ v_35;
assign v_158 = v_157 ^ v_29;
assign v_161 = v_160 ^ v_30;
assign v_173 = v_166 ^ v_36;
assign v_174 = v_169 ^ v_37;
assign v_175 = v_172 ^ v_38;
assign v_177 = ~v_39 ^ v_32;
assign v_178 = v_31 ^ v_40;
assign v_181 = v_25 ^ v_17;
assign v_182 = v_26 ^ v_18;
assign v_183 = v_27 ^ v_19;
assign v_185 = v_28 ^ v_20;
assign v_186 = v_29 ^ v_21;
assign v_187 = v_30 ^ v_22;
assign v_189 = v_31 ^ v_23;
assign v_190 = v_32 ^ v_24;
assign v_192 = v_33 ^ v_17;
assign v_193 = v_34 ^ v_18;
assign v_194 = v_35 ^ v_19;
assign v_196 = v_36 ^ v_20;
assign v_197 = v_37 ^ v_21;
assign v_198 = v_38 ^ v_22;
assign v_200 = v_39 ^ v_23;
assign v_201 = v_40 ^ v_24;
assign x_1 = v_204 | ~v_132;
assign o_1 = x_1;
endmodule
