module formula(i_0,i_1,i_2,i_3, i_4, i_5, i_6, i_7, i_8, i_9, i_10,i_11,i_12,i_13, i_14, i_15, i_16, i_17, i_18, i_19, i_20,i_21,i_22,i_23, i_24, i_25, i_26, i_27, i_28, i_29, i_30,i_31,i_32,i_33, i_34, i_35, i_36, i_37, i_38, i_39, out);
	input i_0, i_1,i_2,i_3, i_4, i_5, i_6, i_7, i_8, i_9, i_10,i_11,i_12,i_13, i_14, i_15, i_16, i_17, i_18, i_19, i_20,i_21,i_22,i_23, i_24, i_25, i_26, i_27, i_28, i_29, i_30,i_31,i_32,i_33, i_34, i_35, i_36, i_37, i_38, i_39;
	output out;
	wire w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20;
	assign w1 = (~i_0 | i_20) & (i_0 | ~i_20);
	assign w2 = (~i_1 | i_21) & (i_1 | ~i_21);
	assign w3 = (~i_2 | i_22) & (i_2 | ~i_22);
	assign w4 = (~i_3 | i_23) & (i_3 | ~i_23);
	assign w5 = (~i_4 | i_24) & (i_4 | ~i_24);
	assign w6 = (~i_5 | i_25) & (i_5 | ~i_25);
	assign w7 = (~i_6 | i_26) & (i_6 | ~i_26);
	assign w8 = (~i_7 | i_27) & (i_7 | ~i_27);
	assign w9 = (~i_8 | i_28) & (i_8 | ~i_28);
	assign w10 = (~i_9 | i_29) & (i_9 | ~i_29);
	assign w11 = (~i_10 | i_30) & (i_10 | ~i_30);
	assign w12 = (~i_11 | i_31) & (i_11 | ~i_31);
	assign w13 = (~i_12 | i_32) & (i_12 | ~i_32);
	assign w14 = (~i_13 | i_33) & (i_13 | ~i_33);
	assign w15 = (~i_14 | i_34) & (i_14 | ~i_34);
	assign w16 = (~i_15 | i_35) & (i_15 | ~i_35);
	assign w17 = (~i_16 | i_36) & (i_16 | ~i_36);
	assign w18 = (~i_17 | i_37) & (i_17 | ~i_37);
	assign w19 = (~i_18 | i_38) & (i_18 | ~i_38);
	assign w20 = (~i_19 | i_39) & (i_19 | ~i_39);
	assign out = w1 & w2 & w3 & w4 & w5 & w6 & w7 & w8 & w9 & w10 & w11 & w12 & w13 & w14 & w15 & w16 & w17 & w18 & w19 & w20;
endmodule
