module SKOLEMFORMULA (i0, i1, i2, );
input i0;
input i1;
output i2;
assign i2 = 1;
endmodule