// Benchmark "SKOLEMFORMULA" written by ABC on Mon May 16 20:30:39 2022

module SKOLEMFORMULA ( 
    i0, i1,
    i2  );
  input  i0, i1;
  output i2;
  assign i2 = 1'b0;
endmodule


