// skolem function for order file variables
// Generated using findDep.cpp 
module small-bug1-fixpoint-10 (v_1, v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_12, v_13, v_14, v_15, v_16, v_17, v_18, v_19, v_20, v_21, v_22, v_23, v_24, v_25, v_26, v_27, v_28, v_29, v_30, v_31, v_32, v_33, v_34, v_35, v_36, v_37, v_38, v_39, v_40, v_41, v_42, v_43, v_44, v_45, v_46, v_47, v_48, v_49, v_50, v_51, v_52, v_53, v_54, v_55, v_56, v_57, v_58, v_59, v_60, v_61, o_1);
input v_1;
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_13;
input v_14;
input v_15;
input v_16;
input v_17;
input v_18;
input v_19;
input v_20;
input v_21;
input v_22;
input v_23;
input v_24;
input v_25;
input v_26;
input v_27;
input v_28;
input v_29;
input v_30;
input v_31;
input v_32;
input v_33;
input v_34;
input v_35;
input v_36;
input v_37;
input v_38;
input v_39;
input v_40;
input v_41;
input v_42;
input v_43;
input v_44;
input v_45;
input v_46;
input v_47;
input v_48;
input v_49;
input v_50;
input v_51;
input v_52;
input v_53;
input v_54;
input v_55;
input v_56;
input v_57;
input v_58;
input v_59;
input v_60;
input v_61;
output o_1;
wire v_62;
wire v_63;
wire v_64;
wire v_65;
wire v_66;
wire v_67;
wire v_68;
wire v_69;
wire v_70;
wire v_71;
wire v_72;
wire v_73;
wire v_74;
wire v_75;
wire v_76;
wire v_77;
wire v_78;
wire v_79;
wire v_80;
wire v_81;
wire v_82;
wire v_83;
wire v_84;
wire v_85;
wire v_86;
wire v_87;
wire v_88;
wire v_89;
wire v_90;
wire v_91;
wire v_92;
wire v_93;
wire v_94;
wire v_95;
wire v_96;
wire v_97;
wire v_98;
wire v_99;
wire v_100;
wire v_101;
wire v_102;
wire v_103;
wire v_104;
wire v_105;
wire v_106;
wire v_107;
wire v_108;
wire v_109;
wire v_110;
wire v_111;
wire v_112;
wire v_113;
wire v_114;
wire v_115;
wire v_116;
wire v_117;
wire v_118;
wire v_119;
wire v_120;
wire v_121;
wire v_122;
wire v_123;
wire v_124;
wire v_125;
wire v_126;
wire v_127;
wire v_128;
wire v_129;
wire v_130;
wire v_131;
wire v_132;
wire v_133;
wire v_134;
wire v_135;
wire v_136;
wire v_137;
wire v_138;
wire v_139;
wire v_140;
wire v_141;
wire v_142;
wire v_143;
wire v_144;
wire v_145;
wire v_146;
wire v_147;
wire v_148;
wire v_149;
wire v_150;
wire v_151;
wire v_152;
wire v_153;
wire v_154;
wire v_155;
wire v_156;
wire v_157;
wire v_158;
wire v_159;
wire v_160;
wire v_161;
wire v_162;
wire v_163;
wire v_164;
wire v_165;
wire v_166;
wire v_167;
wire v_168;
wire v_169;
wire v_170;
wire v_171;
wire v_172;
wire v_173;
wire v_174;
wire v_175;
wire v_176;
wire v_177;
wire v_178;
wire v_179;
wire v_180;
wire v_181;
wire v_182;
wire x_1;
assign v_62 = ~v_1 & v_14;
assign v_63 = ~v_13 & v_62;
assign v_66 = ~v_2 & v_12;
assign v_67 = ~v_16 & v_66;
assign v_70 = ~v_3 & v_15;
assign v_71 = ~v_18 & v_70;
assign v_74 = ~v_4 & v_17;
assign v_75 = ~v_20 & v_74;
assign v_78 = ~v_5 & v_19;
assign v_79 = ~v_22 & v_78;
assign v_82 = ~v_6 & v_21;
assign v_83 = ~v_24 & v_82;
assign v_86 = ~v_7 & v_23;
assign v_87 = ~v_26 & v_86;
assign v_90 = ~v_8 & v_25;
assign v_91 = ~v_28 & v_90;
assign v_94 = ~v_9 & v_27;
assign v_95 = ~v_30 & v_94;
assign v_98 = ~v_10 & v_29;
assign v_99 = ~v_32 & v_98;
assign v_102 = v_172 & v_173 & v_174 & v_175 & v_176;
assign v_103 = ~v_33 & v_45;
assign v_104 = ~v_44 & v_103;
assign v_107 = ~v_34 & v_43;
assign v_108 = ~v_47 & v_107;
assign v_111 = ~v_35 & v_46;
assign v_112 = ~v_49 & v_111;
assign v_115 = ~v_36 & v_48;
assign v_116 = ~v_51 & v_115;
assign v_119 = ~v_37 & v_50;
assign v_120 = ~v_53 & v_119;
assign v_123 = ~v_38 & v_52;
assign v_124 = ~v_55 & v_123;
assign v_127 = ~v_39 & v_54;
assign v_128 = ~v_57 & v_127;
assign v_131 = ~v_40 & v_56;
assign v_132 = ~v_59 & v_131;
assign v_135 = ~v_41 & v_58;
assign v_136 = ~v_61 & v_135;
assign v_139 = v_177 & v_178 & v_179 & v_180;
assign v_142 = ~v_140 & ~v_141;
assign v_145 = ~v_143 & ~v_144;
assign v_148 = ~v_146 & ~v_147;
assign v_151 = ~v_149 & ~v_150;
assign v_154 = ~v_152 & ~v_153;
assign v_157 = ~v_155 & ~v_156;
assign v_160 = ~v_158 & ~v_159;
assign v_163 = ~v_161 & ~v_162;
assign v_166 = ~v_164 & ~v_165;
assign v_169 = ~v_167 & ~v_168;
assign v_171 = v_139 & v_170;
assign v_172 = ~v_1 & ~v_2 & ~v_3 & ~v_4 & ~v_5;
assign v_173 = ~v_6 & ~v_7 & ~v_8 & ~v_9 & ~v_10;
assign v_174 = ~v_11 & ~v_65 & ~v_69 & ~v_73 & ~v_77;
assign v_175 = ~v_81 & ~v_85 & ~v_89 & ~v_93 & ~v_97;
assign v_176 = ~v_101;
assign v_177 = ~v_33 & ~v_34 & ~v_35 & ~v_36 & ~v_37;
assign v_178 = ~v_38 & ~v_39 & ~v_40 & ~v_41 & ~v_42;
assign v_179 = ~v_106 & ~v_110 & ~v_114 & ~v_118 & ~v_122;
assign v_180 = ~v_126 & ~v_130 & ~v_134 & ~v_138;
assign v_64 = v_13 | v_63;
assign v_68 = v_16 | v_67;
assign v_72 = v_18 | v_71;
assign v_76 = v_20 | v_75;
assign v_80 = v_22 | v_79;
assign v_84 = v_24 | v_83;
assign v_88 = v_26 | v_87;
assign v_92 = v_28 | v_91;
assign v_96 = v_30 | v_95;
assign v_100 = v_32 | v_99;
assign v_105 = v_44 | v_104;
assign v_109 = v_47 | v_108;
assign v_113 = v_49 | v_112;
assign v_117 = v_51 | v_116;
assign v_121 = v_53 | v_120;
assign v_125 = v_55 | v_124;
assign v_129 = v_57 | v_128;
assign v_133 = v_59 | v_132;
assign v_137 = v_61 | v_136;
assign v_170 = v_181 | v_182;
assign v_181 = v_142 | v_145 | v_148 | v_151 | v_154;
assign v_182 = v_157 | v_160 | v_163 | v_166 | v_169;
assign v_65 = v_64 ^ v_12;
assign v_69 = v_68 ^ v_15;
assign v_73 = v_72 ^ v_17;
assign v_77 = v_76 ^ v_19;
assign v_81 = v_80 ^ v_21;
assign v_85 = v_84 ^ v_23;
assign v_89 = v_88 ^ v_25;
assign v_93 = v_92 ^ v_27;
assign v_97 = v_96 ^ v_29;
assign v_101 = v_100 ^ v_31;
assign v_106 = v_105 ^ v_43;
assign v_110 = v_109 ^ v_46;
assign v_114 = v_113 ^ v_48;
assign v_118 = v_117 ^ v_50;
assign v_122 = v_121 ^ v_52;
assign v_126 = v_125 ^ v_54;
assign v_130 = v_129 ^ v_56;
assign v_134 = v_133 ^ v_58;
assign v_138 = v_137 ^ v_60;
assign v_140 = v_33 ^ v_11;
assign v_141 = v_45 ^ v_31;
assign v_143 = v_34 ^ v_11;
assign v_144 = v_43 ^ v_31;
assign v_146 = v_35 ^ v_11;
assign v_147 = v_46 ^ v_31;
assign v_149 = v_36 ^ v_11;
assign v_150 = v_48 ^ v_31;
assign v_152 = v_37 ^ v_11;
assign v_153 = v_50 ^ v_31;
assign v_155 = v_38 ^ v_11;
assign v_156 = v_52 ^ v_31;
assign v_158 = v_39 ^ v_11;
assign v_159 = v_54 ^ v_31;
assign v_161 = v_40 ^ v_11;
assign v_162 = v_56 ^ v_31;
assign v_164 = v_41 ^ v_11;
assign v_165 = v_58 ^ v_31;
assign v_167 = v_42 ^ v_11;
assign v_168 = v_60 ^ v_31;
assign x_1 = v_171 | ~v_102;
assign o_1 = x_1;
endmodule
