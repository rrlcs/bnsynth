// Verilog file written by procedure writeCombinationalCircuitInVerilog
//Skolem functions to be generated for i_ variables
module formula ( i_1, i_2, i_3, i_4, i_5, i_6, i_7, i_8, i_9, i_10, i_11, i_12, i_13, i_14, i_15, i_16, i_17, i_18, i_19, i_20, i_21, i_22, i_23, i_24, i_25, i_26, i_27, i_28, i_29, i_30, i_31, i_32, i_33, x_34, x_35, x_36, x_37, x_38, x_39, x_40, x_41, x_42, x_43, x_44, x_45, x_46, x_47, x_48, x_49, x_50, x_51, x_52, x_53, x_54, x_55, x_56, x_57, x_58, x_59, x_60, x_61, x_62, x_63, x_64, x_65, x_66, x_67, x_68, x_69, x_70, x_71, x_72, x_73, x_74, x_75, x_76, x_77, x_78, x_79, x_80, x_81, x_82, x_83, x_84, x_85, x_86, x_87, x_88, x_89, x_90, x_91, x_92, x_93, x_94, x_95, x_96, x_97, x_98, x_99, x_100, x_101, x_102, x_103, o_1 );
input i_1;
input i_2;
input i_3;
input i_4;
input i_5;
input i_6;
input i_7;
input i_8;
input i_9;
input i_10;
input i_11;
input i_12;
input i_13;
input i_14;
input i_15;
input i_16;
input i_17;
input i_18;
input i_19;
input i_20;
input i_21;
input i_22;
input i_23;
input i_24;
input i_25;
input i_26;
input i_27;
input i_28;
input i_29;
input i_30;
input i_31;
input i_32;
input i_33;
input x_34;
input x_35;
input x_36;
input x_37;
input x_38;
input x_39;
input x_40;
input x_41;
input x_42;
input x_43;
input x_44;
input x_45;
input x_46;
input x_47;
input x_48;
input x_49;
input x_50;
input x_51;
input x_52;
input x_53;
input x_54;
input x_55;
input x_56;
input x_57;
input x_58;
input x_59;
input x_60;
input x_61;
input x_62;
input x_63;
input x_64;
input x_65;
input x_66;
input x_67;
input x_68;
input x_69;
input x_70;
input x_71;
input x_72;
input x_73;
input x_74;
input x_75;
input x_76;
input x_77;
input x_78;
input x_79;
input x_80;
input x_81;
input x_82;
input x_83;
input x_84;
input x_85;
input x_86;
input x_87;
input x_88;
input x_89;
input x_90;
input x_91;
input x_92;
input x_93;
input x_94;
input x_95;
input x_96;
input x_97;
input x_98;
input x_99;
input x_100;
input x_101;
input x_102;
input x_103;
output o_1;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire n_53;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_58;
wire n_59;
wire n_60;
wire n_61;
wire n_62;
wire n_63;
wire n_64;
wire n_65;
wire n_66;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;
wire n_95;
wire n_96;
wire n_97;
wire n_98;
wire n_99;
wire n_100;
wire n_101;
wire n_102;
wire n_103;
wire n_104;
wire n_105;
wire n_106;
wire n_107;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_112;
wire n_113;
wire n_114;
wire n_115;
wire n_116;
wire n_117;
wire n_118;
wire n_119;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_124;
wire n_125;
wire n_126;
wire n_127;
wire n_128;
wire n_129;
wire n_130;
wire n_131;
wire n_132;
wire n_133;
wire n_134;
wire n_135;
wire n_136;
wire n_137;
wire n_138;
wire n_139;
wire n_140;
wire n_141;
wire n_142;
wire n_143;
wire n_144;
wire n_145;
wire n_146;
wire n_147;
wire n_148;
wire n_149;
wire n_150;
wire n_151;
wire n_152;
wire n_153;
wire n_154;
wire n_155;
wire n_156;
wire n_157;
wire n_158;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_163;
wire n_164;
wire n_165;
wire n_166;
wire n_167;
wire n_168;
wire n_169;
wire n_170;
wire n_171;
wire n_172;
wire n_173;
wire n_174;
wire n_175;
wire n_176;
wire n_177;
wire n_178;
wire n_179;
wire n_180;
wire n_181;
wire n_182;
wire n_183;
wire n_184;
wire n_185;
wire n_186;
wire n_187;
wire n_188;
wire n_189;
wire n_190;
wire n_191;
wire n_192;
wire n_193;
wire n_194;
wire n_195;
wire n_196;
wire n_197;
wire n_198;
wire n_199;
wire n_200;
wire n_201;
wire n_202;
wire n_203;
wire n_204;
wire n_205;
wire n_206;
wire n_207;
wire n_208;
wire n_209;
wire n_210;
wire n_211;
wire n_212;
wire n_213;
wire n_214;
wire n_215;
wire n_216;
wire n_217;
wire n_218;
wire n_219;
wire n_220;
wire n_221;
wire n_222;
wire n_223;
wire n_224;
wire n_225;
wire n_226;
wire n_227;
wire n_228;
wire n_229;
wire n_230;
wire n_231;
wire n_232;
wire n_233;
wire n_234;
wire n_235;
wire n_236;
wire n_237;
wire n_238;
wire n_239;
wire n_240;
wire n_241;
wire n_242;
wire n_243;
wire n_244;
wire n_245;
wire n_246;
wire n_247;
wire n_248;
wire n_249;
wire n_250;
wire n_251;
wire n_252;
wire n_253;
wire n_254;
wire n_255;
wire n_256;
wire n_257;
wire n_258;
wire n_259;
wire n_260;
wire n_261;
wire n_262;
wire n_263;
wire n_264;
wire n_265;
wire n_266;
wire n_267;
wire n_268;
wire n_269;
wire n_270;
wire n_271;
wire n_272;
wire n_273;
wire n_274;
wire n_275;
wire n_276;
wire n_277;
wire n_278;
wire n_279;
wire n_280;
wire n_281;
wire n_282;
wire n_283;
wire n_284;
wire n_285;
wire n_286;
wire n_287;
wire n_288;
wire n_289;
wire n_290;
wire n_291;
wire n_292;
wire n_293;
wire n_294;
wire n_295;
wire n_296;
wire n_297;
wire n_298;
wire n_299;
wire n_300;
wire n_301;
wire n_302;
wire n_303;
wire n_304;
wire n_305;
wire n_306;
wire n_307;
wire n_308;
wire n_309;
wire n_310;
wire n_311;
wire n_312;
wire n_313;
wire n_314;
wire n_315;
wire n_316;
wire n_317;
wire n_318;
wire n_319;
wire n_320;
wire n_321;
wire n_322;
wire n_323;
wire n_324;
wire n_325;
wire n_326;
wire n_327;
wire n_328;
wire n_329;
wire n_330;
wire n_331;
wire n_332;
wire n_333;
wire n_334;
wire n_335;
wire n_336;
wire n_337;
wire n_338;
wire n_339;
wire n_340;
wire n_341;
wire n_342;
wire n_343;
wire n_344;
wire n_345;
wire n_346;
wire n_347;
wire n_348;
wire n_349;
wire n_350;
wire n_351;
wire n_352;
wire n_353;
wire n_354;
wire n_355;
wire n_356;
wire n_357;
wire n_358;
wire n_359;
wire n_360;
wire n_361;
wire n_362;
wire n_363;
wire n_364;
wire n_365;
wire n_366;
wire n_367;
wire n_368;
wire n_369;
wire n_370;
wire n_371;
wire n_372;
wire n_373;
wire n_374;
wire n_375;
wire n_376;
wire n_377;
wire n_378;
wire n_379;
wire n_380;
wire n_381;
wire n_382;
wire n_383;
wire n_384;
wire n_385;
wire n_386;
wire n_387;
wire n_388;
wire n_389;
wire n_390;
wire n_391;
wire n_392;
wire n_393;
wire n_394;
wire n_395;
wire n_396;
wire n_397;
wire n_398;
wire n_399;
wire n_400;
wire n_401;
wire n_402;
wire n_403;
wire n_404;
wire n_405;
wire n_406;
wire n_407;
wire n_408;
wire n_409;
wire n_410;
wire n_411;
wire n_412;
wire n_413;
wire n_414;
wire n_415;
wire n_416;
wire n_417;
wire n_418;
wire n_419;
wire n_420;
wire n_421;
wire n_422;
wire n_423;
wire n_424;
wire n_425;
wire n_426;
wire n_427;
wire n_428;
wire n_429;
wire n_430;
wire n_431;
wire n_432;
wire n_433;
wire n_434;
wire n_435;
wire n_436;
wire n_437;
wire n_438;
wire n_439;
wire n_440;
wire n_441;
wire n_442;
wire n_443;
wire n_444;
wire n_445;
wire n_446;
wire n_447;
wire n_448;
wire n_449;
wire n_450;
wire n_451;
wire n_452;
wire n_453;
wire n_454;
wire n_455;
wire n_456;
wire n_457;
wire n_458;
wire n_459;
wire n_460;
wire n_461;
wire n_462;
wire n_463;
wire n_464;
wire n_465;
wire n_466;
wire n_467;
wire n_468;
wire n_469;
wire n_470;
wire n_471;
wire n_472;
wire n_473;
wire n_474;
wire n_475;
wire n_476;
wire n_477;
wire n_478;
wire n_479;
wire n_480;
wire n_481;
wire n_482;
wire n_483;
wire n_484;
wire n_485;
wire n_486;
wire n_487;
wire n_488;
wire n_489;
wire n_490;
wire n_491;
wire n_492;
wire n_493;
wire n_494;
wire n_495;
wire n_496;
wire n_497;
wire n_498;
wire n_499;
wire n_500;
wire n_501;
wire n_502;
wire n_503;
wire n_504;
wire n_505;
wire n_506;
wire n_507;
wire n_508;
wire n_509;
wire n_510;
wire n_511;
wire n_512;
wire n_513;
wire n_514;
wire n_515;
wire n_516;
wire n_517;
wire n_518;
wire n_519;
wire n_520;
wire n_521;
wire n_522;
wire n_523;
wire n_524;
wire n_525;
wire n_526;
wire n_527;
wire n_528;
wire n_529;
wire n_530;
wire n_531;
wire n_532;
wire n_533;
wire n_534;
wire n_535;
wire n_536;
wire n_537;
wire n_538;
wire n_539;
wire n_540;
wire n_541;
wire n_542;
wire n_543;
wire n_544;
wire n_545;
wire n_546;
wire n_547;
wire n_548;
wire n_549;
wire n_550;
wire n_551;
wire n_552;
wire n_553;
wire n_554;
wire n_555;
wire n_556;
wire n_557;
wire n_558;
wire n_559;
wire n_560;
wire n_561;
wire n_562;
wire n_563;
wire n_564;
wire n_565;
wire n_566;
wire n_567;
wire n_568;
wire n_569;
wire n_570;
wire n_571;
wire n_572;
wire n_573;
wire n_574;
wire n_575;
wire n_576;
wire n_577;
wire n_578;
wire n_579;
wire n_580;
wire n_581;
wire n_582;
wire n_583;
wire n_584;
wire n_585;
wire n_586;
wire n_587;
wire n_588;
wire n_589;
wire n_590;
wire n_591;
wire n_592;
wire n_593;
wire n_594;
wire n_595;
wire n_596;
wire n_597;
wire n_598;
wire n_599;
assign n_1 = ~i_11 & ~x_44;
assign n_2 =  i_11 &  x_44;
assign n_3 = ~n_1 & ~n_2;
assign n_4 = ~x_58 &  x_60;
assign n_5 = ~x_59 & ~n_4;
assign n_6 =  x_57 & ~n_5;
assign n_7 =  x_56 &  n_4;
assign n_8 = ~x_57 & ~x_59;
assign n_9 = ~n_7 &  n_8;
assign n_10 = ~n_6 & ~n_9;
assign n_11 = ~x_58 & ~x_59;
assign n_12 = ~x_56 & ~x_57;
assign n_13 =  x_60 & ~n_12;
assign n_14 =  n_11 &  n_13;
assign n_15 =  x_58 &  x_59;
assign n_16 = ~x_58 & ~n_12;
assign n_17 = ~x_60 & ~n_16;
assign n_18 = ~n_15 & ~n_17;
assign n_19 = ~n_14 &  n_18;
assign n_20 =  n_10 &  n_19;
assign n_21 = ~x_60 &  n_11;
assign n_22 =  x_57 & ~n_21;
assign n_23 = ~x_57 & ~x_58;
assign n_24 = ~n_22 & ~n_23;
assign n_25 = ~n_15 & ~n_24;
assign n_26 =  x_57 &  n_15;
assign n_27 = ~x_56 & ~n_23;
assign n_28 = ~n_26 &  n_27;
assign n_29 =  n_25 &  n_28;
assign n_30 =  n_20 &  n_29;
assign n_31 =  x_50 &  n_30;
assign n_32 = ~n_31 &  n_3;
assign n_33 =  i_11 &  n_31;
assign n_34 =  x_56 &  n_25;
assign n_35 = ~x_56 & ~n_25;
assign n_36 = ~n_34 & ~n_35;
assign n_37 = ~n_10 &  n_19;
assign n_38 =  x_56 & ~n_22;
assign n_39 = ~x_56 &  n_26;
assign n_40 = ~n_38 & ~n_39;
assign n_41 =  n_37 & ~n_40;
assign n_42 =  n_36 &  n_41;
assign n_43 = ~n_33 & ~n_42;
assign n_44 = ~n_32 &  n_43;
assign n_45 = ~n_10 & ~n_19;
assign n_46 =  n_22 &  n_34;
assign n_47 =  n_45 &  n_46;
assign n_48 = ~x_50 &  x_51;
assign n_49 =  n_3 & ~n_48;
assign n_50 =  i_11 &  n_48;
assign n_51 = ~n_49 & ~n_50;
assign n_52 =  n_42 &  n_51;
assign n_53 = ~n_47 & ~n_52;
assign n_54 = ~n_44 &  n_53;
assign n_55 = ~x_58 &  n_12;
assign n_56 =  n_37 &  n_55;
assign n_57 = ~x_49 & ~x_66;
assign n_58 =  x_36 &  x_44;
assign n_59 = ~n_57 &  n_58;
assign n_60 =  x_37 &  n_59;
assign n_61 =  i_11 &  n_60;
assign n_62 =  x_49 &  x_66;
assign n_63 =  n_60 & ~n_62;
assign n_64 =  n_59 & ~n_62;
assign n_65 = ~n_3 &  n_64;
assign n_66 =  n_3 & ~n_59;
assign n_67 = ~n_65 & ~n_66;
assign n_68 = ~n_63 &  n_67;
assign n_69 = ~n_61 & ~n_68;
assign n_70 =  n_47 &  n_69;
assign n_71 = ~n_56 & ~n_70;
assign n_72 = ~n_54 &  n_71;
assign n_73 =  x_40 &  x_49;
assign n_74 = ~x_40 & ~x_49;
assign n_75 = ~n_73 & ~n_74;
assign n_76 = ~x_63 &  x_64;
assign n_77 =  x_62 &  n_76;
assign n_78 = ~n_75 &  n_77;
assign n_79 = ~i_11 &  n_78;
assign n_80 =  n_74 &  n_77;
assign n_81 = ~n_3 & ~n_80;
assign n_82 = ~n_79 & ~n_81;
assign n_83 =  n_56 & ~n_82;
assign n_84 = ~n_39 & ~n_83;
assign n_85 = ~n_72 &  n_84;
assign n_86 = ~n_25 &  n_28;
assign n_87 =  n_10 & ~n_19;
assign n_88 =  n_86 &  n_87;
assign n_89 = ~x_62 &  n_76;
assign n_90 = ~n_75 &  n_89;
assign n_91 = ~i_11 &  n_90;
assign n_92 =  n_74 &  n_89;
assign n_93 = ~n_3 & ~n_92;
assign n_94 = ~n_91 & ~n_93;
assign n_95 =  n_39 &  n_94;
assign n_96 = ~n_88 & ~n_95;
assign n_97 = ~n_85 &  n_96;
assign n_98 =  n_29 &  n_37;
assign n_99 = ~x_62 &  x_63;
assign n_100 = ~x_64 &  n_99;
assign n_101 = ~x_34 & ~x_49;
assign n_102 =  x_66 &  n_101;
assign n_103 =  n_100 &  n_102;
assign n_104 = ~n_3 & ~n_103;
assign n_105 =  x_34 &  x_49;
assign n_106 = ~n_102 & ~n_105;
assign n_107 =  n_100 & ~n_106;
assign n_108 = ~x_45 &  x_47;
assign n_109 =  x_48 &  x_66;
assign n_110 = ~x_48 & ~x_66;
assign n_111 = ~n_109 & ~n_110;
assign n_112 = ~x_35 & ~n_111;
assign n_113 =  n_108 & ~n_112;
assign n_114 = ~n_3 & ~n_113;
assign n_115 = ~x_35 &  n_110;
assign n_116 =  n_108 & ~n_115;
assign n_117 =  i_11 &  n_116;
assign n_118 = ~n_114 & ~n_117;
assign n_119 = ~x_45 & ~n_118;
assign n_120 = ~n_3 & ~n_111;
assign n_121 =  i_11 & ~n_110;
assign n_122 = ~n_120 & ~n_121;
assign n_123 = ~x_46 &  n_122;
assign n_124 =  x_46 &  n_3;
assign n_125 =  x_45 & ~n_124;
assign n_126 = ~n_123 &  n_125;
assign n_127 = ~n_119 & ~n_126;
assign n_128 =  n_107 & ~n_127;
assign n_129 = ~n_104 & ~n_128;
assign n_130 =  n_88 & ~n_129;
assign n_131 = ~n_98 & ~n_130;
assign n_132 = ~n_97 &  n_131;
assign n_133 = ~n_36 & ~n_40;
assign n_134 =  n_20 &  n_133;
assign n_135 = ~x_39 &  x_62;
assign n_136 = ~x_63 & ~x_64;
assign n_137 =  n_135 &  n_136;
assign n_138 =  n_102 &  n_137;
assign n_139 = ~n_3 & ~n_138;
assign n_140 =  x_45 & ~x_46;
assign n_141 =  n_122 &  n_140;
assign n_142 = ~n_106 &  n_137;
assign n_143 =  n_3 & ~n_140;
assign n_144 =  n_142 & ~n_143;
assign n_145 = ~n_141 &  n_144;
assign n_146 = ~n_139 & ~n_145;
assign n_147 =  n_98 &  n_146;
assign n_148 = ~n_134 & ~n_147;
assign n_149 = ~n_132 &  n_148;
assign n_150 = ~x_38 &  n_3;
assign n_151 =  i_11 &  x_38;
assign n_152 = ~n_150 & ~n_151;
assign n_153 =  n_134 &  n_152;
assign n_154 = ~n_149 & ~n_153;
assign n_155 =  n_37 &  n_86;
assign n_156 = ~i_12 &  x_42;
assign n_157 = ~i_12 & ~x_45;
assign n_158 =  i_12 &  x_45;
assign n_159 = ~n_157 & ~n_158;
assign n_160 = ~x_42 & ~n_159;
assign n_161 = ~n_156 & ~n_160;
assign n_162 =  n_155 &  n_161;
assign n_163 = ~n_31 & ~n_159;
assign n_164 = ~i_12 &  n_31;
assign n_165 = ~n_155 & ~n_164;
assign n_166 = ~n_163 &  n_165;
assign n_167 = ~n_162 & ~n_166;
assign n_168 = ~n_39 & ~n_167;
assign n_169 =  i_13 &  n_90;
assign n_170 = ~i_13 &  x_46;
assign n_171 =  i_13 & ~x_46;
assign n_172 = ~n_170 & ~n_171;
assign n_173 = ~n_92 &  n_172;
assign n_174 = ~n_169 & ~n_173;
assign n_175 =  n_39 & ~n_174;
assign n_176 =  n_47 & ~n_60;
assign n_177 =  n_172 & ~n_176;
assign n_178 = ~n_64 &  n_172;
assign n_179 =  x_45 &  n_170;
assign n_180 =  x_45 &  x_46;
assign n_181 =  i_13 & ~n_180;
assign n_182 =  n_59 & ~n_181;
assign n_183 = ~n_179 &  n_182;
assign n_184 = ~n_178 & ~n_183;
assign n_185 = ~n_63 & ~n_184;
assign n_186 =  n_47 &  n_185;
assign n_187 = ~n_56 & ~n_186;
assign n_188 = ~n_177 &  n_187;
assign n_189 =  i_13 &  n_78;
assign n_190 = ~n_80 &  n_172;
assign n_191 = ~n_189 & ~n_190;
assign n_192 =  n_56 &  n_191;
assign n_193 = ~n_39 & ~n_192;
assign n_194 = ~n_188 &  n_193;
assign n_195 = ~n_175 & ~n_194;
assign n_196 = ~i_12 &  n_90;
assign n_197 = ~n_92 & ~n_159;
assign n_198 = ~n_196 & ~n_197;
assign n_199 =  n_39 &  n_198;
assign n_200 = ~n_88 & ~n_199;
assign n_201 = ~n_195 &  n_200;
assign n_202 = ~n_168 &  n_201;
assign n_203 = ~x_44 & ~x_45;
assign n_204 =  n_107 &  n_203;
assign n_205 =  i_12 &  n_204;
assign n_206 =  n_103 &  n_203;
assign n_207 = ~n_159 & ~n_206;
assign n_208 = ~n_205 & ~n_207;
assign n_209 = ~i_13 &  n_204;
assign n_210 =  n_172 & ~n_206;
assign n_211 = ~n_209 & ~n_210;
assign n_212 =  n_88 & ~n_211;
assign n_213 = ~n_208 &  n_212;
assign n_214 = ~n_202 & ~n_213;
assign n_215 = ~i_17 & ~i_18;
assign n_216 =  n_31 &  n_215;
assign n_217 = ~i_17 &  x_50;
assign n_218 =  i_18 & ~x_51;
assign n_219 = ~i_18 &  x_51;
assign n_220 = ~i_17 & ~n_219;
assign n_221 = ~n_218 &  n_220;
assign n_222 = ~x_50 & ~n_221;
assign n_223 = ~n_217 & ~n_222;
assign n_224 = ~n_31 &  n_223;
assign n_225 = ~n_216 & ~n_224;
assign n_226 = ~n_42 & ~n_225;
assign n_227 = ~x_50 & ~n_215;
assign n_228 = ~n_217 & ~n_227;
assign n_229 =  n_42 &  n_228;
assign n_230 = ~n_226 & ~n_229;
assign n_231 = ~i_20 & ~x_53;
assign n_232 =  i_20 &  x_53;
assign n_233 = ~n_231 & ~n_232;
assign n_234 = ~n_31 &  n_233;
assign n_235 = ~i_20 &  n_31;
assign n_236 = ~n_88 & ~n_235;
assign n_237 = ~n_234 &  n_236;
assign n_238 = ~i_20 &  n_204;
assign n_239 = ~n_206 & ~n_233;
assign n_240 = ~n_238 & ~n_239;
assign n_241 =  n_88 & ~n_240;
assign n_242 = ~n_98 & ~n_241;
assign n_243 = ~n_237 &  n_242;
assign n_244 = ~i_21 & ~x_66;
assign n_245 = ~i_21 & ~x_52;
assign n_246 =  i_21 &  x_52;
assign n_247 = ~n_245 & ~n_246;
assign n_248 =  x_66 &  n_247;
assign n_249 = ~n_244 & ~n_248;
assign n_250 =  n_108 & ~n_249;
assign n_251 =  n_142 &  n_203;
assign n_252 = ~i_21 & ~x_54;
assign n_253 =  i_21 &  x_54;
assign n_254 = ~n_252 & ~n_253;
assign n_255 = ~n_108 &  n_254;
assign n_256 =  n_251 & ~n_255;
assign n_257 = ~n_250 &  n_256;
assign n_258 =  n_138 &  n_203;
assign n_259 = ~n_254 & ~n_258;
assign n_260 =  n_98 & ~n_259;
assign n_261 = ~n_257 &  n_260;
assign n_262 = ~n_233 & ~n_258;
assign n_263 =  i_20 &  n_108;
assign n_264 =  n_251 &  n_263;
assign n_265 = ~n_262 & ~n_264;
assign n_266 =  i_15 & ~x_48;
assign n_267 = ~i_15 &  x_48;
assign n_268 = ~n_266 & ~n_267;
assign n_269 = ~n_265 &  n_268;
assign n_270 =  i_15 & ~x_66;
assign n_271 = ~i_15 &  x_66;
assign n_272 = ~n_270 & ~n_271;
assign n_273 = ~n_108 & ~n_233;
assign n_274 =  n_272 &  n_273;
assign n_275 =  n_251 &  n_274;
assign n_276 =  n_98 & ~n_275;
assign n_277 = ~n_269 &  n_276;
assign n_278 =  i_10 &  x_43;
assign n_279 = ~i_10 & ~x_43;
assign n_280 = ~n_278 & ~n_279;
assign n_281 =  x_67 & ~n_280;
assign n_282 = ~i_16 & ~x_49;
assign n_283 =  i_16 &  x_49;
assign n_284 = ~n_282 & ~n_283;
assign n_285 =  x_54 &  x_66;
assign n_286 = ~x_37 &  n_285;
assign n_287 =  x_52 &  x_66;
assign n_288 = ~x_35 &  n_287;
assign n_289 = ~n_286 & ~n_288;
assign n_290 = ~n_284 &  n_289;
assign n_291 =  n_281 &  n_290;
assign n_292 = ~n_277 &  n_291;
assign n_293 = ~n_261 &  n_292;
assign n_294 = ~n_243 &  n_293;
assign n_295 = ~n_230 &  n_294;
assign n_296 =  i_28 & ~x_61;
assign n_297 = ~i_28 &  x_61;
assign n_298 = ~n_296 & ~n_297;
assign n_299 =  n_107 & ~n_113;
assign n_300 =  n_206 & ~n_299;
assign n_301 =  n_298 & ~n_300;
assign n_302 = ~n_111 &  n_287;
assign n_303 = ~x_48 &  x_66;
assign n_304 = ~i_28 &  n_303;
assign n_305 =  i_28 & ~n_303;
assign n_306 = ~n_304 & ~n_305;
assign n_307 = ~n_112 &  n_306;
assign n_308 = ~n_302 &  n_307;
assign n_309 =  n_116 &  n_204;
assign n_310 = ~n_308 &  n_309;
assign n_311 = ~n_301 & ~n_310;
assign n_312 =  n_88 & ~n_311;
assign n_313 =  n_47 &  n_63;
assign n_314 =  n_298 & ~n_313;
assign n_315 = ~i_28 & ~n_285;
assign n_316 =  n_60 & ~n_315;
assign n_317 =  n_47 &  n_316;
assign n_318 = ~n_314 & ~n_317;
assign n_319 = ~n_88 & ~n_318;
assign n_320 = ~n_312 & ~n_319;
assign n_321 =  x_45 &  n_48;
assign n_322 =  n_42 &  n_321;
assign n_323 = ~n_268 & ~n_322;
assign n_324 = ~i_15 & ~x_43;
assign n_325 =  i_15 &  x_43;
assign n_326 = ~n_324 & ~n_325;
assign n_327 =  n_322 &  n_326;
assign n_328 = ~n_88 & ~n_327;
assign n_329 = ~n_323 &  n_328;
assign n_330 =  n_204 &  n_272;
assign n_331 = ~n_206 &  n_268;
assign n_332 = ~n_330 & ~n_331;
assign n_333 =  n_88 & ~n_332;
assign n_334 = ~n_98 & ~n_333;
assign n_335 = ~n_329 &  n_334;
assign n_336 = ~n_320 & ~n_335;
assign n_337 =  n_295 &  n_336;
assign n_338 = ~i_14 & ~x_47;
assign n_339 =  i_14 &  x_47;
assign n_340 = ~n_338 & ~n_339;
assign n_341 = ~n_258 & ~n_340;
assign n_342 =  i_14 &  n_251;
assign n_343 = ~n_341 & ~n_342;
assign n_344 =  n_98 & ~n_343;
assign n_345 =  x_42 &  n_155;
assign n_346 =  n_340 & ~n_345;
assign n_347 =  i_14 &  n_345;
assign n_348 = ~n_56 & ~n_347;
assign n_349 = ~n_346 &  n_348;
assign n_350 = ~i_14 &  n_78;
assign n_351 = ~n_80 & ~n_340;
assign n_352 = ~n_350 & ~n_351;
assign n_353 =  n_56 & ~n_352;
assign n_354 = ~n_88 & ~n_353;
assign n_355 = ~n_349 &  n_354;
assign n_356 =  i_14 &  n_204;
assign n_357 = ~n_206 & ~n_340;
assign n_358 = ~n_356 & ~n_357;
assign n_359 =  n_88 &  n_358;
assign n_360 = ~n_98 & ~n_359;
assign n_361 = ~n_355 &  n_360;
assign n_362 = ~n_344 & ~n_361;
assign n_363 = ~i_22 & ~x_55;
assign n_364 =  i_22 &  x_55;
assign n_365 = ~n_363 & ~n_364;
assign n_366 = ~x_44 &  n_140;
assign n_367 = ~n_111 & ~n_365;
assign n_368 = ~i_22 & ~n_110;
assign n_369 = ~n_367 & ~n_368;
assign n_370 =  n_366 &  n_369;
assign n_371 =  n_142 & ~n_370;
assign n_372 =  n_138 & ~n_371;
assign n_373 = ~n_365 & ~n_372;
assign n_374 =  n_366 &  n_371;
assign n_375 = ~n_373 & ~n_374;
assign n_376 =  n_98 & ~n_375;
assign n_377 = ~x_44 & ~n_369;
assign n_378 = ~x_46 & ~n_377;
assign n_379 =  x_46 &  n_365;
assign n_380 =  x_45 & ~n_379;
assign n_381 = ~n_378 &  n_380;
assign n_382 =  x_44 & ~n_365;
assign n_383 = ~n_113 & ~n_365;
assign n_384 =  i_22 & ~x_44;
assign n_385 =  n_116 &  n_384;
assign n_386 = ~n_383 & ~n_385;
assign n_387 = ~x_45 & ~n_386;
assign n_388 = ~n_382 & ~n_387;
assign n_389 = ~n_381 &  n_388;
assign n_390 =  n_107 & ~n_389;
assign n_391 = ~n_103 & ~n_365;
assign n_392 =  n_88 & ~n_391;
assign n_393 = ~n_390 &  n_392;
assign n_394 = ~n_176 & ~n_365;
assign n_395 = ~i_22 &  n_59;
assign n_396 = ~n_64 & ~n_365;
assign n_397 = ~n_395 & ~n_396;
assign n_398 = ~n_63 & ~n_397;
assign n_399 =  n_47 &  n_398;
assign n_400 = ~n_88 & ~n_399;
assign n_401 = ~n_394 &  n_400;
assign n_402 = ~n_98 & ~n_401;
assign n_403 = ~n_393 &  n_402;
assign n_404 = ~n_376 & ~n_403;
assign n_405 = ~n_362 & ~n_404;
assign n_406 =  n_337 &  n_405;
assign n_407 =  x_39 &  x_53;
assign n_408 =  n_20 &  n_407;
assign n_409 =  n_46 &  n_408;
assign n_410 = ~x_66 &  n_409;
assign n_411 = ~n_254 & ~n_410;
assign n_412 =  n_244 &  n_409;
assign n_413 = ~n_411 & ~n_412;
assign n_414 = ~n_30 & ~n_413;
assign n_415 = ~x_50 &  n_254;
assign n_416 =  x_43 & ~n_247;
assign n_417 =  i_21 & ~x_43;
assign n_418 =  x_50 & ~n_417;
assign n_419 = ~n_416 &  n_418;
assign n_420 = ~n_415 & ~n_419;
assign n_421 =  n_30 &  n_420;
assign n_422 = ~n_47 & ~n_421;
assign n_423 = ~n_414 &  n_422;
assign n_424 = ~x_66 &  n_59;
assign n_425 = ~n_254 & ~n_424;
assign n_426 =  n_59 &  n_244;
assign n_427 = ~n_425 & ~n_426;
assign n_428 =  n_47 &  n_427;
assign n_429 = ~n_88 & ~n_428;
assign n_430 = ~n_423 &  n_429;
assign n_431 = ~n_206 & ~n_254;
assign n_432 =  x_52 &  x_53;
assign n_433 =  x_48 & ~n_432;
assign n_434 =  n_62 & ~n_433;
assign n_435 =  n_116 &  n_434;
assign n_436 =  i_21 & ~n_435;
assign n_437 = ~i_21 &  n_434;
assign n_438 =  n_113 &  n_437;
assign n_439 =  n_204 & ~n_438;
assign n_440 = ~n_436 &  n_439;
assign n_441 = ~n_431 & ~n_440;
assign n_442 =  n_88 & ~n_441;
assign n_443 = ~n_98 & ~n_442;
assign n_444 = ~n_430 &  n_443;
assign n_445 = ~i_19 & ~x_52;
assign n_446 =  i_19 &  x_52;
assign n_447 = ~n_445 & ~n_446;
assign n_448 = ~x_66 &  n_108;
assign n_449 = ~i_19 &  n_448;
assign n_450 =  n_251 & ~n_449;
assign n_451 =  n_448 &  n_450;
assign n_452 =  n_447 & ~n_451;
assign n_453 =  n_98 & ~n_452;
assign n_454 = ~n_410 &  n_447;
assign n_455 =  i_19 &  n_410;
assign n_456 = ~n_30 & ~n_455;
assign n_457 = ~n_454 &  n_456;
assign n_458 = ~x_43 &  x_50;
assign n_459 = ~i_19 &  n_458;
assign n_460 =  n_447 & ~n_458;
assign n_461 = ~n_459 & ~n_460;
assign n_462 =  n_30 &  n_461;
assign n_463 = ~n_88 & ~n_462;
assign n_464 = ~n_457 &  n_463;
assign n_465 = ~i_19 &  n_204;
assign n_466 = ~n_206 & ~n_447;
assign n_467 = ~n_465 & ~n_466;
assign n_468 =  n_88 &  n_467;
assign n_469 = ~n_98 & ~n_468;
assign n_470 = ~n_464 &  n_469;
assign n_471 = ~n_453 & ~n_470;
assign n_472 = ~n_444 & ~n_471;
assign n_473 =  n_406 &  n_472;
assign n_474 = ~n_214 &  n_473;
assign n_475 = ~n_154 &  n_474;
assign n_476 =  x_68 & ~n_475;
assign n_477 = ~i_11 & ~i_12;
assign n_478 = ~i_13 & ~i_14;
assign n_479 =  n_477 &  n_478;
assign n_480 =  n_215 &  n_479;
assign n_481 =  i_15 &  i_16;
assign n_482 = ~i_15 & ~i_16;
assign n_483 = ~n_481 & ~n_482;
assign n_484 = ~i_19 & ~i_20;
assign n_485 = ~i_21 & ~i_22;
assign n_486 =  n_484 &  n_485;
assign n_487 = ~n_483 &  n_486;
assign n_488 =  n_480 &  n_487;
assign n_489 = ~x_68 & ~n_488;
assign n_490 = ~n_476 & ~n_489;
assign n_491 =  x_67 &  n_490;
assign n_492 = ~x_67 & ~n_490;
assign n_493 = ~n_491 & ~n_492;
assign n_494 =  i_33 &  x_66;
assign n_495 = ~i_33 & ~x_66;
assign n_496 = ~n_494 & ~n_495;
assign n_497 =  i_32 &  x_65;
assign n_498 = ~i_32 & ~x_65;
assign n_499 = ~n_497 & ~n_498;
assign n_500 =  i_31 &  x_64;
assign n_501 = ~i_31 & ~x_64;
assign n_502 = ~n_500 & ~n_501;
assign n_503 =  i_30 &  x_63;
assign n_504 = ~i_30 & ~x_63;
assign n_505 = ~n_503 & ~n_504;
assign n_506 =  i_29 &  x_62;
assign n_507 = ~i_29 & ~x_62;
assign n_508 = ~n_506 & ~n_507;
assign n_509 =  i_28 &  x_61;
assign n_510 = ~i_28 & ~x_61;
assign n_511 = ~n_509 & ~n_510;
assign n_512 =  i_27 &  x_60;
assign n_513 = ~i_27 & ~x_60;
assign n_514 = ~n_512 & ~n_513;
assign n_515 =  i_26 &  x_59;
assign n_516 = ~i_26 & ~x_59;
assign n_517 = ~n_515 & ~n_516;
assign n_518 =  i_25 &  x_58;
assign n_519 = ~i_25 & ~x_58;
assign n_520 = ~n_518 & ~n_519;
assign n_521 =  i_24 &  x_57;
assign n_522 = ~i_24 & ~x_57;
assign n_523 = ~n_521 & ~n_522;
assign n_524 =  i_23 &  x_56;
assign n_525 = ~i_23 & ~x_56;
assign n_526 = ~n_524 & ~n_525;
assign n_527 =  i_18 &  x_51;
assign n_528 = ~i_18 & ~x_51;
assign n_529 = ~n_527 & ~n_528;
assign n_530 =  i_17 &  x_50;
assign n_531 = ~i_17 & ~x_50;
assign n_532 = ~n_530 & ~n_531;
assign n_533 =  i_15 &  x_48;
assign n_534 = ~i_15 & ~x_48;
assign n_535 = ~n_533 & ~n_534;
assign n_536 =  i_13 &  x_46;
assign n_537 = ~i_13 & ~x_46;
assign n_538 = ~n_536 & ~n_537;
assign n_539 =  i_9 &  x_42;
assign n_540 = ~i_9 & ~x_42;
assign n_541 = ~n_539 & ~n_540;
assign n_542 =  i_8 &  x_41;
assign n_543 = ~i_8 & ~x_41;
assign n_544 = ~n_542 & ~n_543;
assign n_545 =  i_7 &  x_40;
assign n_546 = ~i_7 & ~x_40;
assign n_547 = ~n_545 & ~n_546;
assign n_548 =  i_6 &  x_39;
assign n_549 = ~i_6 & ~x_39;
assign n_550 = ~n_548 & ~n_549;
assign n_551 =  i_5 &  x_38;
assign n_552 = ~i_5 & ~x_38;
assign n_553 = ~n_551 & ~n_552;
assign n_554 =  i_4 &  x_37;
assign n_555 = ~i_4 & ~x_37;
assign n_556 = ~n_554 & ~n_555;
assign n_557 =  i_3 &  x_36;
assign n_558 = ~i_3 & ~x_36;
assign n_559 = ~n_557 & ~n_558;
assign n_560 =  i_2 &  x_35;
assign n_561 = ~i_2 & ~x_35;
assign n_562 = ~n_560 & ~n_561;
assign n_563 =  i_1 &  x_34;
assign n_564 = ~i_1 & ~x_34;
assign n_565 = ~n_563 & ~n_564;
assign n_566 = ~n_159 & ~n_233;
assign n_567 = ~n_254 &  n_566;
assign n_568 = ~n_280 &  n_567;
assign n_569 = ~n_284 &  n_568;
assign n_570 = ~n_340 &  n_569;
assign n_571 = ~n_365 &  n_570;
assign n_572 = ~n_447 &  n_571;
assign n_573 = ~n_565 &  n_572;
assign n_574 = ~n_562 &  n_573;
assign n_575 = ~n_559 &  n_574;
assign n_576 = ~n_556 &  n_575;
assign n_577 = ~n_553 &  n_576;
assign n_578 = ~n_550 &  n_577;
assign n_579 = ~n_547 &  n_578;
assign n_580 = ~n_544 &  n_579;
assign n_581 = ~n_541 &  n_580;
assign n_582 = ~n_538 &  n_581;
assign n_583 = ~n_535 &  n_582;
assign n_584 = ~n_532 &  n_583;
assign n_585 = ~n_529 &  n_584;
assign n_586 = ~n_526 &  n_585;
assign n_587 = ~n_523 &  n_586;
assign n_588 = ~n_520 &  n_587;
assign n_589 = ~n_517 &  n_588;
assign n_590 = ~n_514 &  n_589;
assign n_591 = ~n_511 &  n_590;
assign n_592 = ~n_508 &  n_591;
assign n_593 = ~n_505 &  n_592;
assign n_594 = ~n_502 &  n_593;
assign n_595 = ~n_499 &  n_594;
assign n_596 = ~n_496 &  n_595;
assign n_597 = ~n_493 &  n_596;
assign n_598 =  x_68 &  n_597;
assign n_599 = ~n_3 &  n_598;
assign o_1 = ~n_599;
endmodule

