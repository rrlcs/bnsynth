module SKOLEMFORMULA ( 
    inps, outs  );
  input  inps;
  output outs;
  wire net;
  constraint
endmodule