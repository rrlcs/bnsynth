// Benchmark "SKOLEMFORMULA" written by ABC on Tue May 17 20:55:23 2022

module SKOLEMFORMULA ( 
    i0,
    i1  );
  input  i0;
  output i1;
  assign i1 = 1'b1;
endmodule


