// skolem function for order file variables
// Generated using findDep.cpp 
module stmt124_966_965 (v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_12, v_17, v_19, v_21, v_22, v_23, v_26, v_28, v_30, v_31, v_33, v_35, v_37, v_38, v_40, v_42, v_44, v_46, v_48, v_50, v_52, v_55, v_56, v_63, v_65, v_69, v_73, v_75, v_77, v_81, v_88, v_93, v_98, v_101, v_102, v_109, v_110, v_114, v_118, v_119, v_122, v_126, v_130, v_132, v_134, v_136, v_138, v_139, v_143, v_147, v_149, v_153, v_157, v_162, v_164, v_168, v_344, v_345, v_346, v_347, v_348, v_349, v_350, v_351, v_355, v_360, v_362, v_364, v_365, v_366, v_369, v_371, v_373, v_374, v_376, v_378, v_380, v_381, v_383, v_385, v_387, v_389, v_391, v_393, v_395, v_398, v_399, v_406, v_408, v_412, v_416, v_418, v_420, v_424, v_431, v_436, v_441, v_444, v_445, v_452, v_453, v_457, v_461, v_462, v_465, v_469, v_473, v_475, v_477, v_479, v_481, v_482, v_486, v_490, v_492, v_496, v_500, v_505, v_507, v_511, o_1);
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_12;
input v_17;
input v_19;
input v_21;
input v_22;
input v_23;
input v_26;
input v_28;
input v_30;
input v_31;
input v_33;
input v_35;
input v_37;
input v_38;
input v_40;
input v_42;
input v_44;
input v_46;
input v_48;
input v_50;
input v_52;
input v_55;
input v_56;
input v_63;
input v_65;
input v_69;
input v_73;
input v_75;
input v_77;
input v_81;
input v_88;
input v_93;
input v_98;
input v_101;
input v_102;
input v_109;
input v_110;
input v_114;
input v_118;
input v_119;
input v_122;
input v_126;
input v_130;
input v_132;
input v_134;
input v_136;
input v_138;
input v_139;
input v_143;
input v_147;
input v_149;
input v_153;
input v_157;
input v_162;
input v_164;
input v_168;
input v_344;
input v_345;
input v_346;
input v_347;
input v_348;
input v_349;
input v_350;
input v_351;
input v_355;
input v_360;
input v_362;
input v_364;
input v_365;
input v_366;
input v_369;
input v_371;
input v_373;
input v_374;
input v_376;
input v_378;
input v_380;
input v_381;
input v_383;
input v_385;
input v_387;
input v_389;
input v_391;
input v_393;
input v_395;
input v_398;
input v_399;
input v_406;
input v_408;
input v_412;
input v_416;
input v_418;
input v_420;
input v_424;
input v_431;
input v_436;
input v_441;
input v_444;
input v_445;
input v_452;
input v_453;
input v_457;
input v_461;
input v_462;
input v_465;
input v_469;
input v_473;
input v_475;
input v_477;
input v_479;
input v_481;
input v_482;
input v_486;
input v_490;
input v_492;
input v_496;
input v_500;
input v_505;
input v_507;
input v_511;
output o_1;
wire v_1;
wire v_9;
wire v_10;
wire v_11;
wire v_13;
wire v_14;
wire v_15;
wire v_16;
wire v_18;
wire v_20;
wire v_24;
wire v_25;
wire v_27;
wire v_29;
wire v_32;
wire v_34;
wire v_36;
wire v_39;
wire v_41;
wire v_43;
wire v_45;
wire v_47;
wire v_49;
wire v_51;
wire v_53;
wire v_54;
wire v_57;
wire v_58;
wire v_59;
wire v_60;
wire v_61;
wire v_62;
wire v_64;
wire v_66;
wire v_67;
wire v_68;
wire v_70;
wire v_71;
wire v_72;
wire v_74;
wire v_76;
wire v_78;
wire v_79;
wire v_80;
wire v_82;
wire v_83;
wire v_84;
wire v_85;
wire v_86;
wire v_87;
wire v_89;
wire v_90;
wire v_91;
wire v_92;
wire v_94;
wire v_95;
wire v_96;
wire v_97;
wire v_99;
wire v_100;
wire v_103;
wire v_104;
wire v_105;
wire v_106;
wire v_107;
wire v_108;
wire v_111;
wire v_112;
wire v_113;
wire v_115;
wire v_116;
wire v_117;
wire v_120;
wire v_121;
wire v_123;
wire v_124;
wire v_125;
wire v_127;
wire v_128;
wire v_129;
wire v_131;
wire v_133;
wire v_135;
wire v_137;
wire v_140;
wire v_141;
wire v_142;
wire v_144;
wire v_145;
wire v_146;
wire v_148;
wire v_150;
wire v_151;
wire v_152;
wire v_154;
wire v_155;
wire v_156;
wire v_158;
wire v_159;
wire v_160;
wire v_161;
wire v_163;
wire v_165;
wire v_166;
wire v_167;
wire v_169;
wire v_170;
wire v_171;
wire v_172;
wire v_173;
wire v_174;
wire v_175;
wire v_176;
wire v_177;
wire v_178;
wire v_179;
wire v_180;
wire v_181;
wire v_182;
wire v_183;
wire v_184;
wire v_185;
wire v_186;
wire v_187;
wire v_188;
wire v_189;
wire v_190;
wire v_191;
wire v_192;
wire v_193;
wire v_194;
wire v_195;
wire v_196;
wire v_197;
wire v_198;
wire v_199;
wire v_200;
wire v_201;
wire v_202;
wire v_203;
wire v_204;
wire v_205;
wire v_206;
wire v_207;
wire v_208;
wire v_209;
wire v_210;
wire v_211;
wire v_212;
wire v_213;
wire v_214;
wire v_215;
wire v_216;
wire v_217;
wire v_218;
wire v_219;
wire v_220;
wire v_221;
wire v_222;
wire v_223;
wire v_224;
wire v_225;
wire v_226;
wire v_227;
wire v_228;
wire v_229;
wire v_230;
wire v_231;
wire v_232;
wire v_233;
wire v_234;
wire v_235;
wire v_236;
wire v_237;
wire v_238;
wire v_239;
wire v_240;
wire v_241;
wire v_242;
wire v_243;
wire v_244;
wire v_245;
wire v_246;
wire v_247;
wire v_248;
wire v_249;
wire v_250;
wire v_251;
wire v_252;
wire v_253;
wire v_254;
wire v_255;
wire v_256;
wire v_257;
wire v_258;
wire v_259;
wire v_260;
wire v_261;
wire v_262;
wire v_263;
wire v_264;
wire v_265;
wire v_266;
wire v_267;
wire v_268;
wire v_269;
wire v_270;
wire v_271;
wire v_272;
wire v_273;
wire v_274;
wire v_275;
wire v_276;
wire v_277;
wire v_278;
wire v_279;
wire v_280;
wire v_281;
wire v_282;
wire v_283;
wire v_284;
wire v_285;
wire v_286;
wire v_287;
wire v_288;
wire v_289;
wire v_290;
wire v_291;
wire v_292;
wire v_293;
wire v_294;
wire v_295;
wire v_296;
wire v_297;
wire v_298;
wire v_299;
wire v_300;
wire v_301;
wire v_302;
wire v_303;
wire v_304;
wire v_305;
wire v_306;
wire v_307;
wire v_308;
wire v_309;
wire v_310;
wire v_311;
wire v_312;
wire v_313;
wire v_314;
wire v_315;
wire v_316;
wire v_317;
wire v_318;
wire v_319;
wire v_320;
wire v_321;
wire v_322;
wire v_323;
wire v_324;
wire v_325;
wire v_326;
wire v_327;
wire v_328;
wire v_329;
wire v_330;
wire v_331;
wire v_332;
wire v_333;
wire v_334;
wire v_335;
wire v_336;
wire v_337;
wire v_338;
wire v_339;
wire v_340;
wire v_341;
wire v_342;
wire v_343;
wire v_352;
wire v_353;
wire v_354;
wire v_356;
wire v_357;
wire v_358;
wire v_359;
wire v_361;
wire v_363;
wire v_367;
wire v_368;
wire v_370;
wire v_372;
wire v_375;
wire v_377;
wire v_379;
wire v_382;
wire v_384;
wire v_386;
wire v_388;
wire v_390;
wire v_392;
wire v_394;
wire v_396;
wire v_397;
wire v_400;
wire v_401;
wire v_402;
wire v_403;
wire v_404;
wire v_405;
wire v_407;
wire v_409;
wire v_410;
wire v_411;
wire v_413;
wire v_414;
wire v_415;
wire v_417;
wire v_419;
wire v_421;
wire v_422;
wire v_423;
wire v_425;
wire v_426;
wire v_427;
wire v_428;
wire v_429;
wire v_430;
wire v_432;
wire v_433;
wire v_434;
wire v_435;
wire v_437;
wire v_438;
wire v_439;
wire v_440;
wire v_442;
wire v_443;
wire v_446;
wire v_447;
wire v_448;
wire v_449;
wire v_450;
wire v_451;
wire v_454;
wire v_455;
wire v_456;
wire v_458;
wire v_459;
wire v_460;
wire v_463;
wire v_464;
wire v_466;
wire v_467;
wire v_468;
wire v_470;
wire v_471;
wire v_472;
wire v_474;
wire v_476;
wire v_478;
wire v_480;
wire v_483;
wire v_484;
wire v_485;
wire v_487;
wire v_488;
wire v_489;
wire v_491;
wire v_493;
wire v_494;
wire v_495;
wire v_497;
wire v_498;
wire v_499;
wire v_501;
wire v_502;
wire v_503;
wire v_504;
wire v_506;
wire v_508;
wire v_509;
wire v_510;
wire v_512;
wire v_513;
wire v_514;
wire v_515;
wire v_516;
wire v_517;
wire v_518;
wire v_519;
wire v_520;
wire v_521;
wire v_522;
wire v_523;
wire v_524;
wire v_525;
wire v_526;
wire v_527;
wire v_528;
wire v_529;
wire v_530;
wire v_531;
wire v_532;
wire v_533;
wire v_534;
wire v_535;
wire v_536;
wire v_537;
wire v_538;
wire v_539;
wire v_540;
wire v_541;
wire v_542;
wire v_543;
wire v_544;
wire v_545;
wire v_546;
wire v_547;
wire v_548;
wire v_549;
wire v_550;
wire v_551;
wire v_552;
wire v_553;
wire v_554;
wire v_555;
wire v_556;
wire v_557;
wire v_558;
wire v_559;
wire v_560;
wire v_561;
wire v_562;
wire v_563;
wire v_564;
wire v_565;
wire v_566;
wire v_567;
wire v_568;
wire v_569;
wire v_570;
wire v_571;
wire v_572;
wire v_573;
wire v_574;
wire v_575;
wire v_576;
wire v_577;
wire v_578;
wire v_579;
wire v_580;
wire v_581;
wire v_582;
wire v_583;
wire v_584;
wire v_585;
wire v_586;
wire v_587;
wire v_588;
wire v_589;
wire v_590;
wire v_591;
wire v_592;
wire v_593;
wire v_594;
wire v_595;
wire v_596;
wire v_597;
wire v_598;
wire v_599;
wire v_600;
wire v_601;
wire v_602;
wire v_603;
wire v_604;
wire v_605;
wire v_606;
wire v_607;
wire v_608;
wire v_609;
wire v_610;
wire v_611;
wire v_612;
wire v_613;
wire v_614;
wire v_615;
wire v_616;
wire v_617;
wire v_618;
wire v_619;
wire v_620;
wire v_621;
wire v_622;
wire v_623;
wire v_624;
wire v_625;
wire v_626;
wire v_627;
wire v_628;
wire v_629;
wire v_630;
wire v_631;
wire v_632;
wire v_633;
wire v_634;
wire v_635;
wire v_636;
wire v_637;
wire v_638;
wire v_639;
wire v_640;
wire v_641;
wire v_642;
wire v_643;
wire v_644;
wire v_645;
wire v_646;
wire v_647;
wire v_648;
wire v_649;
wire v_650;
wire v_651;
wire v_652;
wire v_653;
wire v_654;
wire v_655;
wire v_656;
wire v_657;
wire v_658;
wire v_659;
wire v_660;
wire v_661;
wire v_662;
wire v_663;
wire v_664;
wire v_665;
wire v_666;
wire v_667;
wire v_668;
wire v_669;
wire v_670;
wire v_671;
wire v_672;
wire v_673;
wire v_674;
wire v_675;
wire v_676;
wire v_677;
wire v_678;
wire v_679;
wire v_680;
wire v_681;
wire v_682;
wire v_683;
wire v_684;
wire v_685;
wire v_686;
wire v_687;
wire v_688;
wire v_689;
wire v_690;
wire v_691;
wire v_692;
wire v_693;
wire v_694;
wire v_695;
wire v_696;
wire v_697;
wire v_698;
wire v_699;
wire v_700;
wire v_701;
wire v_702;
wire v_703;
wire v_704;
wire v_705;
wire v_706;
wire v_707;
wire v_708;
wire v_709;
wire v_710;
wire v_711;
wire v_712;
wire v_713;
wire v_714;
wire v_715;
wire v_716;
wire v_717;
wire v_718;
wire v_719;
wire v_720;
wire v_721;
wire v_722;
wire v_723;
wire v_724;
wire v_725;
wire v_726;
wire v_727;
wire v_728;
wire v_729;
wire v_730;
wire v_731;
wire v_732;
wire v_733;
wire v_734;
wire v_735;
wire v_736;
wire v_737;
wire v_738;
wire v_739;
wire v_740;
wire v_741;
wire v_742;
wire v_743;
wire v_744;
wire v_745;
wire v_746;
wire v_747;
wire v_748;
wire v_749;
wire v_750;
wire v_751;
wire v_752;
wire v_753;
wire v_754;
wire v_755;
wire v_756;
wire v_757;
wire v_758;
wire v_759;
wire v_760;
wire v_761;
wire v_762;
wire v_763;
wire v_764;
wire v_765;
wire v_766;
wire v_767;
wire v_768;
wire v_769;
wire v_770;
wire v_771;
wire v_772;
wire v_773;
wire v_774;
wire v_775;
wire v_776;
wire v_777;
wire v_778;
wire v_779;
wire v_780;
wire v_781;
wire v_782;
wire v_783;
wire v_784;
wire v_785;
wire v_786;
wire v_787;
wire v_788;
wire v_789;
wire v_790;
wire v_791;
wire v_792;
wire v_793;
wire v_794;
wire v_795;
wire v_796;
wire v_797;
wire x_1;
assign v_1 = 1;
assign v_13 = 1;
assign v_18 = 1;
assign v_20 = 1;
assign v_27 = 1;
assign v_32 = 1;
assign v_51 = 1;
assign v_74 = 1;
assign v_78 = 1;
assign v_89 = 1;
assign v_94 = 1;
assign v_99 = 1;
assign v_103 = 1;
assign v_169 = 1;
assign v_171 = 1;
assign v_259 = 1;
assign v_356 = 1;
assign v_361 = 1;
assign v_363 = 1;
assign v_370 = 1;
assign v_375 = 1;
assign v_394 = 1;
assign v_417 = 1;
assign v_421 = 1;
assign v_432 = 1;
assign v_437 = 1;
assign v_442 = 1;
assign v_446 = 1;
assign v_512 = 1;
assign v_516 = 1;
assign v_610 = 1;
assign v_9 = v_7 & v_8;
assign v_10 = v_7 & ~v_8;
assign v_14 = v_6 & v_11;
assign v_15 = ~v_6 & v_11;
assign v_24 = v_22 & ~v_23;
assign v_29 = v_28;
assign v_34 = ~v_33;
assign v_36 = v_33 & v_35;
assign v_39 = v_33 & ~v_35 & v_37 & v_38;
assign v_41 = v_33 & ~v_35 & v_37 & ~v_38 & ~v_40;
assign v_43 = v_33 & ~v_35 & ~v_37 & ~v_42;
assign v_45 = v_33 & ~v_35 & ~v_37 & v_42 & v_44;
assign v_47 = v_704 & v_705;
assign v_49 = v_706 & v_707;
assign v_53 = v_708 & v_709;
assign v_54 = v_710 & v_711;
assign v_57 = v_55 & v_56;
assign v_58 = v_55 & ~v_56;
assign v_60 = v_712 & v_713;
assign v_62 = ~v_28 & ~v_30 & v_61;
assign v_64 = ~v_28 & v_30 & ~v_63;
assign v_66 = ~v_28 & v_30 & v_63 & ~v_65;
assign v_67 = ~v_28 & v_30 & v_63 & v_65;
assign v_70 = v_68 & v_69;
assign v_71 = v_68 & ~v_69;
assign v_76 = v_21 & v_25 & v_72 & v_75;
assign v_79 = v_21 & v_25 & v_72 & ~v_75;
assign v_82 = v_80 & v_81;
assign v_83 = v_80 & ~v_81;
assign v_85 = v_5 & v_16 & v_84;
assign v_86 = ~v_5 & v_16;
assign v_90 = v_4 & v_87;
assign v_91 = ~v_4 & v_87;
assign v_95 = v_3 & v_92;
assign v_96 = ~v_3 & v_92;
assign v_100 = v_2 & v_97;
assign v_104 = v_101 & v_97;
assign v_105 = ~v_101 & v_97;
assign v_107 = ~v_2 & v_106;
assign v_111 = v_109 & v_110;
assign v_112 = v_109 & ~v_110;
assign v_115 = v_113 & v_114;
assign v_116 = v_113 & ~v_114;
assign v_120 = v_117 & ~v_118 & v_119;
assign v_121 = v_117 & ~v_118 & ~v_119;
assign v_123 = v_117 & v_118 & v_122;
assign v_124 = v_117 & v_118 & ~v_122;
assign v_127 = v_125 & v_126;
assign v_128 = v_125 & ~v_126;
assign v_131 = v_129 & v_130;
assign v_133 = v_129 & ~v_130 & v_132;
assign v_135 = v_129 & ~v_130 & ~v_132 & v_134;
assign v_137 = v_129 & ~v_130 & ~v_132 & ~v_134 & v_136;
assign v_140 = v_714 & v_715;
assign v_141 = v_716 & v_717;
assign v_144 = v_142 & v_143;
assign v_145 = v_142 & ~v_143;
assign v_148 = v_146 & v_147;
assign v_150 = v_718 & v_719;
assign v_151 = v_720 & v_721;
assign v_154 = v_152 & v_153;
assign v_155 = v_152 & ~v_153;
assign v_158 = v_156 & v_157;
assign v_159 = v_146 & ~v_147;
assign v_160 = v_156 & ~v_157;
assign v_163 = v_161 & ~v_162;
assign v_165 = v_161 & v_162 & v_164;
assign v_166 = v_161 & v_162 & ~v_164;
assign v_170 = v_108 & v_167;
assign v_172 = v_6;
assign v_174 = v_173 & ~v_21;
assign v_175 = v_173 & v_28;
assign v_176 = v_173 & ~v_28 & v_30 & v_63 & ~v_65;
assign v_177 = v_173 & ~v_28 & v_30 & v_63 & v_65;
assign v_178 = v_173 & ~v_28 & v_30 & ~v_63;
assign v_179 = v_173 & v_31;
assign v_180 = v_173 & ~v_31;
assign v_183 = v_181 & v_182;
assign v_184 = v_722 & v_723;
assign v_186 = v_181 & v_185;
assign v_188 = v_187 & ~v_28 & ~v_30 & v_61;
assign v_190 = v_189 & v_68 & v_69;
assign v_191 = v_189 & v_68 & ~v_69;
assign v_193 = v_192 & v_21 & v_25 & v_72 & v_75;
assign v_194 = v_192 & v_21 & v_25 & v_72 & ~v_75;
assign v_197 = v_195 & v_196;
assign v_199 = v_5 & v_198;
assign v_200 = ~v_5 & v_173;
assign v_202 = v_201 & ~v_88;
assign v_203 = v_201 & v_88;
assign v_205 = v_4 & v_204;
assign v_206 = ~v_4 & v_201;
assign v_208 = v_207 & ~v_93;
assign v_209 = v_207 & v_93;
assign v_211 = v_3 & v_210;
assign v_212 = ~v_3 & v_207;
assign v_214 = v_213 & ~v_98;
assign v_215 = v_213 & v_98;
assign v_217 = v_2 & v_216;
assign v_218 = v_213 & ~v_102;
assign v_219 = v_213 & v_102;
assign v_221 = v_101 & v_220;
assign v_222 = ~v_101 & v_213;
assign v_224 = ~v_2 & v_223;
assign v_226 = v_225 & ~v_109;
assign v_227 = v_225 & v_109 & v_110;
assign v_228 = v_225 & v_109 & ~v_110;
assign v_230 = v_229 & v_113 & v_114;
assign v_231 = v_229 & v_113 & ~v_114;
assign v_233 = v_232 & v_125 & v_126;
assign v_234 = v_232 & v_125 & ~v_126;
assign v_237 = v_235 & v_236;
assign v_238 = v_724 & v_725;
assign v_239 = v_726 & v_727;
assign v_241 = v_240 & v_152 & v_153;
assign v_242 = v_240 & v_152 & ~v_153;
assign v_244 = v_243 & v_156 & v_157;
assign v_245 = v_243 & v_156 & ~v_157;
assign v_246 = v_728 & v_729;
assign v_247 = v_730 & v_731;
assign v_249 = v_248 & v_142 & v_143;
assign v_250 = v_248 & v_142 & ~v_143;
assign v_252 = v_251 & v_146 & v_147;
assign v_253 = v_251 & v_146 & ~v_147;
assign v_257 = v_254 & v_256;
assign v_260 = v_6;
assign v_262 = v_261 & ~v_21;
assign v_263 = v_261 & v_28;
assign v_264 = v_261 & ~v_28 & v_30 & v_63 & ~v_65;
assign v_265 = v_261 & ~v_28 & v_30 & v_63 & v_65;
assign v_266 = v_261 & ~v_28 & v_30 & ~v_63;
assign v_267 = v_261 & v_31;
assign v_268 = v_261 & ~v_31;
assign v_271 = v_269 & v_270;
assign v_272 = v_732 & v_733;
assign v_273 = v_269 & v_185;
assign v_275 = v_274 & ~v_28 & ~v_30 & v_61;
assign v_277 = v_276 & v_68 & v_69;
assign v_278 = v_276 & v_68 & ~v_69;
assign v_280 = v_279 & v_21 & v_25 & v_72 & v_75;
assign v_281 = v_279 & v_21 & v_25 & v_72 & ~v_75;
assign v_283 = v_282 & v_196;
assign v_285 = v_5 & v_284;
assign v_286 = ~v_5 & v_261;
assign v_288 = v_287 & ~v_88;
assign v_289 = v_287 & v_88;
assign v_291 = v_4 & v_290;
assign v_292 = ~v_4 & v_287;
assign v_294 = v_293 & ~v_93;
assign v_295 = v_293 & v_93;
assign v_297 = v_3 & v_296;
assign v_298 = ~v_3 & v_293;
assign v_300 = v_299 & ~v_98;
assign v_301 = v_299 & v_98;
assign v_303 = v_2 & v_302;
assign v_304 = v_299 & ~v_102;
assign v_305 = v_299 & v_102;
assign v_307 = v_101 & v_306;
assign v_308 = ~v_101 & v_299;
assign v_310 = ~v_2 & v_309;
assign v_312 = v_311 & ~v_109;
assign v_313 = v_311 & v_109 & v_110;
assign v_314 = v_311 & v_109 & ~v_110;
assign v_316 = v_315 & v_113 & v_114;
assign v_317 = v_315 & v_113 & ~v_114;
assign v_319 = v_318 & v_125 & v_126;
assign v_320 = v_318 & v_125 & ~v_126;
assign v_323 = v_321 & v_322;
assign v_324 = v_734 & v_735;
assign v_325 = v_736 & v_737;
assign v_327 = v_326 & v_152 & v_153;
assign v_328 = v_326 & v_152 & ~v_153;
assign v_330 = v_329 & v_156 & v_157;
assign v_331 = v_329 & v_156 & ~v_157;
assign v_332 = v_738 & v_739;
assign v_333 = v_740 & v_741;
assign v_335 = v_334 & v_142 & v_143;
assign v_336 = v_334 & v_142 & ~v_143;
assign v_338 = v_337 & v_146 & v_147;
assign v_339 = v_337 & v_146 & ~v_147;
assign v_342 = v_340 & v_341;
assign v_352 = v_350 & v_351;
assign v_353 = v_350 & ~v_351;
assign v_357 = v_349 & v_354;
assign v_358 = ~v_349 & v_354;
assign v_367 = v_365 & ~v_366;
assign v_372 = v_371;
assign v_377 = ~v_376;
assign v_379 = v_376 & v_378;
assign v_382 = v_376 & ~v_378 & v_380 & v_381;
assign v_384 = v_376 & ~v_378 & v_380 & ~v_381 & ~v_383;
assign v_386 = v_376 & ~v_378 & ~v_380 & ~v_385;
assign v_388 = v_376 & ~v_378 & ~v_380 & v_385 & v_387;
assign v_390 = v_742 & v_743;
assign v_392 = v_744 & v_745;
assign v_396 = v_746 & v_747;
assign v_397 = v_748 & v_749;
assign v_400 = v_398 & v_399;
assign v_401 = v_398 & ~v_399;
assign v_403 = v_750 & v_751;
assign v_405 = ~v_371 & ~v_373 & v_404;
assign v_407 = ~v_371 & v_373 & ~v_406;
assign v_409 = ~v_371 & v_373 & v_406 & ~v_408;
assign v_410 = ~v_371 & v_373 & v_406 & v_408;
assign v_413 = v_411 & v_412;
assign v_414 = v_411 & ~v_412;
assign v_419 = v_364 & v_368 & v_415 & v_418;
assign v_422 = v_364 & v_368 & v_415 & ~v_418;
assign v_425 = v_423 & v_424;
assign v_426 = v_423 & ~v_424;
assign v_428 = v_348 & v_359 & v_427;
assign v_429 = ~v_348 & v_359;
assign v_433 = v_347 & v_430;
assign v_434 = ~v_347 & v_430;
assign v_438 = v_346 & v_435;
assign v_439 = ~v_346 & v_435;
assign v_443 = v_345 & v_440;
assign v_447 = v_444 & v_440;
assign v_448 = ~v_444 & v_440;
assign v_450 = ~v_345 & v_449;
assign v_454 = v_452 & v_453;
assign v_455 = v_452 & ~v_453;
assign v_458 = v_456 & v_457;
assign v_459 = v_456 & ~v_457;
assign v_463 = v_460 & ~v_461 & v_462;
assign v_464 = v_460 & ~v_461 & ~v_462;
assign v_466 = v_460 & v_461 & v_465;
assign v_467 = v_460 & v_461 & ~v_465;
assign v_470 = v_468 & v_469;
assign v_471 = v_468 & ~v_469;
assign v_474 = v_472 & v_473;
assign v_476 = v_472 & ~v_473 & v_475;
assign v_478 = v_472 & ~v_473 & ~v_475 & v_477;
assign v_480 = v_472 & ~v_473 & ~v_475 & ~v_477 & v_479;
assign v_483 = v_752 & v_753;
assign v_484 = v_754 & v_755;
assign v_487 = v_485 & v_486;
assign v_488 = v_485 & ~v_486;
assign v_491 = v_489 & v_490;
assign v_493 = v_756 & v_757;
assign v_494 = v_758 & v_759;
assign v_497 = v_495 & v_496;
assign v_498 = v_495 & ~v_496;
assign v_501 = v_499 & v_500;
assign v_502 = v_489 & ~v_490;
assign v_503 = v_499 & ~v_500;
assign v_506 = v_504 & ~v_505;
assign v_508 = v_504 & v_505 & v_507;
assign v_509 = v_504 & v_505 & ~v_507;
assign v_513 = v_344 & v_451 & v_510;
assign v_514 = ~v_344 & v_451 & v_510;
assign v_517 = v_349;
assign v_519 = v_518 & ~v_364;
assign v_520 = v_518 & v_371;
assign v_521 = v_518 & ~v_371 & v_373 & v_406 & ~v_408;
assign v_522 = v_518 & ~v_371 & v_373 & v_406 & v_408;
assign v_523 = v_518 & ~v_371 & v_373 & ~v_406;
assign v_524 = v_518 & v_374;
assign v_525 = v_518 & ~v_374;
assign v_528 = v_526 & v_527;
assign v_529 = v_760 & v_761;
assign v_531 = v_526 & v_530;
assign v_533 = v_532 & ~v_371 & ~v_373 & v_404;
assign v_535 = v_534 & v_411 & v_412;
assign v_536 = v_534 & v_411 & ~v_412;
assign v_538 = v_537 & v_364 & v_368 & v_415 & v_418;
assign v_539 = v_537 & v_364 & v_368 & v_415 & ~v_418;
assign v_542 = v_540 & v_541;
assign v_544 = v_348 & v_543;
assign v_545 = ~v_348 & v_518;
assign v_547 = v_546 & ~v_431;
assign v_548 = v_546 & v_431;
assign v_550 = v_347 & v_549;
assign v_551 = ~v_347 & v_546;
assign v_553 = v_552 & ~v_436;
assign v_554 = v_552 & v_436;
assign v_556 = v_346 & v_555;
assign v_557 = ~v_346 & v_552;
assign v_559 = v_558 & ~v_441;
assign v_560 = v_558 & v_441;
assign v_562 = v_345 & v_561;
assign v_563 = v_558 & ~v_445;
assign v_564 = v_558 & v_445;
assign v_566 = v_444 & v_565;
assign v_567 = ~v_444 & v_558;
assign v_569 = ~v_345 & v_568;
assign v_571 = v_570 & ~v_452;
assign v_572 = v_570 & v_452 & v_453;
assign v_573 = v_570 & v_452 & ~v_453;
assign v_575 = v_574 & v_456 & v_457;
assign v_576 = v_574 & v_456 & ~v_457;
assign v_578 = v_577 & v_468 & v_469;
assign v_579 = v_577 & v_468 & ~v_469;
assign v_582 = v_580 & v_581;
assign v_583 = v_762 & v_763;
assign v_584 = v_764 & v_765;
assign v_586 = v_585 & v_495 & v_496;
assign v_587 = v_585 & v_495 & ~v_496;
assign v_589 = v_588 & v_499 & v_500;
assign v_590 = v_588 & v_499 & ~v_500;
assign v_591 = v_766 & v_767;
assign v_592 = v_768 & v_769;
assign v_594 = v_593 & v_485 & v_486;
assign v_595 = v_593 & v_485 & ~v_486;
assign v_597 = v_596 & v_489 & v_490;
assign v_598 = v_596 & v_489 & ~v_490;
assign v_602 = v_599 & v_601;
assign v_604 = v_603 & ~v_511;
assign v_605 = v_603 & v_511;
assign v_607 = v_344 & v_606;
assign v_608 = ~v_344 & v_603;
assign v_611 = v_349;
assign v_613 = v_612 & ~v_364;
assign v_614 = v_612 & v_371;
assign v_615 = v_612 & ~v_371 & v_373 & v_406 & ~v_408;
assign v_616 = v_612 & ~v_371 & v_373 & v_406 & v_408;
assign v_617 = v_612 & ~v_371 & v_373 & ~v_406;
assign v_618 = v_612 & v_374;
assign v_619 = v_612 & ~v_374;
assign v_622 = v_620 & v_621;
assign v_623 = v_770 & v_771;
assign v_624 = v_620 & v_530;
assign v_626 = v_625 & ~v_371 & ~v_373 & v_404;
assign v_628 = v_627 & v_411 & v_412;
assign v_629 = v_627 & v_411 & ~v_412;
assign v_631 = v_630 & v_364 & v_368 & v_415 & v_418;
assign v_632 = v_630 & v_364 & v_368 & v_415 & ~v_418;
assign v_634 = v_633 & v_541;
assign v_636 = v_348 & v_635;
assign v_637 = ~v_348 & v_612;
assign v_639 = v_638 & ~v_431;
assign v_640 = v_638 & v_431;
assign v_642 = v_347 & v_641;
assign v_643 = ~v_347 & v_638;
assign v_645 = v_644 & ~v_436;
assign v_646 = v_644 & v_436;
assign v_648 = v_346 & v_647;
assign v_649 = ~v_346 & v_644;
assign v_651 = v_650 & ~v_441;
assign v_652 = v_650 & v_441;
assign v_654 = v_345 & v_653;
assign v_655 = v_650 & ~v_445;
assign v_656 = v_650 & v_445;
assign v_658 = v_444 & v_657;
assign v_659 = ~v_444 & v_650;
assign v_661 = ~v_345 & v_660;
assign v_663 = v_662 & ~v_452;
assign v_664 = v_662 & v_452 & v_453;
assign v_665 = v_662 & v_452 & ~v_453;
assign v_667 = v_666 & v_456 & v_457;
assign v_668 = v_666 & v_456 & ~v_457;
assign v_670 = v_669 & v_468 & v_469;
assign v_671 = v_669 & v_468 & ~v_469;
assign v_674 = v_672 & v_673;
assign v_675 = v_772 & v_773;
assign v_676 = v_774 & v_775;
assign v_678 = v_677 & v_495 & v_496;
assign v_679 = v_677 & v_495 & ~v_496;
assign v_681 = v_680 & v_499 & v_500;
assign v_682 = v_680 & v_499 & ~v_500;
assign v_683 = v_776 & v_777;
assign v_684 = v_778 & v_779;
assign v_686 = v_685 & v_485 & v_486;
assign v_687 = v_685 & v_485 & ~v_486;
assign v_689 = v_688 & v_489 & v_490;
assign v_690 = v_688 & v_489 & ~v_490;
assign v_693 = v_691 & v_692;
assign v_695 = v_694 & ~v_511;
assign v_696 = v_694 & v_511;
assign v_698 = v_344 & v_697;
assign v_699 = ~v_344 & v_694;
assign v_703 = ~v_701 & ~v_702 & v_515;
assign v_704 = v_33 & ~v_35 & v_37 & ~v_38 & v_40;
assign v_705 = v_46;
assign v_706 = v_33 & ~v_35 & v_37 & ~v_38 & v_40;
assign v_707 = ~v_46 & v_48;
assign v_708 = v_33 & ~v_35 & ~v_37 & v_42 & ~v_44;
assign v_709 = v_52;
assign v_710 = v_33 & ~v_35 & ~v_37 & v_42 & ~v_44;
assign v_711 = ~v_52;
assign v_712 = v_33 & ~v_35 & v_37 & ~v_38 & v_40;
assign v_713 = ~v_46 & ~v_48 & v_59;
assign v_714 = v_129 & ~v_130 & ~v_132 & ~v_134 & ~v_136;
assign v_715 = v_138 & v_139;
assign v_716 = v_129 & ~v_130 & ~v_132 & ~v_134 & ~v_136;
assign v_717 = v_138 & ~v_139;
assign v_718 = v_129 & ~v_130 & ~v_132 & ~v_134 & ~v_136;
assign v_719 = ~v_138 & v_149;
assign v_720 = v_129 & ~v_130 & ~v_132 & ~v_134 & ~v_136;
assign v_721 = ~v_138 & ~v_149;
assign v_722 = v_181 & v_33 & ~v_35 & v_37 & ~v_38;
assign v_723 = v_40 & ~v_46 & ~v_48 & v_59;
assign v_724 = v_235 & v_129 & ~v_130 & ~v_132 & ~v_134;
assign v_725 = ~v_136 & ~v_138 & v_149;
assign v_726 = v_235 & v_129 & ~v_130 & ~v_132 & ~v_134;
assign v_727 = ~v_136 & ~v_138 & ~v_149;
assign v_728 = v_235 & v_129 & ~v_130 & ~v_132 & ~v_134;
assign v_729 = ~v_136 & v_138 & v_139;
assign v_730 = v_235 & v_129 & ~v_130 & ~v_132 & ~v_134;
assign v_731 = ~v_136 & v_138 & ~v_139;
assign v_732 = v_269 & v_33 & ~v_35 & v_37 & ~v_38;
assign v_733 = v_40 & ~v_46 & ~v_48 & v_59;
assign v_734 = v_321 & v_129 & ~v_130 & ~v_132 & ~v_134;
assign v_735 = ~v_136 & ~v_138 & v_149;
assign v_736 = v_321 & v_129 & ~v_130 & ~v_132 & ~v_134;
assign v_737 = ~v_136 & ~v_138 & ~v_149;
assign v_738 = v_321 & v_129 & ~v_130 & ~v_132 & ~v_134;
assign v_739 = ~v_136 & v_138 & v_139;
assign v_740 = v_321 & v_129 & ~v_130 & ~v_132 & ~v_134;
assign v_741 = ~v_136 & v_138 & ~v_139;
assign v_742 = v_376 & ~v_378 & v_380 & ~v_381 & v_383;
assign v_743 = v_389;
assign v_744 = v_376 & ~v_378 & v_380 & ~v_381 & v_383;
assign v_745 = ~v_389 & v_391;
assign v_746 = v_376 & ~v_378 & ~v_380 & v_385 & ~v_387;
assign v_747 = v_395;
assign v_748 = v_376 & ~v_378 & ~v_380 & v_385 & ~v_387;
assign v_749 = ~v_395;
assign v_750 = v_376 & ~v_378 & v_380 & ~v_381 & v_383;
assign v_751 = ~v_389 & ~v_391 & v_402;
assign v_752 = v_472 & ~v_473 & ~v_475 & ~v_477 & ~v_479;
assign v_753 = v_481 & v_482;
assign v_754 = v_472 & ~v_473 & ~v_475 & ~v_477 & ~v_479;
assign v_755 = v_481 & ~v_482;
assign v_756 = v_472 & ~v_473 & ~v_475 & ~v_477 & ~v_479;
assign v_757 = ~v_481 & v_492;
assign v_758 = v_472 & ~v_473 & ~v_475 & ~v_477 & ~v_479;
assign v_759 = ~v_481 & ~v_492;
assign v_760 = v_526 & v_376 & ~v_378 & v_380 & ~v_381;
assign v_761 = v_383 & ~v_389 & ~v_391 & v_402;
assign v_762 = v_580 & v_472 & ~v_473 & ~v_475 & ~v_477;
assign v_763 = ~v_479 & ~v_481 & v_492;
assign v_764 = v_580 & v_472 & ~v_473 & ~v_475 & ~v_477;
assign v_765 = ~v_479 & ~v_481 & ~v_492;
assign v_766 = v_580 & v_472 & ~v_473 & ~v_475 & ~v_477;
assign v_767 = ~v_479 & v_481 & v_482;
assign v_768 = v_580 & v_472 & ~v_473 & ~v_475 & ~v_477;
assign v_769 = ~v_479 & v_481 & ~v_482;
assign v_770 = v_620 & v_376 & ~v_378 & v_380 & ~v_381;
assign v_771 = v_383 & ~v_389 & ~v_391 & v_402;
assign v_772 = v_672 & v_472 & ~v_473 & ~v_475 & ~v_477;
assign v_773 = ~v_479 & ~v_481 & v_492;
assign v_774 = v_672 & v_472 & ~v_473 & ~v_475 & ~v_477;
assign v_775 = ~v_479 & ~v_481 & ~v_492;
assign v_776 = v_672 & v_472 & ~v_473 & ~v_475 & ~v_477;
assign v_777 = ~v_479 & v_481 & v_482;
assign v_778 = v_672 & v_472 & ~v_473 & ~v_475 & ~v_477;
assign v_779 = ~v_479 & v_481 & ~v_482;
assign v_11 = ~v_7 | v_9 | v_10;
assign v_16 = v_14 | v_15;
assign v_25 = ~v_22 | v_24;
assign v_59 = ~v_55 | v_57 | v_58;
assign v_61 = v_780 | v_781 | v_782;
assign v_68 = v_62 | v_64 | v_66 | v_67;
assign v_72 = v_29 | v_70 | v_71;
assign v_80 = v_76 | v_79;
assign v_84 = ~v_21 | v_82 | v_83;
assign v_87 = v_85 | v_86;
assign v_92 = v_90 | v_91;
assign v_97 = v_95 | v_96;
assign v_106 = v_104 | v_105;
assign v_108 = v_100 | v_107;
assign v_113 = v_111 | v_112;
assign v_117 = v_115 | v_116;
assign v_125 = v_120 | v_121 | v_123 | v_124;
assign v_129 = v_127 | v_128;
assign v_142 = v_140 | v_141;
assign v_146 = v_144 | v_145;
assign v_152 = v_150 | v_151;
assign v_156 = v_154 | v_155;
assign v_161 = v_148 | v_158 | v_159 | v_160;
assign v_167 = v_783 | v_784;
assign v_173 = v_172 | ~v_6;
assign v_181 = v_179 | v_180;
assign v_182 = v_785 | v_786;
assign v_185 = v_53 | v_54;
assign v_187 = v_183 | v_184 | v_186;
assign v_189 = v_176 | v_177 | v_178 | v_188;
assign v_192 = v_175 | v_190 | v_191;
assign v_195 = v_193 | v_194;
assign v_196 = v_82 | v_83;
assign v_198 = v_174 | v_197;
assign v_201 = v_199 | v_200;
assign v_204 = v_202 | v_203;
assign v_207 = v_205 | v_206;
assign v_210 = v_208 | v_209;
assign v_213 = v_211 | v_212;
assign v_216 = v_214 | v_215;
assign v_220 = v_218 | v_219;
assign v_223 = v_221 | v_222;
assign v_225 = v_217 | v_224;
assign v_229 = v_227 | v_228;
assign v_232 = v_230 | v_231;
assign v_235 = v_233 | v_234;
assign v_236 = v_131 | v_133 | v_135 | v_137;
assign v_240 = v_238 | v_239;
assign v_243 = v_241 | v_242;
assign v_248 = v_246 | v_247;
assign v_251 = v_249 | v_250;
assign v_254 = v_244 | v_245 | v_252 | v_253;
assign v_255 = v_165 | v_166;
assign v_256 = v_163 | v_255;
assign v_258 = v_226 | v_237 | v_257;
assign v_261 = v_260 | ~v_6;
assign v_269 = v_267 | v_268;
assign v_270 = v_787 | v_788;
assign v_274 = v_271 | v_272 | v_273;
assign v_276 = v_264 | v_265 | v_266 | v_275;
assign v_279 = v_263 | v_277 | v_278;
assign v_282 = v_280 | v_281;
assign v_284 = v_262 | v_283;
assign v_287 = v_285 | v_286;
assign v_290 = v_288 | v_289;
assign v_293 = v_291 | v_292;
assign v_296 = v_294 | v_295;
assign v_299 = v_297 | v_298;
assign v_302 = v_300 | v_301;
assign v_306 = v_304 | v_305;
assign v_309 = v_307 | v_308;
assign v_311 = v_303 | v_310;
assign v_315 = v_313 | v_314;
assign v_318 = v_316 | v_317;
assign v_321 = v_319 | v_320;
assign v_322 = v_131 | v_133 | v_135 | v_137;
assign v_326 = v_324 | v_325;
assign v_329 = v_327 | v_328;
assign v_334 = v_332 | v_333;
assign v_337 = v_335 | v_336;
assign v_340 = v_330 | v_331 | v_338 | v_339;
assign v_341 = v_163 | v_255;
assign v_343 = v_312 | v_323 | v_342;
assign v_354 = ~v_350 | v_352 | v_353;
assign v_359 = v_357 | v_358;
assign v_368 = ~v_365 | v_367;
assign v_402 = ~v_398 | v_400 | v_401;
assign v_404 = v_789 | v_790 | v_791;
assign v_411 = v_405 | v_407 | v_409 | v_410;
assign v_415 = v_372 | v_413 | v_414;
assign v_423 = v_419 | v_422;
assign v_427 = ~v_364 | v_425 | v_426;
assign v_430 = v_428 | v_429;
assign v_435 = v_433 | v_434;
assign v_440 = v_438 | v_439;
assign v_449 = v_447 | v_448;
assign v_451 = v_443 | v_450;
assign v_456 = v_454 | v_455;
assign v_460 = v_458 | v_459;
assign v_468 = v_463 | v_464 | v_466 | v_467;
assign v_472 = v_470 | v_471;
assign v_485 = v_483 | v_484;
assign v_489 = v_487 | v_488;
assign v_495 = v_493 | v_494;
assign v_499 = v_497 | v_498;
assign v_504 = v_491 | v_501 | v_502 | v_503;
assign v_510 = v_792 | v_793;
assign v_515 = v_513 | v_514;
assign v_518 = v_517 | ~v_349;
assign v_526 = v_524 | v_525;
assign v_527 = v_794 | v_795;
assign v_530 = v_396 | v_397;
assign v_532 = v_528 | v_529 | v_531;
assign v_534 = v_521 | v_522 | v_523 | v_533;
assign v_537 = v_520 | v_535 | v_536;
assign v_540 = v_538 | v_539;
assign v_541 = v_425 | v_426;
assign v_543 = v_519 | v_542;
assign v_546 = v_544 | v_545;
assign v_549 = v_547 | v_548;
assign v_552 = v_550 | v_551;
assign v_555 = v_553 | v_554;
assign v_558 = v_556 | v_557;
assign v_561 = v_559 | v_560;
assign v_565 = v_563 | v_564;
assign v_568 = v_566 | v_567;
assign v_570 = v_562 | v_569;
assign v_574 = v_572 | v_573;
assign v_577 = v_575 | v_576;
assign v_580 = v_578 | v_579;
assign v_581 = v_474 | v_476 | v_478 | v_480;
assign v_585 = v_583 | v_584;
assign v_588 = v_586 | v_587;
assign v_593 = v_591 | v_592;
assign v_596 = v_594 | v_595;
assign v_599 = v_589 | v_590 | v_597 | v_598;
assign v_600 = v_508 | v_509;
assign v_601 = v_506 | v_600;
assign v_603 = v_571 | v_582 | v_602;
assign v_606 = v_604 | v_605;
assign v_609 = v_607 | v_608;
assign v_612 = v_611 | ~v_349;
assign v_620 = v_618 | v_619;
assign v_621 = v_796 | v_797;
assign v_625 = v_622 | v_623 | v_624;
assign v_627 = v_615 | v_616 | v_617 | v_626;
assign v_630 = v_614 | v_628 | v_629;
assign v_633 = v_631 | v_632;
assign v_635 = v_613 | v_634;
assign v_638 = v_636 | v_637;
assign v_641 = v_639 | v_640;
assign v_644 = v_642 | v_643;
assign v_647 = v_645 | v_646;
assign v_650 = v_648 | v_649;
assign v_653 = v_651 | v_652;
assign v_657 = v_655 | v_656;
assign v_660 = v_658 | v_659;
assign v_662 = v_654 | v_661;
assign v_666 = v_664 | v_665;
assign v_669 = v_667 | v_668;
assign v_672 = v_670 | v_671;
assign v_673 = v_474 | v_476 | v_478 | v_480;
assign v_677 = v_675 | v_676;
assign v_680 = v_678 | v_679;
assign v_685 = v_683 | v_684;
assign v_688 = v_686 | v_687;
assign v_691 = v_681 | v_682 | v_689 | v_690;
assign v_692 = v_506 | v_600;
assign v_694 = v_663 | v_674 | v_693;
assign v_697 = v_695 | v_696;
assign v_700 = v_698 | v_699;
assign v_780 = v_34 | v_36 | v_39 | v_41 | v_43;
assign v_781 = v_45 | v_47 | v_49 | v_53 | v_54;
assign v_782 = v_60;
assign v_783 = ~v_109 | v_131 | v_133 | v_135 | v_137;
assign v_784 = v_163 | v_165 | v_166;
assign v_785 = v_34 | v_36 | v_39 | v_41 | v_43;
assign v_786 = v_45 | v_47 | v_49;
assign v_787 = v_34 | v_36 | v_39 | v_41 | v_43;
assign v_788 = v_45 | v_47 | v_49;
assign v_789 = v_377 | v_379 | v_382 | v_384 | v_386;
assign v_790 = v_388 | v_390 | v_392 | v_396 | v_397;
assign v_791 = v_403;
assign v_792 = ~v_452 | v_474 | v_476 | v_478 | v_480;
assign v_793 = v_506 | v_508 | v_509;
assign v_794 = v_377 | v_379 | v_382 | v_384 | v_386;
assign v_795 = v_388 | v_390 | v_392;
assign v_796 = v_377 | v_379 | v_382 | v_384 | v_386;
assign v_797 = v_388 | v_390 | v_392;
assign v_701 = ~v_609 ^ ~v_258;
assign v_702 = ~v_700 ^ ~v_343;
assign x_1 = ~v_170 | v_703;
assign o_1 = x_1;
endmodule
