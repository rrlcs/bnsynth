// Benchmark "SKOLEMFORMULA" written by ABC on Fri May 20 20:57:26 2022

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, i14, i15,
    i16, i17, i18, i19,
    i20, i21, i22, i23, i24, i25, i26, i27, i28, i29, i30, i31, i32, i33,
    i34, i35, i36, i37, i38, i39  );
  input  i0, i1, i2, i3, i4, i5, i6, i7, i8, i9, i10, i11, i12, i13, i14,
    i15, i16, i17, i18, i19;
  output i20, i21, i22, i23, i24, i25, i26, i27, i28, i29, i30, i31, i32, i33,
    i34, i35, i36, i37, i38, i39;
  assign i20 = i0;
  assign i21 = i1;
  assign i22 = i2;
  assign i23 = i3;
  assign i24 = i4;
  assign i25 = i5;
  assign i26 = i6;
  assign i27 = i7;
  assign i28 = i8;
  assign i29 = i9;
  assign i30 = i10;
  assign i31 = i11;
  assign i32 = i12;
  assign i33 = i13;
  assign i34 = i14;
  assign i35 = i15;
  assign i36 = i16;
  assign i37 = i17;
  assign i38 = i18;
  assign i39 = i19;
endmodule


