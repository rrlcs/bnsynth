// Verilog file written by procedure writeCombinationalCircuitInVerilog
//Skolem functions to be generated for i_ variables
module formula ( i_1, i_2, i_3, i_4, i_5, i_6, i_7, i_8, i_9, i_10, i_11, i_12, i_13, i_14, i_15, i_16, i_17, i_18, i_19, i_20, i_21, i_22, i_23, i_24, i_25, i_26, i_27, i_28, i_29, i_30, i_31, i_32, i_33, i_34, i_35, i_36, i_37, i_38, i_39, i_40, i_41, i_42, i_43, i_44, i_45, i_46, i_47, i_48, i_49, i_50, i_51, i_52, i_53, i_54, i_55, i_56, i_57, i_58, i_59, i_60, i_61, i_62, i_63, i_64, i_65, i_66, i_67, i_68, i_69, i_70, i_71, i_72, i_73, i_74, i_75, i_76, i_77, i_78, i_79, i_80, i_81, i_82, i_83, i_84, i_85, i_86, i_87, i_88, i_89, i_90, i_91, i_92, i_93, i_94, i_95, i_96, i_97, i_98, i_99, i_100, i_101, i_102, i_103, i_104, i_105, i_106, i_107, i_108, i_109, i_110, i_111, i_112, i_113, i_114, i_115, i_116, i_117, i_118, i_119, i_120, i_121, i_122, i_123, i_124, i_125, i_126, i_127, i_128, i_129, i_130, i_131, i_132, i_133, i_134, i_135, i_136, i_137, i_138, i_139, i_140, i_141, i_142, i_143, i_144, i_145, i_146, i_147, i_148, i_149, i_150, i_151, i_152, i_153, i_154, i_155, i_156, i_157, i_158, i_159, i_160, i_161, i_162, i_163, i_164, i_165, i_166, i_167, i_168, i_169, i_170, i_171, i_172, i_173, i_174, i_175, i_176, i_177, i_178, i_179, i_180, i_181, i_182, i_183, i_184, i_185, i_186, i_187, i_188, i_189, i_190, i_191, i_192, i_193, i_194, i_195, i_196, i_197, i_198, i_199, i_200, i_201, i_202, i_203, i_204, i_205, i_206, i_207, i_208, i_209, i_210, i_211, i_212, i_213, i_214, i_215, i_216, i_217, i_218, i_219, i_220, i_221, i_222, i_223, i_224, x_225, x_226, x_227, x_228, x_229, x_230, x_231, x_232, x_233, x_234, x_235, x_236, x_237, x_238, x_239, x_240, x_241, x_242, x_243, x_244, x_245, x_246, x_247, x_248, x_249, x_250, x_251, x_252, x_253, x_254, x_255, x_256, x_257, x_258, x_259, x_260, x_261, x_262, x_263, x_264, x_265, x_266, x_267, x_268, x_269, x_270, x_271, x_272, x_273, x_274, x_275, x_276, x_277, x_278, x_279, x_280, x_281, x_282, x_283, x_284, x_285, x_286, x_287, x_288, x_289, x_290, x_291, x_292, x_293, x_294, x_295, x_296, x_297, x_298, x_299, x_300, x_301, x_302, x_303, x_304, x_305, x_306, x_307, x_308, x_309, x_310, x_311, x_312, x_313, x_314, x_315, x_316, x_317, x_318, x_319, x_320, x_321, x_322, x_323, x_324, x_325, x_326, x_327, x_328, x_329, x_330, x_331, x_332, x_333, x_334, x_335, x_336, x_337, x_338, x_339, x_340, x_341, x_342, x_343, x_344, x_345, x_346, x_347, x_348, x_349, x_350, x_351, x_352, x_353, x_354, x_355, x_356, x_357, x_358, x_359, x_360, x_361, x_362, x_363, x_364, x_365, x_366, x_367, x_368, x_369, x_370, x_371, x_372, x_373, x_374, x_375, x_376, x_377, x_378, x_379, x_380, x_381, x_382, x_383, x_384, x_385, x_386, x_387, x_388, x_389, x_390, x_391, x_392, x_393, x_394, x_395, x_396, x_397, x_398, x_399, x_400, x_401, x_402, x_403, x_404, x_405, x_406, x_407, x_408, x_409, x_410, x_411, x_412, x_413, x_414, x_415, x_416, x_417, x_418, x_419, x_420, x_421, x_422, x_423, x_424, x_425, x_426, x_427, x_428, x_429, x_430, x_431, x_432, x_433, x_434, x_435, x_436, x_437, x_438, x_439, x_440, x_441, x_442, x_443, x_444, x_445, x_446, x_447, x_448, x_449, x_450, x_451, x_452, x_453, x_454, x_455, x_456, x_457, x_458, x_459, x_460, x_461, x_462, x_463, x_464, x_465, x_466, x_467, x_468, x_469, x_470, x_471, x_472, x_473, x_474, x_475, x_476, x_477, x_478, x_479, x_480, x_481, x_482, x_483, x_484, x_485, x_486, x_487, x_488, x_489, x_490, x_491, x_492, x_493, x_494, x_495, x_496, x_497, x_498, x_499, x_500, x_501, x_502, x_503, x_504, x_505, x_506, x_507, x_508, x_509, x_510, x_511, x_512, x_513, x_514, x_515, x_516, x_517, x_518, x_519, x_520, x_521, x_522, x_523, x_524, x_525, x_526, x_527, x_528, x_529, x_530, x_531, x_532, x_533, x_534, x_535, x_536, x_537, x_538, x_539, x_540, x_541, x_542, x_543, x_544, x_545, x_546, x_547, x_548, x_549, x_550, x_551, x_552, x_553, x_554, x_555, x_556, x_557, x_558, x_559, x_560, x_561, x_562, x_563, x_564, x_565, x_566, x_567, x_568, x_569, x_570, x_571, x_572, x_573, x_574, x_575, x_576, x_577, x_578, x_579, x_580, x_581, x_582, x_583, x_584, x_585, x_586, x_587, x_588, x_589, x_590, x_591, x_592, x_593, x_594, x_595, x_596, x_597, x_598, x_599, x_600, x_601, x_602, x_603, x_604, x_605, x_606, x_607, x_608, x_609, x_610, x_611, x_612, x_613, x_614, x_615, x_616, x_617, x_618, x_619, x_620, x_621, x_622, x_623, x_624, x_625, x_626, x_627, x_628, x_629, x_630, x_631, x_632, x_633, x_634, x_635, x_636, x_637, x_638, x_639, x_640, x_641, x_642, x_643, x_644, x_645, x_646, x_647, x_648, x_649, x_650, x_651, x_652, x_653, x_654, x_655, x_656, x_657, x_658, x_659, x_660, x_661, x_662, x_663, x_664, x_665, x_666, x_667, x_668, x_669, x_670, x_671, x_672, x_673, x_674, x_675, x_676, x_677, x_678, x_679, x_680, x_681, x_682, x_683, x_684, x_685, x_686, x_687, x_688, x_689, x_690, x_691, x_692, x_693, x_694, x_695, x_696, x_697, x_698, x_699, x_700, x_701, x_702, x_703, x_704, x_705, x_706, x_707, x_708, x_709, x_710, x_711, x_712, x_713, x_714, x_715, x_716, x_717, x_718, x_719, x_720, x_721, x_722, x_723, x_724, x_725, x_726, x_727, x_728, x_729, x_730, x_731, x_732, x_733, x_734, x_735, x_736, x_737, x_738, x_739, x_740, x_741, x_742, x_743, x_744, x_745, x_746, x_747, x_748, x_749, x_750, x_751, x_752, x_753, x_754, x_755, x_756, x_757, x_758, x_759, x_760, x_761, x_762, x_763, x_764, x_765, x_766, x_767, x_768, x_769, x_770, x_771, x_772, x_773, x_774, x_775, x_776, x_777, x_778, x_779, x_780, x_781, x_782, x_783, x_784, x_785, x_786, x_787, x_788, x_789, x_790, x_791, x_792, x_793, x_794, x_795, x_796, x_797, x_798, x_799, x_800, x_801, x_802, x_803, x_804, x_805, x_806, x_807, x_808, x_809, x_810, x_811, x_812, x_813, x_814, x_815, x_816, x_817, x_818, x_819, x_820, x_821, x_822, x_823, x_824, x_825, x_826, x_827, x_828, x_829, x_830, x_831, x_832, x_833, x_834, x_835, x_836, x_837, x_838, x_839, x_840, x_841, x_842, x_843, x_844, x_845, x_846, x_847, x_848, x_849, x_850, x_851, x_852, x_853, x_854, x_855, x_856, x_857, x_858, x_859, x_860, x_861, x_862, x_863, x_864, x_865, x_866, x_867, x_868, x_869, x_870, x_871, x_872, x_873, x_874, x_875, x_876, x_877, x_878, x_879, x_880, x_881, x_882, x_883, x_884, x_885, x_886, x_887, x_888, x_889, x_890, x_891, x_892, x_893, x_894, x_895, x_896, x_897, x_898, x_899, x_900, x_901, x_902, x_903, x_904, x_905, x_906, x_907, x_908, x_909, x_910, x_911, x_912, x_913, x_914, x_915, x_916, x_917, x_918, x_919, x_920, x_921, x_922, x_923, x_924, x_925, x_926, x_927, x_928, x_929, x_930, x_931, x_932, x_933, x_934, x_935, x_936, x_937, x_938, x_939, x_940, x_941, x_942, x_943, x_944, x_945, x_946, x_947, x_948, x_949, x_950, x_951, x_952, x_953, x_954, x_955, x_956, x_957, x_958, x_959, x_960, x_961, x_962, x_963, x_964, x_965, x_966, x_967, x_968, x_969, x_970, x_971, x_972, x_973, x_974, x_975, x_976, x_977, x_978, x_979, x_980, x_981, x_982, x_983, x_984, x_985, x_986, x_987, x_988, x_989, x_990, x_991, x_992, x_993, x_994, x_995, x_996, x_997, x_998, x_999, x_1000, x_1001, x_1002, x_1003, x_1004, x_1005, x_1006, x_1007, x_1008, x_1009, x_1010, x_1011, x_1012, x_1013, x_1014, x_1015, x_1016, x_1017, x_1018, x_1019, x_1020, x_1021, x_1022, x_1023, x_1024, x_1025, x_1026, x_1027, x_1028, x_1029, x_1030, x_1031, x_1032, x_1033, x_1034, x_1035, x_1036, x_1037, x_1038, x_1039, x_1040, x_1041, x_1042, x_1043, x_1044, x_1045, x_1046, x_1047, x_1048, x_1049, x_1050, x_1051, x_1052, x_1053, x_1054, x_1055, x_1056, x_1057, x_1058, x_1059, x_1060, x_1061, x_1062, x_1063, x_1064, x_1065, x_1066, x_1067, x_1068, x_1069, x_1070, x_1071, x_1072, x_1073, x_1074, x_1075, x_1076, x_1077, x_1078, x_1079, x_1080, x_1081, x_1082, x_1083, x_1084, x_1085, x_1086, x_1087, x_1088, x_1089, x_1090, x_1091, x_1092, x_1093, x_1094, x_1095, x_1096, x_1097, x_1098, x_1099, x_1100, x_1101, x_1102, x_1103, x_1104, x_1105, x_1106, x_1107, x_1108, x_1109, x_1110, x_1111, x_1112, x_1113, x_1114, x_1115, x_1116, x_1117, x_1118, x_1119, x_1120, x_1121, x_1122, x_1123, x_1124, x_1125, x_1126, x_1127, x_1128, x_1129, x_1130, x_1131, x_1132, x_1133, x_1134, x_1135, x_1136, x_1137, x_1138, x_1139, x_1140, x_1141, x_1142, x_1143, x_1144, x_1145, x_1146, x_1147, x_1148, x_1149, x_1150, x_1151, x_1152, x_1153, x_1154, x_1155, x_1156, x_1157, x_1158, x_1159, x_1160, x_1161, x_1162, x_1163, x_1164, x_1165, x_1166, x_1167, x_1168, x_1169, x_1170, x_1171, x_1172, x_1173, x_1174, x_1175, x_1176, x_1177, x_1178, x_1179, x_1180, x_1181, x_1182, x_1183, x_1184, x_1185, x_1186, x_1187, x_1188, x_1189, x_1190, x_1191, x_1192, x_1193, x_1194, x_1195, x_1196, x_1197, x_1198, x_1199, x_1200, x_1201, x_1202, x_1203, x_1204, x_1205, x_1206, x_1207, x_1208, x_1209, x_1210, x_1211, x_1212, x_1213, x_1214, x_1215, x_1216, x_1217, x_1218, x_1219, x_1220, x_1221, x_1222, x_1223, x_1224, x_1225, x_1226, x_1227, x_1228, x_1229, x_1230, x_1231, x_1232, x_1233, x_1234, x_1235, x_1236, x_1237, x_1238, x_1239, x_1240, x_1241, x_1242, x_1243, x_1244, x_1245, x_1246, x_1247, x_1248, x_1249, x_1250, x_1251, x_1252, x_1253, x_1254, x_1255, x_1256, x_1257, x_1258, x_1259, x_1260, x_1261, x_1262, x_1263, x_1264, x_1265, x_1266, x_1267, x_1268, x_1269, x_1270, x_1271, x_1272, x_1273, x_1274, x_1275, x_1276, x_1277, x_1278, x_1279, x_1280, x_1281, x_1282, x_1283, x_1284, x_1285, x_1286, x_1287, x_1288, x_1289, x_1290, x_1291, x_1292, x_1293, x_1294, x_1295, x_1296, x_1297, x_1298, x_1299, x_1300, x_1301, x_1302, x_1303, x_1304, x_1305, x_1306, x_1307, x_1308, x_1309, x_1310, x_1311, x_1312, x_1313, x_1314, x_1315, x_1316, x_1317, x_1318, x_1319, x_1320, x_1321, x_1322, x_1323, x_1324, x_1325, x_1326, x_1327, x_1328, x_1329, x_1330, x_1331, x_1332, x_1333, x_1334, x_1335, x_1336, x_1337, x_1338, x_1339, x_1340, x_1341, x_1342, x_1343, x_1344, x_1345, x_1346, x_1347, x_1348, x_1349, x_1350, x_1351, x_1352, x_1353, x_1354, x_1355, x_1356, x_1357, x_1358, x_1359, x_1360, x_1361, x_1362, x_1363, x_1364, x_1365, x_1366, x_1367, x_1368, x_1369, x_1370, x_1371, x_1372, x_1373, x_1374, x_1375, x_1376, x_1377, x_1378, x_1379, x_1380, x_1381, x_1382, x_1383, x_1384, x_1385, x_1386, x_1387, x_1388, x_1389, x_1390, x_1391, x_1392, x_1393, x_1394, x_1395, x_1396, x_1397, x_1398, x_1399, x_1400, x_1401, x_1402, x_1403, x_1404, x_1405, x_1406, x_1407, x_1408, x_1409, x_1410, x_1411, x_1412, x_1413, x_1414, x_1415, x_1416, x_1417, x_1418, x_1419, x_1420, x_1421, x_1422, x_1423, x_1424, x_1425, x_1426, x_1427, x_1428, x_1429, x_1430, x_1431, x_1432, x_1433, x_1434, x_1435, x_1436, x_1437, x_1438, x_1439, x_1440, x_1441, x_1442, x_1443, x_1444, x_1445, x_1446, x_1447, x_1448, x_1449, x_1450, x_1451, x_1452, x_1453, x_1454, x_1455, x_1456, x_1457, x_1458, x_1459, x_1460, x_1461, x_1462, x_1463, x_1464, x_1465, x_1466, x_1467, x_1468, x_1469, x_1470, x_1471, x_1472, x_1473, x_1474, x_1475, x_1476, x_1477, x_1478, x_1479, x_1480, x_1481, x_1482, x_1483, x_1484, x_1485, x_1486, x_1487, x_1488, x_1489, x_1490, x_1491, x_1492, x_1493, x_1494, x_1495, x_1496, x_1497, x_1498, x_1499, x_1500, x_1501, x_1502, x_1503, x_1504, x_1505, x_1506, x_1507, x_1508, x_1509, x_1510, x_1511, x_1512, x_1513, x_1514, x_1515, x_1516, x_1517, x_1518, x_1519, x_1520, x_1521, x_1522, x_1523, x_1524, x_1525, x_1526, x_1527, x_1528, x_1529, x_1530, x_1531, x_1532, x_1533, x_1534, x_1535, x_1536, x_1537, x_1538, x_1539, x_1540, x_1541, x_1542, x_1543, x_1544, x_1545, x_1546, x_1547, x_1548, x_1549, x_1550, x_1551, x_1552, x_1553, x_1554, x_1555, x_1556, x_1557, x_1558, x_1559, x_1560, x_1561, x_1562, x_1563, x_1564, x_1565, x_1566, x_1567, x_1568, x_1569, x_1570, x_1571, x_1572, x_1573, x_1574, x_1575, x_1576, x_1577, x_1578, x_1579, x_1580, x_1581, x_1582, x_1583, x_1584, x_1585, x_1586, x_1587, x_1588, x_1589, x_1590, x_1591, x_1592, x_1593, x_1594, x_1595, x_1596, x_1597, x_1598, x_1599, x_1600, x_1601, x_1602, x_1603, x_1604, x_1605, x_1606, x_1607, x_1608, x_1609, x_1610, x_1611, x_1612, x_1613, x_1614, x_1615, x_1616, x_1617, x_1618, x_1619, x_1620, x_1621, x_1622, x_1623, x_1624, x_1625, x_1626, x_1627, x_1628, x_1629, x_1630, x_1631, x_1632, x_1633, x_1634, x_1635, x_1636, x_1637, x_1638, x_1639, x_1640, x_1641, x_1642, x_1643, x_1644, x_1645, x_1646, x_1647, x_1648, x_1649, x_1650, x_1651, x_1652, x_1653, x_1654, x_1655, x_1656, x_1657, x_1658, x_1659, x_1660, x_1661, x_1662, x_1663, x_1664, x_1665, x_1666, x_1667, x_1668, x_1669, x_1670, x_1671, x_1672, x_1673, x_1674, x_1675, x_1676, x_1677, x_1678, x_1679, x_1680, x_1681, x_1682, x_1683, x_1684, x_1685, x_1686, x_1687, x_1688, x_1689, x_1690, x_1691, x_1692, x_1693, x_1694, x_1695, x_1696, x_1697, x_1698, x_1699, x_1700, x_1701, x_1702, x_1703, x_1704, x_1705, x_1706, x_1707, x_1708, x_1709, x_1710, x_1711, x_1712, x_1713, x_1714, x_1715, x_1716, x_1717, x_1718, x_1719, x_1720, x_1721, x_1722, x_1723, x_1724, x_1725, x_1726, x_1727, x_1728, x_1729, x_1730, x_1731, x_1732, x_1733, x_1734, x_1735, x_1736, x_1737, x_1738, x_1739, x_1740, x_1741, x_1742, x_1743, x_1744, x_1745, x_1746, x_1747, x_1748, x_1749, x_1750, x_1751, x_1752, x_1753, x_1754, x_1755, x_1756, x_1757, x_1758, x_1759, x_1760, x_1761, x_1762, x_1763, x_1764, x_1765, x_1766, x_1767, x_1768, x_1769, x_1770, x_1771, x_1772, x_1773, x_1774, x_1775, x_1776, x_1777, x_1778, x_1779, x_1780, x_1781, x_1782, x_1783, x_1784, x_1785, x_1786, x_1787, x_1788, x_1789, x_1790, x_1791, x_1792, x_1793, x_1794, x_1795, x_1796, x_1797, x_1798, x_1799, x_1800, x_1801, x_1802, x_1803, x_1804, x_1805, x_1806, x_1807, x_1808, x_1809, x_1810, x_1811, x_1812, x_1813, x_1814, x_1815, x_1816, x_1817, x_1818, x_1819, x_1820, x_1821, x_1822, x_1823, x_1824, x_1825, x_1826, x_1827, x_1828, x_1829, x_1830, x_1831, x_1832, x_1833, x_1834, x_1835, x_1836, x_1837, x_1838, x_1839, x_1840, x_1841, x_1842, x_1843, x_1844, x_1845, x_1846, x_1847, x_1848, x_1849, x_1850, x_1851, x_1852, x_1853, x_1854, x_1855, x_1856, x_1857, x_1858, x_1859, x_1860, x_1861, x_1862, x_1863, x_1864, x_1865, x_1866, x_1867, x_1868, x_1869, x_1870, x_1871, x_1872, x_1873, x_1874, x_1875, x_1876, x_1877, x_1878, x_1879, x_1880, x_1881, x_1882, x_1883, x_1884, x_1885, x_1886, x_1887, x_1888, x_1889, x_1890, x_1891, x_1892, x_1893, x_1894, x_1895, x_1896, x_1897, x_1898, x_1899, x_1900, x_1901, x_1902, x_1903, x_1904, x_1905, x_1906, x_1907, x_1908, x_1909, x_1910, x_1911, x_1912, x_1913, x_1914, x_1915, x_1916, x_1917, x_1918, x_1919, x_1920, x_1921, x_1922, x_1923, x_1924, x_1925, x_1926, x_1927, x_1928, x_1929, x_1930, x_1931, x_1932, x_1933, x_1934, x_1935, x_1936, x_1937, x_1938, x_1939, x_1940, x_1941, x_1942, x_1943, x_1944, x_1945, x_1946, x_1947, x_1948, x_1949, x_1950, x_1951, x_1952, x_1953, x_1954, x_1955, x_1956, x_1957, x_1958, x_1959, x_1960, x_1961, x_1962, x_1963, x_1964, x_1965, x_1966, x_1967, x_1968, x_1969, x_1970, x_1971, x_1972, x_1973, x_1974, x_1975, x_1976, x_1977, x_1978, x_1979, x_1980, x_1981, x_1982, x_1983, x_1984, x_1985, x_1986, x_1987, x_1988, x_1989, x_1990, x_1991, x_1992, x_1993, x_1994, x_1995, x_1996, x_1997, x_1998, x_1999, x_2000, x_2001, x_2002, x_2003, x_2004, x_2005, x_2006, x_2007, x_2008, x_2009, x_2010, x_2011, x_2012, x_2013, x_2014, x_2015, x_2016, x_2017, x_2018, x_2019, x_2020, x_2021, x_2022, x_2023, x_2024, x_2025, x_2026, x_2027, x_2028, x_2029, x_2030, x_2031, x_2032, x_2033, x_2034, x_2035, x_2036, x_2037, x_2038, x_2039, x_2040, x_2041, x_2042, x_2043, x_2044, x_2045, x_2046, x_2047, x_2048, x_2049, x_2050, x_2051, x_2052, x_2053, x_2054, x_2055, x_2056, x_2057, x_2058, x_2059, x_2060, x_2061, x_2062, x_2063, x_2064, x_2065, x_2066, x_2067, x_2068, x_2069, x_2070, x_2071, x_2072, x_2073, x_2074, x_2075, x_2076, x_2077, x_2078, x_2079, x_2080, x_2081, x_2082, x_2083, x_2084, x_2085, x_2086, x_2087, x_2088, x_2089, x_2090, x_2091, x_2092, x_2093, x_2094, x_2095, x_2096, x_2097, x_2098, x_2099, x_2100, x_2101, x_2102, x_2103, x_2104, x_2105, x_2106, x_2107, x_2108, x_2109, x_2110, x_2111, x_2112, x_2113, x_2114, x_2115, x_2116, x_2117, x_2118, x_2119, x_2120, x_2121, x_2122, x_2123, x_2124, x_2125, x_2126, x_2127, x_2128, x_2129, x_2130, x_2131, x_2132, x_2133, x_2134, x_2135, x_2136, x_2137, x_2138, x_2139, x_2140, x_2141, x_2142, x_2143, x_2144, x_2145, x_2146, x_2147, x_2148, x_2149, x_2150, x_2151, x_2152, x_2153, x_2154, x_2155, x_2156, x_2157, x_2158, x_2159, x_2160, x_2161, x_2162, x_2163, x_2164, x_2165, x_2166, x_2167, x_2168, x_2169, x_2170, x_2171, x_2172, x_2173, x_2174, x_2175, x_2176, x_2177, x_2178, x_2179, x_2180, x_2181, x_2182, x_2183, x_2184, x_2185, x_2186, x_2187, x_2188, x_2189, x_2190, x_2191, x_2192, x_2193, x_2194, x_2195, x_2196, x_2197, x_2198, x_2199, x_2200, x_2201, x_2202, x_2203, x_2204, x_2205, x_2206, x_2207, x_2208, x_2209, x_2210, x_2211, x_2212, x_2213, x_2214, x_2215, x_2216, x_2217, x_2218, x_2219, x_2220, x_2221, x_2222, x_2223, x_2224, x_2225, x_2226, x_2227, x_2228, x_2229, x_2230, x_2231, x_2232, x_2233, x_2234, x_2235, x_2236, x_2237, x_2238, x_2239, x_2240, x_2241, x_2242, x_2243, x_2244, x_2245, x_2246, x_2247, x_2248, x_2249, x_2250, x_2251, x_2252, x_2253, x_2254, x_2255, x_2256, x_2257, x_2258, x_2259, x_2260, x_2261, x_2262, x_2263, x_2264, x_2265, x_2266, x_2267, x_2268, x_2269, x_2270, x_2271, x_2272, x_2273, x_2274, x_2275, x_2276, x_2277, x_2278, x_2279, x_2280, x_2281, x_2282, x_2283, x_2284, x_2285, x_2286, x_2287, x_2288, x_2289, x_2290, x_2291, x_2292, x_2293, x_2294, x_2295, x_2296, x_2297, x_2298, x_2299, x_2300, x_2301, x_2302, x_2303, x_2304, x_2305, x_2306, x_2307, x_2308, x_2309, x_2310, x_2311, x_2312, x_2313, x_2314, x_2315, x_2316, x_2317, x_2318, x_2319, x_2320, x_2321, x_2322, x_2323, x_2324, x_2325, x_2326, x_2327, x_2328, x_2329, x_2330, x_2331, x_2332, x_2333, x_2334, x_2335, x_2336, x_2337, x_2338, x_2339, x_2340, x_2341, x_2342, x_2343, x_2344, x_2345, x_2346, x_2347, x_2348, x_2349, x_2350, x_2351, x_2352, x_2353, x_2354, x_2355, x_2356, x_2357, x_2358, x_2359, x_2360, x_2361, x_2362, x_2363, x_2364, x_2365, x_2366, x_2367, x_2368, x_2369, x_2370, x_2371, x_2372, x_2373, x_2374, x_2375, x_2376, x_2377, x_2378, x_2379, x_2380, x_2381, x_2382, x_2383, x_2384, x_2385, x_2386, x_2387, x_2388, x_2389, x_2390, x_2391, x_2392, x_2393, x_2394, x_2395, x_2396, x_2397, x_2398, x_2399, x_2400, x_2401, x_2402, x_2403, x_2404, x_2405, x_2406, x_2407, x_2408, x_2409, x_2410, x_2411, x_2412, x_2413, x_2414, x_2415, x_2416, x_2417, x_2418, x_2419, x_2420, x_2421, x_2422, x_2423, x_2424, x_2425, x_2426, x_2427, x_2428, x_2429, x_2430, x_2431, x_2432, x_2433, x_2434, x_2435, x_2436, x_2437, x_2438, x_2439, x_2440, x_2441, x_2442, x_2443, x_2444, x_2445, x_2446, x_2447, x_2448, x_2449, x_2450, x_2451, x_2452, x_2453, x_2454, x_2455, x_2456, x_2457, x_2458, x_2459, x_2460, x_2461, x_2462, x_2463, x_2464, x_2465, x_2466, x_2467, x_2468, x_2469, x_2470, x_2471, x_2472, x_2473, x_2474, x_2475, x_2476, x_2477, x_2478, x_2479, x_2480, x_2481, x_2482, x_2483, x_2484, x_2485, x_2486, x_2487, x_2488, x_2489, x_2490, x_2491, x_2492, x_2493, x_2494, x_2495, x_2496, x_2497, x_2498, x_2499, x_2500, x_2501, x_2502, x_2503, x_2504, x_2505, x_2506, x_2507, x_2508, x_2509, x_2510, x_2511, x_2512, x_2513, x_2514, x_2515, x_2516, x_2517, x_2518, x_2519, x_2520, x_2521, x_2522, x_2523, x_2524, x_2525, x_2526, x_2527, x_2528, x_2529, x_2530, x_2531, x_2532, x_2533, x_2534, x_2535, x_2536, x_2537, x_2538, x_2539, x_2540, x_2541, x_2542, x_2543, x_2544, x_2545, x_2546, x_2547, x_2548, x_2549, x_2550, x_2551, x_2552, x_2553, x_2554, x_2555, x_2556, x_2557, x_2558, x_2559, x_2560, x_2561, x_2562, x_2563, x_2564, x_2565, x_2566, x_2567, x_2568, x_2569, x_2570, x_2571, x_2572, x_2573, x_2574, x_2575, x_2576, x_2577, x_2578, x_2579, x_2580, x_2581, x_2582, x_2583, x_2584, x_2585, x_2586, x_2587, x_2588, x_2589, x_2590, x_2591, x_2592, x_2593, x_2594, x_2595, x_2596, x_2597, x_2598, x_2599, x_2600, x_2601, x_2602, x_2603, x_2604, x_2605, x_2606, x_2607, x_2608, x_2609, x_2610, x_2611, x_2612, x_2613, x_2614, x_2615, x_2616, x_2617, x_2618, x_2619, x_2620, x_2621, x_2622, x_2623, x_2624, x_2625, x_2626, x_2627, x_2628, x_2629, x_2630, x_2631, x_2632, x_2633, x_2634, x_2635, x_2636, x_2637, x_2638, x_2639, x_2640, x_2641, x_2642, x_2643, x_2644, x_2645, x_2646, x_2647, x_2648, x_2649, x_2650, x_2651, x_2652, x_2653, x_2654, x_2655, x_2656, x_2657, x_2658, x_2659, x_2660, x_2661, x_2662, x_2663, x_2664, x_2665, x_2666, x_2667, x_2668, x_2669, x_2670, x_2671, x_2672, x_2673, x_2674, x_2675, x_2676, x_2677, x_2678, x_2679, x_2680, x_2681, x_2682, x_2683, x_2684, x_2685, x_2686, x_2687, x_2688, x_2689, x_2690, x_2691, x_2692, x_2693, x_2694, x_2695, x_2696, x_2697, x_2698, x_2699, x_2700, x_2701, x_2702, x_2703, x_2704, x_2705, x_2706, x_2707, x_2708, x_2709, x_2710, x_2711, x_2712, x_2713, x_2714, x_2715, x_2716, x_2717, x_2718, x_2719, x_2720, x_2721, x_2722, x_2723, x_2724, x_2725, x_2726, x_2727, x_2728, x_2729, x_2730, x_2731, x_2732, x_2733, x_2734, x_2735, x_2736, x_2737, x_2738, x_2739, x_2740, x_2741, x_2742, x_2743, x_2744, x_2745, x_2746, x_2747, x_2748, x_2749, x_2750, x_2751, x_2752, x_2753, x_2754, x_2755, x_2756, x_2757, x_2758, x_2759, x_2760, x_2761, x_2762, x_2763, x_2764, x_2765, x_2766, x_2767, x_2768, x_2769, x_2770, x_2771, x_2772, x_2773, x_2774, x_2775, x_2776, x_2777, x_2778, x_2779, x_2780, x_2781, x_2782, x_2783, x_2784, x_2785, x_2786, x_2787, x_2788, x_2789, x_2790, x_2791, x_2792, x_2793, x_2794, x_2795, x_2796, x_2797, x_2798, x_2799, x_2800, x_2801, x_2802, x_2803, x_2804, x_2805, x_2806, x_2807, x_2808, x_2809, x_2810, x_2811, x_2812, x_2813, x_2814, x_2815, x_2816, x_2817, x_2818, x_2819, x_2820, x_2821, x_2822, x_2823, x_2824, x_2825, x_2826, x_2827, x_2828, x_2829, x_2830, x_2831, x_2832, x_2833, x_2834, x_2835, x_2836, x_2837, x_2838, x_2839, x_2840, x_2841, x_2842, x_2843, x_2844, x_2845, x_2846, x_2847, x_2848, x_2849, x_2850, x_2851, x_2852, x_2853, x_2854, x_2855, x_2856, x_2857, x_2858, x_2859, x_2860, x_2861, x_2862, x_2863, x_2864, x_2865, x_2866, x_2867, x_2868, x_2869, x_2870, x_2871, x_2872, x_2873, x_2874, x_2875, x_2876, x_2877, x_2878, x_2879, x_2880, x_2881, x_2882, x_2883, x_2884, x_2885, x_2886, x_2887, x_2888, x_2889, x_2890, x_2891, x_2892, x_2893, x_2894, x_2895, x_2896, x_2897, x_2898, x_2899, x_2900, x_2901, x_2902, x_2903, x_2904, x_2905, x_2906, x_2907, x_2908, x_2909, x_2910, x_2911, x_2912, x_2913, x_2914, x_2915, x_2916, x_2917, x_2918, x_2919, x_2920, x_2921, x_2922, x_2923, x_2924, x_2925, x_2926, x_2927, x_2928, x_2929, x_2930, x_2931, x_2932, x_2933, x_2934, x_2935, x_2936, x_2937, x_2938, x_2939, x_2940, x_2941, x_2942, x_2943, x_2944, x_2945, x_2946, x_2947, x_2948, x_2949, x_2950, x_2951, x_2952, x_2953, x_2954, x_2955, x_2956, x_2957, x_2958, x_2959, x_2960, x_2961, x_2962, x_2963, x_2964, x_2965, x_2966, x_2967, x_2968, x_2969, x_2970, x_2971, x_2972, x_2973, x_2974, x_2975, x_2976, x_2977, x_2978, x_2979, x_2980, x_2981, x_2982, x_2983, x_2984, x_2985, x_2986, x_2987, x_2988, x_2989, x_2990, x_2991, x_2992, x_2993, x_2994, x_2995, x_2996, x_2997, x_2998, x_2999, x_3000, x_3001, x_3002, x_3003, x_3004, x_3005, x_3006, x_3007, x_3008, x_3009, x_3010, x_3011, x_3012, x_3013, x_3014, x_3015, x_3016, x_3017, x_3018, x_3019, x_3020, x_3021, x_3022, x_3023, x_3024, x_3025, x_3026, x_3027, x_3028, x_3029, x_3030, x_3031, x_3032, x_3033, x_3034, x_3035, x_3036, x_3037, x_3038, x_3039, x_3040, x_3041, x_3042, x_3043, x_3044, x_3045, x_3046, x_3047, x_3048, x_3049, x_3050, x_3051, x_3052, x_3053, x_3054, x_3055, x_3056, x_3057, x_3058, x_3059, x_3060, x_3061, x_3062, x_3063, x_3064, x_3065, x_3066, x_3067, x_3068, x_3069, x_3070, x_3071, x_3072, x_3073, x_3074, x_3075, x_3076, x_3077, x_3078, x_3079, x_3080, x_3081, x_3082, x_3083, x_3084, x_3085, x_3086, x_3087, x_3088, x_3089, x_3090, x_3091, x_3092, x_3093, x_3094, x_3095, x_3096, x_3097, x_3098, x_3099, x_3100, x_3101, x_3102, x_3103, x_3104, x_3105, x_3106, x_3107, x_3108, x_3109, x_3110, x_3111, x_3112, x_3113, x_3114, x_3115, x_3116, x_3117, x_3118, x_3119, x_3120, x_3121, x_3122, x_3123, x_3124, x_3125, x_3126, x_3127, x_3128, x_3129, x_3130, x_3131, x_3132, x_3133, x_3134, x_3135, x_3136, x_3137, x_3138, x_3139, x_3140, x_3141, x_3142, x_3143, x_3144, x_3145, x_3146, x_3147, x_3148, x_3149, x_3150, x_3151, x_3152, x_3153, x_3154, x_3155, x_3156, x_3157, x_3158, x_3159, x_3160, x_3161, x_3162, x_3163, x_3164, x_3165, x_3166, x_3167, x_3168, x_3169, x_3170, x_3171, x_3172, x_3173, x_3174, x_3175, x_3176, x_3177, x_3178, x_3179, x_3180, x_3181, x_3182, x_3183, x_3184, x_3185, x_3186, x_3187, x_3188, x_3189, x_3190, x_3191, x_3192, x_3193, x_3194, x_3195, x_3196, x_3197, x_3198, x_3199, x_3200, x_3201, x_3202, x_3203, x_3204, x_3205, x_3206, x_3207, x_3208, x_3209, x_3210, x_3211, x_3212, x_3213, x_3214, x_3215, x_3216, x_3217, x_3218, x_3219, x_3220, x_3221, x_3222, x_3223, x_3224, x_3225, x_3226, x_3227, x_3228, x_3229, x_3230, x_3231, x_3232, x_3233, x_3234, x_3235, x_3236, x_3237, x_3238, x_3239, x_3240, x_3241, x_3242, x_3243, x_3244, x_3245, x_3246, x_3247, x_3248, x_3249, x_3250, x_3251, x_3252, x_3253, x_3254, x_3255, x_3256, x_3257, x_3258, x_3259, x_3260, x_3261, x_3262, x_3263, x_3264, x_3265, x_3266, x_3267, x_3268, x_3269, x_3270, x_3271, x_3272, x_3273, x_3274, x_3275, x_3276, x_3277, x_3278, x_3279, x_3280, x_3281, x_3282, x_3283, x_3284, x_3285, x_3286, x_3287, x_3288, x_3289, x_3290, x_3291, x_3292, x_3293, x_3294, x_3295, x_3296, x_3297, x_3298, x_3299, x_3300, x_3301, x_3302, x_3303, x_3304, x_3305, x_3306, x_3307, x_3308, x_3309, x_3310, x_3311, x_3312, x_3313, x_3314, x_3315, x_3316, x_3317, x_3318, x_3319, x_3320, x_3321, x_3322, x_3323, x_3324, x_3325, x_3326, x_3327, x_3328, x_3329, x_3330, x_3331, x_3332, x_3333, x_3334, x_3335, x_3336, x_3337, x_3338, x_3339, x_3340, x_3341, x_3342, x_3343, x_3344, x_3345, x_3346, x_3347, x_3348, x_3349, x_3350, x_3351, x_3352, x_3353, x_3354, x_3355, x_3356, x_3357, x_3358, x_3359, x_3360, x_3361, x_3362, x_3363, x_3364, x_3365, x_3366, x_3367, x_3368, x_3369, x_3370, x_3371, x_3372, x_3373, x_3374, x_3375, x_3376, x_3377, x_3378, x_3379, x_3380, x_3381, x_3382, x_3383, x_3384, x_3385, x_3386, x_3387, x_3388, x_3389, x_3390, x_3391, x_3392, x_3393, x_3394, x_3395, x_3396, x_3397, x_3398, x_3399, x_3400, x_3401, x_3402, x_3403, x_3404, x_3405, x_3406, x_3407, x_3408, x_3409, x_3410, x_3411, x_3412, x_3413, x_3414, x_3415, x_3416, x_3417, x_3418, x_3419, x_3420, x_3421, x_3422, x_3423, x_3424, x_3425, x_3426, x_3427, x_3428, x_3429, x_3430, x_3431, x_3432, x_3433, x_3434, x_3435, x_3436, x_3437, x_3438, x_3439, x_3440, x_3441, x_3442, x_3443, x_3444, x_3445, x_3446, x_3447, x_3448, x_3449, x_3450, x_3451, x_3452, x_3453, x_3454, x_3455, x_3456, x_3457, x_3458, x_3459, x_3460, x_3461, x_3462, x_3463, x_3464, x_3465, x_3466, x_3467, x_3468, x_3469, x_3470, x_3471, x_3472, x_3473, x_3474, x_3475, x_3476, x_3477, x_3478, x_3479, x_3480, x_3481, x_3482, x_3483, x_3484, x_3485, x_3486, x_3487, x_3488, x_3489, x_3490, x_3491, x_3492, x_3493, x_3494, x_3495, x_3496, x_3497, x_3498, x_3499, x_3500, x_3501, x_3502, x_3503, x_3504, x_3505, x_3506, x_3507, x_3508, x_3509, x_3510, x_3511, x_3512, x_3513, x_3514, x_3515, x_3516, x_3517, x_3518, x_3519, x_3520, x_3521, x_3522, x_3523, x_3524, x_3525, x_3526, x_3527, x_3528, x_3529, x_3530, x_3531, x_3532, x_3533, x_3534, x_3535, x_3536, x_3537, x_3538, x_3539, x_3540, x_3541, x_3542, x_3543, x_3544, x_3545, x_3546, x_3547, x_3548, x_3549, x_3550, x_3551, x_3552, x_3553, x_3554, x_3555, x_3556, x_3557, x_3558, x_3559, x_3560, x_3561, x_3562, x_3563, x_3564, x_3565, x_3566, x_3567, x_3568, x_3569, x_3570, x_3571, x_3572, x_3573, x_3574, x_3575, x_3576, x_3577, x_3578, x_3579, x_3580, x_3581, x_3582, x_3583, x_3584, x_3585, x_3586, x_3587, x_3588, x_3589, x_3590, x_3591, x_3592, x_3593, x_3594, x_3595, x_3596, x_3597, x_3598, x_3599, x_3600, x_3601, x_3602, x_3603, x_3604, x_3605, x_3606, x_3607, x_3608, x_3609, x_3610, x_3611, x_3612, x_3613, x_3614, x_3615, x_3616, x_3617, x_3618, x_3619, x_3620, x_3621, x_3622, x_3623, x_3624, x_3625, x_3626, x_3627, x_3628, x_3629, x_3630, x_3631, x_3632, x_3633, x_3634, x_3635, x_3636, x_3637, x_3638, x_3639, x_3640, x_3641, x_3642, x_3643, x_3644, x_3645, x_3646, x_3647, x_3648, x_3649, x_3650, x_3651, x_3652, x_3653, x_3654, x_3655, x_3656, x_3657, x_3658, x_3659, x_3660, x_3661, x_3662, x_3663, x_3664, x_3665, x_3666, x_3667, x_3668, x_3669, x_3670, x_3671, x_3672, x_3673, x_3674, x_3675, x_3676, x_3677, x_3678, x_3679, x_3680, x_3681, x_3682, x_3683, x_3684, x_3685, x_3686, x_3687, x_3688, x_3689, x_3690, x_3691, x_3692, x_3693, x_3694, x_3695, x_3696, x_3697, x_3698, x_3699, x_3700, x_3701, x_3702, x_3703, x_3704, x_3705, x_3706, x_3707, x_3708, x_3709, x_3710, x_3711, x_3712, x_3713, x_3714, x_3715, x_3716, x_3717, x_3718, x_3719, x_3720, x_3721, x_3722, x_3723, x_3724, x_3725, x_3726, x_3727, x_3728, x_3729, x_3730, x_3731, x_3732, x_3733, x_3734, x_3735, x_3736, x_3737, x_3738, x_3739, x_3740, x_3741, x_3742, x_3743, x_3744, x_3745, x_3746, x_3747, x_3748, x_3749, x_3750, x_3751, x_3752, x_3753, x_3754, x_3755, x_3756, x_3757, x_3758, x_3759, x_3760, x_3761, x_3762, x_3763, x_3764, x_3765, x_3766, x_3767, x_3768, x_3769, x_3770, x_3771, x_3772, x_3773, x_3774, x_3775, x_3776, x_3777, x_3778, x_3779, x_3780, x_3781, x_3782, x_3783, x_3784, x_3785, x_3786, x_3787, x_3788, x_3789, x_3790, x_3791, x_3792, x_3793, x_3794, x_3795, x_3796, x_3797, x_3798, x_3799, x_3800, x_3801, x_3802, x_3803, x_3804, x_3805, x_3806, x_3807, x_3808, x_3809, x_3810, x_3811, x_3812, x_3813, x_3814, x_3815, x_3816, x_3817, x_3818, x_3819, x_3820, x_3821, x_3822, x_3823, x_3824, x_3825, x_3826, x_3827, x_3828, x_3829, x_3830, x_3831, x_3832, x_3833, x_3834, x_3835, x_3836, x_3837, x_3838, x_3839, x_3840, x_3841, x_3842, x_3843, x_3844, x_3845, x_3846, x_3847, x_3848, x_3849, x_3850, x_3851, x_3852, x_3853, x_3854, x_3855, x_3856, x_3857, x_3858, x_3859, x_3860, x_3861, x_3862, x_3863, x_3864, x_3865, x_3866, x_3867, x_3868, x_3869, x_3870, x_3871, x_3872, x_3873, x_3874, x_3875, x_3876, x_3877, x_3878, x_3879, x_3880, x_3881, x_3882, x_3883, x_3884, x_3885, x_3886, x_3887, x_3888, x_3889, x_3890, x_3891, x_3892, x_3893, x_3894, x_3895, x_3896, x_3897, x_3898, x_3899, x_3900, x_3901, x_3902, x_3903, x_3904, x_3905, x_3906, x_3907, x_3908, x_3909, x_3910, x_3911, x_3912, x_3913, x_3914, x_3915, x_3916, x_3917, x_3918, x_3919, x_3920, x_3921, x_3922, x_3923, x_3924, x_3925, x_3926, x_3927, x_3928, x_3929, x_3930, x_3931, x_3932, x_3933, x_3934, x_3935, x_3936, x_3937, x_3938, x_3939, x_3940, x_3941, x_3942, x_3943, x_3944, x_3945, x_3946, x_3947, x_3948, x_3949, x_3950, x_3951, x_3952, x_3953, x_3954, x_3955, x_3956, x_3957, x_3958, x_3959, x_3960, x_3961, x_3962, x_3963, x_3964, x_3965, x_3966, x_3967, x_3968, x_3969, x_3970, x_3971, x_3972, x_3973, x_3974, x_3975, x_3976, x_3977, x_3978, x_3979, x_3980, x_3981, x_3982, x_3983, x_3984, x_3985, x_3986, x_3987, x_3988, x_3989, x_3990, x_3991, x_3992, x_3993, x_3994, x_3995, x_3996, x_3997, x_3998, x_3999, x_4000, x_4001, x_4002, x_4003, x_4004, x_4005, x_4006, x_4007, x_4008, x_4009, x_4010, x_4011, x_4012, x_4013, x_4014, x_4015, x_4016, x_4017, x_4018, x_4019, x_4020, x_4021, x_4022, x_4023, x_4024, x_4025, x_4026, x_4027, x_4028, x_4029, x_4030, x_4031, x_4032, x_4033, x_4034, x_4035, x_4036, x_4037, x_4038, x_4039, x_4040, x_4041, x_4042, x_4043, x_4044, x_4045, x_4046, x_4047, x_4048, x_4049, x_4050, x_4051, x_4052, x_4053, x_4054, x_4055, x_4056, x_4057, x_4058, x_4059, x_4060, x_4061, x_4062, x_4063, x_4064, x_4065, x_4066, x_4067, x_4068, x_4069, x_4070, x_4071, x_4072, x_4073, x_4074, x_4075, x_4076, x_4077, x_4078, x_4079, x_4080, x_4081, x_4082, x_4083, x_4084, x_4085, x_4086, x_4087, x_4088, x_4089, x_4090, x_4091, x_4092, x_4093, x_4094, x_4095, x_4096, x_4097, x_4098, x_4099, x_4100, x_4101, x_4102, x_4103, x_4104, x_4105, x_4106, x_4107, x_4108, x_4109, x_4110, x_4111, x_4112, x_4113, x_4114, x_4115, x_4116, x_4117, x_4118, x_4119, x_4120, x_4121, x_4122, x_4123, x_4124, x_4125, x_4126, x_4127, x_4128, x_4129, x_4130, x_4131, x_4132, x_4133, x_4134, x_4135, x_4136, x_4137, x_4138, x_4139, x_4140, x_4141, x_4142, x_4143, x_4144, x_4145, x_4146, x_4147, x_4148, x_4149, x_4150, x_4151, x_4152, x_4153, x_4154, x_4155, x_4156, x_4157, x_4158, x_4159, x_4160, x_4161, x_4162, x_4163, x_4164, x_4165, x_4166, x_4167, x_4168, x_4169, x_4170, x_4171, x_4172, x_4173, x_4174, x_4175, x_4176, x_4177, x_4178, x_4179, x_4180, x_4181, x_4182, x_4183, x_4184, x_4185, x_4186, x_4187, x_4188, x_4189, x_4190, x_4191, x_4192, x_4193, x_4194, x_4195, x_4196, x_4197, x_4198, x_4199, x_4200, x_4201, x_4202, x_4203, x_4204, x_4205, x_4206, x_4207, x_4208, x_4209, x_4210, x_4211, x_4212, x_4213, x_4214, x_4215, x_4216, x_4217, x_4218, x_4219, x_4220, x_4221, x_4222, x_4223, x_4224, x_4225, x_4226, x_4227, x_4228, x_4229, x_4230, x_4231, x_4232, x_4233, x_4234, x_4235, x_4236, x_4237, x_4238, x_4239, x_4240, x_4241, x_4242, x_4243, x_4244, x_4245, x_4246, x_4247, x_4248, x_4249, x_4250, x_4251, x_4252, x_4253, x_4254, x_4255, x_4256, x_4257, x_4258, x_4259, x_4260, x_4261, x_4262, x_4263, x_4264, x_4265, x_4266, x_4267, x_4268, x_4269, x_4270, x_4271, x_4272, x_4273, x_4274, x_4275, x_4276, x_4277, x_4278, x_4279, x_4280, x_4281, x_4282, x_4283, x_4284, x_4285, x_4286, x_4287, x_4288, x_4289, x_4290, x_4291, x_4292, x_4293, x_4294, x_4295, x_4296, x_4297, x_4298, x_4299, x_4300, x_4301, x_4302, x_4303, x_4304, x_4305, x_4306, x_4307, x_4308, x_4309, x_4310, x_4311, x_4312, x_4313, x_4314, x_4315, x_4316, x_4317, x_4318, x_4319, x_4320, x_4321, x_4322, x_4323, x_4324, x_4325, x_4326, x_4327, x_4328, x_4329, x_4330, x_4331, x_4332, x_4333, x_4334, x_4335, x_4336, x_4337, x_4338, x_4339, x_4340, x_4341, x_4342, x_4343, x_4344, x_4345, x_4346, x_4347, x_4348, x_4349, x_4350, x_4351, x_4352, x_4353, x_4354, x_4355, x_4356, x_4357, x_4358, x_4359, x_4360, x_4361, x_4362, x_4363, x_4364, x_4365, x_4366, x_4367, x_4368, x_4369, x_4370, x_4371, x_4372, x_4373, x_4374, x_4375, x_4376, x_4377, x_4378, x_4379, x_4380, x_4381, x_4382, x_4383, x_4384, x_4385, x_4386, x_4387, x_4388, x_4389, x_4390, x_4391, x_4392, x_4393, x_4394, x_4395, x_4396, x_4397, x_4398, x_4399, x_4400, x_4401, x_4402, x_4403, x_4404, x_4405, x_4406, x_4407, x_4408, x_4409, x_4410, x_4411, x_4412, x_4413, x_4414, x_4415, x_4416, x_4417, x_4418, x_4419, x_4420, x_4421, x_4422, x_4423, x_4424, x_4425, x_4426, x_4427, x_4428, x_4429, x_4430, x_4431, x_4432, x_4433, x_4434, x_4435, x_4436, x_4437, x_4438, x_4439, x_4440, x_4441, x_4442, x_4443, x_4444, x_4445, x_4446, x_4447, x_4448, x_4449, x_4450, x_4451, x_4452, x_4453, x_4454, x_4455, x_4456, x_4457, x_4458, x_4459, x_4460, x_4461, x_4462, x_4463, x_4464, x_4465, x_4466, x_4467, x_4468, x_4469, x_4470, x_4471, x_4472, x_4473, x_4474, x_4475, x_4476, x_4477, x_4478, x_4479, x_4480, x_4481, x_4482, x_4483, x_4484, x_4485, x_4486, x_4487, x_4488, x_4489, x_4490, x_4491, x_4492, x_4493, x_4494, x_4495, x_4496, x_4497, x_4498, x_4499, x_4500, x_4501, x_4502, x_4503, x_4504, x_4505, x_4506, x_4507, x_4508, x_4509, x_4510, x_4511, x_4512, x_4513, x_4514, x_4515, x_4516, x_4517, x_4518, x_4519, x_4520, x_4521, x_4522, x_4523, x_4524, x_4525, x_4526, x_4527, x_4528, x_4529, x_4530, x_4531, x_4532, x_4533, x_4534, x_4535, x_4536, x_4537, x_4538, x_4539, x_4540, x_4541, x_4542, x_4543, x_4544, x_4545, x_4546, x_4547, x_4548, x_4549, x_4550, x_4551, x_4552, x_4553, x_4554, x_4555, x_4556, x_4557, x_4558, x_4559, x_4560, x_4561, x_4562, x_4563, x_4564, x_4565, x_4566, x_4567, x_4568, x_4569, x_4570, x_4571, x_4572, x_4573, x_4574, x_4575, x_4576, x_4577, x_4578, x_4579, x_4580, x_4581, x_4582, x_4583, x_4584, x_4585, x_4586, x_4587, x_4588, x_4589, x_4590, x_4591, x_4592, x_4593, x_4594, x_4595, x_4596, x_4597, x_4598, x_4599, x_4600, x_4601, x_4602, x_4603, x_4604, x_4605, x_4606, x_4607, x_4608, x_4609, x_4610, x_4611, x_4612, x_4613, x_4614, x_4615, x_4616, x_4617, x_4618, x_4619, x_4620, x_4621, x_4622, x_4623, x_4624, x_4625, x_4626, x_4627, x_4628, x_4629, x_4630, x_4631, x_4632, x_4633, x_4634, x_4635, x_4636, x_4637, x_4638, x_4639, x_4640, x_4641, x_4642, x_4643, x_4644, x_4645, x_4646, x_4647, x_4648, x_4649, x_4650, x_4651, x_4652, x_4653, x_4654, x_4655, x_4656, x_4657, x_4658, x_4659, x_4660, x_4661, x_4662, x_4663, x_4664, x_4665, x_4666, x_4667, x_4668, x_4669, x_4670, x_4671, x_4672, x_4673, x_4674, x_4675, x_4676, x_4677, x_4678, x_4679, x_4680, x_4681, x_4682, x_4683, x_4684, x_4685, x_4686, x_4687, x_4688, x_4689, x_4690, x_4691, x_4692, x_4693, x_4694, x_4695, x_4696, x_4697, x_4698, x_4699, x_4700, x_4701, x_4702, x_4703, x_4704, x_4705, x_4706, x_4707, x_4708, x_4709, x_4710, x_4711, x_4712, x_4713, x_4714, x_4715, x_4716, x_4717, x_4718, x_4719, x_4720, x_4721, x_4722, x_4723, x_4724, x_4725, x_4726, x_4727, x_4728, x_4729, x_4730, x_4731, x_4732, x_4733, x_4734, x_4735, x_4736, x_4737, x_4738, x_4739, x_4740, x_4741, x_4742, x_4743, x_4744, x_4745, x_4746, x_4747, x_4748, x_4749, x_4750, x_4751, x_4752, x_4753, x_4754, x_4755, x_4756, x_4757, x_4758, x_4759, x_4760, x_4761, x_4762, x_4763, x_4764, x_4765, x_4766, x_4767, x_4768, x_4769, x_4770, x_4771, x_4772, x_4773, x_4774, x_4775, x_4776, x_4777, x_4778, x_4779, x_4780, x_4781, x_4782, x_4783, x_4784, x_4785, x_4786, x_4787, x_4788, x_4789, x_4790, x_4791, x_4792, x_4793, x_4794, x_4795, x_4796, x_4797, x_4798, x_4799, x_4800, x_4801, x_4802, x_4803, x_4804, x_4805, x_4806, x_4807, x_4808, x_4809, x_4810, x_4811, x_4812, x_4813, x_4814, x_4815, x_4816, x_4817, x_4818, x_4819, x_4820, x_4821, x_4822, x_4823, x_4824, x_4825, x_4826, x_4827, x_4828, x_4829, x_4830, x_4831, x_4832, x_4833, x_4834, x_4835, x_4836, x_4837, x_4838, x_4839, x_4840, x_4841, x_4842, x_4843, x_4844, x_4845, x_4846, x_4847, x_4848, x_4849, x_4850, x_4851, x_4852, x_4853, x_4854, x_4855, x_4856, x_4857, x_4858, x_4859, x_4860, x_4861, x_4862, x_4863, x_4864, x_4865, x_4866, x_4867, x_4868, x_4869, x_4870, x_4871, x_4872, x_4873, x_4874, x_4875, x_4876, x_4877, x_4878, x_4879, x_4880, x_4881, x_4882, x_4883, x_4884, x_4885, x_4886, x_4887, x_4888, x_4889, x_4890, x_4891, x_4892, x_4893, x_4894, x_4895, x_4896, x_4897, x_4898, x_4899, x_4900, x_4901, x_4902, x_4903, x_4904, x_4905, x_4906, x_4907, x_4908, x_4909, x_4910, x_4911, x_4912, x_4913, x_4914, x_4915, x_4916, x_4917, x_4918, x_4919, x_4920, x_4921, x_4922, x_4923, x_4924, x_4925, x_4926, x_4927, x_4928, x_4929, x_4930, x_4931, x_4932, x_4933, x_4934, x_4935, x_4936, x_4937, x_4938, x_4939, x_4940, x_4941, x_4942, x_4943, x_4944, x_4945, x_4946, x_4947, x_4948, x_4949, x_4950, x_4951, x_4952, x_4953, x_4954, x_4955, x_4956, x_4957, x_4958, x_4959, x_4960, x_4961, x_4962, x_4963, x_4964, x_4965, x_4966, x_4967, x_4968, x_4969, x_4970, x_4971, x_4972, x_4973, x_4974, x_4975, x_4976, x_4977, x_4978, x_4979, x_4980, x_4981, x_4982, x_4983, x_4984, x_4985, x_4986, x_4987, x_4988, x_4989, x_4990, x_4991, x_4992, x_4993, x_4994, x_4995, x_4996, x_4997, x_4998, x_4999, x_5000, x_5001, x_5002, x_5003, x_5004, x_5005, x_5006, x_5007, x_5008, x_5009, x_5010, x_5011, x_5012, x_5013, x_5014, x_5015, x_5016, x_5017, x_5018, x_5019, x_5020, x_5021, x_5022, x_5023, x_5024, x_5025, x_5026, x_5027, x_5028, x_5029, x_5030, x_5031, x_5032, x_5033, x_5034, x_5035, x_5036, x_5037, x_5038, x_5039, x_5040, x_5041, x_5042, x_5043, x_5044, x_5045, x_5046, x_5047, x_5048, x_5049, x_5050, x_5051, x_5052, x_5053, x_5054, x_5055, x_5056, x_5057, x_5058, x_5059, x_5060, x_5061, x_5062, x_5063, x_5064, x_5065, x_5066, x_5067, x_5068, x_5069, x_5070, x_5071, x_5072, x_5073, x_5074, x_5075, x_5076, x_5077, x_5078, x_5079, x_5080, x_5081, x_5082, x_5083, x_5084, x_5085, x_5086, x_5087, x_5088, x_5089, x_5090, x_5091, x_5092, x_5093, x_5094, x_5095, x_5096, x_5097, x_5098, x_5099, x_5100, x_5101, x_5102, x_5103, x_5104, x_5105, x_5106, x_5107, x_5108, x_5109, x_5110, x_5111, x_5112, x_5113, x_5114, x_5115, x_5116, x_5117, x_5118, x_5119, x_5120, x_5121, x_5122, x_5123, x_5124, x_5125, x_5126, x_5127, x_5128, x_5129, x_5130, x_5131, x_5132, x_5133, x_5134, x_5135, x_5136, x_5137, x_5138, x_5139, x_5140, x_5141, x_5142, x_5143, x_5144, x_5145, x_5146, x_5147, x_5148, x_5149, x_5150, x_5151, x_5152, x_5153, x_5154, x_5155, x_5156, x_5157, x_5158, x_5159, x_5160, x_5161, x_5162, x_5163, x_5164, x_5165, x_5166, x_5167, x_5168, x_5169, x_5170, x_5171, x_5172, x_5173, x_5174, x_5175, x_5176, x_5177, x_5178, x_5179, x_5180, x_5181, x_5182, x_5183, x_5184, x_5185, x_5186, x_5187, x_5188, x_5189, x_5190, x_5191, x_5192, x_5193, x_5194, x_5195, x_5196, x_5197, x_5198, x_5199, x_5200, x_5201, x_5202, x_5203, x_5204, x_5205, x_5206, x_5207, x_5208, x_5209, x_5210, x_5211, x_5212, x_5213, x_5214, x_5215, x_5216, x_5217, x_5218, x_5219, x_5220, x_5221, x_5222, x_5223, x_5224, x_5225, x_5226, x_5227, x_5228, x_5229, x_5230, x_5231, x_5232, x_5233, x_5234, x_5235, x_5236, x_5237, x_5238, x_5239, x_5240, x_5241, x_5242, x_5243, x_5244, x_5245, x_5246, x_5247, x_5248, x_5249, x_5250, x_5251, x_5252, x_5253, x_5254, x_5255, x_5256, x_5257, x_5258, x_5259, x_5260, x_5261, x_5262, x_5263, x_5264, x_5265, x_5266, x_5267, x_5268, x_5269, x_5270, x_5271, x_5272, x_5273, x_5274, x_5275, x_5276, x_5277, x_5278, x_5279, x_5280, x_5281, x_5282, x_5283, x_5284, x_5285, x_5286, x_5287, x_5288, x_5289, x_5290, x_5291, x_5292, x_5293, x_5294, x_5295, x_5296, x_5297, x_5298, x_5299, x_5300, x_5301, x_5302, x_5303, x_5304, x_5305, x_5306, x_5307, x_5308, x_5309, x_5310, x_5311, x_5312, x_5313, x_5314, x_5315, x_5316, x_5317, x_5318, x_5319, x_5320, x_5321, x_5322, x_5323, x_5324, x_5325, x_5326, x_5327, x_5328, x_5329, x_5330, x_5331, x_5332, x_5333, x_5334, x_5335, x_5336, x_5337, x_5338, x_5339, x_5340, x_5341, x_5342, x_5343, x_5344, x_5345, x_5346, x_5347, x_5348, x_5349, x_5350, x_5351, x_5352, x_5353, x_5354, x_5355, x_5356, x_5357, x_5358, x_5359, x_5360, x_5361, x_5362, x_5363, x_5364, x_5365, x_5366, x_5367, x_5368, x_5369, x_5370, x_5371, x_5372, x_5373, x_5374, x_5375, x_5376, x_5377, x_5378, x_5379, x_5380, x_5381, x_5382, x_5383, x_5384, x_5385, x_5386, x_5387, x_5388, x_5389, x_5390, x_5391, x_5392, x_5393, x_5394, x_5395, x_5396, x_5397, x_5398, x_5399, x_5400, x_5401, x_5402, x_5403, x_5404, x_5405, x_5406, x_5407, x_5408, x_5409, x_5410, x_5411, x_5412, x_5413, x_5414, x_5415, x_5416, x_5417, x_5418, x_5419, x_5420, x_5421, x_5422, x_5423, x_5424, x_5425, x_5426, x_5427, x_5428, x_5429, x_5430, x_5431, x_5432, x_5433, x_5434, x_5435, x_5436, x_5437, x_5438, x_5439, x_5440, x_5441, x_5442, x_5443, x_5444, x_5445, x_5446, x_5447, x_5448, x_5449, x_5450, x_5451, x_5452, x_5453, x_5454, x_5455, x_5456, x_5457, x_5458, x_5459, x_5460, x_5461, x_5462, x_5463, x_5464, x_5465, x_5466, x_5467, x_5468, x_5469, x_5470, x_5471, x_5472, x_5473, x_5474, x_5475, x_5476, x_5477, x_5478, x_5479, x_5480, x_5481, x_5482, x_5483, x_5484, x_5485, x_5486, x_5487, x_5488, x_5489, x_5490, x_5491, x_5492, x_5493, x_5494, x_5495, x_5496, x_5497, x_5498, x_5499, x_5500, x_5501, x_5502, x_5503, x_5504, x_5505, x_5506, x_5507, x_5508, x_5509, x_5510, x_5511, x_5512, x_5513, x_5514, x_5515, x_5516, x_5517, x_5518, x_5519, x_5520, x_5521, x_5522, x_5523, x_5524, x_5525, x_5526, x_5527, x_5528, x_5529, x_5530, x_5531, x_5532, x_5533, x_5534, x_5535, x_5536, x_5537, x_5538, x_5539, x_5540, x_5541, x_5542, x_5543, x_5544, x_5545, x_5546, x_5547, x_5548, x_5549, x_5550, x_5551, x_5552, x_5553, x_5554, x_5555, x_5556, x_5557, x_5558, x_5559, x_5560, x_5561, x_5562, x_5563, x_5564, x_5565, x_5566, x_5567, x_5568, x_5569, x_5570, x_5571, x_5572, x_5573, x_5574, x_5575, x_5576, x_5577, x_5578, x_5579, x_5580, x_5581, x_5582, x_5583, x_5584, x_5585, x_5586, x_5587, x_5588, x_5589, x_5590, x_5591, x_5592, x_5593, x_5594, x_5595, x_5596, x_5597, x_5598, x_5599, x_5600, x_5601, x_5602, x_5603, x_5604, x_5605, x_5606, x_5607, x_5608, x_5609, x_5610, x_5611, x_5612, x_5613, x_5614, x_5615, x_5616, x_5617, x_5618, x_5619, x_5620, x_5621, x_5622, x_5623, x_5624, x_5625, x_5626, x_5627, x_5628, x_5629, x_5630, x_5631, x_5632, x_5633, x_5634, x_5635, x_5636, x_5637, x_5638, x_5639, x_5640, x_5641, x_5642, x_5643, x_5644, x_5645, x_5646, x_5647, x_5648, x_5649, x_5650, x_5651, x_5652, x_5653, x_5654, x_5655, x_5656, x_5657, x_5658, x_5659, x_5660, x_5661, x_5662, x_5663, x_5664, x_5665, x_5666, x_5667, x_5668, x_5669, x_5670, x_5671, x_5672, x_5673, x_5674, x_5675, x_5676, x_5677, x_5678, x_5679, x_5680, x_5681, x_5682, x_5683, x_5684, x_5685, x_5686, x_5687, x_5688, x_5689, x_5690, x_5691, x_5692, x_5693, x_5694, x_5695, x_5696, x_5697, x_5698, x_5699, x_5700, x_5701, x_5702, x_5703, x_5704, x_5705, x_5706, x_5707, x_5708, x_5709, x_5710, x_5711, x_5712, x_5713, x_5714, x_5715, x_5716, x_5717, x_5718, x_5719, x_5720, x_5721, x_5722, x_5723, x_5724, x_5725, x_5726, x_5727, x_5728, x_5729, x_5730, x_5731, x_5732, x_5733, x_5734, x_5735, x_5736, x_5737, x_5738, x_5739, x_5740, x_5741, x_5742, x_5743, x_5744, x_5745, x_5746, x_5747, x_5748, x_5749, x_5750, x_5751, x_5752, x_5753, x_5754, x_5755, x_5756, x_5757, x_5758, x_5759, x_5760, x_5761, x_5762, x_5763, x_5764, x_5765, x_5766, x_5767, x_5768, x_5769, x_5770, x_5771, x_5772, x_5773, x_5774, x_5775, x_5776, x_5777, x_5778, x_5779, x_5780, x_5781, x_5782, x_5783, x_5784, x_5785, x_5786, x_5787, x_5788, x_5789, x_5790, x_5791, x_5792, x_5793, x_5794, x_5795, x_5796, x_5797, x_5798, x_5799, x_5800, x_5801, x_5802, x_5803, x_5804, x_5805, x_5806, x_5807, x_5808, x_5809, x_5810, x_5811, x_5812, x_5813, x_5814, x_5815, x_5816, x_5817, x_5818, x_5819, x_5820, x_5821, x_5822, x_5823, x_5824, x_5825, x_5826, x_5827, x_5828, x_5829, x_5830, x_5831, x_5832, x_5833, x_5834, x_5835, x_5836, x_5837, x_5838, x_5839, x_5840, x_5841, x_5842, x_5843, x_5844, x_5845, x_5846, x_5847, x_5848, x_5849, x_5850, x_5851, x_5852, x_5853, x_5854, x_5855, x_5856, x_5857, x_5858, x_5859, x_5860, x_5861, x_5862, x_5863, x_5864, x_5865, x_5866, x_5867, x_5868, x_5869, x_5870, x_5871, x_5872, x_5873, x_5874, x_5875, x_5876, x_5877, x_5878, x_5879, x_5880, x_5881, x_5882, x_5883, x_5884, x_5885, x_5886, x_5887, x_5888, x_5889, x_5890, x_5891, x_5892, x_5893, x_5894, x_5895, x_5896, x_5897, x_5898, x_5899, x_5900, x_5901, x_5902, x_5903, x_5904, x_5905, x_5906, x_5907, x_5908, x_5909, x_5910, x_5911, x_5912, x_5913, x_5914, x_5915, x_5916, x_5917, x_5918, x_5919, x_5920, x_5921, x_5922, x_5923, x_5924, x_5925, x_5926, x_5927, x_5928, x_5929, x_5930, x_5931, x_5932, x_5933, x_5934, x_5935, x_5936, x_5937, x_5938, x_5939, x_5940, x_5941, x_5942, x_5943, x_5944, x_5945, x_5946, x_5947, x_5948, x_5949, x_5950, x_5951, x_5952, x_5953, x_5954, x_5955, x_5956, x_5957, x_5958, x_5959, x_5960, x_5961, x_5962, x_5963, x_5964, x_5965, x_5966, x_5967, x_5968, x_5969, x_5970, x_5971, x_5972, x_5973, x_5974, x_5975, x_5976, x_5977, x_5978, x_5979, x_5980, x_5981, x_5982, x_5983, x_5984, x_5985, x_5986, x_5987, x_5988, x_5989, x_5990, x_5991, x_5992, x_5993, x_5994, x_5995, x_5996, x_5997, x_5998, x_5999, x_6000, x_6001, x_6002, x_6003, x_6004, x_6005, x_6006, x_6007, x_6008, x_6009, x_6010, x_6011, x_6012, x_6013, x_6014, x_6015, x_6016, x_6017, x_6018, x_6019, x_6020, x_6021, x_6022, x_6023, x_6024, x_6025, x_6026, x_6027, x_6028, x_6029, x_6030, x_6031, x_6032, x_6033, x_6034, x_6035, x_6036, x_6037, x_6038, x_6039, x_6040, x_6041, x_6042, x_6043, x_6044, x_6045, x_6046, x_6047, x_6048, x_6049, x_6050, x_6051, x_6052, x_6053, x_6054, x_6055, x_6056, x_6057, x_6058, x_6059, x_6060, x_6061, x_6062, x_6063, x_6064, x_6065, x_6066, x_6067, x_6068, x_6069, x_6070, x_6071, x_6072, x_6073, x_6074, x_6075, x_6076, x_6077, x_6078, x_6079, x_6080, x_6081, x_6082, x_6083, x_6084, x_6085, x_6086, x_6087, x_6088, x_6089, x_6090, x_6091, x_6092, x_6093, x_6094, x_6095, x_6096, x_6097, x_6098, x_6099, x_6100, x_6101, x_6102, x_6103, x_6104, x_6105, x_6106, x_6107, x_6108, x_6109, x_6110, x_6111, x_6112, x_6113, x_6114, x_6115, x_6116, x_6117, x_6118, x_6119, x_6120, x_6121, x_6122, x_6123, x_6124, x_6125, x_6126, x_6127, x_6128, x_6129, x_6130, x_6131, x_6132, x_6133, x_6134, x_6135, x_6136, x_6137, x_6138, x_6139, x_6140, x_6141, x_6142, x_6143, x_6144, x_6145, x_6146, x_6147, x_6148, x_6149, x_6150, x_6151, x_6152, x_6153, x_6154, x_6155, x_6156, x_6157, x_6158, x_6159, x_6160, x_6161, x_6162, x_6163, x_6164, x_6165, x_6166, x_6167, x_6168, x_6169, x_6170, x_6171, x_6172, x_6173, x_6174, x_6175, x_6176, x_6177, x_6178, x_6179, x_6180, x_6181, x_6182, x_6183, x_6184, x_6185, x_6186, x_6187, x_6188, x_6189, x_6190, x_6191, x_6192, x_6193, x_6194, x_6195, x_6196, x_6197, x_6198, x_6199, x_6200, x_6201, x_6202, x_6203, x_6204, x_6205, x_6206, x_6207, x_6208, x_6209, x_6210, x_6211, x_6212, x_6213, x_6214, x_6215, x_6216, x_6217, x_6218, x_6219, x_6220, x_6221, x_6222, x_6223, x_6224, x_6225, x_6226, x_6227, x_6228, x_6229, x_6230, x_6231, x_6232, x_6233, x_6234, x_6235, x_6236, x_6237, x_6238, x_6239, x_6240, x_6241, x_6242, x_6243, x_6244, x_6245, x_6246, x_6247, x_6248, x_6249, x_6250, x_6251, x_6252, x_6253, x_6254, o_1 );
input i_1;
input i_2;
input i_3;
input i_4;
input i_5;
input i_6;
input i_7;
input i_8;
input i_9;
input i_10;
input i_11;
input i_12;
input i_13;
input i_14;
input i_15;
input i_16;
input i_17;
input i_18;
input i_19;
input i_20;
input i_21;
input i_22;
input i_23;
input i_24;
input i_25;
input i_26;
input i_27;
input i_28;
input i_29;
input i_30;
input i_31;
input i_32;
input i_33;
input i_34;
input i_35;
input i_36;
input i_37;
input i_38;
input i_39;
input i_40;
input i_41;
input i_42;
input i_43;
input i_44;
input i_45;
input i_46;
input i_47;
input i_48;
input i_49;
input i_50;
input i_51;
input i_52;
input i_53;
input i_54;
input i_55;
input i_56;
input i_57;
input i_58;
input i_59;
input i_60;
input i_61;
input i_62;
input i_63;
input i_64;
input i_65;
input i_66;
input i_67;
input i_68;
input i_69;
input i_70;
input i_71;
input i_72;
input i_73;
input i_74;
input i_75;
input i_76;
input i_77;
input i_78;
input i_79;
input i_80;
input i_81;
input i_82;
input i_83;
input i_84;
input i_85;
input i_86;
input i_87;
input i_88;
input i_89;
input i_90;
input i_91;
input i_92;
input i_93;
input i_94;
input i_95;
input i_96;
input i_97;
input i_98;
input i_99;
input i_100;
input i_101;
input i_102;
input i_103;
input i_104;
input i_105;
input i_106;
input i_107;
input i_108;
input i_109;
input i_110;
input i_111;
input i_112;
input i_113;
input i_114;
input i_115;
input i_116;
input i_117;
input i_118;
input i_119;
input i_120;
input i_121;
input i_122;
input i_123;
input i_124;
input i_125;
input i_126;
input i_127;
input i_128;
input i_129;
input i_130;
input i_131;
input i_132;
input i_133;
input i_134;
input i_135;
input i_136;
input i_137;
input i_138;
input i_139;
input i_140;
input i_141;
input i_142;
input i_143;
input i_144;
input i_145;
input i_146;
input i_147;
input i_148;
input i_149;
input i_150;
input i_151;
input i_152;
input i_153;
input i_154;
input i_155;
input i_156;
input i_157;
input i_158;
input i_159;
input i_160;
input i_161;
input i_162;
input i_163;
input i_164;
input i_165;
input i_166;
input i_167;
input i_168;
input i_169;
input i_170;
input i_171;
input i_172;
input i_173;
input i_174;
input i_175;
input i_176;
input i_177;
input i_178;
input i_179;
input i_180;
input i_181;
input i_182;
input i_183;
input i_184;
input i_185;
input i_186;
input i_187;
input i_188;
input i_189;
input i_190;
input i_191;
input i_192;
input i_193;
input i_194;
input i_195;
input i_196;
input i_197;
input i_198;
input i_199;
input i_200;
input i_201;
input i_202;
input i_203;
input i_204;
input i_205;
input i_206;
input i_207;
input i_208;
input i_209;
input i_210;
input i_211;
input i_212;
input i_213;
input i_214;
input i_215;
input i_216;
input i_217;
input i_218;
input i_219;
input i_220;
input i_221;
input i_222;
input i_223;
input i_224;
input x_225;
input x_226;
input x_227;
input x_228;
input x_229;
input x_230;
input x_231;
input x_232;
input x_233;
input x_234;
input x_235;
input x_236;
input x_237;
input x_238;
input x_239;
input x_240;
input x_241;
input x_242;
input x_243;
input x_244;
input x_245;
input x_246;
input x_247;
input x_248;
input x_249;
input x_250;
input x_251;
input x_252;
input x_253;
input x_254;
input x_255;
input x_256;
input x_257;
input x_258;
input x_259;
input x_260;
input x_261;
input x_262;
input x_263;
input x_264;
input x_265;
input x_266;
input x_267;
input x_268;
input x_269;
input x_270;
input x_271;
input x_272;
input x_273;
input x_274;
input x_275;
input x_276;
input x_277;
input x_278;
input x_279;
input x_280;
input x_281;
input x_282;
input x_283;
input x_284;
input x_285;
input x_286;
input x_287;
input x_288;
input x_289;
input x_290;
input x_291;
input x_292;
input x_293;
input x_294;
input x_295;
input x_296;
input x_297;
input x_298;
input x_299;
input x_300;
input x_301;
input x_302;
input x_303;
input x_304;
input x_305;
input x_306;
input x_307;
input x_308;
input x_309;
input x_310;
input x_311;
input x_312;
input x_313;
input x_314;
input x_315;
input x_316;
input x_317;
input x_318;
input x_319;
input x_320;
input x_321;
input x_322;
input x_323;
input x_324;
input x_325;
input x_326;
input x_327;
input x_328;
input x_329;
input x_330;
input x_331;
input x_332;
input x_333;
input x_334;
input x_335;
input x_336;
input x_337;
input x_338;
input x_339;
input x_340;
input x_341;
input x_342;
input x_343;
input x_344;
input x_345;
input x_346;
input x_347;
input x_348;
input x_349;
input x_350;
input x_351;
input x_352;
input x_353;
input x_354;
input x_355;
input x_356;
input x_357;
input x_358;
input x_359;
input x_360;
input x_361;
input x_362;
input x_363;
input x_364;
input x_365;
input x_366;
input x_367;
input x_368;
input x_369;
input x_370;
input x_371;
input x_372;
input x_373;
input x_374;
input x_375;
input x_376;
input x_377;
input x_378;
input x_379;
input x_380;
input x_381;
input x_382;
input x_383;
input x_384;
input x_385;
input x_386;
input x_387;
input x_388;
input x_389;
input x_390;
input x_391;
input x_392;
input x_393;
input x_394;
input x_395;
input x_396;
input x_397;
input x_398;
input x_399;
input x_400;
input x_401;
input x_402;
input x_403;
input x_404;
input x_405;
input x_406;
input x_407;
input x_408;
input x_409;
input x_410;
input x_411;
input x_412;
input x_413;
input x_414;
input x_415;
input x_416;
input x_417;
input x_418;
input x_419;
input x_420;
input x_421;
input x_422;
input x_423;
input x_424;
input x_425;
input x_426;
input x_427;
input x_428;
input x_429;
input x_430;
input x_431;
input x_432;
input x_433;
input x_434;
input x_435;
input x_436;
input x_437;
input x_438;
input x_439;
input x_440;
input x_441;
input x_442;
input x_443;
input x_444;
input x_445;
input x_446;
input x_447;
input x_448;
input x_449;
input x_450;
input x_451;
input x_452;
input x_453;
input x_454;
input x_455;
input x_456;
input x_457;
input x_458;
input x_459;
input x_460;
input x_461;
input x_462;
input x_463;
input x_464;
input x_465;
input x_466;
input x_467;
input x_468;
input x_469;
input x_470;
input x_471;
input x_472;
input x_473;
input x_474;
input x_475;
input x_476;
input x_477;
input x_478;
input x_479;
input x_480;
input x_481;
input x_482;
input x_483;
input x_484;
input x_485;
input x_486;
input x_487;
input x_488;
input x_489;
input x_490;
input x_491;
input x_492;
input x_493;
input x_494;
input x_495;
input x_496;
input x_497;
input x_498;
input x_499;
input x_500;
input x_501;
input x_502;
input x_503;
input x_504;
input x_505;
input x_506;
input x_507;
input x_508;
input x_509;
input x_510;
input x_511;
input x_512;
input x_513;
input x_514;
input x_515;
input x_516;
input x_517;
input x_518;
input x_519;
input x_520;
input x_521;
input x_522;
input x_523;
input x_524;
input x_525;
input x_526;
input x_527;
input x_528;
input x_529;
input x_530;
input x_531;
input x_532;
input x_533;
input x_534;
input x_535;
input x_536;
input x_537;
input x_538;
input x_539;
input x_540;
input x_541;
input x_542;
input x_543;
input x_544;
input x_545;
input x_546;
input x_547;
input x_548;
input x_549;
input x_550;
input x_551;
input x_552;
input x_553;
input x_554;
input x_555;
input x_556;
input x_557;
input x_558;
input x_559;
input x_560;
input x_561;
input x_562;
input x_563;
input x_564;
input x_565;
input x_566;
input x_567;
input x_568;
input x_569;
input x_570;
input x_571;
input x_572;
input x_573;
input x_574;
input x_575;
input x_576;
input x_577;
input x_578;
input x_579;
input x_580;
input x_581;
input x_582;
input x_583;
input x_584;
input x_585;
input x_586;
input x_587;
input x_588;
input x_589;
input x_590;
input x_591;
input x_592;
input x_593;
input x_594;
input x_595;
input x_596;
input x_597;
input x_598;
input x_599;
input x_600;
input x_601;
input x_602;
input x_603;
input x_604;
input x_605;
input x_606;
input x_607;
input x_608;
input x_609;
input x_610;
input x_611;
input x_612;
input x_613;
input x_614;
input x_615;
input x_616;
input x_617;
input x_618;
input x_619;
input x_620;
input x_621;
input x_622;
input x_623;
input x_624;
input x_625;
input x_626;
input x_627;
input x_628;
input x_629;
input x_630;
input x_631;
input x_632;
input x_633;
input x_634;
input x_635;
input x_636;
input x_637;
input x_638;
input x_639;
input x_640;
input x_641;
input x_642;
input x_643;
input x_644;
input x_645;
input x_646;
input x_647;
input x_648;
input x_649;
input x_650;
input x_651;
input x_652;
input x_653;
input x_654;
input x_655;
input x_656;
input x_657;
input x_658;
input x_659;
input x_660;
input x_661;
input x_662;
input x_663;
input x_664;
input x_665;
input x_666;
input x_667;
input x_668;
input x_669;
input x_670;
input x_671;
input x_672;
input x_673;
input x_674;
input x_675;
input x_676;
input x_677;
input x_678;
input x_679;
input x_680;
input x_681;
input x_682;
input x_683;
input x_684;
input x_685;
input x_686;
input x_687;
input x_688;
input x_689;
input x_690;
input x_691;
input x_692;
input x_693;
input x_694;
input x_695;
input x_696;
input x_697;
input x_698;
input x_699;
input x_700;
input x_701;
input x_702;
input x_703;
input x_704;
input x_705;
input x_706;
input x_707;
input x_708;
input x_709;
input x_710;
input x_711;
input x_712;
input x_713;
input x_714;
input x_715;
input x_716;
input x_717;
input x_718;
input x_719;
input x_720;
input x_721;
input x_722;
input x_723;
input x_724;
input x_725;
input x_726;
input x_727;
input x_728;
input x_729;
input x_730;
input x_731;
input x_732;
input x_733;
input x_734;
input x_735;
input x_736;
input x_737;
input x_738;
input x_739;
input x_740;
input x_741;
input x_742;
input x_743;
input x_744;
input x_745;
input x_746;
input x_747;
input x_748;
input x_749;
input x_750;
input x_751;
input x_752;
input x_753;
input x_754;
input x_755;
input x_756;
input x_757;
input x_758;
input x_759;
input x_760;
input x_761;
input x_762;
input x_763;
input x_764;
input x_765;
input x_766;
input x_767;
input x_768;
input x_769;
input x_770;
input x_771;
input x_772;
input x_773;
input x_774;
input x_775;
input x_776;
input x_777;
input x_778;
input x_779;
input x_780;
input x_781;
input x_782;
input x_783;
input x_784;
input x_785;
input x_786;
input x_787;
input x_788;
input x_789;
input x_790;
input x_791;
input x_792;
input x_793;
input x_794;
input x_795;
input x_796;
input x_797;
input x_798;
input x_799;
input x_800;
input x_801;
input x_802;
input x_803;
input x_804;
input x_805;
input x_806;
input x_807;
input x_808;
input x_809;
input x_810;
input x_811;
input x_812;
input x_813;
input x_814;
input x_815;
input x_816;
input x_817;
input x_818;
input x_819;
input x_820;
input x_821;
input x_822;
input x_823;
input x_824;
input x_825;
input x_826;
input x_827;
input x_828;
input x_829;
input x_830;
input x_831;
input x_832;
input x_833;
input x_834;
input x_835;
input x_836;
input x_837;
input x_838;
input x_839;
input x_840;
input x_841;
input x_842;
input x_843;
input x_844;
input x_845;
input x_846;
input x_847;
input x_848;
input x_849;
input x_850;
input x_851;
input x_852;
input x_853;
input x_854;
input x_855;
input x_856;
input x_857;
input x_858;
input x_859;
input x_860;
input x_861;
input x_862;
input x_863;
input x_864;
input x_865;
input x_866;
input x_867;
input x_868;
input x_869;
input x_870;
input x_871;
input x_872;
input x_873;
input x_874;
input x_875;
input x_876;
input x_877;
input x_878;
input x_879;
input x_880;
input x_881;
input x_882;
input x_883;
input x_884;
input x_885;
input x_886;
input x_887;
input x_888;
input x_889;
input x_890;
input x_891;
input x_892;
input x_893;
input x_894;
input x_895;
input x_896;
input x_897;
input x_898;
input x_899;
input x_900;
input x_901;
input x_902;
input x_903;
input x_904;
input x_905;
input x_906;
input x_907;
input x_908;
input x_909;
input x_910;
input x_911;
input x_912;
input x_913;
input x_914;
input x_915;
input x_916;
input x_917;
input x_918;
input x_919;
input x_920;
input x_921;
input x_922;
input x_923;
input x_924;
input x_925;
input x_926;
input x_927;
input x_928;
input x_929;
input x_930;
input x_931;
input x_932;
input x_933;
input x_934;
input x_935;
input x_936;
input x_937;
input x_938;
input x_939;
input x_940;
input x_941;
input x_942;
input x_943;
input x_944;
input x_945;
input x_946;
input x_947;
input x_948;
input x_949;
input x_950;
input x_951;
input x_952;
input x_953;
input x_954;
input x_955;
input x_956;
input x_957;
input x_958;
input x_959;
input x_960;
input x_961;
input x_962;
input x_963;
input x_964;
input x_965;
input x_966;
input x_967;
input x_968;
input x_969;
input x_970;
input x_971;
input x_972;
input x_973;
input x_974;
input x_975;
input x_976;
input x_977;
input x_978;
input x_979;
input x_980;
input x_981;
input x_982;
input x_983;
input x_984;
input x_985;
input x_986;
input x_987;
input x_988;
input x_989;
input x_990;
input x_991;
input x_992;
input x_993;
input x_994;
input x_995;
input x_996;
input x_997;
input x_998;
input x_999;
input x_1000;
input x_1001;
input x_1002;
input x_1003;
input x_1004;
input x_1005;
input x_1006;
input x_1007;
input x_1008;
input x_1009;
input x_1010;
input x_1011;
input x_1012;
input x_1013;
input x_1014;
input x_1015;
input x_1016;
input x_1017;
input x_1018;
input x_1019;
input x_1020;
input x_1021;
input x_1022;
input x_1023;
input x_1024;
input x_1025;
input x_1026;
input x_1027;
input x_1028;
input x_1029;
input x_1030;
input x_1031;
input x_1032;
input x_1033;
input x_1034;
input x_1035;
input x_1036;
input x_1037;
input x_1038;
input x_1039;
input x_1040;
input x_1041;
input x_1042;
input x_1043;
input x_1044;
input x_1045;
input x_1046;
input x_1047;
input x_1048;
input x_1049;
input x_1050;
input x_1051;
input x_1052;
input x_1053;
input x_1054;
input x_1055;
input x_1056;
input x_1057;
input x_1058;
input x_1059;
input x_1060;
input x_1061;
input x_1062;
input x_1063;
input x_1064;
input x_1065;
input x_1066;
input x_1067;
input x_1068;
input x_1069;
input x_1070;
input x_1071;
input x_1072;
input x_1073;
input x_1074;
input x_1075;
input x_1076;
input x_1077;
input x_1078;
input x_1079;
input x_1080;
input x_1081;
input x_1082;
input x_1083;
input x_1084;
input x_1085;
input x_1086;
input x_1087;
input x_1088;
input x_1089;
input x_1090;
input x_1091;
input x_1092;
input x_1093;
input x_1094;
input x_1095;
input x_1096;
input x_1097;
input x_1098;
input x_1099;
input x_1100;
input x_1101;
input x_1102;
input x_1103;
input x_1104;
input x_1105;
input x_1106;
input x_1107;
input x_1108;
input x_1109;
input x_1110;
input x_1111;
input x_1112;
input x_1113;
input x_1114;
input x_1115;
input x_1116;
input x_1117;
input x_1118;
input x_1119;
input x_1120;
input x_1121;
input x_1122;
input x_1123;
input x_1124;
input x_1125;
input x_1126;
input x_1127;
input x_1128;
input x_1129;
input x_1130;
input x_1131;
input x_1132;
input x_1133;
input x_1134;
input x_1135;
input x_1136;
input x_1137;
input x_1138;
input x_1139;
input x_1140;
input x_1141;
input x_1142;
input x_1143;
input x_1144;
input x_1145;
input x_1146;
input x_1147;
input x_1148;
input x_1149;
input x_1150;
input x_1151;
input x_1152;
input x_1153;
input x_1154;
input x_1155;
input x_1156;
input x_1157;
input x_1158;
input x_1159;
input x_1160;
input x_1161;
input x_1162;
input x_1163;
input x_1164;
input x_1165;
input x_1166;
input x_1167;
input x_1168;
input x_1169;
input x_1170;
input x_1171;
input x_1172;
input x_1173;
input x_1174;
input x_1175;
input x_1176;
input x_1177;
input x_1178;
input x_1179;
input x_1180;
input x_1181;
input x_1182;
input x_1183;
input x_1184;
input x_1185;
input x_1186;
input x_1187;
input x_1188;
input x_1189;
input x_1190;
input x_1191;
input x_1192;
input x_1193;
input x_1194;
input x_1195;
input x_1196;
input x_1197;
input x_1198;
input x_1199;
input x_1200;
input x_1201;
input x_1202;
input x_1203;
input x_1204;
input x_1205;
input x_1206;
input x_1207;
input x_1208;
input x_1209;
input x_1210;
input x_1211;
input x_1212;
input x_1213;
input x_1214;
input x_1215;
input x_1216;
input x_1217;
input x_1218;
input x_1219;
input x_1220;
input x_1221;
input x_1222;
input x_1223;
input x_1224;
input x_1225;
input x_1226;
input x_1227;
input x_1228;
input x_1229;
input x_1230;
input x_1231;
input x_1232;
input x_1233;
input x_1234;
input x_1235;
input x_1236;
input x_1237;
input x_1238;
input x_1239;
input x_1240;
input x_1241;
input x_1242;
input x_1243;
input x_1244;
input x_1245;
input x_1246;
input x_1247;
input x_1248;
input x_1249;
input x_1250;
input x_1251;
input x_1252;
input x_1253;
input x_1254;
input x_1255;
input x_1256;
input x_1257;
input x_1258;
input x_1259;
input x_1260;
input x_1261;
input x_1262;
input x_1263;
input x_1264;
input x_1265;
input x_1266;
input x_1267;
input x_1268;
input x_1269;
input x_1270;
input x_1271;
input x_1272;
input x_1273;
input x_1274;
input x_1275;
input x_1276;
input x_1277;
input x_1278;
input x_1279;
input x_1280;
input x_1281;
input x_1282;
input x_1283;
input x_1284;
input x_1285;
input x_1286;
input x_1287;
input x_1288;
input x_1289;
input x_1290;
input x_1291;
input x_1292;
input x_1293;
input x_1294;
input x_1295;
input x_1296;
input x_1297;
input x_1298;
input x_1299;
input x_1300;
input x_1301;
input x_1302;
input x_1303;
input x_1304;
input x_1305;
input x_1306;
input x_1307;
input x_1308;
input x_1309;
input x_1310;
input x_1311;
input x_1312;
input x_1313;
input x_1314;
input x_1315;
input x_1316;
input x_1317;
input x_1318;
input x_1319;
input x_1320;
input x_1321;
input x_1322;
input x_1323;
input x_1324;
input x_1325;
input x_1326;
input x_1327;
input x_1328;
input x_1329;
input x_1330;
input x_1331;
input x_1332;
input x_1333;
input x_1334;
input x_1335;
input x_1336;
input x_1337;
input x_1338;
input x_1339;
input x_1340;
input x_1341;
input x_1342;
input x_1343;
input x_1344;
input x_1345;
input x_1346;
input x_1347;
input x_1348;
input x_1349;
input x_1350;
input x_1351;
input x_1352;
input x_1353;
input x_1354;
input x_1355;
input x_1356;
input x_1357;
input x_1358;
input x_1359;
input x_1360;
input x_1361;
input x_1362;
input x_1363;
input x_1364;
input x_1365;
input x_1366;
input x_1367;
input x_1368;
input x_1369;
input x_1370;
input x_1371;
input x_1372;
input x_1373;
input x_1374;
input x_1375;
input x_1376;
input x_1377;
input x_1378;
input x_1379;
input x_1380;
input x_1381;
input x_1382;
input x_1383;
input x_1384;
input x_1385;
input x_1386;
input x_1387;
input x_1388;
input x_1389;
input x_1390;
input x_1391;
input x_1392;
input x_1393;
input x_1394;
input x_1395;
input x_1396;
input x_1397;
input x_1398;
input x_1399;
input x_1400;
input x_1401;
input x_1402;
input x_1403;
input x_1404;
input x_1405;
input x_1406;
input x_1407;
input x_1408;
input x_1409;
input x_1410;
input x_1411;
input x_1412;
input x_1413;
input x_1414;
input x_1415;
input x_1416;
input x_1417;
input x_1418;
input x_1419;
input x_1420;
input x_1421;
input x_1422;
input x_1423;
input x_1424;
input x_1425;
input x_1426;
input x_1427;
input x_1428;
input x_1429;
input x_1430;
input x_1431;
input x_1432;
input x_1433;
input x_1434;
input x_1435;
input x_1436;
input x_1437;
input x_1438;
input x_1439;
input x_1440;
input x_1441;
input x_1442;
input x_1443;
input x_1444;
input x_1445;
input x_1446;
input x_1447;
input x_1448;
input x_1449;
input x_1450;
input x_1451;
input x_1452;
input x_1453;
input x_1454;
input x_1455;
input x_1456;
input x_1457;
input x_1458;
input x_1459;
input x_1460;
input x_1461;
input x_1462;
input x_1463;
input x_1464;
input x_1465;
input x_1466;
input x_1467;
input x_1468;
input x_1469;
input x_1470;
input x_1471;
input x_1472;
input x_1473;
input x_1474;
input x_1475;
input x_1476;
input x_1477;
input x_1478;
input x_1479;
input x_1480;
input x_1481;
input x_1482;
input x_1483;
input x_1484;
input x_1485;
input x_1486;
input x_1487;
input x_1488;
input x_1489;
input x_1490;
input x_1491;
input x_1492;
input x_1493;
input x_1494;
input x_1495;
input x_1496;
input x_1497;
input x_1498;
input x_1499;
input x_1500;
input x_1501;
input x_1502;
input x_1503;
input x_1504;
input x_1505;
input x_1506;
input x_1507;
input x_1508;
input x_1509;
input x_1510;
input x_1511;
input x_1512;
input x_1513;
input x_1514;
input x_1515;
input x_1516;
input x_1517;
input x_1518;
input x_1519;
input x_1520;
input x_1521;
input x_1522;
input x_1523;
input x_1524;
input x_1525;
input x_1526;
input x_1527;
input x_1528;
input x_1529;
input x_1530;
input x_1531;
input x_1532;
input x_1533;
input x_1534;
input x_1535;
input x_1536;
input x_1537;
input x_1538;
input x_1539;
input x_1540;
input x_1541;
input x_1542;
input x_1543;
input x_1544;
input x_1545;
input x_1546;
input x_1547;
input x_1548;
input x_1549;
input x_1550;
input x_1551;
input x_1552;
input x_1553;
input x_1554;
input x_1555;
input x_1556;
input x_1557;
input x_1558;
input x_1559;
input x_1560;
input x_1561;
input x_1562;
input x_1563;
input x_1564;
input x_1565;
input x_1566;
input x_1567;
input x_1568;
input x_1569;
input x_1570;
input x_1571;
input x_1572;
input x_1573;
input x_1574;
input x_1575;
input x_1576;
input x_1577;
input x_1578;
input x_1579;
input x_1580;
input x_1581;
input x_1582;
input x_1583;
input x_1584;
input x_1585;
input x_1586;
input x_1587;
input x_1588;
input x_1589;
input x_1590;
input x_1591;
input x_1592;
input x_1593;
input x_1594;
input x_1595;
input x_1596;
input x_1597;
input x_1598;
input x_1599;
input x_1600;
input x_1601;
input x_1602;
input x_1603;
input x_1604;
input x_1605;
input x_1606;
input x_1607;
input x_1608;
input x_1609;
input x_1610;
input x_1611;
input x_1612;
input x_1613;
input x_1614;
input x_1615;
input x_1616;
input x_1617;
input x_1618;
input x_1619;
input x_1620;
input x_1621;
input x_1622;
input x_1623;
input x_1624;
input x_1625;
input x_1626;
input x_1627;
input x_1628;
input x_1629;
input x_1630;
input x_1631;
input x_1632;
input x_1633;
input x_1634;
input x_1635;
input x_1636;
input x_1637;
input x_1638;
input x_1639;
input x_1640;
input x_1641;
input x_1642;
input x_1643;
input x_1644;
input x_1645;
input x_1646;
input x_1647;
input x_1648;
input x_1649;
input x_1650;
input x_1651;
input x_1652;
input x_1653;
input x_1654;
input x_1655;
input x_1656;
input x_1657;
input x_1658;
input x_1659;
input x_1660;
input x_1661;
input x_1662;
input x_1663;
input x_1664;
input x_1665;
input x_1666;
input x_1667;
input x_1668;
input x_1669;
input x_1670;
input x_1671;
input x_1672;
input x_1673;
input x_1674;
input x_1675;
input x_1676;
input x_1677;
input x_1678;
input x_1679;
input x_1680;
input x_1681;
input x_1682;
input x_1683;
input x_1684;
input x_1685;
input x_1686;
input x_1687;
input x_1688;
input x_1689;
input x_1690;
input x_1691;
input x_1692;
input x_1693;
input x_1694;
input x_1695;
input x_1696;
input x_1697;
input x_1698;
input x_1699;
input x_1700;
input x_1701;
input x_1702;
input x_1703;
input x_1704;
input x_1705;
input x_1706;
input x_1707;
input x_1708;
input x_1709;
input x_1710;
input x_1711;
input x_1712;
input x_1713;
input x_1714;
input x_1715;
input x_1716;
input x_1717;
input x_1718;
input x_1719;
input x_1720;
input x_1721;
input x_1722;
input x_1723;
input x_1724;
input x_1725;
input x_1726;
input x_1727;
input x_1728;
input x_1729;
input x_1730;
input x_1731;
input x_1732;
input x_1733;
input x_1734;
input x_1735;
input x_1736;
input x_1737;
input x_1738;
input x_1739;
input x_1740;
input x_1741;
input x_1742;
input x_1743;
input x_1744;
input x_1745;
input x_1746;
input x_1747;
input x_1748;
input x_1749;
input x_1750;
input x_1751;
input x_1752;
input x_1753;
input x_1754;
input x_1755;
input x_1756;
input x_1757;
input x_1758;
input x_1759;
input x_1760;
input x_1761;
input x_1762;
input x_1763;
input x_1764;
input x_1765;
input x_1766;
input x_1767;
input x_1768;
input x_1769;
input x_1770;
input x_1771;
input x_1772;
input x_1773;
input x_1774;
input x_1775;
input x_1776;
input x_1777;
input x_1778;
input x_1779;
input x_1780;
input x_1781;
input x_1782;
input x_1783;
input x_1784;
input x_1785;
input x_1786;
input x_1787;
input x_1788;
input x_1789;
input x_1790;
input x_1791;
input x_1792;
input x_1793;
input x_1794;
input x_1795;
input x_1796;
input x_1797;
input x_1798;
input x_1799;
input x_1800;
input x_1801;
input x_1802;
input x_1803;
input x_1804;
input x_1805;
input x_1806;
input x_1807;
input x_1808;
input x_1809;
input x_1810;
input x_1811;
input x_1812;
input x_1813;
input x_1814;
input x_1815;
input x_1816;
input x_1817;
input x_1818;
input x_1819;
input x_1820;
input x_1821;
input x_1822;
input x_1823;
input x_1824;
input x_1825;
input x_1826;
input x_1827;
input x_1828;
input x_1829;
input x_1830;
input x_1831;
input x_1832;
input x_1833;
input x_1834;
input x_1835;
input x_1836;
input x_1837;
input x_1838;
input x_1839;
input x_1840;
input x_1841;
input x_1842;
input x_1843;
input x_1844;
input x_1845;
input x_1846;
input x_1847;
input x_1848;
input x_1849;
input x_1850;
input x_1851;
input x_1852;
input x_1853;
input x_1854;
input x_1855;
input x_1856;
input x_1857;
input x_1858;
input x_1859;
input x_1860;
input x_1861;
input x_1862;
input x_1863;
input x_1864;
input x_1865;
input x_1866;
input x_1867;
input x_1868;
input x_1869;
input x_1870;
input x_1871;
input x_1872;
input x_1873;
input x_1874;
input x_1875;
input x_1876;
input x_1877;
input x_1878;
input x_1879;
input x_1880;
input x_1881;
input x_1882;
input x_1883;
input x_1884;
input x_1885;
input x_1886;
input x_1887;
input x_1888;
input x_1889;
input x_1890;
input x_1891;
input x_1892;
input x_1893;
input x_1894;
input x_1895;
input x_1896;
input x_1897;
input x_1898;
input x_1899;
input x_1900;
input x_1901;
input x_1902;
input x_1903;
input x_1904;
input x_1905;
input x_1906;
input x_1907;
input x_1908;
input x_1909;
input x_1910;
input x_1911;
input x_1912;
input x_1913;
input x_1914;
input x_1915;
input x_1916;
input x_1917;
input x_1918;
input x_1919;
input x_1920;
input x_1921;
input x_1922;
input x_1923;
input x_1924;
input x_1925;
input x_1926;
input x_1927;
input x_1928;
input x_1929;
input x_1930;
input x_1931;
input x_1932;
input x_1933;
input x_1934;
input x_1935;
input x_1936;
input x_1937;
input x_1938;
input x_1939;
input x_1940;
input x_1941;
input x_1942;
input x_1943;
input x_1944;
input x_1945;
input x_1946;
input x_1947;
input x_1948;
input x_1949;
input x_1950;
input x_1951;
input x_1952;
input x_1953;
input x_1954;
input x_1955;
input x_1956;
input x_1957;
input x_1958;
input x_1959;
input x_1960;
input x_1961;
input x_1962;
input x_1963;
input x_1964;
input x_1965;
input x_1966;
input x_1967;
input x_1968;
input x_1969;
input x_1970;
input x_1971;
input x_1972;
input x_1973;
input x_1974;
input x_1975;
input x_1976;
input x_1977;
input x_1978;
input x_1979;
input x_1980;
input x_1981;
input x_1982;
input x_1983;
input x_1984;
input x_1985;
input x_1986;
input x_1987;
input x_1988;
input x_1989;
input x_1990;
input x_1991;
input x_1992;
input x_1993;
input x_1994;
input x_1995;
input x_1996;
input x_1997;
input x_1998;
input x_1999;
input x_2000;
input x_2001;
input x_2002;
input x_2003;
input x_2004;
input x_2005;
input x_2006;
input x_2007;
input x_2008;
input x_2009;
input x_2010;
input x_2011;
input x_2012;
input x_2013;
input x_2014;
input x_2015;
input x_2016;
input x_2017;
input x_2018;
input x_2019;
input x_2020;
input x_2021;
input x_2022;
input x_2023;
input x_2024;
input x_2025;
input x_2026;
input x_2027;
input x_2028;
input x_2029;
input x_2030;
input x_2031;
input x_2032;
input x_2033;
input x_2034;
input x_2035;
input x_2036;
input x_2037;
input x_2038;
input x_2039;
input x_2040;
input x_2041;
input x_2042;
input x_2043;
input x_2044;
input x_2045;
input x_2046;
input x_2047;
input x_2048;
input x_2049;
input x_2050;
input x_2051;
input x_2052;
input x_2053;
input x_2054;
input x_2055;
input x_2056;
input x_2057;
input x_2058;
input x_2059;
input x_2060;
input x_2061;
input x_2062;
input x_2063;
input x_2064;
input x_2065;
input x_2066;
input x_2067;
input x_2068;
input x_2069;
input x_2070;
input x_2071;
input x_2072;
input x_2073;
input x_2074;
input x_2075;
input x_2076;
input x_2077;
input x_2078;
input x_2079;
input x_2080;
input x_2081;
input x_2082;
input x_2083;
input x_2084;
input x_2085;
input x_2086;
input x_2087;
input x_2088;
input x_2089;
input x_2090;
input x_2091;
input x_2092;
input x_2093;
input x_2094;
input x_2095;
input x_2096;
input x_2097;
input x_2098;
input x_2099;
input x_2100;
input x_2101;
input x_2102;
input x_2103;
input x_2104;
input x_2105;
input x_2106;
input x_2107;
input x_2108;
input x_2109;
input x_2110;
input x_2111;
input x_2112;
input x_2113;
input x_2114;
input x_2115;
input x_2116;
input x_2117;
input x_2118;
input x_2119;
input x_2120;
input x_2121;
input x_2122;
input x_2123;
input x_2124;
input x_2125;
input x_2126;
input x_2127;
input x_2128;
input x_2129;
input x_2130;
input x_2131;
input x_2132;
input x_2133;
input x_2134;
input x_2135;
input x_2136;
input x_2137;
input x_2138;
input x_2139;
input x_2140;
input x_2141;
input x_2142;
input x_2143;
input x_2144;
input x_2145;
input x_2146;
input x_2147;
input x_2148;
input x_2149;
input x_2150;
input x_2151;
input x_2152;
input x_2153;
input x_2154;
input x_2155;
input x_2156;
input x_2157;
input x_2158;
input x_2159;
input x_2160;
input x_2161;
input x_2162;
input x_2163;
input x_2164;
input x_2165;
input x_2166;
input x_2167;
input x_2168;
input x_2169;
input x_2170;
input x_2171;
input x_2172;
input x_2173;
input x_2174;
input x_2175;
input x_2176;
input x_2177;
input x_2178;
input x_2179;
input x_2180;
input x_2181;
input x_2182;
input x_2183;
input x_2184;
input x_2185;
input x_2186;
input x_2187;
input x_2188;
input x_2189;
input x_2190;
input x_2191;
input x_2192;
input x_2193;
input x_2194;
input x_2195;
input x_2196;
input x_2197;
input x_2198;
input x_2199;
input x_2200;
input x_2201;
input x_2202;
input x_2203;
input x_2204;
input x_2205;
input x_2206;
input x_2207;
input x_2208;
input x_2209;
input x_2210;
input x_2211;
input x_2212;
input x_2213;
input x_2214;
input x_2215;
input x_2216;
input x_2217;
input x_2218;
input x_2219;
input x_2220;
input x_2221;
input x_2222;
input x_2223;
input x_2224;
input x_2225;
input x_2226;
input x_2227;
input x_2228;
input x_2229;
input x_2230;
input x_2231;
input x_2232;
input x_2233;
input x_2234;
input x_2235;
input x_2236;
input x_2237;
input x_2238;
input x_2239;
input x_2240;
input x_2241;
input x_2242;
input x_2243;
input x_2244;
input x_2245;
input x_2246;
input x_2247;
input x_2248;
input x_2249;
input x_2250;
input x_2251;
input x_2252;
input x_2253;
input x_2254;
input x_2255;
input x_2256;
input x_2257;
input x_2258;
input x_2259;
input x_2260;
input x_2261;
input x_2262;
input x_2263;
input x_2264;
input x_2265;
input x_2266;
input x_2267;
input x_2268;
input x_2269;
input x_2270;
input x_2271;
input x_2272;
input x_2273;
input x_2274;
input x_2275;
input x_2276;
input x_2277;
input x_2278;
input x_2279;
input x_2280;
input x_2281;
input x_2282;
input x_2283;
input x_2284;
input x_2285;
input x_2286;
input x_2287;
input x_2288;
input x_2289;
input x_2290;
input x_2291;
input x_2292;
input x_2293;
input x_2294;
input x_2295;
input x_2296;
input x_2297;
input x_2298;
input x_2299;
input x_2300;
input x_2301;
input x_2302;
input x_2303;
input x_2304;
input x_2305;
input x_2306;
input x_2307;
input x_2308;
input x_2309;
input x_2310;
input x_2311;
input x_2312;
input x_2313;
input x_2314;
input x_2315;
input x_2316;
input x_2317;
input x_2318;
input x_2319;
input x_2320;
input x_2321;
input x_2322;
input x_2323;
input x_2324;
input x_2325;
input x_2326;
input x_2327;
input x_2328;
input x_2329;
input x_2330;
input x_2331;
input x_2332;
input x_2333;
input x_2334;
input x_2335;
input x_2336;
input x_2337;
input x_2338;
input x_2339;
input x_2340;
input x_2341;
input x_2342;
input x_2343;
input x_2344;
input x_2345;
input x_2346;
input x_2347;
input x_2348;
input x_2349;
input x_2350;
input x_2351;
input x_2352;
input x_2353;
input x_2354;
input x_2355;
input x_2356;
input x_2357;
input x_2358;
input x_2359;
input x_2360;
input x_2361;
input x_2362;
input x_2363;
input x_2364;
input x_2365;
input x_2366;
input x_2367;
input x_2368;
input x_2369;
input x_2370;
input x_2371;
input x_2372;
input x_2373;
input x_2374;
input x_2375;
input x_2376;
input x_2377;
input x_2378;
input x_2379;
input x_2380;
input x_2381;
input x_2382;
input x_2383;
input x_2384;
input x_2385;
input x_2386;
input x_2387;
input x_2388;
input x_2389;
input x_2390;
input x_2391;
input x_2392;
input x_2393;
input x_2394;
input x_2395;
input x_2396;
input x_2397;
input x_2398;
input x_2399;
input x_2400;
input x_2401;
input x_2402;
input x_2403;
input x_2404;
input x_2405;
input x_2406;
input x_2407;
input x_2408;
input x_2409;
input x_2410;
input x_2411;
input x_2412;
input x_2413;
input x_2414;
input x_2415;
input x_2416;
input x_2417;
input x_2418;
input x_2419;
input x_2420;
input x_2421;
input x_2422;
input x_2423;
input x_2424;
input x_2425;
input x_2426;
input x_2427;
input x_2428;
input x_2429;
input x_2430;
input x_2431;
input x_2432;
input x_2433;
input x_2434;
input x_2435;
input x_2436;
input x_2437;
input x_2438;
input x_2439;
input x_2440;
input x_2441;
input x_2442;
input x_2443;
input x_2444;
input x_2445;
input x_2446;
input x_2447;
input x_2448;
input x_2449;
input x_2450;
input x_2451;
input x_2452;
input x_2453;
input x_2454;
input x_2455;
input x_2456;
input x_2457;
input x_2458;
input x_2459;
input x_2460;
input x_2461;
input x_2462;
input x_2463;
input x_2464;
input x_2465;
input x_2466;
input x_2467;
input x_2468;
input x_2469;
input x_2470;
input x_2471;
input x_2472;
input x_2473;
input x_2474;
input x_2475;
input x_2476;
input x_2477;
input x_2478;
input x_2479;
input x_2480;
input x_2481;
input x_2482;
input x_2483;
input x_2484;
input x_2485;
input x_2486;
input x_2487;
input x_2488;
input x_2489;
input x_2490;
input x_2491;
input x_2492;
input x_2493;
input x_2494;
input x_2495;
input x_2496;
input x_2497;
input x_2498;
input x_2499;
input x_2500;
input x_2501;
input x_2502;
input x_2503;
input x_2504;
input x_2505;
input x_2506;
input x_2507;
input x_2508;
input x_2509;
input x_2510;
input x_2511;
input x_2512;
input x_2513;
input x_2514;
input x_2515;
input x_2516;
input x_2517;
input x_2518;
input x_2519;
input x_2520;
input x_2521;
input x_2522;
input x_2523;
input x_2524;
input x_2525;
input x_2526;
input x_2527;
input x_2528;
input x_2529;
input x_2530;
input x_2531;
input x_2532;
input x_2533;
input x_2534;
input x_2535;
input x_2536;
input x_2537;
input x_2538;
input x_2539;
input x_2540;
input x_2541;
input x_2542;
input x_2543;
input x_2544;
input x_2545;
input x_2546;
input x_2547;
input x_2548;
input x_2549;
input x_2550;
input x_2551;
input x_2552;
input x_2553;
input x_2554;
input x_2555;
input x_2556;
input x_2557;
input x_2558;
input x_2559;
input x_2560;
input x_2561;
input x_2562;
input x_2563;
input x_2564;
input x_2565;
input x_2566;
input x_2567;
input x_2568;
input x_2569;
input x_2570;
input x_2571;
input x_2572;
input x_2573;
input x_2574;
input x_2575;
input x_2576;
input x_2577;
input x_2578;
input x_2579;
input x_2580;
input x_2581;
input x_2582;
input x_2583;
input x_2584;
input x_2585;
input x_2586;
input x_2587;
input x_2588;
input x_2589;
input x_2590;
input x_2591;
input x_2592;
input x_2593;
input x_2594;
input x_2595;
input x_2596;
input x_2597;
input x_2598;
input x_2599;
input x_2600;
input x_2601;
input x_2602;
input x_2603;
input x_2604;
input x_2605;
input x_2606;
input x_2607;
input x_2608;
input x_2609;
input x_2610;
input x_2611;
input x_2612;
input x_2613;
input x_2614;
input x_2615;
input x_2616;
input x_2617;
input x_2618;
input x_2619;
input x_2620;
input x_2621;
input x_2622;
input x_2623;
input x_2624;
input x_2625;
input x_2626;
input x_2627;
input x_2628;
input x_2629;
input x_2630;
input x_2631;
input x_2632;
input x_2633;
input x_2634;
input x_2635;
input x_2636;
input x_2637;
input x_2638;
input x_2639;
input x_2640;
input x_2641;
input x_2642;
input x_2643;
input x_2644;
input x_2645;
input x_2646;
input x_2647;
input x_2648;
input x_2649;
input x_2650;
input x_2651;
input x_2652;
input x_2653;
input x_2654;
input x_2655;
input x_2656;
input x_2657;
input x_2658;
input x_2659;
input x_2660;
input x_2661;
input x_2662;
input x_2663;
input x_2664;
input x_2665;
input x_2666;
input x_2667;
input x_2668;
input x_2669;
input x_2670;
input x_2671;
input x_2672;
input x_2673;
input x_2674;
input x_2675;
input x_2676;
input x_2677;
input x_2678;
input x_2679;
input x_2680;
input x_2681;
input x_2682;
input x_2683;
input x_2684;
input x_2685;
input x_2686;
input x_2687;
input x_2688;
input x_2689;
input x_2690;
input x_2691;
input x_2692;
input x_2693;
input x_2694;
input x_2695;
input x_2696;
input x_2697;
input x_2698;
input x_2699;
input x_2700;
input x_2701;
input x_2702;
input x_2703;
input x_2704;
input x_2705;
input x_2706;
input x_2707;
input x_2708;
input x_2709;
input x_2710;
input x_2711;
input x_2712;
input x_2713;
input x_2714;
input x_2715;
input x_2716;
input x_2717;
input x_2718;
input x_2719;
input x_2720;
input x_2721;
input x_2722;
input x_2723;
input x_2724;
input x_2725;
input x_2726;
input x_2727;
input x_2728;
input x_2729;
input x_2730;
input x_2731;
input x_2732;
input x_2733;
input x_2734;
input x_2735;
input x_2736;
input x_2737;
input x_2738;
input x_2739;
input x_2740;
input x_2741;
input x_2742;
input x_2743;
input x_2744;
input x_2745;
input x_2746;
input x_2747;
input x_2748;
input x_2749;
input x_2750;
input x_2751;
input x_2752;
input x_2753;
input x_2754;
input x_2755;
input x_2756;
input x_2757;
input x_2758;
input x_2759;
input x_2760;
input x_2761;
input x_2762;
input x_2763;
input x_2764;
input x_2765;
input x_2766;
input x_2767;
input x_2768;
input x_2769;
input x_2770;
input x_2771;
input x_2772;
input x_2773;
input x_2774;
input x_2775;
input x_2776;
input x_2777;
input x_2778;
input x_2779;
input x_2780;
input x_2781;
input x_2782;
input x_2783;
input x_2784;
input x_2785;
input x_2786;
input x_2787;
input x_2788;
input x_2789;
input x_2790;
input x_2791;
input x_2792;
input x_2793;
input x_2794;
input x_2795;
input x_2796;
input x_2797;
input x_2798;
input x_2799;
input x_2800;
input x_2801;
input x_2802;
input x_2803;
input x_2804;
input x_2805;
input x_2806;
input x_2807;
input x_2808;
input x_2809;
input x_2810;
input x_2811;
input x_2812;
input x_2813;
input x_2814;
input x_2815;
input x_2816;
input x_2817;
input x_2818;
input x_2819;
input x_2820;
input x_2821;
input x_2822;
input x_2823;
input x_2824;
input x_2825;
input x_2826;
input x_2827;
input x_2828;
input x_2829;
input x_2830;
input x_2831;
input x_2832;
input x_2833;
input x_2834;
input x_2835;
input x_2836;
input x_2837;
input x_2838;
input x_2839;
input x_2840;
input x_2841;
input x_2842;
input x_2843;
input x_2844;
input x_2845;
input x_2846;
input x_2847;
input x_2848;
input x_2849;
input x_2850;
input x_2851;
input x_2852;
input x_2853;
input x_2854;
input x_2855;
input x_2856;
input x_2857;
input x_2858;
input x_2859;
input x_2860;
input x_2861;
input x_2862;
input x_2863;
input x_2864;
input x_2865;
input x_2866;
input x_2867;
input x_2868;
input x_2869;
input x_2870;
input x_2871;
input x_2872;
input x_2873;
input x_2874;
input x_2875;
input x_2876;
input x_2877;
input x_2878;
input x_2879;
input x_2880;
input x_2881;
input x_2882;
input x_2883;
input x_2884;
input x_2885;
input x_2886;
input x_2887;
input x_2888;
input x_2889;
input x_2890;
input x_2891;
input x_2892;
input x_2893;
input x_2894;
input x_2895;
input x_2896;
input x_2897;
input x_2898;
input x_2899;
input x_2900;
input x_2901;
input x_2902;
input x_2903;
input x_2904;
input x_2905;
input x_2906;
input x_2907;
input x_2908;
input x_2909;
input x_2910;
input x_2911;
input x_2912;
input x_2913;
input x_2914;
input x_2915;
input x_2916;
input x_2917;
input x_2918;
input x_2919;
input x_2920;
input x_2921;
input x_2922;
input x_2923;
input x_2924;
input x_2925;
input x_2926;
input x_2927;
input x_2928;
input x_2929;
input x_2930;
input x_2931;
input x_2932;
input x_2933;
input x_2934;
input x_2935;
input x_2936;
input x_2937;
input x_2938;
input x_2939;
input x_2940;
input x_2941;
input x_2942;
input x_2943;
input x_2944;
input x_2945;
input x_2946;
input x_2947;
input x_2948;
input x_2949;
input x_2950;
input x_2951;
input x_2952;
input x_2953;
input x_2954;
input x_2955;
input x_2956;
input x_2957;
input x_2958;
input x_2959;
input x_2960;
input x_2961;
input x_2962;
input x_2963;
input x_2964;
input x_2965;
input x_2966;
input x_2967;
input x_2968;
input x_2969;
input x_2970;
input x_2971;
input x_2972;
input x_2973;
input x_2974;
input x_2975;
input x_2976;
input x_2977;
input x_2978;
input x_2979;
input x_2980;
input x_2981;
input x_2982;
input x_2983;
input x_2984;
input x_2985;
input x_2986;
input x_2987;
input x_2988;
input x_2989;
input x_2990;
input x_2991;
input x_2992;
input x_2993;
input x_2994;
input x_2995;
input x_2996;
input x_2997;
input x_2998;
input x_2999;
input x_3000;
input x_3001;
input x_3002;
input x_3003;
input x_3004;
input x_3005;
input x_3006;
input x_3007;
input x_3008;
input x_3009;
input x_3010;
input x_3011;
input x_3012;
input x_3013;
input x_3014;
input x_3015;
input x_3016;
input x_3017;
input x_3018;
input x_3019;
input x_3020;
input x_3021;
input x_3022;
input x_3023;
input x_3024;
input x_3025;
input x_3026;
input x_3027;
input x_3028;
input x_3029;
input x_3030;
input x_3031;
input x_3032;
input x_3033;
input x_3034;
input x_3035;
input x_3036;
input x_3037;
input x_3038;
input x_3039;
input x_3040;
input x_3041;
input x_3042;
input x_3043;
input x_3044;
input x_3045;
input x_3046;
input x_3047;
input x_3048;
input x_3049;
input x_3050;
input x_3051;
input x_3052;
input x_3053;
input x_3054;
input x_3055;
input x_3056;
input x_3057;
input x_3058;
input x_3059;
input x_3060;
input x_3061;
input x_3062;
input x_3063;
input x_3064;
input x_3065;
input x_3066;
input x_3067;
input x_3068;
input x_3069;
input x_3070;
input x_3071;
input x_3072;
input x_3073;
input x_3074;
input x_3075;
input x_3076;
input x_3077;
input x_3078;
input x_3079;
input x_3080;
input x_3081;
input x_3082;
input x_3083;
input x_3084;
input x_3085;
input x_3086;
input x_3087;
input x_3088;
input x_3089;
input x_3090;
input x_3091;
input x_3092;
input x_3093;
input x_3094;
input x_3095;
input x_3096;
input x_3097;
input x_3098;
input x_3099;
input x_3100;
input x_3101;
input x_3102;
input x_3103;
input x_3104;
input x_3105;
input x_3106;
input x_3107;
input x_3108;
input x_3109;
input x_3110;
input x_3111;
input x_3112;
input x_3113;
input x_3114;
input x_3115;
input x_3116;
input x_3117;
input x_3118;
input x_3119;
input x_3120;
input x_3121;
input x_3122;
input x_3123;
input x_3124;
input x_3125;
input x_3126;
input x_3127;
input x_3128;
input x_3129;
input x_3130;
input x_3131;
input x_3132;
input x_3133;
input x_3134;
input x_3135;
input x_3136;
input x_3137;
input x_3138;
input x_3139;
input x_3140;
input x_3141;
input x_3142;
input x_3143;
input x_3144;
input x_3145;
input x_3146;
input x_3147;
input x_3148;
input x_3149;
input x_3150;
input x_3151;
input x_3152;
input x_3153;
input x_3154;
input x_3155;
input x_3156;
input x_3157;
input x_3158;
input x_3159;
input x_3160;
input x_3161;
input x_3162;
input x_3163;
input x_3164;
input x_3165;
input x_3166;
input x_3167;
input x_3168;
input x_3169;
input x_3170;
input x_3171;
input x_3172;
input x_3173;
input x_3174;
input x_3175;
input x_3176;
input x_3177;
input x_3178;
input x_3179;
input x_3180;
input x_3181;
input x_3182;
input x_3183;
input x_3184;
input x_3185;
input x_3186;
input x_3187;
input x_3188;
input x_3189;
input x_3190;
input x_3191;
input x_3192;
input x_3193;
input x_3194;
input x_3195;
input x_3196;
input x_3197;
input x_3198;
input x_3199;
input x_3200;
input x_3201;
input x_3202;
input x_3203;
input x_3204;
input x_3205;
input x_3206;
input x_3207;
input x_3208;
input x_3209;
input x_3210;
input x_3211;
input x_3212;
input x_3213;
input x_3214;
input x_3215;
input x_3216;
input x_3217;
input x_3218;
input x_3219;
input x_3220;
input x_3221;
input x_3222;
input x_3223;
input x_3224;
input x_3225;
input x_3226;
input x_3227;
input x_3228;
input x_3229;
input x_3230;
input x_3231;
input x_3232;
input x_3233;
input x_3234;
input x_3235;
input x_3236;
input x_3237;
input x_3238;
input x_3239;
input x_3240;
input x_3241;
input x_3242;
input x_3243;
input x_3244;
input x_3245;
input x_3246;
input x_3247;
input x_3248;
input x_3249;
input x_3250;
input x_3251;
input x_3252;
input x_3253;
input x_3254;
input x_3255;
input x_3256;
input x_3257;
input x_3258;
input x_3259;
input x_3260;
input x_3261;
input x_3262;
input x_3263;
input x_3264;
input x_3265;
input x_3266;
input x_3267;
input x_3268;
input x_3269;
input x_3270;
input x_3271;
input x_3272;
input x_3273;
input x_3274;
input x_3275;
input x_3276;
input x_3277;
input x_3278;
input x_3279;
input x_3280;
input x_3281;
input x_3282;
input x_3283;
input x_3284;
input x_3285;
input x_3286;
input x_3287;
input x_3288;
input x_3289;
input x_3290;
input x_3291;
input x_3292;
input x_3293;
input x_3294;
input x_3295;
input x_3296;
input x_3297;
input x_3298;
input x_3299;
input x_3300;
input x_3301;
input x_3302;
input x_3303;
input x_3304;
input x_3305;
input x_3306;
input x_3307;
input x_3308;
input x_3309;
input x_3310;
input x_3311;
input x_3312;
input x_3313;
input x_3314;
input x_3315;
input x_3316;
input x_3317;
input x_3318;
input x_3319;
input x_3320;
input x_3321;
input x_3322;
input x_3323;
input x_3324;
input x_3325;
input x_3326;
input x_3327;
input x_3328;
input x_3329;
input x_3330;
input x_3331;
input x_3332;
input x_3333;
input x_3334;
input x_3335;
input x_3336;
input x_3337;
input x_3338;
input x_3339;
input x_3340;
input x_3341;
input x_3342;
input x_3343;
input x_3344;
input x_3345;
input x_3346;
input x_3347;
input x_3348;
input x_3349;
input x_3350;
input x_3351;
input x_3352;
input x_3353;
input x_3354;
input x_3355;
input x_3356;
input x_3357;
input x_3358;
input x_3359;
input x_3360;
input x_3361;
input x_3362;
input x_3363;
input x_3364;
input x_3365;
input x_3366;
input x_3367;
input x_3368;
input x_3369;
input x_3370;
input x_3371;
input x_3372;
input x_3373;
input x_3374;
input x_3375;
input x_3376;
input x_3377;
input x_3378;
input x_3379;
input x_3380;
input x_3381;
input x_3382;
input x_3383;
input x_3384;
input x_3385;
input x_3386;
input x_3387;
input x_3388;
input x_3389;
input x_3390;
input x_3391;
input x_3392;
input x_3393;
input x_3394;
input x_3395;
input x_3396;
input x_3397;
input x_3398;
input x_3399;
input x_3400;
input x_3401;
input x_3402;
input x_3403;
input x_3404;
input x_3405;
input x_3406;
input x_3407;
input x_3408;
input x_3409;
input x_3410;
input x_3411;
input x_3412;
input x_3413;
input x_3414;
input x_3415;
input x_3416;
input x_3417;
input x_3418;
input x_3419;
input x_3420;
input x_3421;
input x_3422;
input x_3423;
input x_3424;
input x_3425;
input x_3426;
input x_3427;
input x_3428;
input x_3429;
input x_3430;
input x_3431;
input x_3432;
input x_3433;
input x_3434;
input x_3435;
input x_3436;
input x_3437;
input x_3438;
input x_3439;
input x_3440;
input x_3441;
input x_3442;
input x_3443;
input x_3444;
input x_3445;
input x_3446;
input x_3447;
input x_3448;
input x_3449;
input x_3450;
input x_3451;
input x_3452;
input x_3453;
input x_3454;
input x_3455;
input x_3456;
input x_3457;
input x_3458;
input x_3459;
input x_3460;
input x_3461;
input x_3462;
input x_3463;
input x_3464;
input x_3465;
input x_3466;
input x_3467;
input x_3468;
input x_3469;
input x_3470;
input x_3471;
input x_3472;
input x_3473;
input x_3474;
input x_3475;
input x_3476;
input x_3477;
input x_3478;
input x_3479;
input x_3480;
input x_3481;
input x_3482;
input x_3483;
input x_3484;
input x_3485;
input x_3486;
input x_3487;
input x_3488;
input x_3489;
input x_3490;
input x_3491;
input x_3492;
input x_3493;
input x_3494;
input x_3495;
input x_3496;
input x_3497;
input x_3498;
input x_3499;
input x_3500;
input x_3501;
input x_3502;
input x_3503;
input x_3504;
input x_3505;
input x_3506;
input x_3507;
input x_3508;
input x_3509;
input x_3510;
input x_3511;
input x_3512;
input x_3513;
input x_3514;
input x_3515;
input x_3516;
input x_3517;
input x_3518;
input x_3519;
input x_3520;
input x_3521;
input x_3522;
input x_3523;
input x_3524;
input x_3525;
input x_3526;
input x_3527;
input x_3528;
input x_3529;
input x_3530;
input x_3531;
input x_3532;
input x_3533;
input x_3534;
input x_3535;
input x_3536;
input x_3537;
input x_3538;
input x_3539;
input x_3540;
input x_3541;
input x_3542;
input x_3543;
input x_3544;
input x_3545;
input x_3546;
input x_3547;
input x_3548;
input x_3549;
input x_3550;
input x_3551;
input x_3552;
input x_3553;
input x_3554;
input x_3555;
input x_3556;
input x_3557;
input x_3558;
input x_3559;
input x_3560;
input x_3561;
input x_3562;
input x_3563;
input x_3564;
input x_3565;
input x_3566;
input x_3567;
input x_3568;
input x_3569;
input x_3570;
input x_3571;
input x_3572;
input x_3573;
input x_3574;
input x_3575;
input x_3576;
input x_3577;
input x_3578;
input x_3579;
input x_3580;
input x_3581;
input x_3582;
input x_3583;
input x_3584;
input x_3585;
input x_3586;
input x_3587;
input x_3588;
input x_3589;
input x_3590;
input x_3591;
input x_3592;
input x_3593;
input x_3594;
input x_3595;
input x_3596;
input x_3597;
input x_3598;
input x_3599;
input x_3600;
input x_3601;
input x_3602;
input x_3603;
input x_3604;
input x_3605;
input x_3606;
input x_3607;
input x_3608;
input x_3609;
input x_3610;
input x_3611;
input x_3612;
input x_3613;
input x_3614;
input x_3615;
input x_3616;
input x_3617;
input x_3618;
input x_3619;
input x_3620;
input x_3621;
input x_3622;
input x_3623;
input x_3624;
input x_3625;
input x_3626;
input x_3627;
input x_3628;
input x_3629;
input x_3630;
input x_3631;
input x_3632;
input x_3633;
input x_3634;
input x_3635;
input x_3636;
input x_3637;
input x_3638;
input x_3639;
input x_3640;
input x_3641;
input x_3642;
input x_3643;
input x_3644;
input x_3645;
input x_3646;
input x_3647;
input x_3648;
input x_3649;
input x_3650;
input x_3651;
input x_3652;
input x_3653;
input x_3654;
input x_3655;
input x_3656;
input x_3657;
input x_3658;
input x_3659;
input x_3660;
input x_3661;
input x_3662;
input x_3663;
input x_3664;
input x_3665;
input x_3666;
input x_3667;
input x_3668;
input x_3669;
input x_3670;
input x_3671;
input x_3672;
input x_3673;
input x_3674;
input x_3675;
input x_3676;
input x_3677;
input x_3678;
input x_3679;
input x_3680;
input x_3681;
input x_3682;
input x_3683;
input x_3684;
input x_3685;
input x_3686;
input x_3687;
input x_3688;
input x_3689;
input x_3690;
input x_3691;
input x_3692;
input x_3693;
input x_3694;
input x_3695;
input x_3696;
input x_3697;
input x_3698;
input x_3699;
input x_3700;
input x_3701;
input x_3702;
input x_3703;
input x_3704;
input x_3705;
input x_3706;
input x_3707;
input x_3708;
input x_3709;
input x_3710;
input x_3711;
input x_3712;
input x_3713;
input x_3714;
input x_3715;
input x_3716;
input x_3717;
input x_3718;
input x_3719;
input x_3720;
input x_3721;
input x_3722;
input x_3723;
input x_3724;
input x_3725;
input x_3726;
input x_3727;
input x_3728;
input x_3729;
input x_3730;
input x_3731;
input x_3732;
input x_3733;
input x_3734;
input x_3735;
input x_3736;
input x_3737;
input x_3738;
input x_3739;
input x_3740;
input x_3741;
input x_3742;
input x_3743;
input x_3744;
input x_3745;
input x_3746;
input x_3747;
input x_3748;
input x_3749;
input x_3750;
input x_3751;
input x_3752;
input x_3753;
input x_3754;
input x_3755;
input x_3756;
input x_3757;
input x_3758;
input x_3759;
input x_3760;
input x_3761;
input x_3762;
input x_3763;
input x_3764;
input x_3765;
input x_3766;
input x_3767;
input x_3768;
input x_3769;
input x_3770;
input x_3771;
input x_3772;
input x_3773;
input x_3774;
input x_3775;
input x_3776;
input x_3777;
input x_3778;
input x_3779;
input x_3780;
input x_3781;
input x_3782;
input x_3783;
input x_3784;
input x_3785;
input x_3786;
input x_3787;
input x_3788;
input x_3789;
input x_3790;
input x_3791;
input x_3792;
input x_3793;
input x_3794;
input x_3795;
input x_3796;
input x_3797;
input x_3798;
input x_3799;
input x_3800;
input x_3801;
input x_3802;
input x_3803;
input x_3804;
input x_3805;
input x_3806;
input x_3807;
input x_3808;
input x_3809;
input x_3810;
input x_3811;
input x_3812;
input x_3813;
input x_3814;
input x_3815;
input x_3816;
input x_3817;
input x_3818;
input x_3819;
input x_3820;
input x_3821;
input x_3822;
input x_3823;
input x_3824;
input x_3825;
input x_3826;
input x_3827;
input x_3828;
input x_3829;
input x_3830;
input x_3831;
input x_3832;
input x_3833;
input x_3834;
input x_3835;
input x_3836;
input x_3837;
input x_3838;
input x_3839;
input x_3840;
input x_3841;
input x_3842;
input x_3843;
input x_3844;
input x_3845;
input x_3846;
input x_3847;
input x_3848;
input x_3849;
input x_3850;
input x_3851;
input x_3852;
input x_3853;
input x_3854;
input x_3855;
input x_3856;
input x_3857;
input x_3858;
input x_3859;
input x_3860;
input x_3861;
input x_3862;
input x_3863;
input x_3864;
input x_3865;
input x_3866;
input x_3867;
input x_3868;
input x_3869;
input x_3870;
input x_3871;
input x_3872;
input x_3873;
input x_3874;
input x_3875;
input x_3876;
input x_3877;
input x_3878;
input x_3879;
input x_3880;
input x_3881;
input x_3882;
input x_3883;
input x_3884;
input x_3885;
input x_3886;
input x_3887;
input x_3888;
input x_3889;
input x_3890;
input x_3891;
input x_3892;
input x_3893;
input x_3894;
input x_3895;
input x_3896;
input x_3897;
input x_3898;
input x_3899;
input x_3900;
input x_3901;
input x_3902;
input x_3903;
input x_3904;
input x_3905;
input x_3906;
input x_3907;
input x_3908;
input x_3909;
input x_3910;
input x_3911;
input x_3912;
input x_3913;
input x_3914;
input x_3915;
input x_3916;
input x_3917;
input x_3918;
input x_3919;
input x_3920;
input x_3921;
input x_3922;
input x_3923;
input x_3924;
input x_3925;
input x_3926;
input x_3927;
input x_3928;
input x_3929;
input x_3930;
input x_3931;
input x_3932;
input x_3933;
input x_3934;
input x_3935;
input x_3936;
input x_3937;
input x_3938;
input x_3939;
input x_3940;
input x_3941;
input x_3942;
input x_3943;
input x_3944;
input x_3945;
input x_3946;
input x_3947;
input x_3948;
input x_3949;
input x_3950;
input x_3951;
input x_3952;
input x_3953;
input x_3954;
input x_3955;
input x_3956;
input x_3957;
input x_3958;
input x_3959;
input x_3960;
input x_3961;
input x_3962;
input x_3963;
input x_3964;
input x_3965;
input x_3966;
input x_3967;
input x_3968;
input x_3969;
input x_3970;
input x_3971;
input x_3972;
input x_3973;
input x_3974;
input x_3975;
input x_3976;
input x_3977;
input x_3978;
input x_3979;
input x_3980;
input x_3981;
input x_3982;
input x_3983;
input x_3984;
input x_3985;
input x_3986;
input x_3987;
input x_3988;
input x_3989;
input x_3990;
input x_3991;
input x_3992;
input x_3993;
input x_3994;
input x_3995;
input x_3996;
input x_3997;
input x_3998;
input x_3999;
input x_4000;
input x_4001;
input x_4002;
input x_4003;
input x_4004;
input x_4005;
input x_4006;
input x_4007;
input x_4008;
input x_4009;
input x_4010;
input x_4011;
input x_4012;
input x_4013;
input x_4014;
input x_4015;
input x_4016;
input x_4017;
input x_4018;
input x_4019;
input x_4020;
input x_4021;
input x_4022;
input x_4023;
input x_4024;
input x_4025;
input x_4026;
input x_4027;
input x_4028;
input x_4029;
input x_4030;
input x_4031;
input x_4032;
input x_4033;
input x_4034;
input x_4035;
input x_4036;
input x_4037;
input x_4038;
input x_4039;
input x_4040;
input x_4041;
input x_4042;
input x_4043;
input x_4044;
input x_4045;
input x_4046;
input x_4047;
input x_4048;
input x_4049;
input x_4050;
input x_4051;
input x_4052;
input x_4053;
input x_4054;
input x_4055;
input x_4056;
input x_4057;
input x_4058;
input x_4059;
input x_4060;
input x_4061;
input x_4062;
input x_4063;
input x_4064;
input x_4065;
input x_4066;
input x_4067;
input x_4068;
input x_4069;
input x_4070;
input x_4071;
input x_4072;
input x_4073;
input x_4074;
input x_4075;
input x_4076;
input x_4077;
input x_4078;
input x_4079;
input x_4080;
input x_4081;
input x_4082;
input x_4083;
input x_4084;
input x_4085;
input x_4086;
input x_4087;
input x_4088;
input x_4089;
input x_4090;
input x_4091;
input x_4092;
input x_4093;
input x_4094;
input x_4095;
input x_4096;
input x_4097;
input x_4098;
input x_4099;
input x_4100;
input x_4101;
input x_4102;
input x_4103;
input x_4104;
input x_4105;
input x_4106;
input x_4107;
input x_4108;
input x_4109;
input x_4110;
input x_4111;
input x_4112;
input x_4113;
input x_4114;
input x_4115;
input x_4116;
input x_4117;
input x_4118;
input x_4119;
input x_4120;
input x_4121;
input x_4122;
input x_4123;
input x_4124;
input x_4125;
input x_4126;
input x_4127;
input x_4128;
input x_4129;
input x_4130;
input x_4131;
input x_4132;
input x_4133;
input x_4134;
input x_4135;
input x_4136;
input x_4137;
input x_4138;
input x_4139;
input x_4140;
input x_4141;
input x_4142;
input x_4143;
input x_4144;
input x_4145;
input x_4146;
input x_4147;
input x_4148;
input x_4149;
input x_4150;
input x_4151;
input x_4152;
input x_4153;
input x_4154;
input x_4155;
input x_4156;
input x_4157;
input x_4158;
input x_4159;
input x_4160;
input x_4161;
input x_4162;
input x_4163;
input x_4164;
input x_4165;
input x_4166;
input x_4167;
input x_4168;
input x_4169;
input x_4170;
input x_4171;
input x_4172;
input x_4173;
input x_4174;
input x_4175;
input x_4176;
input x_4177;
input x_4178;
input x_4179;
input x_4180;
input x_4181;
input x_4182;
input x_4183;
input x_4184;
input x_4185;
input x_4186;
input x_4187;
input x_4188;
input x_4189;
input x_4190;
input x_4191;
input x_4192;
input x_4193;
input x_4194;
input x_4195;
input x_4196;
input x_4197;
input x_4198;
input x_4199;
input x_4200;
input x_4201;
input x_4202;
input x_4203;
input x_4204;
input x_4205;
input x_4206;
input x_4207;
input x_4208;
input x_4209;
input x_4210;
input x_4211;
input x_4212;
input x_4213;
input x_4214;
input x_4215;
input x_4216;
input x_4217;
input x_4218;
input x_4219;
input x_4220;
input x_4221;
input x_4222;
input x_4223;
input x_4224;
input x_4225;
input x_4226;
input x_4227;
input x_4228;
input x_4229;
input x_4230;
input x_4231;
input x_4232;
input x_4233;
input x_4234;
input x_4235;
input x_4236;
input x_4237;
input x_4238;
input x_4239;
input x_4240;
input x_4241;
input x_4242;
input x_4243;
input x_4244;
input x_4245;
input x_4246;
input x_4247;
input x_4248;
input x_4249;
input x_4250;
input x_4251;
input x_4252;
input x_4253;
input x_4254;
input x_4255;
input x_4256;
input x_4257;
input x_4258;
input x_4259;
input x_4260;
input x_4261;
input x_4262;
input x_4263;
input x_4264;
input x_4265;
input x_4266;
input x_4267;
input x_4268;
input x_4269;
input x_4270;
input x_4271;
input x_4272;
input x_4273;
input x_4274;
input x_4275;
input x_4276;
input x_4277;
input x_4278;
input x_4279;
input x_4280;
input x_4281;
input x_4282;
input x_4283;
input x_4284;
input x_4285;
input x_4286;
input x_4287;
input x_4288;
input x_4289;
input x_4290;
input x_4291;
input x_4292;
input x_4293;
input x_4294;
input x_4295;
input x_4296;
input x_4297;
input x_4298;
input x_4299;
input x_4300;
input x_4301;
input x_4302;
input x_4303;
input x_4304;
input x_4305;
input x_4306;
input x_4307;
input x_4308;
input x_4309;
input x_4310;
input x_4311;
input x_4312;
input x_4313;
input x_4314;
input x_4315;
input x_4316;
input x_4317;
input x_4318;
input x_4319;
input x_4320;
input x_4321;
input x_4322;
input x_4323;
input x_4324;
input x_4325;
input x_4326;
input x_4327;
input x_4328;
input x_4329;
input x_4330;
input x_4331;
input x_4332;
input x_4333;
input x_4334;
input x_4335;
input x_4336;
input x_4337;
input x_4338;
input x_4339;
input x_4340;
input x_4341;
input x_4342;
input x_4343;
input x_4344;
input x_4345;
input x_4346;
input x_4347;
input x_4348;
input x_4349;
input x_4350;
input x_4351;
input x_4352;
input x_4353;
input x_4354;
input x_4355;
input x_4356;
input x_4357;
input x_4358;
input x_4359;
input x_4360;
input x_4361;
input x_4362;
input x_4363;
input x_4364;
input x_4365;
input x_4366;
input x_4367;
input x_4368;
input x_4369;
input x_4370;
input x_4371;
input x_4372;
input x_4373;
input x_4374;
input x_4375;
input x_4376;
input x_4377;
input x_4378;
input x_4379;
input x_4380;
input x_4381;
input x_4382;
input x_4383;
input x_4384;
input x_4385;
input x_4386;
input x_4387;
input x_4388;
input x_4389;
input x_4390;
input x_4391;
input x_4392;
input x_4393;
input x_4394;
input x_4395;
input x_4396;
input x_4397;
input x_4398;
input x_4399;
input x_4400;
input x_4401;
input x_4402;
input x_4403;
input x_4404;
input x_4405;
input x_4406;
input x_4407;
input x_4408;
input x_4409;
input x_4410;
input x_4411;
input x_4412;
input x_4413;
input x_4414;
input x_4415;
input x_4416;
input x_4417;
input x_4418;
input x_4419;
input x_4420;
input x_4421;
input x_4422;
input x_4423;
input x_4424;
input x_4425;
input x_4426;
input x_4427;
input x_4428;
input x_4429;
input x_4430;
input x_4431;
input x_4432;
input x_4433;
input x_4434;
input x_4435;
input x_4436;
input x_4437;
input x_4438;
input x_4439;
input x_4440;
input x_4441;
input x_4442;
input x_4443;
input x_4444;
input x_4445;
input x_4446;
input x_4447;
input x_4448;
input x_4449;
input x_4450;
input x_4451;
input x_4452;
input x_4453;
input x_4454;
input x_4455;
input x_4456;
input x_4457;
input x_4458;
input x_4459;
input x_4460;
input x_4461;
input x_4462;
input x_4463;
input x_4464;
input x_4465;
input x_4466;
input x_4467;
input x_4468;
input x_4469;
input x_4470;
input x_4471;
input x_4472;
input x_4473;
input x_4474;
input x_4475;
input x_4476;
input x_4477;
input x_4478;
input x_4479;
input x_4480;
input x_4481;
input x_4482;
input x_4483;
input x_4484;
input x_4485;
input x_4486;
input x_4487;
input x_4488;
input x_4489;
input x_4490;
input x_4491;
input x_4492;
input x_4493;
input x_4494;
input x_4495;
input x_4496;
input x_4497;
input x_4498;
input x_4499;
input x_4500;
input x_4501;
input x_4502;
input x_4503;
input x_4504;
input x_4505;
input x_4506;
input x_4507;
input x_4508;
input x_4509;
input x_4510;
input x_4511;
input x_4512;
input x_4513;
input x_4514;
input x_4515;
input x_4516;
input x_4517;
input x_4518;
input x_4519;
input x_4520;
input x_4521;
input x_4522;
input x_4523;
input x_4524;
input x_4525;
input x_4526;
input x_4527;
input x_4528;
input x_4529;
input x_4530;
input x_4531;
input x_4532;
input x_4533;
input x_4534;
input x_4535;
input x_4536;
input x_4537;
input x_4538;
input x_4539;
input x_4540;
input x_4541;
input x_4542;
input x_4543;
input x_4544;
input x_4545;
input x_4546;
input x_4547;
input x_4548;
input x_4549;
input x_4550;
input x_4551;
input x_4552;
input x_4553;
input x_4554;
input x_4555;
input x_4556;
input x_4557;
input x_4558;
input x_4559;
input x_4560;
input x_4561;
input x_4562;
input x_4563;
input x_4564;
input x_4565;
input x_4566;
input x_4567;
input x_4568;
input x_4569;
input x_4570;
input x_4571;
input x_4572;
input x_4573;
input x_4574;
input x_4575;
input x_4576;
input x_4577;
input x_4578;
input x_4579;
input x_4580;
input x_4581;
input x_4582;
input x_4583;
input x_4584;
input x_4585;
input x_4586;
input x_4587;
input x_4588;
input x_4589;
input x_4590;
input x_4591;
input x_4592;
input x_4593;
input x_4594;
input x_4595;
input x_4596;
input x_4597;
input x_4598;
input x_4599;
input x_4600;
input x_4601;
input x_4602;
input x_4603;
input x_4604;
input x_4605;
input x_4606;
input x_4607;
input x_4608;
input x_4609;
input x_4610;
input x_4611;
input x_4612;
input x_4613;
input x_4614;
input x_4615;
input x_4616;
input x_4617;
input x_4618;
input x_4619;
input x_4620;
input x_4621;
input x_4622;
input x_4623;
input x_4624;
input x_4625;
input x_4626;
input x_4627;
input x_4628;
input x_4629;
input x_4630;
input x_4631;
input x_4632;
input x_4633;
input x_4634;
input x_4635;
input x_4636;
input x_4637;
input x_4638;
input x_4639;
input x_4640;
input x_4641;
input x_4642;
input x_4643;
input x_4644;
input x_4645;
input x_4646;
input x_4647;
input x_4648;
input x_4649;
input x_4650;
input x_4651;
input x_4652;
input x_4653;
input x_4654;
input x_4655;
input x_4656;
input x_4657;
input x_4658;
input x_4659;
input x_4660;
input x_4661;
input x_4662;
input x_4663;
input x_4664;
input x_4665;
input x_4666;
input x_4667;
input x_4668;
input x_4669;
input x_4670;
input x_4671;
input x_4672;
input x_4673;
input x_4674;
input x_4675;
input x_4676;
input x_4677;
input x_4678;
input x_4679;
input x_4680;
input x_4681;
input x_4682;
input x_4683;
input x_4684;
input x_4685;
input x_4686;
input x_4687;
input x_4688;
input x_4689;
input x_4690;
input x_4691;
input x_4692;
input x_4693;
input x_4694;
input x_4695;
input x_4696;
input x_4697;
input x_4698;
input x_4699;
input x_4700;
input x_4701;
input x_4702;
input x_4703;
input x_4704;
input x_4705;
input x_4706;
input x_4707;
input x_4708;
input x_4709;
input x_4710;
input x_4711;
input x_4712;
input x_4713;
input x_4714;
input x_4715;
input x_4716;
input x_4717;
input x_4718;
input x_4719;
input x_4720;
input x_4721;
input x_4722;
input x_4723;
input x_4724;
input x_4725;
input x_4726;
input x_4727;
input x_4728;
input x_4729;
input x_4730;
input x_4731;
input x_4732;
input x_4733;
input x_4734;
input x_4735;
input x_4736;
input x_4737;
input x_4738;
input x_4739;
input x_4740;
input x_4741;
input x_4742;
input x_4743;
input x_4744;
input x_4745;
input x_4746;
input x_4747;
input x_4748;
input x_4749;
input x_4750;
input x_4751;
input x_4752;
input x_4753;
input x_4754;
input x_4755;
input x_4756;
input x_4757;
input x_4758;
input x_4759;
input x_4760;
input x_4761;
input x_4762;
input x_4763;
input x_4764;
input x_4765;
input x_4766;
input x_4767;
input x_4768;
input x_4769;
input x_4770;
input x_4771;
input x_4772;
input x_4773;
input x_4774;
input x_4775;
input x_4776;
input x_4777;
input x_4778;
input x_4779;
input x_4780;
input x_4781;
input x_4782;
input x_4783;
input x_4784;
input x_4785;
input x_4786;
input x_4787;
input x_4788;
input x_4789;
input x_4790;
input x_4791;
input x_4792;
input x_4793;
input x_4794;
input x_4795;
input x_4796;
input x_4797;
input x_4798;
input x_4799;
input x_4800;
input x_4801;
input x_4802;
input x_4803;
input x_4804;
input x_4805;
input x_4806;
input x_4807;
input x_4808;
input x_4809;
input x_4810;
input x_4811;
input x_4812;
input x_4813;
input x_4814;
input x_4815;
input x_4816;
input x_4817;
input x_4818;
input x_4819;
input x_4820;
input x_4821;
input x_4822;
input x_4823;
input x_4824;
input x_4825;
input x_4826;
input x_4827;
input x_4828;
input x_4829;
input x_4830;
input x_4831;
input x_4832;
input x_4833;
input x_4834;
input x_4835;
input x_4836;
input x_4837;
input x_4838;
input x_4839;
input x_4840;
input x_4841;
input x_4842;
input x_4843;
input x_4844;
input x_4845;
input x_4846;
input x_4847;
input x_4848;
input x_4849;
input x_4850;
input x_4851;
input x_4852;
input x_4853;
input x_4854;
input x_4855;
input x_4856;
input x_4857;
input x_4858;
input x_4859;
input x_4860;
input x_4861;
input x_4862;
input x_4863;
input x_4864;
input x_4865;
input x_4866;
input x_4867;
input x_4868;
input x_4869;
input x_4870;
input x_4871;
input x_4872;
input x_4873;
input x_4874;
input x_4875;
input x_4876;
input x_4877;
input x_4878;
input x_4879;
input x_4880;
input x_4881;
input x_4882;
input x_4883;
input x_4884;
input x_4885;
input x_4886;
input x_4887;
input x_4888;
input x_4889;
input x_4890;
input x_4891;
input x_4892;
input x_4893;
input x_4894;
input x_4895;
input x_4896;
input x_4897;
input x_4898;
input x_4899;
input x_4900;
input x_4901;
input x_4902;
input x_4903;
input x_4904;
input x_4905;
input x_4906;
input x_4907;
input x_4908;
input x_4909;
input x_4910;
input x_4911;
input x_4912;
input x_4913;
input x_4914;
input x_4915;
input x_4916;
input x_4917;
input x_4918;
input x_4919;
input x_4920;
input x_4921;
input x_4922;
input x_4923;
input x_4924;
input x_4925;
input x_4926;
input x_4927;
input x_4928;
input x_4929;
input x_4930;
input x_4931;
input x_4932;
input x_4933;
input x_4934;
input x_4935;
input x_4936;
input x_4937;
input x_4938;
input x_4939;
input x_4940;
input x_4941;
input x_4942;
input x_4943;
input x_4944;
input x_4945;
input x_4946;
input x_4947;
input x_4948;
input x_4949;
input x_4950;
input x_4951;
input x_4952;
input x_4953;
input x_4954;
input x_4955;
input x_4956;
input x_4957;
input x_4958;
input x_4959;
input x_4960;
input x_4961;
input x_4962;
input x_4963;
input x_4964;
input x_4965;
input x_4966;
input x_4967;
input x_4968;
input x_4969;
input x_4970;
input x_4971;
input x_4972;
input x_4973;
input x_4974;
input x_4975;
input x_4976;
input x_4977;
input x_4978;
input x_4979;
input x_4980;
input x_4981;
input x_4982;
input x_4983;
input x_4984;
input x_4985;
input x_4986;
input x_4987;
input x_4988;
input x_4989;
input x_4990;
input x_4991;
input x_4992;
input x_4993;
input x_4994;
input x_4995;
input x_4996;
input x_4997;
input x_4998;
input x_4999;
input x_5000;
input x_5001;
input x_5002;
input x_5003;
input x_5004;
input x_5005;
input x_5006;
input x_5007;
input x_5008;
input x_5009;
input x_5010;
input x_5011;
input x_5012;
input x_5013;
input x_5014;
input x_5015;
input x_5016;
input x_5017;
input x_5018;
input x_5019;
input x_5020;
input x_5021;
input x_5022;
input x_5023;
input x_5024;
input x_5025;
input x_5026;
input x_5027;
input x_5028;
input x_5029;
input x_5030;
input x_5031;
input x_5032;
input x_5033;
input x_5034;
input x_5035;
input x_5036;
input x_5037;
input x_5038;
input x_5039;
input x_5040;
input x_5041;
input x_5042;
input x_5043;
input x_5044;
input x_5045;
input x_5046;
input x_5047;
input x_5048;
input x_5049;
input x_5050;
input x_5051;
input x_5052;
input x_5053;
input x_5054;
input x_5055;
input x_5056;
input x_5057;
input x_5058;
input x_5059;
input x_5060;
input x_5061;
input x_5062;
input x_5063;
input x_5064;
input x_5065;
input x_5066;
input x_5067;
input x_5068;
input x_5069;
input x_5070;
input x_5071;
input x_5072;
input x_5073;
input x_5074;
input x_5075;
input x_5076;
input x_5077;
input x_5078;
input x_5079;
input x_5080;
input x_5081;
input x_5082;
input x_5083;
input x_5084;
input x_5085;
input x_5086;
input x_5087;
input x_5088;
input x_5089;
input x_5090;
input x_5091;
input x_5092;
input x_5093;
input x_5094;
input x_5095;
input x_5096;
input x_5097;
input x_5098;
input x_5099;
input x_5100;
input x_5101;
input x_5102;
input x_5103;
input x_5104;
input x_5105;
input x_5106;
input x_5107;
input x_5108;
input x_5109;
input x_5110;
input x_5111;
input x_5112;
input x_5113;
input x_5114;
input x_5115;
input x_5116;
input x_5117;
input x_5118;
input x_5119;
input x_5120;
input x_5121;
input x_5122;
input x_5123;
input x_5124;
input x_5125;
input x_5126;
input x_5127;
input x_5128;
input x_5129;
input x_5130;
input x_5131;
input x_5132;
input x_5133;
input x_5134;
input x_5135;
input x_5136;
input x_5137;
input x_5138;
input x_5139;
input x_5140;
input x_5141;
input x_5142;
input x_5143;
input x_5144;
input x_5145;
input x_5146;
input x_5147;
input x_5148;
input x_5149;
input x_5150;
input x_5151;
input x_5152;
input x_5153;
input x_5154;
input x_5155;
input x_5156;
input x_5157;
input x_5158;
input x_5159;
input x_5160;
input x_5161;
input x_5162;
input x_5163;
input x_5164;
input x_5165;
input x_5166;
input x_5167;
input x_5168;
input x_5169;
input x_5170;
input x_5171;
input x_5172;
input x_5173;
input x_5174;
input x_5175;
input x_5176;
input x_5177;
input x_5178;
input x_5179;
input x_5180;
input x_5181;
input x_5182;
input x_5183;
input x_5184;
input x_5185;
input x_5186;
input x_5187;
input x_5188;
input x_5189;
input x_5190;
input x_5191;
input x_5192;
input x_5193;
input x_5194;
input x_5195;
input x_5196;
input x_5197;
input x_5198;
input x_5199;
input x_5200;
input x_5201;
input x_5202;
input x_5203;
input x_5204;
input x_5205;
input x_5206;
input x_5207;
input x_5208;
input x_5209;
input x_5210;
input x_5211;
input x_5212;
input x_5213;
input x_5214;
input x_5215;
input x_5216;
input x_5217;
input x_5218;
input x_5219;
input x_5220;
input x_5221;
input x_5222;
input x_5223;
input x_5224;
input x_5225;
input x_5226;
input x_5227;
input x_5228;
input x_5229;
input x_5230;
input x_5231;
input x_5232;
input x_5233;
input x_5234;
input x_5235;
input x_5236;
input x_5237;
input x_5238;
input x_5239;
input x_5240;
input x_5241;
input x_5242;
input x_5243;
input x_5244;
input x_5245;
input x_5246;
input x_5247;
input x_5248;
input x_5249;
input x_5250;
input x_5251;
input x_5252;
input x_5253;
input x_5254;
input x_5255;
input x_5256;
input x_5257;
input x_5258;
input x_5259;
input x_5260;
input x_5261;
input x_5262;
input x_5263;
input x_5264;
input x_5265;
input x_5266;
input x_5267;
input x_5268;
input x_5269;
input x_5270;
input x_5271;
input x_5272;
input x_5273;
input x_5274;
input x_5275;
input x_5276;
input x_5277;
input x_5278;
input x_5279;
input x_5280;
input x_5281;
input x_5282;
input x_5283;
input x_5284;
input x_5285;
input x_5286;
input x_5287;
input x_5288;
input x_5289;
input x_5290;
input x_5291;
input x_5292;
input x_5293;
input x_5294;
input x_5295;
input x_5296;
input x_5297;
input x_5298;
input x_5299;
input x_5300;
input x_5301;
input x_5302;
input x_5303;
input x_5304;
input x_5305;
input x_5306;
input x_5307;
input x_5308;
input x_5309;
input x_5310;
input x_5311;
input x_5312;
input x_5313;
input x_5314;
input x_5315;
input x_5316;
input x_5317;
input x_5318;
input x_5319;
input x_5320;
input x_5321;
input x_5322;
input x_5323;
input x_5324;
input x_5325;
input x_5326;
input x_5327;
input x_5328;
input x_5329;
input x_5330;
input x_5331;
input x_5332;
input x_5333;
input x_5334;
input x_5335;
input x_5336;
input x_5337;
input x_5338;
input x_5339;
input x_5340;
input x_5341;
input x_5342;
input x_5343;
input x_5344;
input x_5345;
input x_5346;
input x_5347;
input x_5348;
input x_5349;
input x_5350;
input x_5351;
input x_5352;
input x_5353;
input x_5354;
input x_5355;
input x_5356;
input x_5357;
input x_5358;
input x_5359;
input x_5360;
input x_5361;
input x_5362;
input x_5363;
input x_5364;
input x_5365;
input x_5366;
input x_5367;
input x_5368;
input x_5369;
input x_5370;
input x_5371;
input x_5372;
input x_5373;
input x_5374;
input x_5375;
input x_5376;
input x_5377;
input x_5378;
input x_5379;
input x_5380;
input x_5381;
input x_5382;
input x_5383;
input x_5384;
input x_5385;
input x_5386;
input x_5387;
input x_5388;
input x_5389;
input x_5390;
input x_5391;
input x_5392;
input x_5393;
input x_5394;
input x_5395;
input x_5396;
input x_5397;
input x_5398;
input x_5399;
input x_5400;
input x_5401;
input x_5402;
input x_5403;
input x_5404;
input x_5405;
input x_5406;
input x_5407;
input x_5408;
input x_5409;
input x_5410;
input x_5411;
input x_5412;
input x_5413;
input x_5414;
input x_5415;
input x_5416;
input x_5417;
input x_5418;
input x_5419;
input x_5420;
input x_5421;
input x_5422;
input x_5423;
input x_5424;
input x_5425;
input x_5426;
input x_5427;
input x_5428;
input x_5429;
input x_5430;
input x_5431;
input x_5432;
input x_5433;
input x_5434;
input x_5435;
input x_5436;
input x_5437;
input x_5438;
input x_5439;
input x_5440;
input x_5441;
input x_5442;
input x_5443;
input x_5444;
input x_5445;
input x_5446;
input x_5447;
input x_5448;
input x_5449;
input x_5450;
input x_5451;
input x_5452;
input x_5453;
input x_5454;
input x_5455;
input x_5456;
input x_5457;
input x_5458;
input x_5459;
input x_5460;
input x_5461;
input x_5462;
input x_5463;
input x_5464;
input x_5465;
input x_5466;
input x_5467;
input x_5468;
input x_5469;
input x_5470;
input x_5471;
input x_5472;
input x_5473;
input x_5474;
input x_5475;
input x_5476;
input x_5477;
input x_5478;
input x_5479;
input x_5480;
input x_5481;
input x_5482;
input x_5483;
input x_5484;
input x_5485;
input x_5486;
input x_5487;
input x_5488;
input x_5489;
input x_5490;
input x_5491;
input x_5492;
input x_5493;
input x_5494;
input x_5495;
input x_5496;
input x_5497;
input x_5498;
input x_5499;
input x_5500;
input x_5501;
input x_5502;
input x_5503;
input x_5504;
input x_5505;
input x_5506;
input x_5507;
input x_5508;
input x_5509;
input x_5510;
input x_5511;
input x_5512;
input x_5513;
input x_5514;
input x_5515;
input x_5516;
input x_5517;
input x_5518;
input x_5519;
input x_5520;
input x_5521;
input x_5522;
input x_5523;
input x_5524;
input x_5525;
input x_5526;
input x_5527;
input x_5528;
input x_5529;
input x_5530;
input x_5531;
input x_5532;
input x_5533;
input x_5534;
input x_5535;
input x_5536;
input x_5537;
input x_5538;
input x_5539;
input x_5540;
input x_5541;
input x_5542;
input x_5543;
input x_5544;
input x_5545;
input x_5546;
input x_5547;
input x_5548;
input x_5549;
input x_5550;
input x_5551;
input x_5552;
input x_5553;
input x_5554;
input x_5555;
input x_5556;
input x_5557;
input x_5558;
input x_5559;
input x_5560;
input x_5561;
input x_5562;
input x_5563;
input x_5564;
input x_5565;
input x_5566;
input x_5567;
input x_5568;
input x_5569;
input x_5570;
input x_5571;
input x_5572;
input x_5573;
input x_5574;
input x_5575;
input x_5576;
input x_5577;
input x_5578;
input x_5579;
input x_5580;
input x_5581;
input x_5582;
input x_5583;
input x_5584;
input x_5585;
input x_5586;
input x_5587;
input x_5588;
input x_5589;
input x_5590;
input x_5591;
input x_5592;
input x_5593;
input x_5594;
input x_5595;
input x_5596;
input x_5597;
input x_5598;
input x_5599;
input x_5600;
input x_5601;
input x_5602;
input x_5603;
input x_5604;
input x_5605;
input x_5606;
input x_5607;
input x_5608;
input x_5609;
input x_5610;
input x_5611;
input x_5612;
input x_5613;
input x_5614;
input x_5615;
input x_5616;
input x_5617;
input x_5618;
input x_5619;
input x_5620;
input x_5621;
input x_5622;
input x_5623;
input x_5624;
input x_5625;
input x_5626;
input x_5627;
input x_5628;
input x_5629;
input x_5630;
input x_5631;
input x_5632;
input x_5633;
input x_5634;
input x_5635;
input x_5636;
input x_5637;
input x_5638;
input x_5639;
input x_5640;
input x_5641;
input x_5642;
input x_5643;
input x_5644;
input x_5645;
input x_5646;
input x_5647;
input x_5648;
input x_5649;
input x_5650;
input x_5651;
input x_5652;
input x_5653;
input x_5654;
input x_5655;
input x_5656;
input x_5657;
input x_5658;
input x_5659;
input x_5660;
input x_5661;
input x_5662;
input x_5663;
input x_5664;
input x_5665;
input x_5666;
input x_5667;
input x_5668;
input x_5669;
input x_5670;
input x_5671;
input x_5672;
input x_5673;
input x_5674;
input x_5675;
input x_5676;
input x_5677;
input x_5678;
input x_5679;
input x_5680;
input x_5681;
input x_5682;
input x_5683;
input x_5684;
input x_5685;
input x_5686;
input x_5687;
input x_5688;
input x_5689;
input x_5690;
input x_5691;
input x_5692;
input x_5693;
input x_5694;
input x_5695;
input x_5696;
input x_5697;
input x_5698;
input x_5699;
input x_5700;
input x_5701;
input x_5702;
input x_5703;
input x_5704;
input x_5705;
input x_5706;
input x_5707;
input x_5708;
input x_5709;
input x_5710;
input x_5711;
input x_5712;
input x_5713;
input x_5714;
input x_5715;
input x_5716;
input x_5717;
input x_5718;
input x_5719;
input x_5720;
input x_5721;
input x_5722;
input x_5723;
input x_5724;
input x_5725;
input x_5726;
input x_5727;
input x_5728;
input x_5729;
input x_5730;
input x_5731;
input x_5732;
input x_5733;
input x_5734;
input x_5735;
input x_5736;
input x_5737;
input x_5738;
input x_5739;
input x_5740;
input x_5741;
input x_5742;
input x_5743;
input x_5744;
input x_5745;
input x_5746;
input x_5747;
input x_5748;
input x_5749;
input x_5750;
input x_5751;
input x_5752;
input x_5753;
input x_5754;
input x_5755;
input x_5756;
input x_5757;
input x_5758;
input x_5759;
input x_5760;
input x_5761;
input x_5762;
input x_5763;
input x_5764;
input x_5765;
input x_5766;
input x_5767;
input x_5768;
input x_5769;
input x_5770;
input x_5771;
input x_5772;
input x_5773;
input x_5774;
input x_5775;
input x_5776;
input x_5777;
input x_5778;
input x_5779;
input x_5780;
input x_5781;
input x_5782;
input x_5783;
input x_5784;
input x_5785;
input x_5786;
input x_5787;
input x_5788;
input x_5789;
input x_5790;
input x_5791;
input x_5792;
input x_5793;
input x_5794;
input x_5795;
input x_5796;
input x_5797;
input x_5798;
input x_5799;
input x_5800;
input x_5801;
input x_5802;
input x_5803;
input x_5804;
input x_5805;
input x_5806;
input x_5807;
input x_5808;
input x_5809;
input x_5810;
input x_5811;
input x_5812;
input x_5813;
input x_5814;
input x_5815;
input x_5816;
input x_5817;
input x_5818;
input x_5819;
input x_5820;
input x_5821;
input x_5822;
input x_5823;
input x_5824;
input x_5825;
input x_5826;
input x_5827;
input x_5828;
input x_5829;
input x_5830;
input x_5831;
input x_5832;
input x_5833;
input x_5834;
input x_5835;
input x_5836;
input x_5837;
input x_5838;
input x_5839;
input x_5840;
input x_5841;
input x_5842;
input x_5843;
input x_5844;
input x_5845;
input x_5846;
input x_5847;
input x_5848;
input x_5849;
input x_5850;
input x_5851;
input x_5852;
input x_5853;
input x_5854;
input x_5855;
input x_5856;
input x_5857;
input x_5858;
input x_5859;
input x_5860;
input x_5861;
input x_5862;
input x_5863;
input x_5864;
input x_5865;
input x_5866;
input x_5867;
input x_5868;
input x_5869;
input x_5870;
input x_5871;
input x_5872;
input x_5873;
input x_5874;
input x_5875;
input x_5876;
input x_5877;
input x_5878;
input x_5879;
input x_5880;
input x_5881;
input x_5882;
input x_5883;
input x_5884;
input x_5885;
input x_5886;
input x_5887;
input x_5888;
input x_5889;
input x_5890;
input x_5891;
input x_5892;
input x_5893;
input x_5894;
input x_5895;
input x_5896;
input x_5897;
input x_5898;
input x_5899;
input x_5900;
input x_5901;
input x_5902;
input x_5903;
input x_5904;
input x_5905;
input x_5906;
input x_5907;
input x_5908;
input x_5909;
input x_5910;
input x_5911;
input x_5912;
input x_5913;
input x_5914;
input x_5915;
input x_5916;
input x_5917;
input x_5918;
input x_5919;
input x_5920;
input x_5921;
input x_5922;
input x_5923;
input x_5924;
input x_5925;
input x_5926;
input x_5927;
input x_5928;
input x_5929;
input x_5930;
input x_5931;
input x_5932;
input x_5933;
input x_5934;
input x_5935;
input x_5936;
input x_5937;
input x_5938;
input x_5939;
input x_5940;
input x_5941;
input x_5942;
input x_5943;
input x_5944;
input x_5945;
input x_5946;
input x_5947;
input x_5948;
input x_5949;
input x_5950;
input x_5951;
input x_5952;
input x_5953;
input x_5954;
input x_5955;
input x_5956;
input x_5957;
input x_5958;
input x_5959;
input x_5960;
input x_5961;
input x_5962;
input x_5963;
input x_5964;
input x_5965;
input x_5966;
input x_5967;
input x_5968;
input x_5969;
input x_5970;
input x_5971;
input x_5972;
input x_5973;
input x_5974;
input x_5975;
input x_5976;
input x_5977;
input x_5978;
input x_5979;
input x_5980;
input x_5981;
input x_5982;
input x_5983;
input x_5984;
input x_5985;
input x_5986;
input x_5987;
input x_5988;
input x_5989;
input x_5990;
input x_5991;
input x_5992;
input x_5993;
input x_5994;
input x_5995;
input x_5996;
input x_5997;
input x_5998;
input x_5999;
input x_6000;
input x_6001;
input x_6002;
input x_6003;
input x_6004;
input x_6005;
input x_6006;
input x_6007;
input x_6008;
input x_6009;
input x_6010;
input x_6011;
input x_6012;
input x_6013;
input x_6014;
input x_6015;
input x_6016;
input x_6017;
input x_6018;
input x_6019;
input x_6020;
input x_6021;
input x_6022;
input x_6023;
input x_6024;
input x_6025;
input x_6026;
input x_6027;
input x_6028;
input x_6029;
input x_6030;
input x_6031;
input x_6032;
input x_6033;
input x_6034;
input x_6035;
input x_6036;
input x_6037;
input x_6038;
input x_6039;
input x_6040;
input x_6041;
input x_6042;
input x_6043;
input x_6044;
input x_6045;
input x_6046;
input x_6047;
input x_6048;
input x_6049;
input x_6050;
input x_6051;
input x_6052;
input x_6053;
input x_6054;
input x_6055;
input x_6056;
input x_6057;
input x_6058;
input x_6059;
input x_6060;
input x_6061;
input x_6062;
input x_6063;
input x_6064;
input x_6065;
input x_6066;
input x_6067;
input x_6068;
input x_6069;
input x_6070;
input x_6071;
input x_6072;
input x_6073;
input x_6074;
input x_6075;
input x_6076;
input x_6077;
input x_6078;
input x_6079;
input x_6080;
input x_6081;
input x_6082;
input x_6083;
input x_6084;
input x_6085;
input x_6086;
input x_6087;
input x_6088;
input x_6089;
input x_6090;
input x_6091;
input x_6092;
input x_6093;
input x_6094;
input x_6095;
input x_6096;
input x_6097;
input x_6098;
input x_6099;
input x_6100;
input x_6101;
input x_6102;
input x_6103;
input x_6104;
input x_6105;
input x_6106;
input x_6107;
input x_6108;
input x_6109;
input x_6110;
input x_6111;
input x_6112;
input x_6113;
input x_6114;
input x_6115;
input x_6116;
input x_6117;
input x_6118;
input x_6119;
input x_6120;
input x_6121;
input x_6122;
input x_6123;
input x_6124;
input x_6125;
input x_6126;
input x_6127;
input x_6128;
input x_6129;
input x_6130;
input x_6131;
input x_6132;
input x_6133;
input x_6134;
input x_6135;
input x_6136;
input x_6137;
input x_6138;
input x_6139;
input x_6140;
input x_6141;
input x_6142;
input x_6143;
input x_6144;
input x_6145;
input x_6146;
input x_6147;
input x_6148;
input x_6149;
input x_6150;
input x_6151;
input x_6152;
input x_6153;
input x_6154;
input x_6155;
input x_6156;
input x_6157;
input x_6158;
input x_6159;
input x_6160;
input x_6161;
input x_6162;
input x_6163;
input x_6164;
input x_6165;
input x_6166;
input x_6167;
input x_6168;
input x_6169;
input x_6170;
input x_6171;
input x_6172;
input x_6173;
input x_6174;
input x_6175;
input x_6176;
input x_6177;
input x_6178;
input x_6179;
input x_6180;
input x_6181;
input x_6182;
input x_6183;
input x_6184;
input x_6185;
input x_6186;
input x_6187;
input x_6188;
input x_6189;
input x_6190;
input x_6191;
input x_6192;
input x_6193;
input x_6194;
input x_6195;
input x_6196;
input x_6197;
input x_6198;
input x_6199;
input x_6200;
input x_6201;
input x_6202;
input x_6203;
input x_6204;
input x_6205;
input x_6206;
input x_6207;
input x_6208;
input x_6209;
input x_6210;
input x_6211;
input x_6212;
input x_6213;
input x_6214;
input x_6215;
input x_6216;
input x_6217;
input x_6218;
input x_6219;
input x_6220;
input x_6221;
input x_6222;
input x_6223;
input x_6224;
input x_6225;
input x_6226;
input x_6227;
input x_6228;
input x_6229;
input x_6230;
input x_6231;
input x_6232;
input x_6233;
input x_6234;
input x_6235;
input x_6236;
input x_6237;
input x_6238;
input x_6239;
input x_6240;
input x_6241;
input x_6242;
input x_6243;
input x_6244;
input x_6245;
input x_6246;
input x_6247;
input x_6248;
input x_6249;
input x_6250;
input x_6251;
input x_6252;
input x_6253;
input x_6254;
output o_1;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire n_53;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_58;
wire n_59;
wire n_60;
wire n_61;
wire n_62;
wire n_63;
wire n_64;
wire n_65;
wire n_66;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;
wire n_95;
wire n_96;
wire n_97;
wire n_98;
wire n_99;
wire n_100;
wire n_101;
wire n_102;
wire n_103;
wire n_104;
wire n_105;
wire n_106;
wire n_107;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_112;
wire n_113;
wire n_114;
wire n_115;
wire n_116;
wire n_117;
wire n_118;
wire n_119;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_124;
wire n_125;
wire n_126;
wire n_127;
wire n_128;
wire n_129;
wire n_130;
wire n_131;
wire n_132;
wire n_133;
wire n_134;
wire n_135;
wire n_136;
wire n_137;
wire n_138;
wire n_139;
wire n_140;
wire n_141;
wire n_142;
wire n_143;
wire n_144;
wire n_145;
wire n_146;
wire n_147;
wire n_148;
wire n_149;
wire n_150;
wire n_151;
wire n_152;
wire n_153;
wire n_154;
wire n_155;
wire n_156;
wire n_157;
wire n_158;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_163;
wire n_164;
wire n_165;
wire n_166;
wire n_167;
wire n_168;
wire n_169;
wire n_170;
wire n_171;
wire n_172;
wire n_173;
wire n_174;
wire n_175;
wire n_176;
wire n_177;
wire n_178;
wire n_179;
wire n_180;
wire n_181;
wire n_182;
wire n_183;
wire n_184;
wire n_185;
wire n_186;
wire n_187;
wire n_188;
wire n_189;
wire n_190;
wire n_191;
wire n_192;
wire n_193;
wire n_194;
wire n_195;
wire n_196;
wire n_197;
wire n_198;
wire n_199;
wire n_200;
wire n_201;
wire n_202;
wire n_203;
wire n_204;
wire n_205;
wire n_206;
wire n_207;
wire n_208;
wire n_209;
wire n_210;
wire n_211;
wire n_212;
wire n_213;
wire n_214;
wire n_215;
wire n_216;
wire n_217;
wire n_218;
wire n_219;
wire n_220;
wire n_221;
wire n_222;
wire n_223;
wire n_224;
wire n_225;
wire n_226;
wire n_227;
wire n_228;
wire n_229;
wire n_230;
wire n_231;
wire n_232;
wire n_233;
wire n_234;
wire n_235;
wire n_236;
wire n_237;
wire n_238;
wire n_239;
wire n_240;
wire n_241;
wire n_242;
wire n_243;
wire n_244;
wire n_245;
wire n_246;
wire n_247;
wire n_248;
wire n_249;
wire n_250;
wire n_251;
wire n_252;
wire n_253;
wire n_254;
wire n_255;
wire n_256;
wire n_257;
wire n_258;
wire n_259;
wire n_260;
wire n_261;
wire n_262;
wire n_263;
wire n_264;
wire n_265;
wire n_266;
wire n_267;
wire n_268;
wire n_269;
wire n_270;
wire n_271;
wire n_272;
wire n_273;
wire n_274;
wire n_275;
wire n_276;
wire n_277;
wire n_278;
wire n_279;
wire n_280;
wire n_281;
wire n_282;
wire n_283;
wire n_284;
wire n_285;
wire n_286;
wire n_287;
wire n_288;
wire n_289;
wire n_290;
wire n_291;
wire n_292;
wire n_293;
wire n_294;
wire n_295;
wire n_296;
wire n_297;
wire n_298;
wire n_299;
wire n_300;
wire n_301;
wire n_302;
wire n_303;
wire n_304;
wire n_305;
wire n_306;
wire n_307;
wire n_308;
wire n_309;
wire n_310;
wire n_311;
wire n_312;
wire n_313;
wire n_314;
wire n_315;
wire n_316;
wire n_317;
wire n_318;
wire n_319;
wire n_320;
wire n_321;
wire n_322;
wire n_323;
wire n_324;
wire n_325;
wire n_326;
wire n_327;
wire n_328;
wire n_329;
wire n_330;
wire n_331;
wire n_332;
wire n_333;
wire n_334;
wire n_335;
wire n_336;
wire n_337;
wire n_338;
wire n_339;
wire n_340;
wire n_341;
wire n_342;
wire n_343;
wire n_344;
wire n_345;
wire n_346;
wire n_347;
wire n_348;
wire n_349;
wire n_350;
wire n_351;
wire n_352;
wire n_353;
wire n_354;
wire n_355;
wire n_356;
wire n_357;
wire n_358;
wire n_359;
wire n_360;
wire n_361;
wire n_362;
wire n_363;
wire n_364;
wire n_365;
wire n_366;
wire n_367;
wire n_368;
wire n_369;
wire n_370;
wire n_371;
wire n_372;
wire n_373;
wire n_374;
wire n_375;
wire n_376;
wire n_377;
wire n_378;
wire n_379;
wire n_380;
wire n_381;
wire n_382;
wire n_383;
wire n_384;
wire n_385;
wire n_386;
wire n_387;
wire n_388;
wire n_389;
wire n_390;
wire n_391;
wire n_392;
wire n_393;
wire n_394;
wire n_395;
wire n_396;
wire n_397;
wire n_398;
wire n_399;
wire n_400;
wire n_401;
wire n_402;
wire n_403;
wire n_404;
wire n_405;
wire n_406;
wire n_407;
wire n_408;
wire n_409;
wire n_410;
wire n_411;
wire n_412;
wire n_413;
wire n_414;
wire n_415;
wire n_416;
wire n_417;
wire n_418;
wire n_419;
wire n_420;
wire n_421;
wire n_422;
wire n_423;
wire n_424;
wire n_425;
wire n_426;
wire n_427;
wire n_428;
wire n_429;
wire n_430;
wire n_431;
wire n_432;
wire n_433;
wire n_434;
wire n_435;
wire n_436;
wire n_437;
wire n_438;
wire n_439;
wire n_440;
wire n_441;
wire n_442;
wire n_443;
wire n_444;
wire n_445;
wire n_446;
wire n_447;
wire n_448;
wire n_449;
wire n_450;
wire n_451;
wire n_452;
wire n_453;
wire n_454;
wire n_455;
wire n_456;
wire n_457;
wire n_458;
wire n_459;
wire n_460;
wire n_461;
wire n_462;
wire n_463;
wire n_464;
wire n_465;
wire n_466;
wire n_467;
wire n_468;
wire n_469;
wire n_470;
wire n_471;
wire n_472;
wire n_473;
wire n_474;
wire n_475;
wire n_476;
wire n_477;
wire n_478;
wire n_479;
wire n_480;
wire n_481;
wire n_482;
wire n_483;
wire n_484;
wire n_485;
wire n_486;
wire n_487;
wire n_488;
wire n_489;
wire n_490;
wire n_491;
wire n_492;
wire n_493;
wire n_494;
wire n_495;
wire n_496;
wire n_497;
wire n_498;
wire n_499;
wire n_500;
wire n_501;
wire n_502;
wire n_503;
wire n_504;
wire n_505;
wire n_506;
wire n_507;
wire n_508;
wire n_509;
wire n_510;
wire n_511;
wire n_512;
wire n_513;
wire n_514;
wire n_515;
wire n_516;
wire n_517;
wire n_518;
wire n_519;
wire n_520;
wire n_521;
wire n_522;
wire n_523;
wire n_524;
wire n_525;
wire n_526;
wire n_527;
wire n_528;
wire n_529;
wire n_530;
wire n_531;
wire n_532;
wire n_533;
wire n_534;
wire n_535;
wire n_536;
wire n_537;
wire n_538;
wire n_539;
wire n_540;
wire n_541;
wire n_542;
wire n_543;
wire n_544;
wire n_545;
wire n_546;
wire n_547;
wire n_548;
wire n_549;
wire n_550;
wire n_551;
wire n_552;
wire n_553;
wire n_554;
wire n_555;
wire n_556;
wire n_557;
wire n_558;
wire n_559;
wire n_560;
wire n_561;
wire n_562;
wire n_563;
wire n_564;
wire n_565;
wire n_566;
wire n_567;
wire n_568;
wire n_569;
wire n_570;
wire n_571;
wire n_572;
wire n_573;
wire n_574;
wire n_575;
wire n_576;
wire n_577;
wire n_578;
wire n_579;
wire n_580;
wire n_581;
wire n_582;
wire n_583;
wire n_584;
wire n_585;
wire n_586;
wire n_587;
wire n_588;
wire n_589;
wire n_590;
wire n_591;
wire n_592;
wire n_593;
wire n_594;
wire n_595;
wire n_596;
wire n_597;
wire n_598;
wire n_599;
wire n_600;
wire n_601;
wire n_602;
wire n_603;
wire n_604;
wire n_605;
wire n_606;
wire n_607;
wire n_608;
wire n_609;
wire n_610;
wire n_611;
wire n_612;
wire n_613;
wire n_614;
wire n_615;
wire n_616;
wire n_617;
wire n_618;
wire n_619;
wire n_620;
wire n_621;
wire n_622;
wire n_623;
wire n_624;
wire n_625;
wire n_626;
wire n_627;
wire n_628;
wire n_629;
wire n_630;
wire n_631;
wire n_632;
wire n_633;
wire n_634;
wire n_635;
wire n_636;
wire n_637;
wire n_638;
wire n_639;
wire n_640;
wire n_641;
wire n_642;
wire n_643;
wire n_644;
wire n_645;
wire n_646;
wire n_647;
wire n_648;
wire n_649;
wire n_650;
wire n_651;
wire n_652;
wire n_653;
wire n_654;
wire n_655;
wire n_656;
wire n_657;
wire n_658;
wire n_659;
wire n_660;
wire n_661;
wire n_662;
wire n_663;
wire n_664;
wire n_665;
wire n_666;
wire n_667;
wire n_668;
wire n_669;
wire n_670;
wire n_671;
wire n_672;
wire n_673;
wire n_674;
wire n_675;
wire n_676;
wire n_677;
wire n_678;
wire n_679;
wire n_680;
wire n_681;
wire n_682;
wire n_683;
wire n_684;
wire n_685;
wire n_686;
wire n_687;
wire n_688;
wire n_689;
wire n_690;
wire n_691;
wire n_692;
wire n_693;
wire n_694;
wire n_695;
wire n_696;
wire n_697;
wire n_698;
wire n_699;
wire n_700;
wire n_701;
wire n_702;
wire n_703;
wire n_704;
wire n_705;
wire n_706;
wire n_707;
wire n_708;
wire n_709;
wire n_710;
wire n_711;
wire n_712;
wire n_713;
wire n_714;
wire n_715;
wire n_716;
wire n_717;
wire n_718;
wire n_719;
wire n_720;
wire n_721;
wire n_722;
wire n_723;
wire n_724;
wire n_725;
wire n_726;
wire n_727;
wire n_728;
wire n_729;
wire n_730;
wire n_731;
wire n_732;
wire n_733;
wire n_734;
wire n_735;
wire n_736;
wire n_737;
wire n_738;
wire n_739;
wire n_740;
wire n_741;
wire n_742;
wire n_743;
wire n_744;
wire n_745;
wire n_746;
wire n_747;
wire n_748;
wire n_749;
wire n_750;
wire n_751;
wire n_752;
wire n_753;
wire n_754;
wire n_755;
wire n_756;
wire n_757;
wire n_758;
wire n_759;
wire n_760;
wire n_761;
wire n_762;
wire n_763;
wire n_764;
wire n_765;
wire n_766;
wire n_767;
wire n_768;
wire n_769;
wire n_770;
wire n_771;
wire n_772;
wire n_773;
wire n_774;
wire n_775;
wire n_776;
wire n_777;
wire n_778;
wire n_779;
wire n_780;
wire n_781;
wire n_782;
wire n_783;
wire n_784;
wire n_785;
wire n_786;
wire n_787;
wire n_788;
wire n_789;
wire n_790;
wire n_791;
wire n_792;
wire n_793;
wire n_794;
wire n_795;
wire n_796;
wire n_797;
wire n_798;
wire n_799;
wire n_800;
wire n_801;
wire n_802;
wire n_803;
wire n_804;
wire n_805;
wire n_806;
wire n_807;
wire n_808;
wire n_809;
wire n_810;
wire n_811;
wire n_812;
wire n_813;
wire n_814;
wire n_815;
wire n_816;
wire n_817;
wire n_818;
wire n_819;
wire n_820;
wire n_821;
wire n_822;
wire n_823;
wire n_824;
wire n_825;
wire n_826;
wire n_827;
wire n_828;
wire n_829;
wire n_830;
wire n_831;
wire n_832;
wire n_833;
wire n_834;
wire n_835;
wire n_836;
wire n_837;
wire n_838;
wire n_839;
wire n_840;
wire n_841;
wire n_842;
wire n_843;
wire n_844;
wire n_845;
wire n_846;
wire n_847;
wire n_848;
wire n_849;
wire n_850;
wire n_851;
wire n_852;
wire n_853;
wire n_854;
wire n_855;
wire n_856;
wire n_857;
wire n_858;
wire n_859;
wire n_860;
wire n_861;
wire n_862;
wire n_863;
wire n_864;
wire n_865;
wire n_866;
wire n_867;
wire n_868;
wire n_869;
wire n_870;
wire n_871;
wire n_872;
wire n_873;
wire n_874;
wire n_875;
wire n_876;
wire n_877;
wire n_878;
wire n_879;
wire n_880;
wire n_881;
wire n_882;
wire n_883;
wire n_884;
wire n_885;
wire n_886;
wire n_887;
wire n_888;
wire n_889;
wire n_890;
wire n_891;
wire n_892;
wire n_893;
wire n_894;
wire n_895;
wire n_896;
wire n_897;
wire n_898;
wire n_899;
wire n_900;
wire n_901;
wire n_902;
wire n_903;
wire n_904;
wire n_905;
wire n_906;
wire n_907;
wire n_908;
wire n_909;
wire n_910;
wire n_911;
wire n_912;
wire n_913;
wire n_914;
wire n_915;
wire n_916;
wire n_917;
wire n_918;
wire n_919;
wire n_920;
wire n_921;
wire n_922;
wire n_923;
wire n_924;
wire n_925;
wire n_926;
wire n_927;
wire n_928;
wire n_929;
wire n_930;
wire n_931;
wire n_932;
wire n_933;
wire n_934;
wire n_935;
wire n_936;
wire n_937;
wire n_938;
wire n_939;
wire n_940;
wire n_941;
wire n_942;
wire n_943;
wire n_944;
wire n_945;
wire n_946;
wire n_947;
wire n_948;
wire n_949;
wire n_950;
wire n_951;
wire n_952;
wire n_953;
wire n_954;
wire n_955;
wire n_956;
wire n_957;
wire n_958;
wire n_959;
wire n_960;
wire n_961;
wire n_962;
wire n_963;
wire n_964;
wire n_965;
wire n_966;
wire n_967;
wire n_968;
wire n_969;
wire n_970;
wire n_971;
wire n_972;
wire n_973;
wire n_974;
wire n_975;
wire n_976;
wire n_977;
wire n_978;
wire n_979;
wire n_980;
wire n_981;
wire n_982;
wire n_983;
wire n_984;
wire n_985;
wire n_986;
wire n_987;
wire n_988;
wire n_989;
wire n_990;
wire n_991;
wire n_992;
wire n_993;
wire n_994;
wire n_995;
wire n_996;
wire n_997;
wire n_998;
wire n_999;
wire n_1000;
wire n_1001;
wire n_1002;
wire n_1003;
wire n_1004;
wire n_1005;
wire n_1006;
wire n_1007;
wire n_1008;
wire n_1009;
wire n_1010;
wire n_1011;
wire n_1012;
wire n_1013;
wire n_1014;
wire n_1015;
wire n_1016;
wire n_1017;
wire n_1018;
wire n_1019;
wire n_1020;
wire n_1021;
wire n_1022;
wire n_1023;
wire n_1024;
wire n_1025;
wire n_1026;
wire n_1027;
wire n_1028;
wire n_1029;
wire n_1030;
wire n_1031;
wire n_1032;
wire n_1033;
wire n_1034;
wire n_1035;
wire n_1036;
wire n_1037;
wire n_1038;
wire n_1039;
wire n_1040;
wire n_1041;
wire n_1042;
wire n_1043;
wire n_1044;
wire n_1045;
wire n_1046;
wire n_1047;
wire n_1048;
wire n_1049;
wire n_1050;
wire n_1051;
wire n_1052;
wire n_1053;
wire n_1054;
wire n_1055;
wire n_1056;
wire n_1057;
wire n_1058;
wire n_1059;
wire n_1060;
wire n_1061;
wire n_1062;
wire n_1063;
wire n_1064;
wire n_1065;
wire n_1066;
wire n_1067;
wire n_1068;
wire n_1069;
wire n_1070;
wire n_1071;
wire n_1072;
wire n_1073;
wire n_1074;
wire n_1075;
wire n_1076;
wire n_1077;
wire n_1078;
wire n_1079;
wire n_1080;
wire n_1081;
wire n_1082;
wire n_1083;
wire n_1084;
wire n_1085;
wire n_1086;
wire n_1087;
wire n_1088;
wire n_1089;
wire n_1090;
wire n_1091;
wire n_1092;
wire n_1093;
wire n_1094;
wire n_1095;
wire n_1096;
wire n_1097;
wire n_1098;
wire n_1099;
wire n_1100;
wire n_1101;
wire n_1102;
wire n_1103;
wire n_1104;
wire n_1105;
wire n_1106;
wire n_1107;
wire n_1108;
wire n_1109;
wire n_1110;
wire n_1111;
wire n_1112;
wire n_1113;
wire n_1114;
wire n_1115;
wire n_1116;
wire n_1117;
wire n_1118;
wire n_1119;
wire n_1120;
wire n_1121;
wire n_1122;
wire n_1123;
wire n_1124;
wire n_1125;
wire n_1126;
wire n_1127;
wire n_1128;
wire n_1129;
wire n_1130;
wire n_1131;
wire n_1132;
wire n_1133;
wire n_1134;
wire n_1135;
wire n_1136;
wire n_1137;
wire n_1138;
wire n_1139;
wire n_1140;
wire n_1141;
wire n_1142;
wire n_1143;
wire n_1144;
wire n_1145;
wire n_1146;
wire n_1147;
wire n_1148;
wire n_1149;
wire n_1150;
wire n_1151;
wire n_1152;
wire n_1153;
wire n_1154;
wire n_1155;
wire n_1156;
wire n_1157;
wire n_1158;
wire n_1159;
wire n_1160;
wire n_1161;
wire n_1162;
wire n_1163;
wire n_1164;
wire n_1165;
wire n_1166;
wire n_1167;
wire n_1168;
wire n_1169;
wire n_1170;
wire n_1171;
wire n_1172;
wire n_1173;
wire n_1174;
wire n_1175;
wire n_1176;
wire n_1177;
wire n_1178;
wire n_1179;
wire n_1180;
wire n_1181;
wire n_1182;
wire n_1183;
wire n_1184;
wire n_1185;
wire n_1186;
wire n_1187;
wire n_1188;
wire n_1189;
wire n_1190;
wire n_1191;
wire n_1192;
wire n_1193;
wire n_1194;
wire n_1195;
wire n_1196;
wire n_1197;
wire n_1198;
wire n_1199;
wire n_1200;
wire n_1201;
wire n_1202;
wire n_1203;
wire n_1204;
wire n_1205;
wire n_1206;
wire n_1207;
wire n_1208;
wire n_1209;
wire n_1210;
wire n_1211;
wire n_1212;
wire n_1213;
wire n_1214;
wire n_1215;
wire n_1216;
wire n_1217;
wire n_1218;
wire n_1219;
wire n_1220;
wire n_1221;
wire n_1222;
wire n_1223;
wire n_1224;
wire n_1225;
wire n_1226;
wire n_1227;
wire n_1228;
wire n_1229;
wire n_1230;
wire n_1231;
wire n_1232;
wire n_1233;
wire n_1234;
wire n_1235;
wire n_1236;
wire n_1237;
wire n_1238;
wire n_1239;
wire n_1240;
wire n_1241;
wire n_1242;
wire n_1243;
wire n_1244;
wire n_1245;
wire n_1246;
wire n_1247;
wire n_1248;
wire n_1249;
wire n_1250;
wire n_1251;
wire n_1252;
wire n_1253;
wire n_1254;
wire n_1255;
wire n_1256;
wire n_1257;
wire n_1258;
wire n_1259;
wire n_1260;
wire n_1261;
wire n_1262;
wire n_1263;
wire n_1264;
wire n_1265;
wire n_1266;
wire n_1267;
wire n_1268;
wire n_1269;
wire n_1270;
wire n_1271;
wire n_1272;
wire n_1273;
wire n_1274;
wire n_1275;
wire n_1276;
wire n_1277;
wire n_1278;
wire n_1279;
wire n_1280;
wire n_1281;
wire n_1282;
wire n_1283;
wire n_1284;
wire n_1285;
wire n_1286;
wire n_1287;
wire n_1288;
wire n_1289;
wire n_1290;
wire n_1291;
wire n_1292;
wire n_1293;
wire n_1294;
wire n_1295;
wire n_1296;
wire n_1297;
wire n_1298;
wire n_1299;
wire n_1300;
wire n_1301;
wire n_1302;
wire n_1303;
wire n_1304;
wire n_1305;
wire n_1306;
wire n_1307;
wire n_1308;
wire n_1309;
wire n_1310;
wire n_1311;
wire n_1312;
wire n_1313;
wire n_1314;
wire n_1315;
wire n_1316;
wire n_1317;
wire n_1318;
wire n_1319;
wire n_1320;
wire n_1321;
wire n_1322;
wire n_1323;
wire n_1324;
wire n_1325;
wire n_1326;
wire n_1327;
wire n_1328;
wire n_1329;
wire n_1330;
wire n_1331;
wire n_1332;
wire n_1333;
wire n_1334;
wire n_1335;
wire n_1336;
wire n_1337;
wire n_1338;
wire n_1339;
wire n_1340;
wire n_1341;
wire n_1342;
wire n_1343;
wire n_1344;
wire n_1345;
wire n_1346;
wire n_1347;
wire n_1348;
wire n_1349;
wire n_1350;
wire n_1351;
wire n_1352;
wire n_1353;
wire n_1354;
wire n_1355;
wire n_1356;
wire n_1357;
wire n_1358;
wire n_1359;
wire n_1360;
wire n_1361;
wire n_1362;
wire n_1363;
wire n_1364;
wire n_1365;
wire n_1366;
wire n_1367;
wire n_1368;
wire n_1369;
wire n_1370;
wire n_1371;
wire n_1372;
wire n_1373;
wire n_1374;
wire n_1375;
wire n_1376;
wire n_1377;
wire n_1378;
wire n_1379;
wire n_1380;
wire n_1381;
wire n_1382;
wire n_1383;
wire n_1384;
wire n_1385;
wire n_1386;
wire n_1387;
wire n_1388;
wire n_1389;
wire n_1390;
wire n_1391;
wire n_1392;
wire n_1393;
wire n_1394;
wire n_1395;
wire n_1396;
wire n_1397;
wire n_1398;
wire n_1399;
wire n_1400;
wire n_1401;
wire n_1402;
wire n_1403;
wire n_1404;
wire n_1405;
wire n_1406;
wire n_1407;
wire n_1408;
wire n_1409;
wire n_1410;
wire n_1411;
wire n_1412;
wire n_1413;
wire n_1414;
wire n_1415;
wire n_1416;
wire n_1417;
wire n_1418;
wire n_1419;
wire n_1420;
wire n_1421;
wire n_1422;
wire n_1423;
wire n_1424;
wire n_1425;
wire n_1426;
wire n_1427;
wire n_1428;
wire n_1429;
wire n_1430;
wire n_1431;
wire n_1432;
wire n_1433;
wire n_1434;
wire n_1435;
wire n_1436;
wire n_1437;
wire n_1438;
wire n_1439;
wire n_1440;
wire n_1441;
wire n_1442;
wire n_1443;
wire n_1444;
wire n_1445;
wire n_1446;
wire n_1447;
wire n_1448;
wire n_1449;
wire n_1450;
wire n_1451;
wire n_1452;
wire n_1453;
wire n_1454;
wire n_1455;
wire n_1456;
wire n_1457;
wire n_1458;
wire n_1459;
wire n_1460;
wire n_1461;
wire n_1462;
wire n_1463;
wire n_1464;
wire n_1465;
wire n_1466;
wire n_1467;
wire n_1468;
wire n_1469;
wire n_1470;
wire n_1471;
wire n_1472;
wire n_1473;
wire n_1474;
wire n_1475;
wire n_1476;
wire n_1477;
wire n_1478;
wire n_1479;
wire n_1480;
wire n_1481;
wire n_1482;
wire n_1483;
wire n_1484;
wire n_1485;
wire n_1486;
wire n_1487;
wire n_1488;
wire n_1489;
wire n_1490;
wire n_1491;
wire n_1492;
wire n_1493;
wire n_1494;
wire n_1495;
wire n_1496;
wire n_1497;
wire n_1498;
wire n_1499;
wire n_1500;
wire n_1501;
wire n_1502;
wire n_1503;
wire n_1504;
wire n_1505;
wire n_1506;
wire n_1507;
wire n_1508;
wire n_1509;
wire n_1510;
wire n_1511;
wire n_1512;
wire n_1513;
wire n_1514;
wire n_1515;
wire n_1516;
wire n_1517;
wire n_1518;
wire n_1519;
wire n_1520;
wire n_1521;
wire n_1522;
wire n_1523;
wire n_1524;
wire n_1525;
wire n_1526;
wire n_1527;
wire n_1528;
wire n_1529;
wire n_1530;
wire n_1531;
wire n_1532;
wire n_1533;
wire n_1534;
wire n_1535;
wire n_1536;
wire n_1537;
wire n_1538;
wire n_1539;
wire n_1540;
wire n_1541;
wire n_1542;
wire n_1543;
wire n_1544;
wire n_1545;
wire n_1546;
wire n_1547;
wire n_1548;
wire n_1549;
wire n_1550;
wire n_1551;
wire n_1552;
wire n_1553;
wire n_1554;
wire n_1555;
wire n_1556;
wire n_1557;
wire n_1558;
wire n_1559;
wire n_1560;
wire n_1561;
wire n_1562;
wire n_1563;
wire n_1564;
wire n_1565;
wire n_1566;
wire n_1567;
wire n_1568;
wire n_1569;
wire n_1570;
wire n_1571;
wire n_1572;
wire n_1573;
wire n_1574;
wire n_1575;
wire n_1576;
wire n_1577;
wire n_1578;
wire n_1579;
wire n_1580;
wire n_1581;
wire n_1582;
wire n_1583;
wire n_1584;
wire n_1585;
wire n_1586;
wire n_1587;
wire n_1588;
wire n_1589;
wire n_1590;
wire n_1591;
wire n_1592;
wire n_1593;
wire n_1594;
wire n_1595;
wire n_1596;
wire n_1597;
wire n_1598;
wire n_1599;
wire n_1600;
wire n_1601;
wire n_1602;
wire n_1603;
wire n_1604;
wire n_1605;
wire n_1606;
wire n_1607;
wire n_1608;
wire n_1609;
wire n_1610;
wire n_1611;
wire n_1612;
wire n_1613;
wire n_1614;
wire n_1615;
wire n_1616;
wire n_1617;
wire n_1618;
wire n_1619;
wire n_1620;
wire n_1621;
wire n_1622;
wire n_1623;
wire n_1624;
wire n_1625;
wire n_1626;
wire n_1627;
wire n_1628;
wire n_1629;
wire n_1630;
wire n_1631;
wire n_1632;
wire n_1633;
wire n_1634;
wire n_1635;
wire n_1636;
wire n_1637;
wire n_1638;
wire n_1639;
wire n_1640;
wire n_1641;
wire n_1642;
wire n_1643;
wire n_1644;
wire n_1645;
wire n_1646;
wire n_1647;
wire n_1648;
wire n_1649;
wire n_1650;
wire n_1651;
wire n_1652;
wire n_1653;
wire n_1654;
wire n_1655;
wire n_1656;
wire n_1657;
wire n_1658;
wire n_1659;
wire n_1660;
wire n_1661;
wire n_1662;
wire n_1663;
wire n_1664;
wire n_1665;
wire n_1666;
wire n_1667;
wire n_1668;
wire n_1669;
wire n_1670;
wire n_1671;
wire n_1672;
wire n_1673;
wire n_1674;
wire n_1675;
wire n_1676;
wire n_1677;
wire n_1678;
wire n_1679;
wire n_1680;
wire n_1681;
wire n_1682;
wire n_1683;
wire n_1684;
wire n_1685;
wire n_1686;
wire n_1687;
wire n_1688;
wire n_1689;
wire n_1690;
wire n_1691;
wire n_1692;
wire n_1693;
wire n_1694;
wire n_1695;
wire n_1696;
wire n_1697;
wire n_1698;
wire n_1699;
wire n_1700;
wire n_1701;
wire n_1702;
wire n_1703;
wire n_1704;
wire n_1705;
wire n_1706;
wire n_1707;
wire n_1708;
wire n_1709;
wire n_1710;
wire n_1711;
wire n_1712;
wire n_1713;
wire n_1714;
wire n_1715;
wire n_1716;
wire n_1717;
wire n_1718;
wire n_1719;
wire n_1720;
wire n_1721;
wire n_1722;
wire n_1723;
wire n_1724;
wire n_1725;
wire n_1726;
wire n_1727;
wire n_1728;
wire n_1729;
wire n_1730;
wire n_1731;
wire n_1732;
wire n_1733;
wire n_1734;
wire n_1735;
wire n_1736;
wire n_1737;
wire n_1738;
wire n_1739;
wire n_1740;
wire n_1741;
wire n_1742;
wire n_1743;
wire n_1744;
wire n_1745;
wire n_1746;
wire n_1747;
wire n_1748;
wire n_1749;
wire n_1750;
wire n_1751;
wire n_1752;
wire n_1753;
wire n_1754;
wire n_1755;
wire n_1756;
wire n_1757;
wire n_1758;
wire n_1759;
wire n_1760;
wire n_1761;
wire n_1762;
wire n_1763;
wire n_1764;
wire n_1765;
wire n_1766;
wire n_1767;
wire n_1768;
wire n_1769;
wire n_1770;
wire n_1771;
wire n_1772;
wire n_1773;
wire n_1774;
wire n_1775;
wire n_1776;
wire n_1777;
wire n_1778;
wire n_1779;
wire n_1780;
wire n_1781;
wire n_1782;
wire n_1783;
wire n_1784;
wire n_1785;
wire n_1786;
wire n_1787;
wire n_1788;
wire n_1789;
wire n_1790;
wire n_1791;
wire n_1792;
wire n_1793;
wire n_1794;
wire n_1795;
wire n_1796;
wire n_1797;
wire n_1798;
wire n_1799;
wire n_1800;
wire n_1801;
wire n_1802;
wire n_1803;
wire n_1804;
wire n_1805;
wire n_1806;
wire n_1807;
wire n_1808;
wire n_1809;
wire n_1810;
wire n_1811;
wire n_1812;
wire n_1813;
wire n_1814;
wire n_1815;
wire n_1816;
wire n_1817;
wire n_1818;
wire n_1819;
wire n_1820;
wire n_1821;
wire n_1822;
wire n_1823;
wire n_1824;
wire n_1825;
wire n_1826;
wire n_1827;
wire n_1828;
wire n_1829;
wire n_1830;
wire n_1831;
wire n_1832;
wire n_1833;
wire n_1834;
wire n_1835;
wire n_1836;
wire n_1837;
wire n_1838;
wire n_1839;
wire n_1840;
wire n_1841;
wire n_1842;
wire n_1843;
wire n_1844;
wire n_1845;
wire n_1846;
wire n_1847;
wire n_1848;
wire n_1849;
wire n_1850;
wire n_1851;
wire n_1852;
wire n_1853;
wire n_1854;
wire n_1855;
wire n_1856;
wire n_1857;
wire n_1858;
wire n_1859;
wire n_1860;
wire n_1861;
wire n_1862;
wire n_1863;
wire n_1864;
wire n_1865;
wire n_1866;
wire n_1867;
wire n_1868;
wire n_1869;
wire n_1870;
wire n_1871;
wire n_1872;
wire n_1873;
wire n_1874;
wire n_1875;
wire n_1876;
wire n_1877;
wire n_1878;
wire n_1879;
wire n_1880;
wire n_1881;
wire n_1882;
wire n_1883;
wire n_1884;
wire n_1885;
wire n_1886;
wire n_1887;
wire n_1888;
wire n_1889;
wire n_1890;
wire n_1891;
wire n_1892;
wire n_1893;
wire n_1894;
wire n_1895;
wire n_1896;
wire n_1897;
wire n_1898;
wire n_1899;
wire n_1900;
wire n_1901;
wire n_1902;
wire n_1903;
wire n_1904;
wire n_1905;
wire n_1906;
wire n_1907;
wire n_1908;
wire n_1909;
wire n_1910;
wire n_1911;
wire n_1912;
wire n_1913;
wire n_1914;
wire n_1915;
wire n_1916;
wire n_1917;
wire n_1918;
wire n_1919;
wire n_1920;
wire n_1921;
wire n_1922;
wire n_1923;
wire n_1924;
wire n_1925;
wire n_1926;
wire n_1927;
wire n_1928;
wire n_1929;
wire n_1930;
wire n_1931;
wire n_1932;
wire n_1933;
wire n_1934;
wire n_1935;
wire n_1936;
wire n_1937;
wire n_1938;
wire n_1939;
wire n_1940;
wire n_1941;
wire n_1942;
wire n_1943;
wire n_1944;
wire n_1945;
wire n_1946;
wire n_1947;
wire n_1948;
wire n_1949;
wire n_1950;
wire n_1951;
wire n_1952;
wire n_1953;
wire n_1954;
wire n_1955;
wire n_1956;
wire n_1957;
wire n_1958;
wire n_1959;
wire n_1960;
wire n_1961;
wire n_1962;
wire n_1963;
wire n_1964;
wire n_1965;
wire n_1966;
wire n_1967;
wire n_1968;
wire n_1969;
wire n_1970;
wire n_1971;
wire n_1972;
wire n_1973;
wire n_1974;
wire n_1975;
wire n_1976;
wire n_1977;
wire n_1978;
wire n_1979;
wire n_1980;
wire n_1981;
wire n_1982;
wire n_1983;
wire n_1984;
wire n_1985;
wire n_1986;
wire n_1987;
wire n_1988;
wire n_1989;
wire n_1990;
wire n_1991;
wire n_1992;
wire n_1993;
wire n_1994;
wire n_1995;
wire n_1996;
wire n_1997;
wire n_1998;
wire n_1999;
wire n_2000;
wire n_2001;
wire n_2002;
wire n_2003;
wire n_2004;
wire n_2005;
wire n_2006;
wire n_2007;
wire n_2008;
wire n_2009;
wire n_2010;
wire n_2011;
wire n_2012;
wire n_2013;
wire n_2014;
wire n_2015;
wire n_2016;
wire n_2017;
wire n_2018;
wire n_2019;
wire n_2020;
wire n_2021;
wire n_2022;
wire n_2023;
wire n_2024;
wire n_2025;
wire n_2026;
wire n_2027;
wire n_2028;
wire n_2029;
wire n_2030;
wire n_2031;
wire n_2032;
wire n_2033;
wire n_2034;
wire n_2035;
wire n_2036;
wire n_2037;
wire n_2038;
wire n_2039;
wire n_2040;
wire n_2041;
wire n_2042;
wire n_2043;
wire n_2044;
wire n_2045;
wire n_2046;
wire n_2047;
wire n_2048;
wire n_2049;
wire n_2050;
wire n_2051;
wire n_2052;
wire n_2053;
wire n_2054;
wire n_2055;
wire n_2056;
wire n_2057;
wire n_2058;
wire n_2059;
wire n_2060;
wire n_2061;
wire n_2062;
wire n_2063;
wire n_2064;
wire n_2065;
wire n_2066;
wire n_2067;
wire n_2068;
wire n_2069;
wire n_2070;
wire n_2071;
wire n_2072;
wire n_2073;
wire n_2074;
wire n_2075;
wire n_2076;
wire n_2077;
wire n_2078;
wire n_2079;
wire n_2080;
wire n_2081;
wire n_2082;
wire n_2083;
wire n_2084;
wire n_2085;
wire n_2086;
wire n_2087;
wire n_2088;
wire n_2089;
wire n_2090;
wire n_2091;
wire n_2092;
wire n_2093;
wire n_2094;
wire n_2095;
wire n_2096;
wire n_2097;
wire n_2098;
wire n_2099;
wire n_2100;
wire n_2101;
wire n_2102;
wire n_2103;
wire n_2104;
wire n_2105;
wire n_2106;
wire n_2107;
wire n_2108;
wire n_2109;
wire n_2110;
wire n_2111;
wire n_2112;
wire n_2113;
wire n_2114;
wire n_2115;
wire n_2116;
wire n_2117;
wire n_2118;
wire n_2119;
wire n_2120;
wire n_2121;
wire n_2122;
wire n_2123;
wire n_2124;
wire n_2125;
wire n_2126;
wire n_2127;
wire n_2128;
wire n_2129;
wire n_2130;
wire n_2131;
wire n_2132;
wire n_2133;
wire n_2134;
wire n_2135;
wire n_2136;
wire n_2137;
wire n_2138;
wire n_2139;
wire n_2140;
wire n_2141;
wire n_2142;
wire n_2143;
wire n_2144;
wire n_2145;
wire n_2146;
wire n_2147;
wire n_2148;
wire n_2149;
wire n_2150;
wire n_2151;
wire n_2152;
wire n_2153;
wire n_2154;
wire n_2155;
wire n_2156;
wire n_2157;
wire n_2158;
wire n_2159;
wire n_2160;
wire n_2161;
wire n_2162;
wire n_2163;
wire n_2164;
wire n_2165;
wire n_2166;
wire n_2167;
wire n_2168;
wire n_2169;
wire n_2170;
wire n_2171;
wire n_2172;
wire n_2173;
wire n_2174;
wire n_2175;
wire n_2176;
wire n_2177;
wire n_2178;
wire n_2179;
wire n_2180;
wire n_2181;
wire n_2182;
wire n_2183;
wire n_2184;
wire n_2185;
wire n_2186;
wire n_2187;
wire n_2188;
wire n_2189;
wire n_2190;
wire n_2191;
wire n_2192;
wire n_2193;
wire n_2194;
wire n_2195;
wire n_2196;
wire n_2197;
wire n_2198;
wire n_2199;
wire n_2200;
wire n_2201;
wire n_2202;
wire n_2203;
wire n_2204;
wire n_2205;
wire n_2206;
wire n_2207;
wire n_2208;
wire n_2209;
wire n_2210;
wire n_2211;
wire n_2212;
wire n_2213;
wire n_2214;
wire n_2215;
wire n_2216;
wire n_2217;
wire n_2218;
wire n_2219;
wire n_2220;
wire n_2221;
wire n_2222;
wire n_2223;
wire n_2224;
wire n_2225;
wire n_2226;
wire n_2227;
wire n_2228;
wire n_2229;
wire n_2230;
wire n_2231;
wire n_2232;
wire n_2233;
wire n_2234;
wire n_2235;
wire n_2236;
wire n_2237;
wire n_2238;
wire n_2239;
wire n_2240;
wire n_2241;
wire n_2242;
wire n_2243;
wire n_2244;
wire n_2245;
wire n_2246;
wire n_2247;
wire n_2248;
wire n_2249;
wire n_2250;
wire n_2251;
wire n_2252;
wire n_2253;
wire n_2254;
wire n_2255;
wire n_2256;
wire n_2257;
wire n_2258;
wire n_2259;
wire n_2260;
wire n_2261;
wire n_2262;
wire n_2263;
wire n_2264;
wire n_2265;
wire n_2266;
wire n_2267;
wire n_2268;
wire n_2269;
wire n_2270;
wire n_2271;
wire n_2272;
wire n_2273;
wire n_2274;
wire n_2275;
wire n_2276;
wire n_2277;
wire n_2278;
wire n_2279;
wire n_2280;
wire n_2281;
wire n_2282;
wire n_2283;
wire n_2284;
wire n_2285;
wire n_2286;
wire n_2287;
wire n_2288;
wire n_2289;
wire n_2290;
wire n_2291;
wire n_2292;
wire n_2293;
wire n_2294;
wire n_2295;
wire n_2296;
wire n_2297;
wire n_2298;
wire n_2299;
wire n_2300;
wire n_2301;
wire n_2302;
wire n_2303;
wire n_2304;
wire n_2305;
wire n_2306;
wire n_2307;
wire n_2308;
wire n_2309;
wire n_2310;
wire n_2311;
wire n_2312;
wire n_2313;
wire n_2314;
wire n_2315;
wire n_2316;
wire n_2317;
wire n_2318;
wire n_2319;
wire n_2320;
wire n_2321;
wire n_2322;
wire n_2323;
wire n_2324;
wire n_2325;
wire n_2326;
wire n_2327;
wire n_2328;
wire n_2329;
wire n_2330;
wire n_2331;
wire n_2332;
wire n_2333;
wire n_2334;
wire n_2335;
wire n_2336;
wire n_2337;
wire n_2338;
wire n_2339;
wire n_2340;
wire n_2341;
wire n_2342;
wire n_2343;
wire n_2344;
wire n_2345;
wire n_2346;
wire n_2347;
wire n_2348;
wire n_2349;
wire n_2350;
wire n_2351;
wire n_2352;
wire n_2353;
wire n_2354;
wire n_2355;
wire n_2356;
wire n_2357;
wire n_2358;
wire n_2359;
wire n_2360;
wire n_2361;
wire n_2362;
wire n_2363;
wire n_2364;
wire n_2365;
wire n_2366;
wire n_2367;
wire n_2368;
wire n_2369;
wire n_2370;
wire n_2371;
wire n_2372;
wire n_2373;
wire n_2374;
wire n_2375;
wire n_2376;
wire n_2377;
wire n_2378;
wire n_2379;
wire n_2380;
wire n_2381;
wire n_2382;
wire n_2383;
wire n_2384;
wire n_2385;
wire n_2386;
wire n_2387;
wire n_2388;
wire n_2389;
wire n_2390;
wire n_2391;
wire n_2392;
wire n_2393;
wire n_2394;
wire n_2395;
wire n_2396;
wire n_2397;
wire n_2398;
wire n_2399;
wire n_2400;
wire n_2401;
wire n_2402;
wire n_2403;
wire n_2404;
wire n_2405;
wire n_2406;
wire n_2407;
wire n_2408;
wire n_2409;
wire n_2410;
wire n_2411;
wire n_2412;
wire n_2413;
wire n_2414;
wire n_2415;
wire n_2416;
wire n_2417;
wire n_2418;
wire n_2419;
wire n_2420;
wire n_2421;
wire n_2422;
wire n_2423;
wire n_2424;
wire n_2425;
wire n_2426;
wire n_2427;
wire n_2428;
wire n_2429;
wire n_2430;
wire n_2431;
wire n_2432;
wire n_2433;
wire n_2434;
wire n_2435;
wire n_2436;
wire n_2437;
wire n_2438;
wire n_2439;
wire n_2440;
wire n_2441;
wire n_2442;
wire n_2443;
wire n_2444;
wire n_2445;
wire n_2446;
wire n_2447;
wire n_2448;
wire n_2449;
wire n_2450;
wire n_2451;
wire n_2452;
wire n_2453;
wire n_2454;
wire n_2455;
wire n_2456;
wire n_2457;
wire n_2458;
wire n_2459;
wire n_2460;
wire n_2461;
wire n_2462;
wire n_2463;
wire n_2464;
wire n_2465;
wire n_2466;
wire n_2467;
wire n_2468;
wire n_2469;
wire n_2470;
wire n_2471;
wire n_2472;
wire n_2473;
wire n_2474;
wire n_2475;
wire n_2476;
wire n_2477;
wire n_2478;
wire n_2479;
wire n_2480;
wire n_2481;
wire n_2482;
wire n_2483;
wire n_2484;
wire n_2485;
wire n_2486;
wire n_2487;
wire n_2488;
wire n_2489;
wire n_2490;
wire n_2491;
wire n_2492;
wire n_2493;
wire n_2494;
wire n_2495;
wire n_2496;
wire n_2497;
wire n_2498;
wire n_2499;
wire n_2500;
wire n_2501;
wire n_2502;
wire n_2503;
wire n_2504;
wire n_2505;
wire n_2506;
wire n_2507;
wire n_2508;
wire n_2509;
wire n_2510;
wire n_2511;
wire n_2512;
wire n_2513;
wire n_2514;
wire n_2515;
wire n_2516;
wire n_2517;
wire n_2518;
wire n_2519;
wire n_2520;
wire n_2521;
wire n_2522;
wire n_2523;
wire n_2524;
wire n_2525;
wire n_2526;
wire n_2527;
wire n_2528;
wire n_2529;
wire n_2530;
wire n_2531;
wire n_2532;
wire n_2533;
wire n_2534;
wire n_2535;
wire n_2536;
wire n_2537;
wire n_2538;
wire n_2539;
wire n_2540;
wire n_2541;
wire n_2542;
wire n_2543;
wire n_2544;
wire n_2545;
wire n_2546;
wire n_2547;
wire n_2548;
wire n_2549;
wire n_2550;
wire n_2551;
wire n_2552;
wire n_2553;
wire n_2554;
wire n_2555;
wire n_2556;
wire n_2557;
wire n_2558;
wire n_2559;
wire n_2560;
wire n_2561;
wire n_2562;
wire n_2563;
wire n_2564;
wire n_2565;
wire n_2566;
wire n_2567;
wire n_2568;
wire n_2569;
wire n_2570;
wire n_2571;
wire n_2572;
wire n_2573;
wire n_2574;
wire n_2575;
wire n_2576;
wire n_2577;
wire n_2578;
wire n_2579;
wire n_2580;
wire n_2581;
wire n_2582;
wire n_2583;
wire n_2584;
wire n_2585;
wire n_2586;
wire n_2587;
wire n_2588;
wire n_2589;
wire n_2590;
wire n_2591;
wire n_2592;
wire n_2593;
wire n_2594;
wire n_2595;
wire n_2596;
wire n_2597;
wire n_2598;
wire n_2599;
wire n_2600;
wire n_2601;
wire n_2602;
wire n_2603;
wire n_2604;
wire n_2605;
wire n_2606;
wire n_2607;
wire n_2608;
wire n_2609;
wire n_2610;
wire n_2611;
wire n_2612;
wire n_2613;
wire n_2614;
wire n_2615;
wire n_2616;
wire n_2617;
wire n_2618;
wire n_2619;
wire n_2620;
wire n_2621;
wire n_2622;
wire n_2623;
wire n_2624;
wire n_2625;
wire n_2626;
wire n_2627;
wire n_2628;
wire n_2629;
wire n_2630;
wire n_2631;
wire n_2632;
wire n_2633;
wire n_2634;
wire n_2635;
wire n_2636;
wire n_2637;
wire n_2638;
wire n_2639;
wire n_2640;
wire n_2641;
wire n_2642;
wire n_2643;
wire n_2644;
wire n_2645;
wire n_2646;
wire n_2647;
wire n_2648;
wire n_2649;
wire n_2650;
wire n_2651;
wire n_2652;
wire n_2653;
wire n_2654;
wire n_2655;
wire n_2656;
wire n_2657;
wire n_2658;
wire n_2659;
wire n_2660;
wire n_2661;
wire n_2662;
wire n_2663;
wire n_2664;
wire n_2665;
wire n_2666;
wire n_2667;
wire n_2668;
wire n_2669;
wire n_2670;
wire n_2671;
wire n_2672;
wire n_2673;
wire n_2674;
wire n_2675;
wire n_2676;
wire n_2677;
wire n_2678;
wire n_2679;
wire n_2680;
wire n_2681;
wire n_2682;
wire n_2683;
wire n_2684;
wire n_2685;
wire n_2686;
wire n_2687;
wire n_2688;
wire n_2689;
wire n_2690;
wire n_2691;
wire n_2692;
wire n_2693;
wire n_2694;
wire n_2695;
wire n_2696;
wire n_2697;
wire n_2698;
wire n_2699;
wire n_2700;
wire n_2701;
wire n_2702;
wire n_2703;
wire n_2704;
wire n_2705;
wire n_2706;
wire n_2707;
wire n_2708;
wire n_2709;
wire n_2710;
wire n_2711;
wire n_2712;
wire n_2713;
wire n_2714;
wire n_2715;
wire n_2716;
wire n_2717;
wire n_2718;
wire n_2719;
wire n_2720;
wire n_2721;
wire n_2722;
wire n_2723;
wire n_2724;
wire n_2725;
wire n_2726;
wire n_2727;
wire n_2728;
wire n_2729;
wire n_2730;
wire n_2731;
wire n_2732;
wire n_2733;
wire n_2734;
wire n_2735;
wire n_2736;
wire n_2737;
wire n_2738;
wire n_2739;
wire n_2740;
wire n_2741;
wire n_2742;
wire n_2743;
wire n_2744;
wire n_2745;
wire n_2746;
wire n_2747;
wire n_2748;
wire n_2749;
wire n_2750;
wire n_2751;
wire n_2752;
wire n_2753;
wire n_2754;
wire n_2755;
wire n_2756;
wire n_2757;
wire n_2758;
wire n_2759;
wire n_2760;
wire n_2761;
wire n_2762;
wire n_2763;
wire n_2764;
wire n_2765;
wire n_2766;
wire n_2767;
wire n_2768;
wire n_2769;
wire n_2770;
wire n_2771;
wire n_2772;
wire n_2773;
wire n_2774;
wire n_2775;
wire n_2776;
wire n_2777;
wire n_2778;
wire n_2779;
wire n_2780;
wire n_2781;
wire n_2782;
wire n_2783;
wire n_2784;
wire n_2785;
wire n_2786;
wire n_2787;
wire n_2788;
wire n_2789;
wire n_2790;
wire n_2791;
wire n_2792;
wire n_2793;
wire n_2794;
wire n_2795;
wire n_2796;
wire n_2797;
wire n_2798;
wire n_2799;
wire n_2800;
wire n_2801;
wire n_2802;
wire n_2803;
wire n_2804;
wire n_2805;
wire n_2806;
wire n_2807;
wire n_2808;
wire n_2809;
wire n_2810;
wire n_2811;
wire n_2812;
wire n_2813;
wire n_2814;
wire n_2815;
wire n_2816;
wire n_2817;
wire n_2818;
wire n_2819;
wire n_2820;
wire n_2821;
wire n_2822;
wire n_2823;
wire n_2824;
wire n_2825;
wire n_2826;
wire n_2827;
wire n_2828;
wire n_2829;
wire n_2830;
wire n_2831;
wire n_2832;
wire n_2833;
wire n_2834;
wire n_2835;
wire n_2836;
wire n_2837;
wire n_2838;
wire n_2839;
wire n_2840;
wire n_2841;
wire n_2842;
wire n_2843;
wire n_2844;
wire n_2845;
wire n_2846;
wire n_2847;
wire n_2848;
wire n_2849;
wire n_2850;
wire n_2851;
wire n_2852;
wire n_2853;
wire n_2854;
wire n_2855;
wire n_2856;
wire n_2857;
wire n_2858;
wire n_2859;
wire n_2860;
wire n_2861;
wire n_2862;
wire n_2863;
wire n_2864;
wire n_2865;
wire n_2866;
wire n_2867;
wire n_2868;
wire n_2869;
wire n_2870;
wire n_2871;
wire n_2872;
wire n_2873;
wire n_2874;
wire n_2875;
wire n_2876;
wire n_2877;
wire n_2878;
wire n_2879;
wire n_2880;
wire n_2881;
wire n_2882;
wire n_2883;
wire n_2884;
wire n_2885;
wire n_2886;
wire n_2887;
wire n_2888;
wire n_2889;
wire n_2890;
wire n_2891;
wire n_2892;
wire n_2893;
wire n_2894;
wire n_2895;
wire n_2896;
wire n_2897;
wire n_2898;
wire n_2899;
wire n_2900;
wire n_2901;
wire n_2902;
wire n_2903;
wire n_2904;
wire n_2905;
wire n_2906;
wire n_2907;
wire n_2908;
wire n_2909;
wire n_2910;
wire n_2911;
wire n_2912;
wire n_2913;
wire n_2914;
wire n_2915;
wire n_2916;
wire n_2917;
wire n_2918;
wire n_2919;
wire n_2920;
wire n_2921;
wire n_2922;
wire n_2923;
wire n_2924;
wire n_2925;
wire n_2926;
wire n_2927;
wire n_2928;
wire n_2929;
wire n_2930;
wire n_2931;
wire n_2932;
wire n_2933;
wire n_2934;
wire n_2935;
wire n_2936;
wire n_2937;
wire n_2938;
wire n_2939;
wire n_2940;
wire n_2941;
wire n_2942;
wire n_2943;
wire n_2944;
wire n_2945;
wire n_2946;
wire n_2947;
wire n_2948;
wire n_2949;
wire n_2950;
wire n_2951;
wire n_2952;
wire n_2953;
wire n_2954;
wire n_2955;
wire n_2956;
wire n_2957;
wire n_2958;
wire n_2959;
wire n_2960;
wire n_2961;
wire n_2962;
wire n_2963;
wire n_2964;
wire n_2965;
wire n_2966;
wire n_2967;
wire n_2968;
wire n_2969;
wire n_2970;
wire n_2971;
wire n_2972;
wire n_2973;
wire n_2974;
wire n_2975;
wire n_2976;
wire n_2977;
wire n_2978;
wire n_2979;
wire n_2980;
wire n_2981;
wire n_2982;
wire n_2983;
wire n_2984;
wire n_2985;
wire n_2986;
wire n_2987;
wire n_2988;
wire n_2989;
wire n_2990;
wire n_2991;
wire n_2992;
wire n_2993;
wire n_2994;
wire n_2995;
wire n_2996;
wire n_2997;
wire n_2998;
wire n_2999;
wire n_3000;
wire n_3001;
wire n_3002;
wire n_3003;
wire n_3004;
wire n_3005;
wire n_3006;
wire n_3007;
wire n_3008;
wire n_3009;
wire n_3010;
wire n_3011;
wire n_3012;
wire n_3013;
wire n_3014;
wire n_3015;
wire n_3016;
wire n_3017;
wire n_3018;
wire n_3019;
wire n_3020;
wire n_3021;
wire n_3022;
wire n_3023;
wire n_3024;
wire n_3025;
wire n_3026;
wire n_3027;
wire n_3028;
wire n_3029;
wire n_3030;
wire n_3031;
wire n_3032;
wire n_3033;
wire n_3034;
wire n_3035;
wire n_3036;
wire n_3037;
wire n_3038;
wire n_3039;
wire n_3040;
wire n_3041;
wire n_3042;
wire n_3043;
wire n_3044;
wire n_3045;
wire n_3046;
wire n_3047;
wire n_3048;
wire n_3049;
wire n_3050;
wire n_3051;
wire n_3052;
wire n_3053;
wire n_3054;
wire n_3055;
wire n_3056;
wire n_3057;
wire n_3058;
wire n_3059;
wire n_3060;
wire n_3061;
wire n_3062;
wire n_3063;
wire n_3064;
wire n_3065;
wire n_3066;
wire n_3067;
wire n_3068;
wire n_3069;
wire n_3070;
wire n_3071;
wire n_3072;
wire n_3073;
wire n_3074;
wire n_3075;
wire n_3076;
wire n_3077;
wire n_3078;
wire n_3079;
wire n_3080;
wire n_3081;
wire n_3082;
wire n_3083;
wire n_3084;
wire n_3085;
wire n_3086;
wire n_3087;
wire n_3088;
wire n_3089;
wire n_3090;
wire n_3091;
wire n_3092;
wire n_3093;
wire n_3094;
wire n_3095;
wire n_3096;
wire n_3097;
wire n_3098;
wire n_3099;
wire n_3100;
wire n_3101;
wire n_3102;
wire n_3103;
wire n_3104;
wire n_3105;
wire n_3106;
wire n_3107;
wire n_3108;
wire n_3109;
wire n_3110;
wire n_3111;
wire n_3112;
wire n_3113;
wire n_3114;
wire n_3115;
wire n_3116;
wire n_3117;
wire n_3118;
wire n_3119;
wire n_3120;
wire n_3121;
wire n_3122;
wire n_3123;
wire n_3124;
wire n_3125;
wire n_3126;
wire n_3127;
wire n_3128;
wire n_3129;
wire n_3130;
wire n_3131;
wire n_3132;
wire n_3133;
wire n_3134;
wire n_3135;
wire n_3136;
wire n_3137;
wire n_3138;
wire n_3139;
wire n_3140;
wire n_3141;
wire n_3142;
wire n_3143;
wire n_3144;
wire n_3145;
wire n_3146;
wire n_3147;
wire n_3148;
wire n_3149;
wire n_3150;
wire n_3151;
wire n_3152;
wire n_3153;
wire n_3154;
wire n_3155;
wire n_3156;
wire n_3157;
wire n_3158;
wire n_3159;
wire n_3160;
wire n_3161;
wire n_3162;
wire n_3163;
wire n_3164;
wire n_3165;
wire n_3166;
wire n_3167;
wire n_3168;
wire n_3169;
wire n_3170;
wire n_3171;
wire n_3172;
wire n_3173;
wire n_3174;
wire n_3175;
wire n_3176;
wire n_3177;
wire n_3178;
wire n_3179;
wire n_3180;
wire n_3181;
wire n_3182;
wire n_3183;
wire n_3184;
wire n_3185;
wire n_3186;
wire n_3187;
wire n_3188;
wire n_3189;
wire n_3190;
wire n_3191;
wire n_3192;
wire n_3193;
wire n_3194;
wire n_3195;
wire n_3196;
wire n_3197;
wire n_3198;
wire n_3199;
wire n_3200;
wire n_3201;
wire n_3202;
wire n_3203;
wire n_3204;
wire n_3205;
wire n_3206;
wire n_3207;
wire n_3208;
wire n_3209;
wire n_3210;
wire n_3211;
wire n_3212;
wire n_3213;
wire n_3214;
wire n_3215;
wire n_3216;
wire n_3217;
wire n_3218;
wire n_3219;
wire n_3220;
wire n_3221;
wire n_3222;
wire n_3223;
wire n_3224;
wire n_3225;
wire n_3226;
wire n_3227;
wire n_3228;
wire n_3229;
wire n_3230;
wire n_3231;
wire n_3232;
wire n_3233;
wire n_3234;
wire n_3235;
wire n_3236;
wire n_3237;
wire n_3238;
wire n_3239;
wire n_3240;
wire n_3241;
wire n_3242;
wire n_3243;
wire n_3244;
wire n_3245;
wire n_3246;
wire n_3247;
wire n_3248;
wire n_3249;
wire n_3250;
wire n_3251;
wire n_3252;
wire n_3253;
wire n_3254;
wire n_3255;
wire n_3256;
wire n_3257;
wire n_3258;
wire n_3259;
wire n_3260;
wire n_3261;
wire n_3262;
wire n_3263;
wire n_3264;
wire n_3265;
wire n_3266;
wire n_3267;
wire n_3268;
wire n_3269;
wire n_3270;
wire n_3271;
wire n_3272;
wire n_3273;
wire n_3274;
wire n_3275;
wire n_3276;
wire n_3277;
wire n_3278;
wire n_3279;
wire n_3280;
wire n_3281;
wire n_3282;
wire n_3283;
wire n_3284;
wire n_3285;
wire n_3286;
wire n_3287;
wire n_3288;
wire n_3289;
wire n_3290;
wire n_3291;
wire n_3292;
wire n_3293;
wire n_3294;
wire n_3295;
wire n_3296;
wire n_3297;
wire n_3298;
wire n_3299;
wire n_3300;
wire n_3301;
wire n_3302;
wire n_3303;
wire n_3304;
wire n_3305;
wire n_3306;
wire n_3307;
wire n_3308;
wire n_3309;
wire n_3310;
wire n_3311;
wire n_3312;
wire n_3313;
wire n_3314;
wire n_3315;
wire n_3316;
wire n_3317;
wire n_3318;
wire n_3319;
wire n_3320;
wire n_3321;
wire n_3322;
wire n_3323;
wire n_3324;
wire n_3325;
wire n_3326;
wire n_3327;
wire n_3328;
wire n_3329;
wire n_3330;
wire n_3331;
wire n_3332;
wire n_3333;
wire n_3334;
wire n_3335;
wire n_3336;
wire n_3337;
wire n_3338;
wire n_3339;
wire n_3340;
wire n_3341;
wire n_3342;
wire n_3343;
wire n_3344;
wire n_3345;
wire n_3346;
wire n_3347;
wire n_3348;
wire n_3349;
wire n_3350;
wire n_3351;
wire n_3352;
wire n_3353;
wire n_3354;
wire n_3355;
wire n_3356;
wire n_3357;
wire n_3358;
wire n_3359;
wire n_3360;
wire n_3361;
wire n_3362;
wire n_3363;
wire n_3364;
wire n_3365;
wire n_3366;
wire n_3367;
wire n_3368;
wire n_3369;
wire n_3370;
wire n_3371;
wire n_3372;
wire n_3373;
wire n_3374;
wire n_3375;
wire n_3376;
wire n_3377;
wire n_3378;
wire n_3379;
wire n_3380;
wire n_3381;
wire n_3382;
wire n_3383;
wire n_3384;
wire n_3385;
wire n_3386;
wire n_3387;
wire n_3388;
wire n_3389;
wire n_3390;
wire n_3391;
wire n_3392;
wire n_3393;
wire n_3394;
wire n_3395;
wire n_3396;
wire n_3397;
wire n_3398;
wire n_3399;
wire n_3400;
wire n_3401;
wire n_3402;
wire n_3403;
wire n_3404;
wire n_3405;
wire n_3406;
wire n_3407;
wire n_3408;
wire n_3409;
wire n_3410;
wire n_3411;
wire n_3412;
wire n_3413;
wire n_3414;
wire n_3415;
wire n_3416;
wire n_3417;
wire n_3418;
wire n_3419;
wire n_3420;
wire n_3421;
wire n_3422;
wire n_3423;
wire n_3424;
wire n_3425;
wire n_3426;
wire n_3427;
wire n_3428;
wire n_3429;
wire n_3430;
wire n_3431;
wire n_3432;
wire n_3433;
wire n_3434;
wire n_3435;
wire n_3436;
wire n_3437;
wire n_3438;
wire n_3439;
wire n_3440;
wire n_3441;
wire n_3442;
wire n_3443;
wire n_3444;
wire n_3445;
wire n_3446;
wire n_3447;
wire n_3448;
wire n_3449;
wire n_3450;
wire n_3451;
wire n_3452;
wire n_3453;
wire n_3454;
wire n_3455;
wire n_3456;
wire n_3457;
wire n_3458;
wire n_3459;
wire n_3460;
wire n_3461;
wire n_3462;
wire n_3463;
wire n_3464;
wire n_3465;
wire n_3466;
wire n_3467;
wire n_3468;
wire n_3469;
wire n_3470;
wire n_3471;
wire n_3472;
wire n_3473;
wire n_3474;
wire n_3475;
wire n_3476;
wire n_3477;
wire n_3478;
wire n_3479;
wire n_3480;
wire n_3481;
wire n_3482;
wire n_3483;
wire n_3484;
wire n_3485;
wire n_3486;
wire n_3487;
wire n_3488;
wire n_3489;
wire n_3490;
wire n_3491;
wire n_3492;
wire n_3493;
wire n_3494;
wire n_3495;
wire n_3496;
wire n_3497;
wire n_3498;
wire n_3499;
wire n_3500;
wire n_3501;
wire n_3502;
wire n_3503;
wire n_3504;
wire n_3505;
wire n_3506;
wire n_3507;
wire n_3508;
wire n_3509;
wire n_3510;
wire n_3511;
wire n_3512;
wire n_3513;
wire n_3514;
wire n_3515;
wire n_3516;
wire n_3517;
wire n_3518;
wire n_3519;
wire n_3520;
wire n_3521;
wire n_3522;
wire n_3523;
wire n_3524;
wire n_3525;
wire n_3526;
wire n_3527;
wire n_3528;
wire n_3529;
wire n_3530;
wire n_3531;
wire n_3532;
wire n_3533;
wire n_3534;
wire n_3535;
wire n_3536;
wire n_3537;
wire n_3538;
wire n_3539;
wire n_3540;
wire n_3541;
wire n_3542;
wire n_3543;
wire n_3544;
wire n_3545;
wire n_3546;
wire n_3547;
wire n_3548;
wire n_3549;
wire n_3550;
wire n_3551;
wire n_3552;
wire n_3553;
wire n_3554;
wire n_3555;
wire n_3556;
wire n_3557;
wire n_3558;
wire n_3559;
wire n_3560;
wire n_3561;
wire n_3562;
wire n_3563;
wire n_3564;
wire n_3565;
wire n_3566;
wire n_3567;
wire n_3568;
wire n_3569;
wire n_3570;
wire n_3571;
wire n_3572;
wire n_3573;
wire n_3574;
wire n_3575;
wire n_3576;
wire n_3577;
wire n_3578;
wire n_3579;
wire n_3580;
wire n_3581;
wire n_3582;
wire n_3583;
wire n_3584;
wire n_3585;
wire n_3586;
wire n_3587;
wire n_3588;
wire n_3589;
wire n_3590;
wire n_3591;
wire n_3592;
wire n_3593;
wire n_3594;
wire n_3595;
wire n_3596;
wire n_3597;
wire n_3598;
wire n_3599;
wire n_3600;
wire n_3601;
wire n_3602;
wire n_3603;
wire n_3604;
wire n_3605;
wire n_3606;
wire n_3607;
wire n_3608;
wire n_3609;
wire n_3610;
wire n_3611;
wire n_3612;
wire n_3613;
wire n_3614;
wire n_3615;
wire n_3616;
wire n_3617;
wire n_3618;
wire n_3619;
wire n_3620;
wire n_3621;
wire n_3622;
wire n_3623;
wire n_3624;
wire n_3625;
wire n_3626;
wire n_3627;
wire n_3628;
wire n_3629;
wire n_3630;
wire n_3631;
wire n_3632;
wire n_3633;
wire n_3634;
wire n_3635;
wire n_3636;
wire n_3637;
wire n_3638;
wire n_3639;
wire n_3640;
wire n_3641;
wire n_3642;
wire n_3643;
wire n_3644;
wire n_3645;
wire n_3646;
wire n_3647;
wire n_3648;
wire n_3649;
wire n_3650;
wire n_3651;
wire n_3652;
wire n_3653;
wire n_3654;
wire n_3655;
wire n_3656;
wire n_3657;
wire n_3658;
wire n_3659;
wire n_3660;
wire n_3661;
wire n_3662;
wire n_3663;
wire n_3664;
wire n_3665;
wire n_3666;
wire n_3667;
wire n_3668;
wire n_3669;
wire n_3670;
wire n_3671;
wire n_3672;
wire n_3673;
wire n_3674;
wire n_3675;
wire n_3676;
wire n_3677;
wire n_3678;
wire n_3679;
wire n_3680;
wire n_3681;
wire n_3682;
wire n_3683;
wire n_3684;
wire n_3685;
wire n_3686;
wire n_3687;
wire n_3688;
wire n_3689;
wire n_3690;
wire n_3691;
wire n_3692;
wire n_3693;
wire n_3694;
wire n_3695;
wire n_3696;
wire n_3697;
wire n_3698;
wire n_3699;
wire n_3700;
wire n_3701;
wire n_3702;
wire n_3703;
wire n_3704;
wire n_3705;
wire n_3706;
wire n_3707;
wire n_3708;
wire n_3709;
wire n_3710;
wire n_3711;
wire n_3712;
wire n_3713;
wire n_3714;
wire n_3715;
wire n_3716;
wire n_3717;
wire n_3718;
wire n_3719;
wire n_3720;
wire n_3721;
wire n_3722;
wire n_3723;
wire n_3724;
wire n_3725;
wire n_3726;
wire n_3727;
wire n_3728;
wire n_3729;
wire n_3730;
wire n_3731;
wire n_3732;
wire n_3733;
wire n_3734;
wire n_3735;
wire n_3736;
wire n_3737;
wire n_3738;
wire n_3739;
wire n_3740;
wire n_3741;
wire n_3742;
wire n_3743;
wire n_3744;
wire n_3745;
wire n_3746;
wire n_3747;
wire n_3748;
wire n_3749;
wire n_3750;
wire n_3751;
wire n_3752;
wire n_3753;
wire n_3754;
wire n_3755;
wire n_3756;
wire n_3757;
wire n_3758;
wire n_3759;
wire n_3760;
wire n_3761;
wire n_3762;
wire n_3763;
wire n_3764;
wire n_3765;
wire n_3766;
wire n_3767;
wire n_3768;
wire n_3769;
wire n_3770;
wire n_3771;
wire n_3772;
wire n_3773;
wire n_3774;
wire n_3775;
wire n_3776;
wire n_3777;
wire n_3778;
wire n_3779;
wire n_3780;
wire n_3781;
wire n_3782;
wire n_3783;
wire n_3784;
wire n_3785;
wire n_3786;
wire n_3787;
wire n_3788;
wire n_3789;
wire n_3790;
wire n_3791;
wire n_3792;
wire n_3793;
wire n_3794;
wire n_3795;
wire n_3796;
wire n_3797;
wire n_3798;
wire n_3799;
wire n_3800;
wire n_3801;
wire n_3802;
wire n_3803;
wire n_3804;
wire n_3805;
wire n_3806;
wire n_3807;
wire n_3808;
wire n_3809;
wire n_3810;
wire n_3811;
wire n_3812;
wire n_3813;
wire n_3814;
wire n_3815;
wire n_3816;
wire n_3817;
wire n_3818;
wire n_3819;
wire n_3820;
wire n_3821;
wire n_3822;
wire n_3823;
wire n_3824;
wire n_3825;
wire n_3826;
wire n_3827;
wire n_3828;
wire n_3829;
wire n_3830;
wire n_3831;
wire n_3832;
wire n_3833;
wire n_3834;
wire n_3835;
wire n_3836;
wire n_3837;
wire n_3838;
wire n_3839;
wire n_3840;
wire n_3841;
wire n_3842;
wire n_3843;
wire n_3844;
wire n_3845;
wire n_3846;
wire n_3847;
wire n_3848;
wire n_3849;
wire n_3850;
wire n_3851;
wire n_3852;
wire n_3853;
wire n_3854;
wire n_3855;
wire n_3856;
wire n_3857;
wire n_3858;
wire n_3859;
wire n_3860;
wire n_3861;
wire n_3862;
wire n_3863;
wire n_3864;
wire n_3865;
wire n_3866;
wire n_3867;
wire n_3868;
wire n_3869;
wire n_3870;
wire n_3871;
wire n_3872;
wire n_3873;
wire n_3874;
wire n_3875;
wire n_3876;
wire n_3877;
wire n_3878;
wire n_3879;
wire n_3880;
wire n_3881;
wire n_3882;
wire n_3883;
wire n_3884;
wire n_3885;
wire n_3886;
wire n_3887;
wire n_3888;
wire n_3889;
wire n_3890;
wire n_3891;
wire n_3892;
wire n_3893;
wire n_3894;
wire n_3895;
wire n_3896;
wire n_3897;
wire n_3898;
wire n_3899;
wire n_3900;
wire n_3901;
wire n_3902;
wire n_3903;
wire n_3904;
wire n_3905;
wire n_3906;
wire n_3907;
wire n_3908;
wire n_3909;
wire n_3910;
wire n_3911;
wire n_3912;
wire n_3913;
wire n_3914;
wire n_3915;
wire n_3916;
wire n_3917;
wire n_3918;
wire n_3919;
wire n_3920;
wire n_3921;
wire n_3922;
wire n_3923;
wire n_3924;
wire n_3925;
wire n_3926;
wire n_3927;
wire n_3928;
wire n_3929;
wire n_3930;
wire n_3931;
wire n_3932;
wire n_3933;
wire n_3934;
wire n_3935;
wire n_3936;
wire n_3937;
wire n_3938;
wire n_3939;
wire n_3940;
wire n_3941;
wire n_3942;
wire n_3943;
wire n_3944;
wire n_3945;
wire n_3946;
wire n_3947;
wire n_3948;
wire n_3949;
wire n_3950;
wire n_3951;
wire n_3952;
wire n_3953;
wire n_3954;
wire n_3955;
wire n_3956;
wire n_3957;
wire n_3958;
wire n_3959;
wire n_3960;
wire n_3961;
wire n_3962;
wire n_3963;
wire n_3964;
wire n_3965;
wire n_3966;
wire n_3967;
wire n_3968;
wire n_3969;
wire n_3970;
wire n_3971;
wire n_3972;
wire n_3973;
wire n_3974;
wire n_3975;
wire n_3976;
wire n_3977;
wire n_3978;
wire n_3979;
wire n_3980;
wire n_3981;
wire n_3982;
wire n_3983;
wire n_3984;
wire n_3985;
wire n_3986;
wire n_3987;
wire n_3988;
wire n_3989;
wire n_3990;
wire n_3991;
wire n_3992;
wire n_3993;
wire n_3994;
wire n_3995;
wire n_3996;
wire n_3997;
wire n_3998;
wire n_3999;
wire n_4000;
wire n_4001;
wire n_4002;
wire n_4003;
wire n_4004;
wire n_4005;
wire n_4006;
wire n_4007;
wire n_4008;
wire n_4009;
wire n_4010;
wire n_4011;
wire n_4012;
wire n_4013;
wire n_4014;
wire n_4015;
wire n_4016;
wire n_4017;
wire n_4018;
wire n_4019;
wire n_4020;
wire n_4021;
wire n_4022;
wire n_4023;
wire n_4024;
wire n_4025;
wire n_4026;
wire n_4027;
wire n_4028;
wire n_4029;
wire n_4030;
wire n_4031;
wire n_4032;
wire n_4033;
wire n_4034;
wire n_4035;
wire n_4036;
wire n_4037;
wire n_4038;
wire n_4039;
wire n_4040;
wire n_4041;
wire n_4042;
wire n_4043;
wire n_4044;
wire n_4045;
wire n_4046;
wire n_4047;
wire n_4048;
wire n_4049;
wire n_4050;
wire n_4051;
wire n_4052;
wire n_4053;
wire n_4054;
wire n_4055;
wire n_4056;
wire n_4057;
wire n_4058;
wire n_4059;
wire n_4060;
wire n_4061;
wire n_4062;
wire n_4063;
wire n_4064;
wire n_4065;
wire n_4066;
wire n_4067;
wire n_4068;
wire n_4069;
wire n_4070;
wire n_4071;
wire n_4072;
wire n_4073;
wire n_4074;
wire n_4075;
wire n_4076;
wire n_4077;
wire n_4078;
wire n_4079;
wire n_4080;
wire n_4081;
wire n_4082;
wire n_4083;
wire n_4084;
wire n_4085;
wire n_4086;
wire n_4087;
wire n_4088;
wire n_4089;
wire n_4090;
wire n_4091;
wire n_4092;
wire n_4093;
wire n_4094;
wire n_4095;
wire n_4096;
wire n_4097;
wire n_4098;
wire n_4099;
wire n_4100;
wire n_4101;
wire n_4102;
wire n_4103;
wire n_4104;
wire n_4105;
wire n_4106;
wire n_4107;
wire n_4108;
wire n_4109;
wire n_4110;
wire n_4111;
wire n_4112;
wire n_4113;
wire n_4114;
wire n_4115;
wire n_4116;
wire n_4117;
wire n_4118;
wire n_4119;
wire n_4120;
wire n_4121;
wire n_4122;
wire n_4123;
wire n_4124;
wire n_4125;
wire n_4126;
wire n_4127;
wire n_4128;
wire n_4129;
wire n_4130;
wire n_4131;
wire n_4132;
wire n_4133;
wire n_4134;
wire n_4135;
wire n_4136;
wire n_4137;
wire n_4138;
wire n_4139;
wire n_4140;
wire n_4141;
wire n_4142;
wire n_4143;
wire n_4144;
wire n_4145;
wire n_4146;
wire n_4147;
wire n_4148;
wire n_4149;
wire n_4150;
wire n_4151;
wire n_4152;
wire n_4153;
wire n_4154;
wire n_4155;
wire n_4156;
wire n_4157;
wire n_4158;
wire n_4159;
wire n_4160;
wire n_4161;
wire n_4162;
wire n_4163;
wire n_4164;
wire n_4165;
wire n_4166;
wire n_4167;
wire n_4168;
wire n_4169;
wire n_4170;
wire n_4171;
wire n_4172;
wire n_4173;
wire n_4174;
wire n_4175;
wire n_4176;
wire n_4177;
wire n_4178;
wire n_4179;
wire n_4180;
wire n_4181;
wire n_4182;
wire n_4183;
wire n_4184;
wire n_4185;
wire n_4186;
wire n_4187;
wire n_4188;
wire n_4189;
wire n_4190;
wire n_4191;
wire n_4192;
wire n_4193;
wire n_4194;
wire n_4195;
wire n_4196;
wire n_4197;
wire n_4198;
wire n_4199;
wire n_4200;
wire n_4201;
wire n_4202;
wire n_4203;
wire n_4204;
wire n_4205;
wire n_4206;
wire n_4207;
wire n_4208;
wire n_4209;
wire n_4210;
wire n_4211;
wire n_4212;
wire n_4213;
wire n_4214;
wire n_4215;
wire n_4216;
wire n_4217;
wire n_4218;
wire n_4219;
wire n_4220;
wire n_4221;
wire n_4222;
wire n_4223;
wire n_4224;
wire n_4225;
wire n_4226;
wire n_4227;
wire n_4228;
wire n_4229;
wire n_4230;
wire n_4231;
wire n_4232;
wire n_4233;
wire n_4234;
wire n_4235;
wire n_4236;
wire n_4237;
wire n_4238;
wire n_4239;
wire n_4240;
wire n_4241;
wire n_4242;
wire n_4243;
wire n_4244;
wire n_4245;
wire n_4246;
wire n_4247;
wire n_4248;
wire n_4249;
wire n_4250;
wire n_4251;
wire n_4252;
wire n_4253;
wire n_4254;
wire n_4255;
wire n_4256;
wire n_4257;
wire n_4258;
wire n_4259;
wire n_4260;
wire n_4261;
wire n_4262;
wire n_4263;
wire n_4264;
wire n_4265;
wire n_4266;
wire n_4267;
wire n_4268;
wire n_4269;
wire n_4270;
wire n_4271;
wire n_4272;
wire n_4273;
wire n_4274;
wire n_4275;
wire n_4276;
wire n_4277;
wire n_4278;
wire n_4279;
wire n_4280;
wire n_4281;
wire n_4282;
wire n_4283;
wire n_4284;
wire n_4285;
wire n_4286;
wire n_4287;
wire n_4288;
wire n_4289;
wire n_4290;
wire n_4291;
wire n_4292;
wire n_4293;
wire n_4294;
wire n_4295;
wire n_4296;
wire n_4297;
wire n_4298;
wire n_4299;
wire n_4300;
wire n_4301;
wire n_4302;
wire n_4303;
wire n_4304;
wire n_4305;
wire n_4306;
wire n_4307;
wire n_4308;
wire n_4309;
wire n_4310;
wire n_4311;
wire n_4312;
wire n_4313;
wire n_4314;
wire n_4315;
wire n_4316;
wire n_4317;
wire n_4318;
wire n_4319;
wire n_4320;
wire n_4321;
wire n_4322;
wire n_4323;
wire n_4324;
wire n_4325;
wire n_4326;
wire n_4327;
wire n_4328;
wire n_4329;
wire n_4330;
wire n_4331;
wire n_4332;
wire n_4333;
wire n_4334;
wire n_4335;
wire n_4336;
wire n_4337;
wire n_4338;
wire n_4339;
wire n_4340;
wire n_4341;
wire n_4342;
wire n_4343;
wire n_4344;
wire n_4345;
wire n_4346;
wire n_4347;
wire n_4348;
wire n_4349;
wire n_4350;
wire n_4351;
wire n_4352;
wire n_4353;
wire n_4354;
wire n_4355;
wire n_4356;
wire n_4357;
wire n_4358;
wire n_4359;
wire n_4360;
wire n_4361;
wire n_4362;
wire n_4363;
wire n_4364;
wire n_4365;
wire n_4366;
wire n_4367;
wire n_4368;
wire n_4369;
wire n_4370;
wire n_4371;
wire n_4372;
wire n_4373;
wire n_4374;
wire n_4375;
wire n_4376;
wire n_4377;
wire n_4378;
wire n_4379;
wire n_4380;
wire n_4381;
wire n_4382;
wire n_4383;
wire n_4384;
wire n_4385;
wire n_4386;
wire n_4387;
wire n_4388;
wire n_4389;
wire n_4390;
wire n_4391;
wire n_4392;
wire n_4393;
wire n_4394;
wire n_4395;
wire n_4396;
wire n_4397;
wire n_4398;
wire n_4399;
wire n_4400;
wire n_4401;
wire n_4402;
wire n_4403;
wire n_4404;
wire n_4405;
wire n_4406;
wire n_4407;
wire n_4408;
wire n_4409;
wire n_4410;
wire n_4411;
wire n_4412;
wire n_4413;
wire n_4414;
wire n_4415;
wire n_4416;
wire n_4417;
wire n_4418;
wire n_4419;
wire n_4420;
wire n_4421;
wire n_4422;
wire n_4423;
wire n_4424;
wire n_4425;
wire n_4426;
wire n_4427;
wire n_4428;
wire n_4429;
wire n_4430;
wire n_4431;
wire n_4432;
wire n_4433;
wire n_4434;
wire n_4435;
wire n_4436;
wire n_4437;
wire n_4438;
wire n_4439;
wire n_4440;
wire n_4441;
wire n_4442;
wire n_4443;
wire n_4444;
wire n_4445;
wire n_4446;
wire n_4447;
wire n_4448;
wire n_4449;
wire n_4450;
wire n_4451;
wire n_4452;
wire n_4453;
wire n_4454;
wire n_4455;
wire n_4456;
wire n_4457;
wire n_4458;
wire n_4459;
wire n_4460;
wire n_4461;
wire n_4462;
wire n_4463;
wire n_4464;
wire n_4465;
wire n_4466;
wire n_4467;
wire n_4468;
wire n_4469;
wire n_4470;
wire n_4471;
wire n_4472;
wire n_4473;
wire n_4474;
wire n_4475;
wire n_4476;
wire n_4477;
wire n_4478;
wire n_4479;
wire n_4480;
wire n_4481;
wire n_4482;
wire n_4483;
wire n_4484;
wire n_4485;
wire n_4486;
wire n_4487;
wire n_4488;
wire n_4489;
wire n_4490;
wire n_4491;
wire n_4492;
wire n_4493;
wire n_4494;
wire n_4495;
wire n_4496;
wire n_4497;
wire n_4498;
wire n_4499;
wire n_4500;
wire n_4501;
wire n_4502;
wire n_4503;
wire n_4504;
wire n_4505;
wire n_4506;
wire n_4507;
wire n_4508;
wire n_4509;
wire n_4510;
wire n_4511;
wire n_4512;
wire n_4513;
wire n_4514;
wire n_4515;
wire n_4516;
wire n_4517;
wire n_4518;
wire n_4519;
wire n_4520;
wire n_4521;
wire n_4522;
wire n_4523;
wire n_4524;
wire n_4525;
wire n_4526;
wire n_4527;
wire n_4528;
wire n_4529;
wire n_4530;
wire n_4531;
wire n_4532;
wire n_4533;
wire n_4534;
wire n_4535;
wire n_4536;
wire n_4537;
wire n_4538;
wire n_4539;
wire n_4540;
wire n_4541;
wire n_4542;
wire n_4543;
wire n_4544;
wire n_4545;
wire n_4546;
wire n_4547;
wire n_4548;
wire n_4549;
wire n_4550;
wire n_4551;
wire n_4552;
wire n_4553;
wire n_4554;
wire n_4555;
wire n_4556;
wire n_4557;
wire n_4558;
wire n_4559;
wire n_4560;
wire n_4561;
wire n_4562;
wire n_4563;
wire n_4564;
wire n_4565;
wire n_4566;
wire n_4567;
wire n_4568;
wire n_4569;
wire n_4570;
wire n_4571;
wire n_4572;
wire n_4573;
wire n_4574;
wire n_4575;
wire n_4576;
wire n_4577;
wire n_4578;
wire n_4579;
wire n_4580;
wire n_4581;
wire n_4582;
wire n_4583;
wire n_4584;
wire n_4585;
wire n_4586;
wire n_4587;
wire n_4588;
wire n_4589;
wire n_4590;
wire n_4591;
wire n_4592;
wire n_4593;
wire n_4594;
wire n_4595;
wire n_4596;
wire n_4597;
wire n_4598;
wire n_4599;
wire n_4600;
wire n_4601;
wire n_4602;
wire n_4603;
wire n_4604;
wire n_4605;
wire n_4606;
wire n_4607;
wire n_4608;
wire n_4609;
wire n_4610;
wire n_4611;
wire n_4612;
wire n_4613;
wire n_4614;
wire n_4615;
wire n_4616;
wire n_4617;
wire n_4618;
wire n_4619;
wire n_4620;
wire n_4621;
wire n_4622;
wire n_4623;
wire n_4624;
wire n_4625;
wire n_4626;
wire n_4627;
wire n_4628;
wire n_4629;
wire n_4630;
wire n_4631;
wire n_4632;
wire n_4633;
wire n_4634;
wire n_4635;
wire n_4636;
wire n_4637;
wire n_4638;
wire n_4639;
wire n_4640;
wire n_4641;
wire n_4642;
wire n_4643;
wire n_4644;
wire n_4645;
wire n_4646;
wire n_4647;
wire n_4648;
wire n_4649;
wire n_4650;
wire n_4651;
wire n_4652;
wire n_4653;
wire n_4654;
wire n_4655;
wire n_4656;
wire n_4657;
wire n_4658;
wire n_4659;
wire n_4660;
wire n_4661;
wire n_4662;
wire n_4663;
wire n_4664;
wire n_4665;
wire n_4666;
wire n_4667;
wire n_4668;
wire n_4669;
wire n_4670;
wire n_4671;
wire n_4672;
wire n_4673;
wire n_4674;
wire n_4675;
wire n_4676;
wire n_4677;
wire n_4678;
wire n_4679;
wire n_4680;
wire n_4681;
wire n_4682;
wire n_4683;
wire n_4684;
wire n_4685;
wire n_4686;
wire n_4687;
wire n_4688;
wire n_4689;
wire n_4690;
wire n_4691;
wire n_4692;
wire n_4693;
wire n_4694;
wire n_4695;
wire n_4696;
wire n_4697;
wire n_4698;
wire n_4699;
wire n_4700;
wire n_4701;
wire n_4702;
wire n_4703;
wire n_4704;
wire n_4705;
wire n_4706;
wire n_4707;
wire n_4708;
wire n_4709;
wire n_4710;
wire n_4711;
wire n_4712;
wire n_4713;
wire n_4714;
wire n_4715;
wire n_4716;
wire n_4717;
wire n_4718;
wire n_4719;
wire n_4720;
wire n_4721;
wire n_4722;
wire n_4723;
wire n_4724;
wire n_4725;
wire n_4726;
wire n_4727;
wire n_4728;
wire n_4729;
wire n_4730;
wire n_4731;
wire n_4732;
wire n_4733;
wire n_4734;
wire n_4735;
wire n_4736;
wire n_4737;
wire n_4738;
wire n_4739;
wire n_4740;
wire n_4741;
wire n_4742;
wire n_4743;
wire n_4744;
wire n_4745;
wire n_4746;
wire n_4747;
wire n_4748;
wire n_4749;
wire n_4750;
wire n_4751;
wire n_4752;
wire n_4753;
wire n_4754;
wire n_4755;
wire n_4756;
wire n_4757;
wire n_4758;
wire n_4759;
wire n_4760;
wire n_4761;
wire n_4762;
wire n_4763;
wire n_4764;
wire n_4765;
wire n_4766;
wire n_4767;
wire n_4768;
wire n_4769;
wire n_4770;
wire n_4771;
wire n_4772;
wire n_4773;
wire n_4774;
wire n_4775;
wire n_4776;
wire n_4777;
wire n_4778;
wire n_4779;
wire n_4780;
wire n_4781;
wire n_4782;
wire n_4783;
wire n_4784;
wire n_4785;
wire n_4786;
wire n_4787;
wire n_4788;
wire n_4789;
wire n_4790;
wire n_4791;
wire n_4792;
wire n_4793;
wire n_4794;
wire n_4795;
wire n_4796;
wire n_4797;
wire n_4798;
wire n_4799;
wire n_4800;
wire n_4801;
wire n_4802;
wire n_4803;
wire n_4804;
wire n_4805;
wire n_4806;
wire n_4807;
wire n_4808;
wire n_4809;
wire n_4810;
wire n_4811;
wire n_4812;
wire n_4813;
wire n_4814;
wire n_4815;
wire n_4816;
wire n_4817;
wire n_4818;
wire n_4819;
wire n_4820;
wire n_4821;
wire n_4822;
wire n_4823;
wire n_4824;
wire n_4825;
wire n_4826;
wire n_4827;
wire n_4828;
wire n_4829;
wire n_4830;
wire n_4831;
wire n_4832;
wire n_4833;
wire n_4834;
wire n_4835;
wire n_4836;
wire n_4837;
wire n_4838;
wire n_4839;
wire n_4840;
wire n_4841;
wire n_4842;
wire n_4843;
wire n_4844;
wire n_4845;
wire n_4846;
wire n_4847;
wire n_4848;
wire n_4849;
wire n_4850;
wire n_4851;
wire n_4852;
wire n_4853;
wire n_4854;
wire n_4855;
wire n_4856;
wire n_4857;
wire n_4858;
wire n_4859;
wire n_4860;
wire n_4861;
wire n_4862;
wire n_4863;
wire n_4864;
wire n_4865;
wire n_4866;
wire n_4867;
wire n_4868;
wire n_4869;
wire n_4870;
wire n_4871;
wire n_4872;
wire n_4873;
wire n_4874;
wire n_4875;
wire n_4876;
wire n_4877;
wire n_4878;
wire n_4879;
wire n_4880;
wire n_4881;
wire n_4882;
wire n_4883;
wire n_4884;
wire n_4885;
wire n_4886;
wire n_4887;
wire n_4888;
wire n_4889;
wire n_4890;
wire n_4891;
wire n_4892;
wire n_4893;
wire n_4894;
wire n_4895;
wire n_4896;
wire n_4897;
wire n_4898;
wire n_4899;
wire n_4900;
wire n_4901;
wire n_4902;
wire n_4903;
wire n_4904;
wire n_4905;
wire n_4906;
wire n_4907;
wire n_4908;
wire n_4909;
wire n_4910;
wire n_4911;
wire n_4912;
wire n_4913;
wire n_4914;
wire n_4915;
wire n_4916;
wire n_4917;
wire n_4918;
wire n_4919;
wire n_4920;
wire n_4921;
wire n_4922;
wire n_4923;
wire n_4924;
wire n_4925;
wire n_4926;
wire n_4927;
wire n_4928;
wire n_4929;
wire n_4930;
wire n_4931;
wire n_4932;
wire n_4933;
wire n_4934;
wire n_4935;
wire n_4936;
wire n_4937;
wire n_4938;
wire n_4939;
wire n_4940;
wire n_4941;
wire n_4942;
wire n_4943;
wire n_4944;
wire n_4945;
wire n_4946;
wire n_4947;
wire n_4948;
wire n_4949;
wire n_4950;
wire n_4951;
wire n_4952;
wire n_4953;
wire n_4954;
wire n_4955;
wire n_4956;
wire n_4957;
wire n_4958;
wire n_4959;
wire n_4960;
wire n_4961;
wire n_4962;
wire n_4963;
wire n_4964;
wire n_4965;
wire n_4966;
wire n_4967;
wire n_4968;
wire n_4969;
wire n_4970;
wire n_4971;
wire n_4972;
wire n_4973;
wire n_4974;
wire n_4975;
wire n_4976;
wire n_4977;
wire n_4978;
wire n_4979;
wire n_4980;
wire n_4981;
wire n_4982;
wire n_4983;
wire n_4984;
wire n_4985;
wire n_4986;
wire n_4987;
wire n_4988;
wire n_4989;
wire n_4990;
wire n_4991;
wire n_4992;
wire n_4993;
wire n_4994;
wire n_4995;
wire n_4996;
wire n_4997;
wire n_4998;
wire n_4999;
wire n_5000;
wire n_5001;
wire n_5002;
wire n_5003;
wire n_5004;
wire n_5005;
wire n_5006;
wire n_5007;
wire n_5008;
wire n_5009;
wire n_5010;
wire n_5011;
wire n_5012;
wire n_5013;
wire n_5014;
wire n_5015;
wire n_5016;
wire n_5017;
wire n_5018;
wire n_5019;
wire n_5020;
wire n_5021;
wire n_5022;
wire n_5023;
wire n_5024;
wire n_5025;
wire n_5026;
wire n_5027;
wire n_5028;
wire n_5029;
wire n_5030;
wire n_5031;
wire n_5032;
wire n_5033;
wire n_5034;
wire n_5035;
wire n_5036;
wire n_5037;
wire n_5038;
wire n_5039;
wire n_5040;
wire n_5041;
wire n_5042;
wire n_5043;
wire n_5044;
wire n_5045;
wire n_5046;
wire n_5047;
wire n_5048;
wire n_5049;
wire n_5050;
wire n_5051;
wire n_5052;
wire n_5053;
wire n_5054;
wire n_5055;
wire n_5056;
wire n_5057;
wire n_5058;
wire n_5059;
wire n_5060;
wire n_5061;
wire n_5062;
wire n_5063;
wire n_5064;
wire n_5065;
wire n_5066;
wire n_5067;
wire n_5068;
wire n_5069;
wire n_5070;
wire n_5071;
wire n_5072;
wire n_5073;
wire n_5074;
wire n_5075;
wire n_5076;
wire n_5077;
wire n_5078;
wire n_5079;
wire n_5080;
wire n_5081;
wire n_5082;
wire n_5083;
wire n_5084;
wire n_5085;
wire n_5086;
wire n_5087;
wire n_5088;
wire n_5089;
wire n_5090;
wire n_5091;
wire n_5092;
wire n_5093;
wire n_5094;
wire n_5095;
wire n_5096;
wire n_5097;
wire n_5098;
wire n_5099;
wire n_5100;
wire n_5101;
wire n_5102;
wire n_5103;
wire n_5104;
wire n_5105;
wire n_5106;
wire n_5107;
wire n_5108;
wire n_5109;
wire n_5110;
wire n_5111;
wire n_5112;
wire n_5113;
wire n_5114;
wire n_5115;
wire n_5116;
wire n_5117;
wire n_5118;
wire n_5119;
wire n_5120;
wire n_5121;
wire n_5122;
wire n_5123;
wire n_5124;
wire n_5125;
wire n_5126;
wire n_5127;
wire n_5128;
wire n_5129;
wire n_5130;
wire n_5131;
wire n_5132;
wire n_5133;
wire n_5134;
wire n_5135;
wire n_5136;
wire n_5137;
wire n_5138;
wire n_5139;
wire n_5140;
wire n_5141;
wire n_5142;
wire n_5143;
wire n_5144;
wire n_5145;
wire n_5146;
wire n_5147;
wire n_5148;
wire n_5149;
wire n_5150;
wire n_5151;
wire n_5152;
wire n_5153;
wire n_5154;
wire n_5155;
wire n_5156;
wire n_5157;
wire n_5158;
wire n_5159;
wire n_5160;
wire n_5161;
wire n_5162;
wire n_5163;
wire n_5164;
wire n_5165;
wire n_5166;
wire n_5167;
wire n_5168;
wire n_5169;
wire n_5170;
wire n_5171;
wire n_5172;
wire n_5173;
wire n_5174;
wire n_5175;
wire n_5176;
wire n_5177;
wire n_5178;
wire n_5179;
wire n_5180;
wire n_5181;
wire n_5182;
wire n_5183;
wire n_5184;
wire n_5185;
wire n_5186;
wire n_5187;
wire n_5188;
wire n_5189;
wire n_5190;
wire n_5191;
wire n_5192;
wire n_5193;
wire n_5194;
wire n_5195;
wire n_5196;
wire n_5197;
wire n_5198;
wire n_5199;
wire n_5200;
wire n_5201;
wire n_5202;
wire n_5203;
wire n_5204;
wire n_5205;
wire n_5206;
wire n_5207;
wire n_5208;
wire n_5209;
wire n_5210;
wire n_5211;
wire n_5212;
wire n_5213;
wire n_5214;
wire n_5215;
wire n_5216;
wire n_5217;
wire n_5218;
wire n_5219;
wire n_5220;
wire n_5221;
wire n_5222;
wire n_5223;
wire n_5224;
wire n_5225;
wire n_5226;
wire n_5227;
wire n_5228;
wire n_5229;
wire n_5230;
wire n_5231;
wire n_5232;
wire n_5233;
wire n_5234;
wire n_5235;
wire n_5236;
wire n_5237;
wire n_5238;
wire n_5239;
wire n_5240;
wire n_5241;
wire n_5242;
wire n_5243;
wire n_5244;
wire n_5245;
wire n_5246;
wire n_5247;
wire n_5248;
wire n_5249;
wire n_5250;
wire n_5251;
wire n_5252;
wire n_5253;
wire n_5254;
wire n_5255;
wire n_5256;
wire n_5257;
wire n_5258;
wire n_5259;
wire n_5260;
wire n_5261;
wire n_5262;
wire n_5263;
wire n_5264;
wire n_5265;
wire n_5266;
wire n_5267;
wire n_5268;
wire n_5269;
wire n_5270;
wire n_5271;
wire n_5272;
wire n_5273;
wire n_5274;
wire n_5275;
wire n_5276;
wire n_5277;
wire n_5278;
wire n_5279;
wire n_5280;
wire n_5281;
wire n_5282;
wire n_5283;
wire n_5284;
wire n_5285;
wire n_5286;
wire n_5287;
wire n_5288;
wire n_5289;
wire n_5290;
wire n_5291;
wire n_5292;
wire n_5293;
wire n_5294;
wire n_5295;
wire n_5296;
wire n_5297;
wire n_5298;
wire n_5299;
wire n_5300;
wire n_5301;
wire n_5302;
wire n_5303;
wire n_5304;
wire n_5305;
wire n_5306;
wire n_5307;
wire n_5308;
wire n_5309;
wire n_5310;
wire n_5311;
wire n_5312;
wire n_5313;
wire n_5314;
wire n_5315;
wire n_5316;
wire n_5317;
wire n_5318;
wire n_5319;
wire n_5320;
wire n_5321;
wire n_5322;
wire n_5323;
wire n_5324;
wire n_5325;
wire n_5326;
wire n_5327;
wire n_5328;
wire n_5329;
wire n_5330;
wire n_5331;
wire n_5332;
wire n_5333;
wire n_5334;
wire n_5335;
wire n_5336;
wire n_5337;
wire n_5338;
wire n_5339;
wire n_5340;
wire n_5341;
wire n_5342;
wire n_5343;
wire n_5344;
wire n_5345;
wire n_5346;
wire n_5347;
wire n_5348;
wire n_5349;
wire n_5350;
wire n_5351;
wire n_5352;
wire n_5353;
wire n_5354;
wire n_5355;
wire n_5356;
wire n_5357;
wire n_5358;
wire n_5359;
wire n_5360;
wire n_5361;
wire n_5362;
wire n_5363;
wire n_5364;
wire n_5365;
wire n_5366;
wire n_5367;
wire n_5368;
wire n_5369;
wire n_5370;
wire n_5371;
wire n_5372;
wire n_5373;
wire n_5374;
wire n_5375;
wire n_5376;
wire n_5377;
wire n_5378;
wire n_5379;
wire n_5380;
wire n_5381;
wire n_5382;
wire n_5383;
wire n_5384;
wire n_5385;
wire n_5386;
wire n_5387;
wire n_5388;
wire n_5389;
wire n_5390;
wire n_5391;
wire n_5392;
wire n_5393;
wire n_5394;
wire n_5395;
wire n_5396;
wire n_5397;
wire n_5398;
wire n_5399;
wire n_5400;
wire n_5401;
wire n_5402;
wire n_5403;
wire n_5404;
wire n_5405;
wire n_5406;
wire n_5407;
wire n_5408;
wire n_5409;
wire n_5410;
wire n_5411;
wire n_5412;
wire n_5413;
wire n_5414;
wire n_5415;
wire n_5416;
wire n_5417;
wire n_5418;
wire n_5419;
wire n_5420;
wire n_5421;
wire n_5422;
wire n_5423;
wire n_5424;
wire n_5425;
wire n_5426;
wire n_5427;
wire n_5428;
wire n_5429;
wire n_5430;
wire n_5431;
wire n_5432;
wire n_5433;
wire n_5434;
wire n_5435;
wire n_5436;
wire n_5437;
wire n_5438;
wire n_5439;
wire n_5440;
wire n_5441;
wire n_5442;
wire n_5443;
wire n_5444;
wire n_5445;
wire n_5446;
wire n_5447;
wire n_5448;
wire n_5449;
wire n_5450;
wire n_5451;
wire n_5452;
wire n_5453;
wire n_5454;
wire n_5455;
wire n_5456;
wire n_5457;
wire n_5458;
wire n_5459;
wire n_5460;
wire n_5461;
wire n_5462;
wire n_5463;
wire n_5464;
wire n_5465;
wire n_5466;
wire n_5467;
wire n_5468;
wire n_5469;
wire n_5470;
wire n_5471;
wire n_5472;
wire n_5473;
wire n_5474;
wire n_5475;
wire n_5476;
wire n_5477;
wire n_5478;
wire n_5479;
wire n_5480;
wire n_5481;
wire n_5482;
wire n_5483;
wire n_5484;
wire n_5485;
wire n_5486;
wire n_5487;
wire n_5488;
wire n_5489;
wire n_5490;
wire n_5491;
wire n_5492;
wire n_5493;
wire n_5494;
wire n_5495;
wire n_5496;
wire n_5497;
wire n_5498;
wire n_5499;
wire n_5500;
wire n_5501;
wire n_5502;
wire n_5503;
wire n_5504;
wire n_5505;
wire n_5506;
wire n_5507;
wire n_5508;
wire n_5509;
wire n_5510;
wire n_5511;
wire n_5512;
wire n_5513;
wire n_5514;
wire n_5515;
wire n_5516;
wire n_5517;
wire n_5518;
wire n_5519;
wire n_5520;
wire n_5521;
wire n_5522;
wire n_5523;
wire n_5524;
wire n_5525;
wire n_5526;
wire n_5527;
wire n_5528;
wire n_5529;
wire n_5530;
wire n_5531;
wire n_5532;
wire n_5533;
wire n_5534;
wire n_5535;
wire n_5536;
wire n_5537;
wire n_5538;
wire n_5539;
wire n_5540;
wire n_5541;
wire n_5542;
wire n_5543;
wire n_5544;
wire n_5545;
wire n_5546;
wire n_5547;
wire n_5548;
wire n_5549;
wire n_5550;
wire n_5551;
wire n_5552;
wire n_5553;
wire n_5554;
wire n_5555;
wire n_5556;
wire n_5557;
wire n_5558;
wire n_5559;
wire n_5560;
wire n_5561;
wire n_5562;
wire n_5563;
wire n_5564;
wire n_5565;
wire n_5566;
wire n_5567;
wire n_5568;
wire n_5569;
wire n_5570;
wire n_5571;
wire n_5572;
wire n_5573;
wire n_5574;
wire n_5575;
wire n_5576;
wire n_5577;
wire n_5578;
wire n_5579;
wire n_5580;
wire n_5581;
wire n_5582;
wire n_5583;
wire n_5584;
wire n_5585;
wire n_5586;
wire n_5587;
wire n_5588;
wire n_5589;
wire n_5590;
wire n_5591;
wire n_5592;
wire n_5593;
wire n_5594;
wire n_5595;
wire n_5596;
wire n_5597;
wire n_5598;
wire n_5599;
wire n_5600;
wire n_5601;
wire n_5602;
wire n_5603;
wire n_5604;
wire n_5605;
wire n_5606;
wire n_5607;
wire n_5608;
wire n_5609;
wire n_5610;
wire n_5611;
wire n_5612;
wire n_5613;
wire n_5614;
wire n_5615;
wire n_5616;
wire n_5617;
wire n_5618;
wire n_5619;
wire n_5620;
wire n_5621;
wire n_5622;
wire n_5623;
wire n_5624;
wire n_5625;
wire n_5626;
wire n_5627;
wire n_5628;
wire n_5629;
wire n_5630;
wire n_5631;
wire n_5632;
wire n_5633;
wire n_5634;
wire n_5635;
wire n_5636;
wire n_5637;
wire n_5638;
wire n_5639;
wire n_5640;
wire n_5641;
wire n_5642;
wire n_5643;
wire n_5644;
wire n_5645;
wire n_5646;
wire n_5647;
wire n_5648;
wire n_5649;
wire n_5650;
wire n_5651;
wire n_5652;
wire n_5653;
wire n_5654;
wire n_5655;
wire n_5656;
wire n_5657;
wire n_5658;
wire n_5659;
wire n_5660;
wire n_5661;
wire n_5662;
wire n_5663;
wire n_5664;
wire n_5665;
wire n_5666;
wire n_5667;
wire n_5668;
wire n_5669;
wire n_5670;
wire n_5671;
wire n_5672;
wire n_5673;
wire n_5674;
wire n_5675;
wire n_5676;
wire n_5677;
wire n_5678;
wire n_5679;
wire n_5680;
wire n_5681;
wire n_5682;
wire n_5683;
wire n_5684;
wire n_5685;
wire n_5686;
wire n_5687;
wire n_5688;
wire n_5689;
wire n_5690;
wire n_5691;
wire n_5692;
wire n_5693;
wire n_5694;
wire n_5695;
wire n_5696;
wire n_5697;
wire n_5698;
wire n_5699;
wire n_5700;
wire n_5701;
wire n_5702;
wire n_5703;
wire n_5704;
wire n_5705;
wire n_5706;
wire n_5707;
wire n_5708;
wire n_5709;
wire n_5710;
wire n_5711;
wire n_5712;
wire n_5713;
wire n_5714;
wire n_5715;
wire n_5716;
wire n_5717;
wire n_5718;
wire n_5719;
wire n_5720;
wire n_5721;
wire n_5722;
wire n_5723;
wire n_5724;
wire n_5725;
wire n_5726;
wire n_5727;
wire n_5728;
wire n_5729;
wire n_5730;
wire n_5731;
wire n_5732;
wire n_5733;
wire n_5734;
wire n_5735;
wire n_5736;
wire n_5737;
wire n_5738;
wire n_5739;
wire n_5740;
wire n_5741;
wire n_5742;
wire n_5743;
wire n_5744;
wire n_5745;
wire n_5746;
wire n_5747;
wire n_5748;
wire n_5749;
wire n_5750;
wire n_5751;
wire n_5752;
wire n_5753;
wire n_5754;
wire n_5755;
wire n_5756;
wire n_5757;
wire n_5758;
wire n_5759;
wire n_5760;
wire n_5761;
wire n_5762;
wire n_5763;
wire n_5764;
wire n_5765;
wire n_5766;
wire n_5767;
wire n_5768;
wire n_5769;
wire n_5770;
wire n_5771;
wire n_5772;
wire n_5773;
wire n_5774;
wire n_5775;
wire n_5776;
wire n_5777;
wire n_5778;
wire n_5779;
wire n_5780;
wire n_5781;
wire n_5782;
wire n_5783;
wire n_5784;
wire n_5785;
wire n_5786;
wire n_5787;
wire n_5788;
wire n_5789;
wire n_5790;
wire n_5791;
wire n_5792;
wire n_5793;
wire n_5794;
wire n_5795;
wire n_5796;
wire n_5797;
wire n_5798;
wire n_5799;
wire n_5800;
wire n_5801;
wire n_5802;
wire n_5803;
wire n_5804;
wire n_5805;
wire n_5806;
wire n_5807;
wire n_5808;
wire n_5809;
wire n_5810;
wire n_5811;
wire n_5812;
wire n_5813;
wire n_5814;
wire n_5815;
wire n_5816;
wire n_5817;
wire n_5818;
wire n_5819;
wire n_5820;
wire n_5821;
wire n_5822;
wire n_5823;
wire n_5824;
wire n_5825;
wire n_5826;
wire n_5827;
wire n_5828;
wire n_5829;
wire n_5830;
wire n_5831;
wire n_5832;
wire n_5833;
wire n_5834;
wire n_5835;
wire n_5836;
wire n_5837;
wire n_5838;
wire n_5839;
wire n_5840;
wire n_5841;
wire n_5842;
wire n_5843;
wire n_5844;
wire n_5845;
wire n_5846;
wire n_5847;
wire n_5848;
wire n_5849;
wire n_5850;
wire n_5851;
wire n_5852;
wire n_5853;
wire n_5854;
wire n_5855;
wire n_5856;
wire n_5857;
wire n_5858;
wire n_5859;
wire n_5860;
wire n_5861;
wire n_5862;
wire n_5863;
wire n_5864;
wire n_5865;
wire n_5866;
wire n_5867;
wire n_5868;
wire n_5869;
wire n_5870;
wire n_5871;
wire n_5872;
wire n_5873;
wire n_5874;
wire n_5875;
wire n_5876;
wire n_5877;
wire n_5878;
wire n_5879;
wire n_5880;
wire n_5881;
wire n_5882;
wire n_5883;
wire n_5884;
wire n_5885;
wire n_5886;
wire n_5887;
wire n_5888;
wire n_5889;
wire n_5890;
wire n_5891;
wire n_5892;
wire n_5893;
wire n_5894;
wire n_5895;
wire n_5896;
wire n_5897;
wire n_5898;
wire n_5899;
wire n_5900;
wire n_5901;
wire n_5902;
wire n_5903;
wire n_5904;
wire n_5905;
wire n_5906;
wire n_5907;
wire n_5908;
wire n_5909;
wire n_5910;
wire n_5911;
wire n_5912;
wire n_5913;
wire n_5914;
wire n_5915;
wire n_5916;
wire n_5917;
wire n_5918;
wire n_5919;
wire n_5920;
wire n_5921;
wire n_5922;
wire n_5923;
wire n_5924;
wire n_5925;
wire n_5926;
wire n_5927;
wire n_5928;
wire n_5929;
wire n_5930;
wire n_5931;
wire n_5932;
wire n_5933;
wire n_5934;
wire n_5935;
wire n_5936;
wire n_5937;
wire n_5938;
wire n_5939;
wire n_5940;
wire n_5941;
wire n_5942;
wire n_5943;
wire n_5944;
wire n_5945;
wire n_5946;
wire n_5947;
wire n_5948;
wire n_5949;
wire n_5950;
wire n_5951;
wire n_5952;
wire n_5953;
wire n_5954;
wire n_5955;
wire n_5956;
wire n_5957;
wire n_5958;
wire n_5959;
wire n_5960;
wire n_5961;
wire n_5962;
wire n_5963;
wire n_5964;
wire n_5965;
wire n_5966;
wire n_5967;
wire n_5968;
wire n_5969;
wire n_5970;
wire n_5971;
wire n_5972;
wire n_5973;
wire n_5974;
wire n_5975;
wire n_5976;
wire n_5977;
wire n_5978;
wire n_5979;
wire n_5980;
wire n_5981;
wire n_5982;
wire n_5983;
wire n_5984;
wire n_5985;
wire n_5986;
wire n_5987;
wire n_5988;
wire n_5989;
wire n_5990;
wire n_5991;
wire n_5992;
wire n_5993;
wire n_5994;
wire n_5995;
wire n_5996;
wire n_5997;
wire n_5998;
wire n_5999;
wire n_6000;
wire n_6001;
wire n_6002;
wire n_6003;
wire n_6004;
wire n_6005;
wire n_6006;
wire n_6007;
wire n_6008;
wire n_6009;
wire n_6010;
wire n_6011;
wire n_6012;
wire n_6013;
wire n_6014;
wire n_6015;
wire n_6016;
wire n_6017;
wire n_6018;
wire n_6019;
wire n_6020;
wire n_6021;
wire n_6022;
wire n_6023;
wire n_6024;
wire n_6025;
wire n_6026;
wire n_6027;
wire n_6028;
wire n_6029;
wire n_6030;
wire n_6031;
wire n_6032;
wire n_6033;
wire n_6034;
wire n_6035;
wire n_6036;
wire n_6037;
wire n_6038;
wire n_6039;
wire n_6040;
wire n_6041;
wire n_6042;
wire n_6043;
wire n_6044;
wire n_6045;
wire n_6046;
wire n_6047;
wire n_6048;
wire n_6049;
wire n_6050;
wire n_6051;
wire n_6052;
wire n_6053;
wire n_6054;
wire n_6055;
wire n_6056;
wire n_6057;
wire n_6058;
wire n_6059;
wire n_6060;
wire n_6061;
wire n_6062;
wire n_6063;
wire n_6064;
wire n_6065;
wire n_6066;
wire n_6067;
wire n_6068;
wire n_6069;
wire n_6070;
wire n_6071;
wire n_6072;
wire n_6073;
wire n_6074;
wire n_6075;
wire n_6076;
wire n_6077;
wire n_6078;
wire n_6079;
wire n_6080;
wire n_6081;
wire n_6082;
wire n_6083;
wire n_6084;
wire n_6085;
wire n_6086;
wire n_6087;
wire n_6088;
wire n_6089;
wire n_6090;
wire n_6091;
wire n_6092;
wire n_6093;
wire n_6094;
wire n_6095;
wire n_6096;
wire n_6097;
wire n_6098;
wire n_6099;
wire n_6100;
wire n_6101;
wire n_6102;
wire n_6103;
wire n_6104;
wire n_6105;
wire n_6106;
wire n_6107;
wire n_6108;
wire n_6109;
wire n_6110;
wire n_6111;
wire n_6112;
wire n_6113;
wire n_6114;
wire n_6115;
wire n_6116;
wire n_6117;
wire n_6118;
wire n_6119;
wire n_6120;
wire n_6121;
wire n_6122;
wire n_6123;
wire n_6124;
wire n_6125;
wire n_6126;
wire n_6127;
wire n_6128;
wire n_6129;
wire n_6130;
wire n_6131;
wire n_6132;
wire n_6133;
wire n_6134;
wire n_6135;
wire n_6136;
wire n_6137;
wire n_6138;
wire n_6139;
wire n_6140;
wire n_6141;
wire n_6142;
wire n_6143;
wire n_6144;
wire n_6145;
wire n_6146;
wire n_6147;
wire n_6148;
wire n_6149;
wire n_6150;
wire n_6151;
wire n_6152;
wire n_6153;
wire n_6154;
wire n_6155;
wire n_6156;
wire n_6157;
wire n_6158;
wire n_6159;
wire n_6160;
wire n_6161;
wire n_6162;
wire n_6163;
wire n_6164;
wire n_6165;
wire n_6166;
wire n_6167;
wire n_6168;
wire n_6169;
wire n_6170;
wire n_6171;
wire n_6172;
wire n_6173;
wire n_6174;
wire n_6175;
wire n_6176;
wire n_6177;
wire n_6178;
wire n_6179;
wire n_6180;
wire n_6181;
wire n_6182;
wire n_6183;
wire n_6184;
wire n_6185;
wire n_6186;
wire n_6187;
wire n_6188;
wire n_6189;
wire n_6190;
wire n_6191;
wire n_6192;
wire n_6193;
wire n_6194;
wire n_6195;
wire n_6196;
wire n_6197;
wire n_6198;
wire n_6199;
wire n_6200;
wire n_6201;
wire n_6202;
wire n_6203;
wire n_6204;
wire n_6205;
wire n_6206;
wire n_6207;
wire n_6208;
wire n_6209;
wire n_6210;
wire n_6211;
wire n_6212;
wire n_6213;
wire n_6214;
wire n_6215;
wire n_6216;
wire n_6217;
wire n_6218;
wire n_6219;
wire n_6220;
wire n_6221;
wire n_6222;
wire n_6223;
wire n_6224;
wire n_6225;
wire n_6226;
wire n_6227;
wire n_6228;
wire n_6229;
wire n_6230;
wire n_6231;
wire n_6232;
wire n_6233;
wire n_6234;
wire n_6235;
wire n_6236;
wire n_6237;
wire n_6238;
wire n_6239;
wire n_6240;
wire n_6241;
wire n_6242;
wire n_6243;
wire n_6244;
wire n_6245;
wire n_6246;
wire n_6247;
wire n_6248;
wire n_6249;
wire n_6250;
wire n_6251;
wire n_6252;
wire n_6253;
wire n_6254;
wire n_6255;
wire n_6256;
wire n_6257;
wire n_6258;
wire n_6259;
wire n_6260;
wire n_6261;
wire n_6262;
wire n_6263;
wire n_6264;
wire n_6265;
wire n_6266;
wire n_6267;
wire n_6268;
wire n_6269;
wire n_6270;
wire n_6271;
wire n_6272;
wire n_6273;
wire n_6274;
wire n_6275;
wire n_6276;
wire n_6277;
wire n_6278;
wire n_6279;
wire n_6280;
wire n_6281;
wire n_6282;
wire n_6283;
wire n_6284;
wire n_6285;
wire n_6286;
wire n_6287;
wire n_6288;
wire n_6289;
wire n_6290;
wire n_6291;
wire n_6292;
wire n_6293;
wire n_6294;
wire n_6295;
wire n_6296;
wire n_6297;
wire n_6298;
wire n_6299;
wire n_6300;
wire n_6301;
wire n_6302;
wire n_6303;
wire n_6304;
wire n_6305;
wire n_6306;
wire n_6307;
wire n_6308;
wire n_6309;
wire n_6310;
wire n_6311;
wire n_6312;
wire n_6313;
wire n_6314;
wire n_6315;
wire n_6316;
wire n_6317;
wire n_6318;
wire n_6319;
wire n_6320;
wire n_6321;
wire n_6322;
wire n_6323;
wire n_6324;
wire n_6325;
wire n_6326;
wire n_6327;
wire n_6328;
wire n_6329;
wire n_6330;
wire n_6331;
wire n_6332;
wire n_6333;
wire n_6334;
wire n_6335;
wire n_6336;
wire n_6337;
wire n_6338;
wire n_6339;
wire n_6340;
wire n_6341;
wire n_6342;
wire n_6343;
wire n_6344;
wire n_6345;
wire n_6346;
wire n_6347;
wire n_6348;
wire n_6349;
wire n_6350;
wire n_6351;
wire n_6352;
wire n_6353;
wire n_6354;
wire n_6355;
wire n_6356;
wire n_6357;
wire n_6358;
wire n_6359;
wire n_6360;
wire n_6361;
wire n_6362;
wire n_6363;
wire n_6364;
wire n_6365;
wire n_6366;
wire n_6367;
wire n_6368;
wire n_6369;
wire n_6370;
wire n_6371;
wire n_6372;
wire n_6373;
wire n_6374;
wire n_6375;
wire n_6376;
wire n_6377;
wire n_6378;
wire n_6379;
wire n_6380;
wire n_6381;
wire n_6382;
wire n_6383;
wire n_6384;
wire n_6385;
wire n_6386;
wire n_6387;
wire n_6388;
wire n_6389;
wire n_6390;
wire n_6391;
wire n_6392;
wire n_6393;
wire n_6394;
wire n_6395;
wire n_6396;
wire n_6397;
wire n_6398;
wire n_6399;
wire n_6400;
wire n_6401;
wire n_6402;
wire n_6403;
wire n_6404;
wire n_6405;
wire n_6406;
wire n_6407;
wire n_6408;
wire n_6409;
wire n_6410;
wire n_6411;
wire n_6412;
wire n_6413;
wire n_6414;
wire n_6415;
wire n_6416;
wire n_6417;
wire n_6418;
wire n_6419;
wire n_6420;
wire n_6421;
wire n_6422;
wire n_6423;
wire n_6424;
wire n_6425;
wire n_6426;
wire n_6427;
wire n_6428;
wire n_6429;
wire n_6430;
wire n_6431;
wire n_6432;
wire n_6433;
wire n_6434;
wire n_6435;
wire n_6436;
wire n_6437;
wire n_6438;
wire n_6439;
wire n_6440;
wire n_6441;
wire n_6442;
wire n_6443;
wire n_6444;
wire n_6445;
wire n_6446;
wire n_6447;
wire n_6448;
wire n_6449;
wire n_6450;
wire n_6451;
wire n_6452;
wire n_6453;
wire n_6454;
wire n_6455;
wire n_6456;
wire n_6457;
wire n_6458;
wire n_6459;
wire n_6460;
wire n_6461;
wire n_6462;
wire n_6463;
wire n_6464;
wire n_6465;
wire n_6466;
wire n_6467;
wire n_6468;
wire n_6469;
wire n_6470;
wire n_6471;
wire n_6472;
wire n_6473;
wire n_6474;
wire n_6475;
wire n_6476;
wire n_6477;
wire n_6478;
wire n_6479;
wire n_6480;
wire n_6481;
wire n_6482;
wire n_6483;
wire n_6484;
wire n_6485;
wire n_6486;
wire n_6487;
wire n_6488;
wire n_6489;
wire n_6490;
wire n_6491;
wire n_6492;
wire n_6493;
wire n_6494;
wire n_6495;
wire n_6496;
wire n_6497;
wire n_6498;
wire n_6499;
wire n_6500;
wire n_6501;
wire n_6502;
wire n_6503;
wire n_6504;
wire n_6505;
wire n_6506;
wire n_6507;
wire n_6508;
wire n_6509;
wire n_6510;
wire n_6511;
wire n_6512;
wire n_6513;
wire n_6514;
wire n_6515;
wire n_6516;
wire n_6517;
wire n_6518;
wire n_6519;
wire n_6520;
wire n_6521;
wire n_6522;
wire n_6523;
wire n_6524;
wire n_6525;
wire n_6526;
wire n_6527;
wire n_6528;
wire n_6529;
wire n_6530;
wire n_6531;
wire n_6532;
wire n_6533;
wire n_6534;
wire n_6535;
wire n_6536;
wire n_6537;
wire n_6538;
wire n_6539;
wire n_6540;
wire n_6541;
wire n_6542;
wire n_6543;
wire n_6544;
wire n_6545;
wire n_6546;
wire n_6547;
wire n_6548;
wire n_6549;
wire n_6550;
wire n_6551;
wire n_6552;
wire n_6553;
wire n_6554;
wire n_6555;
wire n_6556;
wire n_6557;
wire n_6558;
wire n_6559;
wire n_6560;
wire n_6561;
wire n_6562;
wire n_6563;
wire n_6564;
wire n_6565;
wire n_6566;
wire n_6567;
wire n_6568;
wire n_6569;
wire n_6570;
wire n_6571;
wire n_6572;
wire n_6573;
wire n_6574;
wire n_6575;
wire n_6576;
wire n_6577;
wire n_6578;
wire n_6579;
wire n_6580;
wire n_6581;
wire n_6582;
wire n_6583;
wire n_6584;
wire n_6585;
wire n_6586;
wire n_6587;
wire n_6588;
wire n_6589;
wire n_6590;
wire n_6591;
wire n_6592;
wire n_6593;
wire n_6594;
wire n_6595;
wire n_6596;
wire n_6597;
wire n_6598;
wire n_6599;
wire n_6600;
wire n_6601;
wire n_6602;
wire n_6603;
wire n_6604;
wire n_6605;
wire n_6606;
wire n_6607;
wire n_6608;
wire n_6609;
wire n_6610;
wire n_6611;
wire n_6612;
wire n_6613;
wire n_6614;
wire n_6615;
wire n_6616;
wire n_6617;
wire n_6618;
wire n_6619;
wire n_6620;
wire n_6621;
wire n_6622;
wire n_6623;
wire n_6624;
wire n_6625;
wire n_6626;
wire n_6627;
wire n_6628;
wire n_6629;
wire n_6630;
wire n_6631;
wire n_6632;
wire n_6633;
wire n_6634;
wire n_6635;
wire n_6636;
wire n_6637;
wire n_6638;
wire n_6639;
wire n_6640;
wire n_6641;
wire n_6642;
wire n_6643;
wire n_6644;
wire n_6645;
wire n_6646;
wire n_6647;
wire n_6648;
wire n_6649;
wire n_6650;
wire n_6651;
wire n_6652;
wire n_6653;
wire n_6654;
wire n_6655;
wire n_6656;
wire n_6657;
wire n_6658;
wire n_6659;
wire n_6660;
wire n_6661;
wire n_6662;
wire n_6663;
wire n_6664;
wire n_6665;
wire n_6666;
wire n_6667;
wire n_6668;
wire n_6669;
wire n_6670;
wire n_6671;
wire n_6672;
wire n_6673;
wire n_6674;
wire n_6675;
wire n_6676;
wire n_6677;
wire n_6678;
wire n_6679;
wire n_6680;
wire n_6681;
wire n_6682;
wire n_6683;
wire n_6684;
wire n_6685;
wire n_6686;
wire n_6687;
wire n_6688;
wire n_6689;
wire n_6690;
wire n_6691;
wire n_6692;
wire n_6693;
wire n_6694;
wire n_6695;
wire n_6696;
wire n_6697;
wire n_6698;
wire n_6699;
wire n_6700;
wire n_6701;
wire n_6702;
wire n_6703;
wire n_6704;
wire n_6705;
wire n_6706;
wire n_6707;
wire n_6708;
wire n_6709;
wire n_6710;
wire n_6711;
wire n_6712;
wire n_6713;
wire n_6714;
wire n_6715;
wire n_6716;
wire n_6717;
wire n_6718;
wire n_6719;
wire n_6720;
wire n_6721;
wire n_6722;
wire n_6723;
wire n_6724;
wire n_6725;
wire n_6726;
wire n_6727;
wire n_6728;
wire n_6729;
wire n_6730;
wire n_6731;
wire n_6732;
wire n_6733;
wire n_6734;
wire n_6735;
wire n_6736;
wire n_6737;
wire n_6738;
wire n_6739;
wire n_6740;
wire n_6741;
wire n_6742;
wire n_6743;
wire n_6744;
wire n_6745;
wire n_6746;
wire n_6747;
wire n_6748;
wire n_6749;
wire n_6750;
wire n_6751;
wire n_6752;
wire n_6753;
wire n_6754;
wire n_6755;
wire n_6756;
wire n_6757;
wire n_6758;
wire n_6759;
wire n_6760;
wire n_6761;
wire n_6762;
wire n_6763;
wire n_6764;
wire n_6765;
wire n_6766;
wire n_6767;
wire n_6768;
wire n_6769;
wire n_6770;
wire n_6771;
wire n_6772;
wire n_6773;
wire n_6774;
wire n_6775;
wire n_6776;
wire n_6777;
wire n_6778;
wire n_6779;
wire n_6780;
wire n_6781;
wire n_6782;
wire n_6783;
wire n_6784;
wire n_6785;
wire n_6786;
wire n_6787;
wire n_6788;
wire n_6789;
wire n_6790;
wire n_6791;
wire n_6792;
wire n_6793;
wire n_6794;
wire n_6795;
wire n_6796;
wire n_6797;
wire n_6798;
wire n_6799;
wire n_6800;
wire n_6801;
wire n_6802;
wire n_6803;
wire n_6804;
wire n_6805;
wire n_6806;
wire n_6807;
wire n_6808;
wire n_6809;
wire n_6810;
wire n_6811;
wire n_6812;
wire n_6813;
wire n_6814;
wire n_6815;
wire n_6816;
wire n_6817;
wire n_6818;
wire n_6819;
wire n_6820;
wire n_6821;
wire n_6822;
wire n_6823;
wire n_6824;
wire n_6825;
wire n_6826;
wire n_6827;
wire n_6828;
wire n_6829;
wire n_6830;
wire n_6831;
wire n_6832;
wire n_6833;
wire n_6834;
wire n_6835;
wire n_6836;
wire n_6837;
wire n_6838;
wire n_6839;
wire n_6840;
wire n_6841;
wire n_6842;
wire n_6843;
wire n_6844;
wire n_6845;
wire n_6846;
wire n_6847;
wire n_6848;
wire n_6849;
wire n_6850;
wire n_6851;
wire n_6852;
wire n_6853;
wire n_6854;
wire n_6855;
wire n_6856;
wire n_6857;
wire n_6858;
wire n_6859;
wire n_6860;
wire n_6861;
wire n_6862;
wire n_6863;
wire n_6864;
wire n_6865;
wire n_6866;
wire n_6867;
wire n_6868;
wire n_6869;
wire n_6870;
wire n_6871;
wire n_6872;
wire n_6873;
wire n_6874;
wire n_6875;
wire n_6876;
wire n_6877;
wire n_6878;
wire n_6879;
wire n_6880;
wire n_6881;
wire n_6882;
wire n_6883;
wire n_6884;
wire n_6885;
wire n_6886;
wire n_6887;
wire n_6888;
wire n_6889;
wire n_6890;
wire n_6891;
wire n_6892;
wire n_6893;
wire n_6894;
wire n_6895;
wire n_6896;
wire n_6897;
wire n_6898;
wire n_6899;
wire n_6900;
wire n_6901;
wire n_6902;
wire n_6903;
wire n_6904;
wire n_6905;
wire n_6906;
wire n_6907;
wire n_6908;
wire n_6909;
wire n_6910;
wire n_6911;
wire n_6912;
wire n_6913;
wire n_6914;
wire n_6915;
wire n_6916;
wire n_6917;
wire n_6918;
wire n_6919;
wire n_6920;
wire n_6921;
wire n_6922;
wire n_6923;
wire n_6924;
wire n_6925;
wire n_6926;
wire n_6927;
wire n_6928;
wire n_6929;
wire n_6930;
wire n_6931;
wire n_6932;
wire n_6933;
wire n_6934;
wire n_6935;
wire n_6936;
wire n_6937;
wire n_6938;
wire n_6939;
wire n_6940;
wire n_6941;
wire n_6942;
wire n_6943;
wire n_6944;
wire n_6945;
wire n_6946;
wire n_6947;
wire n_6948;
wire n_6949;
wire n_6950;
wire n_6951;
wire n_6952;
wire n_6953;
wire n_6954;
wire n_6955;
wire n_6956;
wire n_6957;
wire n_6958;
wire n_6959;
wire n_6960;
wire n_6961;
wire n_6962;
wire n_6963;
wire n_6964;
wire n_6965;
wire n_6966;
wire n_6967;
wire n_6968;
wire n_6969;
wire n_6970;
wire n_6971;
wire n_6972;
wire n_6973;
wire n_6974;
wire n_6975;
wire n_6976;
wire n_6977;
wire n_6978;
wire n_6979;
wire n_6980;
wire n_6981;
wire n_6982;
wire n_6983;
wire n_6984;
wire n_6985;
wire n_6986;
wire n_6987;
wire n_6988;
wire n_6989;
wire n_6990;
wire n_6991;
wire n_6992;
wire n_6993;
wire n_6994;
wire n_6995;
wire n_6996;
wire n_6997;
wire n_6998;
wire n_6999;
wire n_7000;
wire n_7001;
wire n_7002;
wire n_7003;
wire n_7004;
wire n_7005;
wire n_7006;
wire n_7007;
wire n_7008;
wire n_7009;
wire n_7010;
wire n_7011;
wire n_7012;
wire n_7013;
wire n_7014;
wire n_7015;
wire n_7016;
wire n_7017;
wire n_7018;
wire n_7019;
wire n_7020;
wire n_7021;
wire n_7022;
wire n_7023;
wire n_7024;
wire n_7025;
wire n_7026;
wire n_7027;
wire n_7028;
wire n_7029;
wire n_7030;
wire n_7031;
wire n_7032;
wire n_7033;
wire n_7034;
wire n_7035;
wire n_7036;
wire n_7037;
wire n_7038;
wire n_7039;
wire n_7040;
wire n_7041;
wire n_7042;
wire n_7043;
wire n_7044;
wire n_7045;
wire n_7046;
wire n_7047;
wire n_7048;
wire n_7049;
wire n_7050;
wire n_7051;
wire n_7052;
wire n_7053;
wire n_7054;
wire n_7055;
wire n_7056;
wire n_7057;
wire n_7058;
wire n_7059;
wire n_7060;
wire n_7061;
wire n_7062;
wire n_7063;
wire n_7064;
wire n_7065;
wire n_7066;
wire n_7067;
wire n_7068;
wire n_7069;
wire n_7070;
wire n_7071;
wire n_7072;
wire n_7073;
wire n_7074;
wire n_7075;
wire n_7076;
wire n_7077;
wire n_7078;
wire n_7079;
wire n_7080;
wire n_7081;
wire n_7082;
wire n_7083;
wire n_7084;
wire n_7085;
wire n_7086;
wire n_7087;
wire n_7088;
wire n_7089;
wire n_7090;
wire n_7091;
wire n_7092;
wire n_7093;
wire n_7094;
wire n_7095;
wire n_7096;
wire n_7097;
wire n_7098;
wire n_7099;
wire n_7100;
wire n_7101;
wire n_7102;
wire n_7103;
wire n_7104;
wire n_7105;
wire n_7106;
wire n_7107;
wire n_7108;
wire n_7109;
wire n_7110;
wire n_7111;
wire n_7112;
wire n_7113;
wire n_7114;
wire n_7115;
wire n_7116;
wire n_7117;
wire n_7118;
wire n_7119;
wire n_7120;
wire n_7121;
wire n_7122;
wire n_7123;
wire n_7124;
wire n_7125;
wire n_7126;
wire n_7127;
wire n_7128;
wire n_7129;
wire n_7130;
wire n_7131;
wire n_7132;
wire n_7133;
wire n_7134;
wire n_7135;
wire n_7136;
wire n_7137;
wire n_7138;
wire n_7139;
wire n_7140;
wire n_7141;
wire n_7142;
wire n_7143;
wire n_7144;
wire n_7145;
wire n_7146;
wire n_7147;
wire n_7148;
wire n_7149;
wire n_7150;
wire n_7151;
wire n_7152;
wire n_7153;
wire n_7154;
wire n_7155;
wire n_7156;
wire n_7157;
wire n_7158;
wire n_7159;
wire n_7160;
wire n_7161;
wire n_7162;
wire n_7163;
wire n_7164;
wire n_7165;
wire n_7166;
wire n_7167;
wire n_7168;
wire n_7169;
wire n_7170;
wire n_7171;
wire n_7172;
wire n_7173;
wire n_7174;
wire n_7175;
wire n_7176;
wire n_7177;
wire n_7178;
wire n_7179;
wire n_7180;
wire n_7181;
wire n_7182;
wire n_7183;
wire n_7184;
wire n_7185;
wire n_7186;
wire n_7187;
wire n_7188;
wire n_7189;
wire n_7190;
wire n_7191;
wire n_7192;
wire n_7193;
wire n_7194;
wire n_7195;
wire n_7196;
wire n_7197;
wire n_7198;
wire n_7199;
wire n_7200;
wire n_7201;
wire n_7202;
wire n_7203;
wire n_7204;
wire n_7205;
wire n_7206;
wire n_7207;
wire n_7208;
wire n_7209;
wire n_7210;
wire n_7211;
wire n_7212;
wire n_7213;
wire n_7214;
wire n_7215;
wire n_7216;
wire n_7217;
wire n_7218;
wire n_7219;
wire n_7220;
wire n_7221;
wire n_7222;
wire n_7223;
wire n_7224;
wire n_7225;
wire n_7226;
wire n_7227;
wire n_7228;
wire n_7229;
wire n_7230;
wire n_7231;
wire n_7232;
wire n_7233;
wire n_7234;
wire n_7235;
wire n_7236;
wire n_7237;
wire n_7238;
wire n_7239;
wire n_7240;
wire n_7241;
wire n_7242;
wire n_7243;
wire n_7244;
wire n_7245;
wire n_7246;
wire n_7247;
wire n_7248;
wire n_7249;
wire n_7250;
wire n_7251;
wire n_7252;
wire n_7253;
wire n_7254;
wire n_7255;
wire n_7256;
wire n_7257;
wire n_7258;
wire n_7259;
wire n_7260;
wire n_7261;
wire n_7262;
wire n_7263;
wire n_7264;
wire n_7265;
wire n_7266;
wire n_7267;
wire n_7268;
wire n_7269;
wire n_7270;
wire n_7271;
wire n_7272;
wire n_7273;
wire n_7274;
wire n_7275;
wire n_7276;
wire n_7277;
wire n_7278;
wire n_7279;
wire n_7280;
wire n_7281;
wire n_7282;
wire n_7283;
wire n_7284;
wire n_7285;
wire n_7286;
wire n_7287;
wire n_7288;
wire n_7289;
wire n_7290;
wire n_7291;
wire n_7292;
wire n_7293;
wire n_7294;
wire n_7295;
wire n_7296;
wire n_7297;
wire n_7298;
wire n_7299;
wire n_7300;
wire n_7301;
wire n_7302;
wire n_7303;
wire n_7304;
wire n_7305;
wire n_7306;
wire n_7307;
wire n_7308;
wire n_7309;
wire n_7310;
wire n_7311;
wire n_7312;
wire n_7313;
wire n_7314;
wire n_7315;
wire n_7316;
wire n_7317;
wire n_7318;
wire n_7319;
wire n_7320;
wire n_7321;
wire n_7322;
wire n_7323;
wire n_7324;
wire n_7325;
wire n_7326;
wire n_7327;
wire n_7328;
wire n_7329;
wire n_7330;
wire n_7331;
wire n_7332;
wire n_7333;
wire n_7334;
wire n_7335;
wire n_7336;
wire n_7337;
wire n_7338;
wire n_7339;
wire n_7340;
wire n_7341;
wire n_7342;
wire n_7343;
wire n_7344;
wire n_7345;
wire n_7346;
wire n_7347;
wire n_7348;
wire n_7349;
wire n_7350;
wire n_7351;
wire n_7352;
wire n_7353;
wire n_7354;
wire n_7355;
wire n_7356;
wire n_7357;
wire n_7358;
wire n_7359;
wire n_7360;
wire n_7361;
wire n_7362;
wire n_7363;
wire n_7364;
wire n_7365;
wire n_7366;
wire n_7367;
wire n_7368;
wire n_7369;
wire n_7370;
wire n_7371;
wire n_7372;
wire n_7373;
wire n_7374;
wire n_7375;
wire n_7376;
wire n_7377;
wire n_7378;
wire n_7379;
wire n_7380;
wire n_7381;
wire n_7382;
wire n_7383;
wire n_7384;
wire n_7385;
wire n_7386;
wire n_7387;
wire n_7388;
wire n_7389;
wire n_7390;
wire n_7391;
wire n_7392;
wire n_7393;
wire n_7394;
wire n_7395;
wire n_7396;
wire n_7397;
wire n_7398;
wire n_7399;
wire n_7400;
wire n_7401;
wire n_7402;
wire n_7403;
wire n_7404;
wire n_7405;
wire n_7406;
wire n_7407;
wire n_7408;
wire n_7409;
wire n_7410;
wire n_7411;
wire n_7412;
wire n_7413;
wire n_7414;
wire n_7415;
wire n_7416;
wire n_7417;
wire n_7418;
wire n_7419;
wire n_7420;
wire n_7421;
wire n_7422;
wire n_7423;
wire n_7424;
wire n_7425;
wire n_7426;
wire n_7427;
wire n_7428;
wire n_7429;
wire n_7430;
wire n_7431;
wire n_7432;
wire n_7433;
wire n_7434;
wire n_7435;
wire n_7436;
wire n_7437;
wire n_7438;
wire n_7439;
wire n_7440;
wire n_7441;
wire n_7442;
wire n_7443;
wire n_7444;
wire n_7445;
wire n_7446;
wire n_7447;
wire n_7448;
wire n_7449;
wire n_7450;
wire n_7451;
wire n_7452;
wire n_7453;
wire n_7454;
wire n_7455;
wire n_7456;
wire n_7457;
wire n_7458;
wire n_7459;
wire n_7460;
wire n_7461;
wire n_7462;
wire n_7463;
wire n_7464;
wire n_7465;
wire n_7466;
wire n_7467;
wire n_7468;
wire n_7469;
wire n_7470;
wire n_7471;
wire n_7472;
wire n_7473;
wire n_7474;
wire n_7475;
wire n_7476;
wire n_7477;
wire n_7478;
wire n_7479;
wire n_7480;
wire n_7481;
wire n_7482;
wire n_7483;
wire n_7484;
wire n_7485;
wire n_7486;
wire n_7487;
wire n_7488;
wire n_7489;
wire n_7490;
wire n_7491;
wire n_7492;
wire n_7493;
wire n_7494;
wire n_7495;
wire n_7496;
wire n_7497;
wire n_7498;
wire n_7499;
wire n_7500;
wire n_7501;
wire n_7502;
wire n_7503;
wire n_7504;
wire n_7505;
wire n_7506;
wire n_7507;
wire n_7508;
wire n_7509;
wire n_7510;
wire n_7511;
wire n_7512;
wire n_7513;
wire n_7514;
wire n_7515;
wire n_7516;
wire n_7517;
wire n_7518;
wire n_7519;
wire n_7520;
wire n_7521;
wire n_7522;
wire n_7523;
wire n_7524;
wire n_7525;
wire n_7526;
wire n_7527;
wire n_7528;
wire n_7529;
wire n_7530;
wire n_7531;
wire n_7532;
wire n_7533;
wire n_7534;
wire n_7535;
wire n_7536;
wire n_7537;
wire n_7538;
wire n_7539;
wire n_7540;
wire n_7541;
wire n_7542;
wire n_7543;
wire n_7544;
wire n_7545;
wire n_7546;
wire n_7547;
wire n_7548;
wire n_7549;
wire n_7550;
wire n_7551;
wire n_7552;
wire n_7553;
wire n_7554;
wire n_7555;
wire n_7556;
wire n_7557;
wire n_7558;
wire n_7559;
wire n_7560;
wire n_7561;
wire n_7562;
wire n_7563;
wire n_7564;
wire n_7565;
wire n_7566;
wire n_7567;
wire n_7568;
wire n_7569;
wire n_7570;
wire n_7571;
wire n_7572;
wire n_7573;
wire n_7574;
wire n_7575;
wire n_7576;
wire n_7577;
wire n_7578;
wire n_7579;
wire n_7580;
wire n_7581;
wire n_7582;
wire n_7583;
wire n_7584;
wire n_7585;
wire n_7586;
wire n_7587;
wire n_7588;
wire n_7589;
wire n_7590;
wire n_7591;
wire n_7592;
wire n_7593;
wire n_7594;
wire n_7595;
wire n_7596;
wire n_7597;
wire n_7598;
wire n_7599;
wire n_7600;
wire n_7601;
wire n_7602;
wire n_7603;
wire n_7604;
wire n_7605;
wire n_7606;
wire n_7607;
wire n_7608;
wire n_7609;
wire n_7610;
wire n_7611;
wire n_7612;
wire n_7613;
wire n_7614;
wire n_7615;
wire n_7616;
wire n_7617;
wire n_7618;
wire n_7619;
wire n_7620;
wire n_7621;
wire n_7622;
wire n_7623;
wire n_7624;
wire n_7625;
wire n_7626;
wire n_7627;
wire n_7628;
wire n_7629;
wire n_7630;
wire n_7631;
wire n_7632;
wire n_7633;
wire n_7634;
wire n_7635;
wire n_7636;
wire n_7637;
wire n_7638;
wire n_7639;
wire n_7640;
wire n_7641;
wire n_7642;
wire n_7643;
wire n_7644;
wire n_7645;
wire n_7646;
wire n_7647;
wire n_7648;
wire n_7649;
wire n_7650;
wire n_7651;
wire n_7652;
wire n_7653;
wire n_7654;
wire n_7655;
wire n_7656;
wire n_7657;
wire n_7658;
wire n_7659;
wire n_7660;
wire n_7661;
wire n_7662;
wire n_7663;
wire n_7664;
wire n_7665;
wire n_7666;
wire n_7667;
wire n_7668;
wire n_7669;
wire n_7670;
wire n_7671;
wire n_7672;
wire n_7673;
wire n_7674;
wire n_7675;
wire n_7676;
wire n_7677;
wire n_7678;
wire n_7679;
wire n_7680;
wire n_7681;
wire n_7682;
wire n_7683;
wire n_7684;
wire n_7685;
wire n_7686;
wire n_7687;
wire n_7688;
wire n_7689;
wire n_7690;
wire n_7691;
wire n_7692;
wire n_7693;
wire n_7694;
wire n_7695;
wire n_7696;
wire n_7697;
wire n_7698;
wire n_7699;
wire n_7700;
wire n_7701;
wire n_7702;
wire n_7703;
wire n_7704;
wire n_7705;
wire n_7706;
wire n_7707;
wire n_7708;
wire n_7709;
wire n_7710;
wire n_7711;
wire n_7712;
wire n_7713;
wire n_7714;
wire n_7715;
wire n_7716;
wire n_7717;
wire n_7718;
wire n_7719;
wire n_7720;
wire n_7721;
wire n_7722;
wire n_7723;
wire n_7724;
wire n_7725;
wire n_7726;
wire n_7727;
wire n_7728;
wire n_7729;
wire n_7730;
wire n_7731;
wire n_7732;
wire n_7733;
wire n_7734;
wire n_7735;
wire n_7736;
wire n_7737;
wire n_7738;
wire n_7739;
wire n_7740;
wire n_7741;
wire n_7742;
wire n_7743;
wire n_7744;
wire n_7745;
wire n_7746;
wire n_7747;
wire n_7748;
wire n_7749;
wire n_7750;
wire n_7751;
wire n_7752;
wire n_7753;
wire n_7754;
wire n_7755;
wire n_7756;
wire n_7757;
wire n_7758;
wire n_7759;
wire n_7760;
wire n_7761;
wire n_7762;
wire n_7763;
wire n_7764;
wire n_7765;
wire n_7766;
wire n_7767;
wire n_7768;
wire n_7769;
wire n_7770;
wire n_7771;
wire n_7772;
wire n_7773;
wire n_7774;
wire n_7775;
wire n_7776;
wire n_7777;
wire n_7778;
wire n_7779;
wire n_7780;
wire n_7781;
wire n_7782;
wire n_7783;
wire n_7784;
wire n_7785;
wire n_7786;
wire n_7787;
wire n_7788;
wire n_7789;
wire n_7790;
wire n_7791;
wire n_7792;
wire n_7793;
wire n_7794;
wire n_7795;
wire n_7796;
wire n_7797;
wire n_7798;
wire n_7799;
wire n_7800;
wire n_7801;
wire n_7802;
wire n_7803;
wire n_7804;
wire n_7805;
wire n_7806;
wire n_7807;
wire n_7808;
wire n_7809;
wire n_7810;
wire n_7811;
wire n_7812;
wire n_7813;
wire n_7814;
wire n_7815;
wire n_7816;
wire n_7817;
wire n_7818;
wire n_7819;
wire n_7820;
wire n_7821;
wire n_7822;
wire n_7823;
wire n_7824;
wire n_7825;
wire n_7826;
wire n_7827;
wire n_7828;
wire n_7829;
wire n_7830;
wire n_7831;
wire n_7832;
wire n_7833;
wire n_7834;
wire n_7835;
wire n_7836;
wire n_7837;
wire n_7838;
wire n_7839;
wire n_7840;
wire n_7841;
wire n_7842;
wire n_7843;
wire n_7844;
wire n_7845;
wire n_7846;
wire n_7847;
wire n_7848;
wire n_7849;
wire n_7850;
wire n_7851;
wire n_7852;
wire n_7853;
wire n_7854;
wire n_7855;
wire n_7856;
wire n_7857;
wire n_7858;
wire n_7859;
wire n_7860;
wire n_7861;
wire n_7862;
wire n_7863;
wire n_7864;
wire n_7865;
wire n_7866;
wire n_7867;
wire n_7868;
wire n_7869;
wire n_7870;
wire n_7871;
wire n_7872;
wire n_7873;
wire n_7874;
wire n_7875;
wire n_7876;
wire n_7877;
wire n_7878;
wire n_7879;
wire n_7880;
wire n_7881;
wire n_7882;
wire n_7883;
wire n_7884;
wire n_7885;
wire n_7886;
wire n_7887;
wire n_7888;
wire n_7889;
wire n_7890;
wire n_7891;
wire n_7892;
wire n_7893;
wire n_7894;
wire n_7895;
wire n_7896;
wire n_7897;
wire n_7898;
wire n_7899;
wire n_7900;
wire n_7901;
wire n_7902;
wire n_7903;
wire n_7904;
wire n_7905;
wire n_7906;
wire n_7907;
wire n_7908;
wire n_7909;
wire n_7910;
wire n_7911;
wire n_7912;
wire n_7913;
wire n_7914;
wire n_7915;
wire n_7916;
wire n_7917;
wire n_7918;
wire n_7919;
wire n_7920;
wire n_7921;
wire n_7922;
wire n_7923;
wire n_7924;
wire n_7925;
wire n_7926;
wire n_7927;
wire n_7928;
wire n_7929;
wire n_7930;
wire n_7931;
wire n_7932;
wire n_7933;
wire n_7934;
wire n_7935;
wire n_7936;
wire n_7937;
wire n_7938;
wire n_7939;
wire n_7940;
wire n_7941;
wire n_7942;
wire n_7943;
wire n_7944;
wire n_7945;
wire n_7946;
wire n_7947;
wire n_7948;
wire n_7949;
wire n_7950;
wire n_7951;
wire n_7952;
wire n_7953;
wire n_7954;
wire n_7955;
wire n_7956;
wire n_7957;
wire n_7958;
wire n_7959;
wire n_7960;
wire n_7961;
wire n_7962;
wire n_7963;
wire n_7964;
wire n_7965;
wire n_7966;
wire n_7967;
wire n_7968;
wire n_7969;
wire n_7970;
wire n_7971;
wire n_7972;
wire n_7973;
wire n_7974;
wire n_7975;
wire n_7976;
wire n_7977;
wire n_7978;
wire n_7979;
wire n_7980;
wire n_7981;
wire n_7982;
wire n_7983;
wire n_7984;
wire n_7985;
wire n_7986;
wire n_7987;
wire n_7988;
wire n_7989;
wire n_7990;
wire n_7991;
wire n_7992;
wire n_7993;
wire n_7994;
wire n_7995;
wire n_7996;
wire n_7997;
wire n_7998;
wire n_7999;
wire n_8000;
wire n_8001;
wire n_8002;
wire n_8003;
wire n_8004;
wire n_8005;
wire n_8006;
wire n_8007;
wire n_8008;
wire n_8009;
wire n_8010;
wire n_8011;
wire n_8012;
wire n_8013;
wire n_8014;
wire n_8015;
wire n_8016;
wire n_8017;
wire n_8018;
wire n_8019;
wire n_8020;
wire n_8021;
wire n_8022;
wire n_8023;
wire n_8024;
wire n_8025;
wire n_8026;
wire n_8027;
wire n_8028;
wire n_8029;
wire n_8030;
wire n_8031;
wire n_8032;
wire n_8033;
wire n_8034;
wire n_8035;
wire n_8036;
wire n_8037;
wire n_8038;
wire n_8039;
wire n_8040;
wire n_8041;
wire n_8042;
wire n_8043;
wire n_8044;
wire n_8045;
wire n_8046;
wire n_8047;
wire n_8048;
wire n_8049;
wire n_8050;
wire n_8051;
wire n_8052;
wire n_8053;
wire n_8054;
wire n_8055;
wire n_8056;
wire n_8057;
wire n_8058;
wire n_8059;
wire n_8060;
wire n_8061;
wire n_8062;
wire n_8063;
wire n_8064;
wire n_8065;
wire n_8066;
wire n_8067;
wire n_8068;
wire n_8069;
wire n_8070;
wire n_8071;
wire n_8072;
wire n_8073;
wire n_8074;
wire n_8075;
wire n_8076;
wire n_8077;
wire n_8078;
wire n_8079;
wire n_8080;
wire n_8081;
wire n_8082;
wire n_8083;
wire n_8084;
wire n_8085;
wire n_8086;
wire n_8087;
wire n_8088;
wire n_8089;
wire n_8090;
wire n_8091;
wire n_8092;
wire n_8093;
wire n_8094;
wire n_8095;
wire n_8096;
wire n_8097;
wire n_8098;
wire n_8099;
wire n_8100;
wire n_8101;
wire n_8102;
wire n_8103;
wire n_8104;
wire n_8105;
wire n_8106;
wire n_8107;
wire n_8108;
wire n_8109;
wire n_8110;
wire n_8111;
wire n_8112;
wire n_8113;
wire n_8114;
wire n_8115;
wire n_8116;
wire n_8117;
wire n_8118;
wire n_8119;
wire n_8120;
wire n_8121;
wire n_8122;
wire n_8123;
wire n_8124;
wire n_8125;
wire n_8126;
wire n_8127;
wire n_8128;
wire n_8129;
wire n_8130;
wire n_8131;
wire n_8132;
wire n_8133;
wire n_8134;
wire n_8135;
wire n_8136;
wire n_8137;
wire n_8138;
wire n_8139;
wire n_8140;
wire n_8141;
wire n_8142;
wire n_8143;
wire n_8144;
wire n_8145;
wire n_8146;
wire n_8147;
wire n_8148;
wire n_8149;
wire n_8150;
wire n_8151;
wire n_8152;
wire n_8153;
wire n_8154;
wire n_8155;
wire n_8156;
wire n_8157;
wire n_8158;
wire n_8159;
wire n_8160;
wire n_8161;
wire n_8162;
wire n_8163;
wire n_8164;
wire n_8165;
wire n_8166;
wire n_8167;
wire n_8168;
wire n_8169;
wire n_8170;
wire n_8171;
wire n_8172;
wire n_8173;
wire n_8174;
wire n_8175;
wire n_8176;
wire n_8177;
wire n_8178;
wire n_8179;
wire n_8180;
wire n_8181;
wire n_8182;
wire n_8183;
wire n_8184;
wire n_8185;
wire n_8186;
wire n_8187;
wire n_8188;
wire n_8189;
wire n_8190;
wire n_8191;
wire n_8192;
wire n_8193;
wire n_8194;
wire n_8195;
wire n_8196;
wire n_8197;
wire n_8198;
wire n_8199;
wire n_8200;
wire n_8201;
wire n_8202;
wire n_8203;
wire n_8204;
wire n_8205;
wire n_8206;
wire n_8207;
wire n_8208;
wire n_8209;
wire n_8210;
wire n_8211;
wire n_8212;
wire n_8213;
wire n_8214;
wire n_8215;
wire n_8216;
wire n_8217;
wire n_8218;
wire n_8219;
wire n_8220;
wire n_8221;
wire n_8222;
wire n_8223;
wire n_8224;
wire n_8225;
wire n_8226;
wire n_8227;
wire n_8228;
wire n_8229;
wire n_8230;
wire n_8231;
wire n_8232;
wire n_8233;
wire n_8234;
wire n_8235;
wire n_8236;
wire n_8237;
wire n_8238;
wire n_8239;
wire n_8240;
wire n_8241;
wire n_8242;
wire n_8243;
wire n_8244;
wire n_8245;
wire n_8246;
wire n_8247;
wire n_8248;
wire n_8249;
wire n_8250;
wire n_8251;
wire n_8252;
wire n_8253;
wire n_8254;
wire n_8255;
wire n_8256;
wire n_8257;
wire n_8258;
wire n_8259;
wire n_8260;
wire n_8261;
wire n_8262;
wire n_8263;
wire n_8264;
wire n_8265;
wire n_8266;
wire n_8267;
wire n_8268;
wire n_8269;
wire n_8270;
wire n_8271;
wire n_8272;
wire n_8273;
wire n_8274;
wire n_8275;
wire n_8276;
wire n_8277;
wire n_8278;
wire n_8279;
wire n_8280;
wire n_8281;
wire n_8282;
wire n_8283;
wire n_8284;
wire n_8285;
wire n_8286;
wire n_8287;
wire n_8288;
wire n_8289;
wire n_8290;
wire n_8291;
wire n_8292;
wire n_8293;
wire n_8294;
wire n_8295;
wire n_8296;
wire n_8297;
wire n_8298;
wire n_8299;
wire n_8300;
wire n_8301;
wire n_8302;
wire n_8303;
wire n_8304;
wire n_8305;
wire n_8306;
wire n_8307;
wire n_8308;
wire n_8309;
wire n_8310;
wire n_8311;
wire n_8312;
wire n_8313;
wire n_8314;
wire n_8315;
wire n_8316;
wire n_8317;
wire n_8318;
wire n_8319;
wire n_8320;
wire n_8321;
wire n_8322;
wire n_8323;
wire n_8324;
wire n_8325;
wire n_8326;
wire n_8327;
wire n_8328;
wire n_8329;
wire n_8330;
wire n_8331;
wire n_8332;
wire n_8333;
wire n_8334;
wire n_8335;
wire n_8336;
wire n_8337;
wire n_8338;
wire n_8339;
wire n_8340;
wire n_8341;
wire n_8342;
wire n_8343;
wire n_8344;
wire n_8345;
wire n_8346;
wire n_8347;
wire n_8348;
wire n_8349;
wire n_8350;
wire n_8351;
wire n_8352;
wire n_8353;
wire n_8354;
wire n_8355;
wire n_8356;
wire n_8357;
wire n_8358;
wire n_8359;
wire n_8360;
wire n_8361;
wire n_8362;
wire n_8363;
wire n_8364;
wire n_8365;
wire n_8366;
wire n_8367;
wire n_8368;
wire n_8369;
wire n_8370;
wire n_8371;
wire n_8372;
wire n_8373;
wire n_8374;
wire n_8375;
wire n_8376;
wire n_8377;
wire n_8378;
wire n_8379;
wire n_8380;
wire n_8381;
wire n_8382;
wire n_8383;
wire n_8384;
wire n_8385;
wire n_8386;
wire n_8387;
wire n_8388;
wire n_8389;
wire n_8390;
wire n_8391;
wire n_8392;
wire n_8393;
wire n_8394;
wire n_8395;
wire n_8396;
wire n_8397;
wire n_8398;
wire n_8399;
wire n_8400;
wire n_8401;
wire n_8402;
wire n_8403;
wire n_8404;
wire n_8405;
wire n_8406;
wire n_8407;
wire n_8408;
wire n_8409;
wire n_8410;
wire n_8411;
wire n_8412;
wire n_8413;
wire n_8414;
wire n_8415;
wire n_8416;
wire n_8417;
wire n_8418;
wire n_8419;
wire n_8420;
wire n_8421;
wire n_8422;
wire n_8423;
wire n_8424;
wire n_8425;
wire n_8426;
wire n_8427;
wire n_8428;
wire n_8429;
wire n_8430;
wire n_8431;
wire n_8432;
wire n_8433;
wire n_8434;
wire n_8435;
wire n_8436;
wire n_8437;
wire n_8438;
wire n_8439;
wire n_8440;
wire n_8441;
wire n_8442;
wire n_8443;
wire n_8444;
wire n_8445;
wire n_8446;
wire n_8447;
wire n_8448;
wire n_8449;
wire n_8450;
wire n_8451;
wire n_8452;
wire n_8453;
wire n_8454;
wire n_8455;
wire n_8456;
wire n_8457;
wire n_8458;
wire n_8459;
wire n_8460;
wire n_8461;
wire n_8462;
wire n_8463;
wire n_8464;
wire n_8465;
wire n_8466;
wire n_8467;
wire n_8468;
wire n_8469;
wire n_8470;
wire n_8471;
wire n_8472;
wire n_8473;
wire n_8474;
wire n_8475;
wire n_8476;
wire n_8477;
wire n_8478;
wire n_8479;
wire n_8480;
wire n_8481;
wire n_8482;
wire n_8483;
wire n_8484;
wire n_8485;
wire n_8486;
wire n_8487;
wire n_8488;
wire n_8489;
wire n_8490;
wire n_8491;
wire n_8492;
wire n_8493;
wire n_8494;
wire n_8495;
wire n_8496;
wire n_8497;
wire n_8498;
wire n_8499;
wire n_8500;
wire n_8501;
wire n_8502;
wire n_8503;
wire n_8504;
wire n_8505;
wire n_8506;
wire n_8507;
wire n_8508;
wire n_8509;
wire n_8510;
wire n_8511;
wire n_8512;
wire n_8513;
wire n_8514;
wire n_8515;
wire n_8516;
wire n_8517;
wire n_8518;
wire n_8519;
wire n_8520;
wire n_8521;
wire n_8522;
wire n_8523;
wire n_8524;
wire n_8525;
wire n_8526;
wire n_8527;
wire n_8528;
wire n_8529;
wire n_8530;
wire n_8531;
wire n_8532;
wire n_8533;
wire n_8534;
wire n_8535;
wire n_8536;
wire n_8537;
wire n_8538;
wire n_8539;
wire n_8540;
wire n_8541;
wire n_8542;
wire n_8543;
wire n_8544;
wire n_8545;
wire n_8546;
wire n_8547;
wire n_8548;
wire n_8549;
wire n_8550;
wire n_8551;
wire n_8552;
wire n_8553;
wire n_8554;
wire n_8555;
wire n_8556;
wire n_8557;
wire n_8558;
wire n_8559;
wire n_8560;
wire n_8561;
wire n_8562;
wire n_8563;
wire n_8564;
wire n_8565;
wire n_8566;
wire n_8567;
wire n_8568;
wire n_8569;
wire n_8570;
wire n_8571;
wire n_8572;
wire n_8573;
wire n_8574;
wire n_8575;
wire n_8576;
wire n_8577;
wire n_8578;
wire n_8579;
wire n_8580;
wire n_8581;
wire n_8582;
wire n_8583;
wire n_8584;
wire n_8585;
wire n_8586;
wire n_8587;
wire n_8588;
wire n_8589;
wire n_8590;
wire n_8591;
wire n_8592;
wire n_8593;
wire n_8594;
wire n_8595;
wire n_8596;
wire n_8597;
wire n_8598;
wire n_8599;
wire n_8600;
wire n_8601;
wire n_8602;
wire n_8603;
wire n_8604;
wire n_8605;
wire n_8606;
wire n_8607;
wire n_8608;
wire n_8609;
wire n_8610;
wire n_8611;
wire n_8612;
wire n_8613;
wire n_8614;
wire n_8615;
wire n_8616;
wire n_8617;
wire n_8618;
wire n_8619;
wire n_8620;
wire n_8621;
wire n_8622;
wire n_8623;
wire n_8624;
wire n_8625;
wire n_8626;
wire n_8627;
wire n_8628;
wire n_8629;
wire n_8630;
wire n_8631;
wire n_8632;
wire n_8633;
wire n_8634;
wire n_8635;
wire n_8636;
wire n_8637;
wire n_8638;
wire n_8639;
wire n_8640;
wire n_8641;
wire n_8642;
wire n_8643;
wire n_8644;
wire n_8645;
wire n_8646;
wire n_8647;
wire n_8648;
wire n_8649;
wire n_8650;
wire n_8651;
wire n_8652;
wire n_8653;
wire n_8654;
wire n_8655;
wire n_8656;
wire n_8657;
wire n_8658;
wire n_8659;
wire n_8660;
wire n_8661;
wire n_8662;
wire n_8663;
wire n_8664;
wire n_8665;
wire n_8666;
wire n_8667;
wire n_8668;
wire n_8669;
wire n_8670;
wire n_8671;
wire n_8672;
wire n_8673;
wire n_8674;
wire n_8675;
wire n_8676;
wire n_8677;
wire n_8678;
wire n_8679;
wire n_8680;
wire n_8681;
wire n_8682;
wire n_8683;
wire n_8684;
wire n_8685;
wire n_8686;
wire n_8687;
wire n_8688;
wire n_8689;
wire n_8690;
wire n_8691;
wire n_8692;
wire n_8693;
wire n_8694;
wire n_8695;
wire n_8696;
wire n_8697;
wire n_8698;
wire n_8699;
wire n_8700;
wire n_8701;
wire n_8702;
wire n_8703;
wire n_8704;
wire n_8705;
wire n_8706;
wire n_8707;
wire n_8708;
wire n_8709;
wire n_8710;
wire n_8711;
wire n_8712;
wire n_8713;
wire n_8714;
wire n_8715;
wire n_8716;
wire n_8717;
wire n_8718;
wire n_8719;
wire n_8720;
wire n_8721;
wire n_8722;
wire n_8723;
wire n_8724;
wire n_8725;
wire n_8726;
wire n_8727;
wire n_8728;
wire n_8729;
wire n_8730;
wire n_8731;
wire n_8732;
wire n_8733;
wire n_8734;
wire n_8735;
wire n_8736;
wire n_8737;
wire n_8738;
wire n_8739;
wire n_8740;
wire n_8741;
wire n_8742;
wire n_8743;
wire n_8744;
wire n_8745;
wire n_8746;
wire n_8747;
wire n_8748;
wire n_8749;
wire n_8750;
wire n_8751;
wire n_8752;
wire n_8753;
wire n_8754;
wire n_8755;
wire n_8756;
wire n_8757;
wire n_8758;
wire n_8759;
wire n_8760;
wire n_8761;
wire n_8762;
wire n_8763;
wire n_8764;
wire n_8765;
wire n_8766;
wire n_8767;
wire n_8768;
wire n_8769;
wire n_8770;
wire n_8771;
wire n_8772;
wire n_8773;
wire n_8774;
wire n_8775;
wire n_8776;
wire n_8777;
wire n_8778;
wire n_8779;
wire n_8780;
wire n_8781;
wire n_8782;
wire n_8783;
wire n_8784;
wire n_8785;
wire n_8786;
wire n_8787;
wire n_8788;
wire n_8789;
wire n_8790;
wire n_8791;
wire n_8792;
wire n_8793;
wire n_8794;
wire n_8795;
wire n_8796;
wire n_8797;
wire n_8798;
wire n_8799;
wire n_8800;
wire n_8801;
wire n_8802;
wire n_8803;
wire n_8804;
wire n_8805;
wire n_8806;
wire n_8807;
wire n_8808;
wire n_8809;
wire n_8810;
wire n_8811;
wire n_8812;
wire n_8813;
wire n_8814;
wire n_8815;
wire n_8816;
wire n_8817;
wire n_8818;
wire n_8819;
wire n_8820;
wire n_8821;
wire n_8822;
wire n_8823;
wire n_8824;
wire n_8825;
wire n_8826;
wire n_8827;
wire n_8828;
wire n_8829;
wire n_8830;
wire n_8831;
wire n_8832;
wire n_8833;
wire n_8834;
wire n_8835;
wire n_8836;
wire n_8837;
wire n_8838;
wire n_8839;
wire n_8840;
wire n_8841;
wire n_8842;
wire n_8843;
wire n_8844;
wire n_8845;
wire n_8846;
wire n_8847;
wire n_8848;
wire n_8849;
wire n_8850;
wire n_8851;
wire n_8852;
wire n_8853;
wire n_8854;
wire n_8855;
wire n_8856;
wire n_8857;
wire n_8858;
wire n_8859;
wire n_8860;
wire n_8861;
wire n_8862;
wire n_8863;
wire n_8864;
wire n_8865;
wire n_8866;
wire n_8867;
wire n_8868;
wire n_8869;
wire n_8870;
wire n_8871;
wire n_8872;
wire n_8873;
wire n_8874;
wire n_8875;
wire n_8876;
wire n_8877;
wire n_8878;
wire n_8879;
wire n_8880;
wire n_8881;
wire n_8882;
wire n_8883;
wire n_8884;
wire n_8885;
wire n_8886;
wire n_8887;
wire n_8888;
wire n_8889;
wire n_8890;
wire n_8891;
wire n_8892;
wire n_8893;
wire n_8894;
wire n_8895;
wire n_8896;
wire n_8897;
wire n_8898;
wire n_8899;
wire n_8900;
wire n_8901;
wire n_8902;
wire n_8903;
wire n_8904;
wire n_8905;
wire n_8906;
wire n_8907;
wire n_8908;
wire n_8909;
wire n_8910;
wire n_8911;
wire n_8912;
wire n_8913;
wire n_8914;
wire n_8915;
wire n_8916;
wire n_8917;
wire n_8918;
wire n_8919;
wire n_8920;
wire n_8921;
wire n_8922;
wire n_8923;
wire n_8924;
wire n_8925;
wire n_8926;
wire n_8927;
wire n_8928;
wire n_8929;
wire n_8930;
wire n_8931;
wire n_8932;
wire n_8933;
wire n_8934;
wire n_8935;
wire n_8936;
wire n_8937;
wire n_8938;
wire n_8939;
wire n_8940;
wire n_8941;
wire n_8942;
wire n_8943;
wire n_8944;
wire n_8945;
wire n_8946;
wire n_8947;
wire n_8948;
wire n_8949;
wire n_8950;
wire n_8951;
wire n_8952;
wire n_8953;
wire n_8954;
wire n_8955;
wire n_8956;
wire n_8957;
wire n_8958;
wire n_8959;
wire n_8960;
wire n_8961;
wire n_8962;
wire n_8963;
wire n_8964;
wire n_8965;
wire n_8966;
wire n_8967;
wire n_8968;
wire n_8969;
wire n_8970;
wire n_8971;
wire n_8972;
wire n_8973;
wire n_8974;
wire n_8975;
wire n_8976;
wire n_8977;
wire n_8978;
wire n_8979;
wire n_8980;
wire n_8981;
wire n_8982;
wire n_8983;
wire n_8984;
wire n_8985;
wire n_8986;
wire n_8987;
wire n_8988;
wire n_8989;
wire n_8990;
wire n_8991;
wire n_8992;
wire n_8993;
wire n_8994;
wire n_8995;
wire n_8996;
wire n_8997;
wire n_8998;
wire n_8999;
wire n_9000;
wire n_9001;
wire n_9002;
wire n_9003;
wire n_9004;
wire n_9005;
wire n_9006;
wire n_9007;
wire n_9008;
wire n_9009;
wire n_9010;
wire n_9011;
wire n_9012;
wire n_9013;
wire n_9014;
wire n_9015;
wire n_9016;
wire n_9017;
wire n_9018;
wire n_9019;
wire n_9020;
wire n_9021;
wire n_9022;
wire n_9023;
wire n_9024;
wire n_9025;
wire n_9026;
wire n_9027;
wire n_9028;
wire n_9029;
wire n_9030;
wire n_9031;
wire n_9032;
wire n_9033;
wire n_9034;
wire n_9035;
wire n_9036;
wire n_9037;
wire n_9038;
wire n_9039;
wire n_9040;
wire n_9041;
wire n_9042;
wire n_9043;
wire n_9044;
wire n_9045;
wire n_9046;
wire n_9047;
wire n_9048;
wire n_9049;
wire n_9050;
wire n_9051;
wire n_9052;
wire n_9053;
wire n_9054;
wire n_9055;
wire n_9056;
wire n_9057;
wire n_9058;
wire n_9059;
wire n_9060;
wire n_9061;
wire n_9062;
wire n_9063;
wire n_9064;
wire n_9065;
wire n_9066;
wire n_9067;
wire n_9068;
wire n_9069;
wire n_9070;
wire n_9071;
wire n_9072;
wire n_9073;
wire n_9074;
wire n_9075;
wire n_9076;
wire n_9077;
wire n_9078;
wire n_9079;
wire n_9080;
wire n_9081;
wire n_9082;
wire n_9083;
wire n_9084;
wire n_9085;
wire n_9086;
wire n_9087;
wire n_9088;
wire n_9089;
wire n_9090;
wire n_9091;
wire n_9092;
wire n_9093;
wire n_9094;
wire n_9095;
wire n_9096;
wire n_9097;
wire n_9098;
wire n_9099;
wire n_9100;
wire n_9101;
wire n_9102;
wire n_9103;
wire n_9104;
wire n_9105;
wire n_9106;
wire n_9107;
wire n_9108;
wire n_9109;
wire n_9110;
wire n_9111;
wire n_9112;
wire n_9113;
wire n_9114;
wire n_9115;
wire n_9116;
wire n_9117;
wire n_9118;
wire n_9119;
wire n_9120;
wire n_9121;
wire n_9122;
wire n_9123;
wire n_9124;
wire n_9125;
wire n_9126;
wire n_9127;
wire n_9128;
wire n_9129;
wire n_9130;
wire n_9131;
wire n_9132;
wire n_9133;
wire n_9134;
wire n_9135;
wire n_9136;
wire n_9137;
wire n_9138;
wire n_9139;
wire n_9140;
wire n_9141;
wire n_9142;
wire n_9143;
wire n_9144;
wire n_9145;
wire n_9146;
wire n_9147;
wire n_9148;
wire n_9149;
wire n_9150;
wire n_9151;
wire n_9152;
wire n_9153;
wire n_9154;
wire n_9155;
wire n_9156;
wire n_9157;
wire n_9158;
wire n_9159;
wire n_9160;
wire n_9161;
wire n_9162;
wire n_9163;
wire n_9164;
wire n_9165;
wire n_9166;
wire n_9167;
wire n_9168;
wire n_9169;
wire n_9170;
wire n_9171;
wire n_9172;
wire n_9173;
wire n_9174;
wire n_9175;
wire n_9176;
wire n_9177;
wire n_9178;
wire n_9179;
wire n_9180;
wire n_9181;
wire n_9182;
wire n_9183;
wire n_9184;
wire n_9185;
wire n_9186;
wire n_9187;
wire n_9188;
wire n_9189;
wire n_9190;
wire n_9191;
wire n_9192;
wire n_9193;
wire n_9194;
wire n_9195;
wire n_9196;
wire n_9197;
wire n_9198;
wire n_9199;
wire n_9200;
wire n_9201;
wire n_9202;
wire n_9203;
wire n_9204;
wire n_9205;
wire n_9206;
wire n_9207;
wire n_9208;
wire n_9209;
wire n_9210;
wire n_9211;
wire n_9212;
wire n_9213;
wire n_9214;
wire n_9215;
wire n_9216;
wire n_9217;
wire n_9218;
wire n_9219;
wire n_9220;
wire n_9221;
wire n_9222;
wire n_9223;
wire n_9224;
wire n_9225;
wire n_9226;
wire n_9227;
wire n_9228;
wire n_9229;
wire n_9230;
wire n_9231;
wire n_9232;
wire n_9233;
wire n_9234;
wire n_9235;
wire n_9236;
wire n_9237;
wire n_9238;
wire n_9239;
wire n_9240;
wire n_9241;
wire n_9242;
wire n_9243;
wire n_9244;
wire n_9245;
wire n_9246;
wire n_9247;
wire n_9248;
wire n_9249;
wire n_9250;
wire n_9251;
wire n_9252;
wire n_9253;
wire n_9254;
wire n_9255;
wire n_9256;
wire n_9257;
wire n_9258;
wire n_9259;
wire n_9260;
wire n_9261;
wire n_9262;
wire n_9263;
wire n_9264;
wire n_9265;
wire n_9266;
wire n_9267;
wire n_9268;
wire n_9269;
wire n_9270;
wire n_9271;
wire n_9272;
wire n_9273;
wire n_9274;
wire n_9275;
wire n_9276;
wire n_9277;
wire n_9278;
wire n_9279;
wire n_9280;
wire n_9281;
wire n_9282;
wire n_9283;
wire n_9284;
wire n_9285;
wire n_9286;
wire n_9287;
wire n_9288;
wire n_9289;
wire n_9290;
wire n_9291;
wire n_9292;
wire n_9293;
wire n_9294;
wire n_9295;
wire n_9296;
wire n_9297;
wire n_9298;
wire n_9299;
wire n_9300;
wire n_9301;
wire n_9302;
wire n_9303;
wire n_9304;
wire n_9305;
wire n_9306;
wire n_9307;
wire n_9308;
wire n_9309;
wire n_9310;
wire n_9311;
wire n_9312;
wire n_9313;
wire n_9314;
wire n_9315;
wire n_9316;
wire n_9317;
wire n_9318;
wire n_9319;
wire n_9320;
wire n_9321;
wire n_9322;
wire n_9323;
wire n_9324;
wire n_9325;
wire n_9326;
wire n_9327;
wire n_9328;
wire n_9329;
wire n_9330;
wire n_9331;
wire n_9332;
wire n_9333;
wire n_9334;
wire n_9335;
wire n_9336;
wire n_9337;
wire n_9338;
wire n_9339;
wire n_9340;
wire n_9341;
wire n_9342;
wire n_9343;
wire n_9344;
wire n_9345;
wire n_9346;
wire n_9347;
wire n_9348;
wire n_9349;
wire n_9350;
wire n_9351;
wire n_9352;
wire n_9353;
wire n_9354;
wire n_9355;
wire n_9356;
wire n_9357;
wire n_9358;
wire n_9359;
wire n_9360;
wire n_9361;
wire n_9362;
wire n_9363;
wire n_9364;
wire n_9365;
wire n_9366;
wire n_9367;
wire n_9368;
wire n_9369;
wire n_9370;
wire n_9371;
wire n_9372;
wire n_9373;
wire n_9374;
wire n_9375;
wire n_9376;
wire n_9377;
wire n_9378;
wire n_9379;
wire n_9380;
wire n_9381;
wire n_9382;
wire n_9383;
wire n_9384;
wire n_9385;
wire n_9386;
wire n_9387;
wire n_9388;
wire n_9389;
wire n_9390;
wire n_9391;
wire n_9392;
wire n_9393;
wire n_9394;
wire n_9395;
wire n_9396;
wire n_9397;
wire n_9398;
wire n_9399;
wire n_9400;
wire n_9401;
wire n_9402;
wire n_9403;
wire n_9404;
wire n_9405;
wire n_9406;
wire n_9407;
wire n_9408;
wire n_9409;
wire n_9410;
wire n_9411;
wire n_9412;
wire n_9413;
wire n_9414;
wire n_9415;
wire n_9416;
wire n_9417;
wire n_9418;
wire n_9419;
wire n_9420;
wire n_9421;
wire n_9422;
wire n_9423;
wire n_9424;
wire n_9425;
wire n_9426;
wire n_9427;
wire n_9428;
wire n_9429;
wire n_9430;
wire n_9431;
wire n_9432;
wire n_9433;
wire n_9434;
wire n_9435;
wire n_9436;
wire n_9437;
wire n_9438;
wire n_9439;
wire n_9440;
wire n_9441;
wire n_9442;
wire n_9443;
wire n_9444;
wire n_9445;
wire n_9446;
wire n_9447;
wire n_9448;
wire n_9449;
wire n_9450;
wire n_9451;
wire n_9452;
wire n_9453;
wire n_9454;
wire n_9455;
wire n_9456;
wire n_9457;
wire n_9458;
wire n_9459;
wire n_9460;
wire n_9461;
wire n_9462;
wire n_9463;
wire n_9464;
wire n_9465;
wire n_9466;
wire n_9467;
wire n_9468;
wire n_9469;
wire n_9470;
wire n_9471;
wire n_9472;
wire n_9473;
wire n_9474;
wire n_9475;
wire n_9476;
wire n_9477;
wire n_9478;
wire n_9479;
wire n_9480;
wire n_9481;
wire n_9482;
wire n_9483;
wire n_9484;
wire n_9485;
wire n_9486;
wire n_9487;
wire n_9488;
wire n_9489;
wire n_9490;
wire n_9491;
wire n_9492;
wire n_9493;
wire n_9494;
wire n_9495;
wire n_9496;
wire n_9497;
wire n_9498;
wire n_9499;
wire n_9500;
wire n_9501;
wire n_9502;
wire n_9503;
wire n_9504;
wire n_9505;
wire n_9506;
wire n_9507;
wire n_9508;
wire n_9509;
wire n_9510;
wire n_9511;
wire n_9512;
wire n_9513;
wire n_9514;
wire n_9515;
wire n_9516;
wire n_9517;
wire n_9518;
wire n_9519;
wire n_9520;
wire n_9521;
wire n_9522;
wire n_9523;
wire n_9524;
wire n_9525;
wire n_9526;
wire n_9527;
wire n_9528;
wire n_9529;
wire n_9530;
wire n_9531;
wire n_9532;
wire n_9533;
wire n_9534;
wire n_9535;
wire n_9536;
wire n_9537;
wire n_9538;
wire n_9539;
wire n_9540;
wire n_9541;
wire n_9542;
wire n_9543;
wire n_9544;
wire n_9545;
wire n_9546;
wire n_9547;
wire n_9548;
wire n_9549;
wire n_9550;
wire n_9551;
wire n_9552;
wire n_9553;
wire n_9554;
wire n_9555;
wire n_9556;
wire n_9557;
wire n_9558;
wire n_9559;
wire n_9560;
wire n_9561;
wire n_9562;
wire n_9563;
wire n_9564;
wire n_9565;
wire n_9566;
wire n_9567;
wire n_9568;
wire n_9569;
wire n_9570;
wire n_9571;
wire n_9572;
wire n_9573;
wire n_9574;
wire n_9575;
wire n_9576;
wire n_9577;
wire n_9578;
wire n_9579;
wire n_9580;
wire n_9581;
wire n_9582;
wire n_9583;
wire n_9584;
wire n_9585;
wire n_9586;
wire n_9587;
wire n_9588;
wire n_9589;
wire n_9590;
wire n_9591;
wire n_9592;
wire n_9593;
wire n_9594;
wire n_9595;
wire n_9596;
wire n_9597;
wire n_9598;
wire n_9599;
wire n_9600;
wire n_9601;
wire n_9602;
wire n_9603;
wire n_9604;
wire n_9605;
wire n_9606;
wire n_9607;
wire n_9608;
wire n_9609;
wire n_9610;
wire n_9611;
wire n_9612;
wire n_9613;
wire n_9614;
wire n_9615;
wire n_9616;
wire n_9617;
wire n_9618;
wire n_9619;
wire n_9620;
wire n_9621;
wire n_9622;
wire n_9623;
wire n_9624;
wire n_9625;
wire n_9626;
wire n_9627;
wire n_9628;
wire n_9629;
wire n_9630;
wire n_9631;
wire n_9632;
wire n_9633;
wire n_9634;
wire n_9635;
wire n_9636;
wire n_9637;
wire n_9638;
wire n_9639;
wire n_9640;
wire n_9641;
wire n_9642;
wire n_9643;
wire n_9644;
wire n_9645;
wire n_9646;
wire n_9647;
wire n_9648;
wire n_9649;
wire n_9650;
wire n_9651;
wire n_9652;
wire n_9653;
wire n_9654;
wire n_9655;
wire n_9656;
wire n_9657;
wire n_9658;
wire n_9659;
wire n_9660;
wire n_9661;
wire n_9662;
wire n_9663;
wire n_9664;
wire n_9665;
wire n_9666;
wire n_9667;
wire n_9668;
wire n_9669;
wire n_9670;
wire n_9671;
wire n_9672;
wire n_9673;
wire n_9674;
wire n_9675;
wire n_9676;
wire n_9677;
wire n_9678;
wire n_9679;
wire n_9680;
wire n_9681;
wire n_9682;
wire n_9683;
wire n_9684;
wire n_9685;
wire n_9686;
wire n_9687;
wire n_9688;
wire n_9689;
wire n_9690;
wire n_9691;
wire n_9692;
wire n_9693;
wire n_9694;
wire n_9695;
wire n_9696;
wire n_9697;
wire n_9698;
wire n_9699;
wire n_9700;
wire n_9701;
wire n_9702;
wire n_9703;
wire n_9704;
wire n_9705;
wire n_9706;
wire n_9707;
wire n_9708;
wire n_9709;
wire n_9710;
wire n_9711;
wire n_9712;
wire n_9713;
wire n_9714;
wire n_9715;
wire n_9716;
wire n_9717;
wire n_9718;
wire n_9719;
wire n_9720;
wire n_9721;
wire n_9722;
wire n_9723;
wire n_9724;
wire n_9725;
wire n_9726;
wire n_9727;
wire n_9728;
wire n_9729;
wire n_9730;
wire n_9731;
wire n_9732;
wire n_9733;
wire n_9734;
wire n_9735;
wire n_9736;
wire n_9737;
wire n_9738;
wire n_9739;
wire n_9740;
wire n_9741;
wire n_9742;
wire n_9743;
wire n_9744;
wire n_9745;
wire n_9746;
wire n_9747;
wire n_9748;
wire n_9749;
wire n_9750;
wire n_9751;
wire n_9752;
wire n_9753;
wire n_9754;
wire n_9755;
wire n_9756;
wire n_9757;
wire n_9758;
wire n_9759;
wire n_9760;
wire n_9761;
wire n_9762;
wire n_9763;
wire n_9764;
wire n_9765;
wire n_9766;
wire n_9767;
wire n_9768;
wire n_9769;
wire n_9770;
wire n_9771;
wire n_9772;
wire n_9773;
wire n_9774;
wire n_9775;
wire n_9776;
wire n_9777;
wire n_9778;
wire n_9779;
wire n_9780;
wire n_9781;
wire n_9782;
wire n_9783;
wire n_9784;
wire n_9785;
wire n_9786;
wire n_9787;
wire n_9788;
wire n_9789;
wire n_9790;
wire n_9791;
wire n_9792;
wire n_9793;
wire n_9794;
wire n_9795;
wire n_9796;
wire n_9797;
wire n_9798;
wire n_9799;
wire n_9800;
wire n_9801;
wire n_9802;
wire n_9803;
wire n_9804;
wire n_9805;
wire n_9806;
wire n_9807;
wire n_9808;
wire n_9809;
wire n_9810;
wire n_9811;
wire n_9812;
wire n_9813;
wire n_9814;
wire n_9815;
wire n_9816;
wire n_9817;
wire n_9818;
wire n_9819;
wire n_9820;
wire n_9821;
wire n_9822;
wire n_9823;
wire n_9824;
wire n_9825;
wire n_9826;
wire n_9827;
wire n_9828;
wire n_9829;
wire n_9830;
wire n_9831;
wire n_9832;
wire n_9833;
wire n_9834;
wire n_9835;
wire n_9836;
wire n_9837;
wire n_9838;
wire n_9839;
wire n_9840;
wire n_9841;
wire n_9842;
wire n_9843;
wire n_9844;
wire n_9845;
wire n_9846;
wire n_9847;
wire n_9848;
wire n_9849;
wire n_9850;
wire n_9851;
wire n_9852;
wire n_9853;
wire n_9854;
wire n_9855;
wire n_9856;
wire n_9857;
wire n_9858;
wire n_9859;
wire n_9860;
wire n_9861;
wire n_9862;
wire n_9863;
wire n_9864;
wire n_9865;
wire n_9866;
wire n_9867;
wire n_9868;
wire n_9869;
wire n_9870;
wire n_9871;
wire n_9872;
wire n_9873;
wire n_9874;
wire n_9875;
wire n_9876;
wire n_9877;
wire n_9878;
wire n_9879;
wire n_9880;
wire n_9881;
wire n_9882;
wire n_9883;
wire n_9884;
wire n_9885;
wire n_9886;
wire n_9887;
wire n_9888;
wire n_9889;
wire n_9890;
wire n_9891;
wire n_9892;
wire n_9893;
wire n_9894;
wire n_9895;
wire n_9896;
wire n_9897;
wire n_9898;
wire n_9899;
wire n_9900;
wire n_9901;
wire n_9902;
wire n_9903;
wire n_9904;
wire n_9905;
wire n_9906;
wire n_9907;
wire n_9908;
wire n_9909;
wire n_9910;
wire n_9911;
wire n_9912;
wire n_9913;
wire n_9914;
wire n_9915;
wire n_9916;
wire n_9917;
wire n_9918;
wire n_9919;
wire n_9920;
wire n_9921;
wire n_9922;
wire n_9923;
wire n_9924;
wire n_9925;
wire n_9926;
wire n_9927;
wire n_9928;
wire n_9929;
wire n_9930;
wire n_9931;
wire n_9932;
wire n_9933;
wire n_9934;
wire n_9935;
wire n_9936;
wire n_9937;
wire n_9938;
wire n_9939;
wire n_9940;
wire n_9941;
wire n_9942;
wire n_9943;
wire n_9944;
wire n_9945;
wire n_9946;
wire n_9947;
wire n_9948;
wire n_9949;
wire n_9950;
wire n_9951;
wire n_9952;
wire n_9953;
wire n_9954;
wire n_9955;
wire n_9956;
wire n_9957;
wire n_9958;
wire n_9959;
wire n_9960;
wire n_9961;
wire n_9962;
wire n_9963;
wire n_9964;
wire n_9965;
wire n_9966;
wire n_9967;
wire n_9968;
wire n_9969;
wire n_9970;
wire n_9971;
wire n_9972;
wire n_9973;
wire n_9974;
wire n_9975;
wire n_9976;
wire n_9977;
wire n_9978;
wire n_9979;
wire n_9980;
wire n_9981;
wire n_9982;
wire n_9983;
wire n_9984;
wire n_9985;
wire n_9986;
wire n_9987;
wire n_9988;
wire n_9989;
wire n_9990;
wire n_9991;
wire n_9992;
wire n_9993;
wire n_9994;
wire n_9995;
wire n_9996;
wire n_9997;
wire n_9998;
wire n_9999;
wire n_10000;
wire n_10001;
wire n_10002;
wire n_10003;
wire n_10004;
wire n_10005;
wire n_10006;
wire n_10007;
wire n_10008;
wire n_10009;
wire n_10010;
wire n_10011;
wire n_10012;
wire n_10013;
wire n_10014;
wire n_10015;
wire n_10016;
wire n_10017;
wire n_10018;
wire n_10019;
wire n_10020;
wire n_10021;
wire n_10022;
wire n_10023;
wire n_10024;
wire n_10025;
wire n_10026;
wire n_10027;
wire n_10028;
wire n_10029;
wire n_10030;
wire n_10031;
wire n_10032;
wire n_10033;
wire n_10034;
wire n_10035;
wire n_10036;
wire n_10037;
wire n_10038;
wire n_10039;
wire n_10040;
wire n_10041;
wire n_10042;
wire n_10043;
wire n_10044;
wire n_10045;
wire n_10046;
wire n_10047;
wire n_10048;
wire n_10049;
wire n_10050;
wire n_10051;
wire n_10052;
wire n_10053;
wire n_10054;
wire n_10055;
wire n_10056;
wire n_10057;
wire n_10058;
wire n_10059;
wire n_10060;
wire n_10061;
wire n_10062;
wire n_10063;
wire n_10064;
wire n_10065;
wire n_10066;
wire n_10067;
wire n_10068;
wire n_10069;
wire n_10070;
wire n_10071;
wire n_10072;
wire n_10073;
wire n_10074;
wire n_10075;
wire n_10076;
wire n_10077;
wire n_10078;
wire n_10079;
wire n_10080;
wire n_10081;
wire n_10082;
wire n_10083;
wire n_10084;
wire n_10085;
wire n_10086;
wire n_10087;
wire n_10088;
wire n_10089;
wire n_10090;
wire n_10091;
wire n_10092;
wire n_10093;
wire n_10094;
wire n_10095;
wire n_10096;
wire n_10097;
wire n_10098;
wire n_10099;
wire n_10100;
wire n_10101;
wire n_10102;
wire n_10103;
wire n_10104;
wire n_10105;
wire n_10106;
wire n_10107;
wire n_10108;
wire n_10109;
wire n_10110;
wire n_10111;
wire n_10112;
wire n_10113;
wire n_10114;
wire n_10115;
wire n_10116;
wire n_10117;
wire n_10118;
wire n_10119;
wire n_10120;
wire n_10121;
wire n_10122;
wire n_10123;
wire n_10124;
wire n_10125;
wire n_10126;
wire n_10127;
wire n_10128;
wire n_10129;
wire n_10130;
wire n_10131;
wire n_10132;
wire n_10133;
wire n_10134;
wire n_10135;
wire n_10136;
wire n_10137;
wire n_10138;
wire n_10139;
wire n_10140;
wire n_10141;
wire n_10142;
wire n_10143;
wire n_10144;
wire n_10145;
wire n_10146;
wire n_10147;
wire n_10148;
wire n_10149;
wire n_10150;
wire n_10151;
wire n_10152;
wire n_10153;
wire n_10154;
wire n_10155;
wire n_10156;
wire n_10157;
wire n_10158;
wire n_10159;
wire n_10160;
wire n_10161;
wire n_10162;
wire n_10163;
wire n_10164;
wire n_10165;
wire n_10166;
wire n_10167;
wire n_10168;
wire n_10169;
wire n_10170;
wire n_10171;
wire n_10172;
wire n_10173;
wire n_10174;
wire n_10175;
wire n_10176;
wire n_10177;
wire n_10178;
wire n_10179;
wire n_10180;
wire n_10181;
wire n_10182;
wire n_10183;
wire n_10184;
wire n_10185;
wire n_10186;
wire n_10187;
wire n_10188;
wire n_10189;
wire n_10190;
wire n_10191;
wire n_10192;
wire n_10193;
wire n_10194;
wire n_10195;
wire n_10196;
wire n_10197;
wire n_10198;
wire n_10199;
wire n_10200;
wire n_10201;
wire n_10202;
wire n_10203;
wire n_10204;
wire n_10205;
wire n_10206;
wire n_10207;
wire n_10208;
wire n_10209;
wire n_10210;
wire n_10211;
wire n_10212;
wire n_10213;
wire n_10214;
wire n_10215;
wire n_10216;
wire n_10217;
wire n_10218;
wire n_10219;
wire n_10220;
wire n_10221;
wire n_10222;
wire n_10223;
wire n_10224;
wire n_10225;
wire n_10226;
wire n_10227;
wire n_10228;
wire n_10229;
wire n_10230;
wire n_10231;
wire n_10232;
wire n_10233;
wire n_10234;
wire n_10235;
wire n_10236;
wire n_10237;
wire n_10238;
wire n_10239;
wire n_10240;
wire n_10241;
wire n_10242;
wire n_10243;
wire n_10244;
wire n_10245;
wire n_10246;
wire n_10247;
wire n_10248;
wire n_10249;
wire n_10250;
wire n_10251;
wire n_10252;
wire n_10253;
wire n_10254;
wire n_10255;
wire n_10256;
wire n_10257;
wire n_10258;
wire n_10259;
wire n_10260;
wire n_10261;
wire n_10262;
wire n_10263;
wire n_10264;
wire n_10265;
wire n_10266;
wire n_10267;
wire n_10268;
wire n_10269;
wire n_10270;
wire n_10271;
wire n_10272;
wire n_10273;
wire n_10274;
wire n_10275;
wire n_10276;
wire n_10277;
wire n_10278;
wire n_10279;
wire n_10280;
wire n_10281;
wire n_10282;
wire n_10283;
wire n_10284;
wire n_10285;
wire n_10286;
wire n_10287;
wire n_10288;
wire n_10289;
wire n_10290;
wire n_10291;
wire n_10292;
wire n_10293;
wire n_10294;
wire n_10295;
wire n_10296;
wire n_10297;
wire n_10298;
wire n_10299;
wire n_10300;
wire n_10301;
wire n_10302;
wire n_10303;
wire n_10304;
wire n_10305;
wire n_10306;
wire n_10307;
wire n_10308;
wire n_10309;
wire n_10310;
wire n_10311;
wire n_10312;
wire n_10313;
wire n_10314;
wire n_10315;
wire n_10316;
wire n_10317;
wire n_10318;
wire n_10319;
wire n_10320;
wire n_10321;
wire n_10322;
wire n_10323;
wire n_10324;
wire n_10325;
wire n_10326;
wire n_10327;
wire n_10328;
wire n_10329;
wire n_10330;
wire n_10331;
wire n_10332;
wire n_10333;
wire n_10334;
wire n_10335;
wire n_10336;
wire n_10337;
wire n_10338;
wire n_10339;
wire n_10340;
wire n_10341;
wire n_10342;
wire n_10343;
wire n_10344;
wire n_10345;
wire n_10346;
wire n_10347;
wire n_10348;
wire n_10349;
wire n_10350;
wire n_10351;
wire n_10352;
wire n_10353;
wire n_10354;
wire n_10355;
wire n_10356;
wire n_10357;
wire n_10358;
wire n_10359;
wire n_10360;
wire n_10361;
wire n_10362;
wire n_10363;
wire n_10364;
wire n_10365;
wire n_10366;
wire n_10367;
wire n_10368;
wire n_10369;
wire n_10370;
wire n_10371;
wire n_10372;
wire n_10373;
wire n_10374;
wire n_10375;
wire n_10376;
wire n_10377;
wire n_10378;
wire n_10379;
wire n_10380;
wire n_10381;
wire n_10382;
wire n_10383;
wire n_10384;
wire n_10385;
wire n_10386;
wire n_10387;
wire n_10388;
wire n_10389;
wire n_10390;
wire n_10391;
wire n_10392;
wire n_10393;
wire n_10394;
wire n_10395;
wire n_10396;
wire n_10397;
wire n_10398;
wire n_10399;
wire n_10400;
wire n_10401;
wire n_10402;
wire n_10403;
wire n_10404;
wire n_10405;
wire n_10406;
wire n_10407;
wire n_10408;
wire n_10409;
wire n_10410;
wire n_10411;
wire n_10412;
wire n_10413;
wire n_10414;
wire n_10415;
wire n_10416;
wire n_10417;
wire n_10418;
wire n_10419;
wire n_10420;
wire n_10421;
wire n_10422;
wire n_10423;
wire n_10424;
wire n_10425;
wire n_10426;
wire n_10427;
wire n_10428;
wire n_10429;
wire n_10430;
wire n_10431;
wire n_10432;
wire n_10433;
wire n_10434;
wire n_10435;
wire n_10436;
wire n_10437;
wire n_10438;
wire n_10439;
wire n_10440;
wire n_10441;
wire n_10442;
wire n_10443;
wire n_10444;
wire n_10445;
wire n_10446;
wire n_10447;
wire n_10448;
wire n_10449;
wire n_10450;
wire n_10451;
wire n_10452;
wire n_10453;
wire n_10454;
wire n_10455;
wire n_10456;
wire n_10457;
wire n_10458;
wire n_10459;
wire n_10460;
wire n_10461;
wire n_10462;
wire n_10463;
wire n_10464;
wire n_10465;
wire n_10466;
wire n_10467;
wire n_10468;
wire n_10469;
wire n_10470;
wire n_10471;
wire n_10472;
wire n_10473;
wire n_10474;
wire n_10475;
wire n_10476;
wire n_10477;
wire n_10478;
wire n_10479;
wire n_10480;
wire n_10481;
wire n_10482;
wire n_10483;
wire n_10484;
wire n_10485;
wire n_10486;
wire n_10487;
wire n_10488;
wire n_10489;
wire n_10490;
wire n_10491;
wire n_10492;
wire n_10493;
wire n_10494;
wire n_10495;
wire n_10496;
wire n_10497;
wire n_10498;
wire n_10499;
wire n_10500;
wire n_10501;
wire n_10502;
wire n_10503;
wire n_10504;
wire n_10505;
wire n_10506;
wire n_10507;
wire n_10508;
wire n_10509;
wire n_10510;
wire n_10511;
wire n_10512;
wire n_10513;
wire n_10514;
wire n_10515;
wire n_10516;
wire n_10517;
wire n_10518;
wire n_10519;
wire n_10520;
wire n_10521;
wire n_10522;
wire n_10523;
wire n_10524;
wire n_10525;
wire n_10526;
wire n_10527;
wire n_10528;
wire n_10529;
wire n_10530;
wire n_10531;
wire n_10532;
wire n_10533;
wire n_10534;
wire n_10535;
wire n_10536;
wire n_10537;
wire n_10538;
wire n_10539;
wire n_10540;
wire n_10541;
wire n_10542;
wire n_10543;
wire n_10544;
wire n_10545;
wire n_10546;
wire n_10547;
wire n_10548;
wire n_10549;
wire n_10550;
wire n_10551;
wire n_10552;
wire n_10553;
wire n_10554;
wire n_10555;
wire n_10556;
wire n_10557;
wire n_10558;
wire n_10559;
wire n_10560;
wire n_10561;
wire n_10562;
wire n_10563;
wire n_10564;
wire n_10565;
wire n_10566;
wire n_10567;
wire n_10568;
wire n_10569;
wire n_10570;
wire n_10571;
wire n_10572;
wire n_10573;
wire n_10574;
wire n_10575;
wire n_10576;
wire n_10577;
wire n_10578;
wire n_10579;
wire n_10580;
wire n_10581;
wire n_10582;
wire n_10583;
wire n_10584;
wire n_10585;
wire n_10586;
wire n_10587;
wire n_10588;
wire n_10589;
wire n_10590;
wire n_10591;
wire n_10592;
wire n_10593;
wire n_10594;
wire n_10595;
wire n_10596;
wire n_10597;
wire n_10598;
wire n_10599;
wire n_10600;
wire n_10601;
wire n_10602;
wire n_10603;
wire n_10604;
wire n_10605;
wire n_10606;
wire n_10607;
wire n_10608;
wire n_10609;
wire n_10610;
wire n_10611;
wire n_10612;
wire n_10613;
wire n_10614;
wire n_10615;
wire n_10616;
wire n_10617;
wire n_10618;
wire n_10619;
wire n_10620;
wire n_10621;
wire n_10622;
wire n_10623;
wire n_10624;
wire n_10625;
wire n_10626;
wire n_10627;
wire n_10628;
wire n_10629;
wire n_10630;
wire n_10631;
wire n_10632;
wire n_10633;
wire n_10634;
wire n_10635;
wire n_10636;
wire n_10637;
wire n_10638;
wire n_10639;
wire n_10640;
wire n_10641;
wire n_10642;
wire n_10643;
wire n_10644;
wire n_10645;
wire n_10646;
wire n_10647;
wire n_10648;
wire n_10649;
wire n_10650;
wire n_10651;
wire n_10652;
wire n_10653;
wire n_10654;
wire n_10655;
wire n_10656;
wire n_10657;
wire n_10658;
wire n_10659;
wire n_10660;
wire n_10661;
wire n_10662;
wire n_10663;
wire n_10664;
wire n_10665;
wire n_10666;
wire n_10667;
wire n_10668;
wire n_10669;
wire n_10670;
wire n_10671;
wire n_10672;
wire n_10673;
wire n_10674;
wire n_10675;
wire n_10676;
wire n_10677;
wire n_10678;
wire n_10679;
wire n_10680;
wire n_10681;
wire n_10682;
wire n_10683;
wire n_10684;
wire n_10685;
wire n_10686;
wire n_10687;
wire n_10688;
wire n_10689;
wire n_10690;
wire n_10691;
wire n_10692;
wire n_10693;
wire n_10694;
wire n_10695;
wire n_10696;
wire n_10697;
wire n_10698;
wire n_10699;
wire n_10700;
wire n_10701;
wire n_10702;
wire n_10703;
wire n_10704;
wire n_10705;
wire n_10706;
wire n_10707;
wire n_10708;
wire n_10709;
wire n_10710;
wire n_10711;
wire n_10712;
wire n_10713;
wire n_10714;
wire n_10715;
wire n_10716;
wire n_10717;
wire n_10718;
wire n_10719;
wire n_10720;
wire n_10721;
wire n_10722;
wire n_10723;
wire n_10724;
wire n_10725;
wire n_10726;
wire n_10727;
wire n_10728;
wire n_10729;
wire n_10730;
wire n_10731;
wire n_10732;
wire n_10733;
wire n_10734;
wire n_10735;
wire n_10736;
wire n_10737;
wire n_10738;
wire n_10739;
wire n_10740;
wire n_10741;
wire n_10742;
wire n_10743;
wire n_10744;
wire n_10745;
wire n_10746;
wire n_10747;
wire n_10748;
wire n_10749;
wire n_10750;
wire n_10751;
wire n_10752;
wire n_10753;
wire n_10754;
wire n_10755;
wire n_10756;
wire n_10757;
wire n_10758;
wire n_10759;
wire n_10760;
wire n_10761;
wire n_10762;
wire n_10763;
wire n_10764;
wire n_10765;
wire n_10766;
wire n_10767;
wire n_10768;
wire n_10769;
wire n_10770;
wire n_10771;
wire n_10772;
wire n_10773;
wire n_10774;
wire n_10775;
wire n_10776;
wire n_10777;
wire n_10778;
wire n_10779;
wire n_10780;
wire n_10781;
wire n_10782;
wire n_10783;
wire n_10784;
wire n_10785;
wire n_10786;
wire n_10787;
wire n_10788;
wire n_10789;
wire n_10790;
wire n_10791;
wire n_10792;
wire n_10793;
wire n_10794;
wire n_10795;
wire n_10796;
wire n_10797;
wire n_10798;
wire n_10799;
wire n_10800;
wire n_10801;
wire n_10802;
wire n_10803;
wire n_10804;
wire n_10805;
wire n_10806;
wire n_10807;
wire n_10808;
wire n_10809;
wire n_10810;
wire n_10811;
wire n_10812;
wire n_10813;
wire n_10814;
wire n_10815;
wire n_10816;
wire n_10817;
wire n_10818;
wire n_10819;
wire n_10820;
wire n_10821;
wire n_10822;
wire n_10823;
wire n_10824;
wire n_10825;
wire n_10826;
wire n_10827;
wire n_10828;
wire n_10829;
wire n_10830;
wire n_10831;
wire n_10832;
wire n_10833;
wire n_10834;
wire n_10835;
wire n_10836;
wire n_10837;
wire n_10838;
wire n_10839;
wire n_10840;
wire n_10841;
wire n_10842;
wire n_10843;
wire n_10844;
wire n_10845;
wire n_10846;
wire n_10847;
wire n_10848;
wire n_10849;
wire n_10850;
wire n_10851;
wire n_10852;
wire n_10853;
wire n_10854;
wire n_10855;
wire n_10856;
wire n_10857;
wire n_10858;
wire n_10859;
wire n_10860;
wire n_10861;
wire n_10862;
wire n_10863;
wire n_10864;
wire n_10865;
wire n_10866;
wire n_10867;
wire n_10868;
wire n_10869;
wire n_10870;
wire n_10871;
wire n_10872;
wire n_10873;
wire n_10874;
wire n_10875;
wire n_10876;
wire n_10877;
wire n_10878;
wire n_10879;
wire n_10880;
wire n_10881;
wire n_10882;
wire n_10883;
wire n_10884;
wire n_10885;
wire n_10886;
wire n_10887;
wire n_10888;
wire n_10889;
wire n_10890;
wire n_10891;
wire n_10892;
wire n_10893;
wire n_10894;
wire n_10895;
wire n_10896;
wire n_10897;
wire n_10898;
wire n_10899;
wire n_10900;
wire n_10901;
wire n_10902;
wire n_10903;
wire n_10904;
wire n_10905;
wire n_10906;
wire n_10907;
wire n_10908;
wire n_10909;
wire n_10910;
wire n_10911;
wire n_10912;
wire n_10913;
wire n_10914;
wire n_10915;
wire n_10916;
wire n_10917;
wire n_10918;
wire n_10919;
wire n_10920;
wire n_10921;
wire n_10922;
wire n_10923;
wire n_10924;
wire n_10925;
wire n_10926;
wire n_10927;
wire n_10928;
wire n_10929;
wire n_10930;
wire n_10931;
wire n_10932;
wire n_10933;
wire n_10934;
wire n_10935;
wire n_10936;
wire n_10937;
wire n_10938;
wire n_10939;
wire n_10940;
wire n_10941;
wire n_10942;
wire n_10943;
wire n_10944;
wire n_10945;
wire n_10946;
wire n_10947;
wire n_10948;
wire n_10949;
wire n_10950;
wire n_10951;
wire n_10952;
wire n_10953;
wire n_10954;
wire n_10955;
wire n_10956;
wire n_10957;
wire n_10958;
wire n_10959;
wire n_10960;
wire n_10961;
wire n_10962;
wire n_10963;
wire n_10964;
wire n_10965;
wire n_10966;
wire n_10967;
wire n_10968;
wire n_10969;
wire n_10970;
wire n_10971;
wire n_10972;
wire n_10973;
wire n_10974;
wire n_10975;
wire n_10976;
wire n_10977;
wire n_10978;
wire n_10979;
wire n_10980;
wire n_10981;
wire n_10982;
wire n_10983;
wire n_10984;
wire n_10985;
wire n_10986;
wire n_10987;
wire n_10988;
wire n_10989;
wire n_10990;
wire n_10991;
wire n_10992;
wire n_10993;
wire n_10994;
wire n_10995;
wire n_10996;
wire n_10997;
wire n_10998;
wire n_10999;
wire n_11000;
wire n_11001;
wire n_11002;
wire n_11003;
wire n_11004;
wire n_11005;
wire n_11006;
wire n_11007;
wire n_11008;
wire n_11009;
wire n_11010;
wire n_11011;
wire n_11012;
wire n_11013;
wire n_11014;
wire n_11015;
wire n_11016;
wire n_11017;
wire n_11018;
wire n_11019;
wire n_11020;
wire n_11021;
wire n_11022;
wire n_11023;
wire n_11024;
wire n_11025;
wire n_11026;
wire n_11027;
wire n_11028;
wire n_11029;
wire n_11030;
wire n_11031;
wire n_11032;
wire n_11033;
wire n_11034;
wire n_11035;
wire n_11036;
wire n_11037;
wire n_11038;
wire n_11039;
wire n_11040;
wire n_11041;
wire n_11042;
wire n_11043;
wire n_11044;
wire n_11045;
wire n_11046;
wire n_11047;
wire n_11048;
wire n_11049;
wire n_11050;
wire n_11051;
wire n_11052;
wire n_11053;
wire n_11054;
wire n_11055;
wire n_11056;
wire n_11057;
wire n_11058;
wire n_11059;
wire n_11060;
wire n_11061;
wire n_11062;
wire n_11063;
wire n_11064;
wire n_11065;
wire n_11066;
wire n_11067;
wire n_11068;
wire n_11069;
wire n_11070;
wire n_11071;
wire n_11072;
wire n_11073;
wire n_11074;
wire n_11075;
wire n_11076;
wire n_11077;
wire n_11078;
wire n_11079;
wire n_11080;
wire n_11081;
wire n_11082;
wire n_11083;
wire n_11084;
wire n_11085;
wire n_11086;
wire n_11087;
wire n_11088;
wire n_11089;
wire n_11090;
wire n_11091;
wire n_11092;
wire n_11093;
wire n_11094;
wire n_11095;
wire n_11096;
wire n_11097;
wire n_11098;
wire n_11099;
wire n_11100;
wire n_11101;
wire n_11102;
wire n_11103;
wire n_11104;
wire n_11105;
wire n_11106;
wire n_11107;
wire n_11108;
wire n_11109;
wire n_11110;
wire n_11111;
wire n_11112;
wire n_11113;
wire n_11114;
wire n_11115;
wire n_11116;
wire n_11117;
wire n_11118;
wire n_11119;
wire n_11120;
wire n_11121;
wire n_11122;
wire n_11123;
wire n_11124;
wire n_11125;
wire n_11126;
wire n_11127;
wire n_11128;
wire n_11129;
wire n_11130;
wire n_11131;
wire n_11132;
wire n_11133;
wire n_11134;
wire n_11135;
wire n_11136;
wire n_11137;
wire n_11138;
wire n_11139;
wire n_11140;
wire n_11141;
wire n_11142;
wire n_11143;
wire n_11144;
wire n_11145;
wire n_11146;
wire n_11147;
wire n_11148;
wire n_11149;
wire n_11150;
wire n_11151;
wire n_11152;
wire n_11153;
wire n_11154;
wire n_11155;
wire n_11156;
wire n_11157;
wire n_11158;
wire n_11159;
wire n_11160;
wire n_11161;
wire n_11162;
wire n_11163;
wire n_11164;
wire n_11165;
wire n_11166;
wire n_11167;
wire n_11168;
wire n_11169;
wire n_11170;
wire n_11171;
wire n_11172;
wire n_11173;
wire n_11174;
wire n_11175;
wire n_11176;
wire n_11177;
wire n_11178;
wire n_11179;
wire n_11180;
wire n_11181;
wire n_11182;
wire n_11183;
wire n_11184;
wire n_11185;
wire n_11186;
wire n_11187;
wire n_11188;
wire n_11189;
wire n_11190;
wire n_11191;
wire n_11192;
wire n_11193;
wire n_11194;
wire n_11195;
wire n_11196;
wire n_11197;
wire n_11198;
wire n_11199;
wire n_11200;
wire n_11201;
wire n_11202;
wire n_11203;
wire n_11204;
wire n_11205;
wire n_11206;
wire n_11207;
wire n_11208;
wire n_11209;
wire n_11210;
wire n_11211;
wire n_11212;
wire n_11213;
wire n_11214;
wire n_11215;
wire n_11216;
wire n_11217;
wire n_11218;
wire n_11219;
wire n_11220;
wire n_11221;
wire n_11222;
wire n_11223;
wire n_11224;
wire n_11225;
wire n_11226;
wire n_11227;
wire n_11228;
wire n_11229;
wire n_11230;
wire n_11231;
wire n_11232;
wire n_11233;
wire n_11234;
wire n_11235;
wire n_11236;
wire n_11237;
wire n_11238;
wire n_11239;
wire n_11240;
wire n_11241;
wire n_11242;
wire n_11243;
wire n_11244;
wire n_11245;
wire n_11246;
wire n_11247;
wire n_11248;
wire n_11249;
wire n_11250;
wire n_11251;
wire n_11252;
wire n_11253;
wire n_11254;
wire n_11255;
wire n_11256;
wire n_11257;
wire n_11258;
wire n_11259;
wire n_11260;
wire n_11261;
wire n_11262;
wire n_11263;
wire n_11264;
wire n_11265;
wire n_11266;
wire n_11267;
wire n_11268;
wire n_11269;
wire n_11270;
wire n_11271;
wire n_11272;
wire n_11273;
wire n_11274;
wire n_11275;
wire n_11276;
wire n_11277;
wire n_11278;
wire n_11279;
wire n_11280;
wire n_11281;
wire n_11282;
wire n_11283;
wire n_11284;
wire n_11285;
wire n_11286;
wire n_11287;
wire n_11288;
wire n_11289;
wire n_11290;
wire n_11291;
wire n_11292;
wire n_11293;
wire n_11294;
wire n_11295;
wire n_11296;
wire n_11297;
wire n_11298;
wire n_11299;
wire n_11300;
wire n_11301;
wire n_11302;
wire n_11303;
wire n_11304;
wire n_11305;
wire n_11306;
wire n_11307;
wire n_11308;
wire n_11309;
wire n_11310;
wire n_11311;
wire n_11312;
wire n_11313;
wire n_11314;
wire n_11315;
wire n_11316;
wire n_11317;
wire n_11318;
wire n_11319;
wire n_11320;
wire n_11321;
wire n_11322;
wire n_11323;
wire n_11324;
wire n_11325;
wire n_11326;
wire n_11327;
wire n_11328;
wire n_11329;
wire n_11330;
wire n_11331;
wire n_11332;
wire n_11333;
wire n_11334;
wire n_11335;
wire n_11336;
wire n_11337;
wire n_11338;
wire n_11339;
wire n_11340;
wire n_11341;
wire n_11342;
wire n_11343;
wire n_11344;
wire n_11345;
wire n_11346;
wire n_11347;
wire n_11348;
wire n_11349;
wire n_11350;
wire n_11351;
wire n_11352;
wire n_11353;
wire n_11354;
wire n_11355;
wire n_11356;
wire n_11357;
wire n_11358;
wire n_11359;
wire n_11360;
wire n_11361;
wire n_11362;
wire n_11363;
wire n_11364;
wire n_11365;
wire n_11366;
wire n_11367;
wire n_11368;
wire n_11369;
wire n_11370;
wire n_11371;
wire n_11372;
wire n_11373;
wire n_11374;
wire n_11375;
wire n_11376;
wire n_11377;
wire n_11378;
wire n_11379;
wire n_11380;
wire n_11381;
wire n_11382;
wire n_11383;
wire n_11384;
wire n_11385;
wire n_11386;
wire n_11387;
wire n_11388;
wire n_11389;
wire n_11390;
wire n_11391;
wire n_11392;
wire n_11393;
wire n_11394;
wire n_11395;
wire n_11396;
wire n_11397;
wire n_11398;
wire n_11399;
wire n_11400;
wire n_11401;
wire n_11402;
wire n_11403;
wire n_11404;
wire n_11405;
wire n_11406;
wire n_11407;
wire n_11408;
wire n_11409;
wire n_11410;
wire n_11411;
wire n_11412;
wire n_11413;
wire n_11414;
wire n_11415;
wire n_11416;
wire n_11417;
wire n_11418;
wire n_11419;
wire n_11420;
wire n_11421;
wire n_11422;
wire n_11423;
wire n_11424;
wire n_11425;
wire n_11426;
wire n_11427;
wire n_11428;
wire n_11429;
wire n_11430;
wire n_11431;
wire n_11432;
wire n_11433;
wire n_11434;
wire n_11435;
wire n_11436;
wire n_11437;
wire n_11438;
wire n_11439;
wire n_11440;
wire n_11441;
wire n_11442;
wire n_11443;
wire n_11444;
wire n_11445;
wire n_11446;
wire n_11447;
wire n_11448;
wire n_11449;
wire n_11450;
wire n_11451;
wire n_11452;
wire n_11453;
wire n_11454;
wire n_11455;
wire n_11456;
wire n_11457;
wire n_11458;
wire n_11459;
wire n_11460;
wire n_11461;
wire n_11462;
wire n_11463;
wire n_11464;
wire n_11465;
wire n_11466;
wire n_11467;
wire n_11468;
wire n_11469;
wire n_11470;
wire n_11471;
wire n_11472;
wire n_11473;
wire n_11474;
wire n_11475;
wire n_11476;
wire n_11477;
wire n_11478;
wire n_11479;
wire n_11480;
wire n_11481;
wire n_11482;
wire n_11483;
wire n_11484;
wire n_11485;
wire n_11486;
wire n_11487;
wire n_11488;
wire n_11489;
wire n_11490;
wire n_11491;
wire n_11492;
wire n_11493;
wire n_11494;
wire n_11495;
wire n_11496;
wire n_11497;
wire n_11498;
wire n_11499;
wire n_11500;
wire n_11501;
wire n_11502;
wire n_11503;
wire n_11504;
wire n_11505;
wire n_11506;
wire n_11507;
wire n_11508;
wire n_11509;
wire n_11510;
wire n_11511;
wire n_11512;
wire n_11513;
wire n_11514;
wire n_11515;
wire n_11516;
wire n_11517;
wire n_11518;
wire n_11519;
wire n_11520;
wire n_11521;
wire n_11522;
wire n_11523;
wire n_11524;
wire n_11525;
wire n_11526;
wire n_11527;
wire n_11528;
wire n_11529;
wire n_11530;
wire n_11531;
wire n_11532;
wire n_11533;
wire n_11534;
wire n_11535;
wire n_11536;
wire n_11537;
wire n_11538;
wire n_11539;
wire n_11540;
wire n_11541;
wire n_11542;
wire n_11543;
wire n_11544;
wire n_11545;
wire n_11546;
wire n_11547;
wire n_11548;
wire n_11549;
wire n_11550;
wire n_11551;
wire n_11552;
wire n_11553;
wire n_11554;
wire n_11555;
wire n_11556;
wire n_11557;
wire n_11558;
wire n_11559;
wire n_11560;
wire n_11561;
wire n_11562;
wire n_11563;
wire n_11564;
wire n_11565;
wire n_11566;
wire n_11567;
wire n_11568;
wire n_11569;
wire n_11570;
wire n_11571;
wire n_11572;
wire n_11573;
wire n_11574;
wire n_11575;
wire n_11576;
wire n_11577;
wire n_11578;
wire n_11579;
wire n_11580;
wire n_11581;
wire n_11582;
wire n_11583;
wire n_11584;
wire n_11585;
wire n_11586;
wire n_11587;
wire n_11588;
wire n_11589;
wire n_11590;
wire n_11591;
wire n_11592;
wire n_11593;
wire n_11594;
wire n_11595;
wire n_11596;
wire n_11597;
wire n_11598;
wire n_11599;
wire n_11600;
wire n_11601;
wire n_11602;
wire n_11603;
wire n_11604;
wire n_11605;
wire n_11606;
wire n_11607;
wire n_11608;
wire n_11609;
wire n_11610;
wire n_11611;
wire n_11612;
wire n_11613;
wire n_11614;
wire n_11615;
wire n_11616;
wire n_11617;
wire n_11618;
wire n_11619;
wire n_11620;
wire n_11621;
wire n_11622;
wire n_11623;
wire n_11624;
wire n_11625;
wire n_11626;
wire n_11627;
wire n_11628;
wire n_11629;
wire n_11630;
wire n_11631;
wire n_11632;
wire n_11633;
wire n_11634;
wire n_11635;
wire n_11636;
wire n_11637;
wire n_11638;
wire n_11639;
wire n_11640;
wire n_11641;
wire n_11642;
wire n_11643;
wire n_11644;
wire n_11645;
wire n_11646;
wire n_11647;
wire n_11648;
wire n_11649;
wire n_11650;
wire n_11651;
wire n_11652;
wire n_11653;
wire n_11654;
wire n_11655;
wire n_11656;
wire n_11657;
wire n_11658;
wire n_11659;
wire n_11660;
wire n_11661;
wire n_11662;
wire n_11663;
wire n_11664;
wire n_11665;
wire n_11666;
wire n_11667;
wire n_11668;
wire n_11669;
wire n_11670;
wire n_11671;
wire n_11672;
wire n_11673;
wire n_11674;
wire n_11675;
wire n_11676;
wire n_11677;
wire n_11678;
wire n_11679;
wire n_11680;
wire n_11681;
wire n_11682;
wire n_11683;
wire n_11684;
wire n_11685;
wire n_11686;
wire n_11687;
wire n_11688;
wire n_11689;
wire n_11690;
wire n_11691;
wire n_11692;
wire n_11693;
wire n_11694;
wire n_11695;
wire n_11696;
wire n_11697;
wire n_11698;
wire n_11699;
wire n_11700;
wire n_11701;
wire n_11702;
wire n_11703;
wire n_11704;
wire n_11705;
wire n_11706;
wire n_11707;
wire n_11708;
wire n_11709;
wire n_11710;
wire n_11711;
wire n_11712;
wire n_11713;
wire n_11714;
wire n_11715;
wire n_11716;
wire n_11717;
wire n_11718;
wire n_11719;
wire n_11720;
wire n_11721;
wire n_11722;
wire n_11723;
wire n_11724;
wire n_11725;
wire n_11726;
wire n_11727;
wire n_11728;
wire n_11729;
wire n_11730;
wire n_11731;
wire n_11732;
wire n_11733;
wire n_11734;
wire n_11735;
wire n_11736;
wire n_11737;
wire n_11738;
wire n_11739;
wire n_11740;
wire n_11741;
wire n_11742;
wire n_11743;
wire n_11744;
wire n_11745;
wire n_11746;
wire n_11747;
wire n_11748;
wire n_11749;
wire n_11750;
wire n_11751;
wire n_11752;
wire n_11753;
wire n_11754;
wire n_11755;
wire n_11756;
wire n_11757;
wire n_11758;
wire n_11759;
wire n_11760;
wire n_11761;
wire n_11762;
wire n_11763;
wire n_11764;
wire n_11765;
wire n_11766;
wire n_11767;
wire n_11768;
wire n_11769;
wire n_11770;
wire n_11771;
wire n_11772;
wire n_11773;
wire n_11774;
wire n_11775;
wire n_11776;
wire n_11777;
wire n_11778;
wire n_11779;
wire n_11780;
wire n_11781;
wire n_11782;
wire n_11783;
wire n_11784;
wire n_11785;
wire n_11786;
wire n_11787;
wire n_11788;
wire n_11789;
wire n_11790;
wire n_11791;
wire n_11792;
wire n_11793;
wire n_11794;
wire n_11795;
wire n_11796;
wire n_11797;
wire n_11798;
wire n_11799;
wire n_11800;
wire n_11801;
wire n_11802;
wire n_11803;
wire n_11804;
wire n_11805;
wire n_11806;
wire n_11807;
wire n_11808;
wire n_11809;
wire n_11810;
wire n_11811;
wire n_11812;
wire n_11813;
wire n_11814;
wire n_11815;
wire n_11816;
wire n_11817;
wire n_11818;
wire n_11819;
wire n_11820;
wire n_11821;
wire n_11822;
wire n_11823;
wire n_11824;
wire n_11825;
wire n_11826;
wire n_11827;
wire n_11828;
wire n_11829;
wire n_11830;
wire n_11831;
wire n_11832;
wire n_11833;
wire n_11834;
wire n_11835;
wire n_11836;
wire n_11837;
wire n_11838;
wire n_11839;
wire n_11840;
wire n_11841;
wire n_11842;
wire n_11843;
wire n_11844;
wire n_11845;
wire n_11846;
wire n_11847;
wire n_11848;
wire n_11849;
wire n_11850;
wire n_11851;
wire n_11852;
wire n_11853;
wire n_11854;
wire n_11855;
wire n_11856;
wire n_11857;
wire n_11858;
wire n_11859;
wire n_11860;
wire n_11861;
wire n_11862;
wire n_11863;
wire n_11864;
wire n_11865;
wire n_11866;
wire n_11867;
wire n_11868;
wire n_11869;
wire n_11870;
wire n_11871;
wire n_11872;
wire n_11873;
wire n_11874;
wire n_11875;
wire n_11876;
wire n_11877;
wire n_11878;
wire n_11879;
wire n_11880;
wire n_11881;
wire n_11882;
wire n_11883;
wire n_11884;
wire n_11885;
wire n_11886;
wire n_11887;
wire n_11888;
wire n_11889;
wire n_11890;
wire n_11891;
wire n_11892;
wire n_11893;
wire n_11894;
wire n_11895;
wire n_11896;
wire n_11897;
wire n_11898;
wire n_11899;
wire n_11900;
wire n_11901;
wire n_11902;
wire n_11903;
wire n_11904;
wire n_11905;
wire n_11906;
wire n_11907;
wire n_11908;
wire n_11909;
wire n_11910;
wire n_11911;
wire n_11912;
wire n_11913;
wire n_11914;
wire n_11915;
wire n_11916;
wire n_11917;
wire n_11918;
wire n_11919;
wire n_11920;
wire n_11921;
wire n_11922;
wire n_11923;
wire n_11924;
wire n_11925;
wire n_11926;
wire n_11927;
wire n_11928;
wire n_11929;
wire n_11930;
wire n_11931;
wire n_11932;
wire n_11933;
wire n_11934;
wire n_11935;
wire n_11936;
wire n_11937;
wire n_11938;
wire n_11939;
wire n_11940;
wire n_11941;
wire n_11942;
wire n_11943;
wire n_11944;
wire n_11945;
wire n_11946;
wire n_11947;
wire n_11948;
wire n_11949;
wire n_11950;
wire n_11951;
wire n_11952;
wire n_11953;
wire n_11954;
wire n_11955;
wire n_11956;
wire n_11957;
wire n_11958;
wire n_11959;
wire n_11960;
wire n_11961;
wire n_11962;
wire n_11963;
wire n_11964;
wire n_11965;
wire n_11966;
wire n_11967;
wire n_11968;
wire n_11969;
wire n_11970;
wire n_11971;
wire n_11972;
wire n_11973;
wire n_11974;
wire n_11975;
wire n_11976;
wire n_11977;
wire n_11978;
wire n_11979;
wire n_11980;
wire n_11981;
wire n_11982;
wire n_11983;
wire n_11984;
wire n_11985;
wire n_11986;
wire n_11987;
wire n_11988;
wire n_11989;
wire n_11990;
wire n_11991;
wire n_11992;
wire n_11993;
wire n_11994;
wire n_11995;
wire n_11996;
wire n_11997;
wire n_11998;
wire n_11999;
wire n_12000;
wire n_12001;
wire n_12002;
wire n_12003;
wire n_12004;
wire n_12005;
wire n_12006;
wire n_12007;
wire n_12008;
wire n_12009;
wire n_12010;
wire n_12011;
wire n_12012;
wire n_12013;
wire n_12014;
wire n_12015;
wire n_12016;
wire n_12017;
wire n_12018;
wire n_12019;
wire n_12020;
wire n_12021;
wire n_12022;
wire n_12023;
wire n_12024;
wire n_12025;
wire n_12026;
wire n_12027;
wire n_12028;
wire n_12029;
wire n_12030;
wire n_12031;
wire n_12032;
wire n_12033;
wire n_12034;
wire n_12035;
wire n_12036;
wire n_12037;
wire n_12038;
wire n_12039;
wire n_12040;
wire n_12041;
wire n_12042;
wire n_12043;
wire n_12044;
wire n_12045;
wire n_12046;
wire n_12047;
wire n_12048;
wire n_12049;
wire n_12050;
wire n_12051;
wire n_12052;
wire n_12053;
wire n_12054;
wire n_12055;
wire n_12056;
wire n_12057;
wire n_12058;
wire n_12059;
wire n_12060;
wire n_12061;
wire n_12062;
wire n_12063;
wire n_12064;
wire n_12065;
wire n_12066;
wire n_12067;
wire n_12068;
wire n_12069;
wire n_12070;
wire n_12071;
wire n_12072;
wire n_12073;
wire n_12074;
wire n_12075;
wire n_12076;
wire n_12077;
wire n_12078;
wire n_12079;
wire n_12080;
wire n_12081;
wire n_12082;
wire n_12083;
wire n_12084;
wire n_12085;
wire n_12086;
wire n_12087;
wire n_12088;
wire n_12089;
wire n_12090;
wire n_12091;
wire n_12092;
wire n_12093;
wire n_12094;
wire n_12095;
wire n_12096;
wire n_12097;
wire n_12098;
wire n_12099;
wire n_12100;
wire n_12101;
wire n_12102;
wire n_12103;
wire n_12104;
wire n_12105;
wire n_12106;
wire n_12107;
wire n_12108;
wire n_12109;
wire n_12110;
wire n_12111;
wire n_12112;
wire n_12113;
wire n_12114;
wire n_12115;
wire n_12116;
wire n_12117;
wire n_12118;
wire n_12119;
wire n_12120;
wire n_12121;
wire n_12122;
wire n_12123;
wire n_12124;
wire n_12125;
wire n_12126;
wire n_12127;
wire n_12128;
wire n_12129;
wire n_12130;
wire n_12131;
wire n_12132;
wire n_12133;
wire n_12134;
wire n_12135;
wire n_12136;
wire n_12137;
wire n_12138;
wire n_12139;
wire n_12140;
wire n_12141;
wire n_12142;
wire n_12143;
wire n_12144;
wire n_12145;
wire n_12146;
wire n_12147;
wire n_12148;
wire n_12149;
wire n_12150;
wire n_12151;
wire n_12152;
wire n_12153;
wire n_12154;
wire n_12155;
wire n_12156;
wire n_12157;
wire n_12158;
wire n_12159;
wire n_12160;
wire n_12161;
wire n_12162;
wire n_12163;
wire n_12164;
wire n_12165;
wire n_12166;
wire n_12167;
wire n_12168;
wire n_12169;
wire n_12170;
wire n_12171;
wire n_12172;
wire n_12173;
wire n_12174;
wire n_12175;
wire n_12176;
wire n_12177;
wire n_12178;
wire n_12179;
wire n_12180;
wire n_12181;
wire n_12182;
wire n_12183;
wire n_12184;
wire n_12185;
wire n_12186;
wire n_12187;
wire n_12188;
wire n_12189;
wire n_12190;
wire n_12191;
wire n_12192;
wire n_12193;
wire n_12194;
wire n_12195;
wire n_12196;
wire n_12197;
wire n_12198;
wire n_12199;
wire n_12200;
wire n_12201;
wire n_12202;
wire n_12203;
wire n_12204;
wire n_12205;
wire n_12206;
wire n_12207;
wire n_12208;
wire n_12209;
wire n_12210;
wire n_12211;
wire n_12212;
wire n_12213;
wire n_12214;
wire n_12215;
wire n_12216;
wire n_12217;
wire n_12218;
wire n_12219;
wire n_12220;
wire n_12221;
wire n_12222;
wire n_12223;
wire n_12224;
wire n_12225;
wire n_12226;
wire n_12227;
wire n_12228;
wire n_12229;
wire n_12230;
wire n_12231;
wire n_12232;
wire n_12233;
wire n_12234;
wire n_12235;
wire n_12236;
wire n_12237;
wire n_12238;
wire n_12239;
wire n_12240;
wire n_12241;
wire n_12242;
wire n_12243;
wire n_12244;
wire n_12245;
wire n_12246;
wire n_12247;
wire n_12248;
wire n_12249;
wire n_12250;
wire n_12251;
wire n_12252;
wire n_12253;
wire n_12254;
wire n_12255;
wire n_12256;
wire n_12257;
wire n_12258;
wire n_12259;
wire n_12260;
wire n_12261;
wire n_12262;
wire n_12263;
wire n_12264;
wire n_12265;
wire n_12266;
wire n_12267;
wire n_12268;
wire n_12269;
wire n_12270;
wire n_12271;
wire n_12272;
wire n_12273;
wire n_12274;
wire n_12275;
wire n_12276;
wire n_12277;
wire n_12278;
wire n_12279;
wire n_12280;
wire n_12281;
wire n_12282;
wire n_12283;
wire n_12284;
wire n_12285;
wire n_12286;
wire n_12287;
wire n_12288;
wire n_12289;
wire n_12290;
wire n_12291;
wire n_12292;
wire n_12293;
wire n_12294;
wire n_12295;
wire n_12296;
wire n_12297;
wire n_12298;
wire n_12299;
wire n_12300;
wire n_12301;
wire n_12302;
wire n_12303;
wire n_12304;
wire n_12305;
wire n_12306;
wire n_12307;
wire n_12308;
wire n_12309;
wire n_12310;
wire n_12311;
wire n_12312;
wire n_12313;
wire n_12314;
wire n_12315;
wire n_12316;
wire n_12317;
wire n_12318;
wire n_12319;
wire n_12320;
wire n_12321;
wire n_12322;
wire n_12323;
wire n_12324;
wire n_12325;
wire n_12326;
wire n_12327;
wire n_12328;
wire n_12329;
wire n_12330;
wire n_12331;
wire n_12332;
wire n_12333;
wire n_12334;
wire n_12335;
wire n_12336;
wire n_12337;
wire n_12338;
wire n_12339;
wire n_12340;
wire n_12341;
wire n_12342;
wire n_12343;
wire n_12344;
wire n_12345;
wire n_12346;
wire n_12347;
wire n_12348;
wire n_12349;
wire n_12350;
wire n_12351;
wire n_12352;
wire n_12353;
wire n_12354;
wire n_12355;
wire n_12356;
wire n_12357;
wire n_12358;
wire n_12359;
wire n_12360;
wire n_12361;
wire n_12362;
wire n_12363;
wire n_12364;
wire n_12365;
wire n_12366;
wire n_12367;
wire n_12368;
wire n_12369;
wire n_12370;
wire n_12371;
wire n_12372;
wire n_12373;
wire n_12374;
wire n_12375;
wire n_12376;
wire n_12377;
wire n_12378;
wire n_12379;
wire n_12380;
wire n_12381;
wire n_12382;
wire n_12383;
wire n_12384;
wire n_12385;
wire n_12386;
wire n_12387;
wire n_12388;
wire n_12389;
wire n_12390;
wire n_12391;
wire n_12392;
wire n_12393;
wire n_12394;
wire n_12395;
wire n_12396;
wire n_12397;
wire n_12398;
wire n_12399;
wire n_12400;
wire n_12401;
wire n_12402;
wire n_12403;
wire n_12404;
wire n_12405;
wire n_12406;
wire n_12407;
wire n_12408;
wire n_12409;
wire n_12410;
wire n_12411;
wire n_12412;
wire n_12413;
wire n_12414;
wire n_12415;
wire n_12416;
wire n_12417;
wire n_12418;
wire n_12419;
wire n_12420;
wire n_12421;
wire n_12422;
wire n_12423;
wire n_12424;
wire n_12425;
wire n_12426;
wire n_12427;
wire n_12428;
wire n_12429;
wire n_12430;
wire n_12431;
wire n_12432;
wire n_12433;
wire n_12434;
wire n_12435;
wire n_12436;
wire n_12437;
wire n_12438;
wire n_12439;
wire n_12440;
wire n_12441;
wire n_12442;
wire n_12443;
wire n_12444;
wire n_12445;
wire n_12446;
wire n_12447;
wire n_12448;
wire n_12449;
wire n_12450;
wire n_12451;
wire n_12452;
wire n_12453;
wire n_12454;
wire n_12455;
wire n_12456;
wire n_12457;
wire n_12458;
wire n_12459;
wire n_12460;
wire n_12461;
wire n_12462;
wire n_12463;
wire n_12464;
wire n_12465;
wire n_12466;
wire n_12467;
wire n_12468;
wire n_12469;
wire n_12470;
wire n_12471;
wire n_12472;
wire n_12473;
wire n_12474;
wire n_12475;
wire n_12476;
wire n_12477;
wire n_12478;
wire n_12479;
wire n_12480;
wire n_12481;
wire n_12482;
wire n_12483;
wire n_12484;
wire n_12485;
wire n_12486;
wire n_12487;
wire n_12488;
wire n_12489;
wire n_12490;
wire n_12491;
wire n_12492;
wire n_12493;
wire n_12494;
wire n_12495;
wire n_12496;
wire n_12497;
wire n_12498;
wire n_12499;
wire n_12500;
wire n_12501;
wire n_12502;
wire n_12503;
wire n_12504;
wire n_12505;
wire n_12506;
wire n_12507;
wire n_12508;
wire n_12509;
wire n_12510;
wire n_12511;
wire n_12512;
wire n_12513;
wire n_12514;
wire n_12515;
wire n_12516;
wire n_12517;
wire n_12518;
wire n_12519;
wire n_12520;
wire n_12521;
wire n_12522;
wire n_12523;
wire n_12524;
wire n_12525;
wire n_12526;
wire n_12527;
wire n_12528;
wire n_12529;
wire n_12530;
wire n_12531;
wire n_12532;
wire n_12533;
wire n_12534;
wire n_12535;
wire n_12536;
wire n_12537;
wire n_12538;
wire n_12539;
wire n_12540;
wire n_12541;
wire n_12542;
wire n_12543;
wire n_12544;
wire n_12545;
wire n_12546;
wire n_12547;
wire n_12548;
wire n_12549;
wire n_12550;
wire n_12551;
wire n_12552;
wire n_12553;
wire n_12554;
wire n_12555;
wire n_12556;
wire n_12557;
wire n_12558;
wire n_12559;
wire n_12560;
wire n_12561;
wire n_12562;
wire n_12563;
wire n_12564;
wire n_12565;
wire n_12566;
wire n_12567;
wire n_12568;
wire n_12569;
wire n_12570;
wire n_12571;
wire n_12572;
wire n_12573;
wire n_12574;
wire n_12575;
wire n_12576;
wire n_12577;
wire n_12578;
wire n_12579;
wire n_12580;
wire n_12581;
wire n_12582;
wire n_12583;
wire n_12584;
wire n_12585;
wire n_12586;
wire n_12587;
wire n_12588;
wire n_12589;
wire n_12590;
wire n_12591;
wire n_12592;
wire n_12593;
wire n_12594;
wire n_12595;
wire n_12596;
wire n_12597;
wire n_12598;
wire n_12599;
wire n_12600;
wire n_12601;
wire n_12602;
wire n_12603;
wire n_12604;
wire n_12605;
wire n_12606;
wire n_12607;
wire n_12608;
wire n_12609;
wire n_12610;
wire n_12611;
wire n_12612;
wire n_12613;
wire n_12614;
wire n_12615;
wire n_12616;
wire n_12617;
wire n_12618;
wire n_12619;
wire n_12620;
wire n_12621;
wire n_12622;
wire n_12623;
wire n_12624;
wire n_12625;
wire n_12626;
wire n_12627;
wire n_12628;
wire n_12629;
wire n_12630;
wire n_12631;
wire n_12632;
wire n_12633;
wire n_12634;
wire n_12635;
wire n_12636;
wire n_12637;
wire n_12638;
wire n_12639;
wire n_12640;
wire n_12641;
wire n_12642;
wire n_12643;
wire n_12644;
wire n_12645;
wire n_12646;
wire n_12647;
wire n_12648;
wire n_12649;
wire n_12650;
wire n_12651;
wire n_12652;
wire n_12653;
wire n_12654;
wire n_12655;
wire n_12656;
wire n_12657;
wire n_12658;
wire n_12659;
wire n_12660;
wire n_12661;
wire n_12662;
wire n_12663;
wire n_12664;
wire n_12665;
wire n_12666;
wire n_12667;
wire n_12668;
wire n_12669;
wire n_12670;
wire n_12671;
wire n_12672;
wire n_12673;
wire n_12674;
wire n_12675;
wire n_12676;
wire n_12677;
wire n_12678;
wire n_12679;
wire n_12680;
wire n_12681;
wire n_12682;
wire n_12683;
wire n_12684;
wire n_12685;
wire n_12686;
wire n_12687;
wire n_12688;
wire n_12689;
wire n_12690;
wire n_12691;
wire n_12692;
wire n_12693;
wire n_12694;
wire n_12695;
wire n_12696;
wire n_12697;
wire n_12698;
wire n_12699;
wire n_12700;
wire n_12701;
wire n_12702;
wire n_12703;
wire n_12704;
wire n_12705;
wire n_12706;
wire n_12707;
wire n_12708;
wire n_12709;
wire n_12710;
wire n_12711;
wire n_12712;
wire n_12713;
wire n_12714;
wire n_12715;
wire n_12716;
wire n_12717;
wire n_12718;
wire n_12719;
wire n_12720;
wire n_12721;
wire n_12722;
wire n_12723;
wire n_12724;
wire n_12725;
wire n_12726;
wire n_12727;
wire n_12728;
wire n_12729;
wire n_12730;
wire n_12731;
wire n_12732;
wire n_12733;
wire n_12734;
wire n_12735;
wire n_12736;
wire n_12737;
wire n_12738;
wire n_12739;
wire n_12740;
wire n_12741;
wire n_12742;
wire n_12743;
wire n_12744;
wire n_12745;
wire n_12746;
wire n_12747;
wire n_12748;
wire n_12749;
wire n_12750;
wire n_12751;
wire n_12752;
wire n_12753;
wire n_12754;
wire n_12755;
wire n_12756;
wire n_12757;
wire n_12758;
wire n_12759;
wire n_12760;
wire n_12761;
wire n_12762;
wire n_12763;
wire n_12764;
wire n_12765;
wire n_12766;
wire n_12767;
wire n_12768;
wire n_12769;
wire n_12770;
wire n_12771;
wire n_12772;
wire n_12773;
wire n_12774;
wire n_12775;
wire n_12776;
wire n_12777;
wire n_12778;
wire n_12779;
wire n_12780;
wire n_12781;
wire n_12782;
wire n_12783;
wire n_12784;
wire n_12785;
wire n_12786;
wire n_12787;
wire n_12788;
wire n_12789;
wire n_12790;
wire n_12791;
wire n_12792;
wire n_12793;
wire n_12794;
wire n_12795;
wire n_12796;
wire n_12797;
wire n_12798;
wire n_12799;
wire n_12800;
wire n_12801;
wire n_12802;
wire n_12803;
wire n_12804;
wire n_12805;
wire n_12806;
wire n_12807;
wire n_12808;
wire n_12809;
wire n_12810;
wire n_12811;
wire n_12812;
wire n_12813;
wire n_12814;
wire n_12815;
wire n_12816;
wire n_12817;
wire n_12818;
wire n_12819;
wire n_12820;
wire n_12821;
wire n_12822;
wire n_12823;
wire n_12824;
wire n_12825;
wire n_12826;
wire n_12827;
wire n_12828;
wire n_12829;
wire n_12830;
wire n_12831;
wire n_12832;
wire n_12833;
wire n_12834;
wire n_12835;
wire n_12836;
wire n_12837;
wire n_12838;
wire n_12839;
wire n_12840;
wire n_12841;
wire n_12842;
wire n_12843;
wire n_12844;
wire n_12845;
wire n_12846;
wire n_12847;
wire n_12848;
wire n_12849;
wire n_12850;
wire n_12851;
wire n_12852;
wire n_12853;
wire n_12854;
wire n_12855;
wire n_12856;
wire n_12857;
wire n_12858;
wire n_12859;
wire n_12860;
wire n_12861;
wire n_12862;
wire n_12863;
wire n_12864;
wire n_12865;
wire n_12866;
wire n_12867;
wire n_12868;
wire n_12869;
wire n_12870;
wire n_12871;
wire n_12872;
wire n_12873;
wire n_12874;
wire n_12875;
wire n_12876;
wire n_12877;
wire n_12878;
wire n_12879;
wire n_12880;
wire n_12881;
wire n_12882;
wire n_12883;
wire n_12884;
wire n_12885;
wire n_12886;
wire n_12887;
wire n_12888;
wire n_12889;
wire n_12890;
wire n_12891;
wire n_12892;
wire n_12893;
wire n_12894;
wire n_12895;
wire n_12896;
wire n_12897;
wire n_12898;
wire n_12899;
wire n_12900;
wire n_12901;
wire n_12902;
wire n_12903;
wire n_12904;
wire n_12905;
wire n_12906;
wire n_12907;
wire n_12908;
wire n_12909;
wire n_12910;
wire n_12911;
wire n_12912;
wire n_12913;
wire n_12914;
wire n_12915;
wire n_12916;
wire n_12917;
wire n_12918;
wire n_12919;
wire n_12920;
wire n_12921;
wire n_12922;
wire n_12923;
wire n_12924;
wire n_12925;
wire n_12926;
wire n_12927;
wire n_12928;
wire n_12929;
wire n_12930;
wire n_12931;
wire n_12932;
wire n_12933;
wire n_12934;
wire n_12935;
wire n_12936;
wire n_12937;
wire n_12938;
wire n_12939;
wire n_12940;
wire n_12941;
wire n_12942;
wire n_12943;
wire n_12944;
wire n_12945;
wire n_12946;
wire n_12947;
wire n_12948;
wire n_12949;
wire n_12950;
wire n_12951;
wire n_12952;
wire n_12953;
wire n_12954;
wire n_12955;
wire n_12956;
wire n_12957;
wire n_12958;
wire n_12959;
wire n_12960;
wire n_12961;
wire n_12962;
wire n_12963;
wire n_12964;
wire n_12965;
wire n_12966;
wire n_12967;
wire n_12968;
wire n_12969;
wire n_12970;
wire n_12971;
wire n_12972;
wire n_12973;
wire n_12974;
wire n_12975;
wire n_12976;
wire n_12977;
wire n_12978;
wire n_12979;
wire n_12980;
wire n_12981;
wire n_12982;
wire n_12983;
wire n_12984;
wire n_12985;
wire n_12986;
wire n_12987;
wire n_12988;
wire n_12989;
wire n_12990;
wire n_12991;
wire n_12992;
wire n_12993;
wire n_12994;
wire n_12995;
wire n_12996;
wire n_12997;
wire n_12998;
wire n_12999;
wire n_13000;
wire n_13001;
wire n_13002;
wire n_13003;
wire n_13004;
wire n_13005;
wire n_13006;
wire n_13007;
wire n_13008;
wire n_13009;
wire n_13010;
wire n_13011;
wire n_13012;
wire n_13013;
wire n_13014;
wire n_13015;
wire n_13016;
wire n_13017;
wire n_13018;
wire n_13019;
wire n_13020;
wire n_13021;
wire n_13022;
wire n_13023;
wire n_13024;
wire n_13025;
wire n_13026;
wire n_13027;
wire n_13028;
wire n_13029;
wire n_13030;
wire n_13031;
wire n_13032;
wire n_13033;
wire n_13034;
wire n_13035;
wire n_13036;
wire n_13037;
wire n_13038;
wire n_13039;
wire n_13040;
wire n_13041;
wire n_13042;
wire n_13043;
wire n_13044;
wire n_13045;
wire n_13046;
wire n_13047;
wire n_13048;
wire n_13049;
wire n_13050;
wire n_13051;
wire n_13052;
wire n_13053;
wire n_13054;
wire n_13055;
wire n_13056;
wire n_13057;
wire n_13058;
wire n_13059;
wire n_13060;
wire n_13061;
wire n_13062;
wire n_13063;
wire n_13064;
wire n_13065;
wire n_13066;
wire n_13067;
wire n_13068;
wire n_13069;
wire n_13070;
wire n_13071;
wire n_13072;
wire n_13073;
wire n_13074;
wire n_13075;
wire n_13076;
wire n_13077;
wire n_13078;
wire n_13079;
wire n_13080;
wire n_13081;
wire n_13082;
wire n_13083;
wire n_13084;
wire n_13085;
wire n_13086;
wire n_13087;
wire n_13088;
wire n_13089;
wire n_13090;
wire n_13091;
wire n_13092;
wire n_13093;
wire n_13094;
wire n_13095;
wire n_13096;
wire n_13097;
wire n_13098;
wire n_13099;
wire n_13100;
wire n_13101;
wire n_13102;
wire n_13103;
wire n_13104;
wire n_13105;
wire n_13106;
wire n_13107;
wire n_13108;
wire n_13109;
wire n_13110;
wire n_13111;
wire n_13112;
wire n_13113;
wire n_13114;
wire n_13115;
wire n_13116;
wire n_13117;
wire n_13118;
wire n_13119;
wire n_13120;
wire n_13121;
wire n_13122;
wire n_13123;
wire n_13124;
wire n_13125;
wire n_13126;
wire n_13127;
wire n_13128;
wire n_13129;
wire n_13130;
wire n_13131;
wire n_13132;
wire n_13133;
wire n_13134;
wire n_13135;
wire n_13136;
wire n_13137;
wire n_13138;
wire n_13139;
wire n_13140;
wire n_13141;
wire n_13142;
wire n_13143;
wire n_13144;
wire n_13145;
wire n_13146;
wire n_13147;
wire n_13148;
wire n_13149;
wire n_13150;
wire n_13151;
wire n_13152;
wire n_13153;
wire n_13154;
wire n_13155;
wire n_13156;
wire n_13157;
wire n_13158;
wire n_13159;
wire n_13160;
wire n_13161;
wire n_13162;
wire n_13163;
wire n_13164;
wire n_13165;
wire n_13166;
wire n_13167;
wire n_13168;
wire n_13169;
wire n_13170;
wire n_13171;
wire n_13172;
wire n_13173;
wire n_13174;
wire n_13175;
wire n_13176;
wire n_13177;
wire n_13178;
wire n_13179;
wire n_13180;
wire n_13181;
wire n_13182;
wire n_13183;
wire n_13184;
wire n_13185;
wire n_13186;
wire n_13187;
wire n_13188;
wire n_13189;
wire n_13190;
wire n_13191;
wire n_13192;
wire n_13193;
wire n_13194;
wire n_13195;
wire n_13196;
wire n_13197;
wire n_13198;
wire n_13199;
wire n_13200;
wire n_13201;
wire n_13202;
wire n_13203;
wire n_13204;
wire n_13205;
wire n_13206;
wire n_13207;
wire n_13208;
wire n_13209;
wire n_13210;
wire n_13211;
wire n_13212;
wire n_13213;
wire n_13214;
wire n_13215;
wire n_13216;
wire n_13217;
wire n_13218;
wire n_13219;
wire n_13220;
wire n_13221;
wire n_13222;
wire n_13223;
wire n_13224;
wire n_13225;
wire n_13226;
wire n_13227;
wire n_13228;
wire n_13229;
wire n_13230;
wire n_13231;
wire n_13232;
wire n_13233;
wire n_13234;
wire n_13235;
wire n_13236;
wire n_13237;
wire n_13238;
wire n_13239;
wire n_13240;
wire n_13241;
wire n_13242;
wire n_13243;
wire n_13244;
wire n_13245;
wire n_13246;
wire n_13247;
wire n_13248;
wire n_13249;
wire n_13250;
wire n_13251;
wire n_13252;
wire n_13253;
wire n_13254;
wire n_13255;
wire n_13256;
wire n_13257;
wire n_13258;
wire n_13259;
wire n_13260;
wire n_13261;
wire n_13262;
wire n_13263;
wire n_13264;
wire n_13265;
wire n_13266;
wire n_13267;
wire n_13268;
wire n_13269;
wire n_13270;
wire n_13271;
wire n_13272;
wire n_13273;
wire n_13274;
wire n_13275;
wire n_13276;
wire n_13277;
wire n_13278;
wire n_13279;
wire n_13280;
wire n_13281;
wire n_13282;
wire n_13283;
wire n_13284;
wire n_13285;
wire n_13286;
wire n_13287;
wire n_13288;
wire n_13289;
wire n_13290;
wire n_13291;
wire n_13292;
wire n_13293;
wire n_13294;
wire n_13295;
wire n_13296;
wire n_13297;
wire n_13298;
wire n_13299;
wire n_13300;
wire n_13301;
wire n_13302;
wire n_13303;
wire n_13304;
wire n_13305;
wire n_13306;
wire n_13307;
wire n_13308;
wire n_13309;
wire n_13310;
wire n_13311;
wire n_13312;
wire n_13313;
wire n_13314;
wire n_13315;
wire n_13316;
wire n_13317;
wire n_13318;
wire n_13319;
wire n_13320;
wire n_13321;
wire n_13322;
wire n_13323;
wire n_13324;
wire n_13325;
wire n_13326;
wire n_13327;
wire n_13328;
wire n_13329;
wire n_13330;
wire n_13331;
wire n_13332;
wire n_13333;
wire n_13334;
wire n_13335;
wire n_13336;
wire n_13337;
wire n_13338;
wire n_13339;
wire n_13340;
wire n_13341;
wire n_13342;
wire n_13343;
wire n_13344;
wire n_13345;
wire n_13346;
wire n_13347;
wire n_13348;
wire n_13349;
wire n_13350;
wire n_13351;
wire n_13352;
wire n_13353;
wire n_13354;
wire n_13355;
wire n_13356;
wire n_13357;
wire n_13358;
wire n_13359;
wire n_13360;
wire n_13361;
wire n_13362;
wire n_13363;
wire n_13364;
wire n_13365;
wire n_13366;
wire n_13367;
wire n_13368;
wire n_13369;
wire n_13370;
wire n_13371;
wire n_13372;
wire n_13373;
wire n_13374;
wire n_13375;
wire n_13376;
wire n_13377;
wire n_13378;
wire n_13379;
wire n_13380;
wire n_13381;
wire n_13382;
wire n_13383;
wire n_13384;
wire n_13385;
wire n_13386;
wire n_13387;
wire n_13388;
wire n_13389;
wire n_13390;
wire n_13391;
wire n_13392;
wire n_13393;
wire n_13394;
wire n_13395;
wire n_13396;
wire n_13397;
wire n_13398;
wire n_13399;
wire n_13400;
wire n_13401;
wire n_13402;
wire n_13403;
wire n_13404;
wire n_13405;
wire n_13406;
wire n_13407;
wire n_13408;
wire n_13409;
wire n_13410;
wire n_13411;
wire n_13412;
wire n_13413;
wire n_13414;
wire n_13415;
wire n_13416;
wire n_13417;
wire n_13418;
wire n_13419;
wire n_13420;
wire n_13421;
wire n_13422;
wire n_13423;
wire n_13424;
wire n_13425;
wire n_13426;
wire n_13427;
wire n_13428;
wire n_13429;
wire n_13430;
wire n_13431;
wire n_13432;
wire n_13433;
wire n_13434;
wire n_13435;
wire n_13436;
wire n_13437;
wire n_13438;
wire n_13439;
wire n_13440;
wire n_13441;
wire n_13442;
wire n_13443;
wire n_13444;
wire n_13445;
wire n_13446;
wire n_13447;
wire n_13448;
wire n_13449;
wire n_13450;
wire n_13451;
wire n_13452;
wire n_13453;
wire n_13454;
wire n_13455;
wire n_13456;
wire n_13457;
wire n_13458;
wire n_13459;
wire n_13460;
wire n_13461;
wire n_13462;
wire n_13463;
wire n_13464;
wire n_13465;
wire n_13466;
wire n_13467;
wire n_13468;
wire n_13469;
wire n_13470;
wire n_13471;
wire n_13472;
wire n_13473;
wire n_13474;
wire n_13475;
wire n_13476;
wire n_13477;
wire n_13478;
wire n_13479;
wire n_13480;
wire n_13481;
wire n_13482;
wire n_13483;
wire n_13484;
wire n_13485;
wire n_13486;
wire n_13487;
wire n_13488;
wire n_13489;
wire n_13490;
wire n_13491;
wire n_13492;
wire n_13493;
wire n_13494;
wire n_13495;
wire n_13496;
wire n_13497;
wire n_13498;
wire n_13499;
wire n_13500;
wire n_13501;
wire n_13502;
wire n_13503;
wire n_13504;
wire n_13505;
wire n_13506;
wire n_13507;
wire n_13508;
wire n_13509;
wire n_13510;
wire n_13511;
wire n_13512;
wire n_13513;
wire n_13514;
wire n_13515;
wire n_13516;
wire n_13517;
wire n_13518;
wire n_13519;
wire n_13520;
wire n_13521;
wire n_13522;
wire n_13523;
wire n_13524;
wire n_13525;
wire n_13526;
wire n_13527;
wire n_13528;
wire n_13529;
wire n_13530;
wire n_13531;
wire n_13532;
wire n_13533;
wire n_13534;
wire n_13535;
wire n_13536;
wire n_13537;
wire n_13538;
wire n_13539;
wire n_13540;
wire n_13541;
wire n_13542;
wire n_13543;
wire n_13544;
wire n_13545;
wire n_13546;
wire n_13547;
wire n_13548;
wire n_13549;
wire n_13550;
wire n_13551;
wire n_13552;
wire n_13553;
wire n_13554;
wire n_13555;
wire n_13556;
wire n_13557;
wire n_13558;
wire n_13559;
wire n_13560;
wire n_13561;
wire n_13562;
wire n_13563;
wire n_13564;
wire n_13565;
wire n_13566;
wire n_13567;
wire n_13568;
wire n_13569;
wire n_13570;
wire n_13571;
wire n_13572;
wire n_13573;
wire n_13574;
wire n_13575;
wire n_13576;
wire n_13577;
wire n_13578;
wire n_13579;
wire n_13580;
wire n_13581;
wire n_13582;
wire n_13583;
wire n_13584;
wire n_13585;
wire n_13586;
wire n_13587;
wire n_13588;
wire n_13589;
wire n_13590;
wire n_13591;
wire n_13592;
wire n_13593;
wire n_13594;
wire n_13595;
wire n_13596;
wire n_13597;
wire n_13598;
wire n_13599;
wire n_13600;
wire n_13601;
wire n_13602;
wire n_13603;
wire n_13604;
wire n_13605;
wire n_13606;
wire n_13607;
wire n_13608;
wire n_13609;
wire n_13610;
wire n_13611;
wire n_13612;
wire n_13613;
wire n_13614;
wire n_13615;
wire n_13616;
wire n_13617;
wire n_13618;
wire n_13619;
wire n_13620;
wire n_13621;
wire n_13622;
wire n_13623;
wire n_13624;
wire n_13625;
wire n_13626;
wire n_13627;
wire n_13628;
wire n_13629;
wire n_13630;
wire n_13631;
wire n_13632;
wire n_13633;
wire n_13634;
wire n_13635;
wire n_13636;
wire n_13637;
wire n_13638;
wire n_13639;
wire n_13640;
wire n_13641;
wire n_13642;
wire n_13643;
wire n_13644;
wire n_13645;
wire n_13646;
wire n_13647;
wire n_13648;
wire n_13649;
wire n_13650;
wire n_13651;
wire n_13652;
wire n_13653;
wire n_13654;
wire n_13655;
wire n_13656;
wire n_13657;
wire n_13658;
wire n_13659;
wire n_13660;
wire n_13661;
wire n_13662;
wire n_13663;
wire n_13664;
wire n_13665;
wire n_13666;
wire n_13667;
wire n_13668;
wire n_13669;
wire n_13670;
wire n_13671;
wire n_13672;
wire n_13673;
wire n_13674;
wire n_13675;
wire n_13676;
wire n_13677;
wire n_13678;
wire n_13679;
wire n_13680;
wire n_13681;
wire n_13682;
wire n_13683;
wire n_13684;
wire n_13685;
wire n_13686;
wire n_13687;
wire n_13688;
wire n_13689;
wire n_13690;
wire n_13691;
wire n_13692;
wire n_13693;
wire n_13694;
wire n_13695;
wire n_13696;
wire n_13697;
wire n_13698;
wire n_13699;
wire n_13700;
wire n_13701;
wire n_13702;
wire n_13703;
wire n_13704;
wire n_13705;
wire n_13706;
wire n_13707;
wire n_13708;
wire n_13709;
wire n_13710;
wire n_13711;
wire n_13712;
wire n_13713;
wire n_13714;
wire n_13715;
wire n_13716;
wire n_13717;
wire n_13718;
wire n_13719;
wire n_13720;
wire n_13721;
wire n_13722;
wire n_13723;
wire n_13724;
wire n_13725;
wire n_13726;
wire n_13727;
wire n_13728;
wire n_13729;
wire n_13730;
wire n_13731;
wire n_13732;
wire n_13733;
wire n_13734;
wire n_13735;
wire n_13736;
wire n_13737;
wire n_13738;
wire n_13739;
wire n_13740;
wire n_13741;
wire n_13742;
wire n_13743;
wire n_13744;
wire n_13745;
wire n_13746;
wire n_13747;
wire n_13748;
wire n_13749;
wire n_13750;
wire n_13751;
wire n_13752;
wire n_13753;
wire n_13754;
wire n_13755;
wire n_13756;
wire n_13757;
wire n_13758;
wire n_13759;
wire n_13760;
wire n_13761;
wire n_13762;
wire n_13763;
wire n_13764;
wire n_13765;
wire n_13766;
wire n_13767;
wire n_13768;
wire n_13769;
wire n_13770;
wire n_13771;
wire n_13772;
wire n_13773;
wire n_13774;
wire n_13775;
wire n_13776;
wire n_13777;
wire n_13778;
wire n_13779;
wire n_13780;
wire n_13781;
wire n_13782;
wire n_13783;
wire n_13784;
wire n_13785;
wire n_13786;
wire n_13787;
wire n_13788;
wire n_13789;
wire n_13790;
wire n_13791;
wire n_13792;
wire n_13793;
wire n_13794;
wire n_13795;
wire n_13796;
wire n_13797;
wire n_13798;
wire n_13799;
wire n_13800;
wire n_13801;
wire n_13802;
wire n_13803;
wire n_13804;
wire n_13805;
wire n_13806;
wire n_13807;
wire n_13808;
wire n_13809;
wire n_13810;
wire n_13811;
wire n_13812;
wire n_13813;
wire n_13814;
wire n_13815;
wire n_13816;
wire n_13817;
wire n_13818;
wire n_13819;
wire n_13820;
wire n_13821;
wire n_13822;
wire n_13823;
wire n_13824;
wire n_13825;
wire n_13826;
wire n_13827;
wire n_13828;
wire n_13829;
wire n_13830;
wire n_13831;
wire n_13832;
wire n_13833;
wire n_13834;
wire n_13835;
wire n_13836;
wire n_13837;
wire n_13838;
wire n_13839;
wire n_13840;
wire n_13841;
wire n_13842;
wire n_13843;
wire n_13844;
wire n_13845;
wire n_13846;
wire n_13847;
wire n_13848;
wire n_13849;
wire n_13850;
wire n_13851;
wire n_13852;
wire n_13853;
wire n_13854;
wire n_13855;
wire n_13856;
wire n_13857;
wire n_13858;
wire n_13859;
wire n_13860;
wire n_13861;
wire n_13862;
wire n_13863;
wire n_13864;
wire n_13865;
wire n_13866;
wire n_13867;
wire n_13868;
wire n_13869;
wire n_13870;
wire n_13871;
wire n_13872;
wire n_13873;
wire n_13874;
wire n_13875;
wire n_13876;
wire n_13877;
wire n_13878;
wire n_13879;
wire n_13880;
wire n_13881;
wire n_13882;
wire n_13883;
wire n_13884;
wire n_13885;
wire n_13886;
wire n_13887;
wire n_13888;
wire n_13889;
wire n_13890;
wire n_13891;
wire n_13892;
wire n_13893;
wire n_13894;
wire n_13895;
wire n_13896;
wire n_13897;
wire n_13898;
wire n_13899;
wire n_13900;
wire n_13901;
wire n_13902;
wire n_13903;
wire n_13904;
wire n_13905;
wire n_13906;
wire n_13907;
wire n_13908;
wire n_13909;
wire n_13910;
wire n_13911;
wire n_13912;
wire n_13913;
wire n_13914;
wire n_13915;
wire n_13916;
wire n_13917;
wire n_13918;
wire n_13919;
wire n_13920;
wire n_13921;
wire n_13922;
wire n_13923;
wire n_13924;
wire n_13925;
wire n_13926;
wire n_13927;
wire n_13928;
wire n_13929;
wire n_13930;
wire n_13931;
wire n_13932;
wire n_13933;
wire n_13934;
wire n_13935;
wire n_13936;
wire n_13937;
wire n_13938;
wire n_13939;
wire n_13940;
wire n_13941;
wire n_13942;
wire n_13943;
wire n_13944;
wire n_13945;
wire n_13946;
wire n_13947;
wire n_13948;
wire n_13949;
wire n_13950;
wire n_13951;
wire n_13952;
wire n_13953;
wire n_13954;
wire n_13955;
wire n_13956;
wire n_13957;
wire n_13958;
wire n_13959;
wire n_13960;
wire n_13961;
wire n_13962;
wire n_13963;
wire n_13964;
wire n_13965;
wire n_13966;
wire n_13967;
wire n_13968;
wire n_13969;
wire n_13970;
wire n_13971;
wire n_13972;
wire n_13973;
wire n_13974;
wire n_13975;
wire n_13976;
wire n_13977;
wire n_13978;
wire n_13979;
wire n_13980;
wire n_13981;
wire n_13982;
wire n_13983;
wire n_13984;
wire n_13985;
wire n_13986;
wire n_13987;
wire n_13988;
wire n_13989;
wire n_13990;
wire n_13991;
wire n_13992;
wire n_13993;
wire n_13994;
wire n_13995;
wire n_13996;
wire n_13997;
wire n_13998;
wire n_13999;
wire n_14000;
wire n_14001;
wire n_14002;
wire n_14003;
wire n_14004;
wire n_14005;
wire n_14006;
wire n_14007;
wire n_14008;
wire n_14009;
wire n_14010;
wire n_14011;
wire n_14012;
wire n_14013;
wire n_14014;
wire n_14015;
wire n_14016;
wire n_14017;
wire n_14018;
wire n_14019;
wire n_14020;
wire n_14021;
wire n_14022;
wire n_14023;
wire n_14024;
wire n_14025;
wire n_14026;
wire n_14027;
wire n_14028;
wire n_14029;
wire n_14030;
wire n_14031;
wire n_14032;
wire n_14033;
wire n_14034;
wire n_14035;
wire n_14036;
wire n_14037;
wire n_14038;
wire n_14039;
wire n_14040;
wire n_14041;
wire n_14042;
wire n_14043;
wire n_14044;
wire n_14045;
wire n_14046;
wire n_14047;
wire n_14048;
wire n_14049;
wire n_14050;
wire n_14051;
wire n_14052;
wire n_14053;
wire n_14054;
wire n_14055;
wire n_14056;
wire n_14057;
wire n_14058;
wire n_14059;
wire n_14060;
wire n_14061;
wire n_14062;
wire n_14063;
wire n_14064;
wire n_14065;
wire n_14066;
wire n_14067;
wire n_14068;
wire n_14069;
wire n_14070;
wire n_14071;
wire n_14072;
wire n_14073;
wire n_14074;
wire n_14075;
wire n_14076;
wire n_14077;
wire n_14078;
wire n_14079;
wire n_14080;
wire n_14081;
wire n_14082;
wire n_14083;
wire n_14084;
wire n_14085;
wire n_14086;
wire n_14087;
wire n_14088;
wire n_14089;
wire n_14090;
wire n_14091;
wire n_14092;
wire n_14093;
wire n_14094;
wire n_14095;
wire n_14096;
wire n_14097;
wire n_14098;
wire n_14099;
wire n_14100;
wire n_14101;
wire n_14102;
wire n_14103;
wire n_14104;
wire n_14105;
wire n_14106;
wire n_14107;
wire n_14108;
wire n_14109;
wire n_14110;
wire n_14111;
wire n_14112;
wire n_14113;
wire n_14114;
wire n_14115;
wire n_14116;
wire n_14117;
wire n_14118;
wire n_14119;
wire n_14120;
wire n_14121;
wire n_14122;
wire n_14123;
wire n_14124;
wire n_14125;
wire n_14126;
wire n_14127;
wire n_14128;
wire n_14129;
wire n_14130;
wire n_14131;
wire n_14132;
wire n_14133;
wire n_14134;
wire n_14135;
wire n_14136;
wire n_14137;
wire n_14138;
wire n_14139;
wire n_14140;
wire n_14141;
wire n_14142;
wire n_14143;
wire n_14144;
wire n_14145;
wire n_14146;
wire n_14147;
wire n_14148;
wire n_14149;
wire n_14150;
wire n_14151;
wire n_14152;
wire n_14153;
wire n_14154;
wire n_14155;
wire n_14156;
wire n_14157;
wire n_14158;
wire n_14159;
wire n_14160;
wire n_14161;
wire n_14162;
wire n_14163;
wire n_14164;
wire n_14165;
wire n_14166;
wire n_14167;
wire n_14168;
wire n_14169;
wire n_14170;
wire n_14171;
wire n_14172;
wire n_14173;
wire n_14174;
wire n_14175;
wire n_14176;
wire n_14177;
wire n_14178;
wire n_14179;
wire n_14180;
wire n_14181;
wire n_14182;
wire n_14183;
wire n_14184;
wire n_14185;
wire n_14186;
wire n_14187;
wire n_14188;
wire n_14189;
wire n_14190;
wire n_14191;
wire n_14192;
wire n_14193;
wire n_14194;
wire n_14195;
wire n_14196;
wire n_14197;
wire n_14198;
wire n_14199;
wire n_14200;
wire n_14201;
wire n_14202;
wire n_14203;
wire n_14204;
wire n_14205;
wire n_14206;
wire n_14207;
wire n_14208;
wire n_14209;
wire n_14210;
wire n_14211;
wire n_14212;
wire n_14213;
wire n_14214;
wire n_14215;
wire n_14216;
wire n_14217;
wire n_14218;
wire n_14219;
wire n_14220;
wire n_14221;
wire n_14222;
wire n_14223;
wire n_14224;
wire n_14225;
wire n_14226;
wire n_14227;
wire n_14228;
wire n_14229;
wire n_14230;
wire n_14231;
wire n_14232;
wire n_14233;
wire n_14234;
wire n_14235;
wire n_14236;
wire n_14237;
wire n_14238;
wire n_14239;
wire n_14240;
wire n_14241;
wire n_14242;
wire n_14243;
wire n_14244;
wire n_14245;
wire n_14246;
wire n_14247;
wire n_14248;
wire n_14249;
wire n_14250;
wire n_14251;
wire n_14252;
wire n_14253;
wire n_14254;
wire n_14255;
wire n_14256;
wire n_14257;
wire n_14258;
wire n_14259;
wire n_14260;
wire n_14261;
wire n_14262;
wire n_14263;
wire n_14264;
wire n_14265;
wire n_14266;
wire n_14267;
wire n_14268;
wire n_14269;
wire n_14270;
wire n_14271;
wire n_14272;
wire n_14273;
wire n_14274;
wire n_14275;
wire n_14276;
wire n_14277;
wire n_14278;
wire n_14279;
wire n_14280;
wire n_14281;
wire n_14282;
wire n_14283;
wire n_14284;
wire n_14285;
wire n_14286;
wire n_14287;
wire n_14288;
wire n_14289;
wire n_14290;
wire n_14291;
wire n_14292;
wire n_14293;
wire n_14294;
wire n_14295;
wire n_14296;
wire n_14297;
wire n_14298;
wire n_14299;
wire n_14300;
wire n_14301;
wire n_14302;
wire n_14303;
wire n_14304;
wire n_14305;
wire n_14306;
wire n_14307;
wire n_14308;
wire n_14309;
wire n_14310;
wire n_14311;
wire n_14312;
wire n_14313;
wire n_14314;
wire n_14315;
wire n_14316;
wire n_14317;
wire n_14318;
wire n_14319;
wire n_14320;
wire n_14321;
wire n_14322;
wire n_14323;
wire n_14324;
wire n_14325;
wire n_14326;
wire n_14327;
wire n_14328;
wire n_14329;
wire n_14330;
wire n_14331;
wire n_14332;
wire n_14333;
wire n_14334;
wire n_14335;
wire n_14336;
wire n_14337;
wire n_14338;
wire n_14339;
wire n_14340;
wire n_14341;
wire n_14342;
wire n_14343;
wire n_14344;
wire n_14345;
wire n_14346;
wire n_14347;
wire n_14348;
wire n_14349;
wire n_14350;
wire n_14351;
wire n_14352;
wire n_14353;
wire n_14354;
wire n_14355;
wire n_14356;
wire n_14357;
wire n_14358;
wire n_14359;
wire n_14360;
wire n_14361;
wire n_14362;
wire n_14363;
wire n_14364;
wire n_14365;
wire n_14366;
wire n_14367;
wire n_14368;
wire n_14369;
wire n_14370;
wire n_14371;
wire n_14372;
wire n_14373;
wire n_14374;
wire n_14375;
wire n_14376;
wire n_14377;
wire n_14378;
wire n_14379;
wire n_14380;
wire n_14381;
wire n_14382;
wire n_14383;
wire n_14384;
wire n_14385;
wire n_14386;
wire n_14387;
wire n_14388;
wire n_14389;
wire n_14390;
wire n_14391;
wire n_14392;
wire n_14393;
wire n_14394;
wire n_14395;
wire n_14396;
wire n_14397;
wire n_14398;
wire n_14399;
wire n_14400;
wire n_14401;
wire n_14402;
wire n_14403;
wire n_14404;
wire n_14405;
wire n_14406;
wire n_14407;
wire n_14408;
wire n_14409;
wire n_14410;
wire n_14411;
wire n_14412;
wire n_14413;
wire n_14414;
wire n_14415;
wire n_14416;
wire n_14417;
wire n_14418;
wire n_14419;
wire n_14420;
wire n_14421;
wire n_14422;
wire n_14423;
wire n_14424;
wire n_14425;
wire n_14426;
wire n_14427;
wire n_14428;
wire n_14429;
wire n_14430;
wire n_14431;
wire n_14432;
wire n_14433;
wire n_14434;
wire n_14435;
wire n_14436;
wire n_14437;
wire n_14438;
wire n_14439;
wire n_14440;
wire n_14441;
wire n_14442;
wire n_14443;
wire n_14444;
wire n_14445;
wire n_14446;
wire n_14447;
wire n_14448;
wire n_14449;
wire n_14450;
wire n_14451;
wire n_14452;
wire n_14453;
wire n_14454;
wire n_14455;
wire n_14456;
wire n_14457;
wire n_14458;
wire n_14459;
wire n_14460;
wire n_14461;
wire n_14462;
wire n_14463;
wire n_14464;
wire n_14465;
wire n_14466;
wire n_14467;
wire n_14468;
wire n_14469;
wire n_14470;
wire n_14471;
wire n_14472;
wire n_14473;
wire n_14474;
wire n_14475;
wire n_14476;
wire n_14477;
wire n_14478;
wire n_14479;
wire n_14480;
wire n_14481;
wire n_14482;
wire n_14483;
wire n_14484;
wire n_14485;
wire n_14486;
wire n_14487;
wire n_14488;
wire n_14489;
wire n_14490;
wire n_14491;
wire n_14492;
wire n_14493;
wire n_14494;
wire n_14495;
wire n_14496;
wire n_14497;
wire n_14498;
wire n_14499;
wire n_14500;
wire n_14501;
wire n_14502;
wire n_14503;
wire n_14504;
wire n_14505;
wire n_14506;
wire n_14507;
wire n_14508;
wire n_14509;
wire n_14510;
wire n_14511;
wire n_14512;
wire n_14513;
wire n_14514;
wire n_14515;
wire n_14516;
wire n_14517;
wire n_14518;
wire n_14519;
wire n_14520;
wire n_14521;
wire n_14522;
wire n_14523;
wire n_14524;
wire n_14525;
wire n_14526;
wire n_14527;
wire n_14528;
wire n_14529;
wire n_14530;
wire n_14531;
wire n_14532;
wire n_14533;
wire n_14534;
wire n_14535;
wire n_14536;
wire n_14537;
wire n_14538;
wire n_14539;
wire n_14540;
wire n_14541;
wire n_14542;
wire n_14543;
wire n_14544;
wire n_14545;
wire n_14546;
wire n_14547;
wire n_14548;
wire n_14549;
wire n_14550;
wire n_14551;
wire n_14552;
wire n_14553;
wire n_14554;
wire n_14555;
wire n_14556;
wire n_14557;
wire n_14558;
wire n_14559;
wire n_14560;
wire n_14561;
wire n_14562;
wire n_14563;
wire n_14564;
wire n_14565;
wire n_14566;
wire n_14567;
wire n_14568;
wire n_14569;
wire n_14570;
wire n_14571;
wire n_14572;
wire n_14573;
wire n_14574;
wire n_14575;
wire n_14576;
wire n_14577;
wire n_14578;
wire n_14579;
wire n_14580;
wire n_14581;
wire n_14582;
wire n_14583;
wire n_14584;
wire n_14585;
wire n_14586;
wire n_14587;
wire n_14588;
wire n_14589;
wire n_14590;
wire n_14591;
wire n_14592;
wire n_14593;
wire n_14594;
wire n_14595;
wire n_14596;
wire n_14597;
wire n_14598;
wire n_14599;
wire n_14600;
wire n_14601;
wire n_14602;
wire n_14603;
wire n_14604;
wire n_14605;
wire n_14606;
wire n_14607;
wire n_14608;
wire n_14609;
wire n_14610;
wire n_14611;
wire n_14612;
wire n_14613;
wire n_14614;
wire n_14615;
wire n_14616;
wire n_14617;
wire n_14618;
wire n_14619;
wire n_14620;
wire n_14621;
wire n_14622;
wire n_14623;
wire n_14624;
wire n_14625;
wire n_14626;
wire n_14627;
wire n_14628;
wire n_14629;
wire n_14630;
wire n_14631;
wire n_14632;
wire n_14633;
wire n_14634;
wire n_14635;
wire n_14636;
wire n_14637;
wire n_14638;
wire n_14639;
wire n_14640;
wire n_14641;
wire n_14642;
wire n_14643;
wire n_14644;
wire n_14645;
wire n_14646;
wire n_14647;
wire n_14648;
wire n_14649;
wire n_14650;
wire n_14651;
wire n_14652;
wire n_14653;
wire n_14654;
wire n_14655;
wire n_14656;
wire n_14657;
wire n_14658;
wire n_14659;
wire n_14660;
wire n_14661;
wire n_14662;
wire n_14663;
wire n_14664;
wire n_14665;
wire n_14666;
wire n_14667;
wire n_14668;
wire n_14669;
wire n_14670;
wire n_14671;
wire n_14672;
wire n_14673;
wire n_14674;
wire n_14675;
wire n_14676;
wire n_14677;
wire n_14678;
wire n_14679;
wire n_14680;
wire n_14681;
wire n_14682;
wire n_14683;
wire n_14684;
wire n_14685;
wire n_14686;
wire n_14687;
wire n_14688;
wire n_14689;
wire n_14690;
wire n_14691;
wire n_14692;
wire n_14693;
wire n_14694;
wire n_14695;
wire n_14696;
wire n_14697;
wire n_14698;
wire n_14699;
wire n_14700;
wire n_14701;
wire n_14702;
wire n_14703;
wire n_14704;
wire n_14705;
wire n_14706;
wire n_14707;
wire n_14708;
wire n_14709;
wire n_14710;
wire n_14711;
wire n_14712;
wire n_14713;
wire n_14714;
wire n_14715;
wire n_14716;
wire n_14717;
wire n_14718;
wire n_14719;
wire n_14720;
wire n_14721;
wire n_14722;
wire n_14723;
wire n_14724;
wire n_14725;
wire n_14726;
wire n_14727;
wire n_14728;
wire n_14729;
wire n_14730;
wire n_14731;
wire n_14732;
wire n_14733;
wire n_14734;
wire n_14735;
wire n_14736;
wire n_14737;
wire n_14738;
wire n_14739;
wire n_14740;
wire n_14741;
wire n_14742;
wire n_14743;
wire n_14744;
wire n_14745;
wire n_14746;
wire n_14747;
wire n_14748;
wire n_14749;
wire n_14750;
wire n_14751;
wire n_14752;
wire n_14753;
wire n_14754;
wire n_14755;
wire n_14756;
wire n_14757;
wire n_14758;
wire n_14759;
wire n_14760;
wire n_14761;
wire n_14762;
wire n_14763;
wire n_14764;
wire n_14765;
wire n_14766;
wire n_14767;
wire n_14768;
wire n_14769;
wire n_14770;
wire n_14771;
wire n_14772;
wire n_14773;
wire n_14774;
wire n_14775;
wire n_14776;
wire n_14777;
wire n_14778;
wire n_14779;
wire n_14780;
wire n_14781;
wire n_14782;
wire n_14783;
wire n_14784;
wire n_14785;
wire n_14786;
wire n_14787;
wire n_14788;
wire n_14789;
wire n_14790;
wire n_14791;
wire n_14792;
wire n_14793;
wire n_14794;
wire n_14795;
wire n_14796;
wire n_14797;
wire n_14798;
wire n_14799;
wire n_14800;
wire n_14801;
wire n_14802;
wire n_14803;
wire n_14804;
wire n_14805;
wire n_14806;
wire n_14807;
wire n_14808;
wire n_14809;
wire n_14810;
wire n_14811;
wire n_14812;
wire n_14813;
wire n_14814;
wire n_14815;
wire n_14816;
wire n_14817;
wire n_14818;
wire n_14819;
wire n_14820;
wire n_14821;
wire n_14822;
wire n_14823;
wire n_14824;
wire n_14825;
wire n_14826;
wire n_14827;
wire n_14828;
wire n_14829;
wire n_14830;
wire n_14831;
wire n_14832;
wire n_14833;
wire n_14834;
wire n_14835;
wire n_14836;
wire n_14837;
wire n_14838;
wire n_14839;
wire n_14840;
wire n_14841;
wire n_14842;
wire n_14843;
wire n_14844;
wire n_14845;
wire n_14846;
wire n_14847;
wire n_14848;
wire n_14849;
wire n_14850;
wire n_14851;
wire n_14852;
wire n_14853;
wire n_14854;
wire n_14855;
wire n_14856;
wire n_14857;
wire n_14858;
wire n_14859;
wire n_14860;
wire n_14861;
wire n_14862;
wire n_14863;
wire n_14864;
wire n_14865;
wire n_14866;
wire n_14867;
wire n_14868;
wire n_14869;
wire n_14870;
wire n_14871;
wire n_14872;
wire n_14873;
wire n_14874;
wire n_14875;
wire n_14876;
wire n_14877;
wire n_14878;
wire n_14879;
wire n_14880;
wire n_14881;
wire n_14882;
wire n_14883;
wire n_14884;
wire n_14885;
wire n_14886;
wire n_14887;
wire n_14888;
wire n_14889;
wire n_14890;
wire n_14891;
wire n_14892;
wire n_14893;
wire n_14894;
wire n_14895;
wire n_14896;
wire n_14897;
wire n_14898;
wire n_14899;
wire n_14900;
wire n_14901;
wire n_14902;
wire n_14903;
wire n_14904;
wire n_14905;
wire n_14906;
wire n_14907;
wire n_14908;
wire n_14909;
wire n_14910;
wire n_14911;
wire n_14912;
wire n_14913;
wire n_14914;
wire n_14915;
wire n_14916;
wire n_14917;
wire n_14918;
wire n_14919;
wire n_14920;
wire n_14921;
wire n_14922;
wire n_14923;
wire n_14924;
wire n_14925;
wire n_14926;
wire n_14927;
wire n_14928;
wire n_14929;
wire n_14930;
wire n_14931;
wire n_14932;
wire n_14933;
wire n_14934;
wire n_14935;
wire n_14936;
wire n_14937;
wire n_14938;
wire n_14939;
wire n_14940;
wire n_14941;
wire n_14942;
wire n_14943;
wire n_14944;
wire n_14945;
wire n_14946;
wire n_14947;
wire n_14948;
wire n_14949;
wire n_14950;
wire n_14951;
wire n_14952;
wire n_14953;
wire n_14954;
wire n_14955;
wire n_14956;
wire n_14957;
wire n_14958;
wire n_14959;
wire n_14960;
wire n_14961;
wire n_14962;
wire n_14963;
wire n_14964;
wire n_14965;
wire n_14966;
wire n_14967;
wire n_14968;
wire n_14969;
wire n_14970;
wire n_14971;
wire n_14972;
wire n_14973;
wire n_14974;
wire n_14975;
wire n_14976;
wire n_14977;
wire n_14978;
wire n_14979;
wire n_14980;
wire n_14981;
wire n_14982;
wire n_14983;
wire n_14984;
wire n_14985;
wire n_14986;
wire n_14987;
wire n_14988;
wire n_14989;
wire n_14990;
wire n_14991;
wire n_14992;
wire n_14993;
wire n_14994;
wire n_14995;
wire n_14996;
wire n_14997;
wire n_14998;
wire n_14999;
wire n_15000;
wire n_15001;
wire n_15002;
wire n_15003;
wire n_15004;
wire n_15005;
wire n_15006;
wire n_15007;
wire n_15008;
wire n_15009;
wire n_15010;
wire n_15011;
wire n_15012;
wire n_15013;
wire n_15014;
wire n_15015;
wire n_15016;
wire n_15017;
wire n_15018;
wire n_15019;
wire n_15020;
wire n_15021;
wire n_15022;
wire n_15023;
wire n_15024;
wire n_15025;
wire n_15026;
wire n_15027;
wire n_15028;
wire n_15029;
wire n_15030;
wire n_15031;
wire n_15032;
wire n_15033;
wire n_15034;
wire n_15035;
wire n_15036;
wire n_15037;
wire n_15038;
wire n_15039;
wire n_15040;
wire n_15041;
wire n_15042;
wire n_15043;
wire n_15044;
wire n_15045;
wire n_15046;
wire n_15047;
wire n_15048;
wire n_15049;
wire n_15050;
wire n_15051;
wire n_15052;
wire n_15053;
wire n_15054;
wire n_15055;
wire n_15056;
wire n_15057;
wire n_15058;
wire n_15059;
wire n_15060;
wire n_15061;
wire n_15062;
wire n_15063;
wire n_15064;
wire n_15065;
wire n_15066;
wire n_15067;
wire n_15068;
wire n_15069;
wire n_15070;
wire n_15071;
wire n_15072;
wire n_15073;
wire n_15074;
wire n_15075;
wire n_15076;
wire n_15077;
wire n_15078;
wire n_15079;
wire n_15080;
wire n_15081;
wire n_15082;
wire n_15083;
wire n_15084;
wire n_15085;
wire n_15086;
wire n_15087;
wire n_15088;
wire n_15089;
wire n_15090;
wire n_15091;
wire n_15092;
wire n_15093;
wire n_15094;
wire n_15095;
wire n_15096;
wire n_15097;
wire n_15098;
wire n_15099;
wire n_15100;
wire n_15101;
wire n_15102;
wire n_15103;
wire n_15104;
wire n_15105;
wire n_15106;
wire n_15107;
wire n_15108;
wire n_15109;
wire n_15110;
wire n_15111;
wire n_15112;
wire n_15113;
wire n_15114;
wire n_15115;
wire n_15116;
wire n_15117;
wire n_15118;
wire n_15119;
wire n_15120;
wire n_15121;
wire n_15122;
wire n_15123;
wire n_15124;
wire n_15125;
wire n_15126;
wire n_15127;
wire n_15128;
wire n_15129;
wire n_15130;
wire n_15131;
wire n_15132;
wire n_15133;
wire n_15134;
wire n_15135;
wire n_15136;
wire n_15137;
wire n_15138;
wire n_15139;
wire n_15140;
wire n_15141;
wire n_15142;
wire n_15143;
wire n_15144;
wire n_15145;
wire n_15146;
wire n_15147;
wire n_15148;
wire n_15149;
wire n_15150;
wire n_15151;
wire n_15152;
wire n_15153;
wire n_15154;
wire n_15155;
wire n_15156;
wire n_15157;
wire n_15158;
wire n_15159;
wire n_15160;
wire n_15161;
wire n_15162;
wire n_15163;
wire n_15164;
wire n_15165;
wire n_15166;
wire n_15167;
wire n_15168;
wire n_15169;
wire n_15170;
wire n_15171;
wire n_15172;
wire n_15173;
wire n_15174;
wire n_15175;
wire n_15176;
wire n_15177;
wire n_15178;
wire n_15179;
wire n_15180;
wire n_15181;
wire n_15182;
wire n_15183;
wire n_15184;
wire n_15185;
wire n_15186;
wire n_15187;
wire n_15188;
wire n_15189;
wire n_15190;
wire n_15191;
wire n_15192;
wire n_15193;
wire n_15194;
wire n_15195;
wire n_15196;
wire n_15197;
wire n_15198;
wire n_15199;
wire n_15200;
wire n_15201;
wire n_15202;
wire n_15203;
wire n_15204;
wire n_15205;
wire n_15206;
wire n_15207;
wire n_15208;
wire n_15209;
wire n_15210;
wire n_15211;
wire n_15212;
wire n_15213;
wire n_15214;
wire n_15215;
wire n_15216;
wire n_15217;
wire n_15218;
wire n_15219;
wire n_15220;
wire n_15221;
wire n_15222;
wire n_15223;
wire n_15224;
wire n_15225;
wire n_15226;
wire n_15227;
wire n_15228;
wire n_15229;
wire n_15230;
wire n_15231;
wire n_15232;
wire n_15233;
wire n_15234;
wire n_15235;
wire n_15236;
wire n_15237;
wire n_15238;
wire n_15239;
wire n_15240;
wire n_15241;
wire n_15242;
wire n_15243;
wire n_15244;
wire n_15245;
wire n_15246;
wire n_15247;
wire n_15248;
wire n_15249;
wire n_15250;
wire n_15251;
wire n_15252;
wire n_15253;
wire n_15254;
wire n_15255;
wire n_15256;
wire n_15257;
wire n_15258;
wire n_15259;
wire n_15260;
wire n_15261;
wire n_15262;
wire n_15263;
wire n_15264;
wire n_15265;
wire n_15266;
wire n_15267;
wire n_15268;
wire n_15269;
wire n_15270;
wire n_15271;
wire n_15272;
wire n_15273;
wire n_15274;
wire n_15275;
wire n_15276;
wire n_15277;
wire n_15278;
wire n_15279;
wire n_15280;
wire n_15281;
wire n_15282;
wire n_15283;
wire n_15284;
wire n_15285;
wire n_15286;
wire n_15287;
wire n_15288;
wire n_15289;
wire n_15290;
wire n_15291;
wire n_15292;
wire n_15293;
wire n_15294;
wire n_15295;
wire n_15296;
wire n_15297;
wire n_15298;
wire n_15299;
wire n_15300;
wire n_15301;
wire n_15302;
wire n_15303;
wire n_15304;
wire n_15305;
wire n_15306;
wire n_15307;
wire n_15308;
wire n_15309;
wire n_15310;
wire n_15311;
wire n_15312;
wire n_15313;
wire n_15314;
wire n_15315;
wire n_15316;
wire n_15317;
wire n_15318;
wire n_15319;
wire n_15320;
wire n_15321;
wire n_15322;
wire n_15323;
wire n_15324;
wire n_15325;
wire n_15326;
wire n_15327;
wire n_15328;
wire n_15329;
wire n_15330;
wire n_15331;
wire n_15332;
wire n_15333;
wire n_15334;
wire n_15335;
wire n_15336;
wire n_15337;
wire n_15338;
wire n_15339;
wire n_15340;
wire n_15341;
wire n_15342;
wire n_15343;
wire n_15344;
wire n_15345;
wire n_15346;
wire n_15347;
wire n_15348;
wire n_15349;
wire n_15350;
wire n_15351;
wire n_15352;
wire n_15353;
wire n_15354;
wire n_15355;
wire n_15356;
wire n_15357;
wire n_15358;
wire n_15359;
wire n_15360;
wire n_15361;
wire n_15362;
wire n_15363;
wire n_15364;
wire n_15365;
wire n_15366;
wire n_15367;
wire n_15368;
wire n_15369;
wire n_15370;
wire n_15371;
wire n_15372;
wire n_15373;
wire n_15374;
wire n_15375;
wire n_15376;
wire n_15377;
wire n_15378;
wire n_15379;
wire n_15380;
wire n_15381;
wire n_15382;
wire n_15383;
wire n_15384;
wire n_15385;
wire n_15386;
wire n_15387;
wire n_15388;
wire n_15389;
wire n_15390;
wire n_15391;
wire n_15392;
wire n_15393;
wire n_15394;
wire n_15395;
wire n_15396;
wire n_15397;
wire n_15398;
wire n_15399;
wire n_15400;
wire n_15401;
wire n_15402;
wire n_15403;
wire n_15404;
wire n_15405;
wire n_15406;
wire n_15407;
wire n_15408;
wire n_15409;
wire n_15410;
wire n_15411;
wire n_15412;
wire n_15413;
wire n_15414;
wire n_15415;
wire n_15416;
wire n_15417;
wire n_15418;
wire n_15419;
wire n_15420;
wire n_15421;
wire n_15422;
wire n_15423;
wire n_15424;
wire n_15425;
wire n_15426;
wire n_15427;
wire n_15428;
wire n_15429;
wire n_15430;
wire n_15431;
wire n_15432;
wire n_15433;
wire n_15434;
wire n_15435;
wire n_15436;
wire n_15437;
wire n_15438;
wire n_15439;
wire n_15440;
wire n_15441;
wire n_15442;
wire n_15443;
wire n_15444;
wire n_15445;
wire n_15446;
wire n_15447;
wire n_15448;
wire n_15449;
wire n_15450;
wire n_15451;
wire n_15452;
wire n_15453;
wire n_15454;
wire n_15455;
wire n_15456;
wire n_15457;
wire n_15458;
wire n_15459;
wire n_15460;
wire n_15461;
wire n_15462;
wire n_15463;
wire n_15464;
wire n_15465;
wire n_15466;
wire n_15467;
wire n_15468;
wire n_15469;
wire n_15470;
wire n_15471;
wire n_15472;
wire n_15473;
wire n_15474;
wire n_15475;
wire n_15476;
wire n_15477;
wire n_15478;
wire n_15479;
wire n_15480;
wire n_15481;
wire n_15482;
wire n_15483;
wire n_15484;
wire n_15485;
wire n_15486;
wire n_15487;
wire n_15488;
wire n_15489;
wire n_15490;
wire n_15491;
wire n_15492;
wire n_15493;
wire n_15494;
wire n_15495;
wire n_15496;
wire n_15497;
wire n_15498;
wire n_15499;
wire n_15500;
wire n_15501;
wire n_15502;
wire n_15503;
wire n_15504;
wire n_15505;
wire n_15506;
wire n_15507;
wire n_15508;
wire n_15509;
wire n_15510;
wire n_15511;
wire n_15512;
wire n_15513;
wire n_15514;
wire n_15515;
wire n_15516;
wire n_15517;
wire n_15518;
wire n_15519;
wire n_15520;
wire n_15521;
wire n_15522;
wire n_15523;
wire n_15524;
wire n_15525;
wire n_15526;
wire n_15527;
wire n_15528;
wire n_15529;
wire n_15530;
wire n_15531;
wire n_15532;
wire n_15533;
wire n_15534;
wire n_15535;
wire n_15536;
wire n_15537;
wire n_15538;
wire n_15539;
wire n_15540;
wire n_15541;
wire n_15542;
wire n_15543;
wire n_15544;
wire n_15545;
wire n_15546;
wire n_15547;
wire n_15548;
wire n_15549;
wire n_15550;
wire n_15551;
wire n_15552;
wire n_15553;
wire n_15554;
wire n_15555;
wire n_15556;
wire n_15557;
wire n_15558;
wire n_15559;
wire n_15560;
wire n_15561;
wire n_15562;
wire n_15563;
wire n_15564;
wire n_15565;
wire n_15566;
wire n_15567;
wire n_15568;
wire n_15569;
wire n_15570;
wire n_15571;
wire n_15572;
wire n_15573;
wire n_15574;
wire n_15575;
wire n_15576;
wire n_15577;
wire n_15578;
wire n_15579;
wire n_15580;
wire n_15581;
wire n_15582;
wire n_15583;
wire n_15584;
wire n_15585;
wire n_15586;
wire n_15587;
wire n_15588;
wire n_15589;
wire n_15590;
wire n_15591;
wire n_15592;
wire n_15593;
wire n_15594;
wire n_15595;
wire n_15596;
wire n_15597;
wire n_15598;
wire n_15599;
wire n_15600;
wire n_15601;
wire n_15602;
wire n_15603;
wire n_15604;
wire n_15605;
wire n_15606;
wire n_15607;
wire n_15608;
wire n_15609;
wire n_15610;
wire n_15611;
wire n_15612;
wire n_15613;
wire n_15614;
wire n_15615;
wire n_15616;
wire n_15617;
wire n_15618;
wire n_15619;
wire n_15620;
wire n_15621;
wire n_15622;
wire n_15623;
wire n_15624;
wire n_15625;
wire n_15626;
wire n_15627;
wire n_15628;
wire n_15629;
wire n_15630;
wire n_15631;
wire n_15632;
wire n_15633;
wire n_15634;
wire n_15635;
wire n_15636;
wire n_15637;
wire n_15638;
wire n_15639;
wire n_15640;
wire n_15641;
wire n_15642;
wire n_15643;
wire n_15644;
wire n_15645;
wire n_15646;
wire n_15647;
wire n_15648;
wire n_15649;
wire n_15650;
wire n_15651;
wire n_15652;
wire n_15653;
wire n_15654;
wire n_15655;
wire n_15656;
wire n_15657;
wire n_15658;
wire n_15659;
wire n_15660;
wire n_15661;
wire n_15662;
wire n_15663;
wire n_15664;
wire n_15665;
wire n_15666;
wire n_15667;
wire n_15668;
wire n_15669;
wire n_15670;
wire n_15671;
wire n_15672;
wire n_15673;
wire n_15674;
wire n_15675;
wire n_15676;
wire n_15677;
wire n_15678;
wire n_15679;
wire n_15680;
wire n_15681;
wire n_15682;
wire n_15683;
wire n_15684;
wire n_15685;
wire n_15686;
wire n_15687;
wire n_15688;
wire n_15689;
wire n_15690;
wire n_15691;
wire n_15692;
wire n_15693;
wire n_15694;
wire n_15695;
wire n_15696;
wire n_15697;
wire n_15698;
wire n_15699;
wire n_15700;
wire n_15701;
wire n_15702;
wire n_15703;
wire n_15704;
wire n_15705;
wire n_15706;
wire n_15707;
wire n_15708;
wire n_15709;
wire n_15710;
wire n_15711;
wire n_15712;
wire n_15713;
wire n_15714;
wire n_15715;
wire n_15716;
wire n_15717;
wire n_15718;
wire n_15719;
wire n_15720;
wire n_15721;
wire n_15722;
wire n_15723;
wire n_15724;
wire n_15725;
wire n_15726;
wire n_15727;
wire n_15728;
wire n_15729;
wire n_15730;
wire n_15731;
wire n_15732;
wire n_15733;
wire n_15734;
wire n_15735;
wire n_15736;
wire n_15737;
wire n_15738;
wire n_15739;
wire n_15740;
wire n_15741;
wire n_15742;
wire n_15743;
wire n_15744;
wire n_15745;
wire n_15746;
wire n_15747;
wire n_15748;
wire n_15749;
wire n_15750;
wire n_15751;
wire n_15752;
wire n_15753;
wire n_15754;
wire n_15755;
wire n_15756;
wire n_15757;
wire n_15758;
wire n_15759;
wire n_15760;
wire n_15761;
wire n_15762;
wire n_15763;
wire n_15764;
wire n_15765;
wire n_15766;
wire n_15767;
wire n_15768;
wire n_15769;
wire n_15770;
wire n_15771;
wire n_15772;
wire n_15773;
wire n_15774;
wire n_15775;
wire n_15776;
wire n_15777;
wire n_15778;
wire n_15779;
wire n_15780;
wire n_15781;
wire n_15782;
wire n_15783;
wire n_15784;
wire n_15785;
wire n_15786;
wire n_15787;
wire n_15788;
wire n_15789;
wire n_15790;
wire n_15791;
wire n_15792;
wire n_15793;
wire n_15794;
wire n_15795;
wire n_15796;
wire n_15797;
wire n_15798;
wire n_15799;
wire n_15800;
wire n_15801;
wire n_15802;
wire n_15803;
wire n_15804;
wire n_15805;
wire n_15806;
wire n_15807;
wire n_15808;
wire n_15809;
wire n_15810;
wire n_15811;
wire n_15812;
wire n_15813;
wire n_15814;
wire n_15815;
wire n_15816;
wire n_15817;
wire n_15818;
wire n_15819;
wire n_15820;
wire n_15821;
wire n_15822;
wire n_15823;
wire n_15824;
wire n_15825;
wire n_15826;
wire n_15827;
wire n_15828;
wire n_15829;
wire n_15830;
wire n_15831;
wire n_15832;
wire n_15833;
wire n_15834;
wire n_15835;
wire n_15836;
wire n_15837;
wire n_15838;
wire n_15839;
wire n_15840;
wire n_15841;
wire n_15842;
wire n_15843;
wire n_15844;
wire n_15845;
wire n_15846;
wire n_15847;
wire n_15848;
wire n_15849;
wire n_15850;
wire n_15851;
wire n_15852;
wire n_15853;
wire n_15854;
wire n_15855;
wire n_15856;
wire n_15857;
wire n_15858;
wire n_15859;
wire n_15860;
wire n_15861;
wire n_15862;
wire n_15863;
wire n_15864;
wire n_15865;
wire n_15866;
wire n_15867;
wire n_15868;
wire n_15869;
wire n_15870;
wire n_15871;
wire n_15872;
wire n_15873;
wire n_15874;
wire n_15875;
wire n_15876;
wire n_15877;
wire n_15878;
wire n_15879;
wire n_15880;
wire n_15881;
wire n_15882;
wire n_15883;
wire n_15884;
wire n_15885;
wire n_15886;
wire n_15887;
wire n_15888;
wire n_15889;
wire n_15890;
wire n_15891;
wire n_15892;
wire n_15893;
wire n_15894;
wire n_15895;
wire n_15896;
wire n_15897;
wire n_15898;
wire n_15899;
wire n_15900;
wire n_15901;
wire n_15902;
wire n_15903;
wire n_15904;
wire n_15905;
wire n_15906;
wire n_15907;
wire n_15908;
wire n_15909;
wire n_15910;
wire n_15911;
wire n_15912;
wire n_15913;
wire n_15914;
wire n_15915;
wire n_15916;
wire n_15917;
wire n_15918;
wire n_15919;
wire n_15920;
wire n_15921;
wire n_15922;
wire n_15923;
wire n_15924;
wire n_15925;
wire n_15926;
wire n_15927;
wire n_15928;
wire n_15929;
wire n_15930;
wire n_15931;
wire n_15932;
wire n_15933;
wire n_15934;
wire n_15935;
wire n_15936;
wire n_15937;
wire n_15938;
wire n_15939;
wire n_15940;
wire n_15941;
wire n_15942;
wire n_15943;
wire n_15944;
wire n_15945;
wire n_15946;
wire n_15947;
wire n_15948;
wire n_15949;
wire n_15950;
wire n_15951;
wire n_15952;
wire n_15953;
wire n_15954;
wire n_15955;
wire n_15956;
wire n_15957;
wire n_15958;
wire n_15959;
wire n_15960;
wire n_15961;
wire n_15962;
wire n_15963;
wire n_15964;
wire n_15965;
wire n_15966;
wire n_15967;
wire n_15968;
wire n_15969;
wire n_15970;
wire n_15971;
wire n_15972;
wire n_15973;
wire n_15974;
wire n_15975;
wire n_15976;
wire n_15977;
wire n_15978;
wire n_15979;
wire n_15980;
wire n_15981;
wire n_15982;
wire n_15983;
wire n_15984;
wire n_15985;
wire n_15986;
wire n_15987;
wire n_15988;
wire n_15989;
wire n_15990;
wire n_15991;
wire n_15992;
wire n_15993;
wire n_15994;
wire n_15995;
wire n_15996;
wire n_15997;
wire n_15998;
wire n_15999;
wire n_16000;
wire n_16001;
wire n_16002;
wire n_16003;
wire n_16004;
wire n_16005;
wire n_16006;
wire n_16007;
wire n_16008;
wire n_16009;
wire n_16010;
wire n_16011;
wire n_16012;
wire n_16013;
wire n_16014;
wire n_16015;
wire n_16016;
wire n_16017;
wire n_16018;
wire n_16019;
wire n_16020;
wire n_16021;
wire n_16022;
wire n_16023;
wire n_16024;
wire n_16025;
wire n_16026;
wire n_16027;
wire n_16028;
wire n_16029;
wire n_16030;
wire n_16031;
wire n_16032;
wire n_16033;
wire n_16034;
wire n_16035;
wire n_16036;
wire n_16037;
wire n_16038;
wire n_16039;
wire n_16040;
wire n_16041;
wire n_16042;
wire n_16043;
wire n_16044;
wire n_16045;
wire n_16046;
wire n_16047;
wire n_16048;
wire n_16049;
wire n_16050;
wire n_16051;
wire n_16052;
wire n_16053;
wire n_16054;
wire n_16055;
wire n_16056;
wire n_16057;
wire n_16058;
wire n_16059;
wire n_16060;
wire n_16061;
wire n_16062;
wire n_16063;
wire n_16064;
wire n_16065;
wire n_16066;
wire n_16067;
wire n_16068;
wire n_16069;
wire n_16070;
wire n_16071;
wire n_16072;
wire n_16073;
wire n_16074;
wire n_16075;
wire n_16076;
wire n_16077;
wire n_16078;
wire n_16079;
wire n_16080;
wire n_16081;
wire n_16082;
wire n_16083;
wire n_16084;
wire n_16085;
wire n_16086;
wire n_16087;
wire n_16088;
wire n_16089;
wire n_16090;
wire n_16091;
wire n_16092;
wire n_16093;
wire n_16094;
wire n_16095;
wire n_16096;
wire n_16097;
wire n_16098;
wire n_16099;
wire n_16100;
wire n_16101;
wire n_16102;
wire n_16103;
wire n_16104;
wire n_16105;
wire n_16106;
wire n_16107;
wire n_16108;
wire n_16109;
wire n_16110;
wire n_16111;
wire n_16112;
wire n_16113;
wire n_16114;
wire n_16115;
wire n_16116;
wire n_16117;
wire n_16118;
wire n_16119;
wire n_16120;
wire n_16121;
wire n_16122;
wire n_16123;
wire n_16124;
wire n_16125;
wire n_16126;
wire n_16127;
wire n_16128;
wire n_16129;
wire n_16130;
wire n_16131;
wire n_16132;
wire n_16133;
wire n_16134;
wire n_16135;
wire n_16136;
wire n_16137;
wire n_16138;
wire n_16139;
wire n_16140;
wire n_16141;
wire n_16142;
wire n_16143;
wire n_16144;
wire n_16145;
wire n_16146;
wire n_16147;
wire n_16148;
wire n_16149;
wire n_16150;
wire n_16151;
wire n_16152;
wire n_16153;
wire n_16154;
wire n_16155;
wire n_16156;
wire n_16157;
wire n_16158;
wire n_16159;
wire n_16160;
wire n_16161;
wire n_16162;
wire n_16163;
wire n_16164;
wire n_16165;
wire n_16166;
wire n_16167;
wire n_16168;
wire n_16169;
wire n_16170;
wire n_16171;
wire n_16172;
wire n_16173;
wire n_16174;
wire n_16175;
wire n_16176;
wire n_16177;
wire n_16178;
wire n_16179;
wire n_16180;
wire n_16181;
wire n_16182;
wire n_16183;
wire n_16184;
wire n_16185;
wire n_16186;
wire n_16187;
wire n_16188;
wire n_16189;
wire n_16190;
wire n_16191;
wire n_16192;
wire n_16193;
wire n_16194;
wire n_16195;
wire n_16196;
wire n_16197;
wire n_16198;
wire n_16199;
wire n_16200;
wire n_16201;
wire n_16202;
wire n_16203;
wire n_16204;
wire n_16205;
wire n_16206;
wire n_16207;
wire n_16208;
wire n_16209;
wire n_16210;
wire n_16211;
wire n_16212;
wire n_16213;
wire n_16214;
wire n_16215;
wire n_16216;
wire n_16217;
wire n_16218;
wire n_16219;
wire n_16220;
wire n_16221;
wire n_16222;
wire n_16223;
wire n_16224;
wire n_16225;
wire n_16226;
wire n_16227;
wire n_16228;
wire n_16229;
wire n_16230;
wire n_16231;
wire n_16232;
wire n_16233;
wire n_16234;
wire n_16235;
wire n_16236;
wire n_16237;
wire n_16238;
wire n_16239;
wire n_16240;
wire n_16241;
wire n_16242;
wire n_16243;
wire n_16244;
wire n_16245;
wire n_16246;
wire n_16247;
wire n_16248;
wire n_16249;
wire n_16250;
wire n_16251;
wire n_16252;
wire n_16253;
wire n_16254;
wire n_16255;
wire n_16256;
wire n_16257;
wire n_16258;
wire n_16259;
wire n_16260;
wire n_16261;
wire n_16262;
wire n_16263;
wire n_16264;
wire n_16265;
wire n_16266;
wire n_16267;
wire n_16268;
wire n_16269;
wire n_16270;
wire n_16271;
wire n_16272;
wire n_16273;
wire n_16274;
wire n_16275;
wire n_16276;
wire n_16277;
wire n_16278;
wire n_16279;
wire n_16280;
wire n_16281;
wire n_16282;
wire n_16283;
wire n_16284;
wire n_16285;
wire n_16286;
wire n_16287;
wire n_16288;
wire n_16289;
wire n_16290;
wire n_16291;
wire n_16292;
wire n_16293;
wire n_16294;
wire n_16295;
wire n_16296;
wire n_16297;
wire n_16298;
wire n_16299;
wire n_16300;
wire n_16301;
wire n_16302;
wire n_16303;
wire n_16304;
wire n_16305;
wire n_16306;
wire n_16307;
wire n_16308;
wire n_16309;
wire n_16310;
wire n_16311;
wire n_16312;
wire n_16313;
wire n_16314;
wire n_16315;
wire n_16316;
wire n_16317;
wire n_16318;
wire n_16319;
wire n_16320;
wire n_16321;
wire n_16322;
wire n_16323;
wire n_16324;
wire n_16325;
wire n_16326;
wire n_16327;
wire n_16328;
wire n_16329;
wire n_16330;
wire n_16331;
wire n_16332;
wire n_16333;
wire n_16334;
wire n_16335;
wire n_16336;
wire n_16337;
wire n_16338;
wire n_16339;
wire n_16340;
wire n_16341;
wire n_16342;
wire n_16343;
wire n_16344;
wire n_16345;
wire n_16346;
wire n_16347;
wire n_16348;
wire n_16349;
wire n_16350;
wire n_16351;
wire n_16352;
wire n_16353;
wire n_16354;
wire n_16355;
wire n_16356;
wire n_16357;
wire n_16358;
wire n_16359;
wire n_16360;
wire n_16361;
wire n_16362;
wire n_16363;
wire n_16364;
wire n_16365;
wire n_16366;
wire n_16367;
wire n_16368;
wire n_16369;
wire n_16370;
wire n_16371;
wire n_16372;
wire n_16373;
wire n_16374;
wire n_16375;
wire n_16376;
wire n_16377;
wire n_16378;
wire n_16379;
wire n_16380;
wire n_16381;
wire n_16382;
wire n_16383;
wire n_16384;
wire n_16385;
wire n_16386;
wire n_16387;
wire n_16388;
wire n_16389;
wire n_16390;
wire n_16391;
wire n_16392;
wire n_16393;
wire n_16394;
wire n_16395;
wire n_16396;
wire n_16397;
wire n_16398;
wire n_16399;
wire n_16400;
wire n_16401;
wire n_16402;
wire n_16403;
wire n_16404;
wire n_16405;
wire n_16406;
wire n_16407;
wire n_16408;
wire n_16409;
wire n_16410;
wire n_16411;
wire n_16412;
wire n_16413;
wire n_16414;
wire n_16415;
wire n_16416;
wire n_16417;
wire n_16418;
wire n_16419;
wire n_16420;
wire n_16421;
wire n_16422;
wire n_16423;
wire n_16424;
wire n_16425;
wire n_16426;
wire n_16427;
wire n_16428;
wire n_16429;
wire n_16430;
wire n_16431;
wire n_16432;
wire n_16433;
wire n_16434;
wire n_16435;
wire n_16436;
wire n_16437;
wire n_16438;
wire n_16439;
wire n_16440;
wire n_16441;
wire n_16442;
wire n_16443;
wire n_16444;
wire n_16445;
wire n_16446;
wire n_16447;
wire n_16448;
wire n_16449;
wire n_16450;
wire n_16451;
wire n_16452;
wire n_16453;
wire n_16454;
wire n_16455;
wire n_16456;
wire n_16457;
wire n_16458;
wire n_16459;
wire n_16460;
wire n_16461;
wire n_16462;
wire n_16463;
wire n_16464;
wire n_16465;
wire n_16466;
wire n_16467;
wire n_16468;
wire n_16469;
wire n_16470;
wire n_16471;
wire n_16472;
wire n_16473;
wire n_16474;
wire n_16475;
wire n_16476;
wire n_16477;
wire n_16478;
wire n_16479;
wire n_16480;
wire n_16481;
wire n_16482;
wire n_16483;
wire n_16484;
wire n_16485;
wire n_16486;
wire n_16487;
wire n_16488;
wire n_16489;
wire n_16490;
wire n_16491;
wire n_16492;
wire n_16493;
wire n_16494;
wire n_16495;
wire n_16496;
wire n_16497;
wire n_16498;
wire n_16499;
wire n_16500;
wire n_16501;
wire n_16502;
wire n_16503;
wire n_16504;
wire n_16505;
wire n_16506;
wire n_16507;
wire n_16508;
wire n_16509;
wire n_16510;
wire n_16511;
wire n_16512;
wire n_16513;
wire n_16514;
wire n_16515;
wire n_16516;
wire n_16517;
wire n_16518;
wire n_16519;
wire n_16520;
wire n_16521;
wire n_16522;
wire n_16523;
wire n_16524;
wire n_16525;
wire n_16526;
wire n_16527;
wire n_16528;
wire n_16529;
wire n_16530;
wire n_16531;
wire n_16532;
wire n_16533;
wire n_16534;
wire n_16535;
wire n_16536;
wire n_16537;
wire n_16538;
wire n_16539;
wire n_16540;
wire n_16541;
wire n_16542;
wire n_16543;
wire n_16544;
wire n_16545;
wire n_16546;
wire n_16547;
wire n_16548;
wire n_16549;
wire n_16550;
wire n_16551;
wire n_16552;
wire n_16553;
wire n_16554;
wire n_16555;
wire n_16556;
wire n_16557;
wire n_16558;
wire n_16559;
wire n_16560;
wire n_16561;
wire n_16562;
wire n_16563;
wire n_16564;
wire n_16565;
wire n_16566;
wire n_16567;
wire n_16568;
wire n_16569;
wire n_16570;
wire n_16571;
wire n_16572;
wire n_16573;
wire n_16574;
wire n_16575;
wire n_16576;
wire n_16577;
wire n_16578;
wire n_16579;
wire n_16580;
wire n_16581;
wire n_16582;
wire n_16583;
wire n_16584;
wire n_16585;
wire n_16586;
wire n_16587;
wire n_16588;
wire n_16589;
wire n_16590;
wire n_16591;
wire n_16592;
wire n_16593;
wire n_16594;
wire n_16595;
wire n_16596;
wire n_16597;
wire n_16598;
wire n_16599;
wire n_16600;
wire n_16601;
wire n_16602;
wire n_16603;
wire n_16604;
wire n_16605;
wire n_16606;
wire n_16607;
wire n_16608;
wire n_16609;
wire n_16610;
wire n_16611;
wire n_16612;
wire n_16613;
wire n_16614;
wire n_16615;
wire n_16616;
wire n_16617;
wire n_16618;
wire n_16619;
wire n_16620;
wire n_16621;
wire n_16622;
wire n_16623;
wire n_16624;
wire n_16625;
wire n_16626;
wire n_16627;
wire n_16628;
wire n_16629;
wire n_16630;
wire n_16631;
wire n_16632;
wire n_16633;
wire n_16634;
wire n_16635;
wire n_16636;
wire n_16637;
wire n_16638;
wire n_16639;
wire n_16640;
wire n_16641;
wire n_16642;
wire n_16643;
wire n_16644;
wire n_16645;
wire n_16646;
wire n_16647;
wire n_16648;
wire n_16649;
wire n_16650;
wire n_16651;
wire n_16652;
wire n_16653;
wire n_16654;
wire n_16655;
wire n_16656;
wire n_16657;
wire n_16658;
wire n_16659;
wire n_16660;
wire n_16661;
wire n_16662;
wire n_16663;
wire n_16664;
wire n_16665;
wire n_16666;
wire n_16667;
wire n_16668;
wire n_16669;
wire n_16670;
wire n_16671;
wire n_16672;
wire n_16673;
wire n_16674;
wire n_16675;
wire n_16676;
wire n_16677;
wire n_16678;
wire n_16679;
wire n_16680;
wire n_16681;
wire n_16682;
wire n_16683;
wire n_16684;
wire n_16685;
wire n_16686;
wire n_16687;
wire n_16688;
wire n_16689;
wire n_16690;
wire n_16691;
wire n_16692;
wire n_16693;
wire n_16694;
wire n_16695;
wire n_16696;
wire n_16697;
wire n_16698;
wire n_16699;
wire n_16700;
wire n_16701;
wire n_16702;
wire n_16703;
wire n_16704;
wire n_16705;
wire n_16706;
wire n_16707;
wire n_16708;
wire n_16709;
wire n_16710;
wire n_16711;
wire n_16712;
wire n_16713;
wire n_16714;
wire n_16715;
wire n_16716;
wire n_16717;
wire n_16718;
wire n_16719;
wire n_16720;
wire n_16721;
wire n_16722;
wire n_16723;
wire n_16724;
wire n_16725;
wire n_16726;
wire n_16727;
wire n_16728;
wire n_16729;
wire n_16730;
wire n_16731;
wire n_16732;
wire n_16733;
wire n_16734;
wire n_16735;
wire n_16736;
wire n_16737;
wire n_16738;
wire n_16739;
wire n_16740;
wire n_16741;
wire n_16742;
wire n_16743;
wire n_16744;
wire n_16745;
wire n_16746;
wire n_16747;
wire n_16748;
wire n_16749;
wire n_16750;
wire n_16751;
wire n_16752;
wire n_16753;
wire n_16754;
wire n_16755;
wire n_16756;
wire n_16757;
wire n_16758;
wire n_16759;
wire n_16760;
wire n_16761;
wire n_16762;
wire n_16763;
wire n_16764;
wire n_16765;
wire n_16766;
wire n_16767;
wire n_16768;
wire n_16769;
wire n_16770;
wire n_16771;
wire n_16772;
wire n_16773;
wire n_16774;
wire n_16775;
wire n_16776;
wire n_16777;
wire n_16778;
wire n_16779;
wire n_16780;
wire n_16781;
wire n_16782;
wire n_16783;
wire n_16784;
wire n_16785;
wire n_16786;
wire n_16787;
wire n_16788;
wire n_16789;
wire n_16790;
wire n_16791;
wire n_16792;
wire n_16793;
wire n_16794;
wire n_16795;
wire n_16796;
wire n_16797;
wire n_16798;
wire n_16799;
wire n_16800;
wire n_16801;
wire n_16802;
wire n_16803;
wire n_16804;
wire n_16805;
wire n_16806;
wire n_16807;
wire n_16808;
wire n_16809;
wire n_16810;
wire n_16811;
wire n_16812;
wire n_16813;
wire n_16814;
wire n_16815;
wire n_16816;
wire n_16817;
wire n_16818;
wire n_16819;
wire n_16820;
wire n_16821;
wire n_16822;
wire n_16823;
wire n_16824;
wire n_16825;
wire n_16826;
wire n_16827;
wire n_16828;
wire n_16829;
wire n_16830;
wire n_16831;
wire n_16832;
wire n_16833;
wire n_16834;
wire n_16835;
wire n_16836;
wire n_16837;
wire n_16838;
wire n_16839;
wire n_16840;
wire n_16841;
wire n_16842;
wire n_16843;
wire n_16844;
wire n_16845;
wire n_16846;
wire n_16847;
wire n_16848;
wire n_16849;
wire n_16850;
wire n_16851;
wire n_16852;
wire n_16853;
wire n_16854;
wire n_16855;
wire n_16856;
wire n_16857;
wire n_16858;
wire n_16859;
wire n_16860;
wire n_16861;
wire n_16862;
wire n_16863;
wire n_16864;
wire n_16865;
wire n_16866;
wire n_16867;
wire n_16868;
wire n_16869;
wire n_16870;
wire n_16871;
wire n_16872;
wire n_16873;
wire n_16874;
wire n_16875;
wire n_16876;
wire n_16877;
wire n_16878;
wire n_16879;
wire n_16880;
wire n_16881;
wire n_16882;
wire n_16883;
wire n_16884;
wire n_16885;
wire n_16886;
wire n_16887;
wire n_16888;
wire n_16889;
wire n_16890;
wire n_16891;
wire n_16892;
wire n_16893;
wire n_16894;
wire n_16895;
wire n_16896;
wire n_16897;
wire n_16898;
wire n_16899;
wire n_16900;
wire n_16901;
wire n_16902;
wire n_16903;
wire n_16904;
wire n_16905;
wire n_16906;
wire n_16907;
wire n_16908;
wire n_16909;
wire n_16910;
wire n_16911;
wire n_16912;
wire n_16913;
wire n_16914;
wire n_16915;
wire n_16916;
wire n_16917;
wire n_16918;
wire n_16919;
wire n_16920;
wire n_16921;
wire n_16922;
wire n_16923;
wire n_16924;
wire n_16925;
wire n_16926;
wire n_16927;
wire n_16928;
wire n_16929;
wire n_16930;
wire n_16931;
wire n_16932;
wire n_16933;
wire n_16934;
wire n_16935;
wire n_16936;
wire n_16937;
wire n_16938;
wire n_16939;
wire n_16940;
wire n_16941;
wire n_16942;
wire n_16943;
wire n_16944;
wire n_16945;
wire n_16946;
wire n_16947;
wire n_16948;
wire n_16949;
wire n_16950;
wire n_16951;
wire n_16952;
wire n_16953;
wire n_16954;
wire n_16955;
wire n_16956;
wire n_16957;
wire n_16958;
wire n_16959;
wire n_16960;
wire n_16961;
wire n_16962;
wire n_16963;
wire n_16964;
wire n_16965;
wire n_16966;
wire n_16967;
wire n_16968;
wire n_16969;
wire n_16970;
wire n_16971;
wire n_16972;
wire n_16973;
wire n_16974;
wire n_16975;
wire n_16976;
wire n_16977;
wire n_16978;
wire n_16979;
wire n_16980;
wire n_16981;
wire n_16982;
wire n_16983;
wire n_16984;
wire n_16985;
wire n_16986;
wire n_16987;
wire n_16988;
wire n_16989;
wire n_16990;
wire n_16991;
wire n_16992;
wire n_16993;
wire n_16994;
wire n_16995;
wire n_16996;
wire n_16997;
wire n_16998;
wire n_16999;
wire n_17000;
wire n_17001;
wire n_17002;
wire n_17003;
wire n_17004;
wire n_17005;
wire n_17006;
wire n_17007;
wire n_17008;
wire n_17009;
wire n_17010;
wire n_17011;
wire n_17012;
wire n_17013;
wire n_17014;
wire n_17015;
wire n_17016;
wire n_17017;
wire n_17018;
wire n_17019;
wire n_17020;
wire n_17021;
wire n_17022;
wire n_17023;
wire n_17024;
wire n_17025;
wire n_17026;
wire n_17027;
wire n_17028;
wire n_17029;
wire n_17030;
wire n_17031;
wire n_17032;
wire n_17033;
wire n_17034;
wire n_17035;
wire n_17036;
wire n_17037;
wire n_17038;
wire n_17039;
wire n_17040;
wire n_17041;
wire n_17042;
wire n_17043;
wire n_17044;
wire n_17045;
wire n_17046;
wire n_17047;
wire n_17048;
wire n_17049;
wire n_17050;
wire n_17051;
wire n_17052;
wire n_17053;
wire n_17054;
wire n_17055;
wire n_17056;
wire n_17057;
wire n_17058;
wire n_17059;
wire n_17060;
wire n_17061;
wire n_17062;
wire n_17063;
wire n_17064;
wire n_17065;
wire n_17066;
wire n_17067;
wire n_17068;
wire n_17069;
wire n_17070;
wire n_17071;
wire n_17072;
wire n_17073;
wire n_17074;
wire n_17075;
wire n_17076;
wire n_17077;
wire n_17078;
wire n_17079;
wire n_17080;
wire n_17081;
wire n_17082;
wire n_17083;
wire n_17084;
wire n_17085;
wire n_17086;
wire n_17087;
wire n_17088;
wire n_17089;
wire n_17090;
wire n_17091;
wire n_17092;
wire n_17093;
wire n_17094;
wire n_17095;
wire n_17096;
wire n_17097;
wire n_17098;
wire n_17099;
wire n_17100;
wire n_17101;
wire n_17102;
wire n_17103;
wire n_17104;
wire n_17105;
wire n_17106;
wire n_17107;
wire n_17108;
wire n_17109;
wire n_17110;
wire n_17111;
wire n_17112;
wire n_17113;
wire n_17114;
wire n_17115;
wire n_17116;
wire n_17117;
wire n_17118;
wire n_17119;
wire n_17120;
wire n_17121;
wire n_17122;
wire n_17123;
wire n_17124;
wire n_17125;
wire n_17126;
wire n_17127;
wire n_17128;
wire n_17129;
wire n_17130;
wire n_17131;
wire n_17132;
wire n_17133;
wire n_17134;
wire n_17135;
wire n_17136;
wire n_17137;
wire n_17138;
wire n_17139;
wire n_17140;
wire n_17141;
wire n_17142;
wire n_17143;
wire n_17144;
wire n_17145;
wire n_17146;
wire n_17147;
wire n_17148;
wire n_17149;
wire n_17150;
wire n_17151;
wire n_17152;
wire n_17153;
wire n_17154;
wire n_17155;
wire n_17156;
wire n_17157;
wire n_17158;
wire n_17159;
wire n_17160;
wire n_17161;
wire n_17162;
wire n_17163;
wire n_17164;
wire n_17165;
wire n_17166;
wire n_17167;
wire n_17168;
wire n_17169;
wire n_17170;
wire n_17171;
wire n_17172;
wire n_17173;
wire n_17174;
wire n_17175;
wire n_17176;
wire n_17177;
wire n_17178;
wire n_17179;
wire n_17180;
wire n_17181;
wire n_17182;
wire n_17183;
wire n_17184;
wire n_17185;
wire n_17186;
wire n_17187;
wire n_17188;
wire n_17189;
wire n_17190;
wire n_17191;
wire n_17192;
wire n_17193;
wire n_17194;
wire n_17195;
wire n_17196;
wire n_17197;
wire n_17198;
wire n_17199;
wire n_17200;
wire n_17201;
wire n_17202;
wire n_17203;
wire n_17204;
wire n_17205;
wire n_17206;
wire n_17207;
wire n_17208;
wire n_17209;
wire n_17210;
wire n_17211;
wire n_17212;
wire n_17213;
wire n_17214;
wire n_17215;
wire n_17216;
wire n_17217;
wire n_17218;
wire n_17219;
wire n_17220;
wire n_17221;
wire n_17222;
wire n_17223;
wire n_17224;
wire n_17225;
wire n_17226;
wire n_17227;
wire n_17228;
wire n_17229;
wire n_17230;
wire n_17231;
wire n_17232;
wire n_17233;
wire n_17234;
wire n_17235;
wire n_17236;
wire n_17237;
wire n_17238;
wire n_17239;
wire n_17240;
wire n_17241;
wire n_17242;
wire n_17243;
wire n_17244;
wire n_17245;
wire n_17246;
wire n_17247;
wire n_17248;
wire n_17249;
wire n_17250;
wire n_17251;
wire n_17252;
wire n_17253;
wire n_17254;
wire n_17255;
wire n_17256;
wire n_17257;
wire n_17258;
wire n_17259;
wire n_17260;
wire n_17261;
wire n_17262;
wire n_17263;
wire n_17264;
wire n_17265;
wire n_17266;
wire n_17267;
wire n_17268;
wire n_17269;
wire n_17270;
wire n_17271;
wire n_17272;
wire n_17273;
wire n_17274;
wire n_17275;
wire n_17276;
wire n_17277;
wire n_17278;
wire n_17279;
wire n_17280;
wire n_17281;
wire n_17282;
wire n_17283;
wire n_17284;
wire n_17285;
wire n_17286;
wire n_17287;
wire n_17288;
wire n_17289;
wire n_17290;
wire n_17291;
wire n_17292;
wire n_17293;
wire n_17294;
wire n_17295;
wire n_17296;
wire n_17297;
wire n_17298;
wire n_17299;
wire n_17300;
wire n_17301;
wire n_17302;
wire n_17303;
wire n_17304;
wire n_17305;
wire n_17306;
wire n_17307;
wire n_17308;
wire n_17309;
wire n_17310;
wire n_17311;
wire n_17312;
wire n_17313;
wire n_17314;
wire n_17315;
wire n_17316;
wire n_17317;
wire n_17318;
wire n_17319;
wire n_17320;
wire n_17321;
wire n_17322;
wire n_17323;
wire n_17324;
wire n_17325;
wire n_17326;
wire n_17327;
wire n_17328;
wire n_17329;
wire n_17330;
wire n_17331;
wire n_17332;
wire n_17333;
wire n_17334;
wire n_17335;
wire n_17336;
wire n_17337;
wire n_17338;
wire n_17339;
wire n_17340;
wire n_17341;
wire n_17342;
wire n_17343;
wire n_17344;
wire n_17345;
wire n_17346;
wire n_17347;
wire n_17348;
wire n_17349;
wire n_17350;
wire n_17351;
wire n_17352;
wire n_17353;
wire n_17354;
wire n_17355;
wire n_17356;
wire n_17357;
wire n_17358;
wire n_17359;
wire n_17360;
wire n_17361;
wire n_17362;
wire n_17363;
wire n_17364;
wire n_17365;
wire n_17366;
wire n_17367;
wire n_17368;
wire n_17369;
wire n_17370;
wire n_17371;
wire n_17372;
wire n_17373;
wire n_17374;
wire n_17375;
wire n_17376;
wire n_17377;
wire n_17378;
wire n_17379;
wire n_17380;
wire n_17381;
wire n_17382;
wire n_17383;
wire n_17384;
wire n_17385;
wire n_17386;
wire n_17387;
wire n_17388;
wire n_17389;
wire n_17390;
wire n_17391;
wire n_17392;
wire n_17393;
wire n_17394;
wire n_17395;
wire n_17396;
wire n_17397;
wire n_17398;
wire n_17399;
wire n_17400;
wire n_17401;
wire n_17402;
wire n_17403;
wire n_17404;
wire n_17405;
wire n_17406;
wire n_17407;
wire n_17408;
wire n_17409;
wire n_17410;
wire n_17411;
wire n_17412;
wire n_17413;
wire n_17414;
wire n_17415;
wire n_17416;
wire n_17417;
wire n_17418;
wire n_17419;
wire n_17420;
wire n_17421;
wire n_17422;
wire n_17423;
wire n_17424;
wire n_17425;
wire n_17426;
wire n_17427;
wire n_17428;
wire n_17429;
wire n_17430;
wire n_17431;
wire n_17432;
wire n_17433;
wire n_17434;
wire n_17435;
wire n_17436;
wire n_17437;
wire n_17438;
wire n_17439;
wire n_17440;
wire n_17441;
wire n_17442;
wire n_17443;
wire n_17444;
wire n_17445;
wire n_17446;
wire n_17447;
wire n_17448;
wire n_17449;
wire n_17450;
wire n_17451;
wire n_17452;
wire n_17453;
wire n_17454;
wire n_17455;
wire n_17456;
wire n_17457;
wire n_17458;
wire n_17459;
wire n_17460;
wire n_17461;
wire n_17462;
wire n_17463;
wire n_17464;
wire n_17465;
wire n_17466;
wire n_17467;
wire n_17468;
wire n_17469;
wire n_17470;
wire n_17471;
wire n_17472;
wire n_17473;
wire n_17474;
wire n_17475;
wire n_17476;
wire n_17477;
wire n_17478;
wire n_17479;
wire n_17480;
wire n_17481;
wire n_17482;
wire n_17483;
wire n_17484;
wire n_17485;
wire n_17486;
wire n_17487;
wire n_17488;
wire n_17489;
wire n_17490;
wire n_17491;
wire n_17492;
wire n_17493;
wire n_17494;
wire n_17495;
wire n_17496;
wire n_17497;
wire n_17498;
wire n_17499;
wire n_17500;
wire n_17501;
wire n_17502;
wire n_17503;
wire n_17504;
wire n_17505;
wire n_17506;
wire n_17507;
wire n_17508;
wire n_17509;
wire n_17510;
wire n_17511;
wire n_17512;
wire n_17513;
wire n_17514;
wire n_17515;
wire n_17516;
wire n_17517;
wire n_17518;
wire n_17519;
wire n_17520;
wire n_17521;
wire n_17522;
wire n_17523;
wire n_17524;
wire n_17525;
wire n_17526;
wire n_17527;
wire n_17528;
wire n_17529;
wire n_17530;
wire n_17531;
wire n_17532;
wire n_17533;
wire n_17534;
wire n_17535;
wire n_17536;
wire n_17537;
wire n_17538;
wire n_17539;
wire n_17540;
wire n_17541;
wire n_17542;
wire n_17543;
wire n_17544;
wire n_17545;
wire n_17546;
wire n_17547;
wire n_17548;
wire n_17549;
wire n_17550;
wire n_17551;
wire n_17552;
wire n_17553;
wire n_17554;
wire n_17555;
wire n_17556;
wire n_17557;
wire n_17558;
wire n_17559;
wire n_17560;
wire n_17561;
wire n_17562;
wire n_17563;
wire n_17564;
wire n_17565;
wire n_17566;
wire n_17567;
wire n_17568;
wire n_17569;
wire n_17570;
wire n_17571;
wire n_17572;
wire n_17573;
wire n_17574;
wire n_17575;
wire n_17576;
wire n_17577;
wire n_17578;
wire n_17579;
wire n_17580;
wire n_17581;
wire n_17582;
wire n_17583;
wire n_17584;
wire n_17585;
wire n_17586;
wire n_17587;
wire n_17588;
wire n_17589;
wire n_17590;
wire n_17591;
wire n_17592;
wire n_17593;
wire n_17594;
wire n_17595;
wire n_17596;
wire n_17597;
wire n_17598;
wire n_17599;
wire n_17600;
wire n_17601;
wire n_17602;
wire n_17603;
wire n_17604;
wire n_17605;
wire n_17606;
wire n_17607;
wire n_17608;
wire n_17609;
wire n_17610;
wire n_17611;
wire n_17612;
wire n_17613;
wire n_17614;
wire n_17615;
wire n_17616;
wire n_17617;
wire n_17618;
wire n_17619;
wire n_17620;
wire n_17621;
wire n_17622;
wire n_17623;
wire n_17624;
wire n_17625;
wire n_17626;
wire n_17627;
wire n_17628;
wire n_17629;
wire n_17630;
wire n_17631;
wire n_17632;
wire n_17633;
wire n_17634;
wire n_17635;
wire n_17636;
wire n_17637;
wire n_17638;
wire n_17639;
wire n_17640;
wire n_17641;
wire n_17642;
wire n_17643;
wire n_17644;
wire n_17645;
wire n_17646;
wire n_17647;
wire n_17648;
wire n_17649;
wire n_17650;
wire n_17651;
wire n_17652;
wire n_17653;
wire n_17654;
wire n_17655;
wire n_17656;
wire n_17657;
wire n_17658;
wire n_17659;
wire n_17660;
wire n_17661;
wire n_17662;
wire n_17663;
wire n_17664;
wire n_17665;
wire n_17666;
wire n_17667;
wire n_17668;
wire n_17669;
wire n_17670;
wire n_17671;
wire n_17672;
wire n_17673;
wire n_17674;
wire n_17675;
wire n_17676;
wire n_17677;
wire n_17678;
wire n_17679;
wire n_17680;
wire n_17681;
wire n_17682;
wire n_17683;
wire n_17684;
wire n_17685;
wire n_17686;
wire n_17687;
wire n_17688;
wire n_17689;
wire n_17690;
wire n_17691;
wire n_17692;
wire n_17693;
wire n_17694;
wire n_17695;
wire n_17696;
wire n_17697;
wire n_17698;
wire n_17699;
wire n_17700;
wire n_17701;
wire n_17702;
wire n_17703;
wire n_17704;
wire n_17705;
wire n_17706;
wire n_17707;
wire n_17708;
wire n_17709;
wire n_17710;
wire n_17711;
wire n_17712;
wire n_17713;
wire n_17714;
wire n_17715;
wire n_17716;
wire n_17717;
wire n_17718;
wire n_17719;
wire n_17720;
wire n_17721;
wire n_17722;
wire n_17723;
wire n_17724;
wire n_17725;
wire n_17726;
wire n_17727;
wire n_17728;
wire n_17729;
wire n_17730;
wire n_17731;
wire n_17732;
wire n_17733;
wire n_17734;
wire n_17735;
wire n_17736;
wire n_17737;
wire n_17738;
wire n_17739;
wire n_17740;
wire n_17741;
wire n_17742;
wire n_17743;
wire n_17744;
wire n_17745;
wire n_17746;
wire n_17747;
wire n_17748;
wire n_17749;
wire n_17750;
wire n_17751;
wire n_17752;
wire n_17753;
wire n_17754;
wire n_17755;
wire n_17756;
wire n_17757;
wire n_17758;
wire n_17759;
wire n_17760;
wire n_17761;
wire n_17762;
wire n_17763;
wire n_17764;
wire n_17765;
wire n_17766;
wire n_17767;
wire n_17768;
wire n_17769;
wire n_17770;
wire n_17771;
wire n_17772;
wire n_17773;
wire n_17774;
wire n_17775;
wire n_17776;
wire n_17777;
wire n_17778;
wire n_17779;
wire n_17780;
wire n_17781;
wire n_17782;
wire n_17783;
wire n_17784;
wire n_17785;
wire n_17786;
wire n_17787;
wire n_17788;
wire n_17789;
wire n_17790;
wire n_17791;
wire n_17792;
wire n_17793;
wire n_17794;
wire n_17795;
wire n_17796;
wire n_17797;
wire n_17798;
wire n_17799;
wire n_17800;
wire n_17801;
wire n_17802;
wire n_17803;
wire n_17804;
wire n_17805;
wire n_17806;
wire n_17807;
wire n_17808;
wire n_17809;
wire n_17810;
wire n_17811;
wire n_17812;
wire n_17813;
wire n_17814;
wire n_17815;
wire n_17816;
wire n_17817;
wire n_17818;
wire n_17819;
wire n_17820;
wire n_17821;
wire n_17822;
wire n_17823;
wire n_17824;
wire n_17825;
wire n_17826;
wire n_17827;
wire n_17828;
wire n_17829;
wire n_17830;
wire n_17831;
wire n_17832;
wire n_17833;
wire n_17834;
wire n_17835;
wire n_17836;
wire n_17837;
wire n_17838;
wire n_17839;
wire n_17840;
wire n_17841;
wire n_17842;
wire n_17843;
wire n_17844;
wire n_17845;
wire n_17846;
wire n_17847;
wire n_17848;
wire n_17849;
wire n_17850;
wire n_17851;
wire n_17852;
wire n_17853;
wire n_17854;
wire n_17855;
wire n_17856;
wire n_17857;
wire n_17858;
wire n_17859;
wire n_17860;
wire n_17861;
wire n_17862;
wire n_17863;
wire n_17864;
wire n_17865;
wire n_17866;
wire n_17867;
wire n_17868;
wire n_17869;
wire n_17870;
wire n_17871;
wire n_17872;
wire n_17873;
wire n_17874;
wire n_17875;
wire n_17876;
wire n_17877;
wire n_17878;
wire n_17879;
wire n_17880;
wire n_17881;
wire n_17882;
wire n_17883;
wire n_17884;
wire n_17885;
wire n_17886;
wire n_17887;
wire n_17888;
wire n_17889;
wire n_17890;
wire n_17891;
wire n_17892;
wire n_17893;
wire n_17894;
wire n_17895;
wire n_17896;
wire n_17897;
wire n_17898;
wire n_17899;
wire n_17900;
wire n_17901;
wire n_17902;
wire n_17903;
wire n_17904;
wire n_17905;
wire n_17906;
wire n_17907;
wire n_17908;
wire n_17909;
wire n_17910;
wire n_17911;
wire n_17912;
wire n_17913;
wire n_17914;
wire n_17915;
wire n_17916;
wire n_17917;
wire n_17918;
wire n_17919;
wire n_17920;
wire n_17921;
wire n_17922;
wire n_17923;
wire n_17924;
wire n_17925;
wire n_17926;
wire n_17927;
wire n_17928;
wire n_17929;
wire n_17930;
wire n_17931;
wire n_17932;
wire n_17933;
wire n_17934;
wire n_17935;
wire n_17936;
wire n_17937;
wire n_17938;
wire n_17939;
wire n_17940;
wire n_17941;
wire n_17942;
wire n_17943;
wire n_17944;
wire n_17945;
wire n_17946;
wire n_17947;
wire n_17948;
wire n_17949;
wire n_17950;
wire n_17951;
wire n_17952;
wire n_17953;
wire n_17954;
wire n_17955;
wire n_17956;
wire n_17957;
wire n_17958;
wire n_17959;
wire n_17960;
wire n_17961;
wire n_17962;
wire n_17963;
wire n_17964;
wire n_17965;
wire n_17966;
wire n_17967;
wire n_17968;
wire n_17969;
wire n_17970;
wire n_17971;
wire n_17972;
wire n_17973;
wire n_17974;
wire n_17975;
wire n_17976;
wire n_17977;
wire n_17978;
wire n_17979;
wire n_17980;
wire n_17981;
wire n_17982;
wire n_17983;
wire n_17984;
wire n_17985;
wire n_17986;
wire n_17987;
wire n_17988;
wire n_17989;
wire n_17990;
wire n_17991;
wire n_17992;
wire n_17993;
wire n_17994;
wire n_17995;
wire n_17996;
wire n_17997;
wire n_17998;
wire n_17999;
wire n_18000;
wire n_18001;
wire n_18002;
wire n_18003;
wire n_18004;
wire n_18005;
wire n_18006;
wire n_18007;
wire n_18008;
wire n_18009;
wire n_18010;
wire n_18011;
wire n_18012;
wire n_18013;
wire n_18014;
wire n_18015;
wire n_18016;
wire n_18017;
wire n_18018;
wire n_18019;
wire n_18020;
wire n_18021;
wire n_18022;
wire n_18023;
wire n_18024;
wire n_18025;
wire n_18026;
wire n_18027;
wire n_18028;
wire n_18029;
wire n_18030;
wire n_18031;
wire n_18032;
wire n_18033;
wire n_18034;
wire n_18035;
wire n_18036;
wire n_18037;
wire n_18038;
wire n_18039;
wire n_18040;
wire n_18041;
wire n_18042;
wire n_18043;
wire n_18044;
wire n_18045;
wire n_18046;
wire n_18047;
wire n_18048;
wire n_18049;
wire n_18050;
wire n_18051;
wire n_18052;
wire n_18053;
wire n_18054;
wire n_18055;
wire n_18056;
wire n_18057;
wire n_18058;
wire n_18059;
wire n_18060;
wire n_18061;
wire n_18062;
wire n_18063;
wire n_18064;
wire n_18065;
wire n_18066;
wire n_18067;
wire n_18068;
wire n_18069;
wire n_18070;
wire n_18071;
wire n_18072;
wire n_18073;
wire n_18074;
wire n_18075;
wire n_18076;
wire n_18077;
wire n_18078;
wire n_18079;
wire n_18080;
wire n_18081;
wire n_18082;
wire n_18083;
wire n_18084;
wire n_18085;
wire n_18086;
wire n_18087;
wire n_18088;
wire n_18089;
wire n_18090;
wire n_18091;
wire n_18092;
wire n_18093;
wire n_18094;
wire n_18095;
wire n_18096;
wire n_18097;
wire n_18098;
wire n_18099;
wire n_18100;
wire n_18101;
wire n_18102;
wire n_18103;
wire n_18104;
wire n_18105;
wire n_18106;
wire n_18107;
wire n_18108;
wire n_18109;
wire n_18110;
wire n_18111;
wire n_18112;
wire n_18113;
wire n_18114;
wire n_18115;
wire n_18116;
wire n_18117;
wire n_18118;
wire n_18119;
wire n_18120;
wire n_18121;
wire n_18122;
wire n_18123;
wire n_18124;
wire n_18125;
wire n_18126;
wire n_18127;
wire n_18128;
wire n_18129;
wire n_18130;
wire n_18131;
wire n_18132;
wire n_18133;
wire n_18134;
wire n_18135;
wire n_18136;
wire n_18137;
wire n_18138;
wire n_18139;
wire n_18140;
wire n_18141;
wire n_18142;
wire n_18143;
wire n_18144;
wire n_18145;
wire n_18146;
wire n_18147;
wire n_18148;
wire n_18149;
wire n_18150;
wire n_18151;
wire n_18152;
wire n_18153;
wire n_18154;
wire n_18155;
wire n_18156;
wire n_18157;
wire n_18158;
wire n_18159;
wire n_18160;
wire n_18161;
wire n_18162;
wire n_18163;
wire n_18164;
wire n_18165;
wire n_18166;
wire n_18167;
wire n_18168;
wire n_18169;
wire n_18170;
wire n_18171;
wire n_18172;
wire n_18173;
wire n_18174;
wire n_18175;
wire n_18176;
wire n_18177;
wire n_18178;
wire n_18179;
wire n_18180;
wire n_18181;
wire n_18182;
wire n_18183;
wire n_18184;
wire n_18185;
wire n_18186;
wire n_18187;
wire n_18188;
wire n_18189;
wire n_18190;
wire n_18191;
wire n_18192;
wire n_18193;
wire n_18194;
wire n_18195;
wire n_18196;
wire n_18197;
wire n_18198;
wire n_18199;
wire n_18200;
wire n_18201;
wire n_18202;
wire n_18203;
wire n_18204;
wire n_18205;
wire n_18206;
wire n_18207;
wire n_18208;
wire n_18209;
wire n_18210;
wire n_18211;
wire n_18212;
wire n_18213;
wire n_18214;
wire n_18215;
wire n_18216;
wire n_18217;
wire n_18218;
wire n_18219;
wire n_18220;
wire n_18221;
wire n_18222;
wire n_18223;
wire n_18224;
wire n_18225;
wire n_18226;
wire n_18227;
wire n_18228;
wire n_18229;
wire n_18230;
wire n_18231;
wire n_18232;
wire n_18233;
wire n_18234;
wire n_18235;
wire n_18236;
wire n_18237;
wire n_18238;
wire n_18239;
wire n_18240;
wire n_18241;
wire n_18242;
wire n_18243;
wire n_18244;
wire n_18245;
wire n_18246;
wire n_18247;
wire n_18248;
wire n_18249;
wire n_18250;
wire n_18251;
wire n_18252;
wire n_18253;
wire n_18254;
wire n_18255;
wire n_18256;
wire n_18257;
wire n_18258;
wire n_18259;
wire n_18260;
wire n_18261;
wire n_18262;
wire n_18263;
wire n_18264;
wire n_18265;
wire n_18266;
wire n_18267;
wire n_18268;
wire n_18269;
wire n_18270;
wire n_18271;
wire n_18272;
wire n_18273;
wire n_18274;
wire n_18275;
wire n_18276;
wire n_18277;
wire n_18278;
wire n_18279;
wire n_18280;
wire n_18281;
wire n_18282;
wire n_18283;
wire n_18284;
wire n_18285;
wire n_18286;
wire n_18287;
wire n_18288;
wire n_18289;
wire n_18290;
wire n_18291;
wire n_18292;
wire n_18293;
wire n_18294;
wire n_18295;
wire n_18296;
wire n_18297;
wire n_18298;
wire n_18299;
wire n_18300;
wire n_18301;
wire n_18302;
wire n_18303;
wire n_18304;
wire n_18305;
wire n_18306;
wire n_18307;
wire n_18308;
wire n_18309;
wire n_18310;
wire n_18311;
wire n_18312;
wire n_18313;
wire n_18314;
wire n_18315;
wire n_18316;
wire n_18317;
wire n_18318;
wire n_18319;
wire n_18320;
wire n_18321;
wire n_18322;
wire n_18323;
wire n_18324;
wire n_18325;
wire n_18326;
wire n_18327;
wire n_18328;
wire n_18329;
wire n_18330;
wire n_18331;
wire n_18332;
wire n_18333;
wire n_18334;
wire n_18335;
wire n_18336;
wire n_18337;
wire n_18338;
wire n_18339;
wire n_18340;
wire n_18341;
wire n_18342;
wire n_18343;
wire n_18344;
wire n_18345;
wire n_18346;
wire n_18347;
wire n_18348;
wire n_18349;
wire n_18350;
wire n_18351;
wire n_18352;
wire n_18353;
wire n_18354;
wire n_18355;
wire n_18356;
wire n_18357;
wire n_18358;
wire n_18359;
wire n_18360;
wire n_18361;
wire n_18362;
wire n_18363;
wire n_18364;
wire n_18365;
wire n_18366;
wire n_18367;
wire n_18368;
wire n_18369;
wire n_18370;
wire n_18371;
wire n_18372;
wire n_18373;
wire n_18374;
wire n_18375;
wire n_18376;
wire n_18377;
wire n_18378;
wire n_18379;
wire n_18380;
wire n_18381;
wire n_18382;
wire n_18383;
wire n_18384;
wire n_18385;
wire n_18386;
wire n_18387;
wire n_18388;
wire n_18389;
wire n_18390;
wire n_18391;
wire n_18392;
wire n_18393;
wire n_18394;
wire n_18395;
wire n_18396;
wire n_18397;
wire n_18398;
wire n_18399;
wire n_18400;
wire n_18401;
wire n_18402;
wire n_18403;
wire n_18404;
wire n_18405;
wire n_18406;
wire n_18407;
wire n_18408;
wire n_18409;
wire n_18410;
wire n_18411;
wire n_18412;
wire n_18413;
wire n_18414;
wire n_18415;
wire n_18416;
wire n_18417;
wire n_18418;
wire n_18419;
wire n_18420;
wire n_18421;
wire n_18422;
wire n_18423;
wire n_18424;
wire n_18425;
wire n_18426;
wire n_18427;
wire n_18428;
wire n_18429;
wire n_18430;
wire n_18431;
wire n_18432;
wire n_18433;
wire n_18434;
wire n_18435;
wire n_18436;
wire n_18437;
wire n_18438;
wire n_18439;
wire n_18440;
wire n_18441;
wire n_18442;
wire n_18443;
wire n_18444;
wire n_18445;
wire n_18446;
wire n_18447;
wire n_18448;
wire n_18449;
wire n_18450;
wire n_18451;
wire n_18452;
wire n_18453;
wire n_18454;
wire n_18455;
wire n_18456;
wire n_18457;
wire n_18458;
wire n_18459;
wire n_18460;
wire n_18461;
wire n_18462;
wire n_18463;
wire n_18464;
wire n_18465;
wire n_18466;
wire n_18467;
wire n_18468;
wire n_18469;
wire n_18470;
wire n_18471;
wire n_18472;
wire n_18473;
wire n_18474;
wire n_18475;
wire n_18476;
wire n_18477;
wire n_18478;
wire n_18479;
wire n_18480;
wire n_18481;
wire n_18482;
wire n_18483;
wire n_18484;
wire n_18485;
wire n_18486;
wire n_18487;
wire n_18488;
wire n_18489;
wire n_18490;
wire n_18491;
wire n_18492;
wire n_18493;
wire n_18494;
wire n_18495;
wire n_18496;
wire n_18497;
wire n_18498;
wire n_18499;
wire n_18500;
wire n_18501;
wire n_18502;
wire n_18503;
wire n_18504;
wire n_18505;
wire n_18506;
wire n_18507;
wire n_18508;
wire n_18509;
wire n_18510;
wire n_18511;
wire n_18512;
wire n_18513;
wire n_18514;
wire n_18515;
wire n_18516;
wire n_18517;
wire n_18518;
wire n_18519;
wire n_18520;
wire n_18521;
wire n_18522;
wire n_18523;
wire n_18524;
wire n_18525;
wire n_18526;
wire n_18527;
wire n_18528;
wire n_18529;
wire n_18530;
wire n_18531;
wire n_18532;
wire n_18533;
wire n_18534;
wire n_18535;
wire n_18536;
wire n_18537;
wire n_18538;
wire n_18539;
wire n_18540;
wire n_18541;
wire n_18542;
wire n_18543;
wire n_18544;
wire n_18545;
wire n_18546;
wire n_18547;
wire n_18548;
wire n_18549;
wire n_18550;
wire n_18551;
wire n_18552;
wire n_18553;
wire n_18554;
wire n_18555;
wire n_18556;
wire n_18557;
wire n_18558;
wire n_18559;
wire n_18560;
wire n_18561;
wire n_18562;
wire n_18563;
wire n_18564;
wire n_18565;
wire n_18566;
wire n_18567;
wire n_18568;
wire n_18569;
wire n_18570;
wire n_18571;
wire n_18572;
wire n_18573;
wire n_18574;
wire n_18575;
wire n_18576;
wire n_18577;
wire n_18578;
wire n_18579;
wire n_18580;
wire n_18581;
wire n_18582;
wire n_18583;
wire n_18584;
wire n_18585;
wire n_18586;
wire n_18587;
wire n_18588;
wire n_18589;
wire n_18590;
wire n_18591;
wire n_18592;
wire n_18593;
wire n_18594;
wire n_18595;
wire n_18596;
wire n_18597;
wire n_18598;
wire n_18599;
wire n_18600;
wire n_18601;
wire n_18602;
wire n_18603;
wire n_18604;
wire n_18605;
wire n_18606;
wire n_18607;
wire n_18608;
wire n_18609;
wire n_18610;
wire n_18611;
wire n_18612;
wire n_18613;
wire n_18614;
wire n_18615;
wire n_18616;
wire n_18617;
wire n_18618;
wire n_18619;
wire n_18620;
wire n_18621;
wire n_18622;
wire n_18623;
wire n_18624;
wire n_18625;
wire n_18626;
wire n_18627;
wire n_18628;
wire n_18629;
wire n_18630;
wire n_18631;
wire n_18632;
wire n_18633;
wire n_18634;
wire n_18635;
wire n_18636;
wire n_18637;
wire n_18638;
wire n_18639;
wire n_18640;
wire n_18641;
wire n_18642;
wire n_18643;
wire n_18644;
wire n_18645;
wire n_18646;
wire n_18647;
wire n_18648;
wire n_18649;
wire n_18650;
wire n_18651;
wire n_18652;
wire n_18653;
wire n_18654;
wire n_18655;
wire n_18656;
wire n_18657;
wire n_18658;
wire n_18659;
wire n_18660;
wire n_18661;
wire n_18662;
wire n_18663;
wire n_18664;
wire n_18665;
wire n_18666;
wire n_18667;
wire n_18668;
wire n_18669;
wire n_18670;
wire n_18671;
wire n_18672;
wire n_18673;
wire n_18674;
wire n_18675;
wire n_18676;
wire n_18677;
wire n_18678;
wire n_18679;
wire n_18680;
wire n_18681;
wire n_18682;
wire n_18683;
wire n_18684;
wire n_18685;
wire n_18686;
wire n_18687;
wire n_18688;
wire n_18689;
wire n_18690;
wire n_18691;
wire n_18692;
wire n_18693;
wire n_18694;
wire n_18695;
wire n_18696;
wire n_18697;
wire n_18698;
wire n_18699;
wire n_18700;
wire n_18701;
wire n_18702;
wire n_18703;
wire n_18704;
wire n_18705;
wire n_18706;
wire n_18707;
wire n_18708;
wire n_18709;
wire n_18710;
wire n_18711;
wire n_18712;
wire n_18713;
wire n_18714;
wire n_18715;
wire n_18716;
wire n_18717;
wire n_18718;
wire n_18719;
wire n_18720;
wire n_18721;
wire n_18722;
wire n_18723;
wire n_18724;
wire n_18725;
wire n_18726;
wire n_18727;
wire n_18728;
wire n_18729;
wire n_18730;
wire n_18731;
wire n_18732;
wire n_18733;
wire n_18734;
wire n_18735;
wire n_18736;
wire n_18737;
wire n_18738;
wire n_18739;
wire n_18740;
wire n_18741;
wire n_18742;
wire n_18743;
wire n_18744;
wire n_18745;
wire n_18746;
wire n_18747;
wire n_18748;
wire n_18749;
wire n_18750;
wire n_18751;
wire n_18752;
wire n_18753;
wire n_18754;
wire n_18755;
wire n_18756;
wire n_18757;
wire n_18758;
wire n_18759;
wire n_18760;
wire n_18761;
wire n_18762;
wire n_18763;
wire n_18764;
wire n_18765;
wire n_18766;
wire n_18767;
wire n_18768;
wire n_18769;
wire n_18770;
wire n_18771;
wire n_18772;
wire n_18773;
wire n_18774;
wire n_18775;
wire n_18776;
wire n_18777;
wire n_18778;
wire n_18779;
wire n_18780;
wire n_18781;
wire n_18782;
wire n_18783;
wire n_18784;
wire n_18785;
wire n_18786;
wire n_18787;
wire n_18788;
wire n_18789;
wire n_18790;
wire n_18791;
wire n_18792;
wire n_18793;
wire n_18794;
wire n_18795;
wire n_18796;
wire n_18797;
wire n_18798;
wire n_18799;
wire n_18800;
wire n_18801;
wire n_18802;
wire n_18803;
wire n_18804;
wire n_18805;
wire n_18806;
wire n_18807;
wire n_18808;
wire n_18809;
wire n_18810;
wire n_18811;
wire n_18812;
wire n_18813;
wire n_18814;
wire n_18815;
wire n_18816;
wire n_18817;
wire n_18818;
wire n_18819;
wire n_18820;
wire n_18821;
wire n_18822;
wire n_18823;
wire n_18824;
wire n_18825;
wire n_18826;
wire n_18827;
wire n_18828;
wire n_18829;
wire n_18830;
wire n_18831;
wire n_18832;
wire n_18833;
wire n_18834;
wire n_18835;
wire n_18836;
wire n_18837;
wire n_18838;
wire n_18839;
wire n_18840;
wire n_18841;
wire n_18842;
wire n_18843;
wire n_18844;
wire n_18845;
wire n_18846;
wire n_18847;
wire n_18848;
wire n_18849;
wire n_18850;
wire n_18851;
wire n_18852;
wire n_18853;
wire n_18854;
wire n_18855;
wire n_18856;
wire n_18857;
wire n_18858;
wire n_18859;
wire n_18860;
wire n_18861;
wire n_18862;
wire n_18863;
wire n_18864;
wire n_18865;
wire n_18866;
wire n_18867;
wire n_18868;
wire n_18869;
wire n_18870;
wire n_18871;
wire n_18872;
wire n_18873;
wire n_18874;
wire n_18875;
wire n_18876;
wire n_18877;
wire n_18878;
wire n_18879;
wire n_18880;
wire n_18881;
wire n_18882;
wire n_18883;
wire n_18884;
wire n_18885;
wire n_18886;
wire n_18887;
wire n_18888;
wire n_18889;
wire n_18890;
wire n_18891;
wire n_18892;
wire n_18893;
wire n_18894;
wire n_18895;
wire n_18896;
wire n_18897;
wire n_18898;
wire n_18899;
wire n_18900;
wire n_18901;
wire n_18902;
wire n_18903;
wire n_18904;
wire n_18905;
wire n_18906;
wire n_18907;
wire n_18908;
wire n_18909;
wire n_18910;
wire n_18911;
wire n_18912;
wire n_18913;
wire n_18914;
wire n_18915;
wire n_18916;
wire n_18917;
wire n_18918;
wire n_18919;
wire n_18920;
wire n_18921;
wire n_18922;
wire n_18923;
wire n_18924;
wire n_18925;
wire n_18926;
wire n_18927;
wire n_18928;
wire n_18929;
wire n_18930;
wire n_18931;
wire n_18932;
wire n_18933;
wire n_18934;
wire n_18935;
wire n_18936;
wire n_18937;
wire n_18938;
wire n_18939;
wire n_18940;
wire n_18941;
wire n_18942;
wire n_18943;
wire n_18944;
wire n_18945;
wire n_18946;
wire n_18947;
wire n_18948;
wire n_18949;
wire n_18950;
wire n_18951;
wire n_18952;
wire n_18953;
wire n_18954;
wire n_18955;
wire n_18956;
wire n_18957;
wire n_18958;
wire n_18959;
wire n_18960;
wire n_18961;
wire n_18962;
wire n_18963;
wire n_18964;
wire n_18965;
wire n_18966;
wire n_18967;
wire n_18968;
wire n_18969;
wire n_18970;
wire n_18971;
wire n_18972;
wire n_18973;
wire n_18974;
wire n_18975;
wire n_18976;
wire n_18977;
wire n_18978;
wire n_18979;
wire n_18980;
wire n_18981;
wire n_18982;
wire n_18983;
wire n_18984;
wire n_18985;
wire n_18986;
wire n_18987;
wire n_18988;
wire n_18989;
wire n_18990;
wire n_18991;
wire n_18992;
wire n_18993;
wire n_18994;
wire n_18995;
wire n_18996;
wire n_18997;
wire n_18998;
wire n_18999;
wire n_19000;
wire n_19001;
wire n_19002;
wire n_19003;
wire n_19004;
wire n_19005;
wire n_19006;
wire n_19007;
wire n_19008;
wire n_19009;
wire n_19010;
wire n_19011;
wire n_19012;
wire n_19013;
wire n_19014;
wire n_19015;
wire n_19016;
wire n_19017;
wire n_19018;
wire n_19019;
wire n_19020;
wire n_19021;
wire n_19022;
wire n_19023;
wire n_19024;
wire n_19025;
wire n_19026;
wire n_19027;
wire n_19028;
wire n_19029;
wire n_19030;
wire n_19031;
wire n_19032;
wire n_19033;
wire n_19034;
wire n_19035;
wire n_19036;
wire n_19037;
wire n_19038;
wire n_19039;
wire n_19040;
wire n_19041;
wire n_19042;
wire n_19043;
wire n_19044;
wire n_19045;
wire n_19046;
wire n_19047;
wire n_19048;
wire n_19049;
wire n_19050;
wire n_19051;
wire n_19052;
wire n_19053;
wire n_19054;
wire n_19055;
wire n_19056;
wire n_19057;
wire n_19058;
wire n_19059;
wire n_19060;
wire n_19061;
wire n_19062;
wire n_19063;
wire n_19064;
wire n_19065;
wire n_19066;
wire n_19067;
wire n_19068;
wire n_19069;
wire n_19070;
wire n_19071;
wire n_19072;
wire n_19073;
wire n_19074;
wire n_19075;
wire n_19076;
wire n_19077;
wire n_19078;
wire n_19079;
wire n_19080;
wire n_19081;
wire n_19082;
wire n_19083;
wire n_19084;
wire n_19085;
wire n_19086;
wire n_19087;
wire n_19088;
wire n_19089;
wire n_19090;
wire n_19091;
wire n_19092;
wire n_19093;
wire n_19094;
wire n_19095;
wire n_19096;
wire n_19097;
wire n_19098;
wire n_19099;
wire n_19100;
wire n_19101;
wire n_19102;
wire n_19103;
wire n_19104;
wire n_19105;
wire n_19106;
wire n_19107;
wire n_19108;
wire n_19109;
wire n_19110;
wire n_19111;
wire n_19112;
wire n_19113;
wire n_19114;
wire n_19115;
wire n_19116;
wire n_19117;
wire n_19118;
wire n_19119;
wire n_19120;
wire n_19121;
wire n_19122;
wire n_19123;
wire n_19124;
wire n_19125;
wire n_19126;
wire n_19127;
wire n_19128;
wire n_19129;
wire n_19130;
wire n_19131;
wire n_19132;
wire n_19133;
wire n_19134;
wire n_19135;
wire n_19136;
wire n_19137;
wire n_19138;
wire n_19139;
wire n_19140;
wire n_19141;
wire n_19142;
wire n_19143;
wire n_19144;
wire n_19145;
wire n_19146;
wire n_19147;
wire n_19148;
wire n_19149;
wire n_19150;
wire n_19151;
wire n_19152;
wire n_19153;
wire n_19154;
wire n_19155;
wire n_19156;
wire n_19157;
wire n_19158;
wire n_19159;
wire n_19160;
wire n_19161;
wire n_19162;
wire n_19163;
wire n_19164;
wire n_19165;
wire n_19166;
wire n_19167;
wire n_19168;
wire n_19169;
wire n_19170;
wire n_19171;
wire n_19172;
wire n_19173;
wire n_19174;
wire n_19175;
wire n_19176;
wire n_19177;
wire n_19178;
wire n_19179;
wire n_19180;
wire n_19181;
wire n_19182;
wire n_19183;
wire n_19184;
wire n_19185;
wire n_19186;
wire n_19187;
wire n_19188;
wire n_19189;
wire n_19190;
wire n_19191;
wire n_19192;
wire n_19193;
wire n_19194;
wire n_19195;
wire n_19196;
wire n_19197;
wire n_19198;
wire n_19199;
wire n_19200;
wire n_19201;
wire n_19202;
wire n_19203;
wire n_19204;
wire n_19205;
wire n_19206;
wire n_19207;
wire n_19208;
wire n_19209;
wire n_19210;
wire n_19211;
wire n_19212;
wire n_19213;
wire n_19214;
wire n_19215;
wire n_19216;
wire n_19217;
wire n_19218;
wire n_19219;
wire n_19220;
wire n_19221;
wire n_19222;
wire n_19223;
wire n_19224;
wire n_19225;
wire n_19226;
wire n_19227;
wire n_19228;
wire n_19229;
wire n_19230;
wire n_19231;
wire n_19232;
wire n_19233;
wire n_19234;
wire n_19235;
wire n_19236;
wire n_19237;
wire n_19238;
wire n_19239;
wire n_19240;
wire n_19241;
wire n_19242;
wire n_19243;
wire n_19244;
wire n_19245;
wire n_19246;
wire n_19247;
wire n_19248;
wire n_19249;
wire n_19250;
wire n_19251;
wire n_19252;
wire n_19253;
wire n_19254;
wire n_19255;
wire n_19256;
wire n_19257;
wire n_19258;
wire n_19259;
wire n_19260;
wire n_19261;
wire n_19262;
wire n_19263;
wire n_19264;
wire n_19265;
wire n_19266;
wire n_19267;
wire n_19268;
wire n_19269;
wire n_19270;
wire n_19271;
wire n_19272;
wire n_19273;
wire n_19274;
wire n_19275;
wire n_19276;
wire n_19277;
wire n_19278;
wire n_19279;
wire n_19280;
wire n_19281;
wire n_19282;
wire n_19283;
wire n_19284;
wire n_19285;
wire n_19286;
wire n_19287;
wire n_19288;
wire n_19289;
wire n_19290;
wire n_19291;
wire n_19292;
wire n_19293;
wire n_19294;
wire n_19295;
wire n_19296;
wire n_19297;
wire n_19298;
wire n_19299;
wire n_19300;
wire n_19301;
wire n_19302;
wire n_19303;
wire n_19304;
wire n_19305;
wire n_19306;
wire n_19307;
wire n_19308;
wire n_19309;
wire n_19310;
wire n_19311;
wire n_19312;
wire n_19313;
wire n_19314;
wire n_19315;
wire n_19316;
wire n_19317;
wire n_19318;
wire n_19319;
wire n_19320;
wire n_19321;
wire n_19322;
wire n_19323;
wire n_19324;
wire n_19325;
wire n_19326;
wire n_19327;
wire n_19328;
wire n_19329;
wire n_19330;
wire n_19331;
wire n_19332;
wire n_19333;
wire n_19334;
wire n_19335;
wire n_19336;
wire n_19337;
wire n_19338;
wire n_19339;
wire n_19340;
wire n_19341;
wire n_19342;
wire n_19343;
wire n_19344;
wire n_19345;
wire n_19346;
wire n_19347;
wire n_19348;
wire n_19349;
wire n_19350;
wire n_19351;
wire n_19352;
wire n_19353;
wire n_19354;
wire n_19355;
wire n_19356;
wire n_19357;
wire n_19358;
wire n_19359;
wire n_19360;
wire n_19361;
wire n_19362;
wire n_19363;
wire n_19364;
wire n_19365;
wire n_19366;
wire n_19367;
wire n_19368;
wire n_19369;
wire n_19370;
wire n_19371;
wire n_19372;
wire n_19373;
wire n_19374;
wire n_19375;
wire n_19376;
wire n_19377;
wire n_19378;
wire n_19379;
wire n_19380;
wire n_19381;
wire n_19382;
wire n_19383;
wire n_19384;
wire n_19385;
wire n_19386;
wire n_19387;
wire n_19388;
wire n_19389;
wire n_19390;
wire n_19391;
wire n_19392;
wire n_19393;
wire n_19394;
wire n_19395;
wire n_19396;
wire n_19397;
wire n_19398;
wire n_19399;
wire n_19400;
wire n_19401;
wire n_19402;
wire n_19403;
wire n_19404;
wire n_19405;
wire n_19406;
wire n_19407;
wire n_19408;
wire n_19409;
wire n_19410;
wire n_19411;
wire n_19412;
wire n_19413;
wire n_19414;
wire n_19415;
wire n_19416;
wire n_19417;
wire n_19418;
wire n_19419;
wire n_19420;
wire n_19421;
wire n_19422;
wire n_19423;
wire n_19424;
wire n_19425;
wire n_19426;
wire n_19427;
wire n_19428;
wire n_19429;
wire n_19430;
wire n_19431;
wire n_19432;
wire n_19433;
wire n_19434;
wire n_19435;
wire n_19436;
wire n_19437;
wire n_19438;
wire n_19439;
wire n_19440;
wire n_19441;
wire n_19442;
wire n_19443;
wire n_19444;
wire n_19445;
wire n_19446;
wire n_19447;
wire n_19448;
wire n_19449;
wire n_19450;
wire n_19451;
wire n_19452;
wire n_19453;
wire n_19454;
wire n_19455;
wire n_19456;
wire n_19457;
wire n_19458;
wire n_19459;
wire n_19460;
wire n_19461;
wire n_19462;
wire n_19463;
wire n_19464;
wire n_19465;
wire n_19466;
wire n_19467;
wire n_19468;
wire n_19469;
wire n_19470;
wire n_19471;
wire n_19472;
wire n_19473;
wire n_19474;
wire n_19475;
wire n_19476;
wire n_19477;
wire n_19478;
wire n_19479;
wire n_19480;
wire n_19481;
wire n_19482;
wire n_19483;
wire n_19484;
wire n_19485;
wire n_19486;
wire n_19487;
wire n_19488;
wire n_19489;
wire n_19490;
wire n_19491;
wire n_19492;
wire n_19493;
wire n_19494;
wire n_19495;
wire n_19496;
wire n_19497;
wire n_19498;
wire n_19499;
wire n_19500;
wire n_19501;
wire n_19502;
wire n_19503;
wire n_19504;
wire n_19505;
wire n_19506;
wire n_19507;
wire n_19508;
wire n_19509;
wire n_19510;
wire n_19511;
wire n_19512;
wire n_19513;
wire n_19514;
wire n_19515;
wire n_19516;
wire n_19517;
wire n_19518;
wire n_19519;
wire n_19520;
wire n_19521;
wire n_19522;
wire n_19523;
wire n_19524;
wire n_19525;
wire n_19526;
wire n_19527;
wire n_19528;
wire n_19529;
wire n_19530;
wire n_19531;
wire n_19532;
wire n_19533;
wire n_19534;
wire n_19535;
wire n_19536;
wire n_19537;
wire n_19538;
wire n_19539;
wire n_19540;
wire n_19541;
wire n_19542;
wire n_19543;
wire n_19544;
wire n_19545;
wire n_19546;
wire n_19547;
wire n_19548;
wire n_19549;
wire n_19550;
wire n_19551;
wire n_19552;
wire n_19553;
wire n_19554;
wire n_19555;
wire n_19556;
wire n_19557;
wire n_19558;
wire n_19559;
wire n_19560;
wire n_19561;
wire n_19562;
wire n_19563;
wire n_19564;
wire n_19565;
wire n_19566;
wire n_19567;
wire n_19568;
wire n_19569;
wire n_19570;
wire n_19571;
wire n_19572;
wire n_19573;
wire n_19574;
wire n_19575;
wire n_19576;
wire n_19577;
wire n_19578;
wire n_19579;
wire n_19580;
wire n_19581;
wire n_19582;
wire n_19583;
wire n_19584;
wire n_19585;
wire n_19586;
wire n_19587;
wire n_19588;
wire n_19589;
wire n_19590;
wire n_19591;
wire n_19592;
wire n_19593;
wire n_19594;
wire n_19595;
wire n_19596;
wire n_19597;
wire n_19598;
wire n_19599;
wire n_19600;
wire n_19601;
wire n_19602;
wire n_19603;
wire n_19604;
wire n_19605;
wire n_19606;
wire n_19607;
wire n_19608;
wire n_19609;
wire n_19610;
wire n_19611;
wire n_19612;
wire n_19613;
wire n_19614;
wire n_19615;
wire n_19616;
wire n_19617;
wire n_19618;
wire n_19619;
wire n_19620;
wire n_19621;
wire n_19622;
wire n_19623;
wire n_19624;
wire n_19625;
wire n_19626;
wire n_19627;
wire n_19628;
wire n_19629;
wire n_19630;
wire n_19631;
wire n_19632;
wire n_19633;
wire n_19634;
wire n_19635;
wire n_19636;
wire n_19637;
wire n_19638;
wire n_19639;
wire n_19640;
wire n_19641;
wire n_19642;
wire n_19643;
wire n_19644;
wire n_19645;
wire n_19646;
wire n_19647;
wire n_19648;
wire n_19649;
wire n_19650;
wire n_19651;
wire n_19652;
wire n_19653;
wire n_19654;
wire n_19655;
wire n_19656;
wire n_19657;
wire n_19658;
wire n_19659;
wire n_19660;
wire n_19661;
wire n_19662;
wire n_19663;
wire n_19664;
wire n_19665;
wire n_19666;
wire n_19667;
wire n_19668;
wire n_19669;
wire n_19670;
wire n_19671;
wire n_19672;
wire n_19673;
wire n_19674;
wire n_19675;
wire n_19676;
wire n_19677;
wire n_19678;
wire n_19679;
wire n_19680;
wire n_19681;
wire n_19682;
wire n_19683;
wire n_19684;
wire n_19685;
wire n_19686;
wire n_19687;
wire n_19688;
wire n_19689;
wire n_19690;
wire n_19691;
wire n_19692;
wire n_19693;
wire n_19694;
wire n_19695;
wire n_19696;
wire n_19697;
wire n_19698;
wire n_19699;
wire n_19700;
wire n_19701;
wire n_19702;
wire n_19703;
wire n_19704;
wire n_19705;
wire n_19706;
wire n_19707;
wire n_19708;
wire n_19709;
wire n_19710;
wire n_19711;
wire n_19712;
wire n_19713;
wire n_19714;
wire n_19715;
wire n_19716;
wire n_19717;
wire n_19718;
wire n_19719;
wire n_19720;
wire n_19721;
wire n_19722;
wire n_19723;
wire n_19724;
wire n_19725;
wire n_19726;
wire n_19727;
wire n_19728;
wire n_19729;
wire n_19730;
wire n_19731;
wire n_19732;
wire n_19733;
wire n_19734;
wire n_19735;
wire n_19736;
wire n_19737;
wire n_19738;
wire n_19739;
wire n_19740;
wire n_19741;
wire n_19742;
wire n_19743;
wire n_19744;
wire n_19745;
wire n_19746;
wire n_19747;
wire n_19748;
wire n_19749;
wire n_19750;
wire n_19751;
wire n_19752;
wire n_19753;
wire n_19754;
wire n_19755;
wire n_19756;
wire n_19757;
wire n_19758;
wire n_19759;
wire n_19760;
wire n_19761;
wire n_19762;
wire n_19763;
wire n_19764;
wire n_19765;
wire n_19766;
wire n_19767;
wire n_19768;
wire n_19769;
wire n_19770;
wire n_19771;
wire n_19772;
wire n_19773;
wire n_19774;
wire n_19775;
wire n_19776;
wire n_19777;
wire n_19778;
wire n_19779;
wire n_19780;
wire n_19781;
wire n_19782;
wire n_19783;
wire n_19784;
wire n_19785;
wire n_19786;
wire n_19787;
wire n_19788;
wire n_19789;
wire n_19790;
wire n_19791;
wire n_19792;
wire n_19793;
wire n_19794;
wire n_19795;
wire n_19796;
wire n_19797;
wire n_19798;
wire n_19799;
wire n_19800;
wire n_19801;
wire n_19802;
wire n_19803;
wire n_19804;
wire n_19805;
wire n_19806;
wire n_19807;
wire n_19808;
wire n_19809;
wire n_19810;
wire n_19811;
wire n_19812;
wire n_19813;
wire n_19814;
wire n_19815;
wire n_19816;
wire n_19817;
wire n_19818;
wire n_19819;
wire n_19820;
wire n_19821;
wire n_19822;
wire n_19823;
wire n_19824;
wire n_19825;
wire n_19826;
wire n_19827;
wire n_19828;
wire n_19829;
wire n_19830;
wire n_19831;
wire n_19832;
wire n_19833;
wire n_19834;
wire n_19835;
wire n_19836;
wire n_19837;
wire n_19838;
wire n_19839;
wire n_19840;
wire n_19841;
wire n_19842;
wire n_19843;
wire n_19844;
wire n_19845;
wire n_19846;
wire n_19847;
wire n_19848;
wire n_19849;
wire n_19850;
wire n_19851;
wire n_19852;
wire n_19853;
wire n_19854;
wire n_19855;
wire n_19856;
wire n_19857;
wire n_19858;
wire n_19859;
wire n_19860;
wire n_19861;
wire n_19862;
wire n_19863;
wire n_19864;
wire n_19865;
wire n_19866;
wire n_19867;
wire n_19868;
wire n_19869;
wire n_19870;
wire n_19871;
wire n_19872;
wire n_19873;
wire n_19874;
wire n_19875;
wire n_19876;
wire n_19877;
wire n_19878;
wire n_19879;
wire n_19880;
wire n_19881;
wire n_19882;
wire n_19883;
wire n_19884;
wire n_19885;
wire n_19886;
wire n_19887;
wire n_19888;
wire n_19889;
wire n_19890;
wire n_19891;
wire n_19892;
wire n_19893;
wire n_19894;
wire n_19895;
wire n_19896;
wire n_19897;
wire n_19898;
wire n_19899;
wire n_19900;
wire n_19901;
wire n_19902;
wire n_19903;
wire n_19904;
wire n_19905;
wire n_19906;
wire n_19907;
wire n_19908;
wire n_19909;
wire n_19910;
wire n_19911;
wire n_19912;
wire n_19913;
wire n_19914;
wire n_19915;
wire n_19916;
wire n_19917;
wire n_19918;
wire n_19919;
wire n_19920;
wire n_19921;
wire n_19922;
wire n_19923;
wire n_19924;
wire n_19925;
wire n_19926;
wire n_19927;
wire n_19928;
wire n_19929;
wire n_19930;
wire n_19931;
wire n_19932;
wire n_19933;
wire n_19934;
wire n_19935;
wire n_19936;
wire n_19937;
wire n_19938;
wire n_19939;
wire n_19940;
wire n_19941;
wire n_19942;
wire n_19943;
wire n_19944;
wire n_19945;
wire n_19946;
wire n_19947;
wire n_19948;
wire n_19949;
wire n_19950;
wire n_19951;
wire n_19952;
wire n_19953;
wire n_19954;
wire n_19955;
wire n_19956;
wire n_19957;
wire n_19958;
wire n_19959;
wire n_19960;
wire n_19961;
wire n_19962;
wire n_19963;
wire n_19964;
wire n_19965;
wire n_19966;
wire n_19967;
wire n_19968;
wire n_19969;
wire n_19970;
wire n_19971;
wire n_19972;
wire n_19973;
wire n_19974;
wire n_19975;
wire n_19976;
wire n_19977;
wire n_19978;
wire n_19979;
wire n_19980;
wire n_19981;
wire n_19982;
wire n_19983;
wire n_19984;
wire n_19985;
wire n_19986;
wire n_19987;
wire n_19988;
wire n_19989;
wire n_19990;
wire n_19991;
wire n_19992;
wire n_19993;
wire n_19994;
wire n_19995;
wire n_19996;
wire n_19997;
wire n_19998;
wire n_19999;
wire n_20000;
wire n_20001;
wire n_20002;
wire n_20003;
wire n_20004;
wire n_20005;
wire n_20006;
wire n_20007;
wire n_20008;
wire n_20009;
wire n_20010;
wire n_20011;
wire n_20012;
wire n_20013;
wire n_20014;
wire n_20015;
wire n_20016;
wire n_20017;
wire n_20018;
wire n_20019;
wire n_20020;
wire n_20021;
wire n_20022;
wire n_20023;
wire n_20024;
wire n_20025;
wire n_20026;
wire n_20027;
wire n_20028;
wire n_20029;
wire n_20030;
wire n_20031;
wire n_20032;
wire n_20033;
wire n_20034;
wire n_20035;
wire n_20036;
wire n_20037;
wire n_20038;
wire n_20039;
wire n_20040;
wire n_20041;
wire n_20042;
wire n_20043;
wire n_20044;
wire n_20045;
wire n_20046;
wire n_20047;
wire n_20048;
wire n_20049;
wire n_20050;
wire n_20051;
wire n_20052;
wire n_20053;
wire n_20054;
wire n_20055;
wire n_20056;
wire n_20057;
wire n_20058;
wire n_20059;
wire n_20060;
wire n_20061;
wire n_20062;
wire n_20063;
wire n_20064;
wire n_20065;
wire n_20066;
wire n_20067;
wire n_20068;
wire n_20069;
wire n_20070;
wire n_20071;
wire n_20072;
wire n_20073;
wire n_20074;
wire n_20075;
wire n_20076;
wire n_20077;
wire n_20078;
wire n_20079;
wire n_20080;
wire n_20081;
wire n_20082;
wire n_20083;
wire n_20084;
wire n_20085;
wire n_20086;
wire n_20087;
wire n_20088;
wire n_20089;
wire n_20090;
wire n_20091;
wire n_20092;
wire n_20093;
wire n_20094;
wire n_20095;
wire n_20096;
wire n_20097;
wire n_20098;
wire n_20099;
wire n_20100;
wire n_20101;
wire n_20102;
wire n_20103;
wire n_20104;
wire n_20105;
wire n_20106;
wire n_20107;
wire n_20108;
wire n_20109;
wire n_20110;
wire n_20111;
wire n_20112;
wire n_20113;
wire n_20114;
wire n_20115;
wire n_20116;
wire n_20117;
wire n_20118;
wire n_20119;
wire n_20120;
wire n_20121;
wire n_20122;
wire n_20123;
wire n_20124;
wire n_20125;
wire n_20126;
wire n_20127;
wire n_20128;
wire n_20129;
wire n_20130;
wire n_20131;
wire n_20132;
wire n_20133;
wire n_20134;
wire n_20135;
wire n_20136;
wire n_20137;
wire n_20138;
wire n_20139;
wire n_20140;
wire n_20141;
wire n_20142;
wire n_20143;
wire n_20144;
wire n_20145;
wire n_20146;
wire n_20147;
wire n_20148;
wire n_20149;
wire n_20150;
wire n_20151;
wire n_20152;
wire n_20153;
wire n_20154;
wire n_20155;
wire n_20156;
wire n_20157;
wire n_20158;
wire n_20159;
wire n_20160;
wire n_20161;
wire n_20162;
wire n_20163;
wire n_20164;
wire n_20165;
wire n_20166;
wire n_20167;
wire n_20168;
wire n_20169;
wire n_20170;
wire n_20171;
wire n_20172;
wire n_20173;
wire n_20174;
wire n_20175;
wire n_20176;
wire n_20177;
wire n_20178;
wire n_20179;
wire n_20180;
wire n_20181;
wire n_20182;
wire n_20183;
wire n_20184;
wire n_20185;
wire n_20186;
wire n_20187;
wire n_20188;
wire n_20189;
wire n_20190;
wire n_20191;
wire n_20192;
wire n_20193;
wire n_20194;
wire n_20195;
wire n_20196;
wire n_20197;
wire n_20198;
wire n_20199;
wire n_20200;
wire n_20201;
wire n_20202;
wire n_20203;
wire n_20204;
wire n_20205;
wire n_20206;
wire n_20207;
wire n_20208;
wire n_20209;
wire n_20210;
wire n_20211;
wire n_20212;
wire n_20213;
wire n_20214;
wire n_20215;
wire n_20216;
wire n_20217;
wire n_20218;
wire n_20219;
wire n_20220;
wire n_20221;
wire n_20222;
wire n_20223;
wire n_20224;
wire n_20225;
wire n_20226;
wire n_20227;
wire n_20228;
wire n_20229;
wire n_20230;
wire n_20231;
wire n_20232;
wire n_20233;
wire n_20234;
wire n_20235;
wire n_20236;
wire n_20237;
wire n_20238;
wire n_20239;
wire n_20240;
wire n_20241;
wire n_20242;
wire n_20243;
wire n_20244;
wire n_20245;
wire n_20246;
wire n_20247;
wire n_20248;
wire n_20249;
wire n_20250;
wire n_20251;
wire n_20252;
wire n_20253;
wire n_20254;
wire n_20255;
wire n_20256;
wire n_20257;
wire n_20258;
wire n_20259;
wire n_20260;
wire n_20261;
wire n_20262;
wire n_20263;
wire n_20264;
wire n_20265;
wire n_20266;
wire n_20267;
wire n_20268;
wire n_20269;
wire n_20270;
wire n_20271;
wire n_20272;
wire n_20273;
wire n_20274;
wire n_20275;
wire n_20276;
wire n_20277;
wire n_20278;
wire n_20279;
wire n_20280;
wire n_20281;
wire n_20282;
wire n_20283;
wire n_20284;
wire n_20285;
wire n_20286;
wire n_20287;
wire n_20288;
wire n_20289;
wire n_20290;
wire n_20291;
wire n_20292;
wire n_20293;
wire n_20294;
wire n_20295;
wire n_20296;
wire n_20297;
wire n_20298;
wire n_20299;
wire n_20300;
wire n_20301;
wire n_20302;
wire n_20303;
wire n_20304;
wire n_20305;
wire n_20306;
wire n_20307;
wire n_20308;
wire n_20309;
wire n_20310;
wire n_20311;
wire n_20312;
wire n_20313;
wire n_20314;
wire n_20315;
wire n_20316;
wire n_20317;
wire n_20318;
wire n_20319;
wire n_20320;
wire n_20321;
wire n_20322;
wire n_20323;
wire n_20324;
wire n_20325;
wire n_20326;
wire n_20327;
wire n_20328;
wire n_20329;
wire n_20330;
wire n_20331;
wire n_20332;
wire n_20333;
wire n_20334;
wire n_20335;
wire n_20336;
wire n_20337;
wire n_20338;
wire n_20339;
wire n_20340;
wire n_20341;
wire n_20342;
wire n_20343;
wire n_20344;
wire n_20345;
wire n_20346;
wire n_20347;
wire n_20348;
wire n_20349;
wire n_20350;
wire n_20351;
wire n_20352;
wire n_20353;
wire n_20354;
wire n_20355;
wire n_20356;
wire n_20357;
wire n_20358;
wire n_20359;
wire n_20360;
wire n_20361;
wire n_20362;
wire n_20363;
wire n_20364;
wire n_20365;
wire n_20366;
wire n_20367;
wire n_20368;
wire n_20369;
wire n_20370;
wire n_20371;
wire n_20372;
wire n_20373;
wire n_20374;
wire n_20375;
wire n_20376;
wire n_20377;
wire n_20378;
wire n_20379;
wire n_20380;
wire n_20381;
wire n_20382;
wire n_20383;
wire n_20384;
wire n_20385;
wire n_20386;
wire n_20387;
wire n_20388;
wire n_20389;
wire n_20390;
wire n_20391;
wire n_20392;
wire n_20393;
wire n_20394;
wire n_20395;
wire n_20396;
wire n_20397;
wire n_20398;
wire n_20399;
wire n_20400;
wire n_20401;
wire n_20402;
wire n_20403;
wire n_20404;
wire n_20405;
wire n_20406;
wire n_20407;
wire n_20408;
wire n_20409;
wire n_20410;
wire n_20411;
wire n_20412;
wire n_20413;
wire n_20414;
wire n_20415;
wire n_20416;
wire n_20417;
wire n_20418;
wire n_20419;
wire n_20420;
wire n_20421;
wire n_20422;
wire n_20423;
wire n_20424;
wire n_20425;
wire n_20426;
wire n_20427;
wire n_20428;
wire n_20429;
wire n_20430;
wire n_20431;
wire n_20432;
wire n_20433;
wire n_20434;
wire n_20435;
wire n_20436;
wire n_20437;
wire n_20438;
wire n_20439;
wire n_20440;
wire n_20441;
wire n_20442;
wire n_20443;
wire n_20444;
wire n_20445;
wire n_20446;
wire n_20447;
wire n_20448;
wire n_20449;
wire n_20450;
wire n_20451;
wire n_20452;
wire n_20453;
wire n_20454;
wire n_20455;
wire n_20456;
wire n_20457;
wire n_20458;
wire n_20459;
wire n_20460;
wire n_20461;
wire n_20462;
wire n_20463;
wire n_20464;
wire n_20465;
wire n_20466;
wire n_20467;
wire n_20468;
wire n_20469;
wire n_20470;
wire n_20471;
wire n_20472;
wire n_20473;
wire n_20474;
wire n_20475;
wire n_20476;
wire n_20477;
wire n_20478;
wire n_20479;
wire n_20480;
wire n_20481;
wire n_20482;
wire n_20483;
wire n_20484;
wire n_20485;
wire n_20486;
wire n_20487;
wire n_20488;
wire n_20489;
wire n_20490;
wire n_20491;
wire n_20492;
wire n_20493;
wire n_20494;
wire n_20495;
wire n_20496;
wire n_20497;
wire n_20498;
wire n_20499;
wire n_20500;
wire n_20501;
wire n_20502;
wire n_20503;
wire n_20504;
wire n_20505;
wire n_20506;
wire n_20507;
wire n_20508;
wire n_20509;
wire n_20510;
wire n_20511;
wire n_20512;
wire n_20513;
wire n_20514;
wire n_20515;
wire n_20516;
wire n_20517;
wire n_20518;
wire n_20519;
wire n_20520;
wire n_20521;
wire n_20522;
wire n_20523;
wire n_20524;
wire n_20525;
wire n_20526;
wire n_20527;
wire n_20528;
wire n_20529;
wire n_20530;
wire n_20531;
wire n_20532;
wire n_20533;
wire n_20534;
wire n_20535;
wire n_20536;
wire n_20537;
wire n_20538;
wire n_20539;
wire n_20540;
wire n_20541;
wire n_20542;
wire n_20543;
wire n_20544;
wire n_20545;
wire n_20546;
wire n_20547;
wire n_20548;
wire n_20549;
wire n_20550;
wire n_20551;
wire n_20552;
wire n_20553;
wire n_20554;
wire n_20555;
wire n_20556;
wire n_20557;
wire n_20558;
wire n_20559;
wire n_20560;
wire n_20561;
wire n_20562;
wire n_20563;
wire n_20564;
wire n_20565;
wire n_20566;
wire n_20567;
wire n_20568;
wire n_20569;
wire n_20570;
wire n_20571;
wire n_20572;
wire n_20573;
wire n_20574;
wire n_20575;
wire n_20576;
wire n_20577;
wire n_20578;
wire n_20579;
wire n_20580;
wire n_20581;
wire n_20582;
wire n_20583;
wire n_20584;
wire n_20585;
wire n_20586;
wire n_20587;
wire n_20588;
wire n_20589;
wire n_20590;
wire n_20591;
wire n_20592;
wire n_20593;
wire n_20594;
wire n_20595;
wire n_20596;
wire n_20597;
wire n_20598;
wire n_20599;
wire n_20600;
wire n_20601;
wire n_20602;
wire n_20603;
wire n_20604;
wire n_20605;
wire n_20606;
wire n_20607;
wire n_20608;
wire n_20609;
wire n_20610;
wire n_20611;
wire n_20612;
wire n_20613;
wire n_20614;
wire n_20615;
wire n_20616;
wire n_20617;
wire n_20618;
wire n_20619;
wire n_20620;
wire n_20621;
wire n_20622;
wire n_20623;
wire n_20624;
wire n_20625;
wire n_20626;
wire n_20627;
wire n_20628;
wire n_20629;
wire n_20630;
wire n_20631;
wire n_20632;
wire n_20633;
wire n_20634;
wire n_20635;
wire n_20636;
wire n_20637;
wire n_20638;
wire n_20639;
wire n_20640;
wire n_20641;
wire n_20642;
wire n_20643;
wire n_20644;
wire n_20645;
wire n_20646;
wire n_20647;
wire n_20648;
wire n_20649;
wire n_20650;
wire n_20651;
wire n_20652;
wire n_20653;
wire n_20654;
wire n_20655;
wire n_20656;
wire n_20657;
wire n_20658;
wire n_20659;
wire n_20660;
wire n_20661;
wire n_20662;
wire n_20663;
wire n_20664;
wire n_20665;
wire n_20666;
wire n_20667;
wire n_20668;
wire n_20669;
wire n_20670;
wire n_20671;
wire n_20672;
wire n_20673;
wire n_20674;
wire n_20675;
wire n_20676;
wire n_20677;
wire n_20678;
wire n_20679;
wire n_20680;
wire n_20681;
wire n_20682;
wire n_20683;
wire n_20684;
wire n_20685;
wire n_20686;
wire n_20687;
wire n_20688;
wire n_20689;
wire n_20690;
wire n_20691;
wire n_20692;
wire n_20693;
wire n_20694;
wire n_20695;
wire n_20696;
wire n_20697;
wire n_20698;
wire n_20699;
wire n_20700;
wire n_20701;
wire n_20702;
wire n_20703;
wire n_20704;
wire n_20705;
wire n_20706;
wire n_20707;
wire n_20708;
wire n_20709;
wire n_20710;
wire n_20711;
wire n_20712;
wire n_20713;
wire n_20714;
wire n_20715;
wire n_20716;
wire n_20717;
wire n_20718;
wire n_20719;
wire n_20720;
wire n_20721;
wire n_20722;
wire n_20723;
wire n_20724;
wire n_20725;
wire n_20726;
wire n_20727;
wire n_20728;
wire n_20729;
wire n_20730;
wire n_20731;
wire n_20732;
wire n_20733;
wire n_20734;
wire n_20735;
wire n_20736;
wire n_20737;
wire n_20738;
wire n_20739;
wire n_20740;
wire n_20741;
wire n_20742;
wire n_20743;
wire n_20744;
wire n_20745;
wire n_20746;
wire n_20747;
wire n_20748;
wire n_20749;
wire n_20750;
wire n_20751;
wire n_20752;
wire n_20753;
wire n_20754;
wire n_20755;
wire n_20756;
wire n_20757;
wire n_20758;
wire n_20759;
wire n_20760;
wire n_20761;
wire n_20762;
wire n_20763;
wire n_20764;
wire n_20765;
wire n_20766;
wire n_20767;
wire n_20768;
wire n_20769;
wire n_20770;
wire n_20771;
wire n_20772;
wire n_20773;
wire n_20774;
wire n_20775;
wire n_20776;
wire n_20777;
wire n_20778;
wire n_20779;
wire n_20780;
wire n_20781;
wire n_20782;
wire n_20783;
wire n_20784;
wire n_20785;
wire n_20786;
wire n_20787;
wire n_20788;
wire n_20789;
wire n_20790;
wire n_20791;
wire n_20792;
wire n_20793;
wire n_20794;
wire n_20795;
wire n_20796;
wire n_20797;
wire n_20798;
wire n_20799;
wire n_20800;
wire n_20801;
wire n_20802;
wire n_20803;
wire n_20804;
wire n_20805;
wire n_20806;
wire n_20807;
wire n_20808;
wire n_20809;
wire n_20810;
wire n_20811;
wire n_20812;
wire n_20813;
wire n_20814;
wire n_20815;
wire n_20816;
wire n_20817;
wire n_20818;
wire n_20819;
wire n_20820;
wire n_20821;
wire n_20822;
wire n_20823;
wire n_20824;
wire n_20825;
wire n_20826;
wire n_20827;
wire n_20828;
wire n_20829;
wire n_20830;
wire n_20831;
wire n_20832;
wire n_20833;
wire n_20834;
wire n_20835;
wire n_20836;
wire n_20837;
wire n_20838;
wire n_20839;
wire n_20840;
wire n_20841;
wire n_20842;
wire n_20843;
wire n_20844;
wire n_20845;
wire n_20846;
wire n_20847;
wire n_20848;
wire n_20849;
wire n_20850;
wire n_20851;
wire n_20852;
wire n_20853;
wire n_20854;
wire n_20855;
wire n_20856;
wire n_20857;
wire n_20858;
wire n_20859;
wire n_20860;
wire n_20861;
wire n_20862;
wire n_20863;
wire n_20864;
wire n_20865;
wire n_20866;
wire n_20867;
wire n_20868;
wire n_20869;
wire n_20870;
wire n_20871;
wire n_20872;
wire n_20873;
wire n_20874;
wire n_20875;
wire n_20876;
wire n_20877;
wire n_20878;
wire n_20879;
wire n_20880;
wire n_20881;
wire n_20882;
wire n_20883;
wire n_20884;
wire n_20885;
wire n_20886;
wire n_20887;
wire n_20888;
wire n_20889;
wire n_20890;
wire n_20891;
wire n_20892;
wire n_20893;
wire n_20894;
wire n_20895;
wire n_20896;
wire n_20897;
wire n_20898;
wire n_20899;
wire n_20900;
wire n_20901;
wire n_20902;
wire n_20903;
wire n_20904;
wire n_20905;
wire n_20906;
wire n_20907;
wire n_20908;
wire n_20909;
wire n_20910;
wire n_20911;
wire n_20912;
wire n_20913;
wire n_20914;
wire n_20915;
wire n_20916;
wire n_20917;
wire n_20918;
wire n_20919;
wire n_20920;
wire n_20921;
wire n_20922;
wire n_20923;
wire n_20924;
wire n_20925;
wire n_20926;
wire n_20927;
wire n_20928;
wire n_20929;
wire n_20930;
wire n_20931;
wire n_20932;
wire n_20933;
wire n_20934;
wire n_20935;
wire n_20936;
wire n_20937;
wire n_20938;
wire n_20939;
wire n_20940;
wire n_20941;
wire n_20942;
wire n_20943;
wire n_20944;
wire n_20945;
wire n_20946;
wire n_20947;
wire n_20948;
wire n_20949;
wire n_20950;
wire n_20951;
wire n_20952;
wire n_20953;
wire n_20954;
wire n_20955;
wire n_20956;
wire n_20957;
wire n_20958;
wire n_20959;
wire n_20960;
wire n_20961;
wire n_20962;
wire n_20963;
wire n_20964;
wire n_20965;
wire n_20966;
wire n_20967;
wire n_20968;
wire n_20969;
wire n_20970;
wire n_20971;
wire n_20972;
wire n_20973;
wire n_20974;
wire n_20975;
wire n_20976;
wire n_20977;
wire n_20978;
wire n_20979;
wire n_20980;
wire n_20981;
wire n_20982;
wire n_20983;
wire n_20984;
wire n_20985;
wire n_20986;
wire n_20987;
wire n_20988;
wire n_20989;
wire n_20990;
wire n_20991;
wire n_20992;
wire n_20993;
wire n_20994;
wire n_20995;
wire n_20996;
wire n_20997;
wire n_20998;
wire n_20999;
wire n_21000;
wire n_21001;
wire n_21002;
wire n_21003;
wire n_21004;
wire n_21005;
wire n_21006;
wire n_21007;
wire n_21008;
wire n_21009;
wire n_21010;
wire n_21011;
wire n_21012;
wire n_21013;
wire n_21014;
wire n_21015;
wire n_21016;
wire n_21017;
wire n_21018;
wire n_21019;
wire n_21020;
wire n_21021;
wire n_21022;
wire n_21023;
wire n_21024;
wire n_21025;
wire n_21026;
wire n_21027;
wire n_21028;
wire n_21029;
wire n_21030;
wire n_21031;
wire n_21032;
wire n_21033;
wire n_21034;
wire n_21035;
wire n_21036;
wire n_21037;
wire n_21038;
wire n_21039;
wire n_21040;
wire n_21041;
wire n_21042;
wire n_21043;
wire n_21044;
wire n_21045;
wire n_21046;
wire n_21047;
wire n_21048;
wire n_21049;
wire n_21050;
wire n_21051;
wire n_21052;
wire n_21053;
wire n_21054;
wire n_21055;
wire n_21056;
wire n_21057;
wire n_21058;
wire n_21059;
wire n_21060;
wire n_21061;
wire n_21062;
wire n_21063;
wire n_21064;
wire n_21065;
wire n_21066;
wire n_21067;
wire n_21068;
wire n_21069;
wire n_21070;
wire n_21071;
wire n_21072;
wire n_21073;
wire n_21074;
wire n_21075;
wire n_21076;
wire n_21077;
wire n_21078;
wire n_21079;
wire n_21080;
wire n_21081;
wire n_21082;
wire n_21083;
wire n_21084;
wire n_21085;
wire n_21086;
wire n_21087;
wire n_21088;
wire n_21089;
wire n_21090;
wire n_21091;
wire n_21092;
wire n_21093;
wire n_21094;
wire n_21095;
wire n_21096;
wire n_21097;
wire n_21098;
wire n_21099;
wire n_21100;
wire n_21101;
wire n_21102;
wire n_21103;
wire n_21104;
wire n_21105;
wire n_21106;
wire n_21107;
wire n_21108;
wire n_21109;
wire n_21110;
wire n_21111;
wire n_21112;
wire n_21113;
wire n_21114;
wire n_21115;
wire n_21116;
wire n_21117;
wire n_21118;
wire n_21119;
wire n_21120;
wire n_21121;
wire n_21122;
wire n_21123;
wire n_21124;
wire n_21125;
wire n_21126;
wire n_21127;
wire n_21128;
wire n_21129;
wire n_21130;
wire n_21131;
wire n_21132;
wire n_21133;
wire n_21134;
wire n_21135;
wire n_21136;
wire n_21137;
wire n_21138;
wire n_21139;
wire n_21140;
wire n_21141;
wire n_21142;
wire n_21143;
wire n_21144;
wire n_21145;
wire n_21146;
wire n_21147;
wire n_21148;
wire n_21149;
wire n_21150;
wire n_21151;
wire n_21152;
wire n_21153;
wire n_21154;
wire n_21155;
wire n_21156;
wire n_21157;
wire n_21158;
wire n_21159;
wire n_21160;
wire n_21161;
wire n_21162;
wire n_21163;
wire n_21164;
wire n_21165;
wire n_21166;
wire n_21167;
wire n_21168;
wire n_21169;
wire n_21170;
wire n_21171;
wire n_21172;
wire n_21173;
wire n_21174;
wire n_21175;
wire n_21176;
wire n_21177;
wire n_21178;
wire n_21179;
wire n_21180;
wire n_21181;
wire n_21182;
wire n_21183;
wire n_21184;
wire n_21185;
wire n_21186;
wire n_21187;
wire n_21188;
wire n_21189;
wire n_21190;
wire n_21191;
wire n_21192;
wire n_21193;
wire n_21194;
wire n_21195;
wire n_21196;
wire n_21197;
wire n_21198;
wire n_21199;
wire n_21200;
wire n_21201;
wire n_21202;
wire n_21203;
wire n_21204;
wire n_21205;
wire n_21206;
wire n_21207;
wire n_21208;
wire n_21209;
wire n_21210;
wire n_21211;
wire n_21212;
wire n_21213;
wire n_21214;
wire n_21215;
wire n_21216;
wire n_21217;
wire n_21218;
wire n_21219;
wire n_21220;
wire n_21221;
wire n_21222;
wire n_21223;
wire n_21224;
wire n_21225;
wire n_21226;
wire n_21227;
wire n_21228;
wire n_21229;
wire n_21230;
wire n_21231;
wire n_21232;
wire n_21233;
wire n_21234;
wire n_21235;
wire n_21236;
wire n_21237;
wire n_21238;
wire n_21239;
wire n_21240;
wire n_21241;
wire n_21242;
wire n_21243;
wire n_21244;
wire n_21245;
wire n_21246;
wire n_21247;
wire n_21248;
wire n_21249;
wire n_21250;
wire n_21251;
wire n_21252;
wire n_21253;
wire n_21254;
wire n_21255;
wire n_21256;
wire n_21257;
wire n_21258;
wire n_21259;
wire n_21260;
wire n_21261;
wire n_21262;
wire n_21263;
wire n_21264;
wire n_21265;
wire n_21266;
wire n_21267;
wire n_21268;
wire n_21269;
wire n_21270;
wire n_21271;
wire n_21272;
wire n_21273;
wire n_21274;
wire n_21275;
wire n_21276;
wire n_21277;
wire n_21278;
wire n_21279;
wire n_21280;
wire n_21281;
wire n_21282;
wire n_21283;
wire n_21284;
wire n_21285;
wire n_21286;
wire n_21287;
wire n_21288;
wire n_21289;
wire n_21290;
wire n_21291;
wire n_21292;
wire n_21293;
wire n_21294;
wire n_21295;
wire n_21296;
wire n_21297;
wire n_21298;
wire n_21299;
wire n_21300;
wire n_21301;
wire n_21302;
wire n_21303;
wire n_21304;
wire n_21305;
wire n_21306;
wire n_21307;
wire n_21308;
wire n_21309;
wire n_21310;
wire n_21311;
wire n_21312;
wire n_21313;
wire n_21314;
wire n_21315;
wire n_21316;
wire n_21317;
wire n_21318;
wire n_21319;
wire n_21320;
wire n_21321;
wire n_21322;
wire n_21323;
wire n_21324;
wire n_21325;
wire n_21326;
wire n_21327;
wire n_21328;
wire n_21329;
wire n_21330;
wire n_21331;
wire n_21332;
wire n_21333;
wire n_21334;
wire n_21335;
wire n_21336;
wire n_21337;
wire n_21338;
wire n_21339;
wire n_21340;
wire n_21341;
wire n_21342;
wire n_21343;
wire n_21344;
wire n_21345;
wire n_21346;
wire n_21347;
wire n_21348;
wire n_21349;
wire n_21350;
wire n_21351;
wire n_21352;
wire n_21353;
wire n_21354;
wire n_21355;
wire n_21356;
wire n_21357;
wire n_21358;
wire n_21359;
wire n_21360;
wire n_21361;
wire n_21362;
wire n_21363;
wire n_21364;
wire n_21365;
wire n_21366;
wire n_21367;
wire n_21368;
wire n_21369;
wire n_21370;
wire n_21371;
wire n_21372;
wire n_21373;
wire n_21374;
wire n_21375;
wire n_21376;
wire n_21377;
wire n_21378;
wire n_21379;
wire n_21380;
wire n_21381;
wire n_21382;
wire n_21383;
wire n_21384;
wire n_21385;
wire n_21386;
wire n_21387;
wire n_21388;
wire n_21389;
wire n_21390;
wire n_21391;
wire n_21392;
wire n_21393;
wire n_21394;
wire n_21395;
wire n_21396;
wire n_21397;
wire n_21398;
wire n_21399;
wire n_21400;
wire n_21401;
wire n_21402;
wire n_21403;
wire n_21404;
wire n_21405;
wire n_21406;
wire n_21407;
wire n_21408;
wire n_21409;
wire n_21410;
wire n_21411;
wire n_21412;
wire n_21413;
wire n_21414;
wire n_21415;
wire n_21416;
wire n_21417;
wire n_21418;
wire n_21419;
wire n_21420;
wire n_21421;
wire n_21422;
wire n_21423;
wire n_21424;
wire n_21425;
wire n_21426;
wire n_21427;
wire n_21428;
wire n_21429;
wire n_21430;
wire n_21431;
wire n_21432;
wire n_21433;
wire n_21434;
wire n_21435;
wire n_21436;
wire n_21437;
wire n_21438;
wire n_21439;
wire n_21440;
wire n_21441;
wire n_21442;
wire n_21443;
wire n_21444;
wire n_21445;
wire n_21446;
wire n_21447;
wire n_21448;
wire n_21449;
wire n_21450;
wire n_21451;
wire n_21452;
wire n_21453;
wire n_21454;
wire n_21455;
wire n_21456;
wire n_21457;
wire n_21458;
wire n_21459;
wire n_21460;
wire n_21461;
wire n_21462;
wire n_21463;
wire n_21464;
wire n_21465;
wire n_21466;
wire n_21467;
wire n_21468;
wire n_21469;
wire n_21470;
wire n_21471;
wire n_21472;
wire n_21473;
wire n_21474;
wire n_21475;
wire n_21476;
wire n_21477;
wire n_21478;
wire n_21479;
wire n_21480;
wire n_21481;
wire n_21482;
wire n_21483;
wire n_21484;
wire n_21485;
wire n_21486;
wire n_21487;
wire n_21488;
wire n_21489;
wire n_21490;
wire n_21491;
wire n_21492;
wire n_21493;
wire n_21494;
wire n_21495;
wire n_21496;
wire n_21497;
wire n_21498;
wire n_21499;
wire n_21500;
wire n_21501;
wire n_21502;
wire n_21503;
wire n_21504;
wire n_21505;
wire n_21506;
wire n_21507;
wire n_21508;
wire n_21509;
wire n_21510;
wire n_21511;
wire n_21512;
wire n_21513;
wire n_21514;
wire n_21515;
wire n_21516;
wire n_21517;
wire n_21518;
wire n_21519;
wire n_21520;
wire n_21521;
wire n_21522;
wire n_21523;
wire n_21524;
wire n_21525;
wire n_21526;
wire n_21527;
wire n_21528;
wire n_21529;
wire n_21530;
wire n_21531;
wire n_21532;
wire n_21533;
wire n_21534;
wire n_21535;
wire n_21536;
wire n_21537;
wire n_21538;
wire n_21539;
wire n_21540;
wire n_21541;
wire n_21542;
wire n_21543;
wire n_21544;
wire n_21545;
wire n_21546;
wire n_21547;
wire n_21548;
wire n_21549;
wire n_21550;
wire n_21551;
wire n_21552;
wire n_21553;
wire n_21554;
wire n_21555;
wire n_21556;
wire n_21557;
wire n_21558;
wire n_21559;
wire n_21560;
wire n_21561;
wire n_21562;
wire n_21563;
wire n_21564;
wire n_21565;
wire n_21566;
wire n_21567;
wire n_21568;
wire n_21569;
wire n_21570;
wire n_21571;
wire n_21572;
wire n_21573;
wire n_21574;
wire n_21575;
wire n_21576;
wire n_21577;
wire n_21578;
wire n_21579;
wire n_21580;
wire n_21581;
wire n_21582;
wire n_21583;
wire n_21584;
wire n_21585;
wire n_21586;
wire n_21587;
wire n_21588;
wire n_21589;
wire n_21590;
wire n_21591;
wire n_21592;
wire n_21593;
wire n_21594;
wire n_21595;
wire n_21596;
wire n_21597;
wire n_21598;
wire n_21599;
wire n_21600;
wire n_21601;
wire n_21602;
wire n_21603;
wire n_21604;
wire n_21605;
wire n_21606;
wire n_21607;
wire n_21608;
wire n_21609;
wire n_21610;
wire n_21611;
wire n_21612;
wire n_21613;
wire n_21614;
wire n_21615;
wire n_21616;
wire n_21617;
wire n_21618;
wire n_21619;
wire n_21620;
wire n_21621;
wire n_21622;
wire n_21623;
wire n_21624;
wire n_21625;
wire n_21626;
wire n_21627;
wire n_21628;
wire n_21629;
wire n_21630;
wire n_21631;
wire n_21632;
wire n_21633;
wire n_21634;
wire n_21635;
wire n_21636;
wire n_21637;
wire n_21638;
wire n_21639;
wire n_21640;
wire n_21641;
wire n_21642;
wire n_21643;
wire n_21644;
wire n_21645;
wire n_21646;
wire n_21647;
wire n_21648;
wire n_21649;
wire n_21650;
wire n_21651;
wire n_21652;
wire n_21653;
wire n_21654;
wire n_21655;
wire n_21656;
wire n_21657;
wire n_21658;
wire n_21659;
wire n_21660;
wire n_21661;
wire n_21662;
wire n_21663;
wire n_21664;
wire n_21665;
wire n_21666;
wire n_21667;
wire n_21668;
wire n_21669;
wire n_21670;
wire n_21671;
wire n_21672;
wire n_21673;
wire n_21674;
wire n_21675;
wire n_21676;
wire n_21677;
wire n_21678;
wire n_21679;
wire n_21680;
wire n_21681;
wire n_21682;
wire n_21683;
wire n_21684;
wire n_21685;
wire n_21686;
wire n_21687;
wire n_21688;
wire n_21689;
wire n_21690;
wire n_21691;
wire n_21692;
wire n_21693;
wire n_21694;
wire n_21695;
wire n_21696;
wire n_21697;
wire n_21698;
wire n_21699;
wire n_21700;
wire n_21701;
wire n_21702;
wire n_21703;
wire n_21704;
wire n_21705;
wire n_21706;
wire n_21707;
wire n_21708;
wire n_21709;
wire n_21710;
wire n_21711;
wire n_21712;
wire n_21713;
wire n_21714;
wire n_21715;
wire n_21716;
wire n_21717;
wire n_21718;
wire n_21719;
wire n_21720;
wire n_21721;
wire n_21722;
wire n_21723;
wire n_21724;
wire n_21725;
wire n_21726;
wire n_21727;
wire n_21728;
wire n_21729;
wire n_21730;
wire n_21731;
wire n_21732;
wire n_21733;
wire n_21734;
wire n_21735;
wire n_21736;
wire n_21737;
wire n_21738;
wire n_21739;
wire n_21740;
wire n_21741;
wire n_21742;
wire n_21743;
wire n_21744;
wire n_21745;
wire n_21746;
wire n_21747;
wire n_21748;
wire n_21749;
wire n_21750;
wire n_21751;
wire n_21752;
wire n_21753;
wire n_21754;
wire n_21755;
wire n_21756;
wire n_21757;
wire n_21758;
wire n_21759;
wire n_21760;
wire n_21761;
wire n_21762;
wire n_21763;
wire n_21764;
wire n_21765;
wire n_21766;
wire n_21767;
wire n_21768;
wire n_21769;
wire n_21770;
wire n_21771;
wire n_21772;
wire n_21773;
wire n_21774;
wire n_21775;
wire n_21776;
wire n_21777;
wire n_21778;
wire n_21779;
wire n_21780;
wire n_21781;
wire n_21782;
wire n_21783;
wire n_21784;
wire n_21785;
wire n_21786;
wire n_21787;
wire n_21788;
wire n_21789;
wire n_21790;
wire n_21791;
wire n_21792;
wire n_21793;
wire n_21794;
wire n_21795;
wire n_21796;
wire n_21797;
wire n_21798;
wire n_21799;
wire n_21800;
wire n_21801;
wire n_21802;
wire n_21803;
wire n_21804;
wire n_21805;
wire n_21806;
wire n_21807;
wire n_21808;
wire n_21809;
wire n_21810;
wire n_21811;
wire n_21812;
wire n_21813;
wire n_21814;
wire n_21815;
wire n_21816;
wire n_21817;
wire n_21818;
wire n_21819;
wire n_21820;
wire n_21821;
wire n_21822;
wire n_21823;
wire n_21824;
wire n_21825;
wire n_21826;
wire n_21827;
wire n_21828;
wire n_21829;
wire n_21830;
wire n_21831;
wire n_21832;
wire n_21833;
wire n_21834;
wire n_21835;
wire n_21836;
wire n_21837;
wire n_21838;
wire n_21839;
wire n_21840;
wire n_21841;
wire n_21842;
wire n_21843;
wire n_21844;
wire n_21845;
wire n_21846;
wire n_21847;
wire n_21848;
wire n_21849;
wire n_21850;
wire n_21851;
wire n_21852;
wire n_21853;
wire n_21854;
wire n_21855;
wire n_21856;
wire n_21857;
wire n_21858;
wire n_21859;
wire n_21860;
wire n_21861;
wire n_21862;
wire n_21863;
wire n_21864;
wire n_21865;
wire n_21866;
wire n_21867;
wire n_21868;
wire n_21869;
wire n_21870;
wire n_21871;
wire n_21872;
wire n_21873;
wire n_21874;
wire n_21875;
wire n_21876;
wire n_21877;
wire n_21878;
wire n_21879;
wire n_21880;
wire n_21881;
wire n_21882;
wire n_21883;
wire n_21884;
wire n_21885;
wire n_21886;
wire n_21887;
wire n_21888;
wire n_21889;
wire n_21890;
wire n_21891;
wire n_21892;
wire n_21893;
wire n_21894;
wire n_21895;
wire n_21896;
wire n_21897;
wire n_21898;
wire n_21899;
wire n_21900;
wire n_21901;
wire n_21902;
wire n_21903;
wire n_21904;
wire n_21905;
wire n_21906;
wire n_21907;
wire n_21908;
wire n_21909;
wire n_21910;
wire n_21911;
wire n_21912;
wire n_21913;
wire n_21914;
wire n_21915;
wire n_21916;
wire n_21917;
wire n_21918;
wire n_21919;
wire n_21920;
wire n_21921;
wire n_21922;
wire n_21923;
wire n_21924;
wire n_21925;
wire n_21926;
wire n_21927;
wire n_21928;
wire n_21929;
wire n_21930;
wire n_21931;
wire n_21932;
wire n_21933;
wire n_21934;
wire n_21935;
wire n_21936;
wire n_21937;
wire n_21938;
wire n_21939;
wire n_21940;
wire n_21941;
wire n_21942;
wire n_21943;
wire n_21944;
wire n_21945;
wire n_21946;
wire n_21947;
wire n_21948;
wire n_21949;
wire n_21950;
wire n_21951;
wire n_21952;
wire n_21953;
wire n_21954;
wire n_21955;
wire n_21956;
wire n_21957;
wire n_21958;
wire n_21959;
wire n_21960;
wire n_21961;
wire n_21962;
wire n_21963;
wire n_21964;
wire n_21965;
wire n_21966;
wire n_21967;
wire n_21968;
wire n_21969;
wire n_21970;
wire n_21971;
wire n_21972;
wire n_21973;
wire n_21974;
wire n_21975;
wire n_21976;
wire n_21977;
wire n_21978;
wire n_21979;
wire n_21980;
wire n_21981;
wire n_21982;
wire n_21983;
wire n_21984;
wire n_21985;
wire n_21986;
wire n_21987;
wire n_21988;
wire n_21989;
wire n_21990;
wire n_21991;
wire n_21992;
wire n_21993;
wire n_21994;
wire n_21995;
wire n_21996;
wire n_21997;
wire n_21998;
wire n_21999;
wire n_22000;
wire n_22001;
wire n_22002;
wire n_22003;
wire n_22004;
wire n_22005;
wire n_22006;
wire n_22007;
wire n_22008;
wire n_22009;
wire n_22010;
wire n_22011;
wire n_22012;
wire n_22013;
wire n_22014;
wire n_22015;
wire n_22016;
wire n_22017;
wire n_22018;
wire n_22019;
wire n_22020;
wire n_22021;
wire n_22022;
wire n_22023;
wire n_22024;
wire n_22025;
wire n_22026;
wire n_22027;
wire n_22028;
wire n_22029;
wire n_22030;
wire n_22031;
wire n_22032;
wire n_22033;
wire n_22034;
wire n_22035;
wire n_22036;
wire n_22037;
wire n_22038;
wire n_22039;
wire n_22040;
wire n_22041;
wire n_22042;
wire n_22043;
wire n_22044;
wire n_22045;
wire n_22046;
wire n_22047;
wire n_22048;
wire n_22049;
wire n_22050;
wire n_22051;
wire n_22052;
wire n_22053;
wire n_22054;
wire n_22055;
wire n_22056;
wire n_22057;
wire n_22058;
wire n_22059;
wire n_22060;
wire n_22061;
wire n_22062;
wire n_22063;
wire n_22064;
wire n_22065;
wire n_22066;
wire n_22067;
wire n_22068;
wire n_22069;
wire n_22070;
wire n_22071;
wire n_22072;
wire n_22073;
wire n_22074;
wire n_22075;
wire n_22076;
wire n_22077;
wire n_22078;
wire n_22079;
wire n_22080;
wire n_22081;
wire n_22082;
wire n_22083;
wire n_22084;
wire n_22085;
wire n_22086;
wire n_22087;
wire n_22088;
wire n_22089;
wire n_22090;
wire n_22091;
wire n_22092;
wire n_22093;
wire n_22094;
wire n_22095;
wire n_22096;
wire n_22097;
wire n_22098;
wire n_22099;
wire n_22100;
wire n_22101;
wire n_22102;
wire n_22103;
wire n_22104;
wire n_22105;
wire n_22106;
wire n_22107;
wire n_22108;
wire n_22109;
wire n_22110;
wire n_22111;
wire n_22112;
wire n_22113;
wire n_22114;
wire n_22115;
wire n_22116;
wire n_22117;
wire n_22118;
wire n_22119;
wire n_22120;
wire n_22121;
wire n_22122;
wire n_22123;
wire n_22124;
wire n_22125;
wire n_22126;
wire n_22127;
wire n_22128;
wire n_22129;
wire n_22130;
wire n_22131;
wire n_22132;
wire n_22133;
wire n_22134;
wire n_22135;
wire n_22136;
wire n_22137;
wire n_22138;
wire n_22139;
wire n_22140;
wire n_22141;
wire n_22142;
wire n_22143;
wire n_22144;
wire n_22145;
wire n_22146;
wire n_22147;
wire n_22148;
wire n_22149;
wire n_22150;
wire n_22151;
wire n_22152;
wire n_22153;
wire n_22154;
wire n_22155;
wire n_22156;
wire n_22157;
wire n_22158;
wire n_22159;
wire n_22160;
wire n_22161;
wire n_22162;
wire n_22163;
wire n_22164;
wire n_22165;
wire n_22166;
wire n_22167;
wire n_22168;
wire n_22169;
wire n_22170;
wire n_22171;
wire n_22172;
wire n_22173;
wire n_22174;
wire n_22175;
wire n_22176;
wire n_22177;
wire n_22178;
wire n_22179;
wire n_22180;
wire n_22181;
wire n_22182;
wire n_22183;
wire n_22184;
wire n_22185;
wire n_22186;
wire n_22187;
wire n_22188;
wire n_22189;
wire n_22190;
wire n_22191;
wire n_22192;
wire n_22193;
wire n_22194;
wire n_22195;
wire n_22196;
wire n_22197;
wire n_22198;
wire n_22199;
wire n_22200;
wire n_22201;
wire n_22202;
wire n_22203;
wire n_22204;
wire n_22205;
wire n_22206;
wire n_22207;
wire n_22208;
wire n_22209;
wire n_22210;
wire n_22211;
wire n_22212;
wire n_22213;
wire n_22214;
wire n_22215;
wire n_22216;
wire n_22217;
wire n_22218;
wire n_22219;
wire n_22220;
wire n_22221;
wire n_22222;
wire n_22223;
wire n_22224;
wire n_22225;
wire n_22226;
wire n_22227;
wire n_22228;
wire n_22229;
wire n_22230;
wire n_22231;
wire n_22232;
wire n_22233;
wire n_22234;
wire n_22235;
wire n_22236;
wire n_22237;
wire n_22238;
wire n_22239;
wire n_22240;
wire n_22241;
wire n_22242;
wire n_22243;
wire n_22244;
wire n_22245;
wire n_22246;
wire n_22247;
wire n_22248;
wire n_22249;
wire n_22250;
wire n_22251;
wire n_22252;
wire n_22253;
wire n_22254;
wire n_22255;
wire n_22256;
wire n_22257;
wire n_22258;
wire n_22259;
wire n_22260;
wire n_22261;
wire n_22262;
wire n_22263;
wire n_22264;
wire n_22265;
wire n_22266;
wire n_22267;
wire n_22268;
wire n_22269;
wire n_22270;
wire n_22271;
wire n_22272;
wire n_22273;
wire n_22274;
wire n_22275;
wire n_22276;
wire n_22277;
wire n_22278;
wire n_22279;
wire n_22280;
wire n_22281;
wire n_22282;
wire n_22283;
wire n_22284;
wire n_22285;
wire n_22286;
wire n_22287;
wire n_22288;
wire n_22289;
wire n_22290;
wire n_22291;
wire n_22292;
wire n_22293;
wire n_22294;
wire n_22295;
wire n_22296;
wire n_22297;
wire n_22298;
wire n_22299;
wire n_22300;
wire n_22301;
wire n_22302;
wire n_22303;
wire n_22304;
wire n_22305;
wire n_22306;
wire n_22307;
wire n_22308;
wire n_22309;
wire n_22310;
wire n_22311;
wire n_22312;
wire n_22313;
wire n_22314;
wire n_22315;
wire n_22316;
wire n_22317;
wire n_22318;
wire n_22319;
wire n_22320;
wire n_22321;
wire n_22322;
wire n_22323;
wire n_22324;
wire n_22325;
wire n_22326;
wire n_22327;
wire n_22328;
wire n_22329;
wire n_22330;
wire n_22331;
wire n_22332;
wire n_22333;
wire n_22334;
wire n_22335;
wire n_22336;
wire n_22337;
wire n_22338;
wire n_22339;
wire n_22340;
wire n_22341;
wire n_22342;
wire n_22343;
wire n_22344;
wire n_22345;
wire n_22346;
wire n_22347;
wire n_22348;
wire n_22349;
wire n_22350;
wire n_22351;
wire n_22352;
wire n_22353;
wire n_22354;
wire n_22355;
wire n_22356;
wire n_22357;
wire n_22358;
wire n_22359;
wire n_22360;
wire n_22361;
wire n_22362;
wire n_22363;
wire n_22364;
wire n_22365;
wire n_22366;
wire n_22367;
wire n_22368;
wire n_22369;
wire n_22370;
wire n_22371;
wire n_22372;
wire n_22373;
wire n_22374;
wire n_22375;
wire n_22376;
wire n_22377;
wire n_22378;
wire n_22379;
wire n_22380;
wire n_22381;
wire n_22382;
wire n_22383;
wire n_22384;
wire n_22385;
wire n_22386;
wire n_22387;
wire n_22388;
wire n_22389;
wire n_22390;
wire n_22391;
wire n_22392;
wire n_22393;
wire n_22394;
wire n_22395;
wire n_22396;
wire n_22397;
wire n_22398;
wire n_22399;
wire n_22400;
wire n_22401;
wire n_22402;
wire n_22403;
wire n_22404;
wire n_22405;
wire n_22406;
wire n_22407;
wire n_22408;
wire n_22409;
wire n_22410;
wire n_22411;
wire n_22412;
wire n_22413;
wire n_22414;
wire n_22415;
wire n_22416;
wire n_22417;
wire n_22418;
wire n_22419;
wire n_22420;
wire n_22421;
wire n_22422;
wire n_22423;
wire n_22424;
wire n_22425;
wire n_22426;
wire n_22427;
wire n_22428;
wire n_22429;
wire n_22430;
wire n_22431;
wire n_22432;
wire n_22433;
wire n_22434;
wire n_22435;
wire n_22436;
wire n_22437;
wire n_22438;
wire n_22439;
wire n_22440;
wire n_22441;
wire n_22442;
wire n_22443;
wire n_22444;
wire n_22445;
wire n_22446;
wire n_22447;
wire n_22448;
wire n_22449;
wire n_22450;
wire n_22451;
wire n_22452;
wire n_22453;
wire n_22454;
wire n_22455;
wire n_22456;
wire n_22457;
wire n_22458;
wire n_22459;
wire n_22460;
wire n_22461;
wire n_22462;
wire n_22463;
wire n_22464;
wire n_22465;
wire n_22466;
wire n_22467;
wire n_22468;
wire n_22469;
wire n_22470;
wire n_22471;
wire n_22472;
wire n_22473;
wire n_22474;
wire n_22475;
wire n_22476;
wire n_22477;
wire n_22478;
wire n_22479;
wire n_22480;
wire n_22481;
wire n_22482;
wire n_22483;
wire n_22484;
wire n_22485;
wire n_22486;
wire n_22487;
wire n_22488;
wire n_22489;
wire n_22490;
wire n_22491;
wire n_22492;
wire n_22493;
wire n_22494;
wire n_22495;
wire n_22496;
wire n_22497;
wire n_22498;
wire n_22499;
wire n_22500;
wire n_22501;
wire n_22502;
wire n_22503;
wire n_22504;
wire n_22505;
wire n_22506;
wire n_22507;
wire n_22508;
wire n_22509;
wire n_22510;
wire n_22511;
wire n_22512;
wire n_22513;
wire n_22514;
wire n_22515;
wire n_22516;
wire n_22517;
wire n_22518;
wire n_22519;
wire n_22520;
wire n_22521;
wire n_22522;
wire n_22523;
wire n_22524;
wire n_22525;
wire n_22526;
wire n_22527;
wire n_22528;
wire n_22529;
wire n_22530;
wire n_22531;
wire n_22532;
wire n_22533;
wire n_22534;
wire n_22535;
wire n_22536;
wire n_22537;
wire n_22538;
wire n_22539;
wire n_22540;
wire n_22541;
wire n_22542;
wire n_22543;
wire n_22544;
wire n_22545;
wire n_22546;
wire n_22547;
wire n_22548;
wire n_22549;
wire n_22550;
wire n_22551;
wire n_22552;
wire n_22553;
wire n_22554;
wire n_22555;
wire n_22556;
wire n_22557;
wire n_22558;
wire n_22559;
wire n_22560;
wire n_22561;
wire n_22562;
wire n_22563;
wire n_22564;
wire n_22565;
wire n_22566;
wire n_22567;
wire n_22568;
wire n_22569;
wire n_22570;
wire n_22571;
wire n_22572;
wire n_22573;
wire n_22574;
wire n_22575;
wire n_22576;
wire n_22577;
wire n_22578;
wire n_22579;
wire n_22580;
wire n_22581;
wire n_22582;
wire n_22583;
wire n_22584;
wire n_22585;
wire n_22586;
wire n_22587;
wire n_22588;
wire n_22589;
wire n_22590;
wire n_22591;
wire n_22592;
wire n_22593;
wire n_22594;
wire n_22595;
wire n_22596;
wire n_22597;
wire n_22598;
wire n_22599;
wire n_22600;
wire n_22601;
wire n_22602;
wire n_22603;
wire n_22604;
wire n_22605;
wire n_22606;
wire n_22607;
wire n_22608;
wire n_22609;
wire n_22610;
wire n_22611;
wire n_22612;
wire n_22613;
wire n_22614;
wire n_22615;
wire n_22616;
wire n_22617;
wire n_22618;
wire n_22619;
wire n_22620;
wire n_22621;
wire n_22622;
wire n_22623;
wire n_22624;
wire n_22625;
wire n_22626;
wire n_22627;
wire n_22628;
wire n_22629;
wire n_22630;
wire n_22631;
wire n_22632;
wire n_22633;
wire n_22634;
wire n_22635;
wire n_22636;
wire n_22637;
wire n_22638;
wire n_22639;
wire n_22640;
wire n_22641;
wire n_22642;
wire n_22643;
wire n_22644;
wire n_22645;
wire n_22646;
wire n_22647;
wire n_22648;
wire n_22649;
wire n_22650;
wire n_22651;
wire n_22652;
wire n_22653;
wire n_22654;
wire n_22655;
wire n_22656;
wire n_22657;
wire n_22658;
wire n_22659;
wire n_22660;
wire n_22661;
wire n_22662;
wire n_22663;
wire n_22664;
wire n_22665;
wire n_22666;
wire n_22667;
wire n_22668;
wire n_22669;
wire n_22670;
wire n_22671;
wire n_22672;
wire n_22673;
wire n_22674;
wire n_22675;
wire n_22676;
wire n_22677;
wire n_22678;
wire n_22679;
wire n_22680;
wire n_22681;
wire n_22682;
wire n_22683;
wire n_22684;
wire n_22685;
wire n_22686;
wire n_22687;
wire n_22688;
wire n_22689;
wire n_22690;
wire n_22691;
wire n_22692;
wire n_22693;
wire n_22694;
wire n_22695;
wire n_22696;
wire n_22697;
wire n_22698;
wire n_22699;
wire n_22700;
wire n_22701;
wire n_22702;
wire n_22703;
wire n_22704;
wire n_22705;
wire n_22706;
wire n_22707;
wire n_22708;
wire n_22709;
wire n_22710;
wire n_22711;
wire n_22712;
wire n_22713;
wire n_22714;
wire n_22715;
wire n_22716;
wire n_22717;
wire n_22718;
wire n_22719;
wire n_22720;
wire n_22721;
wire n_22722;
wire n_22723;
wire n_22724;
wire n_22725;
wire n_22726;
wire n_22727;
wire n_22728;
wire n_22729;
wire n_22730;
wire n_22731;
wire n_22732;
wire n_22733;
wire n_22734;
wire n_22735;
wire n_22736;
wire n_22737;
wire n_22738;
wire n_22739;
wire n_22740;
wire n_22741;
wire n_22742;
wire n_22743;
wire n_22744;
wire n_22745;
wire n_22746;
wire n_22747;
wire n_22748;
wire n_22749;
wire n_22750;
wire n_22751;
wire n_22752;
wire n_22753;
wire n_22754;
wire n_22755;
wire n_22756;
wire n_22757;
wire n_22758;
wire n_22759;
wire n_22760;
wire n_22761;
wire n_22762;
wire n_22763;
wire n_22764;
wire n_22765;
wire n_22766;
wire n_22767;
wire n_22768;
wire n_22769;
wire n_22770;
wire n_22771;
wire n_22772;
wire n_22773;
wire n_22774;
wire n_22775;
wire n_22776;
wire n_22777;
wire n_22778;
wire n_22779;
wire n_22780;
wire n_22781;
wire n_22782;
wire n_22783;
wire n_22784;
wire n_22785;
wire n_22786;
wire n_22787;
wire n_22788;
wire n_22789;
wire n_22790;
wire n_22791;
wire n_22792;
wire n_22793;
wire n_22794;
wire n_22795;
wire n_22796;
wire n_22797;
wire n_22798;
wire n_22799;
wire n_22800;
wire n_22801;
wire n_22802;
wire n_22803;
wire n_22804;
wire n_22805;
wire n_22806;
wire n_22807;
wire n_22808;
wire n_22809;
wire n_22810;
wire n_22811;
wire n_22812;
wire n_22813;
wire n_22814;
wire n_22815;
wire n_22816;
wire n_22817;
wire n_22818;
wire n_22819;
wire n_22820;
wire n_22821;
wire n_22822;
wire n_22823;
wire n_22824;
wire n_22825;
wire n_22826;
wire n_22827;
wire n_22828;
wire n_22829;
wire n_22830;
wire n_22831;
wire n_22832;
wire n_22833;
wire n_22834;
wire n_22835;
wire n_22836;
wire n_22837;
wire n_22838;
wire n_22839;
wire n_22840;
wire n_22841;
wire n_22842;
wire n_22843;
wire n_22844;
wire n_22845;
wire n_22846;
wire n_22847;
wire n_22848;
wire n_22849;
wire n_22850;
wire n_22851;
wire n_22852;
wire n_22853;
wire n_22854;
wire n_22855;
wire n_22856;
wire n_22857;
wire n_22858;
wire n_22859;
wire n_22860;
wire n_22861;
wire n_22862;
wire n_22863;
wire n_22864;
wire n_22865;
wire n_22866;
wire n_22867;
wire n_22868;
wire n_22869;
wire n_22870;
wire n_22871;
wire n_22872;
wire n_22873;
wire n_22874;
wire n_22875;
wire n_22876;
wire n_22877;
wire n_22878;
wire n_22879;
wire n_22880;
wire n_22881;
wire n_22882;
wire n_22883;
wire n_22884;
wire n_22885;
wire n_22886;
wire n_22887;
wire n_22888;
wire n_22889;
wire n_22890;
wire n_22891;
wire n_22892;
wire n_22893;
wire n_22894;
wire n_22895;
wire n_22896;
wire n_22897;
wire n_22898;
wire n_22899;
wire n_22900;
wire n_22901;
wire n_22902;
wire n_22903;
wire n_22904;
wire n_22905;
wire n_22906;
wire n_22907;
wire n_22908;
wire n_22909;
wire n_22910;
wire n_22911;
wire n_22912;
wire n_22913;
wire n_22914;
wire n_22915;
wire n_22916;
wire n_22917;
wire n_22918;
wire n_22919;
wire n_22920;
wire n_22921;
wire n_22922;
wire n_22923;
wire n_22924;
wire n_22925;
wire n_22926;
wire n_22927;
wire n_22928;
wire n_22929;
wire n_22930;
wire n_22931;
wire n_22932;
wire n_22933;
wire n_22934;
wire n_22935;
wire n_22936;
wire n_22937;
wire n_22938;
wire n_22939;
wire n_22940;
wire n_22941;
wire n_22942;
wire n_22943;
wire n_22944;
wire n_22945;
wire n_22946;
wire n_22947;
wire n_22948;
wire n_22949;
wire n_22950;
wire n_22951;
wire n_22952;
wire n_22953;
wire n_22954;
wire n_22955;
wire n_22956;
wire n_22957;
wire n_22958;
wire n_22959;
wire n_22960;
wire n_22961;
wire n_22962;
wire n_22963;
wire n_22964;
wire n_22965;
wire n_22966;
wire n_22967;
wire n_22968;
wire n_22969;
wire n_22970;
wire n_22971;
wire n_22972;
wire n_22973;
wire n_22974;
wire n_22975;
wire n_22976;
wire n_22977;
wire n_22978;
wire n_22979;
wire n_22980;
wire n_22981;
wire n_22982;
wire n_22983;
wire n_22984;
wire n_22985;
wire n_22986;
wire n_22987;
wire n_22988;
wire n_22989;
wire n_22990;
wire n_22991;
wire n_22992;
wire n_22993;
wire n_22994;
wire n_22995;
wire n_22996;
wire n_22997;
wire n_22998;
wire n_22999;
wire n_23000;
wire n_23001;
wire n_23002;
wire n_23003;
wire n_23004;
wire n_23005;
wire n_23006;
wire n_23007;
wire n_23008;
wire n_23009;
wire n_23010;
wire n_23011;
wire n_23012;
wire n_23013;
wire n_23014;
wire n_23015;
wire n_23016;
wire n_23017;
wire n_23018;
wire n_23019;
wire n_23020;
wire n_23021;
wire n_23022;
wire n_23023;
wire n_23024;
wire n_23025;
wire n_23026;
wire n_23027;
wire n_23028;
wire n_23029;
wire n_23030;
wire n_23031;
wire n_23032;
wire n_23033;
wire n_23034;
wire n_23035;
wire n_23036;
wire n_23037;
wire n_23038;
wire n_23039;
wire n_23040;
wire n_23041;
wire n_23042;
wire n_23043;
wire n_23044;
wire n_23045;
wire n_23046;
wire n_23047;
wire n_23048;
wire n_23049;
wire n_23050;
wire n_23051;
wire n_23052;
wire n_23053;
wire n_23054;
wire n_23055;
wire n_23056;
wire n_23057;
wire n_23058;
wire n_23059;
wire n_23060;
wire n_23061;
wire n_23062;
wire n_23063;
wire n_23064;
wire n_23065;
wire n_23066;
wire n_23067;
wire n_23068;
wire n_23069;
wire n_23070;
wire n_23071;
wire n_23072;
wire n_23073;
wire n_23074;
wire n_23075;
wire n_23076;
wire n_23077;
wire n_23078;
wire n_23079;
wire n_23080;
wire n_23081;
wire n_23082;
wire n_23083;
wire n_23084;
wire n_23085;
wire n_23086;
wire n_23087;
wire n_23088;
wire n_23089;
wire n_23090;
wire n_23091;
wire n_23092;
wire n_23093;
wire n_23094;
wire n_23095;
wire n_23096;
wire n_23097;
wire n_23098;
wire n_23099;
wire n_23100;
wire n_23101;
wire n_23102;
wire n_23103;
wire n_23104;
wire n_23105;
wire n_23106;
wire n_23107;
wire n_23108;
wire n_23109;
wire n_23110;
wire n_23111;
wire n_23112;
wire n_23113;
wire n_23114;
wire n_23115;
wire n_23116;
wire n_23117;
wire n_23118;
wire n_23119;
wire n_23120;
wire n_23121;
wire n_23122;
wire n_23123;
wire n_23124;
wire n_23125;
wire n_23126;
wire n_23127;
wire n_23128;
wire n_23129;
wire n_23130;
wire n_23131;
wire n_23132;
wire n_23133;
wire n_23134;
wire n_23135;
wire n_23136;
wire n_23137;
wire n_23138;
wire n_23139;
wire n_23140;
wire n_23141;
wire n_23142;
wire n_23143;
wire n_23144;
wire n_23145;
wire n_23146;
wire n_23147;
wire n_23148;
wire n_23149;
wire n_23150;
wire n_23151;
wire n_23152;
wire n_23153;
wire n_23154;
wire n_23155;
wire n_23156;
wire n_23157;
wire n_23158;
wire n_23159;
wire n_23160;
wire n_23161;
wire n_23162;
wire n_23163;
wire n_23164;
wire n_23165;
wire n_23166;
wire n_23167;
wire n_23168;
wire n_23169;
wire n_23170;
wire n_23171;
wire n_23172;
wire n_23173;
wire n_23174;
wire n_23175;
wire n_23176;
wire n_23177;
wire n_23178;
wire n_23179;
wire n_23180;
wire n_23181;
wire n_23182;
wire n_23183;
wire n_23184;
wire n_23185;
wire n_23186;
wire n_23187;
wire n_23188;
wire n_23189;
wire n_23190;
wire n_23191;
wire n_23192;
wire n_23193;
wire n_23194;
wire n_23195;
wire n_23196;
wire n_23197;
wire n_23198;
wire n_23199;
wire n_23200;
wire n_23201;
wire n_23202;
wire n_23203;
wire n_23204;
wire n_23205;
wire n_23206;
wire n_23207;
wire n_23208;
wire n_23209;
wire n_23210;
wire n_23211;
wire n_23212;
wire n_23213;
wire n_23214;
wire n_23215;
wire n_23216;
wire n_23217;
wire n_23218;
wire n_23219;
wire n_23220;
wire n_23221;
wire n_23222;
wire n_23223;
wire n_23224;
wire n_23225;
wire n_23226;
wire n_23227;
wire n_23228;
wire n_23229;
wire n_23230;
wire n_23231;
wire n_23232;
wire n_23233;
wire n_23234;
wire n_23235;
wire n_23236;
wire n_23237;
wire n_23238;
wire n_23239;
wire n_23240;
wire n_23241;
wire n_23242;
wire n_23243;
wire n_23244;
wire n_23245;
wire n_23246;
wire n_23247;
wire n_23248;
wire n_23249;
wire n_23250;
wire n_23251;
wire n_23252;
wire n_23253;
wire n_23254;
wire n_23255;
wire n_23256;
wire n_23257;
wire n_23258;
wire n_23259;
wire n_23260;
wire n_23261;
wire n_23262;
wire n_23263;
wire n_23264;
wire n_23265;
wire n_23266;
wire n_23267;
wire n_23268;
wire n_23269;
wire n_23270;
wire n_23271;
wire n_23272;
wire n_23273;
wire n_23274;
wire n_23275;
wire n_23276;
wire n_23277;
wire n_23278;
wire n_23279;
wire n_23280;
wire n_23281;
wire n_23282;
wire n_23283;
wire n_23284;
wire n_23285;
wire n_23286;
wire n_23287;
wire n_23288;
wire n_23289;
wire n_23290;
wire n_23291;
wire n_23292;
wire n_23293;
wire n_23294;
wire n_23295;
wire n_23296;
wire n_23297;
wire n_23298;
wire n_23299;
wire n_23300;
wire n_23301;
wire n_23302;
wire n_23303;
wire n_23304;
wire n_23305;
wire n_23306;
wire n_23307;
wire n_23308;
wire n_23309;
wire n_23310;
wire n_23311;
wire n_23312;
wire n_23313;
wire n_23314;
wire n_23315;
wire n_23316;
wire n_23317;
wire n_23318;
wire n_23319;
wire n_23320;
wire n_23321;
wire n_23322;
wire n_23323;
wire n_23324;
wire n_23325;
wire n_23326;
wire n_23327;
wire n_23328;
wire n_23329;
wire n_23330;
wire n_23331;
wire n_23332;
wire n_23333;
wire n_23334;
wire n_23335;
wire n_23336;
wire n_23337;
wire n_23338;
wire n_23339;
wire n_23340;
wire n_23341;
wire n_23342;
wire n_23343;
wire n_23344;
wire n_23345;
wire n_23346;
wire n_23347;
wire n_23348;
wire n_23349;
wire n_23350;
wire n_23351;
wire n_23352;
wire n_23353;
wire n_23354;
wire n_23355;
wire n_23356;
wire n_23357;
wire n_23358;
wire n_23359;
wire n_23360;
wire n_23361;
wire n_23362;
wire n_23363;
wire n_23364;
wire n_23365;
wire n_23366;
wire n_23367;
wire n_23368;
wire n_23369;
wire n_23370;
wire n_23371;
wire n_23372;
wire n_23373;
wire n_23374;
wire n_23375;
wire n_23376;
wire n_23377;
wire n_23378;
wire n_23379;
wire n_23380;
wire n_23381;
wire n_23382;
wire n_23383;
wire n_23384;
wire n_23385;
wire n_23386;
wire n_23387;
wire n_23388;
wire n_23389;
wire n_23390;
wire n_23391;
wire n_23392;
wire n_23393;
wire n_23394;
wire n_23395;
wire n_23396;
wire n_23397;
wire n_23398;
wire n_23399;
wire n_23400;
wire n_23401;
wire n_23402;
wire n_23403;
wire n_23404;
wire n_23405;
wire n_23406;
wire n_23407;
wire n_23408;
wire n_23409;
wire n_23410;
wire n_23411;
wire n_23412;
wire n_23413;
wire n_23414;
wire n_23415;
wire n_23416;
wire n_23417;
wire n_23418;
wire n_23419;
wire n_23420;
wire n_23421;
wire n_23422;
wire n_23423;
wire n_23424;
wire n_23425;
wire n_23426;
wire n_23427;
wire n_23428;
wire n_23429;
wire n_23430;
wire n_23431;
wire n_23432;
wire n_23433;
wire n_23434;
wire n_23435;
wire n_23436;
wire n_23437;
wire n_23438;
wire n_23439;
wire n_23440;
wire n_23441;
wire n_23442;
wire n_23443;
wire n_23444;
wire n_23445;
wire n_23446;
wire n_23447;
wire n_23448;
wire n_23449;
wire n_23450;
wire n_23451;
wire n_23452;
wire n_23453;
wire n_23454;
wire n_23455;
wire n_23456;
wire n_23457;
wire n_23458;
wire n_23459;
wire n_23460;
wire n_23461;
wire n_23462;
wire n_23463;
wire n_23464;
wire n_23465;
wire n_23466;
wire n_23467;
wire n_23468;
wire n_23469;
wire n_23470;
wire n_23471;
wire n_23472;
wire n_23473;
wire n_23474;
wire n_23475;
wire n_23476;
wire n_23477;
wire n_23478;
wire n_23479;
wire n_23480;
wire n_23481;
wire n_23482;
wire n_23483;
wire n_23484;
wire n_23485;
wire n_23486;
wire n_23487;
wire n_23488;
wire n_23489;
wire n_23490;
wire n_23491;
wire n_23492;
wire n_23493;
wire n_23494;
wire n_23495;
wire n_23496;
wire n_23497;
wire n_23498;
wire n_23499;
wire n_23500;
wire n_23501;
wire n_23502;
wire n_23503;
wire n_23504;
wire n_23505;
wire n_23506;
wire n_23507;
wire n_23508;
wire n_23509;
wire n_23510;
wire n_23511;
wire n_23512;
wire n_23513;
wire n_23514;
wire n_23515;
wire n_23516;
wire n_23517;
wire n_23518;
wire n_23519;
wire n_23520;
wire n_23521;
wire n_23522;
wire n_23523;
wire n_23524;
wire n_23525;
wire n_23526;
wire n_23527;
wire n_23528;
wire n_23529;
wire n_23530;
wire n_23531;
wire n_23532;
wire n_23533;
wire n_23534;
wire n_23535;
wire n_23536;
wire n_23537;
wire n_23538;
wire n_23539;
wire n_23540;
wire n_23541;
wire n_23542;
wire n_23543;
wire n_23544;
wire n_23545;
wire n_23546;
wire n_23547;
wire n_23548;
wire n_23549;
wire n_23550;
wire n_23551;
wire n_23552;
wire n_23553;
wire n_23554;
wire n_23555;
wire n_23556;
wire n_23557;
wire n_23558;
wire n_23559;
wire n_23560;
wire n_23561;
wire n_23562;
wire n_23563;
wire n_23564;
wire n_23565;
wire n_23566;
wire n_23567;
wire n_23568;
wire n_23569;
wire n_23570;
wire n_23571;
wire n_23572;
wire n_23573;
wire n_23574;
wire n_23575;
wire n_23576;
wire n_23577;
wire n_23578;
wire n_23579;
wire n_23580;
wire n_23581;
wire n_23582;
wire n_23583;
wire n_23584;
wire n_23585;
wire n_23586;
wire n_23587;
wire n_23588;
wire n_23589;
wire n_23590;
wire n_23591;
wire n_23592;
wire n_23593;
wire n_23594;
wire n_23595;
wire n_23596;
wire n_23597;
wire n_23598;
wire n_23599;
wire n_23600;
wire n_23601;
wire n_23602;
wire n_23603;
wire n_23604;
wire n_23605;
wire n_23606;
wire n_23607;
wire n_23608;
wire n_23609;
wire n_23610;
wire n_23611;
wire n_23612;
wire n_23613;
wire n_23614;
wire n_23615;
wire n_23616;
wire n_23617;
wire n_23618;
wire n_23619;
wire n_23620;
wire n_23621;
wire n_23622;
wire n_23623;
wire n_23624;
wire n_23625;
wire n_23626;
wire n_23627;
wire n_23628;
wire n_23629;
wire n_23630;
wire n_23631;
wire n_23632;
wire n_23633;
wire n_23634;
wire n_23635;
wire n_23636;
wire n_23637;
wire n_23638;
wire n_23639;
wire n_23640;
wire n_23641;
wire n_23642;
wire n_23643;
wire n_23644;
wire n_23645;
wire n_23646;
wire n_23647;
wire n_23648;
wire n_23649;
wire n_23650;
wire n_23651;
wire n_23652;
wire n_23653;
wire n_23654;
wire n_23655;
wire n_23656;
wire n_23657;
wire n_23658;
wire n_23659;
wire n_23660;
wire n_23661;
wire n_23662;
wire n_23663;
wire n_23664;
wire n_23665;
wire n_23666;
wire n_23667;
wire n_23668;
wire n_23669;
wire n_23670;
wire n_23671;
wire n_23672;
wire n_23673;
wire n_23674;
wire n_23675;
wire n_23676;
wire n_23677;
wire n_23678;
wire n_23679;
wire n_23680;
wire n_23681;
wire n_23682;
wire n_23683;
wire n_23684;
wire n_23685;
wire n_23686;
wire n_23687;
wire n_23688;
wire n_23689;
wire n_23690;
wire n_23691;
wire n_23692;
wire n_23693;
wire n_23694;
wire n_23695;
wire n_23696;
wire n_23697;
wire n_23698;
wire n_23699;
wire n_23700;
wire n_23701;
wire n_23702;
wire n_23703;
wire n_23704;
wire n_23705;
wire n_23706;
wire n_23707;
wire n_23708;
wire n_23709;
wire n_23710;
wire n_23711;
wire n_23712;
wire n_23713;
wire n_23714;
wire n_23715;
wire n_23716;
wire n_23717;
wire n_23718;
wire n_23719;
wire n_23720;
wire n_23721;
wire n_23722;
wire n_23723;
wire n_23724;
wire n_23725;
wire n_23726;
wire n_23727;
wire n_23728;
wire n_23729;
wire n_23730;
wire n_23731;
wire n_23732;
wire n_23733;
wire n_23734;
wire n_23735;
wire n_23736;
wire n_23737;
wire n_23738;
wire n_23739;
wire n_23740;
wire n_23741;
wire n_23742;
wire n_23743;
wire n_23744;
wire n_23745;
wire n_23746;
wire n_23747;
wire n_23748;
wire n_23749;
wire n_23750;
wire n_23751;
wire n_23752;
wire n_23753;
wire n_23754;
wire n_23755;
wire n_23756;
wire n_23757;
wire n_23758;
wire n_23759;
wire n_23760;
wire n_23761;
wire n_23762;
wire n_23763;
wire n_23764;
wire n_23765;
wire n_23766;
wire n_23767;
wire n_23768;
wire n_23769;
wire n_23770;
wire n_23771;
wire n_23772;
wire n_23773;
wire n_23774;
wire n_23775;
wire n_23776;
wire n_23777;
wire n_23778;
wire n_23779;
wire n_23780;
wire n_23781;
wire n_23782;
wire n_23783;
wire n_23784;
wire n_23785;
wire n_23786;
wire n_23787;
wire n_23788;
wire n_23789;
wire n_23790;
wire n_23791;
wire n_23792;
wire n_23793;
wire n_23794;
wire n_23795;
wire n_23796;
wire n_23797;
wire n_23798;
wire n_23799;
wire n_23800;
wire n_23801;
wire n_23802;
wire n_23803;
wire n_23804;
wire n_23805;
wire n_23806;
wire n_23807;
wire n_23808;
wire n_23809;
wire n_23810;
wire n_23811;
wire n_23812;
wire n_23813;
wire n_23814;
wire n_23815;
wire n_23816;
wire n_23817;
wire n_23818;
wire n_23819;
wire n_23820;
wire n_23821;
wire n_23822;
wire n_23823;
wire n_23824;
wire n_23825;
wire n_23826;
wire n_23827;
wire n_23828;
wire n_23829;
wire n_23830;
wire n_23831;
wire n_23832;
wire n_23833;
wire n_23834;
wire n_23835;
wire n_23836;
wire n_23837;
wire n_23838;
wire n_23839;
wire n_23840;
wire n_23841;
wire n_23842;
wire n_23843;
wire n_23844;
wire n_23845;
wire n_23846;
wire n_23847;
wire n_23848;
wire n_23849;
wire n_23850;
wire n_23851;
wire n_23852;
wire n_23853;
wire n_23854;
wire n_23855;
wire n_23856;
wire n_23857;
wire n_23858;
wire n_23859;
wire n_23860;
wire n_23861;
wire n_23862;
wire n_23863;
wire n_23864;
wire n_23865;
wire n_23866;
wire n_23867;
wire n_23868;
wire n_23869;
wire n_23870;
wire n_23871;
wire n_23872;
wire n_23873;
wire n_23874;
wire n_23875;
wire n_23876;
wire n_23877;
wire n_23878;
wire n_23879;
wire n_23880;
wire n_23881;
wire n_23882;
wire n_23883;
wire n_23884;
wire n_23885;
wire n_23886;
wire n_23887;
wire n_23888;
wire n_23889;
wire n_23890;
wire n_23891;
wire n_23892;
wire n_23893;
wire n_23894;
wire n_23895;
wire n_23896;
wire n_23897;
wire n_23898;
wire n_23899;
wire n_23900;
wire n_23901;
wire n_23902;
wire n_23903;
wire n_23904;
wire n_23905;
wire n_23906;
wire n_23907;
wire n_23908;
wire n_23909;
wire n_23910;
wire n_23911;
wire n_23912;
wire n_23913;
wire n_23914;
wire n_23915;
wire n_23916;
wire n_23917;
wire n_23918;
wire n_23919;
wire n_23920;
wire n_23921;
wire n_23922;
wire n_23923;
wire n_23924;
wire n_23925;
wire n_23926;
wire n_23927;
wire n_23928;
wire n_23929;
wire n_23930;
wire n_23931;
wire n_23932;
wire n_23933;
wire n_23934;
wire n_23935;
wire n_23936;
wire n_23937;
wire n_23938;
wire n_23939;
wire n_23940;
wire n_23941;
wire n_23942;
wire n_23943;
wire n_23944;
wire n_23945;
wire n_23946;
wire n_23947;
wire n_23948;
wire n_23949;
wire n_23950;
wire n_23951;
wire n_23952;
wire n_23953;
wire n_23954;
wire n_23955;
wire n_23956;
wire n_23957;
wire n_23958;
wire n_23959;
wire n_23960;
wire n_23961;
wire n_23962;
wire n_23963;
wire n_23964;
wire n_23965;
wire n_23966;
wire n_23967;
wire n_23968;
wire n_23969;
wire n_23970;
wire n_23971;
wire n_23972;
wire n_23973;
wire n_23974;
wire n_23975;
wire n_23976;
wire n_23977;
wire n_23978;
wire n_23979;
wire n_23980;
wire n_23981;
wire n_23982;
wire n_23983;
wire n_23984;
wire n_23985;
wire n_23986;
wire n_23987;
wire n_23988;
wire n_23989;
wire n_23990;
wire n_23991;
wire n_23992;
wire n_23993;
wire n_23994;
wire n_23995;
wire n_23996;
wire n_23997;
wire n_23998;
wire n_23999;
wire n_24000;
wire n_24001;
wire n_24002;
wire n_24003;
wire n_24004;
wire n_24005;
wire n_24006;
wire n_24007;
wire n_24008;
wire n_24009;
wire n_24010;
wire n_24011;
wire n_24012;
wire n_24013;
wire n_24014;
wire n_24015;
wire n_24016;
wire n_24017;
wire n_24018;
wire n_24019;
wire n_24020;
wire n_24021;
wire n_24022;
wire n_24023;
wire n_24024;
wire n_24025;
wire n_24026;
wire n_24027;
wire n_24028;
wire n_24029;
wire n_24030;
wire n_24031;
wire n_24032;
wire n_24033;
wire n_24034;
wire n_24035;
wire n_24036;
wire n_24037;
wire n_24038;
wire n_24039;
wire n_24040;
wire n_24041;
wire n_24042;
wire n_24043;
wire n_24044;
wire n_24045;
wire n_24046;
wire n_24047;
wire n_24048;
wire n_24049;
wire n_24050;
wire n_24051;
wire n_24052;
wire n_24053;
wire n_24054;
wire n_24055;
wire n_24056;
wire n_24057;
wire n_24058;
wire n_24059;
wire n_24060;
wire n_24061;
wire n_24062;
wire n_24063;
wire n_24064;
wire n_24065;
wire n_24066;
wire n_24067;
wire n_24068;
wire n_24069;
wire n_24070;
wire n_24071;
wire n_24072;
wire n_24073;
wire n_24074;
wire n_24075;
wire n_24076;
wire n_24077;
wire n_24078;
wire n_24079;
wire n_24080;
wire n_24081;
wire n_24082;
wire n_24083;
wire n_24084;
wire n_24085;
wire n_24086;
wire n_24087;
wire n_24088;
wire n_24089;
wire n_24090;
wire n_24091;
wire n_24092;
wire n_24093;
wire n_24094;
wire n_24095;
wire n_24096;
wire n_24097;
wire n_24098;
wire n_24099;
wire n_24100;
wire n_24101;
wire n_24102;
wire n_24103;
wire n_24104;
wire n_24105;
wire n_24106;
wire n_24107;
wire n_24108;
wire n_24109;
wire n_24110;
wire n_24111;
wire n_24112;
wire n_24113;
wire n_24114;
wire n_24115;
wire n_24116;
wire n_24117;
wire n_24118;
wire n_24119;
wire n_24120;
wire n_24121;
wire n_24122;
wire n_24123;
wire n_24124;
wire n_24125;
wire n_24126;
wire n_24127;
wire n_24128;
wire n_24129;
wire n_24130;
wire n_24131;
wire n_24132;
wire n_24133;
wire n_24134;
wire n_24135;
wire n_24136;
wire n_24137;
wire n_24138;
wire n_24139;
wire n_24140;
wire n_24141;
wire n_24142;
wire n_24143;
wire n_24144;
wire n_24145;
wire n_24146;
wire n_24147;
wire n_24148;
wire n_24149;
wire n_24150;
wire n_24151;
wire n_24152;
wire n_24153;
wire n_24154;
wire n_24155;
wire n_24156;
wire n_24157;
wire n_24158;
wire n_24159;
wire n_24160;
wire n_24161;
wire n_24162;
wire n_24163;
wire n_24164;
wire n_24165;
wire n_24166;
wire n_24167;
wire n_24168;
wire n_24169;
wire n_24170;
wire n_24171;
wire n_24172;
wire n_24173;
wire n_24174;
wire n_24175;
wire n_24176;
wire n_24177;
wire n_24178;
wire n_24179;
wire n_24180;
wire n_24181;
wire n_24182;
wire n_24183;
wire n_24184;
wire n_24185;
wire n_24186;
wire n_24187;
wire n_24188;
wire n_24189;
wire n_24190;
wire n_24191;
wire n_24192;
wire n_24193;
wire n_24194;
wire n_24195;
wire n_24196;
wire n_24197;
wire n_24198;
wire n_24199;
wire n_24200;
wire n_24201;
wire n_24202;
wire n_24203;
wire n_24204;
wire n_24205;
wire n_24206;
wire n_24207;
wire n_24208;
wire n_24209;
wire n_24210;
wire n_24211;
wire n_24212;
wire n_24213;
wire n_24214;
wire n_24215;
wire n_24216;
wire n_24217;
wire n_24218;
wire n_24219;
wire n_24220;
wire n_24221;
wire n_24222;
wire n_24223;
wire n_24224;
wire n_24225;
wire n_24226;
wire n_24227;
wire n_24228;
wire n_24229;
wire n_24230;
wire n_24231;
wire n_24232;
wire n_24233;
wire n_24234;
wire n_24235;
wire n_24236;
wire n_24237;
wire n_24238;
wire n_24239;
wire n_24240;
wire n_24241;
wire n_24242;
wire n_24243;
wire n_24244;
wire n_24245;
wire n_24246;
wire n_24247;
wire n_24248;
wire n_24249;
wire n_24250;
wire n_24251;
wire n_24252;
wire n_24253;
wire n_24254;
wire n_24255;
wire n_24256;
wire n_24257;
wire n_24258;
wire n_24259;
wire n_24260;
wire n_24261;
wire n_24262;
wire n_24263;
wire n_24264;
wire n_24265;
wire n_24266;
wire n_24267;
wire n_24268;
wire n_24269;
wire n_24270;
wire n_24271;
wire n_24272;
wire n_24273;
wire n_24274;
wire n_24275;
wire n_24276;
wire n_24277;
wire n_24278;
wire n_24279;
wire n_24280;
wire n_24281;
wire n_24282;
wire n_24283;
wire n_24284;
wire n_24285;
wire n_24286;
wire n_24287;
wire n_24288;
wire n_24289;
wire n_24290;
wire n_24291;
wire n_24292;
wire n_24293;
wire n_24294;
wire n_24295;
wire n_24296;
wire n_24297;
wire n_24298;
wire n_24299;
wire n_24300;
wire n_24301;
wire n_24302;
wire n_24303;
wire n_24304;
wire n_24305;
wire n_24306;
wire n_24307;
wire n_24308;
wire n_24309;
wire n_24310;
wire n_24311;
wire n_24312;
wire n_24313;
wire n_24314;
wire n_24315;
wire n_24316;
wire n_24317;
wire n_24318;
wire n_24319;
wire n_24320;
wire n_24321;
wire n_24322;
wire n_24323;
wire n_24324;
wire n_24325;
wire n_24326;
wire n_24327;
wire n_24328;
wire n_24329;
wire n_24330;
wire n_24331;
wire n_24332;
wire n_24333;
wire n_24334;
wire n_24335;
wire n_24336;
wire n_24337;
wire n_24338;
wire n_24339;
wire n_24340;
wire n_24341;
wire n_24342;
wire n_24343;
wire n_24344;
wire n_24345;
wire n_24346;
wire n_24347;
wire n_24348;
wire n_24349;
wire n_24350;
wire n_24351;
wire n_24352;
wire n_24353;
wire n_24354;
wire n_24355;
wire n_24356;
wire n_24357;
wire n_24358;
wire n_24359;
wire n_24360;
wire n_24361;
wire n_24362;
wire n_24363;
wire n_24364;
wire n_24365;
wire n_24366;
wire n_24367;
wire n_24368;
wire n_24369;
wire n_24370;
wire n_24371;
wire n_24372;
wire n_24373;
wire n_24374;
wire n_24375;
wire n_24376;
wire n_24377;
wire n_24378;
wire n_24379;
wire n_24380;
wire n_24381;
wire n_24382;
wire n_24383;
wire n_24384;
wire n_24385;
wire n_24386;
wire n_24387;
wire n_24388;
wire n_24389;
wire n_24390;
wire n_24391;
wire n_24392;
wire n_24393;
wire n_24394;
wire n_24395;
wire n_24396;
wire n_24397;
wire n_24398;
wire n_24399;
wire n_24400;
wire n_24401;
wire n_24402;
wire n_24403;
wire n_24404;
wire n_24405;
wire n_24406;
wire n_24407;
wire n_24408;
wire n_24409;
wire n_24410;
wire n_24411;
wire n_24412;
wire n_24413;
wire n_24414;
wire n_24415;
wire n_24416;
wire n_24417;
wire n_24418;
wire n_24419;
wire n_24420;
wire n_24421;
wire n_24422;
wire n_24423;
wire n_24424;
wire n_24425;
wire n_24426;
wire n_24427;
wire n_24428;
wire n_24429;
wire n_24430;
wire n_24431;
wire n_24432;
wire n_24433;
wire n_24434;
wire n_24435;
wire n_24436;
wire n_24437;
wire n_24438;
wire n_24439;
wire n_24440;
wire n_24441;
wire n_24442;
wire n_24443;
wire n_24444;
wire n_24445;
wire n_24446;
wire n_24447;
wire n_24448;
wire n_24449;
wire n_24450;
wire n_24451;
wire n_24452;
wire n_24453;
wire n_24454;
wire n_24455;
wire n_24456;
wire n_24457;
wire n_24458;
wire n_24459;
wire n_24460;
wire n_24461;
wire n_24462;
wire n_24463;
wire n_24464;
wire n_24465;
wire n_24466;
wire n_24467;
wire n_24468;
wire n_24469;
wire n_24470;
wire n_24471;
wire n_24472;
wire n_24473;
wire n_24474;
wire n_24475;
wire n_24476;
wire n_24477;
wire n_24478;
wire n_24479;
wire n_24480;
wire n_24481;
wire n_24482;
wire n_24483;
wire n_24484;
wire n_24485;
wire n_24486;
wire n_24487;
wire n_24488;
wire n_24489;
wire n_24490;
wire n_24491;
wire n_24492;
wire n_24493;
wire n_24494;
wire n_24495;
wire n_24496;
wire n_24497;
wire n_24498;
wire n_24499;
wire n_24500;
wire n_24501;
wire n_24502;
wire n_24503;
wire n_24504;
wire n_24505;
wire n_24506;
wire n_24507;
wire n_24508;
wire n_24509;
wire n_24510;
wire n_24511;
wire n_24512;
wire n_24513;
wire n_24514;
wire n_24515;
wire n_24516;
wire n_24517;
wire n_24518;
wire n_24519;
wire n_24520;
wire n_24521;
wire n_24522;
wire n_24523;
wire n_24524;
wire n_24525;
wire n_24526;
wire n_24527;
wire n_24528;
wire n_24529;
wire n_24530;
wire n_24531;
wire n_24532;
wire n_24533;
wire n_24534;
wire n_24535;
wire n_24536;
wire n_24537;
wire n_24538;
wire n_24539;
wire n_24540;
wire n_24541;
wire n_24542;
wire n_24543;
wire n_24544;
wire n_24545;
wire n_24546;
wire n_24547;
wire n_24548;
wire n_24549;
wire n_24550;
wire n_24551;
wire n_24552;
wire n_24553;
wire n_24554;
wire n_24555;
wire n_24556;
wire n_24557;
wire n_24558;
wire n_24559;
wire n_24560;
wire n_24561;
wire n_24562;
wire n_24563;
wire n_24564;
wire n_24565;
wire n_24566;
wire n_24567;
wire n_24568;
wire n_24569;
wire n_24570;
wire n_24571;
wire n_24572;
wire n_24573;
wire n_24574;
wire n_24575;
wire n_24576;
wire n_24577;
wire n_24578;
wire n_24579;
wire n_24580;
wire n_24581;
wire n_24582;
wire n_24583;
wire n_24584;
wire n_24585;
wire n_24586;
wire n_24587;
wire n_24588;
wire n_24589;
wire n_24590;
wire n_24591;
wire n_24592;
wire n_24593;
wire n_24594;
wire n_24595;
wire n_24596;
wire n_24597;
wire n_24598;
wire n_24599;
wire n_24600;
wire n_24601;
wire n_24602;
wire n_24603;
wire n_24604;
wire n_24605;
wire n_24606;
wire n_24607;
wire n_24608;
wire n_24609;
wire n_24610;
wire n_24611;
wire n_24612;
wire n_24613;
wire n_24614;
wire n_24615;
wire n_24616;
wire n_24617;
wire n_24618;
wire n_24619;
wire n_24620;
wire n_24621;
wire n_24622;
wire n_24623;
wire n_24624;
wire n_24625;
wire n_24626;
wire n_24627;
wire n_24628;
wire n_24629;
wire n_24630;
wire n_24631;
wire n_24632;
wire n_24633;
wire n_24634;
wire n_24635;
wire n_24636;
wire n_24637;
wire n_24638;
wire n_24639;
wire n_24640;
wire n_24641;
wire n_24642;
wire n_24643;
wire n_24644;
wire n_24645;
wire n_24646;
wire n_24647;
wire n_24648;
wire n_24649;
wire n_24650;
wire n_24651;
wire n_24652;
wire n_24653;
wire n_24654;
wire n_24655;
wire n_24656;
wire n_24657;
wire n_24658;
wire n_24659;
wire n_24660;
wire n_24661;
wire n_24662;
wire n_24663;
wire n_24664;
wire n_24665;
wire n_24666;
wire n_24667;
wire n_24668;
wire n_24669;
wire n_24670;
wire n_24671;
wire n_24672;
wire n_24673;
wire n_24674;
wire n_24675;
wire n_24676;
wire n_24677;
wire n_24678;
wire n_24679;
wire n_24680;
wire n_24681;
wire n_24682;
wire n_24683;
wire n_24684;
wire n_24685;
wire n_24686;
wire n_24687;
wire n_24688;
wire n_24689;
wire n_24690;
wire n_24691;
wire n_24692;
wire n_24693;
wire n_24694;
wire n_24695;
wire n_24696;
wire n_24697;
wire n_24698;
wire n_24699;
wire n_24700;
wire n_24701;
wire n_24702;
wire n_24703;
wire n_24704;
wire n_24705;
wire n_24706;
wire n_24707;
wire n_24708;
wire n_24709;
wire n_24710;
wire n_24711;
wire n_24712;
wire n_24713;
wire n_24714;
wire n_24715;
wire n_24716;
wire n_24717;
wire n_24718;
wire n_24719;
wire n_24720;
wire n_24721;
wire n_24722;
wire n_24723;
wire n_24724;
wire n_24725;
wire n_24726;
wire n_24727;
wire n_24728;
wire n_24729;
wire n_24730;
wire n_24731;
wire n_24732;
wire n_24733;
wire n_24734;
wire n_24735;
wire n_24736;
wire n_24737;
wire n_24738;
wire n_24739;
wire n_24740;
wire n_24741;
wire n_24742;
wire n_24743;
wire n_24744;
wire n_24745;
wire n_24746;
wire n_24747;
wire n_24748;
wire n_24749;
wire n_24750;
wire n_24751;
wire n_24752;
wire n_24753;
wire n_24754;
wire n_24755;
wire n_24756;
wire n_24757;
wire n_24758;
wire n_24759;
wire n_24760;
wire n_24761;
wire n_24762;
wire n_24763;
wire n_24764;
wire n_24765;
wire n_24766;
wire n_24767;
wire n_24768;
wire n_24769;
wire n_24770;
wire n_24771;
wire n_24772;
wire n_24773;
wire n_24774;
wire n_24775;
wire n_24776;
wire n_24777;
wire n_24778;
wire n_24779;
wire n_24780;
wire n_24781;
wire n_24782;
wire n_24783;
wire n_24784;
wire n_24785;
wire n_24786;
wire n_24787;
wire n_24788;
wire n_24789;
wire n_24790;
wire n_24791;
wire n_24792;
wire n_24793;
wire n_24794;
wire n_24795;
wire n_24796;
wire n_24797;
wire n_24798;
wire n_24799;
wire n_24800;
wire n_24801;
wire n_24802;
wire n_24803;
wire n_24804;
wire n_24805;
wire n_24806;
wire n_24807;
wire n_24808;
wire n_24809;
wire n_24810;
wire n_24811;
wire n_24812;
wire n_24813;
wire n_24814;
wire n_24815;
wire n_24816;
wire n_24817;
wire n_24818;
wire n_24819;
wire n_24820;
wire n_24821;
wire n_24822;
wire n_24823;
wire n_24824;
wire n_24825;
wire n_24826;
wire n_24827;
wire n_24828;
wire n_24829;
wire n_24830;
wire n_24831;
wire n_24832;
wire n_24833;
wire n_24834;
wire n_24835;
wire n_24836;
wire n_24837;
wire n_24838;
wire n_24839;
wire n_24840;
wire n_24841;
wire n_24842;
wire n_24843;
wire n_24844;
wire n_24845;
wire n_24846;
wire n_24847;
wire n_24848;
wire n_24849;
wire n_24850;
wire n_24851;
wire n_24852;
wire n_24853;
wire n_24854;
wire n_24855;
wire n_24856;
wire n_24857;
wire n_24858;
wire n_24859;
wire n_24860;
wire n_24861;
wire n_24862;
wire n_24863;
wire n_24864;
wire n_24865;
wire n_24866;
wire n_24867;
wire n_24868;
wire n_24869;
wire n_24870;
wire n_24871;
wire n_24872;
wire n_24873;
wire n_24874;
wire n_24875;
wire n_24876;
wire n_24877;
wire n_24878;
wire n_24879;
wire n_24880;
wire n_24881;
wire n_24882;
wire n_24883;
wire n_24884;
wire n_24885;
wire n_24886;
wire n_24887;
wire n_24888;
wire n_24889;
wire n_24890;
wire n_24891;
wire n_24892;
wire n_24893;
wire n_24894;
wire n_24895;
wire n_24896;
wire n_24897;
wire n_24898;
wire n_24899;
wire n_24900;
wire n_24901;
wire n_24902;
wire n_24903;
wire n_24904;
wire n_24905;
wire n_24906;
wire n_24907;
wire n_24908;
wire n_24909;
wire n_24910;
wire n_24911;
wire n_24912;
wire n_24913;
wire n_24914;
wire n_24915;
wire n_24916;
wire n_24917;
wire n_24918;
wire n_24919;
wire n_24920;
wire n_24921;
wire n_24922;
wire n_24923;
wire n_24924;
wire n_24925;
wire n_24926;
wire n_24927;
wire n_24928;
wire n_24929;
wire n_24930;
wire n_24931;
wire n_24932;
wire n_24933;
wire n_24934;
wire n_24935;
wire n_24936;
wire n_24937;
wire n_24938;
wire n_24939;
wire n_24940;
wire n_24941;
wire n_24942;
wire n_24943;
wire n_24944;
wire n_24945;
wire n_24946;
wire n_24947;
wire n_24948;
wire n_24949;
wire n_24950;
wire n_24951;
wire n_24952;
wire n_24953;
wire n_24954;
wire n_24955;
wire n_24956;
wire n_24957;
wire n_24958;
wire n_24959;
wire n_24960;
wire n_24961;
wire n_24962;
wire n_24963;
wire n_24964;
wire n_24965;
wire n_24966;
wire n_24967;
wire n_24968;
wire n_24969;
wire n_24970;
wire n_24971;
wire n_24972;
wire n_24973;
wire n_24974;
wire n_24975;
wire n_24976;
wire n_24977;
wire n_24978;
wire n_24979;
wire n_24980;
wire n_24981;
wire n_24982;
wire n_24983;
wire n_24984;
wire n_24985;
wire n_24986;
wire n_24987;
wire n_24988;
wire n_24989;
wire n_24990;
wire n_24991;
wire n_24992;
wire n_24993;
wire n_24994;
wire n_24995;
wire n_24996;
wire n_24997;
wire n_24998;
wire n_24999;
wire n_25000;
wire n_25001;
wire n_25002;
wire n_25003;
wire n_25004;
wire n_25005;
wire n_25006;
wire n_25007;
wire n_25008;
wire n_25009;
wire n_25010;
wire n_25011;
wire n_25012;
wire n_25013;
wire n_25014;
wire n_25015;
wire n_25016;
wire n_25017;
wire n_25018;
wire n_25019;
wire n_25020;
wire n_25021;
wire n_25022;
wire n_25023;
wire n_25024;
wire n_25025;
wire n_25026;
wire n_25027;
wire n_25028;
wire n_25029;
wire n_25030;
wire n_25031;
wire n_25032;
wire n_25033;
wire n_25034;
wire n_25035;
wire n_25036;
wire n_25037;
wire n_25038;
wire n_25039;
wire n_25040;
wire n_25041;
wire n_25042;
wire n_25043;
wire n_25044;
wire n_25045;
wire n_25046;
wire n_25047;
wire n_25048;
wire n_25049;
wire n_25050;
wire n_25051;
wire n_25052;
wire n_25053;
wire n_25054;
wire n_25055;
wire n_25056;
wire n_25057;
wire n_25058;
wire n_25059;
wire n_25060;
wire n_25061;
wire n_25062;
wire n_25063;
wire n_25064;
wire n_25065;
wire n_25066;
wire n_25067;
wire n_25068;
wire n_25069;
wire n_25070;
wire n_25071;
wire n_25072;
wire n_25073;
wire n_25074;
wire n_25075;
wire n_25076;
wire n_25077;
wire n_25078;
wire n_25079;
wire n_25080;
wire n_25081;
wire n_25082;
wire n_25083;
wire n_25084;
wire n_25085;
wire n_25086;
wire n_25087;
wire n_25088;
wire n_25089;
wire n_25090;
wire n_25091;
wire n_25092;
wire n_25093;
wire n_25094;
wire n_25095;
wire n_25096;
wire n_25097;
wire n_25098;
wire n_25099;
wire n_25100;
wire n_25101;
wire n_25102;
wire n_25103;
wire n_25104;
wire n_25105;
wire n_25106;
wire n_25107;
wire n_25108;
wire n_25109;
wire n_25110;
wire n_25111;
wire n_25112;
wire n_25113;
wire n_25114;
wire n_25115;
wire n_25116;
wire n_25117;
wire n_25118;
wire n_25119;
wire n_25120;
wire n_25121;
wire n_25122;
wire n_25123;
wire n_25124;
wire n_25125;
wire n_25126;
wire n_25127;
wire n_25128;
wire n_25129;
wire n_25130;
wire n_25131;
wire n_25132;
wire n_25133;
wire n_25134;
wire n_25135;
wire n_25136;
wire n_25137;
wire n_25138;
wire n_25139;
wire n_25140;
wire n_25141;
wire n_25142;
wire n_25143;
wire n_25144;
wire n_25145;
wire n_25146;
wire n_25147;
wire n_25148;
wire n_25149;
wire n_25150;
wire n_25151;
wire n_25152;
wire n_25153;
wire n_25154;
wire n_25155;
wire n_25156;
wire n_25157;
wire n_25158;
wire n_25159;
wire n_25160;
wire n_25161;
wire n_25162;
wire n_25163;
wire n_25164;
wire n_25165;
wire n_25166;
wire n_25167;
wire n_25168;
wire n_25169;
wire n_25170;
wire n_25171;
wire n_25172;
wire n_25173;
wire n_25174;
wire n_25175;
wire n_25176;
wire n_25177;
wire n_25178;
wire n_25179;
wire n_25180;
wire n_25181;
wire n_25182;
wire n_25183;
wire n_25184;
wire n_25185;
wire n_25186;
wire n_25187;
wire n_25188;
wire n_25189;
wire n_25190;
wire n_25191;
wire n_25192;
wire n_25193;
wire n_25194;
wire n_25195;
wire n_25196;
wire n_25197;
wire n_25198;
wire n_25199;
wire n_25200;
wire n_25201;
wire n_25202;
wire n_25203;
wire n_25204;
wire n_25205;
wire n_25206;
wire n_25207;
wire n_25208;
wire n_25209;
wire n_25210;
wire n_25211;
wire n_25212;
wire n_25213;
wire n_25214;
wire n_25215;
wire n_25216;
wire n_25217;
wire n_25218;
wire n_25219;
wire n_25220;
wire n_25221;
wire n_25222;
wire n_25223;
wire n_25224;
wire n_25225;
wire n_25226;
wire n_25227;
wire n_25228;
wire n_25229;
wire n_25230;
wire n_25231;
wire n_25232;
wire n_25233;
wire n_25234;
wire n_25235;
wire n_25236;
wire n_25237;
wire n_25238;
wire n_25239;
wire n_25240;
wire n_25241;
wire n_25242;
wire n_25243;
wire n_25244;
wire n_25245;
wire n_25246;
wire n_25247;
wire n_25248;
wire n_25249;
wire n_25250;
wire n_25251;
wire n_25252;
wire n_25253;
wire n_25254;
wire n_25255;
wire n_25256;
wire n_25257;
wire n_25258;
wire n_25259;
wire n_25260;
wire n_25261;
wire n_25262;
wire n_25263;
wire n_25264;
wire n_25265;
wire n_25266;
wire n_25267;
wire n_25268;
wire n_25269;
wire n_25270;
wire n_25271;
wire n_25272;
wire n_25273;
wire n_25274;
wire n_25275;
wire n_25276;
wire n_25277;
wire n_25278;
wire n_25279;
wire n_25280;
wire n_25281;
wire n_25282;
wire n_25283;
wire n_25284;
wire n_25285;
wire n_25286;
wire n_25287;
wire n_25288;
wire n_25289;
wire n_25290;
wire n_25291;
wire n_25292;
wire n_25293;
wire n_25294;
wire n_25295;
wire n_25296;
wire n_25297;
wire n_25298;
wire n_25299;
wire n_25300;
wire n_25301;
wire n_25302;
wire n_25303;
wire n_25304;
wire n_25305;
wire n_25306;
wire n_25307;
wire n_25308;
wire n_25309;
wire n_25310;
wire n_25311;
wire n_25312;
wire n_25313;
wire n_25314;
wire n_25315;
wire n_25316;
wire n_25317;
wire n_25318;
wire n_25319;
wire n_25320;
wire n_25321;
wire n_25322;
wire n_25323;
wire n_25324;
wire n_25325;
wire n_25326;
wire n_25327;
wire n_25328;
wire n_25329;
wire n_25330;
wire n_25331;
wire n_25332;
wire n_25333;
wire n_25334;
wire n_25335;
wire n_25336;
wire n_25337;
wire n_25338;
wire n_25339;
wire n_25340;
wire n_25341;
wire n_25342;
wire n_25343;
wire n_25344;
wire n_25345;
wire n_25346;
wire n_25347;
wire n_25348;
wire n_25349;
wire n_25350;
wire n_25351;
wire n_25352;
wire n_25353;
wire n_25354;
wire n_25355;
wire n_25356;
wire n_25357;
wire n_25358;
wire n_25359;
wire n_25360;
wire n_25361;
wire n_25362;
wire n_25363;
wire n_25364;
wire n_25365;
wire n_25366;
wire n_25367;
wire n_25368;
wire n_25369;
wire n_25370;
wire n_25371;
wire n_25372;
wire n_25373;
wire n_25374;
wire n_25375;
wire n_25376;
wire n_25377;
wire n_25378;
wire n_25379;
wire n_25380;
wire n_25381;
wire n_25382;
wire n_25383;
wire n_25384;
wire n_25385;
wire n_25386;
wire n_25387;
wire n_25388;
wire n_25389;
wire n_25390;
wire n_25391;
wire n_25392;
wire n_25393;
wire n_25394;
wire n_25395;
wire n_25396;
wire n_25397;
wire n_25398;
wire n_25399;
wire n_25400;
wire n_25401;
wire n_25402;
wire n_25403;
wire n_25404;
wire n_25405;
wire n_25406;
wire n_25407;
wire n_25408;
wire n_25409;
wire n_25410;
wire n_25411;
wire n_25412;
wire n_25413;
wire n_25414;
wire n_25415;
wire n_25416;
wire n_25417;
wire n_25418;
wire n_25419;
wire n_25420;
wire n_25421;
wire n_25422;
wire n_25423;
wire n_25424;
wire n_25425;
wire n_25426;
wire n_25427;
wire n_25428;
wire n_25429;
wire n_25430;
wire n_25431;
wire n_25432;
wire n_25433;
wire n_25434;
wire n_25435;
wire n_25436;
wire n_25437;
wire n_25438;
wire n_25439;
wire n_25440;
wire n_25441;
wire n_25442;
wire n_25443;
wire n_25444;
wire n_25445;
wire n_25446;
wire n_25447;
wire n_25448;
wire n_25449;
wire n_25450;
wire n_25451;
wire n_25452;
wire n_25453;
wire n_25454;
wire n_25455;
wire n_25456;
wire n_25457;
wire n_25458;
wire n_25459;
wire n_25460;
wire n_25461;
wire n_25462;
wire n_25463;
wire n_25464;
wire n_25465;
wire n_25466;
wire n_25467;
wire n_25468;
wire n_25469;
wire n_25470;
wire n_25471;
wire n_25472;
wire n_25473;
wire n_25474;
wire n_25475;
wire n_25476;
wire n_25477;
wire n_25478;
wire n_25479;
wire n_25480;
wire n_25481;
wire n_25482;
wire n_25483;
wire n_25484;
wire n_25485;
wire n_25486;
wire n_25487;
wire n_25488;
wire n_25489;
wire n_25490;
wire n_25491;
wire n_25492;
wire n_25493;
wire n_25494;
wire n_25495;
wire n_25496;
wire n_25497;
wire n_25498;
wire n_25499;
wire n_25500;
wire n_25501;
wire n_25502;
wire n_25503;
wire n_25504;
wire n_25505;
wire n_25506;
wire n_25507;
wire n_25508;
wire n_25509;
wire n_25510;
wire n_25511;
wire n_25512;
wire n_25513;
wire n_25514;
wire n_25515;
wire n_25516;
wire n_25517;
wire n_25518;
wire n_25519;
wire n_25520;
wire n_25521;
wire n_25522;
wire n_25523;
wire n_25524;
wire n_25525;
wire n_25526;
wire n_25527;
wire n_25528;
wire n_25529;
wire n_25530;
wire n_25531;
wire n_25532;
wire n_25533;
wire n_25534;
wire n_25535;
wire n_25536;
wire n_25537;
wire n_25538;
wire n_25539;
wire n_25540;
wire n_25541;
wire n_25542;
wire n_25543;
wire n_25544;
wire n_25545;
wire n_25546;
wire n_25547;
wire n_25548;
wire n_25549;
wire n_25550;
wire n_25551;
wire n_25552;
wire n_25553;
wire n_25554;
wire n_25555;
wire n_25556;
wire n_25557;
wire n_25558;
wire n_25559;
wire n_25560;
wire n_25561;
wire n_25562;
wire n_25563;
wire n_25564;
wire n_25565;
wire n_25566;
wire n_25567;
wire n_25568;
wire n_25569;
wire n_25570;
wire n_25571;
wire n_25572;
wire n_25573;
wire n_25574;
wire n_25575;
wire n_25576;
wire n_25577;
wire n_25578;
wire n_25579;
wire n_25580;
wire n_25581;
wire n_25582;
wire n_25583;
wire n_25584;
wire n_25585;
wire n_25586;
wire n_25587;
wire n_25588;
wire n_25589;
wire n_25590;
wire n_25591;
wire n_25592;
wire n_25593;
wire n_25594;
wire n_25595;
wire n_25596;
wire n_25597;
wire n_25598;
wire n_25599;
wire n_25600;
wire n_25601;
wire n_25602;
wire n_25603;
wire n_25604;
wire n_25605;
wire n_25606;
wire n_25607;
wire n_25608;
wire n_25609;
wire n_25610;
wire n_25611;
wire n_25612;
wire n_25613;
wire n_25614;
wire n_25615;
wire n_25616;
wire n_25617;
wire n_25618;
wire n_25619;
wire n_25620;
wire n_25621;
wire n_25622;
wire n_25623;
wire n_25624;
wire n_25625;
wire n_25626;
wire n_25627;
wire n_25628;
wire n_25629;
wire n_25630;
wire n_25631;
wire n_25632;
wire n_25633;
wire n_25634;
wire n_25635;
wire n_25636;
wire n_25637;
wire n_25638;
wire n_25639;
wire n_25640;
wire n_25641;
wire n_25642;
wire n_25643;
wire n_25644;
wire n_25645;
wire n_25646;
wire n_25647;
wire n_25648;
wire n_25649;
wire n_25650;
wire n_25651;
wire n_25652;
wire n_25653;
wire n_25654;
wire n_25655;
wire n_25656;
wire n_25657;
wire n_25658;
wire n_25659;
wire n_25660;
wire n_25661;
wire n_25662;
wire n_25663;
wire n_25664;
wire n_25665;
wire n_25666;
wire n_25667;
wire n_25668;
wire n_25669;
wire n_25670;
wire n_25671;
wire n_25672;
wire n_25673;
wire n_25674;
wire n_25675;
wire n_25676;
wire n_25677;
wire n_25678;
wire n_25679;
wire n_25680;
wire n_25681;
wire n_25682;
wire n_25683;
wire n_25684;
wire n_25685;
wire n_25686;
wire n_25687;
wire n_25688;
wire n_25689;
wire n_25690;
wire n_25691;
wire n_25692;
wire n_25693;
wire n_25694;
wire n_25695;
wire n_25696;
wire n_25697;
wire n_25698;
wire n_25699;
wire n_25700;
wire n_25701;
wire n_25702;
wire n_25703;
wire n_25704;
wire n_25705;
wire n_25706;
wire n_25707;
wire n_25708;
wire n_25709;
wire n_25710;
wire n_25711;
wire n_25712;
wire n_25713;
wire n_25714;
wire n_25715;
wire n_25716;
wire n_25717;
wire n_25718;
wire n_25719;
wire n_25720;
wire n_25721;
wire n_25722;
wire n_25723;
wire n_25724;
wire n_25725;
wire n_25726;
wire n_25727;
wire n_25728;
wire n_25729;
wire n_25730;
wire n_25731;
wire n_25732;
wire n_25733;
wire n_25734;
wire n_25735;
wire n_25736;
wire n_25737;
wire n_25738;
wire n_25739;
wire n_25740;
wire n_25741;
wire n_25742;
wire n_25743;
wire n_25744;
wire n_25745;
wire n_25746;
wire n_25747;
wire n_25748;
wire n_25749;
wire n_25750;
wire n_25751;
wire n_25752;
wire n_25753;
wire n_25754;
wire n_25755;
wire n_25756;
wire n_25757;
wire n_25758;
wire n_25759;
wire n_25760;
wire n_25761;
wire n_25762;
wire n_25763;
wire n_25764;
wire n_25765;
wire n_25766;
wire n_25767;
wire n_25768;
wire n_25769;
wire n_25770;
wire n_25771;
wire n_25772;
wire n_25773;
wire n_25774;
wire n_25775;
wire n_25776;
wire n_25777;
wire n_25778;
wire n_25779;
wire n_25780;
wire n_25781;
wire n_25782;
wire n_25783;
wire n_25784;
wire n_25785;
wire n_25786;
wire n_25787;
wire n_25788;
wire n_25789;
wire n_25790;
wire n_25791;
wire n_25792;
wire n_25793;
wire n_25794;
wire n_25795;
wire n_25796;
wire n_25797;
wire n_25798;
wire n_25799;
wire n_25800;
wire n_25801;
wire n_25802;
wire n_25803;
wire n_25804;
wire n_25805;
wire n_25806;
wire n_25807;
wire n_25808;
wire n_25809;
wire n_25810;
wire n_25811;
wire n_25812;
wire n_25813;
wire n_25814;
wire n_25815;
wire n_25816;
wire n_25817;
wire n_25818;
wire n_25819;
wire n_25820;
wire n_25821;
wire n_25822;
wire n_25823;
wire n_25824;
wire n_25825;
wire n_25826;
wire n_25827;
wire n_25828;
wire n_25829;
wire n_25830;
wire n_25831;
wire n_25832;
wire n_25833;
wire n_25834;
wire n_25835;
wire n_25836;
wire n_25837;
wire n_25838;
wire n_25839;
wire n_25840;
wire n_25841;
wire n_25842;
wire n_25843;
wire n_25844;
wire n_25845;
wire n_25846;
wire n_25847;
wire n_25848;
wire n_25849;
wire n_25850;
wire n_25851;
wire n_25852;
wire n_25853;
wire n_25854;
wire n_25855;
wire n_25856;
wire n_25857;
wire n_25858;
wire n_25859;
wire n_25860;
wire n_25861;
wire n_25862;
wire n_25863;
wire n_25864;
wire n_25865;
wire n_25866;
wire n_25867;
wire n_25868;
wire n_25869;
wire n_25870;
wire n_25871;
wire n_25872;
wire n_25873;
wire n_25874;
wire n_25875;
wire n_25876;
wire n_25877;
wire n_25878;
wire n_25879;
wire n_25880;
wire n_25881;
wire n_25882;
wire n_25883;
wire n_25884;
wire n_25885;
wire n_25886;
wire n_25887;
wire n_25888;
wire n_25889;
wire n_25890;
wire n_25891;
wire n_25892;
wire n_25893;
wire n_25894;
wire n_25895;
wire n_25896;
wire n_25897;
wire n_25898;
wire n_25899;
wire n_25900;
wire n_25901;
wire n_25902;
wire n_25903;
wire n_25904;
wire n_25905;
wire n_25906;
wire n_25907;
wire n_25908;
wire n_25909;
wire n_25910;
wire n_25911;
wire n_25912;
wire n_25913;
wire n_25914;
wire n_25915;
wire n_25916;
wire n_25917;
wire n_25918;
wire n_25919;
wire n_25920;
wire n_25921;
wire n_25922;
wire n_25923;
wire n_25924;
wire n_25925;
wire n_25926;
wire n_25927;
wire n_25928;
wire n_25929;
wire n_25930;
wire n_25931;
wire n_25932;
wire n_25933;
wire n_25934;
wire n_25935;
wire n_25936;
wire n_25937;
wire n_25938;
wire n_25939;
wire n_25940;
wire n_25941;
wire n_25942;
wire n_25943;
wire n_25944;
wire n_25945;
wire n_25946;
wire n_25947;
wire n_25948;
wire n_25949;
wire n_25950;
wire n_25951;
wire n_25952;
wire n_25953;
wire n_25954;
wire n_25955;
wire n_25956;
wire n_25957;
wire n_25958;
wire n_25959;
wire n_25960;
wire n_25961;
wire n_25962;
wire n_25963;
wire n_25964;
wire n_25965;
wire n_25966;
wire n_25967;
wire n_25968;
wire n_25969;
wire n_25970;
wire n_25971;
wire n_25972;
wire n_25973;
wire n_25974;
wire n_25975;
wire n_25976;
wire n_25977;
wire n_25978;
wire n_25979;
wire n_25980;
wire n_25981;
wire n_25982;
wire n_25983;
wire n_25984;
wire n_25985;
wire n_25986;
wire n_25987;
wire n_25988;
wire n_25989;
wire n_25990;
wire n_25991;
wire n_25992;
wire n_25993;
wire n_25994;
wire n_25995;
wire n_25996;
wire n_25997;
wire n_25998;
wire n_25999;
wire n_26000;
wire n_26001;
wire n_26002;
wire n_26003;
wire n_26004;
wire n_26005;
wire n_26006;
wire n_26007;
wire n_26008;
wire n_26009;
wire n_26010;
wire n_26011;
wire n_26012;
wire n_26013;
wire n_26014;
wire n_26015;
wire n_26016;
wire n_26017;
wire n_26018;
wire n_26019;
wire n_26020;
wire n_26021;
wire n_26022;
wire n_26023;
wire n_26024;
wire n_26025;
wire n_26026;
wire n_26027;
wire n_26028;
wire n_26029;
wire n_26030;
wire n_26031;
wire n_26032;
wire n_26033;
wire n_26034;
wire n_26035;
wire n_26036;
wire n_26037;
wire n_26038;
wire n_26039;
wire n_26040;
wire n_26041;
wire n_26042;
wire n_26043;
wire n_26044;
wire n_26045;
wire n_26046;
wire n_26047;
wire n_26048;
wire n_26049;
wire n_26050;
wire n_26051;
wire n_26052;
wire n_26053;
wire n_26054;
wire n_26055;
wire n_26056;
wire n_26057;
wire n_26058;
wire n_26059;
wire n_26060;
wire n_26061;
wire n_26062;
wire n_26063;
wire n_26064;
wire n_26065;
wire n_26066;
wire n_26067;
wire n_26068;
wire n_26069;
wire n_26070;
wire n_26071;
wire n_26072;
wire n_26073;
wire n_26074;
wire n_26075;
wire n_26076;
wire n_26077;
wire n_26078;
wire n_26079;
wire n_26080;
wire n_26081;
wire n_26082;
wire n_26083;
wire n_26084;
wire n_26085;
wire n_26086;
wire n_26087;
wire n_26088;
wire n_26089;
wire n_26090;
wire n_26091;
wire n_26092;
wire n_26093;
wire n_26094;
wire n_26095;
wire n_26096;
wire n_26097;
wire n_26098;
wire n_26099;
wire n_26100;
wire n_26101;
wire n_26102;
wire n_26103;
wire n_26104;
wire n_26105;
wire n_26106;
wire n_26107;
wire n_26108;
wire n_26109;
wire n_26110;
wire n_26111;
wire n_26112;
wire n_26113;
wire n_26114;
wire n_26115;
wire n_26116;
wire n_26117;
wire n_26118;
wire n_26119;
wire n_26120;
wire n_26121;
wire n_26122;
wire n_26123;
wire n_26124;
wire n_26125;
wire n_26126;
wire n_26127;
wire n_26128;
wire n_26129;
wire n_26130;
wire n_26131;
wire n_26132;
wire n_26133;
wire n_26134;
wire n_26135;
wire n_26136;
wire n_26137;
wire n_26138;
wire n_26139;
wire n_26140;
wire n_26141;
wire n_26142;
wire n_26143;
wire n_26144;
wire n_26145;
wire n_26146;
wire n_26147;
wire n_26148;
wire n_26149;
wire n_26150;
wire n_26151;
wire n_26152;
wire n_26153;
wire n_26154;
wire n_26155;
wire n_26156;
wire n_26157;
wire n_26158;
wire n_26159;
wire n_26160;
wire n_26161;
wire n_26162;
wire n_26163;
wire n_26164;
wire n_26165;
wire n_26166;
wire n_26167;
wire n_26168;
wire n_26169;
wire n_26170;
wire n_26171;
wire n_26172;
wire n_26173;
wire n_26174;
wire n_26175;
wire n_26176;
wire n_26177;
wire n_26178;
wire n_26179;
wire n_26180;
wire n_26181;
wire n_26182;
wire n_26183;
wire n_26184;
wire n_26185;
wire n_26186;
wire n_26187;
wire n_26188;
wire n_26189;
wire n_26190;
wire n_26191;
wire n_26192;
wire n_26193;
wire n_26194;
wire n_26195;
wire n_26196;
wire n_26197;
wire n_26198;
wire n_26199;
wire n_26200;
wire n_26201;
wire n_26202;
wire n_26203;
wire n_26204;
wire n_26205;
wire n_26206;
wire n_26207;
wire n_26208;
wire n_26209;
wire n_26210;
wire n_26211;
wire n_26212;
wire n_26213;
wire n_26214;
wire n_26215;
wire n_26216;
wire n_26217;
wire n_26218;
wire n_26219;
wire n_26220;
wire n_26221;
wire n_26222;
wire n_26223;
wire n_26224;
wire n_26225;
wire n_26226;
wire n_26227;
wire n_26228;
wire n_26229;
wire n_26230;
wire n_26231;
wire n_26232;
wire n_26233;
wire n_26234;
wire n_26235;
wire n_26236;
wire n_26237;
wire n_26238;
wire n_26239;
wire n_26240;
wire n_26241;
wire n_26242;
wire n_26243;
wire n_26244;
wire n_26245;
wire n_26246;
wire n_26247;
wire n_26248;
wire n_26249;
wire n_26250;
wire n_26251;
wire n_26252;
wire n_26253;
wire n_26254;
wire n_26255;
wire n_26256;
wire n_26257;
wire n_26258;
wire n_26259;
wire n_26260;
wire n_26261;
wire n_26262;
wire n_26263;
wire n_26264;
wire n_26265;
wire n_26266;
wire n_26267;
wire n_26268;
wire n_26269;
wire n_26270;
wire n_26271;
wire n_26272;
wire n_26273;
wire n_26274;
wire n_26275;
wire n_26276;
wire n_26277;
wire n_26278;
wire n_26279;
wire n_26280;
wire n_26281;
wire n_26282;
wire n_26283;
wire n_26284;
wire n_26285;
wire n_26286;
wire n_26287;
wire n_26288;
wire n_26289;
wire n_26290;
wire n_26291;
wire n_26292;
wire n_26293;
wire n_26294;
wire n_26295;
wire n_26296;
wire n_26297;
wire n_26298;
wire n_26299;
wire n_26300;
wire n_26301;
wire n_26302;
wire n_26303;
wire n_26304;
wire n_26305;
wire n_26306;
wire n_26307;
wire n_26308;
wire n_26309;
wire n_26310;
wire n_26311;
wire n_26312;
wire n_26313;
wire n_26314;
wire n_26315;
wire n_26316;
wire n_26317;
wire n_26318;
wire n_26319;
wire n_26320;
wire n_26321;
wire n_26322;
wire n_26323;
wire n_26324;
wire n_26325;
wire n_26326;
wire n_26327;
wire n_26328;
wire n_26329;
wire n_26330;
wire n_26331;
wire n_26332;
wire n_26333;
wire n_26334;
wire n_26335;
wire n_26336;
wire n_26337;
wire n_26338;
wire n_26339;
wire n_26340;
wire n_26341;
wire n_26342;
wire n_26343;
wire n_26344;
wire n_26345;
wire n_26346;
wire n_26347;
wire n_26348;
wire n_26349;
wire n_26350;
wire n_26351;
wire n_26352;
wire n_26353;
wire n_26354;
wire n_26355;
wire n_26356;
wire n_26357;
wire n_26358;
wire n_26359;
wire n_26360;
wire n_26361;
wire n_26362;
wire n_26363;
wire n_26364;
wire n_26365;
wire n_26366;
wire n_26367;
wire n_26368;
wire n_26369;
wire n_26370;
wire n_26371;
wire n_26372;
wire n_26373;
wire n_26374;
wire n_26375;
wire n_26376;
wire n_26377;
wire n_26378;
wire n_26379;
wire n_26380;
wire n_26381;
wire n_26382;
wire n_26383;
wire n_26384;
wire n_26385;
wire n_26386;
wire n_26387;
wire n_26388;
wire n_26389;
wire n_26390;
wire n_26391;
wire n_26392;
wire n_26393;
wire n_26394;
wire n_26395;
wire n_26396;
wire n_26397;
wire n_26398;
wire n_26399;
wire n_26400;
wire n_26401;
wire n_26402;
wire n_26403;
wire n_26404;
wire n_26405;
wire n_26406;
wire n_26407;
wire n_26408;
wire n_26409;
wire n_26410;
wire n_26411;
wire n_26412;
wire n_26413;
wire n_26414;
wire n_26415;
wire n_26416;
wire n_26417;
wire n_26418;
wire n_26419;
wire n_26420;
wire n_26421;
wire n_26422;
wire n_26423;
wire n_26424;
wire n_26425;
wire n_26426;
wire n_26427;
wire n_26428;
wire n_26429;
wire n_26430;
wire n_26431;
wire n_26432;
wire n_26433;
wire n_26434;
wire n_26435;
wire n_26436;
wire n_26437;
wire n_26438;
wire n_26439;
wire n_26440;
wire n_26441;
wire n_26442;
wire n_26443;
wire n_26444;
wire n_26445;
wire n_26446;
wire n_26447;
wire n_26448;
wire n_26449;
wire n_26450;
wire n_26451;
wire n_26452;
wire n_26453;
wire n_26454;
wire n_26455;
wire n_26456;
wire n_26457;
wire n_26458;
wire n_26459;
wire n_26460;
wire n_26461;
wire n_26462;
wire n_26463;
wire n_26464;
wire n_26465;
wire n_26466;
wire n_26467;
wire n_26468;
wire n_26469;
wire n_26470;
wire n_26471;
wire n_26472;
wire n_26473;
wire n_26474;
wire n_26475;
wire n_26476;
wire n_26477;
wire n_26478;
wire n_26479;
wire n_26480;
wire n_26481;
wire n_26482;
wire n_26483;
wire n_26484;
wire n_26485;
wire n_26486;
wire n_26487;
wire n_26488;
wire n_26489;
wire n_26490;
wire n_26491;
wire n_26492;
wire n_26493;
wire n_26494;
wire n_26495;
wire n_26496;
wire n_26497;
wire n_26498;
wire n_26499;
wire n_26500;
wire n_26501;
wire n_26502;
wire n_26503;
wire n_26504;
wire n_26505;
wire n_26506;
wire n_26507;
wire n_26508;
wire n_26509;
wire n_26510;
wire n_26511;
wire n_26512;
wire n_26513;
wire n_26514;
wire n_26515;
wire n_26516;
wire n_26517;
wire n_26518;
wire n_26519;
wire n_26520;
wire n_26521;
wire n_26522;
wire n_26523;
wire n_26524;
wire n_26525;
wire n_26526;
wire n_26527;
wire n_26528;
wire n_26529;
wire n_26530;
wire n_26531;
wire n_26532;
wire n_26533;
wire n_26534;
wire n_26535;
wire n_26536;
wire n_26537;
wire n_26538;
wire n_26539;
wire n_26540;
wire n_26541;
wire n_26542;
wire n_26543;
wire n_26544;
wire n_26545;
wire n_26546;
wire n_26547;
wire n_26548;
wire n_26549;
wire n_26550;
wire n_26551;
wire n_26552;
wire n_26553;
wire n_26554;
wire n_26555;
wire n_26556;
wire n_26557;
wire n_26558;
wire n_26559;
wire n_26560;
wire n_26561;
wire n_26562;
wire n_26563;
wire n_26564;
wire n_26565;
wire n_26566;
wire n_26567;
wire n_26568;
wire n_26569;
wire n_26570;
wire n_26571;
wire n_26572;
wire n_26573;
wire n_26574;
wire n_26575;
wire n_26576;
wire n_26577;
wire n_26578;
wire n_26579;
wire n_26580;
wire n_26581;
wire n_26582;
wire n_26583;
wire n_26584;
wire n_26585;
wire n_26586;
wire n_26587;
wire n_26588;
wire n_26589;
wire n_26590;
wire n_26591;
wire n_26592;
wire n_26593;
wire n_26594;
wire n_26595;
wire n_26596;
wire n_26597;
wire n_26598;
wire n_26599;
wire n_26600;
wire n_26601;
wire n_26602;
wire n_26603;
wire n_26604;
wire n_26605;
wire n_26606;
wire n_26607;
wire n_26608;
wire n_26609;
wire n_26610;
wire n_26611;
wire n_26612;
wire n_26613;
wire n_26614;
wire n_26615;
wire n_26616;
wire n_26617;
wire n_26618;
wire n_26619;
wire n_26620;
wire n_26621;
wire n_26622;
wire n_26623;
wire n_26624;
wire n_26625;
wire n_26626;
wire n_26627;
wire n_26628;
wire n_26629;
wire n_26630;
wire n_26631;
wire n_26632;
wire n_26633;
wire n_26634;
wire n_26635;
wire n_26636;
wire n_26637;
wire n_26638;
wire n_26639;
wire n_26640;
wire n_26641;
wire n_26642;
wire n_26643;
wire n_26644;
wire n_26645;
wire n_26646;
wire n_26647;
wire n_26648;
wire n_26649;
wire n_26650;
wire n_26651;
wire n_26652;
wire n_26653;
wire n_26654;
wire n_26655;
wire n_26656;
wire n_26657;
wire n_26658;
wire n_26659;
wire n_26660;
wire n_26661;
wire n_26662;
wire n_26663;
wire n_26664;
wire n_26665;
wire n_26666;
wire n_26667;
wire n_26668;
wire n_26669;
wire n_26670;
wire n_26671;
wire n_26672;
wire n_26673;
wire n_26674;
wire n_26675;
wire n_26676;
wire n_26677;
wire n_26678;
wire n_26679;
wire n_26680;
wire n_26681;
wire n_26682;
wire n_26683;
wire n_26684;
wire n_26685;
wire n_26686;
wire n_26687;
wire n_26688;
wire n_26689;
wire n_26690;
wire n_26691;
wire n_26692;
wire n_26693;
wire n_26694;
wire n_26695;
wire n_26696;
wire n_26697;
wire n_26698;
wire n_26699;
wire n_26700;
wire n_26701;
wire n_26702;
wire n_26703;
wire n_26704;
wire n_26705;
wire n_26706;
wire n_26707;
wire n_26708;
wire n_26709;
wire n_26710;
wire n_26711;
wire n_26712;
wire n_26713;
wire n_26714;
wire n_26715;
wire n_26716;
wire n_26717;
wire n_26718;
wire n_26719;
wire n_26720;
wire n_26721;
wire n_26722;
wire n_26723;
wire n_26724;
wire n_26725;
wire n_26726;
wire n_26727;
wire n_26728;
wire n_26729;
wire n_26730;
wire n_26731;
wire n_26732;
wire n_26733;
wire n_26734;
wire n_26735;
wire n_26736;
wire n_26737;
wire n_26738;
wire n_26739;
wire n_26740;
wire n_26741;
wire n_26742;
wire n_26743;
wire n_26744;
wire n_26745;
wire n_26746;
wire n_26747;
wire n_26748;
wire n_26749;
wire n_26750;
wire n_26751;
wire n_26752;
wire n_26753;
wire n_26754;
wire n_26755;
wire n_26756;
wire n_26757;
wire n_26758;
wire n_26759;
wire n_26760;
wire n_26761;
wire n_26762;
wire n_26763;
wire n_26764;
wire n_26765;
wire n_26766;
wire n_26767;
wire n_26768;
wire n_26769;
wire n_26770;
wire n_26771;
wire n_26772;
wire n_26773;
wire n_26774;
wire n_26775;
wire n_26776;
wire n_26777;
wire n_26778;
wire n_26779;
wire n_26780;
wire n_26781;
wire n_26782;
wire n_26783;
wire n_26784;
wire n_26785;
wire n_26786;
wire n_26787;
wire n_26788;
wire n_26789;
wire n_26790;
wire n_26791;
wire n_26792;
wire n_26793;
wire n_26794;
wire n_26795;
wire n_26796;
wire n_26797;
wire n_26798;
wire n_26799;
wire n_26800;
wire n_26801;
wire n_26802;
wire n_26803;
wire n_26804;
wire n_26805;
wire n_26806;
wire n_26807;
wire n_26808;
wire n_26809;
wire n_26810;
wire n_26811;
wire n_26812;
wire n_26813;
wire n_26814;
wire n_26815;
wire n_26816;
wire n_26817;
wire n_26818;
wire n_26819;
wire n_26820;
wire n_26821;
wire n_26822;
wire n_26823;
wire n_26824;
wire n_26825;
wire n_26826;
wire n_26827;
wire n_26828;
wire n_26829;
wire n_26830;
wire n_26831;
wire n_26832;
wire n_26833;
wire n_26834;
wire n_26835;
wire n_26836;
wire n_26837;
wire n_26838;
wire n_26839;
wire n_26840;
wire n_26841;
wire n_26842;
wire n_26843;
wire n_26844;
wire n_26845;
wire n_26846;
wire n_26847;
wire n_26848;
wire n_26849;
wire n_26850;
wire n_26851;
wire n_26852;
wire n_26853;
wire n_26854;
wire n_26855;
wire n_26856;
wire n_26857;
wire n_26858;
wire n_26859;
wire n_26860;
wire n_26861;
wire n_26862;
wire n_26863;
wire n_26864;
wire n_26865;
wire n_26866;
wire n_26867;
wire n_26868;
wire n_26869;
wire n_26870;
wire n_26871;
wire n_26872;
wire n_26873;
wire n_26874;
wire n_26875;
wire n_26876;
wire n_26877;
wire n_26878;
wire n_26879;
wire n_26880;
wire n_26881;
wire n_26882;
wire n_26883;
wire n_26884;
wire n_26885;
wire n_26886;
wire n_26887;
wire n_26888;
wire n_26889;
wire n_26890;
wire n_26891;
wire n_26892;
wire n_26893;
wire n_26894;
wire n_26895;
wire n_26896;
wire n_26897;
wire n_26898;
wire n_26899;
wire n_26900;
wire n_26901;
wire n_26902;
wire n_26903;
wire n_26904;
wire n_26905;
wire n_26906;
wire n_26907;
wire n_26908;
wire n_26909;
wire n_26910;
wire n_26911;
wire n_26912;
wire n_26913;
wire n_26914;
wire n_26915;
wire n_26916;
wire n_26917;
wire n_26918;
wire n_26919;
wire n_26920;
wire n_26921;
wire n_26922;
wire n_26923;
wire n_26924;
wire n_26925;
wire n_26926;
wire n_26927;
wire n_26928;
wire n_26929;
wire n_26930;
wire n_26931;
wire n_26932;
wire n_26933;
wire n_26934;
wire n_26935;
wire n_26936;
wire n_26937;
wire n_26938;
wire n_26939;
wire n_26940;
wire n_26941;
wire n_26942;
wire n_26943;
wire n_26944;
wire n_26945;
wire n_26946;
wire n_26947;
wire n_26948;
wire n_26949;
wire n_26950;
wire n_26951;
wire n_26952;
wire n_26953;
wire n_26954;
wire n_26955;
wire n_26956;
wire n_26957;
wire n_26958;
wire n_26959;
wire n_26960;
wire n_26961;
wire n_26962;
wire n_26963;
wire n_26964;
wire n_26965;
wire n_26966;
wire n_26967;
wire n_26968;
wire n_26969;
wire n_26970;
wire n_26971;
wire n_26972;
wire n_26973;
wire n_26974;
wire n_26975;
wire n_26976;
wire n_26977;
wire n_26978;
wire n_26979;
wire n_26980;
wire n_26981;
wire n_26982;
wire n_26983;
wire n_26984;
wire n_26985;
wire n_26986;
wire n_26987;
wire n_26988;
wire n_26989;
wire n_26990;
wire n_26991;
wire n_26992;
wire n_26993;
wire n_26994;
wire n_26995;
wire n_26996;
wire n_26997;
wire n_26998;
wire n_26999;
wire n_27000;
wire n_27001;
wire n_27002;
wire n_27003;
wire n_27004;
wire n_27005;
wire n_27006;
wire n_27007;
wire n_27008;
wire n_27009;
wire n_27010;
wire n_27011;
wire n_27012;
wire n_27013;
wire n_27014;
wire n_27015;
wire n_27016;
wire n_27017;
wire n_27018;
wire n_27019;
wire n_27020;
wire n_27021;
wire n_27022;
wire n_27023;
wire n_27024;
wire n_27025;
wire n_27026;
wire n_27027;
wire n_27028;
wire n_27029;
wire n_27030;
wire n_27031;
wire n_27032;
wire n_27033;
wire n_27034;
wire n_27035;
wire n_27036;
wire n_27037;
wire n_27038;
wire n_27039;
wire n_27040;
wire n_27041;
wire n_27042;
wire n_27043;
wire n_27044;
wire n_27045;
wire n_27046;
wire n_27047;
wire n_27048;
wire n_27049;
wire n_27050;
wire n_27051;
wire n_27052;
wire n_27053;
wire n_27054;
wire n_27055;
wire n_27056;
wire n_27057;
wire n_27058;
wire n_27059;
wire n_27060;
wire n_27061;
wire n_27062;
wire n_27063;
wire n_27064;
wire n_27065;
wire n_27066;
wire n_27067;
wire n_27068;
wire n_27069;
wire n_27070;
wire n_27071;
wire n_27072;
wire n_27073;
wire n_27074;
wire n_27075;
wire n_27076;
wire n_27077;
wire n_27078;
wire n_27079;
wire n_27080;
wire n_27081;
wire n_27082;
wire n_27083;
wire n_27084;
wire n_27085;
wire n_27086;
wire n_27087;
wire n_27088;
wire n_27089;
wire n_27090;
wire n_27091;
wire n_27092;
wire n_27093;
wire n_27094;
wire n_27095;
wire n_27096;
wire n_27097;
wire n_27098;
wire n_27099;
wire n_27100;
wire n_27101;
wire n_27102;
wire n_27103;
wire n_27104;
wire n_27105;
wire n_27106;
wire n_27107;
wire n_27108;
wire n_27109;
wire n_27110;
wire n_27111;
wire n_27112;
wire n_27113;
wire n_27114;
wire n_27115;
wire n_27116;
wire n_27117;
wire n_27118;
wire n_27119;
wire n_27120;
wire n_27121;
wire n_27122;
wire n_27123;
wire n_27124;
wire n_27125;
wire n_27126;
wire n_27127;
wire n_27128;
wire n_27129;
wire n_27130;
wire n_27131;
wire n_27132;
wire n_27133;
wire n_27134;
wire n_27135;
wire n_27136;
wire n_27137;
wire n_27138;
wire n_27139;
wire n_27140;
wire n_27141;
wire n_27142;
wire n_27143;
wire n_27144;
wire n_27145;
wire n_27146;
wire n_27147;
wire n_27148;
wire n_27149;
wire n_27150;
wire n_27151;
wire n_27152;
wire n_27153;
wire n_27154;
wire n_27155;
wire n_27156;
wire n_27157;
wire n_27158;
wire n_27159;
wire n_27160;
wire n_27161;
wire n_27162;
wire n_27163;
wire n_27164;
wire n_27165;
wire n_27166;
wire n_27167;
wire n_27168;
wire n_27169;
wire n_27170;
wire n_27171;
wire n_27172;
wire n_27173;
wire n_27174;
wire n_27175;
wire n_27176;
wire n_27177;
wire n_27178;
wire n_27179;
wire n_27180;
wire n_27181;
wire n_27182;
wire n_27183;
wire n_27184;
wire n_27185;
wire n_27186;
wire n_27187;
wire n_27188;
wire n_27189;
wire n_27190;
wire n_27191;
wire n_27192;
wire n_27193;
wire n_27194;
wire n_27195;
wire n_27196;
wire n_27197;
wire n_27198;
wire n_27199;
wire n_27200;
wire n_27201;
wire n_27202;
wire n_27203;
wire n_27204;
wire n_27205;
wire n_27206;
wire n_27207;
wire n_27208;
wire n_27209;
wire n_27210;
wire n_27211;
wire n_27212;
wire n_27213;
wire n_27214;
wire n_27215;
wire n_27216;
wire n_27217;
wire n_27218;
wire n_27219;
wire n_27220;
wire n_27221;
wire n_27222;
wire n_27223;
wire n_27224;
wire n_27225;
wire n_27226;
wire n_27227;
wire n_27228;
wire n_27229;
wire n_27230;
wire n_27231;
wire n_27232;
wire n_27233;
wire n_27234;
wire n_27235;
wire n_27236;
wire n_27237;
wire n_27238;
wire n_27239;
wire n_27240;
wire n_27241;
wire n_27242;
wire n_27243;
wire n_27244;
wire n_27245;
wire n_27246;
wire n_27247;
wire n_27248;
wire n_27249;
wire n_27250;
wire n_27251;
wire n_27252;
wire n_27253;
wire n_27254;
wire n_27255;
wire n_27256;
wire n_27257;
wire n_27258;
wire n_27259;
wire n_27260;
wire n_27261;
wire n_27262;
wire n_27263;
wire n_27264;
wire n_27265;
wire n_27266;
wire n_27267;
wire n_27268;
wire n_27269;
wire n_27270;
wire n_27271;
wire n_27272;
wire n_27273;
wire n_27274;
wire n_27275;
wire n_27276;
wire n_27277;
wire n_27278;
wire n_27279;
wire n_27280;
wire n_27281;
wire n_27282;
wire n_27283;
wire n_27284;
wire n_27285;
wire n_27286;
wire n_27287;
wire n_27288;
wire n_27289;
wire n_27290;
wire n_27291;
wire n_27292;
wire n_27293;
wire n_27294;
wire n_27295;
wire n_27296;
wire n_27297;
wire n_27298;
wire n_27299;
wire n_27300;
wire n_27301;
wire n_27302;
wire n_27303;
wire n_27304;
wire n_27305;
wire n_27306;
wire n_27307;
wire n_27308;
wire n_27309;
wire n_27310;
wire n_27311;
wire n_27312;
wire n_27313;
wire n_27314;
wire n_27315;
wire n_27316;
wire n_27317;
wire n_27318;
wire n_27319;
wire n_27320;
wire n_27321;
wire n_27322;
wire n_27323;
wire n_27324;
wire n_27325;
wire n_27326;
wire n_27327;
wire n_27328;
wire n_27329;
wire n_27330;
wire n_27331;
wire n_27332;
wire n_27333;
wire n_27334;
wire n_27335;
wire n_27336;
wire n_27337;
wire n_27338;
wire n_27339;
wire n_27340;
wire n_27341;
wire n_27342;
wire n_27343;
wire n_27344;
wire n_27345;
wire n_27346;
wire n_27347;
wire n_27348;
wire n_27349;
wire n_27350;
wire n_27351;
wire n_27352;
wire n_27353;
wire n_27354;
wire n_27355;
wire n_27356;
wire n_27357;
wire n_27358;
wire n_27359;
wire n_27360;
wire n_27361;
wire n_27362;
wire n_27363;
wire n_27364;
wire n_27365;
wire n_27366;
wire n_27367;
wire n_27368;
wire n_27369;
wire n_27370;
wire n_27371;
wire n_27372;
wire n_27373;
wire n_27374;
wire n_27375;
wire n_27376;
wire n_27377;
wire n_27378;
wire n_27379;
wire n_27380;
wire n_27381;
wire n_27382;
wire n_27383;
wire n_27384;
wire n_27385;
wire n_27386;
wire n_27387;
wire n_27388;
wire n_27389;
wire n_27390;
wire n_27391;
wire n_27392;
wire n_27393;
wire n_27394;
wire n_27395;
wire n_27396;
wire n_27397;
wire n_27398;
wire n_27399;
wire n_27400;
wire n_27401;
wire n_27402;
wire n_27403;
wire n_27404;
wire n_27405;
wire n_27406;
wire n_27407;
wire n_27408;
wire n_27409;
wire n_27410;
wire n_27411;
wire n_27412;
wire n_27413;
wire n_27414;
wire n_27415;
wire n_27416;
wire n_27417;
wire n_27418;
wire n_27419;
wire n_27420;
wire n_27421;
wire n_27422;
wire n_27423;
wire n_27424;
wire n_27425;
wire n_27426;
wire n_27427;
wire n_27428;
wire n_27429;
assign n_1 =  x_398 &  x_1596;
assign n_2 = ~x_398 & ~x_1596;
assign n_3 = ~n_1 & ~n_2;
assign n_4 = ~x_399 &  n_3;
assign n_5 =  x_400 &  n_4;
assign n_6 = ~x_1380 &  n_5;
assign n_7 =  x_399 &  n_3;
assign n_8 =  x_400 &  n_7;
assign n_9 = ~x_1378 &  n_8;
assign n_10 = ~n_6 & ~n_9;
assign n_11 = ~x_400 &  n_7;
assign n_12 = ~x_1382 &  n_11;
assign n_13 = ~x_400 &  n_4;
assign n_14 = ~x_1384 &  n_13;
assign n_15 = ~n_12 & ~n_14;
assign n_16 =  n_10 &  n_15;
assign n_17 =  x_399 &  n_1;
assign n_18 =  x_400 & ~n_17;
assign n_19 = ~x_400 &  n_17;
assign n_20 = ~n_18 & ~n_19;
assign n_21 = ~x_399 & ~n_1;
assign n_22 = ~n_17 & ~n_21;
assign n_23 = ~n_3 & ~n_22;
assign n_24 = ~n_20 &  n_23;
assign n_25 = ~x_1381 &  n_24;
assign n_26 =  n_20 &  n_23;
assign n_27 = ~x_1385 &  n_26;
assign n_28 = ~n_25 & ~n_27;
assign n_29 = ~n_3 &  n_22;
assign n_30 =  x_400 &  n_29;
assign n_31 = ~x_1379 &  n_30;
assign n_32 = ~x_400 &  n_29;
assign n_33 = ~x_1383 &  n_32;
assign n_34 = ~n_31 & ~n_33;
assign n_35 =  n_28 &  n_34;
assign n_36 =  n_16 &  n_35;
assign n_37 =  x_424 &  n_36;
assign n_38 = ~x_424 & ~n_36;
assign n_39 = ~n_37 & ~n_38;
assign n_40 = ~x_1376 &  n_13;
assign n_41 = ~x_1374 &  n_11;
assign n_42 = ~n_40 & ~n_41;
assign n_43 = ~x_1370 &  n_8;
assign n_44 = ~x_1372 &  n_5;
assign n_45 = ~n_43 & ~n_44;
assign n_46 =  n_42 &  n_45;
assign n_47 = ~x_1377 &  n_26;
assign n_48 = ~x_1371 &  n_30;
assign n_49 = ~n_47 & ~n_48;
assign n_50 = ~x_1373 &  n_24;
assign n_51 = ~x_1375 &  n_32;
assign n_52 = ~n_50 & ~n_51;
assign n_53 =  n_49 &  n_52;
assign n_54 =  n_46 &  n_53;
assign n_55 =  x_423 &  n_54;
assign n_56 = ~x_423 & ~n_54;
assign n_57 = ~n_55 & ~n_56;
assign n_58 = ~x_1368 &  n_13;
assign n_59 = ~x_1362 &  n_8;
assign n_60 = ~n_58 & ~n_59;
assign n_61 = ~x_1366 &  n_11;
assign n_62 = ~x_1364 &  n_5;
assign n_63 = ~n_61 & ~n_62;
assign n_64 =  n_60 &  n_63;
assign n_65 = ~x_1365 &  n_24;
assign n_66 = ~x_1369 &  n_26;
assign n_67 = ~n_65 & ~n_66;
assign n_68 = ~x_1363 &  n_30;
assign n_69 = ~x_1367 &  n_32;
assign n_70 = ~n_68 & ~n_69;
assign n_71 =  n_67 &  n_70;
assign n_72 =  n_64 &  n_71;
assign n_73 =  x_422 &  n_72;
assign n_74 = ~x_422 & ~n_72;
assign n_75 = ~n_73 & ~n_74;
assign n_76 = ~x_1354 &  n_8;
assign n_77 = ~x_1356 &  n_5;
assign n_78 = ~n_76 & ~n_77;
assign n_79 = ~x_1358 &  n_11;
assign n_80 = ~x_1360 &  n_13;
assign n_81 = ~n_79 & ~n_80;
assign n_82 =  n_78 &  n_81;
assign n_83 = ~x_1361 &  n_26;
assign n_84 = ~x_1359 &  n_32;
assign n_85 = ~n_83 & ~n_84;
assign n_86 = ~x_1357 &  n_24;
assign n_87 = ~x_1355 &  n_30;
assign n_88 = ~n_86 & ~n_87;
assign n_89 =  n_85 &  n_88;
assign n_90 =  n_82 &  n_89;
assign n_91 =  x_421 &  n_90;
assign n_92 = ~x_421 & ~n_90;
assign n_93 = ~n_91 & ~n_92;
assign n_94 = ~x_1350 &  n_11;
assign n_95 = ~x_1348 &  n_5;
assign n_96 = ~n_94 & ~n_95;
assign n_97 = ~x_1346 &  n_8;
assign n_98 = ~x_1352 &  n_13;
assign n_99 = ~n_97 & ~n_98;
assign n_100 =  n_96 &  n_99;
assign n_101 = ~x_1347 &  n_30;
assign n_102 = ~x_1353 &  n_26;
assign n_103 = ~n_101 & ~n_102;
assign n_104 = ~x_1351 &  n_32;
assign n_105 = ~x_1349 &  n_24;
assign n_106 = ~n_104 & ~n_105;
assign n_107 =  n_103 &  n_106;
assign n_108 =  n_100 &  n_107;
assign n_109 =  x_420 &  n_108;
assign n_110 = ~x_420 & ~n_108;
assign n_111 = ~n_109 & ~n_110;
assign n_112 = ~x_1340 &  n_5;
assign n_113 = ~x_1338 &  n_8;
assign n_114 = ~n_112 & ~n_113;
assign n_115 = ~x_1342 &  n_11;
assign n_116 = ~x_1344 &  n_13;
assign n_117 = ~n_115 & ~n_116;
assign n_118 =  n_114 &  n_117;
assign n_119 = ~x_1341 &  n_24;
assign n_120 = ~x_1345 &  n_26;
assign n_121 = ~n_119 & ~n_120;
assign n_122 = ~x_1339 &  n_30;
assign n_123 = ~x_1343 &  n_32;
assign n_124 = ~n_122 & ~n_123;
assign n_125 =  n_121 &  n_124;
assign n_126 =  n_118 &  n_125;
assign n_127 =  x_419 &  n_126;
assign n_128 = ~x_419 & ~n_126;
assign n_129 = ~n_127 & ~n_128;
assign n_130 = ~x_1332 &  n_5;
assign n_131 = ~x_1334 &  n_11;
assign n_132 = ~n_130 & ~n_131;
assign n_133 = ~x_1330 &  n_8;
assign n_134 = ~x_1336 &  n_13;
assign n_135 = ~n_133 & ~n_134;
assign n_136 =  n_132 &  n_135;
assign n_137 = ~x_1335 &  n_32;
assign n_138 = ~x_1333 &  n_24;
assign n_139 = ~n_137 & ~n_138;
assign n_140 = ~x_1337 &  n_26;
assign n_141 = ~x_1331 &  n_30;
assign n_142 = ~n_140 & ~n_141;
assign n_143 =  n_139 &  n_142;
assign n_144 =  n_136 &  n_143;
assign n_145 =  x_418 &  n_144;
assign n_146 = ~x_418 & ~n_144;
assign n_147 = ~n_145 & ~n_146;
assign n_148 = ~x_1324 &  n_5;
assign n_149 = ~x_1326 &  n_11;
assign n_150 = ~n_148 & ~n_149;
assign n_151 = ~x_1328 &  n_13;
assign n_152 = ~x_1322 &  n_8;
assign n_153 = ~n_151 & ~n_152;
assign n_154 =  n_150 &  n_153;
assign n_155 = ~x_1323 &  n_30;
assign n_156 = ~x_1327 &  n_32;
assign n_157 = ~n_155 & ~n_156;
assign n_158 = ~x_1329 &  n_26;
assign n_159 = ~x_1325 &  n_24;
assign n_160 = ~n_158 & ~n_159;
assign n_161 =  n_157 &  n_160;
assign n_162 =  n_154 &  n_161;
assign n_163 =  x_417 &  n_162;
assign n_164 = ~x_417 & ~n_162;
assign n_165 = ~n_163 & ~n_164;
assign n_166 = ~x_1316 &  n_5;
assign n_167 = ~x_1314 &  n_8;
assign n_168 = ~n_166 & ~n_167;
assign n_169 = ~x_1320 &  n_13;
assign n_170 = ~x_1318 &  n_11;
assign n_171 = ~n_169 & ~n_170;
assign n_172 =  n_168 &  n_171;
assign n_173 = ~x_1317 &  n_24;
assign n_174 = ~x_1315 &  n_30;
assign n_175 = ~n_173 & ~n_174;
assign n_176 = ~x_1319 &  n_32;
assign n_177 = ~x_1321 &  n_26;
assign n_178 = ~n_176 & ~n_177;
assign n_179 =  n_175 &  n_178;
assign n_180 =  n_172 &  n_179;
assign n_181 =  x_416 &  n_180;
assign n_182 = ~x_416 & ~n_180;
assign n_183 = ~n_181 & ~n_182;
assign n_184 = ~x_1308 &  n_5;
assign n_185 = ~x_1306 &  n_8;
assign n_186 = ~n_184 & ~n_185;
assign n_187 = ~x_1312 &  n_13;
assign n_188 = ~x_1310 &  n_11;
assign n_189 = ~n_187 & ~n_188;
assign n_190 =  n_186 &  n_189;
assign n_191 = ~x_1309 &  n_24;
assign n_192 = ~x_1307 &  n_30;
assign n_193 = ~n_191 & ~n_192;
assign n_194 = ~x_1311 &  n_32;
assign n_195 = ~x_1313 &  n_26;
assign n_196 = ~n_194 & ~n_195;
assign n_197 =  n_193 &  n_196;
assign n_198 =  n_190 &  n_197;
assign n_199 =  x_415 &  n_198;
assign n_200 = ~x_415 & ~n_198;
assign n_201 = ~n_199 & ~n_200;
assign n_202 = ~x_1298 &  n_8;
assign n_203 = ~x_1302 &  n_11;
assign n_204 = ~n_202 & ~n_203;
assign n_205 = ~x_1304 &  n_13;
assign n_206 = ~x_1300 &  n_5;
assign n_207 = ~n_205 & ~n_206;
assign n_208 =  n_204 &  n_207;
assign n_209 = ~x_1299 &  n_30;
assign n_210 = ~x_1305 &  n_26;
assign n_211 = ~n_209 & ~n_210;
assign n_212 = ~x_1301 &  n_24;
assign n_213 = ~x_1303 &  n_32;
assign n_214 = ~n_212 & ~n_213;
assign n_215 =  n_211 &  n_214;
assign n_216 =  n_208 &  n_215;
assign n_217 =  x_414 &  n_216;
assign n_218 = ~x_414 & ~n_216;
assign n_219 = ~n_217 & ~n_218;
assign n_220 = ~x_1294 &  n_11;
assign n_221 = ~x_1292 &  n_5;
assign n_222 = ~n_220 & ~n_221;
assign n_223 = ~x_1290 &  n_8;
assign n_224 = ~x_1296 &  n_13;
assign n_225 = ~n_223 & ~n_224;
assign n_226 =  n_222 &  n_225;
assign n_227 = ~x_1297 &  n_26;
assign n_228 = ~x_1291 &  n_30;
assign n_229 = ~n_227 & ~n_228;
assign n_230 = ~x_1295 &  n_32;
assign n_231 = ~x_1293 &  n_24;
assign n_232 = ~n_230 & ~n_231;
assign n_233 =  n_229 &  n_232;
assign n_234 =  n_226 &  n_233;
assign n_235 =  x_413 &  n_234;
assign n_236 = ~x_413 & ~n_234;
assign n_237 = ~n_235 & ~n_236;
assign n_238 = ~x_1286 &  n_11;
assign n_239 = ~x_1284 &  n_5;
assign n_240 = ~n_238 & ~n_239;
assign n_241 = ~x_1282 &  n_8;
assign n_242 = ~x_1288 &  n_13;
assign n_243 = ~n_241 & ~n_242;
assign n_244 =  n_240 &  n_243;
assign n_245 = ~x_1287 &  n_32;
assign n_246 = ~x_1283 &  n_30;
assign n_247 = ~n_245 & ~n_246;
assign n_248 = ~x_1285 &  n_24;
assign n_249 = ~x_1289 &  n_26;
assign n_250 = ~n_248 & ~n_249;
assign n_251 =  n_247 &  n_250;
assign n_252 =  n_244 &  n_251;
assign n_253 =  x_412 &  n_252;
assign n_254 = ~x_412 & ~n_252;
assign n_255 = ~n_253 & ~n_254;
assign n_256 = ~x_1280 &  n_13;
assign n_257 = ~x_1276 &  n_5;
assign n_258 = ~n_256 & ~n_257;
assign n_259 = ~x_1278 &  n_11;
assign n_260 = ~x_1274 &  n_8;
assign n_261 = ~n_259 & ~n_260;
assign n_262 =  n_258 &  n_261;
assign n_263 = ~x_1281 &  n_26;
assign n_264 = ~x_1275 &  n_30;
assign n_265 = ~n_263 & ~n_264;
assign n_266 = ~x_1279 &  n_32;
assign n_267 = ~x_1277 &  n_24;
assign n_268 = ~n_266 & ~n_267;
assign n_269 =  n_265 &  n_268;
assign n_270 =  n_262 &  n_269;
assign n_271 =  x_411 &  n_270;
assign n_272 = ~x_411 & ~n_270;
assign n_273 = ~n_271 & ~n_272;
assign n_274 = ~x_1272 &  n_13;
assign n_275 = ~x_1268 &  n_5;
assign n_276 = ~n_274 & ~n_275;
assign n_277 = ~x_1270 &  n_11;
assign n_278 = ~x_1266 &  n_8;
assign n_279 = ~n_277 & ~n_278;
assign n_280 =  n_276 &  n_279;
assign n_281 = ~x_1271 &  n_32;
assign n_282 = ~x_1273 &  n_26;
assign n_283 = ~n_281 & ~n_282;
assign n_284 = ~x_1269 &  n_24;
assign n_285 = ~x_1267 &  n_30;
assign n_286 = ~n_284 & ~n_285;
assign n_287 =  n_283 &  n_286;
assign n_288 =  n_280 &  n_287;
assign n_289 =  x_410 &  n_288;
assign n_290 = ~x_410 & ~n_288;
assign n_291 = ~n_289 & ~n_290;
assign n_292 = ~x_1260 &  n_5;
assign n_293 = ~x_1262 &  n_11;
assign n_294 = ~n_292 & ~n_293;
assign n_295 = ~x_1264 &  n_13;
assign n_296 = ~x_1258 &  n_8;
assign n_297 = ~n_295 & ~n_296;
assign n_298 =  n_294 &  n_297;
assign n_299 = ~x_1265 &  n_26;
assign n_300 = ~x_1261 &  n_24;
assign n_301 = ~n_299 & ~n_300;
assign n_302 = ~x_1259 &  n_30;
assign n_303 = ~x_1263 &  n_32;
assign n_304 = ~n_302 & ~n_303;
assign n_305 =  n_301 &  n_304;
assign n_306 =  n_298 &  n_305;
assign n_307 =  x_409 &  n_306;
assign n_308 = ~x_409 & ~n_306;
assign n_309 = ~n_307 & ~n_308;
assign n_310 = ~x_1250 &  n_8;
assign n_311 = ~x_1256 &  n_13;
assign n_312 = ~n_310 & ~n_311;
assign n_313 = ~x_1254 &  n_11;
assign n_314 = ~x_1252 &  n_5;
assign n_315 = ~n_313 & ~n_314;
assign n_316 =  n_312 &  n_315;
assign n_317 = ~x_1257 &  n_26;
assign n_318 = ~x_1253 &  n_24;
assign n_319 = ~n_317 & ~n_318;
assign n_320 = ~x_1255 &  n_32;
assign n_321 = ~x_1251 &  n_30;
assign n_322 = ~n_320 & ~n_321;
assign n_323 =  n_319 &  n_322;
assign n_324 =  n_316 &  n_323;
assign n_325 =  x_408 &  n_324;
assign n_326 = ~x_408 & ~n_324;
assign n_327 = ~n_325 & ~n_326;
assign n_328 = ~x_1244 &  n_5;
assign n_329 = ~x_1248 &  n_13;
assign n_330 = ~n_328 & ~n_329;
assign n_331 = ~x_1242 &  n_8;
assign n_332 = ~x_1246 &  n_11;
assign n_333 = ~n_331 & ~n_332;
assign n_334 =  n_330 &  n_333;
assign n_335 = ~x_1249 &  n_26;
assign n_336 = ~x_1245 &  n_24;
assign n_337 = ~n_335 & ~n_336;
assign n_338 = ~x_1243 &  n_30;
assign n_339 = ~x_1247 &  n_32;
assign n_340 = ~n_338 & ~n_339;
assign n_341 =  n_337 &  n_340;
assign n_342 =  n_334 &  n_341;
assign n_343 =  x_407 &  n_342;
assign n_344 = ~x_407 & ~n_342;
assign n_345 = ~n_343 & ~n_344;
assign n_346 = ~x_1234 &  n_8;
assign n_347 = ~x_1238 &  n_11;
assign n_348 = ~n_346 & ~n_347;
assign n_349 = ~x_1240 &  n_13;
assign n_350 = ~x_1236 &  n_5;
assign n_351 = ~n_349 & ~n_350;
assign n_352 =  n_348 &  n_351;
assign n_353 = ~x_1239 &  n_32;
assign n_354 = ~x_1235 &  n_30;
assign n_355 = ~n_353 & ~n_354;
assign n_356 = ~x_1237 &  n_24;
assign n_357 = ~x_1241 &  n_26;
assign n_358 = ~n_356 & ~n_357;
assign n_359 =  n_355 &  n_358;
assign n_360 =  n_352 &  n_359;
assign n_361 =  x_406 &  n_360;
assign n_362 = ~x_406 & ~n_360;
assign n_363 = ~n_361 & ~n_362;
assign n_364 = ~x_1228 &  n_5;
assign n_365 = ~x_1232 &  n_13;
assign n_366 = ~n_364 & ~n_365;
assign n_367 = ~x_1230 &  n_11;
assign n_368 = ~x_1226 &  n_8;
assign n_369 = ~n_367 & ~n_368;
assign n_370 =  n_366 &  n_369;
assign n_371 = ~x_1233 &  n_26;
assign n_372 = ~x_1227 &  n_30;
assign n_373 = ~n_371 & ~n_372;
assign n_374 = ~x_1231 &  n_32;
assign n_375 = ~x_1229 &  n_24;
assign n_376 = ~n_374 & ~n_375;
assign n_377 =  n_373 &  n_376;
assign n_378 =  n_370 &  n_377;
assign n_379 =  x_405 &  n_378;
assign n_380 = ~x_405 & ~n_378;
assign n_381 = ~n_379 & ~n_380;
assign n_382 = ~x_1220 &  n_5;
assign n_383 = ~x_1222 &  n_11;
assign n_384 = ~n_382 & ~n_383;
assign n_385 = ~x_1218 &  n_8;
assign n_386 = ~x_1224 &  n_13;
assign n_387 = ~n_385 & ~n_386;
assign n_388 =  n_384 &  n_387;
assign n_389 = ~x_1219 &  n_30;
assign n_390 = ~x_1225 &  n_26;
assign n_391 = ~n_389 & ~n_390;
assign n_392 = ~x_1223 &  n_32;
assign n_393 = ~x_1221 &  n_24;
assign n_394 = ~n_392 & ~n_393;
assign n_395 =  n_391 &  n_394;
assign n_396 =  n_388 &  n_395;
assign n_397 =  x_404 &  n_396;
assign n_398 = ~x_404 & ~n_396;
assign n_399 = ~n_397 & ~n_398;
assign n_400 = ~x_1216 &  n_13;
assign n_401 = ~x_1212 &  n_5;
assign n_402 = ~n_400 & ~n_401;
assign n_403 = ~x_1210 &  n_8;
assign n_404 = ~x_1214 &  n_11;
assign n_405 = ~n_403 & ~n_404;
assign n_406 =  n_402 &  n_405;
assign n_407 = ~x_1213 &  n_24;
assign n_408 = ~x_1211 &  n_30;
assign n_409 = ~n_407 & ~n_408;
assign n_410 = ~x_1217 &  n_26;
assign n_411 = ~x_1215 &  n_32;
assign n_412 = ~n_410 & ~n_411;
assign n_413 =  n_409 &  n_412;
assign n_414 =  n_406 &  n_413;
assign n_415 =  x_403 &  n_414;
assign n_416 = ~x_403 & ~n_414;
assign n_417 = ~n_415 & ~n_416;
assign n_418 = ~x_1208 &  n_13;
assign n_419 = ~x_1206 &  n_11;
assign n_420 = ~n_418 & ~n_419;
assign n_421 = ~x_1204 &  n_5;
assign n_422 = ~x_1202 &  n_8;
assign n_423 = ~n_421 & ~n_422;
assign n_424 =  n_420 &  n_423;
assign n_425 = ~x_1207 &  n_32;
assign n_426 = ~x_1209 &  n_26;
assign n_427 = ~n_425 & ~n_426;
assign n_428 = ~x_1203 &  n_30;
assign n_429 = ~x_1205 &  n_24;
assign n_430 = ~n_428 & ~n_429;
assign n_431 =  n_427 &  n_430;
assign n_432 =  n_424 &  n_431;
assign n_433 =  x_402 &  n_432;
assign n_434 = ~x_402 & ~n_432;
assign n_435 = ~n_433 & ~n_434;
assign n_436 =  x_320 &  x_1472;
assign n_437 =  x_297 &  x_301;
assign n_438 = ~x_297 & ~x_301;
assign n_439 = ~n_437 & ~n_438;
assign n_440 = ~x_298 &  n_439;
assign n_441 = ~x_299 &  n_440;
assign n_442 = ~x_1606 &  n_441;
assign n_443 =  x_298 &  n_439;
assign n_444 = ~x_299 &  n_443;
assign n_445 = ~x_1609 &  n_444;
assign n_446 = ~n_442 & ~n_445;
assign n_447 =  x_299 &  n_443;
assign n_448 = ~x_1604 &  n_447;
assign n_449 =  x_299 &  n_440;
assign n_450 = ~x_1605 &  n_449;
assign n_451 = ~n_448 & ~n_450;
assign n_452 =  n_446 &  n_451;
assign n_453 =  x_298 &  n_437;
assign n_454 = ~x_298 & ~n_437;
assign n_455 = ~n_453 & ~n_454;
assign n_456 = ~n_439 & ~n_455;
assign n_457 = ~x_299 & ~n_453;
assign n_458 =  x_299 &  n_453;
assign n_459 = ~n_457 & ~n_458;
assign n_460 =  n_456 & ~n_459;
assign n_461 = ~x_1608 &  n_460;
assign n_462 = ~n_439 &  n_455;
assign n_463 =  x_299 &  n_462;
assign n_464 = ~x_1603 &  n_463;
assign n_465 = ~n_461 & ~n_464;
assign n_466 =  n_456 &  n_459;
assign n_467 = ~x_1607 &  n_466;
assign n_468 = ~x_299 &  n_462;
assign n_469 = ~x_1602 &  n_468;
assign n_470 = ~n_467 & ~n_469;
assign n_471 =  n_465 &  n_470;
assign n_472 =  n_452 &  n_471;
assign n_473 =  n_436 & ~n_472;
assign n_474 =  x_305 & ~n_436;
assign n_475 = ~n_473 & ~n_474;
assign n_476 =  x_306 & ~n_436;
assign n_477 = ~x_1615 &  n_449;
assign n_478 = ~x_1617 &  n_444;
assign n_479 = ~n_477 & ~n_478;
assign n_480 = ~x_1612 &  n_447;
assign n_481 = ~x_1613 &  n_441;
assign n_482 = ~n_480 & ~n_481;
assign n_483 =  n_479 &  n_482;
assign n_484 = ~x_1616 &  n_468;
assign n_485 = ~x_1611 &  n_463;
assign n_486 = ~n_484 & ~n_485;
assign n_487 = ~x_1614 &  n_466;
assign n_488 = ~x_1610 &  n_460;
assign n_489 = ~n_487 & ~n_488;
assign n_490 =  n_486 &  n_489;
assign n_491 =  n_483 &  n_490;
assign n_492 =  n_436 & ~n_491;
assign n_493 = ~x_1479 &  n_449;
assign n_494 = ~x_1475 &  n_447;
assign n_495 = ~n_493 & ~n_494;
assign n_496 = ~x_1474 &  n_444;
assign n_497 = ~x_1478 &  n_441;
assign n_498 = ~n_496 & ~n_497;
assign n_499 =  n_495 &  n_498;
assign n_500 = ~x_1480 &  n_463;
assign n_501 = ~x_1477 &  n_468;
assign n_502 = ~n_500 & ~n_501;
assign n_503 = ~x_1476 &  n_460;
assign n_504 = ~x_1473 &  n_466;
assign n_505 = ~n_503 & ~n_504;
assign n_506 =  n_502 &  n_505;
assign n_507 =  n_499 &  n_506;
assign n_508 =  n_492 & ~n_507;
assign n_509 = ~n_476 & ~n_508;
assign n_510 = ~n_475 & ~n_509;
assign n_511 =  x_401 &  n_510;
assign n_512 = ~x_401 & ~n_510;
assign n_513 = ~n_511 & ~n_512;
assign n_514 =  x_400 & ~n_20;
assign n_515 = ~x_400 &  n_20;
assign n_516 = ~n_514 & ~n_515;
assign n_517 =  x_399 &  n_22;
assign n_518 = ~x_399 & ~n_22;
assign n_519 = ~n_517 & ~n_518;
assign n_520 =  x_398 &  n_3;
assign n_521 = ~x_398 & ~n_3;
assign n_522 = ~n_520 & ~n_521;
assign n_523 =  x_317 & ~x_318;
assign n_524 =  x_3140 &  n_523;
assign n_525 =  x_397 &  n_524;
assign n_526 = ~x_397 & ~n_524;
assign n_527 = ~n_525 & ~n_526;
assign n_528 =  x_396 &  x_3233;
assign n_529 = ~x_396 & ~x_3233;
assign n_530 = ~n_528 & ~n_529;
assign n_531 =  x_307 & ~x_1139;
assign n_532 =  x_317 &  x_1468;
assign n_533 =  x_401 & ~x_1725;
assign n_534 =  n_532 &  n_533;
assign n_535 = ~x_307 & ~x_3158;
assign n_536 = ~n_534 &  n_535;
assign n_537 =  x_395 &  n_536;
assign n_538 = ~n_531 & ~n_537;
assign n_539 =  x_395 & ~n_538;
assign n_540 = ~x_395 &  n_538;
assign n_541 = ~n_539 & ~n_540;
assign n_542 =  x_307 & ~x_1138;
assign n_543 =  x_394 &  n_536;
assign n_544 = ~n_542 & ~n_543;
assign n_545 =  x_394 & ~n_544;
assign n_546 = ~x_394 &  n_544;
assign n_547 = ~n_545 & ~n_546;
assign n_548 =  x_307 & ~x_1137;
assign n_549 =  x_393 &  n_536;
assign n_550 = ~n_548 & ~n_549;
assign n_551 =  x_393 & ~n_550;
assign n_552 = ~x_393 &  n_550;
assign n_553 = ~n_551 & ~n_552;
assign n_554 =  x_307 & ~x_1136;
assign n_555 =  x_392 &  n_536;
assign n_556 = ~n_554 & ~n_555;
assign n_557 =  x_392 & ~n_556;
assign n_558 = ~x_392 &  n_556;
assign n_559 = ~n_557 & ~n_558;
assign n_560 =  x_307 & ~x_1135;
assign n_561 =  x_391 &  n_536;
assign n_562 = ~n_560 & ~n_561;
assign n_563 =  x_391 & ~n_562;
assign n_564 = ~x_391 &  n_562;
assign n_565 = ~n_563 & ~n_564;
assign n_566 =  x_307 & ~x_1134;
assign n_567 =  x_390 &  n_536;
assign n_568 = ~n_566 & ~n_567;
assign n_569 =  x_390 & ~n_568;
assign n_570 = ~x_390 &  n_568;
assign n_571 = ~n_569 & ~n_570;
assign n_572 =  x_307 & ~x_1133;
assign n_573 =  x_389 &  n_536;
assign n_574 = ~n_572 & ~n_573;
assign n_575 =  x_389 & ~n_574;
assign n_576 = ~x_389 &  n_574;
assign n_577 = ~n_575 & ~n_576;
assign n_578 = ~x_388 &  n_536;
assign n_579 =  x_296 &  x_316;
assign n_580 = ~x_1852 &  n_441;
assign n_581 = ~x_1848 &  n_449;
assign n_582 = ~n_580 & ~n_581;
assign n_583 = ~x_1850 &  n_444;
assign n_584 = ~x_1846 &  n_447;
assign n_585 = ~n_583 & ~n_584;
assign n_586 =  n_582 &  n_585;
assign n_587 = ~x_1853 &  n_460;
assign n_588 = ~x_1851 &  n_468;
assign n_589 = ~n_587 & ~n_588;
assign n_590 = ~x_1847 &  n_463;
assign n_591 = ~x_1849 &  n_466;
assign n_592 = ~n_590 & ~n_591;
assign n_593 =  n_589 &  n_592;
assign n_594 =  n_586 &  n_593;
assign n_595 = ~x_1854 &  n_447;
assign n_596 = ~x_1856 &  n_449;
assign n_597 = ~n_595 & ~n_596;
assign n_598 = ~x_1860 &  n_441;
assign n_599 = ~x_1858 &  n_444;
assign n_600 = ~n_598 & ~n_599;
assign n_601 =  n_597 &  n_600;
assign n_602 = ~x_1857 &  n_466;
assign n_603 = ~x_1859 &  n_468;
assign n_604 = ~n_602 & ~n_603;
assign n_605 = ~x_1861 &  n_460;
assign n_606 = ~x_1855 &  n_463;
assign n_607 = ~n_605 & ~n_606;
assign n_608 =  n_604 &  n_607;
assign n_609 =  n_601 &  n_608;
assign n_610 = ~n_594 & ~n_609;
assign n_611 =  n_579 & ~n_610;
assign n_612 = ~n_536 & ~n_611;
assign n_613 =  x_307 & ~x_1132;
assign n_614 =  n_612 & ~n_613;
assign n_615 = ~n_578 & ~n_614;
assign n_616 =  x_388 &  n_615;
assign n_617 = ~x_388 & ~n_615;
assign n_618 = ~n_616 & ~n_617;
assign n_619 =  x_307 & ~x_1131;
assign n_620 =  x_387 &  n_536;
assign n_621 = ~n_619 & ~n_620;
assign n_622 =  x_387 & ~n_621;
assign n_623 = ~x_387 &  n_621;
assign n_624 = ~n_622 & ~n_623;
assign n_625 =  x_307 & ~x_1130;
assign n_626 =  x_386 &  n_536;
assign n_627 = ~n_625 & ~n_626;
assign n_628 =  x_386 & ~n_627;
assign n_629 = ~x_386 &  n_627;
assign n_630 = ~n_628 & ~n_629;
assign n_631 =  x_307 & ~x_1129;
assign n_632 =  x_385 &  n_536;
assign n_633 = ~n_631 & ~n_632;
assign n_634 =  x_385 & ~n_633;
assign n_635 = ~x_385 &  n_633;
assign n_636 = ~n_634 & ~n_635;
assign n_637 =  x_307 & ~x_1128;
assign n_638 =  x_384 &  n_536;
assign n_639 = ~n_637 & ~n_638;
assign n_640 =  x_384 & ~n_639;
assign n_641 = ~x_384 &  n_639;
assign n_642 = ~n_640 & ~n_641;
assign n_643 =  x_307 & ~x_1127;
assign n_644 =  x_383 &  n_536;
assign n_645 = ~n_643 & ~n_644;
assign n_646 =  x_383 & ~n_645;
assign n_647 = ~x_383 &  n_645;
assign n_648 = ~n_646 & ~n_647;
assign n_649 =  x_307 & ~x_1126;
assign n_650 =  x_382 &  n_536;
assign n_651 = ~n_649 & ~n_650;
assign n_652 =  x_382 & ~n_651;
assign n_653 = ~x_382 &  n_651;
assign n_654 = ~n_652 & ~n_653;
assign n_655 =  x_307 & ~x_1125;
assign n_656 =  x_381 &  n_536;
assign n_657 = ~n_655 & ~n_656;
assign n_658 =  x_381 & ~n_657;
assign n_659 = ~x_381 &  n_657;
assign n_660 = ~n_658 & ~n_659;
assign n_661 = ~x_380 &  n_536;
assign n_662 =  x_307 & ~x_1124;
assign n_663 =  n_612 & ~n_662;
assign n_664 = ~n_661 & ~n_663;
assign n_665 =  x_380 &  n_664;
assign n_666 = ~x_380 & ~n_664;
assign n_667 = ~n_665 & ~n_666;
assign n_668 =  x_307 & ~x_1123;
assign n_669 =  x_379 &  n_536;
assign n_670 = ~n_668 & ~n_669;
assign n_671 =  x_379 & ~n_670;
assign n_672 = ~x_379 &  n_670;
assign n_673 = ~n_671 & ~n_672;
assign n_674 =  x_307 & ~x_1122;
assign n_675 =  x_378 &  n_536;
assign n_676 = ~n_674 & ~n_675;
assign n_677 =  x_378 & ~n_676;
assign n_678 = ~x_378 &  n_676;
assign n_679 = ~n_677 & ~n_678;
assign n_680 =  x_307 & ~x_1121;
assign n_681 =  x_377 &  n_536;
assign n_682 = ~n_680 & ~n_681;
assign n_683 =  x_377 & ~n_682;
assign n_684 = ~x_377 &  n_682;
assign n_685 = ~n_683 & ~n_684;
assign n_686 =  x_307 & ~x_1120;
assign n_687 =  x_376 &  n_536;
assign n_688 = ~n_686 & ~n_687;
assign n_689 =  x_376 & ~n_688;
assign n_690 = ~x_376 &  n_688;
assign n_691 = ~n_689 & ~n_690;
assign n_692 =  x_307 & ~x_1119;
assign n_693 =  x_375 &  n_536;
assign n_694 = ~n_692 & ~n_693;
assign n_695 =  x_375 & ~n_694;
assign n_696 = ~x_375 &  n_694;
assign n_697 = ~n_695 & ~n_696;
assign n_698 =  x_307 & ~x_1118;
assign n_699 =  x_374 &  n_536;
assign n_700 = ~n_698 & ~n_699;
assign n_701 =  x_374 & ~n_700;
assign n_702 = ~x_374 &  n_700;
assign n_703 = ~n_701 & ~n_702;
assign n_704 =  x_307 & ~x_1117;
assign n_705 =  x_373 &  n_536;
assign n_706 = ~n_704 & ~n_705;
assign n_707 =  x_373 & ~n_706;
assign n_708 = ~x_373 &  n_706;
assign n_709 = ~n_707 & ~n_708;
assign n_710 = ~x_372 &  n_536;
assign n_711 =  x_307 & ~x_1116;
assign n_712 =  n_612 & ~n_711;
assign n_713 = ~n_710 & ~n_712;
assign n_714 =  x_372 &  n_713;
assign n_715 = ~x_372 & ~n_713;
assign n_716 = ~n_714 & ~n_715;
assign n_717 =  x_307 & ~x_1115;
assign n_718 =  x_371 &  n_536;
assign n_719 = ~n_717 & ~n_718;
assign n_720 =  x_371 & ~n_719;
assign n_721 = ~x_371 &  n_719;
assign n_722 = ~n_720 & ~n_721;
assign n_723 =  x_307 & ~x_1114;
assign n_724 =  x_370 &  n_536;
assign n_725 = ~n_723 & ~n_724;
assign n_726 =  x_370 & ~n_725;
assign n_727 = ~x_370 &  n_725;
assign n_728 = ~n_726 & ~n_727;
assign n_729 =  x_307 & ~x_1113;
assign n_730 =  x_369 &  n_536;
assign n_731 = ~n_729 & ~n_730;
assign n_732 =  x_369 & ~n_731;
assign n_733 = ~x_369 &  n_731;
assign n_734 = ~n_732 & ~n_733;
assign n_735 =  x_307 & ~x_1112;
assign n_736 =  x_368 &  n_536;
assign n_737 = ~n_735 & ~n_736;
assign n_738 =  x_368 & ~n_737;
assign n_739 = ~x_368 &  n_737;
assign n_740 = ~n_738 & ~n_739;
assign n_741 =  x_307 & ~x_1111;
assign n_742 =  x_367 &  n_536;
assign n_743 = ~n_741 & ~n_742;
assign n_744 =  x_367 & ~n_743;
assign n_745 = ~x_367 &  n_743;
assign n_746 = ~n_744 & ~n_745;
assign n_747 =  x_307 & ~x_1110;
assign n_748 =  x_366 &  n_536;
assign n_749 = ~n_747 & ~n_748;
assign n_750 =  x_366 & ~n_749;
assign n_751 = ~x_366 &  n_749;
assign n_752 = ~n_750 & ~n_751;
assign n_753 =  x_307 & ~x_1109;
assign n_754 =  x_365 &  n_536;
assign n_755 = ~n_753 & ~n_754;
assign n_756 =  x_365 & ~n_755;
assign n_757 = ~x_365 &  n_755;
assign n_758 = ~n_756 & ~n_757;
assign n_759 = ~x_364 &  n_536;
assign n_760 =  x_307 & ~x_1108;
assign n_761 =  n_612 & ~n_760;
assign n_762 = ~n_759 & ~n_761;
assign n_763 =  x_364 &  n_762;
assign n_764 = ~x_364 & ~n_762;
assign n_765 = ~n_763 & ~n_764;
assign n_766 =  x_307 & ~x_1107;
assign n_767 =  x_363 &  n_536;
assign n_768 = ~n_766 & ~n_767;
assign n_769 =  x_363 & ~n_768;
assign n_770 = ~x_363 &  n_768;
assign n_771 = ~n_769 & ~n_770;
assign n_772 =  x_307 & ~x_1106;
assign n_773 =  x_362 &  n_536;
assign n_774 = ~n_772 & ~n_773;
assign n_775 =  x_362 & ~n_774;
assign n_776 = ~x_362 &  n_774;
assign n_777 = ~n_775 & ~n_776;
assign n_778 =  x_307 & ~x_1105;
assign n_779 =  x_361 &  n_536;
assign n_780 = ~n_778 & ~n_779;
assign n_781 =  x_361 & ~n_780;
assign n_782 = ~x_361 &  n_780;
assign n_783 = ~n_781 & ~n_782;
assign n_784 =  x_307 & ~x_1104;
assign n_785 =  x_360 &  n_536;
assign n_786 = ~n_784 & ~n_785;
assign n_787 =  x_360 & ~n_786;
assign n_788 = ~x_360 &  n_786;
assign n_789 = ~n_787 & ~n_788;
assign n_790 =  x_307 & ~x_1103;
assign n_791 =  x_359 &  n_536;
assign n_792 = ~n_790 & ~n_791;
assign n_793 =  x_359 & ~n_792;
assign n_794 = ~x_359 &  n_792;
assign n_795 = ~n_793 & ~n_794;
assign n_796 =  x_307 & ~x_1102;
assign n_797 =  x_358 &  n_536;
assign n_798 = ~n_796 & ~n_797;
assign n_799 =  x_358 & ~n_798;
assign n_800 = ~x_358 &  n_798;
assign n_801 = ~n_799 & ~n_800;
assign n_802 =  x_307 & ~x_1101;
assign n_803 =  x_357 &  n_536;
assign n_804 = ~n_802 & ~n_803;
assign n_805 =  x_357 & ~n_804;
assign n_806 = ~x_357 &  n_804;
assign n_807 = ~n_805 & ~n_806;
assign n_808 = ~x_356 &  n_536;
assign n_809 =  x_307 & ~x_1100;
assign n_810 =  n_612 & ~n_809;
assign n_811 = ~n_808 & ~n_810;
assign n_812 =  x_356 &  n_811;
assign n_813 = ~x_356 & ~n_811;
assign n_814 = ~n_812 & ~n_813;
assign n_815 =  x_307 & ~x_1099;
assign n_816 =  x_355 &  n_536;
assign n_817 = ~n_815 & ~n_816;
assign n_818 =  x_355 & ~n_817;
assign n_819 = ~x_355 &  n_817;
assign n_820 = ~n_818 & ~n_819;
assign n_821 =  x_307 & ~x_1098;
assign n_822 =  x_354 &  n_536;
assign n_823 = ~n_821 & ~n_822;
assign n_824 =  x_354 & ~n_823;
assign n_825 = ~x_354 &  n_823;
assign n_826 = ~n_824 & ~n_825;
assign n_827 =  x_307 & ~x_1097;
assign n_828 =  x_353 &  n_536;
assign n_829 = ~n_827 & ~n_828;
assign n_830 =  x_353 & ~n_829;
assign n_831 = ~x_353 &  n_829;
assign n_832 = ~n_830 & ~n_831;
assign n_833 =  x_307 & ~x_1096;
assign n_834 =  x_352 &  n_536;
assign n_835 = ~n_833 & ~n_834;
assign n_836 =  x_352 & ~n_835;
assign n_837 = ~x_352 &  n_835;
assign n_838 = ~n_836 & ~n_837;
assign n_839 =  x_307 & ~x_1095;
assign n_840 =  x_351 &  n_536;
assign n_841 = ~n_839 & ~n_840;
assign n_842 =  x_351 & ~n_841;
assign n_843 = ~x_351 &  n_841;
assign n_844 = ~n_842 & ~n_843;
assign n_845 =  x_307 & ~x_1094;
assign n_846 =  x_350 &  n_536;
assign n_847 = ~n_845 & ~n_846;
assign n_848 =  x_350 & ~n_847;
assign n_849 = ~x_350 &  n_847;
assign n_850 = ~n_848 & ~n_849;
assign n_851 =  x_307 & ~x_1093;
assign n_852 =  x_349 &  n_536;
assign n_853 = ~n_851 & ~n_852;
assign n_854 =  x_349 & ~n_853;
assign n_855 = ~x_349 &  n_853;
assign n_856 = ~n_854 & ~n_855;
assign n_857 = ~x_348 &  n_536;
assign n_858 =  x_307 & ~x_1092;
assign n_859 =  n_612 & ~n_858;
assign n_860 = ~n_857 & ~n_859;
assign n_861 =  x_348 &  n_860;
assign n_862 = ~x_348 & ~n_860;
assign n_863 = ~n_861 & ~n_862;
assign n_864 =  x_307 & ~x_1091;
assign n_865 =  x_347 &  n_536;
assign n_866 = ~n_864 & ~n_865;
assign n_867 =  x_347 & ~n_866;
assign n_868 = ~x_347 &  n_866;
assign n_869 = ~n_867 & ~n_868;
assign n_870 =  x_307 & ~x_1090;
assign n_871 =  x_346 &  n_536;
assign n_872 = ~n_870 & ~n_871;
assign n_873 =  x_346 & ~n_872;
assign n_874 = ~x_346 &  n_872;
assign n_875 = ~n_873 & ~n_874;
assign n_876 =  x_307 & ~x_1089;
assign n_877 =  x_345 &  n_536;
assign n_878 = ~n_876 & ~n_877;
assign n_879 =  x_345 & ~n_878;
assign n_880 = ~x_345 &  n_878;
assign n_881 = ~n_879 & ~n_880;
assign n_882 =  x_307 & ~x_1088;
assign n_883 =  x_344 &  n_536;
assign n_884 = ~n_882 & ~n_883;
assign n_885 =  x_344 & ~n_884;
assign n_886 = ~x_344 &  n_884;
assign n_887 = ~n_885 & ~n_886;
assign n_888 =  x_307 & ~x_1087;
assign n_889 =  x_343 &  n_536;
assign n_890 = ~n_888 & ~n_889;
assign n_891 =  x_343 & ~n_890;
assign n_892 = ~x_343 &  n_890;
assign n_893 = ~n_891 & ~n_892;
assign n_894 =  x_307 & ~x_1086;
assign n_895 =  x_342 &  n_536;
assign n_896 = ~n_894 & ~n_895;
assign n_897 =  x_342 & ~n_896;
assign n_898 = ~x_342 &  n_896;
assign n_899 = ~n_897 & ~n_898;
assign n_900 =  x_307 & ~x_1085;
assign n_901 =  x_341 &  n_536;
assign n_902 = ~n_900 & ~n_901;
assign n_903 =  x_341 & ~n_902;
assign n_904 = ~x_341 &  n_902;
assign n_905 = ~n_903 & ~n_904;
assign n_906 = ~x_340 &  n_536;
assign n_907 =  x_307 & ~x_1084;
assign n_908 =  n_612 & ~n_907;
assign n_909 = ~n_906 & ~n_908;
assign n_910 =  x_340 &  n_909;
assign n_911 = ~x_340 & ~n_909;
assign n_912 = ~n_910 & ~n_911;
assign n_913 =  x_339 &  n_536;
assign n_914 =  x_1468 & ~n_536;
assign n_915 =  x_338 &  x_401;
assign n_916 =  x_307 & ~x_1075;
assign n_917 = ~n_915 & ~n_916;
assign n_918 =  n_914 & ~n_917;
assign n_919 = ~n_913 & ~n_918;
assign n_920 =  x_339 & ~n_919;
assign n_921 = ~x_339 &  n_919;
assign n_922 = ~n_920 & ~n_921;
assign n_923 =  x_316 &  x_1725;
assign n_924 = ~n_436 & ~n_923;
assign n_925 =  x_338 &  n_924;
assign n_926 = ~x_1714 &  n_468;
assign n_927 = ~x_1710 &  n_463;
assign n_928 = ~x_1712 &  n_466;
assign n_929 = ~n_927 & ~n_928;
assign n_930 = ~n_926 &  n_929;
assign n_931 = ~x_1715 &  n_441;
assign n_932 = ~x_1711 &  n_449;
assign n_933 = ~x_1713 &  n_444;
assign n_934 = ~n_932 & ~n_933;
assign n_935 = ~n_931 &  n_934;
assign n_936 = ~x_1716 &  n_460;
assign n_937 = ~x_1709 &  n_447;
assign n_938 =  n_436 & ~n_937;
assign n_939 = ~n_936 &  n_938;
assign n_940 =  n_935 &  n_939;
assign n_941 =  n_930 &  n_940;
assign n_942 = ~n_925 & ~n_941;
assign n_943 =  x_338 & ~n_942;
assign n_944 = ~x_338 &  n_942;
assign n_945 = ~n_943 & ~n_944;
assign n_946 =  x_337 &  n_536;
assign n_947 =  x_336 &  x_401;
assign n_948 =  x_307 & ~x_1066;
assign n_949 = ~n_947 & ~n_948;
assign n_950 =  n_914 & ~n_949;
assign n_951 = ~n_946 & ~n_950;
assign n_952 =  x_337 & ~n_951;
assign n_953 = ~x_337 &  n_951;
assign n_954 = ~n_952 & ~n_953;
assign n_955 =  x_336 &  n_924;
assign n_956 = ~x_1704 &  n_466;
assign n_957 = ~x_1708 &  n_460;
assign n_958 = ~x_1702 &  n_463;
assign n_959 = ~n_957 & ~n_958;
assign n_960 = ~n_956 &  n_959;
assign n_961 = ~x_1703 &  n_449;
assign n_962 = ~x_1707 &  n_441;
assign n_963 = ~x_1701 &  n_447;
assign n_964 = ~n_962 & ~n_963;
assign n_965 = ~n_961 &  n_964;
assign n_966 = ~x_1706 &  n_468;
assign n_967 = ~x_1705 &  n_444;
assign n_968 =  n_436 & ~n_967;
assign n_969 = ~n_966 &  n_968;
assign n_970 =  n_965 &  n_969;
assign n_971 =  n_960 &  n_970;
assign n_972 = ~n_955 & ~n_971;
assign n_973 =  x_336 & ~n_972;
assign n_974 = ~x_336 &  n_972;
assign n_975 = ~n_973 & ~n_974;
assign n_976 =  x_335 &  n_536;
assign n_977 =  x_334 &  x_401;
assign n_978 =  x_307 & ~x_1057;
assign n_979 = ~n_977 & ~n_978;
assign n_980 =  n_914 & ~n_979;
assign n_981 = ~n_976 & ~n_980;
assign n_982 =  x_335 & ~n_981;
assign n_983 = ~x_335 &  n_981;
assign n_984 = ~n_982 & ~n_983;
assign n_985 =  x_334 &  n_924;
assign n_986 = ~x_1700 &  n_460;
assign n_987 = ~x_1696 &  n_466;
assign n_988 = ~x_1694 &  n_463;
assign n_989 = ~n_987 & ~n_988;
assign n_990 = ~n_986 &  n_989;
assign n_991 = ~x_1697 &  n_444;
assign n_992 = ~x_1699 &  n_441;
assign n_993 = ~x_1695 &  n_449;
assign n_994 = ~n_992 & ~n_993;
assign n_995 = ~n_991 &  n_994;
assign n_996 = ~x_1698 &  n_468;
assign n_997 = ~x_1693 &  n_447;
assign n_998 =  n_436 & ~n_997;
assign n_999 = ~n_996 &  n_998;
assign n_1000 =  n_995 &  n_999;
assign n_1001 =  n_990 &  n_1000;
assign n_1002 = ~n_985 & ~n_1001;
assign n_1003 =  x_334 & ~n_1002;
assign n_1004 = ~x_334 &  n_1002;
assign n_1005 = ~n_1003 & ~n_1004;
assign n_1006 =  x_333 &  n_536;
assign n_1007 =  x_332 &  x_401;
assign n_1008 =  x_307 & ~x_1048;
assign n_1009 = ~n_1007 & ~n_1008;
assign n_1010 =  n_914 & ~n_1009;
assign n_1011 = ~n_1006 & ~n_1010;
assign n_1012 =  x_333 & ~n_1011;
assign n_1013 = ~x_333 &  n_1011;
assign n_1014 = ~n_1012 & ~n_1013;
assign n_1015 =  x_332 &  n_924;
assign n_1016 = ~x_1690 &  n_468;
assign n_1017 = ~x_1688 &  n_466;
assign n_1018 = ~x_1686 &  n_463;
assign n_1019 = ~n_1017 & ~n_1018;
assign n_1020 = ~n_1016 &  n_1019;
assign n_1021 = ~x_1691 &  n_441;
assign n_1022 = ~x_1689 &  n_444;
assign n_1023 = ~x_1687 &  n_449;
assign n_1024 = ~n_1022 & ~n_1023;
assign n_1025 = ~n_1021 &  n_1024;
assign n_1026 = ~x_1692 &  n_460;
assign n_1027 = ~x_1685 &  n_447;
assign n_1028 =  n_436 & ~n_1027;
assign n_1029 = ~n_1026 &  n_1028;
assign n_1030 =  n_1025 &  n_1029;
assign n_1031 =  n_1020 &  n_1030;
assign n_1032 = ~n_1015 & ~n_1031;
assign n_1033 =  x_332 & ~n_1032;
assign n_1034 = ~x_332 &  n_1032;
assign n_1035 = ~n_1033 & ~n_1034;
assign n_1036 =  x_331 &  n_536;
assign n_1037 =  x_330 &  x_401;
assign n_1038 =  x_307 & ~x_1039;
assign n_1039 = ~n_1037 & ~n_1038;
assign n_1040 =  n_914 & ~n_1039;
assign n_1041 = ~n_1036 & ~n_1040;
assign n_1042 =  x_331 & ~n_1041;
assign n_1043 = ~x_331 &  n_1041;
assign n_1044 = ~n_1042 & ~n_1043;
assign n_1045 =  x_330 &  n_924;
assign n_1046 = ~x_1678 &  n_463;
assign n_1047 = ~x_1682 &  n_468;
assign n_1048 = ~x_1684 &  n_460;
assign n_1049 = ~n_1047 & ~n_1048;
assign n_1050 = ~n_1046 &  n_1049;
assign n_1051 = ~x_1683 &  n_441;
assign n_1052 = ~x_1679 &  n_449;
assign n_1053 = ~x_1677 &  n_447;
assign n_1054 = ~n_1052 & ~n_1053;
assign n_1055 = ~n_1051 &  n_1054;
assign n_1056 = ~x_1680 &  n_466;
assign n_1057 = ~x_1681 &  n_444;
assign n_1058 =  n_436 & ~n_1057;
assign n_1059 = ~n_1056 &  n_1058;
assign n_1060 =  n_1055 &  n_1059;
assign n_1061 =  n_1050 &  n_1060;
assign n_1062 = ~n_1045 & ~n_1061;
assign n_1063 =  x_330 & ~n_1062;
assign n_1064 = ~x_330 &  n_1062;
assign n_1065 = ~n_1063 & ~n_1064;
assign n_1066 =  x_329 &  n_536;
assign n_1067 =  x_328 &  x_401;
assign n_1068 =  x_307 & ~x_1030;
assign n_1069 = ~n_1067 & ~n_1068;
assign n_1070 =  n_914 & ~n_1069;
assign n_1071 = ~n_1066 & ~n_1070;
assign n_1072 =  x_329 & ~n_1071;
assign n_1073 = ~x_329 &  n_1071;
assign n_1074 = ~n_1072 & ~n_1073;
assign n_1075 =  x_328 &  n_924;
assign n_1076 = ~x_1676 &  n_460;
assign n_1077 = ~x_1672 &  n_466;
assign n_1078 = ~x_1670 &  n_463;
assign n_1079 = ~n_1077 & ~n_1078;
assign n_1080 = ~n_1076 &  n_1079;
assign n_1081 = ~x_1675 &  n_441;
assign n_1082 = ~x_1673 &  n_444;
assign n_1083 = ~x_1671 &  n_449;
assign n_1084 = ~n_1082 & ~n_1083;
assign n_1085 = ~n_1081 &  n_1084;
assign n_1086 = ~x_1674 &  n_468;
assign n_1087 = ~x_1669 &  n_447;
assign n_1088 =  n_436 & ~n_1087;
assign n_1089 = ~n_1086 &  n_1088;
assign n_1090 =  n_1085 &  n_1089;
assign n_1091 =  n_1080 &  n_1090;
assign n_1092 = ~n_1075 & ~n_1091;
assign n_1093 =  x_328 & ~n_1092;
assign n_1094 = ~x_328 &  n_1092;
assign n_1095 = ~n_1093 & ~n_1094;
assign n_1096 =  x_327 &  n_536;
assign n_1097 =  x_326 &  x_401;
assign n_1098 =  x_307 &  x_325;
assign n_1099 = ~n_1097 & ~n_1098;
assign n_1100 = ~n_1099 &  n_914;
assign n_1101 = ~n_1096 & ~n_1100;
assign n_1102 =  x_327 & ~n_1101;
assign n_1103 = ~x_327 &  n_1101;
assign n_1104 = ~n_1102 & ~n_1103;
assign n_1105 =  x_326 &  n_924;
assign n_1106 = ~x_1662 &  n_463;
assign n_1107 = ~x_1668 &  n_460;
assign n_1108 = ~x_1664 &  n_466;
assign n_1109 = ~n_1107 & ~n_1108;
assign n_1110 = ~n_1106 &  n_1109;
assign n_1111 = ~x_1665 &  n_444;
assign n_1112 = ~x_1663 &  n_449;
assign n_1113 = ~x_1667 &  n_441;
assign n_1114 = ~n_1112 & ~n_1113;
assign n_1115 = ~n_1111 &  n_1114;
assign n_1116 = ~x_1666 &  n_468;
assign n_1117 = ~x_1661 &  n_447;
assign n_1118 =  n_436 & ~n_1117;
assign n_1119 = ~n_1116 &  n_1118;
assign n_1120 =  n_1115 &  n_1119;
assign n_1121 =  n_1110 &  n_1120;
assign n_1122 = ~n_1105 & ~n_1121;
assign n_1123 =  x_326 & ~n_1122;
assign n_1124 = ~x_326 &  n_1122;
assign n_1125 = ~n_1123 & ~n_1124;
assign n_1126 =  x_1652 & ~n_923;
assign n_1127 =  x_325 &  n_1126;
assign n_1128 = ~x_1652 &  n_609;
assign n_1129 = ~n_1127 & ~n_1128;
assign n_1130 =  x_325 & ~n_1129;
assign n_1131 = ~x_325 &  n_1129;
assign n_1132 = ~n_1130 & ~n_1131;
assign n_1133 = ~x_324 &  n_536;
assign n_1134 =  x_323 &  x_401;
assign n_1135 =  x_307 &  x_322;
assign n_1136 = ~n_1134 & ~n_1135;
assign n_1137 =  x_1468 & ~n_1136;
assign n_1138 = ~n_1137 &  n_612;
assign n_1139 = ~n_1133 & ~n_1138;
assign n_1140 =  x_324 &  n_1139;
assign n_1141 = ~x_324 & ~n_1139;
assign n_1142 = ~n_1140 & ~n_1141;
assign n_1143 =  x_323 &  n_924;
assign n_1144 = ~x_1660 &  n_460;
assign n_1145 = ~x_1658 &  n_468;
assign n_1146 = ~x_1654 &  n_463;
assign n_1147 = ~n_1145 & ~n_1146;
assign n_1148 = ~n_1144 &  n_1147;
assign n_1149 = ~x_1655 &  n_449;
assign n_1150 = ~x_1653 &  n_447;
assign n_1151 = ~x_1657 &  n_444;
assign n_1152 = ~n_1150 & ~n_1151;
assign n_1153 = ~n_1149 &  n_1152;
assign n_1154 = ~x_1656 &  n_466;
assign n_1155 = ~x_1659 &  n_441;
assign n_1156 =  n_436 & ~n_1155;
assign n_1157 = ~n_1154 &  n_1156;
assign n_1158 =  n_1153 &  n_1157;
assign n_1159 =  n_1148 &  n_1158;
assign n_1160 = ~n_1143 & ~n_1159;
assign n_1161 =  x_323 & ~n_1160;
assign n_1162 = ~x_323 &  n_1160;
assign n_1163 = ~n_1161 & ~n_1162;
assign n_1164 =  x_322 &  n_1126;
assign n_1165 = ~x_1652 &  n_594;
assign n_1166 = ~n_1164 & ~n_1165;
assign n_1167 =  x_322 & ~n_1166;
assign n_1168 = ~x_322 &  n_1166;
assign n_1169 = ~n_1167 & ~n_1168;
assign n_1170 = ~x_316 & ~n_532;
assign n_1171 = ~x_1732 &  n_1170;
assign n_1172 = ~x_321 & ~n_532;
assign n_1173 = ~n_579 & ~n_1172;
assign n_1174 = ~n_1171 &  n_1173;
assign n_1175 =  x_321 &  n_1174;
assign n_1176 = ~x_321 & ~n_1174;
assign n_1177 = ~n_1175 & ~n_1176;
assign n_1178 =  x_1472 & ~n_507;
assign n_1179 =  x_320 &  n_1178;
assign n_1180 =  x_401 &  x_1725;
assign n_1181 =  n_532 &  n_1180;
assign n_1182 = ~x_1469 & ~n_1181;
assign n_1183 = ~n_923 &  n_1182;
assign n_1184 = ~x_304 & ~n_923;
assign n_1185 = ~n_1180 &  n_1184;
assign n_1186 = ~n_1183 & ~n_1185;
assign n_1187 = ~n_1179 & ~n_1186;
assign n_1188 =  n_472 & ~n_491;
assign n_1189 =  n_1178 &  n_1188;
assign n_1190 = ~n_1187 & ~n_1189;
assign n_1191 =  x_1745 &  x_1746;
assign n_1192 =  x_1747 &  n_1191;
assign n_1193 = ~x_320 & ~n_1192;
assign n_1194 = ~n_1186 &  n_1193;
assign n_1195 = ~n_1190 & ~n_1194;
assign n_1196 =  x_320 &  n_1195;
assign n_1197 = ~x_320 & ~n_1195;
assign n_1198 = ~n_1196 & ~n_1197;
assign n_1199 =  x_319 &  n_1186;
assign n_1200 = ~x_319 & ~n_1186;
assign n_1201 = ~n_1199 & ~n_1200;
assign n_1202 =  x_296 & ~n_1170;
assign n_1203 =  x_318 & ~n_1171;
assign n_1204 = ~n_1202 & ~n_1203;
assign n_1205 =  x_318 & ~n_1204;
assign n_1206 = ~x_318 &  n_1204;
assign n_1207 = ~n_1205 & ~n_1206;
assign n_1208 = ~x_1481 & ~n_1183;
assign n_1209 = ~x_317 & ~n_1192;
assign n_1210 =  n_1183 &  n_1209;
assign n_1211 = ~n_1208 & ~n_1210;
assign n_1212 =  x_317 &  n_1211;
assign n_1213 = ~x_317 & ~n_1211;
assign n_1214 = ~n_1212 & ~n_1213;
assign n_1215 =  n_491 &  n_1179;
assign n_1216 =  x_296 &  x_317;
assign n_1217 =  x_401 &  n_1216;
assign n_1218 = ~x_316 & ~n_1217;
assign n_1219 = ~x_1725 & ~n_1218;
assign n_1220 = ~n_1215 & ~n_1219;
assign n_1221 =  x_316 & ~n_1220;
assign n_1222 = ~x_316 &  n_1220;
assign n_1223 = ~n_1221 & ~n_1222;
assign n_1224 = ~x_315 & ~n_923;
assign n_1225 = ~n_1181 &  n_1224;
assign n_1226 = ~x_1472 & ~n_1225;
assign n_1227 =  x_315 &  n_1226;
assign n_1228 = ~x_315 & ~n_1226;
assign n_1229 = ~n_1227 & ~n_1228;
assign n_1230 =  x_314 &  x_2550;
assign n_1231 = ~x_314 & ~x_2550;
assign n_1232 = ~n_1230 & ~n_1231;
assign n_1233 =  x_313 &  x_1771;
assign n_1234 = ~x_313 & ~x_1771;
assign n_1235 = ~n_1233 & ~n_1234;
assign n_1236 =  x_312 &  n_1192;
assign n_1237 = ~x_312 & ~n_1192;
assign n_1238 = ~n_1236 & ~n_1237;
assign n_1239 =  x_311 &  x_1764;
assign n_1240 = ~x_311 & ~x_1764;
assign n_1241 = ~n_1239 & ~n_1240;
assign n_1242 =  x_310 &  x_1753;
assign n_1243 = ~x_310 & ~x_1753;
assign n_1244 = ~n_1242 & ~n_1243;
assign n_1245 =  x_309 &  x_1748;
assign n_1246 = ~x_309 & ~x_1748;
assign n_1247 = ~n_1245 & ~n_1246;
assign n_1248 = ~x_307 & ~n_1180;
assign n_1249 = ~n_1182 & ~n_1248;
assign n_1250 = ~x_1472 & ~n_923;
assign n_1251 = ~n_1249 &  n_1250;
assign n_1252 =  x_308 &  n_1251;
assign n_1253 =  n_1179 & ~n_1188;
assign n_1254 = ~x_304 &  x_307;
assign n_1255 = ~n_1254 & ~n_579;
assign n_1256 = ~n_1253 &  n_1255;
assign n_1257 = ~n_1251 & ~n_1256;
assign n_1258 = ~n_1252 & ~n_1257;
assign n_1259 =  x_308 & ~n_1258;
assign n_1260 = ~x_308 &  n_1258;
assign n_1261 = ~n_1259 & ~n_1260;
assign n_1262 = ~x_307 &  x_1469;
assign n_1263 =  x_307 &  n_1262;
assign n_1264 = ~x_307 & ~n_1262;
assign n_1265 = ~n_1263 & ~n_1264;
assign n_1266 = ~n_476 & ~n_492;
assign n_1267 =  x_306 & ~n_1266;
assign n_1268 = ~x_306 &  n_1266;
assign n_1269 = ~n_1267 & ~n_1268;
assign n_1270 =  x_305 & ~n_475;
assign n_1271 = ~x_305 &  n_475;
assign n_1272 = ~n_1270 & ~n_1271;
assign n_1273 =  x_304 &  x_1471;
assign n_1274 = ~x_304 & ~x_1471;
assign n_1275 = ~n_1273 & ~n_1274;
assign n_1276 =  x_300 & ~x_301;
assign n_1277 = ~x_302 & ~x_303;
assign n_1278 =  x_301 & ~n_1277;
assign n_1279 =  x_313 & ~n_1278;
assign n_1280 = ~n_1276 &  n_1279;
assign n_1281 = ~x_300 &  n_1277;
assign n_1282 =  x_301 & ~x_313;
assign n_1283 = ~n_1281 &  n_1282;
assign n_1284 = ~n_1280 & ~n_1283;
assign n_1285 =  x_302 &  x_303;
assign n_1286 = ~n_1285 & ~n_1277;
assign n_1287 =  x_300 &  x_301;
assign n_1288 = ~n_1286 & ~n_1287;
assign n_1289 = ~n_1282 & ~n_1288;
assign n_1290 = ~n_1284 &  n_1289;
assign n_1291 =  x_303 &  n_1284;
assign n_1292 =  n_1283 & ~n_1286;
assign n_1293 = ~n_1291 & ~n_1292;
assign n_1294 = ~n_1290 &  n_1293;
assign n_1295 =  x_303 & ~n_1294;
assign n_1296 = ~x_303 &  n_1294;
assign n_1297 = ~n_1295 & ~n_1296;
assign n_1298 = ~x_302 & ~n_1284;
assign n_1299 =  x_302 &  n_1284;
assign n_1300 = ~n_1298 & ~n_1299;
assign n_1301 =  x_302 & ~n_1300;
assign n_1302 = ~x_302 &  n_1300;
assign n_1303 = ~n_1301 & ~n_1302;
assign n_1304 =  x_301 &  x_320;
assign n_1305 = ~x_301 & ~x_320;
assign n_1306 = ~n_1304 & ~n_1305;
assign n_1307 =  n_1285 &  n_1279;
assign n_1308 = ~n_1276 & ~n_1307;
assign n_1309 =  x_300 & ~n_1308;
assign n_1310 = ~x_300 &  n_1308;
assign n_1311 = ~n_1309 & ~n_1310;
assign n_1312 =  x_299 &  n_459;
assign n_1313 = ~x_299 & ~n_459;
assign n_1314 = ~n_1312 & ~n_1313;
assign n_1315 =  x_298 &  n_455;
assign n_1316 = ~x_298 & ~n_455;
assign n_1317 = ~n_1315 & ~n_1316;
assign n_1318 =  x_297 &  n_439;
assign n_1319 = ~x_297 & ~n_439;
assign n_1320 = ~n_1318 & ~n_1319;
assign n_1321 = ~x_1482 & ~n_1179;
assign n_1322 =  x_296 & ~n_1321;
assign n_1323 = ~x_296 &  n_1321;
assign n_1324 = ~n_1322 & ~n_1323;
assign n_1325 =  i_10 &  x_295;
assign n_1326 =  x_294 &  n_1325;
assign n_1327 =  i_9 &  x_295;
assign n_1328 = ~n_1325 & ~n_1327;
assign n_1329 =  x_228 &  n_1328;
assign n_1330 = ~x_3104 &  n_1329;
assign n_1331 = ~n_1326 & ~n_1330;
assign n_1332 =  x_294 & ~n_1331;
assign n_1333 = ~x_294 &  n_1331;
assign n_1334 = ~n_1332 & ~n_1333;
assign n_1335 =  x_293 &  n_1325;
assign n_1336 = ~x_3103 &  n_1329;
assign n_1337 = ~n_1335 & ~n_1336;
assign n_1338 =  x_293 & ~n_1337;
assign n_1339 = ~x_293 &  n_1337;
assign n_1340 = ~n_1338 & ~n_1339;
assign n_1341 =  x_292 &  n_1325;
assign n_1342 = ~x_3102 &  n_1329;
assign n_1343 = ~n_1341 & ~n_1342;
assign n_1344 =  x_292 & ~n_1343;
assign n_1345 = ~x_292 &  n_1343;
assign n_1346 = ~n_1344 & ~n_1345;
assign n_1347 =  x_291 &  n_1325;
assign n_1348 = ~x_3101 &  n_1329;
assign n_1349 = ~n_1347 & ~n_1348;
assign n_1350 =  x_291 & ~n_1349;
assign n_1351 = ~x_291 &  n_1349;
assign n_1352 = ~n_1350 & ~n_1351;
assign n_1353 =  x_290 &  n_1325;
assign n_1354 = ~x_3100 &  n_1329;
assign n_1355 = ~n_1353 & ~n_1354;
assign n_1356 =  x_290 & ~n_1355;
assign n_1357 = ~x_290 &  n_1355;
assign n_1358 = ~n_1356 & ~n_1357;
assign n_1359 =  x_289 &  n_1325;
assign n_1360 = ~x_3099 &  n_1329;
assign n_1361 = ~n_1359 & ~n_1360;
assign n_1362 =  x_289 & ~n_1361;
assign n_1363 = ~x_289 &  n_1361;
assign n_1364 = ~n_1362 & ~n_1363;
assign n_1365 =  x_288 &  n_1325;
assign n_1366 = ~x_3098 &  n_1329;
assign n_1367 = ~n_1365 & ~n_1366;
assign n_1368 =  x_288 & ~n_1367;
assign n_1369 = ~x_288 &  n_1367;
assign n_1370 = ~n_1368 & ~n_1369;
assign n_1371 =  x_287 &  n_1325;
assign n_1372 = ~x_3097 &  n_1329;
assign n_1373 = ~n_1371 & ~n_1372;
assign n_1374 =  x_287 & ~n_1373;
assign n_1375 = ~x_287 &  n_1373;
assign n_1376 = ~n_1374 & ~n_1375;
assign n_1377 =  x_286 &  n_1325;
assign n_1378 = ~x_3096 &  n_1329;
assign n_1379 = ~n_1377 & ~n_1378;
assign n_1380 =  x_286 & ~n_1379;
assign n_1381 = ~x_286 &  n_1379;
assign n_1382 = ~n_1380 & ~n_1381;
assign n_1383 =  x_285 &  n_1325;
assign n_1384 = ~x_3095 &  n_1329;
assign n_1385 = ~n_1383 & ~n_1384;
assign n_1386 =  x_285 & ~n_1385;
assign n_1387 = ~x_285 &  n_1385;
assign n_1388 = ~n_1386 & ~n_1387;
assign n_1389 =  x_284 &  n_1325;
assign n_1390 = ~x_3094 &  n_1329;
assign n_1391 = ~n_1389 & ~n_1390;
assign n_1392 =  x_284 & ~n_1391;
assign n_1393 = ~x_284 &  n_1391;
assign n_1394 = ~n_1392 & ~n_1393;
assign n_1395 =  x_283 &  n_1325;
assign n_1396 = ~x_3093 &  n_1329;
assign n_1397 = ~n_1395 & ~n_1396;
assign n_1398 =  x_283 & ~n_1397;
assign n_1399 = ~x_283 &  n_1397;
assign n_1400 = ~n_1398 & ~n_1399;
assign n_1401 =  x_282 &  n_1325;
assign n_1402 = ~x_3092 &  n_1329;
assign n_1403 = ~n_1401 & ~n_1402;
assign n_1404 =  x_282 & ~n_1403;
assign n_1405 = ~x_282 &  n_1403;
assign n_1406 = ~n_1404 & ~n_1405;
assign n_1407 =  x_281 &  n_1325;
assign n_1408 = ~x_3091 &  n_1329;
assign n_1409 = ~n_1407 & ~n_1408;
assign n_1410 =  x_281 & ~n_1409;
assign n_1411 = ~x_281 &  n_1409;
assign n_1412 = ~n_1410 & ~n_1411;
assign n_1413 =  x_280 &  n_1325;
assign n_1414 = ~x_3090 &  n_1329;
assign n_1415 = ~n_1413 & ~n_1414;
assign n_1416 =  x_280 & ~n_1415;
assign n_1417 = ~x_280 &  n_1415;
assign n_1418 = ~n_1416 & ~n_1417;
assign n_1419 =  x_279 &  n_1325;
assign n_1420 = ~x_3089 &  n_1329;
assign n_1421 = ~n_1419 & ~n_1420;
assign n_1422 =  x_279 & ~n_1421;
assign n_1423 = ~x_279 &  n_1421;
assign n_1424 = ~n_1422 & ~n_1423;
assign n_1425 =  x_278 &  n_1325;
assign n_1426 = ~x_3088 &  n_1329;
assign n_1427 = ~n_1425 & ~n_1426;
assign n_1428 =  x_278 & ~n_1427;
assign n_1429 = ~x_278 &  n_1427;
assign n_1430 = ~n_1428 & ~n_1429;
assign n_1431 =  x_277 &  n_1325;
assign n_1432 = ~x_3087 &  n_1329;
assign n_1433 = ~n_1431 & ~n_1432;
assign n_1434 =  x_277 & ~n_1433;
assign n_1435 = ~x_277 &  n_1433;
assign n_1436 = ~n_1434 & ~n_1435;
assign n_1437 =  x_276 &  n_1325;
assign n_1438 = ~x_3086 &  n_1329;
assign n_1439 = ~n_1437 & ~n_1438;
assign n_1440 =  x_276 & ~n_1439;
assign n_1441 = ~x_276 &  n_1439;
assign n_1442 = ~n_1440 & ~n_1441;
assign n_1443 =  x_275 &  n_1325;
assign n_1444 = ~x_3085 &  n_1329;
assign n_1445 = ~n_1443 & ~n_1444;
assign n_1446 =  x_275 & ~n_1445;
assign n_1447 = ~x_275 &  n_1445;
assign n_1448 = ~n_1446 & ~n_1447;
assign n_1449 =  x_274 &  n_1325;
assign n_1450 = ~x_3084 &  n_1329;
assign n_1451 = ~n_1449 & ~n_1450;
assign n_1452 =  x_274 & ~n_1451;
assign n_1453 = ~x_274 &  n_1451;
assign n_1454 = ~n_1452 & ~n_1453;
assign n_1455 =  x_273 &  n_1325;
assign n_1456 = ~x_3083 &  n_1329;
assign n_1457 = ~n_1455 & ~n_1456;
assign n_1458 =  x_273 & ~n_1457;
assign n_1459 = ~x_273 &  n_1457;
assign n_1460 = ~n_1458 & ~n_1459;
assign n_1461 =  x_272 &  n_1325;
assign n_1462 = ~x_3082 &  n_1329;
assign n_1463 = ~n_1461 & ~n_1462;
assign n_1464 =  x_272 & ~n_1463;
assign n_1465 = ~x_272 &  n_1463;
assign n_1466 = ~n_1464 & ~n_1465;
assign n_1467 =  x_271 &  n_1325;
assign n_1468 = ~x_3081 &  n_1329;
assign n_1469 = ~n_1467 & ~n_1468;
assign n_1470 =  x_271 & ~n_1469;
assign n_1471 = ~x_271 &  n_1469;
assign n_1472 = ~n_1470 & ~n_1471;
assign n_1473 =  x_270 &  n_1325;
assign n_1474 = ~x_3080 &  n_1329;
assign n_1475 = ~n_1473 & ~n_1474;
assign n_1476 =  x_270 & ~n_1475;
assign n_1477 = ~x_270 &  n_1475;
assign n_1478 = ~n_1476 & ~n_1477;
assign n_1479 =  x_269 &  n_1325;
assign n_1480 = ~x_3079 &  n_1329;
assign n_1481 = ~n_1479 & ~n_1480;
assign n_1482 =  x_269 & ~n_1481;
assign n_1483 = ~x_269 &  n_1481;
assign n_1484 = ~n_1482 & ~n_1483;
assign n_1485 =  x_268 &  n_1325;
assign n_1486 = ~x_3078 &  n_1329;
assign n_1487 = ~n_1485 & ~n_1486;
assign n_1488 =  x_268 & ~n_1487;
assign n_1489 = ~x_268 &  n_1487;
assign n_1490 = ~n_1488 & ~n_1489;
assign n_1491 =  x_267 &  n_1325;
assign n_1492 = ~x_3077 &  n_1329;
assign n_1493 = ~n_1491 & ~n_1492;
assign n_1494 =  x_267 & ~n_1493;
assign n_1495 = ~x_267 &  n_1493;
assign n_1496 = ~n_1494 & ~n_1495;
assign n_1497 =  x_265 &  n_1325;
assign n_1498 = ~x_266 &  n_1329;
assign n_1499 = ~n_1497 & ~n_1498;
assign n_1500 =  x_263 & ~n_1325;
assign n_1501 = ~x_263 & ~n_1328;
assign n_1502 = ~n_1500 & ~n_1501;
assign n_1503 =  x_264 &  n_1325;
assign n_1504 =  x_3076 &  n_1329;
assign n_1505 = ~n_1503 & ~n_1504;
assign n_1506 =  n_1502 & ~n_1505;
assign n_1507 =  n_1499 & ~n_1506;
assign n_1508 = ~n_1499 &  n_1506;
assign n_1509 = ~n_1507 & ~n_1508;
assign n_1510 =  x_266 & ~n_1509;
assign n_1511 = ~x_266 &  n_1509;
assign n_1512 = ~n_1510 & ~n_1511;
assign n_1513 =  x_265 & ~n_1499;
assign n_1514 = ~x_265 &  n_1499;
assign n_1515 = ~n_1513 & ~n_1514;
assign n_1516 =  x_264 & ~n_1505;
assign n_1517 = ~x_264 &  n_1505;
assign n_1518 = ~n_1516 & ~n_1517;
assign n_1519 =  x_263 &  n_1502;
assign n_1520 = ~x_263 & ~n_1502;
assign n_1521 = ~n_1519 & ~n_1520;
assign n_1522 =  i_14 &  x_295;
assign n_1523 =  x_262 &  n_1522;
assign n_1524 =  i_13 &  x_295;
assign n_1525 = ~n_1524 & ~n_1522;
assign n_1526 =  x_225 &  n_1525;
assign n_1527 = ~x_2521 &  n_1526;
assign n_1528 = ~n_1523 & ~n_1527;
assign n_1529 =  x_262 & ~n_1528;
assign n_1530 = ~x_262 &  n_1528;
assign n_1531 = ~n_1529 & ~n_1530;
assign n_1532 =  x_261 &  n_1522;
assign n_1533 = ~x_2520 &  n_1526;
assign n_1534 = ~n_1532 & ~n_1533;
assign n_1535 =  x_261 & ~n_1534;
assign n_1536 = ~x_261 &  n_1534;
assign n_1537 = ~n_1535 & ~n_1536;
assign n_1538 =  x_260 &  n_1522;
assign n_1539 = ~x_2519 &  n_1526;
assign n_1540 = ~n_1538 & ~n_1539;
assign n_1541 =  x_260 & ~n_1540;
assign n_1542 = ~x_260 &  n_1540;
assign n_1543 = ~n_1541 & ~n_1542;
assign n_1544 =  x_259 &  n_1522;
assign n_1545 = ~x_2518 &  n_1526;
assign n_1546 = ~n_1544 & ~n_1545;
assign n_1547 =  x_259 & ~n_1546;
assign n_1548 = ~x_259 &  n_1546;
assign n_1549 = ~n_1547 & ~n_1548;
assign n_1550 =  x_258 &  n_1522;
assign n_1551 = ~x_2517 &  n_1526;
assign n_1552 = ~n_1550 & ~n_1551;
assign n_1553 =  x_258 & ~n_1552;
assign n_1554 = ~x_258 &  n_1552;
assign n_1555 = ~n_1553 & ~n_1554;
assign n_1556 =  x_257 &  n_1522;
assign n_1557 = ~x_2516 &  n_1526;
assign n_1558 = ~n_1556 & ~n_1557;
assign n_1559 =  x_257 & ~n_1558;
assign n_1560 = ~x_257 &  n_1558;
assign n_1561 = ~n_1559 & ~n_1560;
assign n_1562 =  x_256 &  n_1522;
assign n_1563 = ~x_2515 &  n_1526;
assign n_1564 = ~n_1562 & ~n_1563;
assign n_1565 =  x_256 & ~n_1564;
assign n_1566 = ~x_256 &  n_1564;
assign n_1567 = ~n_1565 & ~n_1566;
assign n_1568 =  x_255 &  n_1522;
assign n_1569 = ~x_2514 &  n_1526;
assign n_1570 = ~n_1568 & ~n_1569;
assign n_1571 =  x_255 & ~n_1570;
assign n_1572 = ~x_255 &  n_1570;
assign n_1573 = ~n_1571 & ~n_1572;
assign n_1574 =  x_254 &  n_1522;
assign n_1575 = ~x_2513 &  n_1526;
assign n_1576 = ~n_1574 & ~n_1575;
assign n_1577 =  x_254 & ~n_1576;
assign n_1578 = ~x_254 &  n_1576;
assign n_1579 = ~n_1577 & ~n_1578;
assign n_1580 =  x_253 &  n_1522;
assign n_1581 = ~x_2512 &  n_1526;
assign n_1582 = ~n_1580 & ~n_1581;
assign n_1583 =  x_253 & ~n_1582;
assign n_1584 = ~x_253 &  n_1582;
assign n_1585 = ~n_1583 & ~n_1584;
assign n_1586 =  x_252 &  n_1522;
assign n_1587 = ~x_2511 &  n_1526;
assign n_1588 = ~n_1586 & ~n_1587;
assign n_1589 =  x_252 & ~n_1588;
assign n_1590 = ~x_252 &  n_1588;
assign n_1591 = ~n_1589 & ~n_1590;
assign n_1592 =  x_251 &  n_1522;
assign n_1593 = ~x_2510 &  n_1526;
assign n_1594 = ~n_1592 & ~n_1593;
assign n_1595 =  x_251 & ~n_1594;
assign n_1596 = ~x_251 &  n_1594;
assign n_1597 = ~n_1595 & ~n_1596;
assign n_1598 =  x_250 &  n_1522;
assign n_1599 = ~x_2509 &  n_1526;
assign n_1600 = ~n_1598 & ~n_1599;
assign n_1601 =  x_250 & ~n_1600;
assign n_1602 = ~x_250 &  n_1600;
assign n_1603 = ~n_1601 & ~n_1602;
assign n_1604 =  x_249 &  n_1522;
assign n_1605 = ~x_2508 &  n_1526;
assign n_1606 = ~n_1604 & ~n_1605;
assign n_1607 =  x_249 & ~n_1606;
assign n_1608 = ~x_249 &  n_1606;
assign n_1609 = ~n_1607 & ~n_1608;
assign n_1610 =  x_248 &  n_1522;
assign n_1611 = ~x_2507 &  n_1526;
assign n_1612 = ~n_1610 & ~n_1611;
assign n_1613 =  x_248 & ~n_1612;
assign n_1614 = ~x_248 &  n_1612;
assign n_1615 = ~n_1613 & ~n_1614;
assign n_1616 =  x_247 &  n_1522;
assign n_1617 = ~x_2506 &  n_1526;
assign n_1618 = ~n_1616 & ~n_1617;
assign n_1619 =  x_247 & ~n_1618;
assign n_1620 = ~x_247 &  n_1618;
assign n_1621 = ~n_1619 & ~n_1620;
assign n_1622 =  x_246 &  n_1522;
assign n_1623 = ~x_2505 &  n_1526;
assign n_1624 = ~n_1622 & ~n_1623;
assign n_1625 =  x_246 & ~n_1624;
assign n_1626 = ~x_246 &  n_1624;
assign n_1627 = ~n_1625 & ~n_1626;
assign n_1628 =  x_245 &  n_1522;
assign n_1629 = ~x_2504 &  n_1526;
assign n_1630 = ~n_1628 & ~n_1629;
assign n_1631 =  x_245 & ~n_1630;
assign n_1632 = ~x_245 &  n_1630;
assign n_1633 = ~n_1631 & ~n_1632;
assign n_1634 =  x_244 &  n_1522;
assign n_1635 = ~x_2503 &  n_1526;
assign n_1636 = ~n_1634 & ~n_1635;
assign n_1637 =  x_244 & ~n_1636;
assign n_1638 = ~x_244 &  n_1636;
assign n_1639 = ~n_1637 & ~n_1638;
assign n_1640 =  x_243 &  n_1522;
assign n_1641 = ~x_2502 &  n_1526;
assign n_1642 = ~n_1640 & ~n_1641;
assign n_1643 =  x_243 & ~n_1642;
assign n_1644 = ~x_243 &  n_1642;
assign n_1645 = ~n_1643 & ~n_1644;
assign n_1646 =  x_242 &  n_1522;
assign n_1647 = ~x_2501 &  n_1526;
assign n_1648 = ~n_1646 & ~n_1647;
assign n_1649 =  x_242 & ~n_1648;
assign n_1650 = ~x_242 &  n_1648;
assign n_1651 = ~n_1649 & ~n_1650;
assign n_1652 =  x_241 &  n_1522;
assign n_1653 = ~x_2500 &  n_1526;
assign n_1654 = ~n_1652 & ~n_1653;
assign n_1655 =  x_241 & ~n_1654;
assign n_1656 = ~x_241 &  n_1654;
assign n_1657 = ~n_1655 & ~n_1656;
assign n_1658 =  x_240 &  n_1522;
assign n_1659 = ~x_2499 &  n_1526;
assign n_1660 = ~n_1658 & ~n_1659;
assign n_1661 =  x_240 & ~n_1660;
assign n_1662 = ~x_240 &  n_1660;
assign n_1663 = ~n_1661 & ~n_1662;
assign n_1664 =  x_239 &  n_1522;
assign n_1665 = ~x_2498 &  n_1526;
assign n_1666 = ~n_1664 & ~n_1665;
assign n_1667 =  x_239 & ~n_1666;
assign n_1668 = ~x_239 &  n_1666;
assign n_1669 = ~n_1667 & ~n_1668;
assign n_1670 =  x_238 &  n_1522;
assign n_1671 = ~x_2497 &  n_1526;
assign n_1672 = ~n_1670 & ~n_1671;
assign n_1673 =  x_238 & ~n_1672;
assign n_1674 = ~x_238 &  n_1672;
assign n_1675 = ~n_1673 & ~n_1674;
assign n_1676 =  x_237 &  n_1522;
assign n_1677 = ~x_2496 &  n_1526;
assign n_1678 = ~n_1676 & ~n_1677;
assign n_1679 =  x_237 & ~n_1678;
assign n_1680 = ~x_237 &  n_1678;
assign n_1681 = ~n_1679 & ~n_1680;
assign n_1682 =  x_236 &  n_1522;
assign n_1683 = ~x_2495 &  n_1526;
assign n_1684 = ~n_1682 & ~n_1683;
assign n_1685 =  x_236 & ~n_1684;
assign n_1686 = ~x_236 &  n_1684;
assign n_1687 = ~n_1685 & ~n_1686;
assign n_1688 =  x_235 &  n_1522;
assign n_1689 = ~x_2494 &  n_1526;
assign n_1690 = ~n_1688 & ~n_1689;
assign n_1691 =  x_235 & ~n_1690;
assign n_1692 = ~x_235 &  n_1690;
assign n_1693 = ~n_1691 & ~n_1692;
assign n_1694 =  x_234 &  n_1522;
assign n_1695 = ~x_2493 &  n_1526;
assign n_1696 = ~n_1694 & ~n_1695;
assign n_1697 =  x_234 & ~n_1696;
assign n_1698 = ~x_234 &  n_1696;
assign n_1699 = ~n_1697 & ~n_1698;
assign n_1700 =  x_233 &  n_1522;
assign n_1701 =  x_2492 &  n_1526;
assign n_1702 = ~n_1700 & ~n_1701;
assign n_1703 =  x_233 & ~n_1702;
assign n_1704 = ~x_233 &  n_1702;
assign n_1705 = ~n_1703 & ~n_1704;
assign n_1706 =  x_232 & ~n_1522;
assign n_1707 = ~x_232 & ~n_1525;
assign n_1708 = ~n_1706 & ~n_1707;
assign n_1709 =  x_232 &  n_1708;
assign n_1710 = ~x_232 & ~n_1708;
assign n_1711 = ~n_1709 & ~n_1710;
assign n_1712 = ~n_509 &  n_1211;
assign n_1713 = ~n_1321 &  n_1220;
assign n_1714 =  n_1712 &  n_1713;
assign n_1715 =  n_475 &  n_1714;
assign n_1716 = ~x_229 &  n_1715;
assign n_1717 =  n_1321 & ~n_1219;
assign n_1718 = ~n_1716 & ~n_1717;
assign n_1719 = ~n_1718 &  n_1195;
assign n_1720 =  x_231 &  n_1719;
assign n_1721 = ~x_231 & ~n_1719;
assign n_1722 = ~n_1720 & ~n_1721;
assign n_1723 =  x_1470 &  n_1716;
assign n_1724 = ~n_1262 &  n_1723;
assign n_1725 =  x_230 & ~n_1724;
assign n_1726 = ~x_230 &  n_1724;
assign n_1727 = ~n_1725 & ~n_1726;
assign n_1728 =  x_229 &  n_1724;
assign n_1729 = ~x_229 & ~n_1724;
assign n_1730 = ~n_1728 & ~n_1729;
assign n_1731 = ~x_227 &  n_1325;
assign n_1732 = ~n_1328 & ~n_1731;
assign n_1733 =  x_228 & ~n_1732;
assign n_1734 = ~x_228 &  n_1732;
assign n_1735 = ~n_1733 & ~n_1734;
assign n_1736 =  x_227 &  n_1732;
assign n_1737 = ~x_227 & ~n_1732;
assign n_1738 = ~n_1736 & ~n_1737;
assign n_1739 =  n_1524 & ~n_1522;
assign n_1740 = ~x_225 &  n_1522;
assign n_1741 = ~n_1739 & ~n_1740;
assign n_1742 =  x_226 & ~n_1741;
assign n_1743 = ~x_226 &  n_1741;
assign n_1744 = ~n_1742 & ~n_1743;
assign n_1745 =  x_225 &  n_1741;
assign n_1746 = ~x_225 & ~n_1741;
assign n_1747 = ~n_1745 & ~n_1746;
assign n_1748 =  x_1492 &  x_1771;
assign n_1749 =  x_1493 &  n_1748;
assign n_1750 =  x_1494 &  n_1749;
assign n_1751 =  x_310 &  x_1768;
assign n_1752 =  i_191 &  n_1751;
assign n_1753 =  n_1750 & ~n_1752;
assign n_1754 = ~x_2158 & ~n_1750;
assign n_1755 = ~n_1753 & ~n_1754;
assign n_1756 =  x_2158 &  n_1755;
assign n_1757 = ~x_2158 & ~n_1755;
assign n_1758 = ~n_1756 & ~n_1757;
assign n_1759 = ~x_1492 &  x_1771;
assign n_1760 = ~x_1493 &  n_1759;
assign n_1761 = ~x_1494 &  n_1760;
assign n_1762 =  x_2157 & ~n_1761;
assign n_1763 =  i_190 &  n_1751;
assign n_1764 =  n_1761 &  n_1763;
assign n_1765 = ~n_1762 & ~n_1764;
assign n_1766 =  x_2157 & ~n_1765;
assign n_1767 = ~x_2157 &  n_1765;
assign n_1768 = ~n_1766 & ~n_1767;
assign n_1769 = ~x_1493 &  n_1748;
assign n_1770 = ~x_1494 &  n_1769;
assign n_1771 =  x_2156 & ~n_1770;
assign n_1772 =  n_1770 &  n_1763;
assign n_1773 = ~n_1771 & ~n_1772;
assign n_1774 =  x_2156 & ~n_1773;
assign n_1775 = ~x_2156 &  n_1773;
assign n_1776 = ~n_1774 & ~n_1775;
assign n_1777 =  x_1493 &  n_1759;
assign n_1778 = ~x_1494 &  n_1777;
assign n_1779 =  x_2155 & ~n_1778;
assign n_1780 =  n_1778 &  n_1763;
assign n_1781 = ~n_1779 & ~n_1780;
assign n_1782 =  x_2155 & ~n_1781;
assign n_1783 = ~x_2155 &  n_1781;
assign n_1784 = ~n_1782 & ~n_1783;
assign n_1785 = ~x_1494 &  n_1749;
assign n_1786 =  x_2154 & ~n_1785;
assign n_1787 =  n_1785 &  n_1763;
assign n_1788 = ~n_1786 & ~n_1787;
assign n_1789 =  x_2154 & ~n_1788;
assign n_1790 = ~x_2154 &  n_1788;
assign n_1791 = ~n_1789 & ~n_1790;
assign n_1792 =  x_1494 &  n_1760;
assign n_1793 =  x_2153 & ~n_1792;
assign n_1794 =  n_1792 &  n_1763;
assign n_1795 = ~n_1793 & ~n_1794;
assign n_1796 =  x_2153 & ~n_1795;
assign n_1797 = ~x_2153 &  n_1795;
assign n_1798 = ~n_1796 & ~n_1797;
assign n_1799 =  x_1494 &  n_1769;
assign n_1800 =  x_2152 & ~n_1799;
assign n_1801 =  n_1799 &  n_1763;
assign n_1802 = ~n_1800 & ~n_1801;
assign n_1803 =  x_2152 & ~n_1802;
assign n_1804 = ~x_2152 &  n_1802;
assign n_1805 = ~n_1803 & ~n_1804;
assign n_1806 =  x_1494 &  n_1777;
assign n_1807 =  x_2151 & ~n_1806;
assign n_1808 =  n_1806 &  n_1763;
assign n_1809 = ~n_1807 & ~n_1808;
assign n_1810 =  x_2151 & ~n_1809;
assign n_1811 = ~x_2151 &  n_1809;
assign n_1812 = ~n_1810 & ~n_1811;
assign n_1813 =  n_1750 & ~n_1763;
assign n_1814 = ~x_2150 & ~n_1750;
assign n_1815 = ~n_1813 & ~n_1814;
assign n_1816 =  x_2150 &  n_1815;
assign n_1817 = ~x_2150 & ~n_1815;
assign n_1818 = ~n_1816 & ~n_1817;
assign n_1819 =  x_2149 & ~n_1761;
assign n_1820 =  i_189 &  n_1751;
assign n_1821 =  n_1761 &  n_1820;
assign n_1822 = ~n_1819 & ~n_1821;
assign n_1823 =  x_2149 & ~n_1822;
assign n_1824 = ~x_2149 &  n_1822;
assign n_1825 = ~n_1823 & ~n_1824;
assign n_1826 =  x_2148 & ~n_1770;
assign n_1827 =  n_1770 &  n_1820;
assign n_1828 = ~n_1826 & ~n_1827;
assign n_1829 =  x_2148 & ~n_1828;
assign n_1830 = ~x_2148 &  n_1828;
assign n_1831 = ~n_1829 & ~n_1830;
assign n_1832 =  x_2147 & ~n_1778;
assign n_1833 =  n_1778 &  n_1820;
assign n_1834 = ~n_1832 & ~n_1833;
assign n_1835 =  x_2147 & ~n_1834;
assign n_1836 = ~x_2147 &  n_1834;
assign n_1837 = ~n_1835 & ~n_1836;
assign n_1838 =  x_2146 & ~n_1785;
assign n_1839 =  n_1785 &  n_1820;
assign n_1840 = ~n_1838 & ~n_1839;
assign n_1841 =  x_2146 & ~n_1840;
assign n_1842 = ~x_2146 &  n_1840;
assign n_1843 = ~n_1841 & ~n_1842;
assign n_1844 =  x_2145 & ~n_1792;
assign n_1845 =  n_1792 &  n_1820;
assign n_1846 = ~n_1844 & ~n_1845;
assign n_1847 =  x_2145 & ~n_1846;
assign n_1848 = ~x_2145 &  n_1846;
assign n_1849 = ~n_1847 & ~n_1848;
assign n_1850 =  x_2144 & ~n_1799;
assign n_1851 =  n_1799 &  n_1820;
assign n_1852 = ~n_1850 & ~n_1851;
assign n_1853 =  x_2144 & ~n_1852;
assign n_1854 = ~x_2144 &  n_1852;
assign n_1855 = ~n_1853 & ~n_1854;
assign n_1856 =  x_2143 & ~n_1806;
assign n_1857 =  n_1806 &  n_1820;
assign n_1858 = ~n_1856 & ~n_1857;
assign n_1859 =  x_2143 & ~n_1858;
assign n_1860 = ~x_2143 &  n_1858;
assign n_1861 = ~n_1859 & ~n_1860;
assign n_1862 =  n_1750 & ~n_1820;
assign n_1863 = ~x_2142 & ~n_1750;
assign n_1864 = ~n_1862 & ~n_1863;
assign n_1865 =  x_2142 &  n_1864;
assign n_1866 = ~x_2142 & ~n_1864;
assign n_1867 = ~n_1865 & ~n_1866;
assign n_1868 =  x_2141 & ~n_1761;
assign n_1869 =  i_188 &  n_1751;
assign n_1870 =  n_1761 &  n_1869;
assign n_1871 = ~n_1868 & ~n_1870;
assign n_1872 =  x_2141 & ~n_1871;
assign n_1873 = ~x_2141 &  n_1871;
assign n_1874 = ~n_1872 & ~n_1873;
assign n_1875 =  x_2140 & ~n_1770;
assign n_1876 =  n_1770 &  n_1869;
assign n_1877 = ~n_1875 & ~n_1876;
assign n_1878 =  x_2140 & ~n_1877;
assign n_1879 = ~x_2140 &  n_1877;
assign n_1880 = ~n_1878 & ~n_1879;
assign n_1881 =  x_2139 & ~n_1778;
assign n_1882 =  n_1778 &  n_1869;
assign n_1883 = ~n_1881 & ~n_1882;
assign n_1884 =  x_2139 & ~n_1883;
assign n_1885 = ~x_2139 &  n_1883;
assign n_1886 = ~n_1884 & ~n_1885;
assign n_1887 =  x_2138 & ~n_1785;
assign n_1888 =  n_1785 &  n_1869;
assign n_1889 = ~n_1887 & ~n_1888;
assign n_1890 =  x_2138 & ~n_1889;
assign n_1891 = ~x_2138 &  n_1889;
assign n_1892 = ~n_1890 & ~n_1891;
assign n_1893 =  x_2137 & ~n_1792;
assign n_1894 =  n_1792 &  n_1869;
assign n_1895 = ~n_1893 & ~n_1894;
assign n_1896 =  x_2137 & ~n_1895;
assign n_1897 = ~x_2137 &  n_1895;
assign n_1898 = ~n_1896 & ~n_1897;
assign n_1899 =  x_2136 & ~n_1799;
assign n_1900 =  n_1799 &  n_1869;
assign n_1901 = ~n_1899 & ~n_1900;
assign n_1902 =  x_2136 & ~n_1901;
assign n_1903 = ~x_2136 &  n_1901;
assign n_1904 = ~n_1902 & ~n_1903;
assign n_1905 =  x_2135 & ~n_1806;
assign n_1906 =  n_1806 &  n_1869;
assign n_1907 = ~n_1905 & ~n_1906;
assign n_1908 =  x_2135 & ~n_1907;
assign n_1909 = ~x_2135 &  n_1907;
assign n_1910 = ~n_1908 & ~n_1909;
assign n_1911 =  n_1750 & ~n_1869;
assign n_1912 = ~x_2134 & ~n_1750;
assign n_1913 = ~n_1911 & ~n_1912;
assign n_1914 =  x_2134 &  n_1913;
assign n_1915 = ~x_2134 & ~n_1913;
assign n_1916 = ~n_1914 & ~n_1915;
assign n_1917 =  x_2133 & ~n_1761;
assign n_1918 =  i_187 &  n_1751;
assign n_1919 =  n_1761 &  n_1918;
assign n_1920 = ~n_1917 & ~n_1919;
assign n_1921 =  x_2133 & ~n_1920;
assign n_1922 = ~x_2133 &  n_1920;
assign n_1923 = ~n_1921 & ~n_1922;
assign n_1924 =  x_2132 & ~n_1770;
assign n_1925 =  n_1770 &  n_1918;
assign n_1926 = ~n_1924 & ~n_1925;
assign n_1927 =  x_2132 & ~n_1926;
assign n_1928 = ~x_2132 &  n_1926;
assign n_1929 = ~n_1927 & ~n_1928;
assign n_1930 =  x_2131 & ~n_1778;
assign n_1931 =  n_1778 &  n_1918;
assign n_1932 = ~n_1930 & ~n_1931;
assign n_1933 =  x_2131 & ~n_1932;
assign n_1934 = ~x_2131 &  n_1932;
assign n_1935 = ~n_1933 & ~n_1934;
assign n_1936 =  x_2130 & ~n_1785;
assign n_1937 =  n_1785 &  n_1918;
assign n_1938 = ~n_1936 & ~n_1937;
assign n_1939 =  x_2130 & ~n_1938;
assign n_1940 = ~x_2130 &  n_1938;
assign n_1941 = ~n_1939 & ~n_1940;
assign n_1942 =  x_2129 & ~n_1792;
assign n_1943 =  n_1792 &  n_1918;
assign n_1944 = ~n_1942 & ~n_1943;
assign n_1945 =  x_2129 & ~n_1944;
assign n_1946 = ~x_2129 &  n_1944;
assign n_1947 = ~n_1945 & ~n_1946;
assign n_1948 =  x_2128 & ~n_1799;
assign n_1949 =  n_1799 &  n_1918;
assign n_1950 = ~n_1948 & ~n_1949;
assign n_1951 =  x_2128 & ~n_1950;
assign n_1952 = ~x_2128 &  n_1950;
assign n_1953 = ~n_1951 & ~n_1952;
assign n_1954 =  x_2127 & ~n_1806;
assign n_1955 =  n_1806 &  n_1918;
assign n_1956 = ~n_1954 & ~n_1955;
assign n_1957 =  x_2127 & ~n_1956;
assign n_1958 = ~x_2127 &  n_1956;
assign n_1959 = ~n_1957 & ~n_1958;
assign n_1960 =  n_1750 & ~n_1918;
assign n_1961 = ~x_2126 & ~n_1750;
assign n_1962 = ~n_1960 & ~n_1961;
assign n_1963 =  x_2126 &  n_1962;
assign n_1964 = ~x_2126 & ~n_1962;
assign n_1965 = ~n_1963 & ~n_1964;
assign n_1966 =  x_2125 & ~n_1761;
assign n_1967 =  i_186 &  n_1751;
assign n_1968 =  n_1761 &  n_1967;
assign n_1969 = ~n_1966 & ~n_1968;
assign n_1970 =  x_2125 & ~n_1969;
assign n_1971 = ~x_2125 &  n_1969;
assign n_1972 = ~n_1970 & ~n_1971;
assign n_1973 =  x_2124 & ~n_1770;
assign n_1974 =  n_1770 &  n_1967;
assign n_1975 = ~n_1973 & ~n_1974;
assign n_1976 =  x_2124 & ~n_1975;
assign n_1977 = ~x_2124 &  n_1975;
assign n_1978 = ~n_1976 & ~n_1977;
assign n_1979 =  x_2123 & ~n_1778;
assign n_1980 =  n_1778 &  n_1967;
assign n_1981 = ~n_1979 & ~n_1980;
assign n_1982 =  x_2123 & ~n_1981;
assign n_1983 = ~x_2123 &  n_1981;
assign n_1984 = ~n_1982 & ~n_1983;
assign n_1985 =  x_2122 & ~n_1785;
assign n_1986 =  n_1785 &  n_1967;
assign n_1987 = ~n_1985 & ~n_1986;
assign n_1988 =  x_2122 & ~n_1987;
assign n_1989 = ~x_2122 &  n_1987;
assign n_1990 = ~n_1988 & ~n_1989;
assign n_1991 =  x_2121 & ~n_1792;
assign n_1992 =  n_1792 &  n_1967;
assign n_1993 = ~n_1991 & ~n_1992;
assign n_1994 =  x_2121 & ~n_1993;
assign n_1995 = ~x_2121 &  n_1993;
assign n_1996 = ~n_1994 & ~n_1995;
assign n_1997 =  x_2120 & ~n_1799;
assign n_1998 =  n_1799 &  n_1967;
assign n_1999 = ~n_1997 & ~n_1998;
assign n_2000 =  x_2120 & ~n_1999;
assign n_2001 = ~x_2120 &  n_1999;
assign n_2002 = ~n_2000 & ~n_2001;
assign n_2003 =  x_2119 & ~n_1806;
assign n_2004 =  n_1806 &  n_1967;
assign n_2005 = ~n_2003 & ~n_2004;
assign n_2006 =  x_2119 & ~n_2005;
assign n_2007 = ~x_2119 &  n_2005;
assign n_2008 = ~n_2006 & ~n_2007;
assign n_2009 =  n_1750 & ~n_1967;
assign n_2010 = ~x_2118 & ~n_1750;
assign n_2011 = ~n_2009 & ~n_2010;
assign n_2012 =  x_2118 &  n_2011;
assign n_2013 = ~x_2118 & ~n_2011;
assign n_2014 = ~n_2012 & ~n_2013;
assign n_2015 =  x_2117 & ~n_1761;
assign n_2016 =  i_185 &  n_1751;
assign n_2017 =  n_1761 &  n_2016;
assign n_2018 = ~n_2015 & ~n_2017;
assign n_2019 =  x_2117 & ~n_2018;
assign n_2020 = ~x_2117 &  n_2018;
assign n_2021 = ~n_2019 & ~n_2020;
assign n_2022 =  x_2116 & ~n_1770;
assign n_2023 =  n_1770 &  n_2016;
assign n_2024 = ~n_2022 & ~n_2023;
assign n_2025 =  x_2116 & ~n_2024;
assign n_2026 = ~x_2116 &  n_2024;
assign n_2027 = ~n_2025 & ~n_2026;
assign n_2028 =  x_2115 & ~n_1778;
assign n_2029 =  n_1778 &  n_2016;
assign n_2030 = ~n_2028 & ~n_2029;
assign n_2031 =  x_2115 & ~n_2030;
assign n_2032 = ~x_2115 &  n_2030;
assign n_2033 = ~n_2031 & ~n_2032;
assign n_2034 =  x_2114 & ~n_1785;
assign n_2035 =  n_1785 &  n_2016;
assign n_2036 = ~n_2034 & ~n_2035;
assign n_2037 =  x_2114 & ~n_2036;
assign n_2038 = ~x_2114 &  n_2036;
assign n_2039 = ~n_2037 & ~n_2038;
assign n_2040 =  x_2113 & ~n_1792;
assign n_2041 =  n_1792 &  n_2016;
assign n_2042 = ~n_2040 & ~n_2041;
assign n_2043 =  x_2113 & ~n_2042;
assign n_2044 = ~x_2113 &  n_2042;
assign n_2045 = ~n_2043 & ~n_2044;
assign n_2046 =  x_2112 & ~n_1799;
assign n_2047 =  n_1799 &  n_2016;
assign n_2048 = ~n_2046 & ~n_2047;
assign n_2049 =  x_2112 & ~n_2048;
assign n_2050 = ~x_2112 &  n_2048;
assign n_2051 = ~n_2049 & ~n_2050;
assign n_2052 =  x_2111 & ~n_1806;
assign n_2053 =  n_1806 &  n_2016;
assign n_2054 = ~n_2052 & ~n_2053;
assign n_2055 =  x_2111 & ~n_2054;
assign n_2056 = ~x_2111 &  n_2054;
assign n_2057 = ~n_2055 & ~n_2056;
assign n_2058 =  n_1750 & ~n_2016;
assign n_2059 = ~x_2110 & ~n_1750;
assign n_2060 = ~n_2058 & ~n_2059;
assign n_2061 =  x_2110 &  n_2060;
assign n_2062 = ~x_2110 & ~n_2060;
assign n_2063 = ~n_2061 & ~n_2062;
assign n_2064 =  x_2109 & ~n_1761;
assign n_2065 =  i_184 &  n_1751;
assign n_2066 =  n_1761 &  n_2065;
assign n_2067 = ~n_2064 & ~n_2066;
assign n_2068 =  x_2109 & ~n_2067;
assign n_2069 = ~x_2109 &  n_2067;
assign n_2070 = ~n_2068 & ~n_2069;
assign n_2071 =  x_2108 & ~n_1770;
assign n_2072 =  n_1770 &  n_2065;
assign n_2073 = ~n_2071 & ~n_2072;
assign n_2074 =  x_2108 & ~n_2073;
assign n_2075 = ~x_2108 &  n_2073;
assign n_2076 = ~n_2074 & ~n_2075;
assign n_2077 =  x_2107 & ~n_1778;
assign n_2078 =  n_1778 &  n_2065;
assign n_2079 = ~n_2077 & ~n_2078;
assign n_2080 =  x_2107 & ~n_2079;
assign n_2081 = ~x_2107 &  n_2079;
assign n_2082 = ~n_2080 & ~n_2081;
assign n_2083 =  x_2106 & ~n_1785;
assign n_2084 =  n_1785 &  n_2065;
assign n_2085 = ~n_2083 & ~n_2084;
assign n_2086 =  x_2106 & ~n_2085;
assign n_2087 = ~x_2106 &  n_2085;
assign n_2088 = ~n_2086 & ~n_2087;
assign n_2089 =  x_2105 & ~n_1792;
assign n_2090 =  n_1792 &  n_2065;
assign n_2091 = ~n_2089 & ~n_2090;
assign n_2092 =  x_2105 & ~n_2091;
assign n_2093 = ~x_2105 &  n_2091;
assign n_2094 = ~n_2092 & ~n_2093;
assign n_2095 =  x_2104 & ~n_1799;
assign n_2096 =  n_1799 &  n_2065;
assign n_2097 = ~n_2095 & ~n_2096;
assign n_2098 =  x_2104 & ~n_2097;
assign n_2099 = ~x_2104 &  n_2097;
assign n_2100 = ~n_2098 & ~n_2099;
assign n_2101 =  x_2103 & ~n_1806;
assign n_2102 =  n_1806 &  n_2065;
assign n_2103 = ~n_2101 & ~n_2102;
assign n_2104 =  x_2103 & ~n_2103;
assign n_2105 = ~x_2103 &  n_2103;
assign n_2106 = ~n_2104 & ~n_2105;
assign n_2107 =  n_1750 & ~n_2065;
assign n_2108 = ~x_2102 & ~n_1750;
assign n_2109 = ~n_2107 & ~n_2108;
assign n_2110 =  x_2102 &  n_2109;
assign n_2111 = ~x_2102 & ~n_2109;
assign n_2112 = ~n_2110 & ~n_2111;
assign n_2113 =  x_2101 & ~n_1761;
assign n_2114 =  i_183 &  n_1751;
assign n_2115 =  n_1761 &  n_2114;
assign n_2116 = ~n_2113 & ~n_2115;
assign n_2117 =  x_2101 & ~n_2116;
assign n_2118 = ~x_2101 &  n_2116;
assign n_2119 = ~n_2117 & ~n_2118;
assign n_2120 =  x_2100 & ~n_1770;
assign n_2121 =  n_1770 &  n_2114;
assign n_2122 = ~n_2120 & ~n_2121;
assign n_2123 =  x_2100 & ~n_2122;
assign n_2124 = ~x_2100 &  n_2122;
assign n_2125 = ~n_2123 & ~n_2124;
assign n_2126 =  x_2099 & ~n_1778;
assign n_2127 =  n_1778 &  n_2114;
assign n_2128 = ~n_2126 & ~n_2127;
assign n_2129 =  x_2099 & ~n_2128;
assign n_2130 = ~x_2099 &  n_2128;
assign n_2131 = ~n_2129 & ~n_2130;
assign n_2132 =  x_2098 & ~n_1785;
assign n_2133 =  n_1785 &  n_2114;
assign n_2134 = ~n_2132 & ~n_2133;
assign n_2135 =  x_2098 & ~n_2134;
assign n_2136 = ~x_2098 &  n_2134;
assign n_2137 = ~n_2135 & ~n_2136;
assign n_2138 =  x_2097 & ~n_1792;
assign n_2139 =  n_1792 &  n_2114;
assign n_2140 = ~n_2138 & ~n_2139;
assign n_2141 =  x_2097 & ~n_2140;
assign n_2142 = ~x_2097 &  n_2140;
assign n_2143 = ~n_2141 & ~n_2142;
assign n_2144 =  x_2096 & ~n_1799;
assign n_2145 =  n_1799 &  n_2114;
assign n_2146 = ~n_2144 & ~n_2145;
assign n_2147 =  x_2096 & ~n_2146;
assign n_2148 = ~x_2096 &  n_2146;
assign n_2149 = ~n_2147 & ~n_2148;
assign n_2150 =  x_2095 & ~n_1806;
assign n_2151 =  n_1806 &  n_2114;
assign n_2152 = ~n_2150 & ~n_2151;
assign n_2153 =  x_2095 & ~n_2152;
assign n_2154 = ~x_2095 &  n_2152;
assign n_2155 = ~n_2153 & ~n_2154;
assign n_2156 =  n_1750 & ~n_2114;
assign n_2157 = ~x_2094 & ~n_1750;
assign n_2158 = ~n_2156 & ~n_2157;
assign n_2159 =  x_2094 &  n_2158;
assign n_2160 = ~x_2094 & ~n_2158;
assign n_2161 = ~n_2159 & ~n_2160;
assign n_2162 =  x_2093 & ~n_1761;
assign n_2163 =  i_182 &  n_1751;
assign n_2164 =  n_1761 &  n_2163;
assign n_2165 = ~n_2162 & ~n_2164;
assign n_2166 =  x_2093 & ~n_2165;
assign n_2167 = ~x_2093 &  n_2165;
assign n_2168 = ~n_2166 & ~n_2167;
assign n_2169 =  x_2092 & ~n_1770;
assign n_2170 =  n_1770 &  n_2163;
assign n_2171 = ~n_2169 & ~n_2170;
assign n_2172 =  x_2092 & ~n_2171;
assign n_2173 = ~x_2092 &  n_2171;
assign n_2174 = ~n_2172 & ~n_2173;
assign n_2175 =  x_2091 & ~n_1778;
assign n_2176 =  n_1778 &  n_2163;
assign n_2177 = ~n_2175 & ~n_2176;
assign n_2178 =  x_2091 & ~n_2177;
assign n_2179 = ~x_2091 &  n_2177;
assign n_2180 = ~n_2178 & ~n_2179;
assign n_2181 =  x_2090 & ~n_1785;
assign n_2182 =  n_1785 &  n_2163;
assign n_2183 = ~n_2181 & ~n_2182;
assign n_2184 =  x_2090 & ~n_2183;
assign n_2185 = ~x_2090 &  n_2183;
assign n_2186 = ~n_2184 & ~n_2185;
assign n_2187 =  x_2089 & ~n_1792;
assign n_2188 =  n_1792 &  n_2163;
assign n_2189 = ~n_2187 & ~n_2188;
assign n_2190 =  x_2089 & ~n_2189;
assign n_2191 = ~x_2089 &  n_2189;
assign n_2192 = ~n_2190 & ~n_2191;
assign n_2193 =  x_2088 & ~n_1799;
assign n_2194 =  n_1799 &  n_2163;
assign n_2195 = ~n_2193 & ~n_2194;
assign n_2196 =  x_2088 & ~n_2195;
assign n_2197 = ~x_2088 &  n_2195;
assign n_2198 = ~n_2196 & ~n_2197;
assign n_2199 =  x_2087 & ~n_1806;
assign n_2200 =  n_1806 &  n_2163;
assign n_2201 = ~n_2199 & ~n_2200;
assign n_2202 =  x_2087 & ~n_2201;
assign n_2203 = ~x_2087 &  n_2201;
assign n_2204 = ~n_2202 & ~n_2203;
assign n_2205 =  n_1750 & ~n_2163;
assign n_2206 = ~x_2086 & ~n_1750;
assign n_2207 = ~n_2205 & ~n_2206;
assign n_2208 =  x_2086 &  n_2207;
assign n_2209 = ~x_2086 & ~n_2207;
assign n_2210 = ~n_2208 & ~n_2209;
assign n_2211 =  x_2085 & ~n_1761;
assign n_2212 =  i_181 &  n_1751;
assign n_2213 =  n_1761 &  n_2212;
assign n_2214 = ~n_2211 & ~n_2213;
assign n_2215 =  x_2085 & ~n_2214;
assign n_2216 = ~x_2085 &  n_2214;
assign n_2217 = ~n_2215 & ~n_2216;
assign n_2218 =  x_2084 & ~n_1770;
assign n_2219 =  n_1770 &  n_2212;
assign n_2220 = ~n_2218 & ~n_2219;
assign n_2221 =  x_2084 & ~n_2220;
assign n_2222 = ~x_2084 &  n_2220;
assign n_2223 = ~n_2221 & ~n_2222;
assign n_2224 =  x_2083 & ~n_1778;
assign n_2225 =  n_1778 &  n_2212;
assign n_2226 = ~n_2224 & ~n_2225;
assign n_2227 =  x_2083 & ~n_2226;
assign n_2228 = ~x_2083 &  n_2226;
assign n_2229 = ~n_2227 & ~n_2228;
assign n_2230 =  x_2082 & ~n_1785;
assign n_2231 =  n_1785 &  n_2212;
assign n_2232 = ~n_2230 & ~n_2231;
assign n_2233 =  x_2082 & ~n_2232;
assign n_2234 = ~x_2082 &  n_2232;
assign n_2235 = ~n_2233 & ~n_2234;
assign n_2236 =  x_2081 & ~n_1792;
assign n_2237 =  n_1792 &  n_2212;
assign n_2238 = ~n_2236 & ~n_2237;
assign n_2239 =  x_2081 & ~n_2238;
assign n_2240 = ~x_2081 &  n_2238;
assign n_2241 = ~n_2239 & ~n_2240;
assign n_2242 =  x_2080 & ~n_1799;
assign n_2243 =  n_1799 &  n_2212;
assign n_2244 = ~n_2242 & ~n_2243;
assign n_2245 =  x_2080 & ~n_2244;
assign n_2246 = ~x_2080 &  n_2244;
assign n_2247 = ~n_2245 & ~n_2246;
assign n_2248 =  x_2079 & ~n_1806;
assign n_2249 =  n_1806 &  n_2212;
assign n_2250 = ~n_2248 & ~n_2249;
assign n_2251 =  x_2079 & ~n_2250;
assign n_2252 = ~x_2079 &  n_2250;
assign n_2253 = ~n_2251 & ~n_2252;
assign n_2254 =  n_1750 & ~n_2212;
assign n_2255 = ~x_2078 & ~n_1750;
assign n_2256 = ~n_2254 & ~n_2255;
assign n_2257 =  x_2078 &  n_2256;
assign n_2258 = ~x_2078 & ~n_2256;
assign n_2259 = ~n_2257 & ~n_2258;
assign n_2260 =  x_2077 & ~n_1761;
assign n_2261 =  i_180 &  n_1751;
assign n_2262 =  n_1761 &  n_2261;
assign n_2263 = ~n_2260 & ~n_2262;
assign n_2264 =  x_2077 & ~n_2263;
assign n_2265 = ~x_2077 &  n_2263;
assign n_2266 = ~n_2264 & ~n_2265;
assign n_2267 =  x_2076 & ~n_1770;
assign n_2268 =  n_1770 &  n_2261;
assign n_2269 = ~n_2267 & ~n_2268;
assign n_2270 =  x_2076 & ~n_2269;
assign n_2271 = ~x_2076 &  n_2269;
assign n_2272 = ~n_2270 & ~n_2271;
assign n_2273 =  x_2075 & ~n_1778;
assign n_2274 =  n_1778 &  n_2261;
assign n_2275 = ~n_2273 & ~n_2274;
assign n_2276 =  x_2075 & ~n_2275;
assign n_2277 = ~x_2075 &  n_2275;
assign n_2278 = ~n_2276 & ~n_2277;
assign n_2279 =  x_2074 & ~n_1785;
assign n_2280 =  n_1785 &  n_2261;
assign n_2281 = ~n_2279 & ~n_2280;
assign n_2282 =  x_2074 & ~n_2281;
assign n_2283 = ~x_2074 &  n_2281;
assign n_2284 = ~n_2282 & ~n_2283;
assign n_2285 =  x_2073 & ~n_1792;
assign n_2286 =  n_1792 &  n_2261;
assign n_2287 = ~n_2285 & ~n_2286;
assign n_2288 =  x_2073 & ~n_2287;
assign n_2289 = ~x_2073 &  n_2287;
assign n_2290 = ~n_2288 & ~n_2289;
assign n_2291 =  x_2072 & ~n_1799;
assign n_2292 =  n_1799 &  n_2261;
assign n_2293 = ~n_2291 & ~n_2292;
assign n_2294 =  x_2072 & ~n_2293;
assign n_2295 = ~x_2072 &  n_2293;
assign n_2296 = ~n_2294 & ~n_2295;
assign n_2297 =  x_2071 & ~n_1806;
assign n_2298 =  n_1806 &  n_2261;
assign n_2299 = ~n_2297 & ~n_2298;
assign n_2300 =  x_2071 & ~n_2299;
assign n_2301 = ~x_2071 &  n_2299;
assign n_2302 = ~n_2300 & ~n_2301;
assign n_2303 =  n_1750 & ~n_2261;
assign n_2304 = ~x_2070 & ~n_1750;
assign n_2305 = ~n_2303 & ~n_2304;
assign n_2306 =  x_2070 &  n_2305;
assign n_2307 = ~x_2070 & ~n_2305;
assign n_2308 = ~n_2306 & ~n_2307;
assign n_2309 =  x_2069 & ~n_1761;
assign n_2310 =  i_179 &  n_1751;
assign n_2311 =  n_1761 &  n_2310;
assign n_2312 = ~n_2309 & ~n_2311;
assign n_2313 =  x_2069 & ~n_2312;
assign n_2314 = ~x_2069 &  n_2312;
assign n_2315 = ~n_2313 & ~n_2314;
assign n_2316 =  x_2068 & ~n_1770;
assign n_2317 =  n_1770 &  n_2310;
assign n_2318 = ~n_2316 & ~n_2317;
assign n_2319 =  x_2068 & ~n_2318;
assign n_2320 = ~x_2068 &  n_2318;
assign n_2321 = ~n_2319 & ~n_2320;
assign n_2322 =  x_2067 & ~n_1778;
assign n_2323 =  n_1778 &  n_2310;
assign n_2324 = ~n_2322 & ~n_2323;
assign n_2325 =  x_2067 & ~n_2324;
assign n_2326 = ~x_2067 &  n_2324;
assign n_2327 = ~n_2325 & ~n_2326;
assign n_2328 =  x_2066 & ~n_1785;
assign n_2329 =  n_1785 &  n_2310;
assign n_2330 = ~n_2328 & ~n_2329;
assign n_2331 =  x_2066 & ~n_2330;
assign n_2332 = ~x_2066 &  n_2330;
assign n_2333 = ~n_2331 & ~n_2332;
assign n_2334 =  x_2065 & ~n_1792;
assign n_2335 =  n_1792 &  n_2310;
assign n_2336 = ~n_2334 & ~n_2335;
assign n_2337 =  x_2065 & ~n_2336;
assign n_2338 = ~x_2065 &  n_2336;
assign n_2339 = ~n_2337 & ~n_2338;
assign n_2340 =  x_2064 & ~n_1799;
assign n_2341 =  n_1799 &  n_2310;
assign n_2342 = ~n_2340 & ~n_2341;
assign n_2343 =  x_2064 & ~n_2342;
assign n_2344 = ~x_2064 &  n_2342;
assign n_2345 = ~n_2343 & ~n_2344;
assign n_2346 =  x_2063 & ~n_1806;
assign n_2347 =  n_1806 &  n_2310;
assign n_2348 = ~n_2346 & ~n_2347;
assign n_2349 =  x_2063 & ~n_2348;
assign n_2350 = ~x_2063 &  n_2348;
assign n_2351 = ~n_2349 & ~n_2350;
assign n_2352 =  n_1750 & ~n_2310;
assign n_2353 = ~x_2062 & ~n_1750;
assign n_2354 = ~n_2352 & ~n_2353;
assign n_2355 =  x_2062 &  n_2354;
assign n_2356 = ~x_2062 & ~n_2354;
assign n_2357 = ~n_2355 & ~n_2356;
assign n_2358 =  x_2061 & ~n_1761;
assign n_2359 =  i_178 &  n_1751;
assign n_2360 =  n_1761 &  n_2359;
assign n_2361 = ~n_2358 & ~n_2360;
assign n_2362 =  x_2061 & ~n_2361;
assign n_2363 = ~x_2061 &  n_2361;
assign n_2364 = ~n_2362 & ~n_2363;
assign n_2365 =  x_2060 & ~n_1770;
assign n_2366 =  n_1770 &  n_2359;
assign n_2367 = ~n_2365 & ~n_2366;
assign n_2368 =  x_2060 & ~n_2367;
assign n_2369 = ~x_2060 &  n_2367;
assign n_2370 = ~n_2368 & ~n_2369;
assign n_2371 =  x_2059 & ~n_1778;
assign n_2372 =  n_1778 &  n_2359;
assign n_2373 = ~n_2371 & ~n_2372;
assign n_2374 =  x_2059 & ~n_2373;
assign n_2375 = ~x_2059 &  n_2373;
assign n_2376 = ~n_2374 & ~n_2375;
assign n_2377 =  x_2058 & ~n_1785;
assign n_2378 =  n_1785 &  n_2359;
assign n_2379 = ~n_2377 & ~n_2378;
assign n_2380 =  x_2058 & ~n_2379;
assign n_2381 = ~x_2058 &  n_2379;
assign n_2382 = ~n_2380 & ~n_2381;
assign n_2383 =  x_2057 & ~n_1792;
assign n_2384 =  n_1792 &  n_2359;
assign n_2385 = ~n_2383 & ~n_2384;
assign n_2386 =  x_2057 & ~n_2385;
assign n_2387 = ~x_2057 &  n_2385;
assign n_2388 = ~n_2386 & ~n_2387;
assign n_2389 =  x_2056 & ~n_1799;
assign n_2390 =  n_1799 &  n_2359;
assign n_2391 = ~n_2389 & ~n_2390;
assign n_2392 =  x_2056 & ~n_2391;
assign n_2393 = ~x_2056 &  n_2391;
assign n_2394 = ~n_2392 & ~n_2393;
assign n_2395 =  x_2055 & ~n_1806;
assign n_2396 =  n_1806 &  n_2359;
assign n_2397 = ~n_2395 & ~n_2396;
assign n_2398 =  x_2055 & ~n_2397;
assign n_2399 = ~x_2055 &  n_2397;
assign n_2400 = ~n_2398 & ~n_2399;
assign n_2401 =  n_1750 & ~n_2359;
assign n_2402 = ~x_2054 & ~n_1750;
assign n_2403 = ~n_2401 & ~n_2402;
assign n_2404 =  x_2054 &  n_2403;
assign n_2405 = ~x_2054 & ~n_2403;
assign n_2406 = ~n_2404 & ~n_2405;
assign n_2407 =  x_2053 & ~n_1761;
assign n_2408 =  i_177 &  n_1751;
assign n_2409 =  n_1761 &  n_2408;
assign n_2410 = ~n_2407 & ~n_2409;
assign n_2411 =  x_2053 & ~n_2410;
assign n_2412 = ~x_2053 &  n_2410;
assign n_2413 = ~n_2411 & ~n_2412;
assign n_2414 =  x_2052 & ~n_1770;
assign n_2415 =  n_1770 &  n_2408;
assign n_2416 = ~n_2414 & ~n_2415;
assign n_2417 =  x_2052 & ~n_2416;
assign n_2418 = ~x_2052 &  n_2416;
assign n_2419 = ~n_2417 & ~n_2418;
assign n_2420 =  x_2051 & ~n_1778;
assign n_2421 =  n_1778 &  n_2408;
assign n_2422 = ~n_2420 & ~n_2421;
assign n_2423 =  x_2051 & ~n_2422;
assign n_2424 = ~x_2051 &  n_2422;
assign n_2425 = ~n_2423 & ~n_2424;
assign n_2426 =  x_2050 & ~n_1785;
assign n_2427 =  n_1785 &  n_2408;
assign n_2428 = ~n_2426 & ~n_2427;
assign n_2429 =  x_2050 & ~n_2428;
assign n_2430 = ~x_2050 &  n_2428;
assign n_2431 = ~n_2429 & ~n_2430;
assign n_2432 =  x_2049 & ~n_1792;
assign n_2433 =  n_1792 &  n_2408;
assign n_2434 = ~n_2432 & ~n_2433;
assign n_2435 =  x_2049 & ~n_2434;
assign n_2436 = ~x_2049 &  n_2434;
assign n_2437 = ~n_2435 & ~n_2436;
assign n_2438 =  x_2048 & ~n_1799;
assign n_2439 =  n_1799 &  n_2408;
assign n_2440 = ~n_2438 & ~n_2439;
assign n_2441 =  x_2048 & ~n_2440;
assign n_2442 = ~x_2048 &  n_2440;
assign n_2443 = ~n_2441 & ~n_2442;
assign n_2444 =  x_2047 & ~n_1806;
assign n_2445 =  n_1806 &  n_2408;
assign n_2446 = ~n_2444 & ~n_2445;
assign n_2447 =  x_2047 & ~n_2446;
assign n_2448 = ~x_2047 &  n_2446;
assign n_2449 = ~n_2447 & ~n_2448;
assign n_2450 =  n_1750 & ~n_2408;
assign n_2451 = ~x_2046 & ~n_1750;
assign n_2452 = ~n_2450 & ~n_2451;
assign n_2453 =  x_2046 &  n_2452;
assign n_2454 = ~x_2046 & ~n_2452;
assign n_2455 = ~n_2453 & ~n_2454;
assign n_2456 =  x_2045 & ~n_1761;
assign n_2457 =  i_176 &  n_1751;
assign n_2458 =  n_1761 &  n_2457;
assign n_2459 = ~n_2456 & ~n_2458;
assign n_2460 =  x_2045 & ~n_2459;
assign n_2461 = ~x_2045 &  n_2459;
assign n_2462 = ~n_2460 & ~n_2461;
assign n_2463 =  x_2044 & ~n_1770;
assign n_2464 =  n_1770 &  n_2457;
assign n_2465 = ~n_2463 & ~n_2464;
assign n_2466 =  x_2044 & ~n_2465;
assign n_2467 = ~x_2044 &  n_2465;
assign n_2468 = ~n_2466 & ~n_2467;
assign n_2469 =  x_2043 & ~n_1778;
assign n_2470 =  n_1778 &  n_2457;
assign n_2471 = ~n_2469 & ~n_2470;
assign n_2472 =  x_2043 & ~n_2471;
assign n_2473 = ~x_2043 &  n_2471;
assign n_2474 = ~n_2472 & ~n_2473;
assign n_2475 =  x_2042 & ~n_1785;
assign n_2476 =  n_1785 &  n_2457;
assign n_2477 = ~n_2475 & ~n_2476;
assign n_2478 =  x_2042 & ~n_2477;
assign n_2479 = ~x_2042 &  n_2477;
assign n_2480 = ~n_2478 & ~n_2479;
assign n_2481 =  x_2041 & ~n_1792;
assign n_2482 =  n_1792 &  n_2457;
assign n_2483 = ~n_2481 & ~n_2482;
assign n_2484 =  x_2041 & ~n_2483;
assign n_2485 = ~x_2041 &  n_2483;
assign n_2486 = ~n_2484 & ~n_2485;
assign n_2487 =  x_2040 & ~n_1799;
assign n_2488 =  n_1799 &  n_2457;
assign n_2489 = ~n_2487 & ~n_2488;
assign n_2490 =  x_2040 & ~n_2489;
assign n_2491 = ~x_2040 &  n_2489;
assign n_2492 = ~n_2490 & ~n_2491;
assign n_2493 =  x_2039 & ~n_1806;
assign n_2494 =  n_1806 &  n_2457;
assign n_2495 = ~n_2493 & ~n_2494;
assign n_2496 =  x_2039 & ~n_2495;
assign n_2497 = ~x_2039 &  n_2495;
assign n_2498 = ~n_2496 & ~n_2497;
assign n_2499 =  n_1750 & ~n_2457;
assign n_2500 = ~x_2038 & ~n_1750;
assign n_2501 = ~n_2499 & ~n_2500;
assign n_2502 =  x_2038 &  n_2501;
assign n_2503 = ~x_2038 & ~n_2501;
assign n_2504 = ~n_2502 & ~n_2503;
assign n_2505 =  x_2037 & ~n_1761;
assign n_2506 =  i_175 &  n_1751;
assign n_2507 =  n_1761 &  n_2506;
assign n_2508 = ~n_2505 & ~n_2507;
assign n_2509 =  x_2037 & ~n_2508;
assign n_2510 = ~x_2037 &  n_2508;
assign n_2511 = ~n_2509 & ~n_2510;
assign n_2512 =  x_2036 & ~n_1770;
assign n_2513 =  n_1770 &  n_2506;
assign n_2514 = ~n_2512 & ~n_2513;
assign n_2515 =  x_2036 & ~n_2514;
assign n_2516 = ~x_2036 &  n_2514;
assign n_2517 = ~n_2515 & ~n_2516;
assign n_2518 =  x_2035 & ~n_1778;
assign n_2519 =  n_1778 &  n_2506;
assign n_2520 = ~n_2518 & ~n_2519;
assign n_2521 =  x_2035 & ~n_2520;
assign n_2522 = ~x_2035 &  n_2520;
assign n_2523 = ~n_2521 & ~n_2522;
assign n_2524 =  x_2034 & ~n_1785;
assign n_2525 =  n_1785 &  n_2506;
assign n_2526 = ~n_2524 & ~n_2525;
assign n_2527 =  x_2034 & ~n_2526;
assign n_2528 = ~x_2034 &  n_2526;
assign n_2529 = ~n_2527 & ~n_2528;
assign n_2530 =  x_2033 & ~n_1792;
assign n_2531 =  n_1792 &  n_2506;
assign n_2532 = ~n_2530 & ~n_2531;
assign n_2533 =  x_2033 & ~n_2532;
assign n_2534 = ~x_2033 &  n_2532;
assign n_2535 = ~n_2533 & ~n_2534;
assign n_2536 =  x_2032 & ~n_1799;
assign n_2537 =  n_1799 &  n_2506;
assign n_2538 = ~n_2536 & ~n_2537;
assign n_2539 =  x_2032 & ~n_2538;
assign n_2540 = ~x_2032 &  n_2538;
assign n_2541 = ~n_2539 & ~n_2540;
assign n_2542 =  x_2031 & ~n_1806;
assign n_2543 =  n_1806 &  n_2506;
assign n_2544 = ~n_2542 & ~n_2543;
assign n_2545 =  x_2031 & ~n_2544;
assign n_2546 = ~x_2031 &  n_2544;
assign n_2547 = ~n_2545 & ~n_2546;
assign n_2548 =  n_1750 & ~n_2506;
assign n_2549 = ~x_2030 & ~n_1750;
assign n_2550 = ~n_2548 & ~n_2549;
assign n_2551 =  x_2030 &  n_2550;
assign n_2552 = ~x_2030 & ~n_2550;
assign n_2553 = ~n_2551 & ~n_2552;
assign n_2554 =  x_2029 & ~n_1761;
assign n_2555 =  i_174 &  n_1751;
assign n_2556 =  n_1761 &  n_2555;
assign n_2557 = ~n_2554 & ~n_2556;
assign n_2558 =  x_2029 & ~n_2557;
assign n_2559 = ~x_2029 &  n_2557;
assign n_2560 = ~n_2558 & ~n_2559;
assign n_2561 =  x_2028 & ~n_1770;
assign n_2562 =  n_1770 &  n_2555;
assign n_2563 = ~n_2561 & ~n_2562;
assign n_2564 =  x_2028 & ~n_2563;
assign n_2565 = ~x_2028 &  n_2563;
assign n_2566 = ~n_2564 & ~n_2565;
assign n_2567 =  x_2027 & ~n_1778;
assign n_2568 =  n_1778 &  n_2555;
assign n_2569 = ~n_2567 & ~n_2568;
assign n_2570 =  x_2027 & ~n_2569;
assign n_2571 = ~x_2027 &  n_2569;
assign n_2572 = ~n_2570 & ~n_2571;
assign n_2573 =  x_2026 & ~n_1785;
assign n_2574 =  n_1785 &  n_2555;
assign n_2575 = ~n_2573 & ~n_2574;
assign n_2576 =  x_2026 & ~n_2575;
assign n_2577 = ~x_2026 &  n_2575;
assign n_2578 = ~n_2576 & ~n_2577;
assign n_2579 =  x_2025 & ~n_1792;
assign n_2580 =  n_1792 &  n_2555;
assign n_2581 = ~n_2579 & ~n_2580;
assign n_2582 =  x_2025 & ~n_2581;
assign n_2583 = ~x_2025 &  n_2581;
assign n_2584 = ~n_2582 & ~n_2583;
assign n_2585 =  x_2024 & ~n_1799;
assign n_2586 =  n_1799 &  n_2555;
assign n_2587 = ~n_2585 & ~n_2586;
assign n_2588 =  x_2024 & ~n_2587;
assign n_2589 = ~x_2024 &  n_2587;
assign n_2590 = ~n_2588 & ~n_2589;
assign n_2591 =  x_2023 & ~n_1806;
assign n_2592 =  n_1806 &  n_2555;
assign n_2593 = ~n_2591 & ~n_2592;
assign n_2594 =  x_2023 & ~n_2593;
assign n_2595 = ~x_2023 &  n_2593;
assign n_2596 = ~n_2594 & ~n_2595;
assign n_2597 =  n_1750 & ~n_2555;
assign n_2598 = ~x_2022 & ~n_1750;
assign n_2599 = ~n_2597 & ~n_2598;
assign n_2600 =  x_2022 &  n_2599;
assign n_2601 = ~x_2022 & ~n_2599;
assign n_2602 = ~n_2600 & ~n_2601;
assign n_2603 =  x_2021 & ~n_1761;
assign n_2604 =  i_173 &  n_1751;
assign n_2605 =  n_1761 &  n_2604;
assign n_2606 = ~n_2603 & ~n_2605;
assign n_2607 =  x_2021 & ~n_2606;
assign n_2608 = ~x_2021 &  n_2606;
assign n_2609 = ~n_2607 & ~n_2608;
assign n_2610 =  x_2020 & ~n_1770;
assign n_2611 =  n_1770 &  n_2604;
assign n_2612 = ~n_2610 & ~n_2611;
assign n_2613 =  x_2020 & ~n_2612;
assign n_2614 = ~x_2020 &  n_2612;
assign n_2615 = ~n_2613 & ~n_2614;
assign n_2616 =  x_2019 & ~n_1778;
assign n_2617 =  n_1778 &  n_2604;
assign n_2618 = ~n_2616 & ~n_2617;
assign n_2619 =  x_2019 & ~n_2618;
assign n_2620 = ~x_2019 &  n_2618;
assign n_2621 = ~n_2619 & ~n_2620;
assign n_2622 =  x_2018 & ~n_1785;
assign n_2623 =  n_1785 &  n_2604;
assign n_2624 = ~n_2622 & ~n_2623;
assign n_2625 =  x_2018 & ~n_2624;
assign n_2626 = ~x_2018 &  n_2624;
assign n_2627 = ~n_2625 & ~n_2626;
assign n_2628 =  x_2017 & ~n_1792;
assign n_2629 =  n_1792 &  n_2604;
assign n_2630 = ~n_2628 & ~n_2629;
assign n_2631 =  x_2017 & ~n_2630;
assign n_2632 = ~x_2017 &  n_2630;
assign n_2633 = ~n_2631 & ~n_2632;
assign n_2634 =  x_2016 & ~n_1799;
assign n_2635 =  n_1799 &  n_2604;
assign n_2636 = ~n_2634 & ~n_2635;
assign n_2637 =  x_2016 & ~n_2636;
assign n_2638 = ~x_2016 &  n_2636;
assign n_2639 = ~n_2637 & ~n_2638;
assign n_2640 =  x_2015 & ~n_1806;
assign n_2641 =  n_1806 &  n_2604;
assign n_2642 = ~n_2640 & ~n_2641;
assign n_2643 =  x_2015 & ~n_2642;
assign n_2644 = ~x_2015 &  n_2642;
assign n_2645 = ~n_2643 & ~n_2644;
assign n_2646 =  n_1750 & ~n_2604;
assign n_2647 = ~x_2014 & ~n_1750;
assign n_2648 = ~n_2646 & ~n_2647;
assign n_2649 =  x_2014 &  n_2648;
assign n_2650 = ~x_2014 & ~n_2648;
assign n_2651 = ~n_2649 & ~n_2650;
assign n_2652 =  x_2013 & ~n_1761;
assign n_2653 =  i_172 &  n_1751;
assign n_2654 =  n_1761 &  n_2653;
assign n_2655 = ~n_2652 & ~n_2654;
assign n_2656 =  x_2013 & ~n_2655;
assign n_2657 = ~x_2013 &  n_2655;
assign n_2658 = ~n_2656 & ~n_2657;
assign n_2659 =  x_2012 & ~n_1770;
assign n_2660 =  n_1770 &  n_2653;
assign n_2661 = ~n_2659 & ~n_2660;
assign n_2662 =  x_2012 & ~n_2661;
assign n_2663 = ~x_2012 &  n_2661;
assign n_2664 = ~n_2662 & ~n_2663;
assign n_2665 =  x_2011 & ~n_1778;
assign n_2666 =  n_1778 &  n_2653;
assign n_2667 = ~n_2665 & ~n_2666;
assign n_2668 =  x_2011 & ~n_2667;
assign n_2669 = ~x_2011 &  n_2667;
assign n_2670 = ~n_2668 & ~n_2669;
assign n_2671 =  x_2010 & ~n_1785;
assign n_2672 =  n_1785 &  n_2653;
assign n_2673 = ~n_2671 & ~n_2672;
assign n_2674 =  x_2010 & ~n_2673;
assign n_2675 = ~x_2010 &  n_2673;
assign n_2676 = ~n_2674 & ~n_2675;
assign n_2677 =  x_2009 & ~n_1792;
assign n_2678 =  n_1792 &  n_2653;
assign n_2679 = ~n_2677 & ~n_2678;
assign n_2680 =  x_2009 & ~n_2679;
assign n_2681 = ~x_2009 &  n_2679;
assign n_2682 = ~n_2680 & ~n_2681;
assign n_2683 =  x_2008 & ~n_1799;
assign n_2684 =  n_1799 &  n_2653;
assign n_2685 = ~n_2683 & ~n_2684;
assign n_2686 =  x_2008 & ~n_2685;
assign n_2687 = ~x_2008 &  n_2685;
assign n_2688 = ~n_2686 & ~n_2687;
assign n_2689 =  x_2007 & ~n_1806;
assign n_2690 =  n_1806 &  n_2653;
assign n_2691 = ~n_2689 & ~n_2690;
assign n_2692 =  x_2007 & ~n_2691;
assign n_2693 = ~x_2007 &  n_2691;
assign n_2694 = ~n_2692 & ~n_2693;
assign n_2695 =  n_1750 & ~n_2653;
assign n_2696 = ~x_2006 & ~n_1750;
assign n_2697 = ~n_2695 & ~n_2696;
assign n_2698 =  x_2006 &  n_2697;
assign n_2699 = ~x_2006 & ~n_2697;
assign n_2700 = ~n_2698 & ~n_2699;
assign n_2701 =  x_2005 & ~n_1761;
assign n_2702 =  i_171 &  n_1751;
assign n_2703 =  n_1761 &  n_2702;
assign n_2704 = ~n_2701 & ~n_2703;
assign n_2705 =  x_2005 & ~n_2704;
assign n_2706 = ~x_2005 &  n_2704;
assign n_2707 = ~n_2705 & ~n_2706;
assign n_2708 =  x_2004 & ~n_1770;
assign n_2709 =  n_1770 &  n_2702;
assign n_2710 = ~n_2708 & ~n_2709;
assign n_2711 =  x_2004 & ~n_2710;
assign n_2712 = ~x_2004 &  n_2710;
assign n_2713 = ~n_2711 & ~n_2712;
assign n_2714 =  x_2003 & ~n_1778;
assign n_2715 =  n_1778 &  n_2702;
assign n_2716 = ~n_2714 & ~n_2715;
assign n_2717 =  x_2003 & ~n_2716;
assign n_2718 = ~x_2003 &  n_2716;
assign n_2719 = ~n_2717 & ~n_2718;
assign n_2720 =  x_2002 & ~n_1785;
assign n_2721 =  n_1785 &  n_2702;
assign n_2722 = ~n_2720 & ~n_2721;
assign n_2723 =  x_2002 & ~n_2722;
assign n_2724 = ~x_2002 &  n_2722;
assign n_2725 = ~n_2723 & ~n_2724;
assign n_2726 =  x_2001 & ~n_1792;
assign n_2727 =  n_1792 &  n_2702;
assign n_2728 = ~n_2726 & ~n_2727;
assign n_2729 =  x_2001 & ~n_2728;
assign n_2730 = ~x_2001 &  n_2728;
assign n_2731 = ~n_2729 & ~n_2730;
assign n_2732 =  x_2000 & ~n_1799;
assign n_2733 =  n_1799 &  n_2702;
assign n_2734 = ~n_2732 & ~n_2733;
assign n_2735 =  x_2000 & ~n_2734;
assign n_2736 = ~x_2000 &  n_2734;
assign n_2737 = ~n_2735 & ~n_2736;
assign n_2738 =  x_1999 & ~n_1806;
assign n_2739 =  n_1806 &  n_2702;
assign n_2740 = ~n_2738 & ~n_2739;
assign n_2741 =  x_1999 & ~n_2740;
assign n_2742 = ~x_1999 &  n_2740;
assign n_2743 = ~n_2741 & ~n_2742;
assign n_2744 =  n_1750 & ~n_2702;
assign n_2745 = ~x_1998 & ~n_1750;
assign n_2746 = ~n_2744 & ~n_2745;
assign n_2747 =  x_1998 &  n_2746;
assign n_2748 = ~x_1998 & ~n_2746;
assign n_2749 = ~n_2747 & ~n_2748;
assign n_2750 =  x_1997 & ~n_1761;
assign n_2751 =  i_170 &  n_1751;
assign n_2752 =  n_1761 &  n_2751;
assign n_2753 = ~n_2750 & ~n_2752;
assign n_2754 =  x_1997 & ~n_2753;
assign n_2755 = ~x_1997 &  n_2753;
assign n_2756 = ~n_2754 & ~n_2755;
assign n_2757 =  x_1996 & ~n_1770;
assign n_2758 =  n_1770 &  n_2751;
assign n_2759 = ~n_2757 & ~n_2758;
assign n_2760 =  x_1996 & ~n_2759;
assign n_2761 = ~x_1996 &  n_2759;
assign n_2762 = ~n_2760 & ~n_2761;
assign n_2763 =  x_1995 & ~n_1778;
assign n_2764 =  n_1778 &  n_2751;
assign n_2765 = ~n_2763 & ~n_2764;
assign n_2766 =  x_1995 & ~n_2765;
assign n_2767 = ~x_1995 &  n_2765;
assign n_2768 = ~n_2766 & ~n_2767;
assign n_2769 =  x_1994 & ~n_1785;
assign n_2770 =  n_1785 &  n_2751;
assign n_2771 = ~n_2769 & ~n_2770;
assign n_2772 =  x_1994 & ~n_2771;
assign n_2773 = ~x_1994 &  n_2771;
assign n_2774 = ~n_2772 & ~n_2773;
assign n_2775 =  x_1993 & ~n_1792;
assign n_2776 =  n_1792 &  n_2751;
assign n_2777 = ~n_2775 & ~n_2776;
assign n_2778 =  x_1993 & ~n_2777;
assign n_2779 = ~x_1993 &  n_2777;
assign n_2780 = ~n_2778 & ~n_2779;
assign n_2781 =  x_1992 & ~n_1799;
assign n_2782 =  n_1799 &  n_2751;
assign n_2783 = ~n_2781 & ~n_2782;
assign n_2784 =  x_1992 & ~n_2783;
assign n_2785 = ~x_1992 &  n_2783;
assign n_2786 = ~n_2784 & ~n_2785;
assign n_2787 =  x_1991 & ~n_1806;
assign n_2788 =  n_1806 &  n_2751;
assign n_2789 = ~n_2787 & ~n_2788;
assign n_2790 =  x_1991 & ~n_2789;
assign n_2791 = ~x_1991 &  n_2789;
assign n_2792 = ~n_2790 & ~n_2791;
assign n_2793 =  n_1750 & ~n_2751;
assign n_2794 = ~x_1990 & ~n_1750;
assign n_2795 = ~n_2793 & ~n_2794;
assign n_2796 =  x_1990 &  n_2795;
assign n_2797 = ~x_1990 & ~n_2795;
assign n_2798 = ~n_2796 & ~n_2797;
assign n_2799 =  x_1989 & ~n_1761;
assign n_2800 =  i_169 &  n_1751;
assign n_2801 =  n_1761 &  n_2800;
assign n_2802 = ~n_2799 & ~n_2801;
assign n_2803 =  x_1989 & ~n_2802;
assign n_2804 = ~x_1989 &  n_2802;
assign n_2805 = ~n_2803 & ~n_2804;
assign n_2806 =  x_1988 & ~n_1770;
assign n_2807 =  n_1770 &  n_2800;
assign n_2808 = ~n_2806 & ~n_2807;
assign n_2809 =  x_1988 & ~n_2808;
assign n_2810 = ~x_1988 &  n_2808;
assign n_2811 = ~n_2809 & ~n_2810;
assign n_2812 =  x_1987 & ~n_1778;
assign n_2813 =  n_1778 &  n_2800;
assign n_2814 = ~n_2812 & ~n_2813;
assign n_2815 =  x_1987 & ~n_2814;
assign n_2816 = ~x_1987 &  n_2814;
assign n_2817 = ~n_2815 & ~n_2816;
assign n_2818 =  x_1986 & ~n_1785;
assign n_2819 =  n_1785 &  n_2800;
assign n_2820 = ~n_2818 & ~n_2819;
assign n_2821 =  x_1986 & ~n_2820;
assign n_2822 = ~x_1986 &  n_2820;
assign n_2823 = ~n_2821 & ~n_2822;
assign n_2824 =  x_1985 & ~n_1792;
assign n_2825 =  n_1792 &  n_2800;
assign n_2826 = ~n_2824 & ~n_2825;
assign n_2827 =  x_1985 & ~n_2826;
assign n_2828 = ~x_1985 &  n_2826;
assign n_2829 = ~n_2827 & ~n_2828;
assign n_2830 =  x_1984 & ~n_1799;
assign n_2831 =  n_1799 &  n_2800;
assign n_2832 = ~n_2830 & ~n_2831;
assign n_2833 =  x_1984 & ~n_2832;
assign n_2834 = ~x_1984 &  n_2832;
assign n_2835 = ~n_2833 & ~n_2834;
assign n_2836 =  x_1983 & ~n_1806;
assign n_2837 =  n_1806 &  n_2800;
assign n_2838 = ~n_2836 & ~n_2837;
assign n_2839 =  x_1983 & ~n_2838;
assign n_2840 = ~x_1983 &  n_2838;
assign n_2841 = ~n_2839 & ~n_2840;
assign n_2842 =  n_1750 & ~n_2800;
assign n_2843 = ~x_1982 & ~n_1750;
assign n_2844 = ~n_2842 & ~n_2843;
assign n_2845 =  x_1982 &  n_2844;
assign n_2846 = ~x_1982 & ~n_2844;
assign n_2847 = ~n_2845 & ~n_2846;
assign n_2848 =  x_1981 & ~n_1761;
assign n_2849 =  i_168 &  n_1751;
assign n_2850 =  n_1761 &  n_2849;
assign n_2851 = ~n_2848 & ~n_2850;
assign n_2852 =  x_1981 & ~n_2851;
assign n_2853 = ~x_1981 &  n_2851;
assign n_2854 = ~n_2852 & ~n_2853;
assign n_2855 =  x_1980 & ~n_1770;
assign n_2856 =  n_1770 &  n_2849;
assign n_2857 = ~n_2855 & ~n_2856;
assign n_2858 =  x_1980 & ~n_2857;
assign n_2859 = ~x_1980 &  n_2857;
assign n_2860 = ~n_2858 & ~n_2859;
assign n_2861 =  x_1979 & ~n_1778;
assign n_2862 =  n_1778 &  n_2849;
assign n_2863 = ~n_2861 & ~n_2862;
assign n_2864 =  x_1979 & ~n_2863;
assign n_2865 = ~x_1979 &  n_2863;
assign n_2866 = ~n_2864 & ~n_2865;
assign n_2867 =  x_1978 & ~n_1785;
assign n_2868 =  n_1785 &  n_2849;
assign n_2869 = ~n_2867 & ~n_2868;
assign n_2870 =  x_1978 & ~n_2869;
assign n_2871 = ~x_1978 &  n_2869;
assign n_2872 = ~n_2870 & ~n_2871;
assign n_2873 =  x_1977 & ~n_1792;
assign n_2874 =  n_1792 &  n_2849;
assign n_2875 = ~n_2873 & ~n_2874;
assign n_2876 =  x_1977 & ~n_2875;
assign n_2877 = ~x_1977 &  n_2875;
assign n_2878 = ~n_2876 & ~n_2877;
assign n_2879 =  x_1976 & ~n_1799;
assign n_2880 =  n_1799 &  n_2849;
assign n_2881 = ~n_2879 & ~n_2880;
assign n_2882 =  x_1976 & ~n_2881;
assign n_2883 = ~x_1976 &  n_2881;
assign n_2884 = ~n_2882 & ~n_2883;
assign n_2885 =  x_1975 & ~n_1806;
assign n_2886 =  n_1806 &  n_2849;
assign n_2887 = ~n_2885 & ~n_2886;
assign n_2888 =  x_1975 & ~n_2887;
assign n_2889 = ~x_1975 &  n_2887;
assign n_2890 = ~n_2888 & ~n_2889;
assign n_2891 =  n_1750 & ~n_2849;
assign n_2892 = ~x_1974 & ~n_1750;
assign n_2893 = ~n_2891 & ~n_2892;
assign n_2894 =  x_1974 &  n_2893;
assign n_2895 = ~x_1974 & ~n_2893;
assign n_2896 = ~n_2894 & ~n_2895;
assign n_2897 =  x_1973 & ~n_1761;
assign n_2898 =  i_167 &  n_1751;
assign n_2899 =  n_1761 &  n_2898;
assign n_2900 = ~n_2897 & ~n_2899;
assign n_2901 =  x_1973 & ~n_2900;
assign n_2902 = ~x_1973 &  n_2900;
assign n_2903 = ~n_2901 & ~n_2902;
assign n_2904 =  x_1972 & ~n_1770;
assign n_2905 =  n_1770 &  n_2898;
assign n_2906 = ~n_2904 & ~n_2905;
assign n_2907 =  x_1972 & ~n_2906;
assign n_2908 = ~x_1972 &  n_2906;
assign n_2909 = ~n_2907 & ~n_2908;
assign n_2910 =  x_1971 & ~n_1778;
assign n_2911 =  n_1778 &  n_2898;
assign n_2912 = ~n_2910 & ~n_2911;
assign n_2913 =  x_1971 & ~n_2912;
assign n_2914 = ~x_1971 &  n_2912;
assign n_2915 = ~n_2913 & ~n_2914;
assign n_2916 =  x_1970 & ~n_1785;
assign n_2917 =  n_1785 &  n_2898;
assign n_2918 = ~n_2916 & ~n_2917;
assign n_2919 =  x_1970 & ~n_2918;
assign n_2920 = ~x_1970 &  n_2918;
assign n_2921 = ~n_2919 & ~n_2920;
assign n_2922 =  x_1969 & ~n_1792;
assign n_2923 =  n_1792 &  n_2898;
assign n_2924 = ~n_2922 & ~n_2923;
assign n_2925 =  x_1969 & ~n_2924;
assign n_2926 = ~x_1969 &  n_2924;
assign n_2927 = ~n_2925 & ~n_2926;
assign n_2928 =  x_1968 & ~n_1799;
assign n_2929 =  n_1799 &  n_2898;
assign n_2930 = ~n_2928 & ~n_2929;
assign n_2931 =  x_1968 & ~n_2930;
assign n_2932 = ~x_1968 &  n_2930;
assign n_2933 = ~n_2931 & ~n_2932;
assign n_2934 =  x_1967 & ~n_1806;
assign n_2935 =  n_1806 &  n_2898;
assign n_2936 = ~n_2934 & ~n_2935;
assign n_2937 =  x_1967 & ~n_2936;
assign n_2938 = ~x_1967 &  n_2936;
assign n_2939 = ~n_2937 & ~n_2938;
assign n_2940 =  n_1750 & ~n_2898;
assign n_2941 = ~x_1966 & ~n_1750;
assign n_2942 = ~n_2940 & ~n_2941;
assign n_2943 =  x_1966 &  n_2942;
assign n_2944 = ~x_1966 & ~n_2942;
assign n_2945 = ~n_2943 & ~n_2944;
assign n_2946 =  x_1965 & ~n_1761;
assign n_2947 =  i_166 &  n_1751;
assign n_2948 =  n_1761 &  n_2947;
assign n_2949 = ~n_2946 & ~n_2948;
assign n_2950 =  x_1965 & ~n_2949;
assign n_2951 = ~x_1965 &  n_2949;
assign n_2952 = ~n_2950 & ~n_2951;
assign n_2953 =  x_1964 & ~n_1770;
assign n_2954 =  n_1770 &  n_2947;
assign n_2955 = ~n_2953 & ~n_2954;
assign n_2956 =  x_1964 & ~n_2955;
assign n_2957 = ~x_1964 &  n_2955;
assign n_2958 = ~n_2956 & ~n_2957;
assign n_2959 =  x_1963 & ~n_1778;
assign n_2960 =  n_1778 &  n_2947;
assign n_2961 = ~n_2959 & ~n_2960;
assign n_2962 =  x_1963 & ~n_2961;
assign n_2963 = ~x_1963 &  n_2961;
assign n_2964 = ~n_2962 & ~n_2963;
assign n_2965 =  x_1962 & ~n_1785;
assign n_2966 =  n_1785 &  n_2947;
assign n_2967 = ~n_2965 & ~n_2966;
assign n_2968 =  x_1962 & ~n_2967;
assign n_2969 = ~x_1962 &  n_2967;
assign n_2970 = ~n_2968 & ~n_2969;
assign n_2971 =  x_1961 & ~n_1792;
assign n_2972 =  n_1792 &  n_2947;
assign n_2973 = ~n_2971 & ~n_2972;
assign n_2974 =  x_1961 & ~n_2973;
assign n_2975 = ~x_1961 &  n_2973;
assign n_2976 = ~n_2974 & ~n_2975;
assign n_2977 =  x_1960 & ~n_1799;
assign n_2978 =  n_1799 &  n_2947;
assign n_2979 = ~n_2977 & ~n_2978;
assign n_2980 =  x_1960 & ~n_2979;
assign n_2981 = ~x_1960 &  n_2979;
assign n_2982 = ~n_2980 & ~n_2981;
assign n_2983 =  x_1959 & ~n_1806;
assign n_2984 =  n_1806 &  n_2947;
assign n_2985 = ~n_2983 & ~n_2984;
assign n_2986 =  x_1959 & ~n_2985;
assign n_2987 = ~x_1959 &  n_2985;
assign n_2988 = ~n_2986 & ~n_2987;
assign n_2989 =  n_1750 & ~n_2947;
assign n_2990 = ~x_1958 & ~n_1750;
assign n_2991 = ~n_2989 & ~n_2990;
assign n_2992 =  x_1958 &  n_2991;
assign n_2993 = ~x_1958 & ~n_2991;
assign n_2994 = ~n_2992 & ~n_2993;
assign n_2995 =  x_1957 & ~n_1761;
assign n_2996 =  i_165 &  n_1751;
assign n_2997 =  n_1761 &  n_2996;
assign n_2998 = ~n_2995 & ~n_2997;
assign n_2999 =  x_1957 & ~n_2998;
assign n_3000 = ~x_1957 &  n_2998;
assign n_3001 = ~n_2999 & ~n_3000;
assign n_3002 =  x_1956 & ~n_1770;
assign n_3003 =  n_1770 &  n_2996;
assign n_3004 = ~n_3002 & ~n_3003;
assign n_3005 =  x_1956 & ~n_3004;
assign n_3006 = ~x_1956 &  n_3004;
assign n_3007 = ~n_3005 & ~n_3006;
assign n_3008 =  x_1955 & ~n_1778;
assign n_3009 =  n_1778 &  n_2996;
assign n_3010 = ~n_3008 & ~n_3009;
assign n_3011 =  x_1955 & ~n_3010;
assign n_3012 = ~x_1955 &  n_3010;
assign n_3013 = ~n_3011 & ~n_3012;
assign n_3014 =  x_1954 & ~n_1785;
assign n_3015 =  n_1785 &  n_2996;
assign n_3016 = ~n_3014 & ~n_3015;
assign n_3017 =  x_1954 & ~n_3016;
assign n_3018 = ~x_1954 &  n_3016;
assign n_3019 = ~n_3017 & ~n_3018;
assign n_3020 =  x_1953 & ~n_1792;
assign n_3021 =  n_1792 &  n_2996;
assign n_3022 = ~n_3020 & ~n_3021;
assign n_3023 =  x_1953 & ~n_3022;
assign n_3024 = ~x_1953 &  n_3022;
assign n_3025 = ~n_3023 & ~n_3024;
assign n_3026 =  x_1952 & ~n_1799;
assign n_3027 =  n_1799 &  n_2996;
assign n_3028 = ~n_3026 & ~n_3027;
assign n_3029 =  x_1952 & ~n_3028;
assign n_3030 = ~x_1952 &  n_3028;
assign n_3031 = ~n_3029 & ~n_3030;
assign n_3032 =  x_1951 & ~n_1806;
assign n_3033 =  n_1806 &  n_2996;
assign n_3034 = ~n_3032 & ~n_3033;
assign n_3035 =  x_1951 & ~n_3034;
assign n_3036 = ~x_1951 &  n_3034;
assign n_3037 = ~n_3035 & ~n_3036;
assign n_3038 =  n_1750 & ~n_2996;
assign n_3039 = ~x_1950 & ~n_1750;
assign n_3040 = ~n_3038 & ~n_3039;
assign n_3041 =  x_1950 &  n_3040;
assign n_3042 = ~x_1950 & ~n_3040;
assign n_3043 = ~n_3041 & ~n_3042;
assign n_3044 =  x_1949 & ~n_1761;
assign n_3045 =  i_164 &  n_1751;
assign n_3046 =  n_1761 &  n_3045;
assign n_3047 = ~n_3044 & ~n_3046;
assign n_3048 =  x_1949 & ~n_3047;
assign n_3049 = ~x_1949 &  n_3047;
assign n_3050 = ~n_3048 & ~n_3049;
assign n_3051 =  x_1948 & ~n_1770;
assign n_3052 =  n_1770 &  n_3045;
assign n_3053 = ~n_3051 & ~n_3052;
assign n_3054 =  x_1948 & ~n_3053;
assign n_3055 = ~x_1948 &  n_3053;
assign n_3056 = ~n_3054 & ~n_3055;
assign n_3057 =  x_1947 & ~n_1778;
assign n_3058 =  n_1778 &  n_3045;
assign n_3059 = ~n_3057 & ~n_3058;
assign n_3060 =  x_1947 & ~n_3059;
assign n_3061 = ~x_1947 &  n_3059;
assign n_3062 = ~n_3060 & ~n_3061;
assign n_3063 =  x_1946 & ~n_1785;
assign n_3064 =  n_1785 &  n_3045;
assign n_3065 = ~n_3063 & ~n_3064;
assign n_3066 =  x_1946 & ~n_3065;
assign n_3067 = ~x_1946 &  n_3065;
assign n_3068 = ~n_3066 & ~n_3067;
assign n_3069 =  x_1945 & ~n_1792;
assign n_3070 =  n_1792 &  n_3045;
assign n_3071 = ~n_3069 & ~n_3070;
assign n_3072 =  x_1945 & ~n_3071;
assign n_3073 = ~x_1945 &  n_3071;
assign n_3074 = ~n_3072 & ~n_3073;
assign n_3075 =  x_1944 & ~n_1799;
assign n_3076 =  n_1799 &  n_3045;
assign n_3077 = ~n_3075 & ~n_3076;
assign n_3078 =  x_1944 & ~n_3077;
assign n_3079 = ~x_1944 &  n_3077;
assign n_3080 = ~n_3078 & ~n_3079;
assign n_3081 =  x_1943 & ~n_1806;
assign n_3082 =  n_1806 &  n_3045;
assign n_3083 = ~n_3081 & ~n_3082;
assign n_3084 =  x_1943 & ~n_3083;
assign n_3085 = ~x_1943 &  n_3083;
assign n_3086 = ~n_3084 & ~n_3085;
assign n_3087 =  n_1750 & ~n_3045;
assign n_3088 = ~x_1942 & ~n_1750;
assign n_3089 = ~n_3087 & ~n_3088;
assign n_3090 =  x_1942 &  n_3089;
assign n_3091 = ~x_1942 & ~n_3089;
assign n_3092 = ~n_3090 & ~n_3091;
assign n_3093 =  x_1941 & ~n_1761;
assign n_3094 =  i_163 &  n_1751;
assign n_3095 =  n_1761 &  n_3094;
assign n_3096 = ~n_3093 & ~n_3095;
assign n_3097 =  x_1941 & ~n_3096;
assign n_3098 = ~x_1941 &  n_3096;
assign n_3099 = ~n_3097 & ~n_3098;
assign n_3100 =  x_1940 & ~n_1770;
assign n_3101 =  n_1770 &  n_3094;
assign n_3102 = ~n_3100 & ~n_3101;
assign n_3103 =  x_1940 & ~n_3102;
assign n_3104 = ~x_1940 &  n_3102;
assign n_3105 = ~n_3103 & ~n_3104;
assign n_3106 =  x_1939 & ~n_1778;
assign n_3107 =  n_1778 &  n_3094;
assign n_3108 = ~n_3106 & ~n_3107;
assign n_3109 =  x_1939 & ~n_3108;
assign n_3110 = ~x_1939 &  n_3108;
assign n_3111 = ~n_3109 & ~n_3110;
assign n_3112 =  x_1938 & ~n_1785;
assign n_3113 =  n_1785 &  n_3094;
assign n_3114 = ~n_3112 & ~n_3113;
assign n_3115 =  x_1938 & ~n_3114;
assign n_3116 = ~x_1938 &  n_3114;
assign n_3117 = ~n_3115 & ~n_3116;
assign n_3118 =  x_1937 & ~n_1792;
assign n_3119 =  n_1792 &  n_3094;
assign n_3120 = ~n_3118 & ~n_3119;
assign n_3121 =  x_1937 & ~n_3120;
assign n_3122 = ~x_1937 &  n_3120;
assign n_3123 = ~n_3121 & ~n_3122;
assign n_3124 =  x_1936 & ~n_1799;
assign n_3125 =  n_1799 &  n_3094;
assign n_3126 = ~n_3124 & ~n_3125;
assign n_3127 =  x_1936 & ~n_3126;
assign n_3128 = ~x_1936 &  n_3126;
assign n_3129 = ~n_3127 & ~n_3128;
assign n_3130 =  x_1935 & ~n_1806;
assign n_3131 =  n_1806 &  n_3094;
assign n_3132 = ~n_3130 & ~n_3131;
assign n_3133 =  x_1935 & ~n_3132;
assign n_3134 = ~x_1935 &  n_3132;
assign n_3135 = ~n_3133 & ~n_3134;
assign n_3136 =  n_1750 & ~n_3094;
assign n_3137 = ~x_1934 & ~n_1750;
assign n_3138 = ~n_3136 & ~n_3137;
assign n_3139 =  x_1934 &  n_3138;
assign n_3140 = ~x_1934 & ~n_3138;
assign n_3141 = ~n_3139 & ~n_3140;
assign n_3142 =  x_1933 & ~n_1761;
assign n_3143 =  i_162 &  n_1751;
assign n_3144 =  n_1761 &  n_3143;
assign n_3145 = ~n_3142 & ~n_3144;
assign n_3146 =  x_1933 & ~n_3145;
assign n_3147 = ~x_1933 &  n_3145;
assign n_3148 = ~n_3146 & ~n_3147;
assign n_3149 =  x_1932 & ~n_1770;
assign n_3150 =  n_1770 &  n_3143;
assign n_3151 = ~n_3149 & ~n_3150;
assign n_3152 =  x_1932 & ~n_3151;
assign n_3153 = ~x_1932 &  n_3151;
assign n_3154 = ~n_3152 & ~n_3153;
assign n_3155 =  x_1931 & ~n_1778;
assign n_3156 =  n_1778 &  n_3143;
assign n_3157 = ~n_3155 & ~n_3156;
assign n_3158 =  x_1931 & ~n_3157;
assign n_3159 = ~x_1931 &  n_3157;
assign n_3160 = ~n_3158 & ~n_3159;
assign n_3161 =  x_1930 & ~n_1785;
assign n_3162 =  n_1785 &  n_3143;
assign n_3163 = ~n_3161 & ~n_3162;
assign n_3164 =  x_1930 & ~n_3163;
assign n_3165 = ~x_1930 &  n_3163;
assign n_3166 = ~n_3164 & ~n_3165;
assign n_3167 =  x_1929 & ~n_1792;
assign n_3168 =  n_1792 &  n_3143;
assign n_3169 = ~n_3167 & ~n_3168;
assign n_3170 =  x_1929 & ~n_3169;
assign n_3171 = ~x_1929 &  n_3169;
assign n_3172 = ~n_3170 & ~n_3171;
assign n_3173 =  x_1928 & ~n_1799;
assign n_3174 =  n_1799 &  n_3143;
assign n_3175 = ~n_3173 & ~n_3174;
assign n_3176 =  x_1928 & ~n_3175;
assign n_3177 = ~x_1928 &  n_3175;
assign n_3178 = ~n_3176 & ~n_3177;
assign n_3179 =  x_1927 & ~n_1806;
assign n_3180 =  n_1806 &  n_3143;
assign n_3181 = ~n_3179 & ~n_3180;
assign n_3182 =  x_1927 & ~n_3181;
assign n_3183 = ~x_1927 &  n_3181;
assign n_3184 = ~n_3182 & ~n_3183;
assign n_3185 =  n_1750 & ~n_3143;
assign n_3186 = ~x_1926 & ~n_1750;
assign n_3187 = ~n_3185 & ~n_3186;
assign n_3188 =  x_1926 &  n_3187;
assign n_3189 = ~x_1926 & ~n_3187;
assign n_3190 = ~n_3188 & ~n_3189;
assign n_3191 =  x_1925 & ~n_1761;
assign n_3192 =  i_161 &  n_1751;
assign n_3193 =  n_1761 &  n_3192;
assign n_3194 = ~n_3191 & ~n_3193;
assign n_3195 =  x_1925 & ~n_3194;
assign n_3196 = ~x_1925 &  n_3194;
assign n_3197 = ~n_3195 & ~n_3196;
assign n_3198 =  x_1924 & ~n_1770;
assign n_3199 =  n_1770 &  n_3192;
assign n_3200 = ~n_3198 & ~n_3199;
assign n_3201 =  x_1924 & ~n_3200;
assign n_3202 = ~x_1924 &  n_3200;
assign n_3203 = ~n_3201 & ~n_3202;
assign n_3204 =  x_1923 & ~n_1778;
assign n_3205 =  n_1778 &  n_3192;
assign n_3206 = ~n_3204 & ~n_3205;
assign n_3207 =  x_1923 & ~n_3206;
assign n_3208 = ~x_1923 &  n_3206;
assign n_3209 = ~n_3207 & ~n_3208;
assign n_3210 =  x_1922 & ~n_1785;
assign n_3211 =  n_1785 &  n_3192;
assign n_3212 = ~n_3210 & ~n_3211;
assign n_3213 =  x_1922 & ~n_3212;
assign n_3214 = ~x_1922 &  n_3212;
assign n_3215 = ~n_3213 & ~n_3214;
assign n_3216 =  x_1921 & ~n_1792;
assign n_3217 =  n_1792 &  n_3192;
assign n_3218 = ~n_3216 & ~n_3217;
assign n_3219 =  x_1921 & ~n_3218;
assign n_3220 = ~x_1921 &  n_3218;
assign n_3221 = ~n_3219 & ~n_3220;
assign n_3222 =  x_1920 & ~n_1799;
assign n_3223 =  n_1799 &  n_3192;
assign n_3224 = ~n_3222 & ~n_3223;
assign n_3225 =  x_1920 & ~n_3224;
assign n_3226 = ~x_1920 &  n_3224;
assign n_3227 = ~n_3225 & ~n_3226;
assign n_3228 =  x_1919 & ~n_1806;
assign n_3229 =  n_1806 &  n_3192;
assign n_3230 = ~n_3228 & ~n_3229;
assign n_3231 =  x_1919 & ~n_3230;
assign n_3232 = ~x_1919 &  n_3230;
assign n_3233 = ~n_3231 & ~n_3232;
assign n_3234 =  n_1750 & ~n_3192;
assign n_3235 = ~x_1918 & ~n_1750;
assign n_3236 = ~n_3234 & ~n_3235;
assign n_3237 =  x_1918 &  n_3236;
assign n_3238 = ~x_1918 & ~n_3236;
assign n_3239 = ~n_3237 & ~n_3238;
assign n_3240 = ~x_1745 &  x_1746;
assign n_3241 =  x_1747 &  n_3240;
assign n_3242 =  x_1719 & ~n_3241;
assign n_3243 = ~x_1486 & ~n_3242;
assign n_3244 =  x_1751 & ~x_1752;
assign n_3245 =  x_1763 &  n_3244;
assign n_3246 = ~x_1484 & ~x_1485;
assign n_3247 = ~x_1483 &  n_3246;
assign n_3248 =  x_1761 &  x_1762;
assign n_3249 = ~n_3247 &  n_3248;
assign n_3250 =  n_3245 &  n_3249;
assign n_3251 = ~n_3243 &  n_3250;
assign n_3252 =  x_1751 &  x_1752;
assign n_3253 =  x_1763 &  n_3252;
assign n_3254 =  x_1762 & ~n_3253;
assign n_3255 = ~n_3251 &  n_3254;
assign n_3256 =  x_1745 & ~x_1746;
assign n_3257 =  x_1747 &  n_3256;
assign n_3258 =  n_3247 &  n_3245;
assign n_3259 = ~x_1762 & ~n_3258;
assign n_3260 =  n_3257 & ~n_3259;
assign n_3261 = ~n_3255 &  n_3260;
assign n_3262 = ~i_217 & ~i_218;
assign n_3263 =  x_295 & ~n_3262;
assign n_3264 =  n_1191 & ~n_3263;
assign n_3265 =  n_3240 &  n_3244;
assign n_3266 = ~x_1747 & ~x_1748;
assign n_3267 =  x_311 &  n_3266;
assign n_3268 = ~x_1747 &  n_3256;
assign n_3269 = ~n_3267 & ~n_3268;
assign n_3270 = ~n_3265 &  n_3269;
assign n_3271 = ~n_3264 &  n_3270;
assign n_3272 = ~n_3261 &  n_3271;
assign n_3273 = ~x_1747 &  n_3272;
assign n_3274 = ~n_3243 &  n_3256;
assign n_3275 = ~n_3246 &  n_3274;
assign n_3276 = ~x_1747 & ~n_3240;
assign n_3277 = ~n_3275 &  n_3276;
assign n_3278 = ~n_3251 &  n_3257;
assign n_3279 = ~x_1747 &  x_1753;
assign n_3280 =  n_3265 &  n_3279;
assign n_3281 =  x_1751 & ~x_1763;
assign n_3282 = ~x_1748 & ~n_3281;
assign n_3283 = ~n_3280 & ~n_3282;
assign n_3284 = ~n_3278 &  n_3283;
assign n_3285 = ~n_3277 &  n_3284;
assign n_3286 = ~n_3273 & ~n_3285;
assign n_3287 =  x_1749 &  x_1751;
assign n_3288 = ~n_3287 &  n_3272;
assign n_3289 = ~n_1192 & ~n_3241;
assign n_3290 =  n_3288 &  n_3289;
assign n_3291 = ~x_1745 &  n_3290;
assign n_3292 =  n_3240 & ~n_3258;
assign n_3293 = ~x_1745 &  x_1747;
assign n_3294 = ~x_1747 &  n_1191;
assign n_3295 = ~n_3293 & ~n_3294;
assign n_3296 = ~n_3292 &  n_3295;
assign n_3297 = ~n_3290 &  n_3296;
assign n_3298 = ~n_3291 & ~n_3297;
assign n_3299 = ~x_1746 &  n_3288;
assign n_3300 =  n_3247 &  n_3280;
assign n_3301 = ~n_3241 & ~n_3256;
assign n_3302 = ~n_3294 &  n_3301;
assign n_3303 = ~n_3300 &  n_3302;
assign n_3304 = ~n_3290 &  n_3303;
assign n_3305 = ~n_3299 & ~n_3304;
assign n_3306 = ~n_3298 & ~n_3305;
assign n_3307 =  n_3286 &  n_3306;
assign n_3308 = ~n_1192 & ~n_3307;
assign n_3309 =  x_1917 &  n_3308;
assign n_3310 =  x_450 &  n_3307;
assign n_3311 = ~n_3309 & ~n_3310;
assign n_3312 =  x_1917 & ~n_3311;
assign n_3313 = ~x_1917 &  n_3311;
assign n_3314 = ~n_3312 & ~n_3313;
assign n_3315 =  x_1916 & ~n_1761;
assign n_3316 =  i_160 &  n_1751;
assign n_3317 =  n_1761 &  n_3316;
assign n_3318 = ~n_3315 & ~n_3317;
assign n_3319 =  x_1916 & ~n_3318;
assign n_3320 = ~x_1916 &  n_3318;
assign n_3321 = ~n_3319 & ~n_3320;
assign n_3322 =  x_1915 & ~n_1770;
assign n_3323 =  n_1770 &  n_3316;
assign n_3324 = ~n_3322 & ~n_3323;
assign n_3325 =  x_1915 & ~n_3324;
assign n_3326 = ~x_1915 &  n_3324;
assign n_3327 = ~n_3325 & ~n_3326;
assign n_3328 =  x_1914 & ~n_1778;
assign n_3329 =  n_1778 &  n_3316;
assign n_3330 = ~n_3328 & ~n_3329;
assign n_3331 =  x_1914 & ~n_3330;
assign n_3332 = ~x_1914 &  n_3330;
assign n_3333 = ~n_3331 & ~n_3332;
assign n_3334 =  x_1913 & ~n_1785;
assign n_3335 =  n_1785 &  n_3316;
assign n_3336 = ~n_3334 & ~n_3335;
assign n_3337 =  x_1913 & ~n_3336;
assign n_3338 = ~x_1913 &  n_3336;
assign n_3339 = ~n_3337 & ~n_3338;
assign n_3340 =  x_1912 & ~n_1792;
assign n_3341 =  n_1792 &  n_3316;
assign n_3342 = ~n_3340 & ~n_3341;
assign n_3343 =  x_1912 & ~n_3342;
assign n_3344 = ~x_1912 &  n_3342;
assign n_3345 = ~n_3343 & ~n_3344;
assign n_3346 =  x_1911 & ~n_1799;
assign n_3347 =  n_1799 &  n_3316;
assign n_3348 = ~n_3346 & ~n_3347;
assign n_3349 =  x_1911 & ~n_3348;
assign n_3350 = ~x_1911 &  n_3348;
assign n_3351 = ~n_3349 & ~n_3350;
assign n_3352 =  x_1910 & ~n_1806;
assign n_3353 =  n_1806 &  n_3316;
assign n_3354 = ~n_3352 & ~n_3353;
assign n_3355 =  x_1910 & ~n_3354;
assign n_3356 = ~x_1910 &  n_3354;
assign n_3357 = ~n_3355 & ~n_3356;
assign n_3358 =  n_1750 & ~n_3316;
assign n_3359 = ~x_1909 & ~n_1750;
assign n_3360 = ~n_3358 & ~n_3359;
assign n_3361 =  x_1909 &  n_3360;
assign n_3362 = ~x_1909 & ~n_3360;
assign n_3363 = ~n_3361 & ~n_3362;
assign n_3364 =  x_1908 &  n_3308;
assign n_3365 = ~x_446 &  n_3307;
assign n_3366 = ~n_3364 & ~n_3365;
assign n_3367 =  x_1908 & ~n_3366;
assign n_3368 = ~x_1908 &  n_3366;
assign n_3369 = ~n_3367 & ~n_3368;
assign n_3370 =  x_1907 & ~n_1761;
assign n_3371 =  i_159 &  n_1751;
assign n_3372 =  n_1761 &  n_3371;
assign n_3373 = ~n_3370 & ~n_3372;
assign n_3374 =  x_1907 & ~n_3373;
assign n_3375 = ~x_1907 &  n_3373;
assign n_3376 = ~n_3374 & ~n_3375;
assign n_3377 =  x_1906 & ~n_1770;
assign n_3378 =  n_1770 &  n_3371;
assign n_3379 = ~n_3377 & ~n_3378;
assign n_3380 =  x_1906 & ~n_3379;
assign n_3381 = ~x_1906 &  n_3379;
assign n_3382 = ~n_3380 & ~n_3381;
assign n_3383 =  x_1905 & ~n_1778;
assign n_3384 =  n_1778 &  n_3371;
assign n_3385 = ~n_3383 & ~n_3384;
assign n_3386 =  x_1905 & ~n_3385;
assign n_3387 = ~x_1905 &  n_3385;
assign n_3388 = ~n_3386 & ~n_3387;
assign n_3389 =  x_1904 & ~n_1785;
assign n_3390 =  n_1785 &  n_3371;
assign n_3391 = ~n_3389 & ~n_3390;
assign n_3392 =  x_1904 & ~n_3391;
assign n_3393 = ~x_1904 &  n_3391;
assign n_3394 = ~n_3392 & ~n_3393;
assign n_3395 =  x_1903 & ~n_1792;
assign n_3396 =  n_1792 &  n_3371;
assign n_3397 = ~n_3395 & ~n_3396;
assign n_3398 =  x_1903 & ~n_3397;
assign n_3399 = ~x_1903 &  n_3397;
assign n_3400 = ~n_3398 & ~n_3399;
assign n_3401 =  x_1902 & ~n_1799;
assign n_3402 =  n_1799 &  n_3371;
assign n_3403 = ~n_3401 & ~n_3402;
assign n_3404 =  x_1902 & ~n_3403;
assign n_3405 = ~x_1902 &  n_3403;
assign n_3406 = ~n_3404 & ~n_3405;
assign n_3407 =  x_1901 & ~n_1806;
assign n_3408 =  n_1806 &  n_3371;
assign n_3409 = ~n_3407 & ~n_3408;
assign n_3410 =  x_1901 & ~n_3409;
assign n_3411 = ~x_1901 &  n_3409;
assign n_3412 = ~n_3410 & ~n_3411;
assign n_3413 =  n_1750 & ~n_3371;
assign n_3414 = ~x_1900 & ~n_1750;
assign n_3415 = ~n_3413 & ~n_3414;
assign n_3416 =  x_1900 &  n_3415;
assign n_3417 = ~x_1900 & ~n_3415;
assign n_3418 = ~n_3416 & ~n_3417;
assign n_3419 =  x_1899 &  n_3308;
assign n_3420 =  x_449 &  n_3307;
assign n_3421 = ~n_3419 & ~n_3420;
assign n_3422 =  x_1899 & ~n_3421;
assign n_3423 = ~x_1899 &  n_3421;
assign n_3424 = ~n_3422 & ~n_3423;
assign n_3425 =  x_1898 & ~n_1761;
assign n_3426 =  i_158 &  n_1751;
assign n_3427 =  n_1761 &  n_3426;
assign n_3428 = ~n_3425 & ~n_3427;
assign n_3429 =  x_1898 & ~n_3428;
assign n_3430 = ~x_1898 &  n_3428;
assign n_3431 = ~n_3429 & ~n_3430;
assign n_3432 =  x_1897 & ~n_1770;
assign n_3433 =  n_1770 &  n_3426;
assign n_3434 = ~n_3432 & ~n_3433;
assign n_3435 =  x_1897 & ~n_3434;
assign n_3436 = ~x_1897 &  n_3434;
assign n_3437 = ~n_3435 & ~n_3436;
assign n_3438 =  x_1896 & ~n_1778;
assign n_3439 =  n_1778 &  n_3426;
assign n_3440 = ~n_3438 & ~n_3439;
assign n_3441 =  x_1896 & ~n_3440;
assign n_3442 = ~x_1896 &  n_3440;
assign n_3443 = ~n_3441 & ~n_3442;
assign n_3444 =  x_1895 & ~n_1785;
assign n_3445 =  n_1785 &  n_3426;
assign n_3446 = ~n_3444 & ~n_3445;
assign n_3447 =  x_1895 & ~n_3446;
assign n_3448 = ~x_1895 &  n_3446;
assign n_3449 = ~n_3447 & ~n_3448;
assign n_3450 =  x_1894 & ~n_1792;
assign n_3451 =  n_1792 &  n_3426;
assign n_3452 = ~n_3450 & ~n_3451;
assign n_3453 =  x_1894 & ~n_3452;
assign n_3454 = ~x_1894 &  n_3452;
assign n_3455 = ~n_3453 & ~n_3454;
assign n_3456 =  x_1893 & ~n_1799;
assign n_3457 =  n_1799 &  n_3426;
assign n_3458 = ~n_3456 & ~n_3457;
assign n_3459 =  x_1893 & ~n_3458;
assign n_3460 = ~x_1893 &  n_3458;
assign n_3461 = ~n_3459 & ~n_3460;
assign n_3462 =  x_1892 & ~n_1806;
assign n_3463 =  n_1806 &  n_3426;
assign n_3464 = ~n_3462 & ~n_3463;
assign n_3465 =  x_1892 & ~n_3464;
assign n_3466 = ~x_1892 &  n_3464;
assign n_3467 = ~n_3465 & ~n_3466;
assign n_3468 =  n_1750 & ~n_3426;
assign n_3469 = ~x_1891 & ~n_1750;
assign n_3470 = ~n_3468 & ~n_3469;
assign n_3471 =  x_1891 &  n_3470;
assign n_3472 = ~x_1891 & ~n_3470;
assign n_3473 = ~n_3471 & ~n_3472;
assign n_3474 =  x_1890 &  n_3308;
assign n_3475 = ~x_445 &  n_3307;
assign n_3476 = ~n_3474 & ~n_3475;
assign n_3477 =  x_1890 & ~n_3476;
assign n_3478 = ~x_1890 &  n_3476;
assign n_3479 = ~n_3477 & ~n_3478;
assign n_3480 =  x_1889 & ~n_1761;
assign n_3481 =  i_157 &  n_1751;
assign n_3482 =  n_1761 &  n_3481;
assign n_3483 = ~n_3480 & ~n_3482;
assign n_3484 =  x_1889 & ~n_3483;
assign n_3485 = ~x_1889 &  n_3483;
assign n_3486 = ~n_3484 & ~n_3485;
assign n_3487 =  x_1888 & ~n_1770;
assign n_3488 =  n_1770 &  n_3481;
assign n_3489 = ~n_3487 & ~n_3488;
assign n_3490 =  x_1888 & ~n_3489;
assign n_3491 = ~x_1888 &  n_3489;
assign n_3492 = ~n_3490 & ~n_3491;
assign n_3493 =  x_1887 & ~n_1778;
assign n_3494 =  n_1778 &  n_3481;
assign n_3495 = ~n_3493 & ~n_3494;
assign n_3496 =  x_1887 & ~n_3495;
assign n_3497 = ~x_1887 &  n_3495;
assign n_3498 = ~n_3496 & ~n_3497;
assign n_3499 =  x_1886 & ~n_1785;
assign n_3500 =  n_1785 &  n_3481;
assign n_3501 = ~n_3499 & ~n_3500;
assign n_3502 =  x_1886 & ~n_3501;
assign n_3503 = ~x_1886 &  n_3501;
assign n_3504 = ~n_3502 & ~n_3503;
assign n_3505 =  x_1885 & ~n_1792;
assign n_3506 =  n_1792 &  n_3481;
assign n_3507 = ~n_3505 & ~n_3506;
assign n_3508 =  x_1885 & ~n_3507;
assign n_3509 = ~x_1885 &  n_3507;
assign n_3510 = ~n_3508 & ~n_3509;
assign n_3511 =  x_1884 & ~n_1799;
assign n_3512 =  n_1799 &  n_3481;
assign n_3513 = ~n_3511 & ~n_3512;
assign n_3514 =  x_1884 & ~n_3513;
assign n_3515 = ~x_1884 &  n_3513;
assign n_3516 = ~n_3514 & ~n_3515;
assign n_3517 =  n_1391 &  n_1385;
assign n_3518 =  n_1379 &  n_1373;
assign n_3519 =  n_3517 &  n_3518;
assign n_3520 =  n_1415 &  n_1409;
assign n_3521 =  n_1403 &  n_1397;
assign n_3522 =  n_3520 &  n_3521;
assign n_3523 =  n_3519 &  n_3522;
assign n_3524 =  n_1343 &  n_1337;
assign n_3525 =  x_3105 &  n_1325;
assign n_3526 = ~x_3106 &  n_1329;
assign n_3527 = ~n_3525 & ~n_3526;
assign n_3528 =  n_1331 &  n_3527;
assign n_3529 =  n_3524 &  n_3528;
assign n_3530 =  n_1367 &  n_1361;
assign n_3531 =  n_1355 &  n_1349;
assign n_3532 =  n_3530 &  n_3531;
assign n_3533 =  n_3529 &  n_3532;
assign n_3534 =  n_3523 &  n_3533;
assign n_3535 =  n_1487 &  n_1481;
assign n_3536 =  n_1475 &  n_1469;
assign n_3537 =  n_3535 &  n_3536;
assign n_3538 = ~n_1732 &  n_1505;
assign n_3539 =  n_1499 &  n_1493;
assign n_3540 =  n_3538 &  n_3539;
assign n_3541 =  n_3537 &  n_3540;
assign n_3542 =  n_1439 &  n_1433;
assign n_3543 =  n_1427 &  n_1421;
assign n_3544 =  n_3542 &  n_3543;
assign n_3545 =  n_1463 &  n_1457;
assign n_3546 =  n_1451 &  n_1445;
assign n_3547 =  n_3545 &  n_3546;
assign n_3548 =  n_3544 &  n_3547;
assign n_3549 =  n_3541 &  n_3548;
assign n_3550 =  n_3534 &  n_3549;
assign n_3551 =  x_3239 &  n_3550;
assign n_3552 = ~x_3239 & ~n_3550;
assign n_3553 = ~n_3551 & ~n_3552;
assign n_3554 = ~x_2435 & ~x_2437;
assign n_3555 = ~x_2436 &  n_3554;
assign n_3556 =  x_2435 & ~x_2436;
assign n_3557 = ~x_2437 &  n_3556;
assign n_3558 = ~x_2439 & ~n_3557;
assign n_3559 = ~x_1761 & ~x_1768;
assign n_3560 = ~x_1768 &  x_2440;
assign n_3561 = ~n_3559 & ~n_3560;
assign n_3562 =  i_219 & ~i_220;
assign n_3563 =  x_295 &  n_3562;
assign n_3564 = ~i_218 &  n_3563;
assign n_3565 =  i_217 &  x_295;
assign n_3566 =  x_1768 &  n_3565;
assign n_3567 =  n_3564 & ~n_3566;
assign n_3568 =  n_3561 & ~n_3567;
assign n_3569 =  i_220 &  x_295;
assign n_3570 = ~n_3563 & ~n_3569;
assign n_3571 = ~n_3263 &  n_3570;
assign n_3572 = ~i_223 & ~i_224;
assign n_3573 = ~n_3563 &  n_3572;
assign n_3574 = ~n_3571 & ~n_3573;
assign n_3575 = ~n_3568 &  n_3574;
assign n_3576 = ~n_3558 &  n_3575;
assign n_3577 = ~x_2436 &  x_2437;
assign n_3578 =  x_2436 & ~x_2441;
assign n_3579 =  n_3578 &  n_3554;
assign n_3580 = ~n_3577 & ~n_3579;
assign n_3581 =  n_3571 & ~n_3572;
assign n_3582 = ~n_3580 & ~n_3581;
assign n_3583 = ~x_2438 & ~n_3575;
assign n_3584 =  n_3582 &  n_3583;
assign n_3585 =  n_3558 & ~n_3584;
assign n_3586 =  x_2442 &  n_3568;
assign n_3587 = ~x_2435 &  x_2441;
assign n_3588 = ~n_3586 &  n_3587;
assign n_3589 =  x_2435 &  x_2437;
assign n_3590 =  n_3578 & ~n_3554;
assign n_3591 = ~n_3589 &  n_3590;
assign n_3592 =  n_3567 &  n_3591;
assign n_3593 = ~x_2438 & ~n_3580;
assign n_3594 =  n_3561 & ~n_3593;
assign n_3595 = ~n_3592 &  n_3594;
assign n_3596 = ~n_3588 &  n_3595;
assign n_3597 =  n_3585 & ~n_3596;
assign n_3598 = ~n_3576 & ~n_3597;
assign n_3599 = ~n_3555 &  n_3598;
assign n_3600 = ~n_3561 & ~n_3567;
assign n_3601 = ~n_3571 &  n_3600;
assign n_3602 =  n_3593 & ~n_3601;
assign n_3603 = ~x_2442 &  n_3592;
assign n_3604 = ~n_3561 & ~n_3603;
assign n_3605 = ~n_3602 &  n_3604;
assign n_3606 =  n_3585 &  n_3605;
assign n_3607 = ~n_3581 & ~n_3601;
assign n_3608 = ~n_3558 & ~n_3573;
assign n_3609 = ~n_3607 &  n_3608;
assign n_3610 = ~n_3555 & ~n_3609;
assign n_3611 = ~n_3606 &  n_3610;
assign n_3612 = ~n_3599 & ~n_3611;
assign n_3613 =  x_2443 & ~n_3612;
assign n_3614 =  n_3555 & ~n_3560;
assign n_3615 = ~n_3560 & ~n_3586;
assign n_3616 = ~n_3564 &  n_3615;
assign n_3617 =  n_3564 &  n_3566;
assign n_3618 = ~n_3616 & ~n_3617;
assign n_3619 =  n_3574 & ~n_3618;
assign n_3620 = ~n_3557 & ~n_3582;
assign n_3621 = ~n_3619 & ~n_3620;
assign n_3622 = ~x_2442 & ~n_3618;
assign n_3623 =  x_2442 &  n_3559;
assign n_3624 =  n_3591 & ~n_3623;
assign n_3625 = ~n_3622 &  n_3624;
assign n_3626 =  n_3578 &  n_3589;
assign n_3627 = ~n_3559 &  n_3626;
assign n_3628 =  n_3615 & ~n_3627;
assign n_3629 = ~n_3625 &  n_3628;
assign n_3630 = ~n_3556 & ~n_3579;
assign n_3631 = ~n_3629 &  n_3630;
assign n_3632 = ~n_3621 & ~n_3631;
assign n_3633 = ~n_3614 & ~n_3632;
assign n_3634 =  n_3633 &  n_3612;
assign n_3635 =  i_151 & ~i_152;
assign n_3636 =  x_295 &  n_3635;
assign n_3637 =  x_1758 &  n_3636;
assign n_3638 =  x_1489 &  n_3637;
assign n_3639 =  n_3634 & ~n_3638;
assign n_3640 = ~n_3613 & ~n_3639;
assign n_3641 =  x_2444 & ~n_3634;
assign n_3642 =  x_1761 & ~x_1768;
assign n_3643 = ~x_2366 &  n_3642;
assign n_3644 =  x_309 & ~x_310;
assign n_3645 =  x_1768 &  n_3644;
assign n_3646 =  x_1770 & ~x_2400;
assign n_3647 =  n_3645 &  n_3646;
assign n_3648 = ~n_3643 & ~n_3647;
assign n_3649 =  n_3634 & ~n_3648;
assign n_3650 = ~n_3641 & ~n_3649;
assign n_3651 = ~n_3640 & ~n_3650;
assign n_3652 =  x_2445 & ~n_3634;
assign n_3653 =  x_1770 & ~x_2401;
assign n_3654 =  n_3645 & ~n_3653;
assign n_3655 =  x_2367 &  n_3642;
assign n_3656 = ~n_3654 & ~n_3655;
assign n_3657 =  n_3634 & ~n_3656;
assign n_3658 = ~n_3652 & ~n_3657;
assign n_3659 =  x_2446 & ~n_3634;
assign n_3660 =  x_1770 & ~x_2402;
assign n_3661 =  n_3645 & ~n_3660;
assign n_3662 =  x_2368 &  n_3642;
assign n_3663 = ~n_3661 & ~n_3662;
assign n_3664 =  n_3634 & ~n_3663;
assign n_3665 = ~n_3659 & ~n_3664;
assign n_3666 =  n_3658 &  n_3665;
assign n_3667 =  n_3651 &  n_3666;
assign n_3668 = ~x_1761 &  x_1768;
assign n_3669 =  x_2442 & ~n_3612;
assign n_3670 = ~n_3668 & ~n_3669;
assign n_3671 =  n_3617 &  n_3670;
assign n_3672 =  n_3667 &  n_3671;
assign n_3673 = ~n_1325 &  n_1327;
assign n_3674 =  x_1721 &  x_1722;
assign n_3675 =  x_308 &  n_3674;
assign n_3676 =  i_12 &  x_295;
assign n_3677 = ~x_1721 &  x_1722;
assign n_3678 = ~n_3676 &  n_3677;
assign n_3679 =  i_11 &  x_295;
assign n_3680 =  x_1724 & ~n_3679;
assign n_3681 =  x_1723 &  n_3680;
assign n_3682 =  n_3678 &  n_3681;
assign n_3683 = ~n_3675 & ~n_3682;
assign n_3684 =  x_1729 & ~n_3683;
assign n_3685 = ~n_3676 &  n_3679;
assign n_3686 = ~x_1727 & ~x_1728;
assign n_3687 =  x_308 &  n_3686;
assign n_3688 = ~n_3685 &  n_3687;
assign n_3689 = ~n_3684 & ~n_3688;
assign n_3690 = ~n_3673 & ~n_3689;
assign n_3691 =  x_1721 & ~x_1722;
assign n_3692 =  x_1723 &  x_1724;
assign n_3693 =  n_3691 &  n_3692;
assign n_3694 =  n_1328 &  n_3693;
assign n_3695 = ~n_3675 & ~n_3694;
assign n_3696 =  x_1726 & ~n_3685;
assign n_3697 = ~n_3695 &  n_3696;
assign n_3698 = ~n_3690 & ~n_3697;
assign n_3699 = ~x_1725 & ~n_3698;
assign n_3700 = ~x_308 &  n_1257;
assign n_3701 =  x_3153 &  n_3700;
assign n_3702 =  x_3153 &  n_1258;
assign n_3703 = ~x_3154 &  n_3702;
assign n_3704 = ~n_3701 & ~n_3703;
assign n_3705 = ~n_3699 & ~n_3704;
assign n_3706 = ~x_3153 & ~n_3700;
assign n_3707 =  n_3706 &  n_3699;
assign n_3708 = ~n_3705 & ~n_3707;
assign n_3709 = ~n_3672 &  n_3708;
assign n_3710 =  x_3238 & ~n_3709;
assign n_3711 = ~x_3238 &  n_3709;
assign n_3712 = ~n_3710 & ~n_3711;
assign n_3713 =  x_2449 & ~n_3634;
assign n_3714 = ~n_3639 & ~n_3713;
assign n_3715 =  x_310 &  n_3637;
assign n_3716 =  n_3634 &  n_3715;
assign n_3717 = ~x_1755 & ~n_3636;
assign n_3718 =  x_1757 & ~n_3717;
assign n_3719 =  x_309 &  x_1758;
assign n_3720 =  n_3718 &  n_3719;
assign n_3721 =  n_3716 &  n_3720;
assign n_3722 =  n_3714 &  n_3721;
assign n_3723 =  x_3237 &  n_3722;
assign n_3724 = ~x_3237 & ~n_3722;
assign n_3725 = ~n_3723 & ~n_3724;
assign n_3726 =  x_227 &  n_3673;
assign n_3727 =  x_3107 &  n_3726;
assign n_3728 =  x_3108 &  x_3109;
assign n_3729 =  x_3110 &  n_3728;
assign n_3730 =  x_3111 &  n_3729;
assign n_3731 =  x_3112 &  n_3730;
assign n_3732 =  x_3113 &  n_3731;
assign n_3733 =  x_3114 &  n_3732;
assign n_3734 =  x_3115 &  n_3733;
assign n_3735 =  x_3116 &  n_3734;
assign n_3736 =  x_3117 &  n_3735;
assign n_3737 =  x_3118 &  n_3736;
assign n_3738 =  x_3119 &  n_3737;
assign n_3739 =  x_3120 &  n_3738;
assign n_3740 =  x_3121 &  n_3739;
assign n_3741 =  x_3122 &  n_3740;
assign n_3742 =  x_3123 &  n_3741;
assign n_3743 =  x_3124 &  n_3742;
assign n_3744 =  x_3125 &  n_3743;
assign n_3745 =  x_3126 &  n_3744;
assign n_3746 =  x_3127 &  n_3745;
assign n_3747 =  x_3128 &  n_3746;
assign n_3748 =  x_3129 &  n_3747;
assign n_3749 =  x_3130 &  n_3748;
assign n_3750 =  x_3131 &  n_3749;
assign n_3751 =  x_3132 &  n_3750;
assign n_3752 =  x_3133 &  n_3751;
assign n_3753 =  x_3134 &  n_3752;
assign n_3754 =  x_3135 &  n_3753;
assign n_3755 =  x_3136 &  n_3754;
assign n_3756 =  x_3137 &  n_3755;
assign n_3757 =  x_3138 &  n_3756;
assign n_3758 =  n_3727 & ~n_3757;
assign n_3759 = ~n_1325 & ~n_3758;
assign n_3760 =  x_3139 & ~n_3759;
assign n_3761 = ~x_3139 &  n_3727;
assign n_3762 =  n_3757 &  n_3761;
assign n_3763 = ~n_3760 & ~n_3762;
assign n_3764 =  x_3138 & ~n_3759;
assign n_3765 =  n_3756 &  n_3758;
assign n_3766 = ~n_3764 & ~n_3765;
assign n_3767 =  x_3137 &  n_1325;
assign n_3768 = ~x_3137 & ~n_3755;
assign n_3769 =  n_3727 & ~n_3756;
assign n_3770 = ~n_3768 &  n_3769;
assign n_3771 = ~n_3767 & ~n_3770;
assign n_3772 =  x_3136 &  n_1325;
assign n_3773 = ~x_3136 & ~n_3754;
assign n_3774 =  n_3727 & ~n_3755;
assign n_3775 = ~n_3773 &  n_3774;
assign n_3776 = ~n_3772 & ~n_3775;
assign n_3777 =  x_3135 &  n_1325;
assign n_3778 = ~x_3135 & ~n_3753;
assign n_3779 =  n_3727 & ~n_3754;
assign n_3780 = ~n_3778 &  n_3779;
assign n_3781 = ~n_3777 & ~n_3780;
assign n_3782 =  x_3134 &  n_1325;
assign n_3783 = ~x_3134 & ~n_3752;
assign n_3784 =  n_3727 & ~n_3753;
assign n_3785 = ~n_3783 &  n_3784;
assign n_3786 = ~n_3782 & ~n_3785;
assign n_3787 =  x_3133 &  n_1325;
assign n_3788 = ~x_3133 & ~n_3751;
assign n_3789 =  n_3727 & ~n_3752;
assign n_3790 = ~n_3788 &  n_3789;
assign n_3791 = ~n_3787 & ~n_3790;
assign n_3792 =  x_3132 &  n_1325;
assign n_3793 = ~x_3132 & ~n_3750;
assign n_3794 =  n_3727 & ~n_3751;
assign n_3795 = ~n_3793 &  n_3794;
assign n_3796 = ~n_3792 & ~n_3795;
assign n_3797 =  x_3131 &  n_1325;
assign n_3798 = ~x_3131 & ~n_3749;
assign n_3799 =  n_3727 & ~n_3750;
assign n_3800 = ~n_3798 &  n_3799;
assign n_3801 = ~n_3797 & ~n_3800;
assign n_3802 =  x_3130 &  n_1325;
assign n_3803 = ~x_3130 & ~n_3748;
assign n_3804 =  n_3727 & ~n_3749;
assign n_3805 = ~n_3803 &  n_3804;
assign n_3806 = ~n_3802 & ~n_3805;
assign n_3807 =  x_3129 &  n_1325;
assign n_3808 = ~x_3129 & ~n_3747;
assign n_3809 =  n_3727 & ~n_3748;
assign n_3810 = ~n_3808 &  n_3809;
assign n_3811 = ~n_3807 & ~n_3810;
assign n_3812 =  x_3128 &  n_1325;
assign n_3813 = ~x_3128 & ~n_3746;
assign n_3814 =  n_3727 & ~n_3747;
assign n_3815 = ~n_3813 &  n_3814;
assign n_3816 = ~n_3812 & ~n_3815;
assign n_3817 =  x_3127 &  n_1325;
assign n_3818 = ~x_3127 & ~n_3745;
assign n_3819 =  n_3727 & ~n_3746;
assign n_3820 = ~n_3818 &  n_3819;
assign n_3821 = ~n_3817 & ~n_3820;
assign n_3822 =  x_3126 &  n_1325;
assign n_3823 = ~x_3126 & ~n_3744;
assign n_3824 =  n_3727 & ~n_3745;
assign n_3825 = ~n_3823 &  n_3824;
assign n_3826 = ~n_3822 & ~n_3825;
assign n_3827 =  x_3125 &  n_1325;
assign n_3828 = ~x_3125 & ~n_3743;
assign n_3829 =  n_3727 & ~n_3744;
assign n_3830 = ~n_3828 &  n_3829;
assign n_3831 = ~n_3827 & ~n_3830;
assign n_3832 =  x_3124 &  n_1325;
assign n_3833 = ~x_3124 & ~n_3742;
assign n_3834 =  n_3727 & ~n_3743;
assign n_3835 = ~n_3833 &  n_3834;
assign n_3836 = ~n_3832 & ~n_3835;
assign n_3837 =  x_3123 &  n_1325;
assign n_3838 = ~x_3123 & ~n_3741;
assign n_3839 =  n_3727 & ~n_3742;
assign n_3840 = ~n_3838 &  n_3839;
assign n_3841 = ~n_3837 & ~n_3840;
assign n_3842 =  x_3122 &  n_1325;
assign n_3843 = ~x_3122 & ~n_3740;
assign n_3844 =  n_3727 & ~n_3741;
assign n_3845 = ~n_3843 &  n_3844;
assign n_3846 = ~n_3842 & ~n_3845;
assign n_3847 =  x_3121 &  n_1325;
assign n_3848 = ~x_3121 & ~n_3739;
assign n_3849 =  n_3727 & ~n_3740;
assign n_3850 = ~n_3848 &  n_3849;
assign n_3851 = ~n_3847 & ~n_3850;
assign n_3852 =  x_3120 &  n_1325;
assign n_3853 = ~x_3120 & ~n_3738;
assign n_3854 =  n_3727 & ~n_3739;
assign n_3855 = ~n_3853 &  n_3854;
assign n_3856 = ~n_3852 & ~n_3855;
assign n_3857 =  x_3119 &  n_1325;
assign n_3858 = ~x_3119 & ~n_3737;
assign n_3859 =  n_3727 & ~n_3738;
assign n_3860 = ~n_3858 &  n_3859;
assign n_3861 = ~n_3857 & ~n_3860;
assign n_3862 =  x_3118 &  n_1325;
assign n_3863 = ~x_3118 & ~n_3736;
assign n_3864 =  n_3727 & ~n_3737;
assign n_3865 = ~n_3863 &  n_3864;
assign n_3866 = ~n_3862 & ~n_3865;
assign n_3867 =  x_3117 &  n_1325;
assign n_3868 = ~x_3117 & ~n_3735;
assign n_3869 =  n_3727 & ~n_3736;
assign n_3870 = ~n_3868 &  n_3869;
assign n_3871 = ~n_3867 & ~n_3870;
assign n_3872 =  x_3116 &  n_1325;
assign n_3873 = ~x_3116 & ~n_3734;
assign n_3874 =  n_3727 & ~n_3735;
assign n_3875 = ~n_3873 &  n_3874;
assign n_3876 = ~n_3872 & ~n_3875;
assign n_3877 =  x_3115 &  n_1325;
assign n_3878 = ~x_3115 & ~n_3733;
assign n_3879 =  n_3727 & ~n_3878;
assign n_3880 = ~n_3734 &  n_3879;
assign n_3881 = ~n_3877 & ~n_3880;
assign n_3882 =  x_3114 &  n_1325;
assign n_3883 = ~x_3114 & ~n_3732;
assign n_3884 =  n_3727 & ~n_3733;
assign n_3885 = ~n_3883 &  n_3884;
assign n_3886 = ~n_3882 & ~n_3885;
assign n_3887 =  x_3113 &  n_1325;
assign n_3888 = ~x_3113 & ~n_3731;
assign n_3889 =  n_3727 & ~n_3732;
assign n_3890 = ~n_3888 &  n_3889;
assign n_3891 = ~n_3887 & ~n_3890;
assign n_3892 =  x_3112 &  n_1325;
assign n_3893 = ~x_3112 & ~n_3730;
assign n_3894 =  n_3727 & ~n_3893;
assign n_3895 = ~n_3731 &  n_3894;
assign n_3896 = ~n_3892 & ~n_3895;
assign n_3897 =  x_3111 &  n_1325;
assign n_3898 = ~x_3111 & ~n_3729;
assign n_3899 = ~n_3898 & ~n_3730;
assign n_3900 =  n_3727 &  n_3899;
assign n_3901 = ~n_3897 & ~n_3900;
assign n_3902 =  x_3110 &  n_1325;
assign n_3903 = ~x_3110 & ~n_3728;
assign n_3904 = ~n_3903 & ~n_3729;
assign n_3905 =  n_3727 &  n_3904;
assign n_3906 = ~n_3902 & ~n_3905;
assign n_3907 =  x_3109 &  n_1325;
assign n_3908 = ~x_3108 & ~x_3109;
assign n_3909 = ~n_3908 & ~n_3728;
assign n_3910 =  n_3726 &  n_3909;
assign n_3911 = ~n_3907 & ~n_3910;
assign n_3912 =  n_1732 &  n_3911;
assign n_3913 =  n_3906 &  n_3912;
assign n_3914 =  n_3901 &  n_3913;
assign n_3915 =  n_3896 &  n_3914;
assign n_3916 =  n_3891 &  n_3915;
assign n_3917 =  n_3886 &  n_3916;
assign n_3918 =  n_3881 &  n_3917;
assign n_3919 =  n_3876 &  n_3918;
assign n_3920 =  n_3871 &  n_3919;
assign n_3921 =  n_3866 &  n_3920;
assign n_3922 =  n_3861 &  n_3921;
assign n_3923 =  n_3856 &  n_3922;
assign n_3924 =  n_3851 &  n_3923;
assign n_3925 =  n_3846 &  n_3924;
assign n_3926 =  n_3841 &  n_3925;
assign n_3927 =  n_3836 &  n_3926;
assign n_3928 =  n_3831 &  n_3927;
assign n_3929 =  n_3826 &  n_3928;
assign n_3930 =  n_3821 &  n_3929;
assign n_3931 =  n_3816 &  n_3930;
assign n_3932 =  n_3811 &  n_3931;
assign n_3933 =  n_3806 &  n_3932;
assign n_3934 =  n_3801 &  n_3933;
assign n_3935 =  n_3796 &  n_3934;
assign n_3936 =  n_3791 &  n_3935;
assign n_3937 =  n_3786 &  n_3936;
assign n_3938 =  n_3781 &  n_3937;
assign n_3939 =  n_3776 &  n_3938;
assign n_3940 =  n_3771 &  n_3939;
assign n_3941 =  n_3766 &  n_3940;
assign n_3942 =  n_3763 &  n_3941;
assign n_3943 =  x_3236 &  n_3942;
assign n_3944 = ~x_3236 & ~n_3942;
assign n_3945 = ~n_3943 & ~n_3944;
assign n_3946 =  x_2522 &  n_1522;
assign n_3947 = ~x_2523 &  n_1526;
assign n_3948 = ~n_3946 & ~n_3947;
assign n_3949 =  n_1534 &  n_1528;
assign n_3950 =  n_3948 &  n_3949;
assign n_3951 =  n_1558 &  n_1552;
assign n_3952 =  n_1546 &  n_1540;
assign n_3953 =  n_3951 &  n_3952;
assign n_3954 =  n_1582 &  n_1576;
assign n_3955 =  n_1570 &  n_1564;
assign n_3956 =  n_3954 &  n_3955;
assign n_3957 =  n_3953 &  n_3956;
assign n_3958 =  n_3950 &  n_3957;
assign n_3959 = ~n_1708 &  n_1702;
assign n_3960 =  n_1741 &  n_1696;
assign n_3961 =  n_1690 &  n_1684;
assign n_3962 =  n_3960 &  n_3961;
assign n_3963 =  n_3959 &  n_3962;
assign n_3964 =  n_1654 &  n_1648;
assign n_3965 =  n_1642 &  n_1636;
assign n_3966 =  n_3964 &  n_3965;
assign n_3967 =  n_1678 &  n_1672;
assign n_3968 =  n_1666 &  n_1660;
assign n_3969 =  n_3967 &  n_3968;
assign n_3970 =  n_3966 &  n_3969;
assign n_3971 =  n_1606 &  n_1600;
assign n_3972 =  n_1594 &  n_1588;
assign n_3973 =  n_3971 &  n_3972;
assign n_3974 =  n_1630 &  n_1624;
assign n_3975 =  n_1618 &  n_1612;
assign n_3976 =  n_3974 &  n_3975;
assign n_3977 =  n_3973 &  n_3976;
assign n_3978 =  n_3970 &  n_3977;
assign n_3979 =  n_3963 &  n_3978;
assign n_3980 =  n_3958 &  n_3979;
assign n_3981 =  x_3235 &  n_3980;
assign n_3982 = ~x_3235 & ~n_3980;
assign n_3983 = ~n_3981 & ~n_3982;
assign n_3984 = ~n_3263 & ~n_3667;
assign n_3985 =  x_3234 & ~n_3984;
assign n_3986 = ~x_3234 &  n_3984;
assign n_3987 = ~n_3985 & ~n_3986;
assign n_3988 =  n_1101 &  n_1041;
assign n_3989 =  n_981 &  n_919;
assign n_3990 =  n_3988 &  n_3989;
assign n_3991 =  n_574 &  n_562;
assign n_3992 =  n_550 &  n_538;
assign n_3993 =  n_3991 &  n_3992;
assign n_3994 =  n_627 & ~n_3993;
assign n_3995 =  n_657 &  n_645;
assign n_3996 =  n_633 &  n_621;
assign n_3997 =  n_3995 &  n_3996;
assign n_3998 = ~n_3994 &  n_3997;
assign n_3999 =  n_676 & ~n_3998;
assign n_4000 =  n_706 &  n_694;
assign n_4001 =  n_682 &  n_670;
assign n_4002 =  n_4000 &  n_4001;
assign n_4003 = ~n_3999 &  n_4002;
assign n_4004 =  n_725 & ~n_4003;
assign n_4005 =  n_755 &  n_743;
assign n_4006 =  n_731 &  n_719;
assign n_4007 =  n_4005 &  n_4006;
assign n_4008 = ~n_4004 &  n_4007;
assign n_4009 =  n_774 & ~n_4008;
assign n_4010 =  n_804 &  n_792;
assign n_4011 =  n_780 &  n_768;
assign n_4012 =  n_4010 &  n_4011;
assign n_4013 = ~n_4009 &  n_4012;
assign n_4014 =  n_823 & ~n_4013;
assign n_4015 =  n_902 &  n_890;
assign n_4016 =  n_878 &  n_866;
assign n_4017 =  n_4015 &  n_4016;
assign n_4018 =  n_853 &  n_841;
assign n_4019 =  n_829 &  n_817;
assign n_4020 =  n_4018 &  n_4019;
assign n_4021 =  n_4017 &  n_4020;
assign n_4022 = ~n_4014 &  n_4021;
assign n_4023 = ~n_872 &  n_4017;
assign n_4024 =  n_951 & ~n_4023;
assign n_4025 = ~n_4022 &  n_4024;
assign n_4026 =  n_3990 & ~n_4025;
assign n_4027 = ~x_3227 & ~n_4026;
assign n_4028 = ~x_3222 & ~x_3224;
assign n_4029 = ~x_3226 & ~x_3228;
assign n_4030 =  n_4028 &  n_4029;
assign n_4031 = ~n_4027 &  n_4030;
assign n_4032 = ~x_3218 & ~n_4031;
assign n_4033 = ~x_3213 & ~x_3215;
assign n_4034 = ~x_3217 & ~x_3219;
assign n_4035 =  n_4033 &  n_4034;
assign n_4036 = ~n_4032 &  n_4035;
assign n_4037 = ~x_3209 & ~n_4036;
assign n_4038 = ~x_3204 & ~x_3206;
assign n_4039 = ~x_3208 & ~x_3210;
assign n_4040 =  n_4038 &  n_4039;
assign n_4041 = ~n_4037 &  n_4040;
assign n_4042 = ~x_3200 & ~n_4041;
assign n_4043 = ~x_3195 & ~x_3197;
assign n_4044 = ~x_3199 & ~x_3201;
assign n_4045 =  n_4043 &  n_4044;
assign n_4046 = ~n_4042 &  n_4045;
assign n_4047 = ~x_3191 & ~n_4046;
assign n_4048 = ~x_3186 & ~x_3188;
assign n_4049 = ~x_3190 & ~x_3192;
assign n_4050 =  n_4048 &  n_4049;
assign n_4051 = ~n_4047 &  n_4050;
assign n_4052 = ~x_3182 & ~n_4051;
assign n_4053 = ~x_3177 & ~x_3179;
assign n_4054 = ~x_3181 & ~x_3183;
assign n_4055 =  n_4053 &  n_4054;
assign n_4056 = ~x_3161 & ~x_3163;
assign n_4057 = ~x_3168 & ~x_3170;
assign n_4058 = ~x_3172 & ~x_3174;
assign n_4059 =  n_4057 &  n_4058;
assign n_4060 =  n_4056 &  n_4059;
assign n_4061 =  n_4055 &  n_4060;
assign n_4062 = ~n_4052 &  n_4061;
assign n_4063 = ~x_3164 & ~n_4062;
assign n_4064 = ~x_3165 & ~n_4063;
assign n_4065 =  n_713 &  n_706;
assign n_4066 = ~x_3159 & ~n_611;
assign n_4067 =  x_3194 &  n_4066;
assign n_4068 =  x_3193 & ~n_4067;
assign n_4069 = ~x_3195 &  n_4068;
assign n_4070 = ~n_4065 & ~n_4069;
assign n_4071 =  x_3212 &  n_4066;
assign n_4072 =  x_3211 & ~n_4071;
assign n_4073 = ~x_3213 &  n_4072;
assign n_4074 =  n_811 &  n_804;
assign n_4075 = ~n_4073 & ~n_4074;
assign n_4076 =  n_4070 &  n_4075;
assign n_4077 =  n_1139 &  n_1101;
assign n_4078 = ~n_823 &  n_817;
assign n_4079 = ~n_896 &  n_890;
assign n_4080 = ~n_4078 & ~n_4079;
assign n_4081 = ~n_847 &  n_841;
assign n_4082 = ~n_798 &  n_792;
assign n_4083 = ~n_4081 & ~n_4082;
assign n_4084 =  n_4080 &  n_4083;
assign n_4085 = ~n_676 &  n_670;
assign n_4086 = ~n_556 &  n_550;
assign n_4087 = ~n_4085 & ~n_4086;
assign n_4088 = ~n_627 &  n_621;
assign n_4089 = ~n_568 &  n_562;
assign n_4090 = ~n_4088 & ~n_4089;
assign n_4091 =  n_4087 &  n_4090;
assign n_4092 = ~n_737 &  n_731;
assign n_4093 = ~n_639 &  n_633;
assign n_4094 = ~n_4092 & ~n_4093;
assign n_4095 = ~n_651 &  n_645;
assign n_4096 = ~n_872 &  n_866;
assign n_4097 = ~n_4095 & ~n_4096;
assign n_4098 =  n_4094 &  n_4097;
assign n_4099 =  n_4091 &  n_4098;
assign n_4100 =  n_4084 &  n_4099;
assign n_4101 = ~n_951 &  n_919;
assign n_4102 = ~n_544 &  n_538;
assign n_4103 =  x_3189 & ~x_3190;
assign n_4104 =  x_3162 & ~x_3163;
assign n_4105 = ~n_4103 & ~n_4104;
assign n_4106 =  x_3173 & ~x_3174;
assign n_4107 =  x_3214 & ~x_3215;
assign n_4108 = ~n_4106 & ~n_4107;
assign n_4109 =  n_4105 &  n_4108;
assign n_4110 =  x_3198 & ~x_3199;
assign n_4111 =  x_3216 & ~x_3217;
assign n_4112 = ~n_4110 & ~n_4111;
assign n_4113 =  x_3225 & ~x_3226;
assign n_4114 =  x_3196 & ~x_3197;
assign n_4115 = ~n_4113 & ~n_4114;
assign n_4116 =  n_4112 &  n_4115;
assign n_4117 =  n_4109 &  n_4116;
assign n_4118 =  x_3182 & ~x_3183;
assign n_4119 =  x_3209 & ~x_3210;
assign n_4120 = ~n_4118 & ~n_4119;
assign n_4121 =  x_3191 & ~x_3192;
assign n_4122 =  x_3169 & ~x_3170;
assign n_4123 = ~n_4121 & ~n_4122;
assign n_4124 =  n_4120 &  n_4123;
assign n_4125 =  x_3171 & ~x_3172;
assign n_4126 =  x_3227 & ~x_3228;
assign n_4127 = ~n_4125 & ~n_4126;
assign n_4128 =  x_3187 & ~x_3188;
assign n_4129 =  x_3218 & ~x_3219;
assign n_4130 = ~n_4128 & ~n_4129;
assign n_4131 =  n_4127 &  n_4130;
assign n_4132 =  n_4124 &  n_4131;
assign n_4133 =  x_3178 & ~x_3179;
assign n_4134 =  x_3200 & ~x_3201;
assign n_4135 =  x_3207 & ~x_3208;
assign n_4136 = ~n_4134 & ~n_4135;
assign n_4137 = ~n_4133 &  n_4136;
assign n_4138 =  x_3205 & ~x_3206;
assign n_4139 =  x_3160 & ~x_3161;
assign n_4140 = ~n_4138 & ~n_4139;
assign n_4141 =  x_3223 & ~x_3224;
assign n_4142 =  x_3180 & ~x_3181;
assign n_4143 = ~n_4141 & ~n_4142;
assign n_4144 =  n_4140 &  n_4143;
assign n_4145 =  n_4137 &  n_4144;
assign n_4146 =  n_4132 &  n_4145;
assign n_4147 =  n_4117 &  n_4146;
assign n_4148 = ~n_4102 &  n_4147;
assign n_4149 = ~n_4101 &  n_4148;
assign n_4150 = ~n_1071 &  n_1041;
assign n_4151 = ~n_1011 &  n_981;
assign n_4152 = ~n_4150 & ~n_4151;
assign n_4153 =  n_4149 &  n_4152;
assign n_4154 = ~n_688 &  n_682;
assign n_4155 = ~n_700 &  n_694;
assign n_4156 = ~n_4154 & ~n_4155;
assign n_4157 = ~n_835 &  n_829;
assign n_4158 = ~n_884 &  n_878;
assign n_4159 = ~n_4157 & ~n_4158;
assign n_4160 =  n_4156 &  n_4159;
assign n_4161 = ~n_749 &  n_743;
assign n_4162 = ~n_786 &  n_780;
assign n_4163 = ~n_4161 & ~n_4162;
assign n_4164 = ~n_725 &  n_719;
assign n_4165 = ~n_774 &  n_768;
assign n_4166 = ~n_4164 & ~n_4165;
assign n_4167 =  n_4163 &  n_4166;
assign n_4168 =  n_4160 &  n_4167;
assign n_4169 =  n_4153 &  n_4168;
assign n_4170 =  n_4100 &  n_4169;
assign n_4171 = ~n_4077 &  n_4170;
assign n_4172 =  n_909 &  n_902;
assign n_4173 =  n_860 &  n_853;
assign n_4174 = ~n_4172 & ~n_4173;
assign n_4175 =  n_4171 &  n_4174;
assign n_4176 =  n_4076 &  n_4175;
assign n_4177 =  x_3185 &  n_4066;
assign n_4178 =  x_3184 & ~n_4177;
assign n_4179 = ~x_3186 &  n_4178;
assign n_4180 =  x_3221 &  n_4066;
assign n_4181 =  x_3220 & ~n_4180;
assign n_4182 = ~x_3222 &  n_4181;
assign n_4183 = ~n_4179 & ~n_4182;
assign n_4184 =  n_664 &  n_657;
assign n_4185 =  n_762 &  n_755;
assign n_4186 = ~n_4184 & ~n_4185;
assign n_4187 =  n_4183 &  n_4186;
assign n_4188 =  x_3167 &  n_4066;
assign n_4189 =  x_3166 & ~n_4188;
assign n_4190 = ~x_3168 &  n_4189;
assign n_4191 =  x_3203 &  n_4066;
assign n_4192 =  x_3202 & ~n_4191;
assign n_4193 = ~x_3204 &  n_4192;
assign n_4194 = ~n_4190 & ~n_4193;
assign n_4195 =  n_615 &  n_574;
assign n_4196 =  x_3176 &  n_4066;
assign n_4197 =  x_3175 & ~n_4196;
assign n_4198 = ~x_3177 &  n_4197;
assign n_4199 = ~n_4195 & ~n_4198;
assign n_4200 =  n_4194 &  n_4199;
assign n_4201 =  n_4187 &  n_4200;
assign n_4202 =  n_4176 &  n_4201;
assign n_4203 = ~n_4064 &  n_4202;
assign n_4204 = ~n_811 & ~n_762;
assign n_4205 = ~n_713 & ~n_664;
assign n_4206 =  n_4204 &  n_4205;
assign n_4207 =  n_1071 &  n_1011;
assign n_4208 =  n_951 &  n_4207;
assign n_4209 =  n_3990 &  n_4208;
assign n_4210 =  n_4021 &  n_4209;
assign n_4211 =  n_4002 &  n_4007;
assign n_4212 =  n_4012 &  n_4211;
assign n_4213 =  n_568 &  n_556;
assign n_4214 =  n_544 &  n_4213;
assign n_4215 =  n_676 &  n_651;
assign n_4216 =  n_639 &  n_627;
assign n_4217 =  n_4215 &  n_4216;
assign n_4218 =  n_4214 &  n_4217;
assign n_4219 =  n_3993 &  n_3997;
assign n_4220 =  n_4218 &  n_4219;
assign n_4221 =  n_872 &  n_847;
assign n_4222 =  n_835 &  n_823;
assign n_4223 =  n_4221 &  n_4222;
assign n_4224 = ~x_3209 & ~x_3214;
assign n_4225 = ~x_3216 & ~x_3218;
assign n_4226 =  n_4224 &  n_4225;
assign n_4227 = ~x_3198 & ~x_3200;
assign n_4228 = ~x_3205 & ~x_3207;
assign n_4229 =  n_4227 &  n_4228;
assign n_4230 =  n_4226 &  n_4229;
assign n_4231 = ~x_3223 & ~x_3225;
assign n_4232 = ~x_3227 &  n_4231;
assign n_4233 =  n_4030 &  n_4232;
assign n_4234 =  n_4230 &  n_4233;
assign n_4235 = ~x_3160 & ~x_3162;
assign n_4236 = ~x_3164 & ~x_3165;
assign n_4237 = ~x_3169 & ~x_3171;
assign n_4238 =  n_4236 &  n_4237;
assign n_4239 =  n_4235 &  n_4238;
assign n_4240 = ~x_3187 & ~x_3189;
assign n_4241 = ~x_3191 & ~x_3196;
assign n_4242 =  n_4240 &  n_4241;
assign n_4243 = ~x_3173 & ~x_3178;
assign n_4244 = ~x_3180 & ~x_3182;
assign n_4245 =  n_4243 &  n_4244;
assign n_4246 =  n_4242 &  n_4245;
assign n_4247 =  n_4239 &  n_4246;
assign n_4248 =  n_4234 &  n_4247;
assign n_4249 =  n_4035 &  n_4040;
assign n_4250 =  n_4045 &  n_4050;
assign n_4251 =  n_4249 &  n_4250;
assign n_4252 =  n_4061 &  n_4251;
assign n_4253 =  n_4248 &  n_4252;
assign n_4254 =  n_896 &  n_884;
assign n_4255 =  n_4253 &  n_4254;
assign n_4256 =  n_4223 &  n_4255;
assign n_4257 =  n_737 &  n_725;
assign n_4258 =  n_700 &  n_688;
assign n_4259 =  n_4257 &  n_4258;
assign n_4260 =  n_798 &  n_786;
assign n_4261 =  n_774 &  n_749;
assign n_4262 =  n_4260 &  n_4261;
assign n_4263 =  n_4259 &  n_4262;
assign n_4264 =  n_4256 &  n_4263;
assign n_4265 =  n_4220 &  n_4264;
assign n_4266 =  n_4212 &  n_4265;
assign n_4267 =  n_4210 &  n_4266;
assign n_4268 = ~n_1139 &  n_4267;
assign n_4269 = ~n_909 & ~n_860;
assign n_4270 =  n_4268 &  n_4269;
assign n_4271 =  n_4206 &  n_4270;
assign n_4272 = ~n_4068 & ~n_4192;
assign n_4273 = ~n_4072 & ~n_4181;
assign n_4274 =  n_4272 &  n_4273;
assign n_4275 = ~n_615 & ~n_4189;
assign n_4276 = ~n_4197 & ~n_4178;
assign n_4277 =  n_4275 &  n_4276;
assign n_4278 =  n_4274 &  n_4277;
assign n_4279 =  n_4271 &  n_4278;
assign n_4280 = ~x_308 &  x_1725;
assign n_4281 = ~x_1723 & ~n_1325;
assign n_4282 =  n_3691 &  n_4281;
assign n_4283 =  n_3678 & ~n_3680;
assign n_4284 =  n_3673 &  n_3691;
assign n_4285 = ~n_4283 & ~n_4284;
assign n_4286 = ~n_4282 &  n_4285;
assign n_4287 = ~x_1721 & ~x_1722;
assign n_4288 =  n_4286 & ~n_4287;
assign n_4289 =  n_4280 & ~n_4288;
assign n_4290 =  x_1725 & ~n_4289;
assign n_4291 = ~n_4290 &  n_3698;
assign n_4292 = ~x_1471 & ~x_1597;
assign n_4293 = ~n_1226 &  n_4292;
assign n_4294 = ~n_4291 & ~n_4293;
assign n_4295 = ~n_1204 & ~n_1173;
assign n_4296 =  n_4294 &  n_4295;
assign n_4297 = ~n_4279 &  n_4296;
assign n_4298 = ~n_4203 &  n_4297;
assign n_4299 =  x_3233 &  n_4298;
assign n_4300 = ~x_3233 & ~n_4298;
assign n_4301 = ~n_4299 & ~n_4300;
assign n_4302 =  x_319 &  x_3140;
assign n_4303 =  n_1739 &  n_4302;
assign n_4304 =  i_146 &  x_295;
assign n_4305 = ~x_3149 & ~n_4304;
assign n_4306 =  x_3149 &  n_4304;
assign n_4307 = ~n_4305 & ~n_4306;
assign n_4308 = ~i_145 &  x_3150;
assign n_4309 =  i_145 & ~x_3150;
assign n_4310 = ~n_4308 & ~n_4309;
assign n_4311 =  i_143 & ~x_3152;
assign n_4312 = ~i_143 &  x_3152;
assign n_4313 = ~n_4311 & ~n_4312;
assign n_4314 =  n_4310 &  n_4313;
assign n_4315 =  i_148 &  x_295;
assign n_4316 =  x_3146 & ~n_4315;
assign n_4317 =  i_150 &  x_295;
assign n_4318 = ~x_3148 &  n_4317;
assign n_4319 = ~n_4316 & ~n_4318;
assign n_4320 =  n_4314 &  n_4319;
assign n_4321 = ~n_4307 &  n_4320;
assign n_4322 =  x_3148 & ~n_4317;
assign n_4323 =  i_147 &  x_295;
assign n_4324 =  x_3151 & ~n_4323;
assign n_4325 = ~n_4322 & ~n_4324;
assign n_4326 =  i_149 &  x_295;
assign n_4327 = ~x_3145 &  n_4326;
assign n_4328 =  i_144 &  x_295;
assign n_4329 = ~x_3147 &  n_4328;
assign n_4330 = ~n_4327 & ~n_4329;
assign n_4331 =  n_4325 &  n_4330;
assign n_4332 = ~x_3146 &  n_4315;
assign n_4333 =  x_3145 & ~n_4326;
assign n_4334 = ~n_4332 & ~n_4333;
assign n_4335 = ~x_3151 &  n_4323;
assign n_4336 =  x_3147 & ~n_4328;
assign n_4337 = ~n_4335 & ~n_4336;
assign n_4338 =  n_4334 &  n_4337;
assign n_4339 =  n_4331 &  n_4338;
assign n_4340 =  n_4321 &  n_4339;
assign n_4341 =  n_4303 & ~n_4340;
assign n_4342 =  x_3144 &  n_4341;
assign n_4343 =  x_3232 &  n_4342;
assign n_4344 = ~x_3232 & ~n_4342;
assign n_4345 = ~n_4343 & ~n_4344;
assign n_4346 = ~i_2 & ~i_4;
assign n_4347 = ~i_6 & ~i_8;
assign n_4348 =  n_4346 &  n_4347;
assign n_4349 =  x_295 & ~n_4348;
assign n_4350 =  i_7 &  x_295;
assign n_4351 = ~i_8 &  n_4350;
assign n_4352 = ~i_5 & ~i_6;
assign n_4353 =  x_295 & ~n_4352;
assign n_4354 = ~n_4351 &  n_4353;
assign n_4355 = ~i_3 & ~i_4;
assign n_4356 =  n_4354 & ~n_4355;
assign n_4357 =  i_1 &  x_295;
assign n_4358 = ~i_2 &  n_4357;
assign n_4359 =  x_3140 & ~n_4358;
assign n_4360 =  n_4356 &  n_4359;
assign n_4361 = ~n_4349 &  n_4360;
assign n_4362 =  x_3141 &  n_4361;
assign n_4363 =  x_3142 & ~x_3143;
assign n_4364 =  n_4362 & ~n_4363;
assign n_4365 =  x_3231 &  n_4364;
assign n_4366 = ~x_3231 & ~n_4364;
assign n_4367 = ~n_4365 & ~n_4366;
assign n_4368 = ~x_1725 & ~x_1726;
assign n_4369 = ~x_1729 &  n_4368;
assign n_4370 = ~x_1499 & ~n_4369;
assign n_4371 = ~x_2547 & ~x_2548;
assign n_4372 = ~x_2546 &  n_4371;
assign n_4373 = ~x_2545 &  n_4372;
assign n_4374 = ~x_2544 &  n_4373;
assign n_4375 = ~n_4370 &  n_4374;
assign n_4376 =  x_1557 &  n_4375;
assign n_4377 = ~x_314 &  x_2549;
assign n_4378 = ~x_2551 &  x_2552;
assign n_4379 =  n_4377 &  n_4378;
assign n_4380 = ~x_3063 &  n_4379;
assign n_4381 =  x_314 &  x_2549;
assign n_4382 =  x_2551 & ~x_2552;
assign n_4383 =  n_4381 &  n_4382;
assign n_4384 = ~x_3061 &  n_4383;
assign n_4385 = ~n_4380 & ~n_4384;
assign n_4386 =  x_2551 &  x_2552;
assign n_4387 =  n_4386 &  n_4381;
assign n_4388 = ~x_3053 &  n_4387;
assign n_4389 =  n_4377 &  n_4386;
assign n_4390 = ~x_3067 &  n_4389;
assign n_4391 = ~n_4388 & ~n_4390;
assign n_4392 =  n_4385 &  n_4391;
assign n_4393 = ~x_2551 & ~x_2552;
assign n_4394 = ~x_2549 & ~x_2550;
assign n_4395 =  n_4393 &  n_4394;
assign n_4396 = ~x_3054 &  n_4395;
assign n_4397 =  n_4386 &  n_4394;
assign n_4398 = ~x_3066 &  n_4397;
assign n_4399 = ~n_4396 & ~n_4398;
assign n_4400 =  n_4394 &  n_4378;
assign n_4401 = ~x_3062 &  n_4400;
assign n_4402 = ~x_2549 &  x_2550;
assign n_4403 =  n_4393 &  n_4402;
assign n_4404 = ~x_3056 &  n_4403;
assign n_4405 = ~n_4401 & ~n_4404;
assign n_4406 =  n_4399 &  n_4405;
assign n_4407 =  n_4392 &  n_4406;
assign n_4408 =  n_4394 &  n_4382;
assign n_4409 = ~x_3058 &  n_4408;
assign n_4410 =  n_4377 &  n_4393;
assign n_4411 = ~x_3055 &  n_4410;
assign n_4412 = ~n_4409 & ~n_4411;
assign n_4413 =  n_4402 &  n_4382;
assign n_4414 = ~x_3060 &  n_4413;
assign n_4415 =  n_4386 &  n_4402;
assign n_4416 = ~x_3068 &  n_4415;
assign n_4417 = ~n_4414 & ~n_4416;
assign n_4418 =  n_4412 &  n_4417;
assign n_4419 =  n_4381 &  n_4378;
assign n_4420 = ~x_3065 &  n_4419;
assign n_4421 =  n_4377 &  n_4382;
assign n_4422 = ~x_3059 &  n_4421;
assign n_4423 = ~n_4420 & ~n_4422;
assign n_4424 =  n_4393 &  n_4381;
assign n_4425 = ~x_3057 &  n_4424;
assign n_4426 =  n_4402 &  n_4378;
assign n_4427 = ~x_3064 &  n_4426;
assign n_4428 = ~n_4425 & ~n_4427;
assign n_4429 =  n_4423 &  n_4428;
assign n_4430 =  n_4418 &  n_4429;
assign n_4431 =  n_4407 &  n_4430;
assign n_4432 = ~x_1559 &  n_4431;
assign n_4433 =  x_1559 & ~n_4431;
assign n_4434 = ~n_4432 & ~n_4433;
assign n_4435 = ~x_3048 &  n_4426;
assign n_4436 = ~x_3047 &  n_4379;
assign n_4437 = ~n_4435 & ~n_4436;
assign n_4438 = ~x_3037 &  n_4387;
assign n_4439 = ~x_3043 &  n_4421;
assign n_4440 = ~n_4438 & ~n_4439;
assign n_4441 =  n_4437 &  n_4440;
assign n_4442 = ~x_3045 &  n_4383;
assign n_4443 = ~x_3042 &  n_4408;
assign n_4444 = ~n_4442 & ~n_4443;
assign n_4445 = ~x_3039 &  n_4410;
assign n_4446 = ~x_3049 &  n_4419;
assign n_4447 = ~n_4445 & ~n_4446;
assign n_4448 =  n_4444 &  n_4447;
assign n_4449 =  n_4441 &  n_4448;
assign n_4450 = ~x_3038 &  n_4395;
assign n_4451 = ~x_3046 &  n_4400;
assign n_4452 = ~n_4450 & ~n_4451;
assign n_4453 = ~x_3044 &  n_4413;
assign n_4454 = ~x_3040 &  n_4403;
assign n_4455 = ~n_4453 & ~n_4454;
assign n_4456 =  n_4452 &  n_4455;
assign n_4457 = ~x_3050 &  n_4397;
assign n_4458 = ~x_3051 &  n_4389;
assign n_4459 = ~n_4457 & ~n_4458;
assign n_4460 = ~x_3052 &  n_4415;
assign n_4461 = ~x_3041 &  n_4424;
assign n_4462 = ~n_4460 & ~n_4461;
assign n_4463 =  n_4459 &  n_4462;
assign n_4464 =  n_4456 &  n_4463;
assign n_4465 =  n_4449 &  n_4464;
assign n_4466 =  x_1558 & ~n_4465;
assign n_4467 = ~x_1558 &  n_4465;
assign n_4468 = ~n_4466 & ~n_4467;
assign n_4469 = ~x_3023 &  n_4410;
assign n_4470 = ~x_3036 &  n_4415;
assign n_4471 = ~n_4469 & ~n_4470;
assign n_4472 = ~x_3021 &  n_4387;
assign n_4473 = ~x_3026 &  n_4408;
assign n_4474 = ~n_4472 & ~n_4473;
assign n_4475 =  n_4471 &  n_4474;
assign n_4476 = ~x_3031 &  n_4379;
assign n_4477 = ~x_3025 &  n_4424;
assign n_4478 = ~n_4476 & ~n_4477;
assign n_4479 = ~x_3035 &  n_4389;
assign n_4480 = ~x_3024 &  n_4403;
assign n_4481 = ~n_4479 & ~n_4480;
assign n_4482 =  n_4478 &  n_4481;
assign n_4483 =  n_4475 &  n_4482;
assign n_4484 = ~x_3034 &  n_4397;
assign n_4485 = ~x_3022 &  n_4395;
assign n_4486 = ~n_4484 & ~n_4485;
assign n_4487 = ~x_3033 &  n_4419;
assign n_4488 = ~x_3028 &  n_4413;
assign n_4489 = ~n_4487 & ~n_4488;
assign n_4490 =  n_4486 &  n_4489;
assign n_4491 = ~x_3027 &  n_4421;
assign n_4492 = ~x_3030 &  n_4400;
assign n_4493 = ~n_4491 & ~n_4492;
assign n_4494 = ~x_3032 &  n_4426;
assign n_4495 = ~x_3029 &  n_4383;
assign n_4496 = ~n_4494 & ~n_4495;
assign n_4497 =  n_4493 &  n_4496;
assign n_4498 =  n_4490 &  n_4497;
assign n_4499 =  n_4483 &  n_4498;
assign n_4500 =  x_1501 & ~n_4499;
assign n_4501 = ~x_1501 &  n_4499;
assign n_4502 = ~n_4500 & ~n_4501;
assign n_4503 = ~x_3015 &  n_4379;
assign n_4504 = ~x_3007 &  n_4410;
assign n_4505 = ~n_4503 & ~n_4504;
assign n_4506 = ~x_3005 &  n_4387;
assign n_4507 = ~x_3010 &  n_4408;
assign n_4508 = ~n_4506 & ~n_4507;
assign n_4509 =  n_4505 &  n_4508;
assign n_4510 = ~x_3020 &  n_4415;
assign n_4511 = ~x_3019 &  n_4389;
assign n_4512 = ~n_4510 & ~n_4511;
assign n_4513 = ~x_3012 &  n_4413;
assign n_4514 = ~x_3011 &  n_4421;
assign n_4515 = ~n_4513 & ~n_4514;
assign n_4516 =  n_4512 &  n_4515;
assign n_4517 =  n_4509 &  n_4516;
assign n_4518 = ~x_3018 &  n_4397;
assign n_4519 = ~x_3014 &  n_4400;
assign n_4520 = ~n_4518 & ~n_4519;
assign n_4521 = ~x_3009 &  n_4424;
assign n_4522 = ~x_3006 &  n_4395;
assign n_4523 = ~n_4521 & ~n_4522;
assign n_4524 =  n_4520 &  n_4523;
assign n_4525 = ~x_3008 &  n_4403;
assign n_4526 = ~x_3016 &  n_4426;
assign n_4527 = ~n_4525 & ~n_4526;
assign n_4528 = ~x_3013 &  n_4383;
assign n_4529 = ~x_3017 &  n_4419;
assign n_4530 = ~n_4528 & ~n_4529;
assign n_4531 =  n_4527 &  n_4530;
assign n_4532 =  n_4524 &  n_4531;
assign n_4533 =  n_4517 &  n_4532;
assign n_4534 =  x_1502 & ~n_4533;
assign n_4535 = ~x_1502 &  n_4533;
assign n_4536 = ~n_4534 & ~n_4535;
assign n_4537 = ~x_2992 &  n_4403;
assign n_4538 = ~x_2997 &  n_4383;
assign n_4539 = ~n_4537 & ~n_4538;
assign n_4540 = ~x_2989 &  n_4387;
assign n_4541 = ~x_2996 &  n_4413;
assign n_4542 = ~n_4540 & ~n_4541;
assign n_4543 =  n_4539 &  n_4542;
assign n_4544 = ~x_3001 &  n_4419;
assign n_4545 = ~x_2999 &  n_4379;
assign n_4546 = ~n_4544 & ~n_4545;
assign n_4547 = ~x_2990 &  n_4395;
assign n_4548 = ~x_2994 &  n_4408;
assign n_4549 = ~n_4547 & ~n_4548;
assign n_4550 =  n_4546 &  n_4549;
assign n_4551 =  n_4543 &  n_4550;
assign n_4552 = ~x_2995 &  n_4421;
assign n_4553 = ~x_3003 &  n_4389;
assign n_4554 = ~n_4552 & ~n_4553;
assign n_4555 = ~x_2998 &  n_4400;
assign n_4556 = ~x_2993 &  n_4424;
assign n_4557 = ~n_4555 & ~n_4556;
assign n_4558 =  n_4554 &  n_4557;
assign n_4559 = ~x_3000 &  n_4426;
assign n_4560 = ~x_2991 &  n_4410;
assign n_4561 = ~n_4559 & ~n_4560;
assign n_4562 = ~x_3004 &  n_4415;
assign n_4563 = ~x_3002 &  n_4397;
assign n_4564 = ~n_4562 & ~n_4563;
assign n_4565 =  n_4561 &  n_4564;
assign n_4566 =  n_4558 &  n_4565;
assign n_4567 =  n_4551 &  n_4566;
assign n_4568 =  x_1503 & ~n_4567;
assign n_4569 = ~x_1503 &  n_4567;
assign n_4570 = ~n_4568 & ~n_4569;
assign n_4571 = ~x_2983 &  n_4379;
assign n_4572 = ~x_2980 &  n_4413;
assign n_4573 = ~n_4571 & ~n_4572;
assign n_4574 = ~x_2973 &  n_4387;
assign n_4575 = ~x_2986 &  n_4397;
assign n_4576 = ~n_4574 & ~n_4575;
assign n_4577 =  n_4573 &  n_4576;
assign n_4578 = ~x_2982 &  n_4400;
assign n_4579 = ~x_2974 &  n_4395;
assign n_4580 = ~n_4578 & ~n_4579;
assign n_4581 = ~x_2987 &  n_4389;
assign n_4582 = ~x_2978 &  n_4408;
assign n_4583 = ~n_4581 & ~n_4582;
assign n_4584 =  n_4580 &  n_4583;
assign n_4585 =  n_4577 &  n_4584;
assign n_4586 = ~x_2984 &  n_4426;
assign n_4587 = ~x_2979 &  n_4421;
assign n_4588 = ~n_4586 & ~n_4587;
assign n_4589 = ~x_2976 &  n_4403;
assign n_4590 = ~x_2981 &  n_4383;
assign n_4591 = ~n_4589 & ~n_4590;
assign n_4592 =  n_4588 &  n_4591;
assign n_4593 = ~x_2977 &  n_4424;
assign n_4594 = ~x_2975 &  n_4410;
assign n_4595 = ~n_4593 & ~n_4594;
assign n_4596 = ~x_2985 &  n_4419;
assign n_4597 = ~x_2988 &  n_4415;
assign n_4598 = ~n_4596 & ~n_4597;
assign n_4599 =  n_4595 &  n_4598;
assign n_4600 =  n_4592 &  n_4599;
assign n_4601 =  n_4585 &  n_4600;
assign n_4602 =  x_1504 & ~n_4601;
assign n_4603 = ~x_1504 &  n_4601;
assign n_4604 = ~n_4602 & ~n_4603;
assign n_4605 = ~x_2968 &  n_4426;
assign n_4606 = ~x_2967 &  n_4379;
assign n_4607 = ~n_4605 & ~n_4606;
assign n_4608 = ~x_2957 &  n_4387;
assign n_4609 = ~x_2959 &  n_4410;
assign n_4610 = ~n_4608 & ~n_4609;
assign n_4611 =  n_4607 &  n_4610;
assign n_4612 = ~x_2971 &  n_4389;
assign n_4613 = ~x_2963 &  n_4421;
assign n_4614 = ~n_4612 & ~n_4613;
assign n_4615 = ~x_2969 &  n_4419;
assign n_4616 = ~x_2964 &  n_4413;
assign n_4617 = ~n_4615 & ~n_4616;
assign n_4618 =  n_4614 &  n_4617;
assign n_4619 =  n_4611 &  n_4618;
assign n_4620 = ~x_2958 &  n_4395;
assign n_4621 = ~x_2970 &  n_4397;
assign n_4622 = ~n_4620 & ~n_4621;
assign n_4623 = ~x_2960 &  n_4403;
assign n_4624 = ~x_2965 &  n_4383;
assign n_4625 = ~n_4623 & ~n_4624;
assign n_4626 =  n_4622 &  n_4625;
assign n_4627 = ~x_2961 &  n_4424;
assign n_4628 = ~x_2962 &  n_4408;
assign n_4629 = ~n_4627 & ~n_4628;
assign n_4630 = ~x_2966 &  n_4400;
assign n_4631 = ~x_2972 &  n_4415;
assign n_4632 = ~n_4630 & ~n_4631;
assign n_4633 =  n_4629 &  n_4632;
assign n_4634 =  n_4626 &  n_4633;
assign n_4635 =  n_4619 &  n_4634;
assign n_4636 =  x_1505 & ~n_4635;
assign n_4637 = ~x_1505 &  n_4635;
assign n_4638 = ~n_4636 & ~n_4637;
assign n_4639 = ~x_2953 &  n_4419;
assign n_4640 = ~x_2951 &  n_4379;
assign n_4641 = ~n_4639 & ~n_4640;
assign n_4642 = ~x_2941 &  n_4387;
assign n_4643 = ~x_2946 &  n_4408;
assign n_4644 = ~n_4642 & ~n_4643;
assign n_4645 =  n_4641 &  n_4644;
assign n_4646 = ~x_2955 &  n_4389;
assign n_4647 = ~x_2952 &  n_4426;
assign n_4648 = ~n_4646 & ~n_4647;
assign n_4649 = ~x_2947 &  n_4421;
assign n_4650 = ~x_2944 &  n_4403;
assign n_4651 = ~n_4649 & ~n_4650;
assign n_4652 =  n_4648 &  n_4651;
assign n_4653 =  n_4645 &  n_4652;
assign n_4654 = ~x_2943 &  n_4410;
assign n_4655 = ~x_2954 &  n_4397;
assign n_4656 = ~n_4654 & ~n_4655;
assign n_4657 = ~x_2948 &  n_4413;
assign n_4658 = ~x_2942 &  n_4395;
assign n_4659 = ~n_4657 & ~n_4658;
assign n_4660 =  n_4656 &  n_4659;
assign n_4661 = ~x_2950 &  n_4400;
assign n_4662 = ~x_2949 &  n_4383;
assign n_4663 = ~n_4661 & ~n_4662;
assign n_4664 = ~x_2945 &  n_4424;
assign n_4665 = ~x_2956 &  n_4415;
assign n_4666 = ~n_4664 & ~n_4665;
assign n_4667 =  n_4663 &  n_4666;
assign n_4668 =  n_4660 &  n_4667;
assign n_4669 =  n_4653 &  n_4668;
assign n_4670 =  x_1506 & ~n_4669;
assign n_4671 = ~x_1506 &  n_4669;
assign n_4672 = ~n_4670 & ~n_4671;
assign n_4673 = ~x_2927 &  n_4410;
assign n_4674 = ~x_2933 &  n_4383;
assign n_4675 = ~n_4673 & ~n_4674;
assign n_4676 = ~x_2925 &  n_4387;
assign n_4677 = ~x_2932 &  n_4413;
assign n_4678 = ~n_4676 & ~n_4677;
assign n_4679 =  n_4675 &  n_4678;
assign n_4680 = ~x_2939 &  n_4389;
assign n_4681 = ~x_2934 &  n_4400;
assign n_4682 = ~n_4680 & ~n_4681;
assign n_4683 = ~x_2937 &  n_4419;
assign n_4684 = ~x_2931 &  n_4421;
assign n_4685 = ~n_4683 & ~n_4684;
assign n_4686 =  n_4682 &  n_4685;
assign n_4687 =  n_4679 &  n_4686;
assign n_4688 = ~x_2938 &  n_4397;
assign n_4689 = ~x_2935 &  n_4379;
assign n_4690 = ~n_4688 & ~n_4689;
assign n_4691 = ~x_2936 &  n_4426;
assign n_4692 = ~x_2930 &  n_4408;
assign n_4693 = ~n_4691 & ~n_4692;
assign n_4694 =  n_4690 &  n_4693;
assign n_4695 = ~x_2940 &  n_4415;
assign n_4696 = ~x_2926 &  n_4395;
assign n_4697 = ~n_4695 & ~n_4696;
assign n_4698 = ~x_2929 &  n_4424;
assign n_4699 = ~x_2928 &  n_4403;
assign n_4700 = ~n_4698 & ~n_4699;
assign n_4701 =  n_4697 &  n_4700;
assign n_4702 =  n_4694 &  n_4701;
assign n_4703 =  n_4687 &  n_4702;
assign n_4704 =  x_1507 & ~n_4703;
assign n_4705 = ~x_1507 &  n_4703;
assign n_4706 = ~n_4704 & ~n_4705;
assign n_4707 = ~x_2916 &  n_4413;
assign n_4708 = ~x_2923 &  n_4389;
assign n_4709 = ~n_4707 & ~n_4708;
assign n_4710 = ~x_2909 &  n_4387;
assign n_4711 = ~x_2914 &  n_4408;
assign n_4712 = ~n_4710 & ~n_4711;
assign n_4713 =  n_4709 &  n_4712;
assign n_4714 = ~x_2922 &  n_4397;
assign n_4715 = ~x_2918 &  n_4400;
assign n_4716 = ~n_4714 & ~n_4715;
assign n_4717 = ~x_2921 &  n_4419;
assign n_4718 = ~x_2912 &  n_4403;
assign n_4719 = ~n_4717 & ~n_4718;
assign n_4720 =  n_4716 &  n_4719;
assign n_4721 =  n_4713 &  n_4720;
assign n_4722 = ~x_2919 &  n_4379;
assign n_4723 = ~x_2915 &  n_4421;
assign n_4724 = ~n_4722 & ~n_4723;
assign n_4725 = ~x_2911 &  n_4410;
assign n_4726 = ~x_2913 &  n_4424;
assign n_4727 = ~n_4725 & ~n_4726;
assign n_4728 =  n_4724 &  n_4727;
assign n_4729 = ~x_2924 &  n_4415;
assign n_4730 = ~x_2910 &  n_4395;
assign n_4731 = ~n_4729 & ~n_4730;
assign n_4732 = ~x_2920 &  n_4426;
assign n_4733 = ~x_2917 &  n_4383;
assign n_4734 = ~n_4732 & ~n_4733;
assign n_4735 =  n_4731 &  n_4734;
assign n_4736 =  n_4728 &  n_4735;
assign n_4737 =  n_4721 &  n_4736;
assign n_4738 =  x_1508 & ~n_4737;
assign n_4739 = ~x_1508 &  n_4737;
assign n_4740 = ~n_4738 & ~n_4739;
assign n_4741 = ~x_2905 &  n_4419;
assign n_4742 = ~x_2900 &  n_4413;
assign n_4743 = ~n_4741 & ~n_4742;
assign n_4744 = ~x_2893 &  n_4387;
assign n_4745 = ~x_2899 &  n_4421;
assign n_4746 = ~n_4744 & ~n_4745;
assign n_4747 =  n_4743 &  n_4746;
assign n_4748 = ~x_2901 &  n_4383;
assign n_4749 = ~x_2902 &  n_4400;
assign n_4750 = ~n_4748 & ~n_4749;
assign n_4751 = ~x_2906 &  n_4397;
assign n_4752 = ~x_2897 &  n_4424;
assign n_4753 = ~n_4751 & ~n_4752;
assign n_4754 =  n_4750 &  n_4753;
assign n_4755 =  n_4747 &  n_4754;
assign n_4756 = ~x_2898 &  n_4408;
assign n_4757 = ~x_2903 &  n_4379;
assign n_4758 = ~n_4756 & ~n_4757;
assign n_4759 = ~x_2896 &  n_4403;
assign n_4760 = ~x_2908 &  n_4415;
assign n_4761 = ~n_4759 & ~n_4760;
assign n_4762 =  n_4758 &  n_4761;
assign n_4763 = ~x_2894 &  n_4395;
assign n_4764 = ~x_2907 &  n_4389;
assign n_4765 = ~n_4763 & ~n_4764;
assign n_4766 = ~x_2895 &  n_4410;
assign n_4767 = ~x_2904 &  n_4426;
assign n_4768 = ~n_4766 & ~n_4767;
assign n_4769 =  n_4765 &  n_4768;
assign n_4770 =  n_4762 &  n_4769;
assign n_4771 =  n_4755 &  n_4770;
assign n_4772 =  x_1509 & ~n_4771;
assign n_4773 = ~x_1509 &  n_4771;
assign n_4774 = ~n_4772 & ~n_4773;
assign n_4775 = ~x_2889 &  n_4419;
assign n_4776 = ~x_2892 &  n_4415;
assign n_4777 = ~n_4775 & ~n_4776;
assign n_4778 = ~x_2877 &  n_4387;
assign n_4779 = ~x_2883 &  n_4421;
assign n_4780 = ~n_4778 & ~n_4779;
assign n_4781 =  n_4777 &  n_4780;
assign n_4782 = ~x_2891 &  n_4389;
assign n_4783 = ~x_2887 &  n_4379;
assign n_4784 = ~n_4782 & ~n_4783;
assign n_4785 = ~x_2884 &  n_4413;
assign n_4786 = ~x_2879 &  n_4410;
assign n_4787 = ~n_4785 & ~n_4786;
assign n_4788 =  n_4784 &  n_4787;
assign n_4789 =  n_4781 &  n_4788;
assign n_4790 = ~x_2886 &  n_4400;
assign n_4791 = ~x_2888 &  n_4426;
assign n_4792 = ~n_4790 & ~n_4791;
assign n_4793 = ~x_2880 &  n_4403;
assign n_4794 = ~x_2890 &  n_4397;
assign n_4795 = ~n_4793 & ~n_4794;
assign n_4796 =  n_4792 &  n_4795;
assign n_4797 = ~x_2885 &  n_4383;
assign n_4798 = ~x_2878 &  n_4395;
assign n_4799 = ~n_4797 & ~n_4798;
assign n_4800 = ~x_2881 &  n_4424;
assign n_4801 = ~x_2882 &  n_4408;
assign n_4802 = ~n_4800 & ~n_4801;
assign n_4803 =  n_4799 &  n_4802;
assign n_4804 =  n_4796 &  n_4803;
assign n_4805 =  n_4789 &  n_4804;
assign n_4806 =  x_1510 & ~n_4805;
assign n_4807 = ~x_1510 &  n_4805;
assign n_4808 = ~n_4806 & ~n_4807;
assign n_4809 = ~x_2868 &  n_4413;
assign n_4810 = ~x_2869 &  n_4383;
assign n_4811 = ~n_4809 & ~n_4810;
assign n_4812 = ~x_2861 &  n_4387;
assign n_4813 = ~x_2876 &  n_4415;
assign n_4814 = ~n_4812 & ~n_4813;
assign n_4815 =  n_4811 &  n_4814;
assign n_4816 = ~x_2870 &  n_4400;
assign n_4817 = ~x_2863 &  n_4410;
assign n_4818 = ~n_4816 & ~n_4817;
assign n_4819 = ~x_2867 &  n_4421;
assign n_4820 = ~x_2862 &  n_4395;
assign n_4821 = ~n_4819 & ~n_4820;
assign n_4822 =  n_4818 &  n_4821;
assign n_4823 =  n_4815 &  n_4822;
assign n_4824 = ~x_2866 &  n_4408;
assign n_4825 = ~x_2871 &  n_4379;
assign n_4826 = ~n_4824 & ~n_4825;
assign n_4827 = ~x_2874 &  n_4397;
assign n_4828 = ~x_2872 &  n_4426;
assign n_4829 = ~n_4827 & ~n_4828;
assign n_4830 =  n_4826 &  n_4829;
assign n_4831 = ~x_2865 &  n_4424;
assign n_4832 = ~x_2875 &  n_4389;
assign n_4833 = ~n_4831 & ~n_4832;
assign n_4834 = ~x_2864 &  n_4403;
assign n_4835 = ~x_2873 &  n_4419;
assign n_4836 = ~n_4834 & ~n_4835;
assign n_4837 =  n_4833 &  n_4836;
assign n_4838 =  n_4830 &  n_4837;
assign n_4839 =  n_4823 &  n_4838;
assign n_4840 =  x_1511 & ~n_4839;
assign n_4841 = ~x_1511 &  n_4839;
assign n_4842 = ~n_4840 & ~n_4841;
assign n_4843 = ~x_2853 &  n_4383;
assign n_4844 = ~x_2860 &  n_4415;
assign n_4845 = ~n_4843 & ~n_4844;
assign n_4846 = ~x_2845 &  n_4387;
assign n_4847 = ~x_2859 &  n_4389;
assign n_4848 = ~n_4846 & ~n_4847;
assign n_4849 =  n_4845 &  n_4848;
assign n_4850 = ~x_2850 &  n_4408;
assign n_4851 = ~x_2847 &  n_4410;
assign n_4852 = ~n_4850 & ~n_4851;
assign n_4853 = ~x_2855 &  n_4379;
assign n_4854 = ~x_2851 &  n_4421;
assign n_4855 = ~n_4853 & ~n_4854;
assign n_4856 =  n_4852 &  n_4855;
assign n_4857 =  n_4849 &  n_4856;
assign n_4858 = ~x_2854 &  n_4400;
assign n_4859 = ~x_2858 &  n_4397;
assign n_4860 = ~n_4858 & ~n_4859;
assign n_4861 = ~x_2856 &  n_4426;
assign n_4862 = ~x_2848 &  n_4403;
assign n_4863 = ~n_4861 & ~n_4862;
assign n_4864 =  n_4860 &  n_4863;
assign n_4865 = ~x_2857 &  n_4419;
assign n_4866 = ~x_2846 &  n_4395;
assign n_4867 = ~n_4865 & ~n_4866;
assign n_4868 = ~x_2849 &  n_4424;
assign n_4869 = ~x_2852 &  n_4413;
assign n_4870 = ~n_4868 & ~n_4869;
assign n_4871 =  n_4867 &  n_4870;
assign n_4872 =  n_4864 &  n_4871;
assign n_4873 =  n_4857 &  n_4872;
assign n_4874 =  x_1512 & ~n_4873;
assign n_4875 = ~x_1512 &  n_4873;
assign n_4876 = ~n_4874 & ~n_4875;
assign n_4877 = ~x_2837 &  n_4383;
assign n_4878 = ~x_2843 &  n_4389;
assign n_4879 = ~n_4877 & ~n_4878;
assign n_4880 = ~x_2829 &  n_4387;
assign n_4881 = ~x_2842 &  n_4397;
assign n_4882 = ~n_4880 & ~n_4881;
assign n_4883 =  n_4879 &  n_4882;
assign n_4884 = ~x_2836 &  n_4413;
assign n_4885 = ~x_2834 &  n_4408;
assign n_4886 = ~n_4884 & ~n_4885;
assign n_4887 = ~x_2832 &  n_4403;
assign n_4888 = ~x_2840 &  n_4426;
assign n_4889 = ~n_4887 & ~n_4888;
assign n_4890 =  n_4886 &  n_4889;
assign n_4891 =  n_4883 &  n_4890;
assign n_4892 = ~x_2831 &  n_4410;
assign n_4893 = ~x_2838 &  n_4400;
assign n_4894 = ~n_4892 & ~n_4893;
assign n_4895 = ~x_2839 &  n_4379;
assign n_4896 = ~x_2844 &  n_4415;
assign n_4897 = ~n_4895 & ~n_4896;
assign n_4898 =  n_4894 &  n_4897;
assign n_4899 = ~x_2835 &  n_4421;
assign n_4900 = ~x_2830 &  n_4395;
assign n_4901 = ~n_4899 & ~n_4900;
assign n_4902 = ~x_2841 &  n_4419;
assign n_4903 = ~x_2833 &  n_4424;
assign n_4904 = ~n_4902 & ~n_4903;
assign n_4905 =  n_4901 &  n_4904;
assign n_4906 =  n_4898 &  n_4905;
assign n_4907 =  n_4891 &  n_4906;
assign n_4908 =  x_1513 & ~n_4907;
assign n_4909 = ~x_1513 &  n_4907;
assign n_4910 = ~n_4908 & ~n_4909;
assign n_4911 = ~x_2828 &  n_4415;
assign n_4912 = ~x_2818 &  n_4408;
assign n_4913 = ~n_4911 & ~n_4912;
assign n_4914 = ~x_2813 &  n_4387;
assign n_4915 = ~x_2823 &  n_4379;
assign n_4916 = ~n_4914 & ~n_4915;
assign n_4917 =  n_4913 &  n_4916;
assign n_4918 = ~x_2822 &  n_4400;
assign n_4919 = ~x_2814 &  n_4395;
assign n_4920 = ~n_4918 & ~n_4919;
assign n_4921 = ~x_2824 &  n_4426;
assign n_4922 = ~x_2826 &  n_4397;
assign n_4923 = ~n_4921 & ~n_4922;
assign n_4924 =  n_4920 &  n_4923;
assign n_4925 =  n_4917 &  n_4924;
assign n_4926 = ~x_2827 &  n_4389;
assign n_4927 = ~x_2819 &  n_4421;
assign n_4928 = ~n_4926 & ~n_4927;
assign n_4929 = ~x_2816 &  n_4403;
assign n_4930 = ~x_2821 &  n_4383;
assign n_4931 = ~n_4929 & ~n_4930;
assign n_4932 =  n_4928 &  n_4931;
assign n_4933 = ~x_2825 &  n_4419;
assign n_4934 = ~x_2815 &  n_4410;
assign n_4935 = ~n_4933 & ~n_4934;
assign n_4936 = ~x_2820 &  n_4413;
assign n_4937 = ~x_2817 &  n_4424;
assign n_4938 = ~n_4936 & ~n_4937;
assign n_4939 =  n_4935 &  n_4938;
assign n_4940 =  n_4932 &  n_4939;
assign n_4941 =  n_4925 &  n_4940;
assign n_4942 =  x_1514 & ~n_4941;
assign n_4943 = ~x_1514 &  n_4941;
assign n_4944 = ~n_4942 & ~n_4943;
assign n_4945 = ~x_2806 &  n_4400;
assign n_4946 = ~x_2804 &  n_4413;
assign n_4947 = ~n_4945 & ~n_4946;
assign n_4948 = ~x_2797 &  n_4387;
assign n_4949 = ~x_2798 &  n_4395;
assign n_4950 = ~n_4948 & ~n_4949;
assign n_4951 =  n_4947 &  n_4950;
assign n_4952 = ~x_2803 &  n_4421;
assign n_4953 = ~x_2809 &  n_4419;
assign n_4954 = ~n_4952 & ~n_4953;
assign n_4955 = ~x_2802 &  n_4408;
assign n_4956 = ~x_2800 &  n_4403;
assign n_4957 = ~n_4955 & ~n_4956;
assign n_4958 =  n_4954 &  n_4957;
assign n_4959 =  n_4951 &  n_4958;
assign n_4960 = ~x_2810 &  n_4397;
assign n_4961 = ~x_2807 &  n_4379;
assign n_4962 = ~n_4960 & ~n_4961;
assign n_4963 = ~x_2801 &  n_4424;
assign n_4964 = ~x_2799 &  n_4410;
assign n_4965 = ~n_4963 & ~n_4964;
assign n_4966 =  n_4962 &  n_4965;
assign n_4967 = ~x_2811 &  n_4389;
assign n_4968 = ~x_2808 &  n_4426;
assign n_4969 = ~n_4967 & ~n_4968;
assign n_4970 = ~x_2812 &  n_4415;
assign n_4971 = ~x_2805 &  n_4383;
assign n_4972 = ~n_4970 & ~n_4971;
assign n_4973 =  n_4969 &  n_4972;
assign n_4974 =  n_4966 &  n_4973;
assign n_4975 =  n_4959 &  n_4974;
assign n_4976 =  x_1515 & ~n_4975;
assign n_4977 = ~x_1515 &  n_4975;
assign n_4978 = ~n_4976 & ~n_4977;
assign n_4979 = ~x_2788 &  n_4413;
assign n_4980 = ~x_2793 &  n_4419;
assign n_4981 = ~n_4979 & ~n_4980;
assign n_4982 = ~x_2781 &  n_4387;
assign n_4983 = ~x_2786 &  n_4408;
assign n_4984 = ~n_4982 & ~n_4983;
assign n_4985 =  n_4981 &  n_4984;
assign n_4986 = ~x_2791 &  n_4379;
assign n_4987 = ~x_2795 &  n_4389;
assign n_4988 = ~n_4986 & ~n_4987;
assign n_4989 = ~x_2794 &  n_4397;
assign n_4990 = ~x_2784 &  n_4403;
assign n_4991 = ~n_4989 & ~n_4990;
assign n_4992 =  n_4988 &  n_4991;
assign n_4993 =  n_4985 &  n_4992;
assign n_4994 = ~x_2790 &  n_4400;
assign n_4995 = ~x_2787 &  n_4421;
assign n_4996 = ~n_4994 & ~n_4995;
assign n_4997 = ~x_2783 &  n_4410;
assign n_4998 = ~x_2785 &  n_4424;
assign n_4999 = ~n_4997 & ~n_4998;
assign n_5000 =  n_4996 &  n_4999;
assign n_5001 = ~x_2796 &  n_4415;
assign n_5002 = ~x_2782 &  n_4395;
assign n_5003 = ~n_5001 & ~n_5002;
assign n_5004 = ~x_2789 &  n_4383;
assign n_5005 = ~x_2792 &  n_4426;
assign n_5006 = ~n_5004 & ~n_5005;
assign n_5007 =  n_5003 &  n_5006;
assign n_5008 =  n_5000 &  n_5007;
assign n_5009 =  n_4993 &  n_5008;
assign n_5010 =  x_1516 & ~n_5009;
assign n_5011 = ~x_1516 &  n_5009;
assign n_5012 = ~n_5010 & ~n_5011;
assign n_5013 = ~x_2773 &  n_4383;
assign n_5014 = ~x_2776 &  n_4426;
assign n_5015 = ~n_5013 & ~n_5014;
assign n_5016 = ~x_2765 &  n_4387;
assign n_5017 = ~x_2779 &  n_4389;
assign n_5018 = ~n_5016 & ~n_5017;
assign n_5019 =  n_5015 &  n_5018;
assign n_5020 = ~x_2774 &  n_4400;
assign n_5021 = ~x_2766 &  n_4395;
assign n_5022 = ~n_5020 & ~n_5021;
assign n_5023 = ~x_2775 &  n_4379;
assign n_5024 = ~x_2772 &  n_4413;
assign n_5025 = ~n_5023 & ~n_5024;
assign n_5026 =  n_5022 &  n_5025;
assign n_5027 =  n_5019 &  n_5026;
assign n_5028 = ~x_2767 &  n_4410;
assign n_5029 = ~x_2770 &  n_4408;
assign n_5030 = ~n_5028 & ~n_5029;
assign n_5031 = ~x_2777 &  n_4419;
assign n_5032 = ~x_2768 &  n_4403;
assign n_5033 = ~n_5031 & ~n_5032;
assign n_5034 =  n_5030 &  n_5033;
assign n_5035 = ~x_2769 &  n_4424;
assign n_5036 = ~x_2771 &  n_4421;
assign n_5037 = ~n_5035 & ~n_5036;
assign n_5038 = ~x_2778 &  n_4397;
assign n_5039 = ~x_2780 &  n_4415;
assign n_5040 = ~n_5038 & ~n_5039;
assign n_5041 =  n_5037 &  n_5040;
assign n_5042 =  n_5034 &  n_5041;
assign n_5043 =  n_5027 &  n_5042;
assign n_5044 =  x_1517 & ~n_5043;
assign n_5045 = ~x_1517 &  n_5043;
assign n_5046 = ~n_5044 & ~n_5045;
assign n_5047 = ~x_2761 &  n_4419;
assign n_5048 = ~x_2757 &  n_4383;
assign n_5049 = ~n_5047 & ~n_5048;
assign n_5050 = ~x_2749 &  n_4387;
assign n_5051 = ~x_2763 &  n_4389;
assign n_5052 = ~n_5050 & ~n_5051;
assign n_5053 =  n_5049 &  n_5052;
assign n_5054 = ~x_2759 &  n_4379;
assign n_5055 = ~x_2750 &  n_4395;
assign n_5056 = ~n_5054 & ~n_5055;
assign n_5057 = ~x_2751 &  n_4410;
assign n_5058 = ~x_2754 &  n_4408;
assign n_5059 = ~n_5057 & ~n_5058;
assign n_5060 =  n_5056 &  n_5059;
assign n_5061 =  n_5053 &  n_5060;
assign n_5062 = ~x_2762 &  n_4397;
assign n_5063 = ~x_2755 &  n_4421;
assign n_5064 = ~n_5062 & ~n_5063;
assign n_5065 = ~x_2756 &  n_4413;
assign n_5066 = ~x_2752 &  n_4403;
assign n_5067 = ~n_5065 & ~n_5066;
assign n_5068 =  n_5064 &  n_5067;
assign n_5069 = ~x_2764 &  n_4415;
assign n_5070 = ~x_2758 &  n_4400;
assign n_5071 = ~n_5069 & ~n_5070;
assign n_5072 = ~x_2753 &  n_4424;
assign n_5073 = ~x_2760 &  n_4426;
assign n_5074 = ~n_5072 & ~n_5073;
assign n_5075 =  n_5071 &  n_5074;
assign n_5076 =  n_5068 &  n_5075;
assign n_5077 =  n_5061 &  n_5076;
assign n_5078 =  x_1518 & ~n_5077;
assign n_5079 = ~x_1518 &  n_5077;
assign n_5080 = ~n_5078 & ~n_5079;
assign n_5081 = ~x_2742 &  n_4400;
assign n_5082 = ~x_2740 &  n_4413;
assign n_5083 = ~n_5081 & ~n_5082;
assign n_5084 = ~x_2733 &  n_4387;
assign n_5085 = ~x_2736 &  n_4403;
assign n_5086 = ~n_5084 & ~n_5085;
assign n_5087 =  n_5083 &  n_5086;
assign n_5088 = ~x_2743 &  n_4379;
assign n_5089 = ~x_2746 &  n_4397;
assign n_5090 = ~n_5088 & ~n_5089;
assign n_5091 = ~x_2748 &  n_4415;
assign n_5092 = ~x_2737 &  n_4424;
assign n_5093 = ~n_5091 & ~n_5092;
assign n_5094 =  n_5090 &  n_5093;
assign n_5095 =  n_5087 &  n_5094;
assign n_5096 = ~x_2747 &  n_4389;
assign n_5097 = ~x_2744 &  n_4426;
assign n_5098 = ~n_5096 & ~n_5097;
assign n_5099 = ~x_2734 &  n_4395;
assign n_5100 = ~x_2739 &  n_4421;
assign n_5101 = ~n_5099 & ~n_5100;
assign n_5102 =  n_5098 &  n_5101;
assign n_5103 = ~x_2741 &  n_4383;
assign n_5104 = ~x_2735 &  n_4410;
assign n_5105 = ~n_5103 & ~n_5104;
assign n_5106 = ~x_2738 &  n_4408;
assign n_5107 = ~x_2745 &  n_4419;
assign n_5108 = ~n_5106 & ~n_5107;
assign n_5109 =  n_5105 &  n_5108;
assign n_5110 =  n_5102 &  n_5109;
assign n_5111 =  n_5095 &  n_5110;
assign n_5112 =  x_1519 & ~n_5111;
assign n_5113 = ~x_1519 &  n_5111;
assign n_5114 = ~n_5112 & ~n_5113;
assign n_5115 = ~x_2718 &  n_4395;
assign n_5116 = ~x_2721 &  n_4424;
assign n_5117 = ~n_5115 & ~n_5116;
assign n_5118 = ~x_2717 &  n_4387;
assign n_5119 = ~x_2730 &  n_4397;
assign n_5120 = ~n_5118 & ~n_5119;
assign n_5121 =  n_5117 &  n_5120;
assign n_5122 = ~x_2731 &  n_4389;
assign n_5123 = ~x_2719 &  n_4410;
assign n_5124 = ~n_5122 & ~n_5123;
assign n_5125 = ~x_2724 &  n_4413;
assign n_5126 = ~x_2728 &  n_4426;
assign n_5127 = ~n_5125 & ~n_5126;
assign n_5128 =  n_5124 &  n_5127;
assign n_5129 =  n_5121 &  n_5128;
assign n_5130 = ~x_2727 &  n_4379;
assign n_5131 = ~x_2722 &  n_4408;
assign n_5132 = ~n_5130 & ~n_5131;
assign n_5133 = ~x_2726 &  n_4400;
assign n_5134 = ~x_2729 &  n_4419;
assign n_5135 = ~n_5133 & ~n_5134;
assign n_5136 =  n_5132 &  n_5135;
assign n_5137 = ~x_2732 &  n_4415;
assign n_5138 = ~x_2723 &  n_4421;
assign n_5139 = ~n_5137 & ~n_5138;
assign n_5140 = ~x_2725 &  n_4383;
assign n_5141 = ~x_2720 &  n_4403;
assign n_5142 = ~n_5140 & ~n_5141;
assign n_5143 =  n_5139 &  n_5142;
assign n_5144 =  n_5136 &  n_5143;
assign n_5145 =  n_5129 &  n_5144;
assign n_5146 =  x_1520 & ~n_5145;
assign n_5147 = ~x_1520 &  n_5145;
assign n_5148 = ~n_5146 & ~n_5147;
assign n_5149 = ~x_2709 &  n_4383;
assign n_5150 = ~x_2706 &  n_4408;
assign n_5151 = ~n_5149 & ~n_5150;
assign n_5152 = ~x_2701 &  n_4387;
assign n_5153 = ~x_2711 &  n_4379;
assign n_5154 = ~n_5152 & ~n_5153;
assign n_5155 =  n_5151 &  n_5154;
assign n_5156 = ~x_2702 &  n_4395;
assign n_5157 = ~x_2703 &  n_4410;
assign n_5158 = ~n_5156 & ~n_5157;
assign n_5159 = ~x_2712 &  n_4426;
assign n_5160 = ~x_2708 &  n_4413;
assign n_5161 = ~n_5159 & ~n_5160;
assign n_5162 =  n_5158 &  n_5161;
assign n_5163 =  n_5155 &  n_5162;
assign n_5164 = ~x_2714 &  n_4397;
assign n_5165 = ~x_2715 &  n_4389;
assign n_5166 = ~n_5164 & ~n_5165;
assign n_5167 = ~x_2705 &  n_4424;
assign n_5168 = ~x_2710 &  n_4400;
assign n_5169 = ~n_5167 & ~n_5168;
assign n_5170 =  n_5166 &  n_5169;
assign n_5171 = ~x_2704 &  n_4403;
assign n_5172 = ~x_2707 &  n_4421;
assign n_5173 = ~n_5171 & ~n_5172;
assign n_5174 = ~x_2713 &  n_4419;
assign n_5175 = ~x_2716 &  n_4415;
assign n_5176 = ~n_5174 & ~n_5175;
assign n_5177 =  n_5173 &  n_5176;
assign n_5178 =  n_5170 &  n_5177;
assign n_5179 =  n_5163 &  n_5178;
assign n_5180 =  x_1521 & ~n_5179;
assign n_5181 = ~x_1521 &  n_5179;
assign n_5182 = ~n_5180 & ~n_5181;
assign n_5183 = ~x_2689 &  n_4424;
assign n_5184 = ~x_2700 &  n_4415;
assign n_5185 = ~n_5183 & ~n_5184;
assign n_5186 = ~x_2685 &  n_4387;
assign n_5187 = ~x_2691 &  n_4421;
assign n_5188 = ~n_5186 & ~n_5187;
assign n_5189 =  n_5185 &  n_5188;
assign n_5190 = ~x_2699 &  n_4389;
assign n_5191 = ~x_2687 &  n_4410;
assign n_5192 = ~n_5190 & ~n_5191;
assign n_5193 = ~x_2694 &  n_4400;
assign n_5194 = ~x_2690 &  n_4408;
assign n_5195 = ~n_5193 & ~n_5194;
assign n_5196 =  n_5192 &  n_5195;
assign n_5197 =  n_5189 &  n_5196;
assign n_5198 = ~x_2697 &  n_4419;
assign n_5199 = ~x_2686 &  n_4395;
assign n_5200 = ~n_5198 & ~n_5199;
assign n_5201 = ~x_2688 &  n_4403;
assign n_5202 = ~x_2696 &  n_4426;
assign n_5203 = ~n_5201 & ~n_5202;
assign n_5204 =  n_5200 &  n_5203;
assign n_5205 = ~x_2692 &  n_4413;
assign n_5206 = ~x_2698 &  n_4397;
assign n_5207 = ~n_5205 & ~n_5206;
assign n_5208 = ~x_2695 &  n_4379;
assign n_5209 = ~x_2693 &  n_4383;
assign n_5210 = ~n_5208 & ~n_5209;
assign n_5211 =  n_5207 &  n_5210;
assign n_5212 =  n_5204 &  n_5211;
assign n_5213 =  n_5197 &  n_5212;
assign n_5214 =  x_1522 & ~n_5213;
assign n_5215 = ~x_1522 &  n_5213;
assign n_5216 = ~n_5214 & ~n_5215;
assign n_5217 = ~x_2675 &  n_4421;
assign n_5218 = ~x_2680 &  n_4426;
assign n_5219 = ~n_5217 & ~n_5218;
assign n_5220 = ~x_2669 &  n_4387;
assign n_5221 = ~x_2673 &  n_4424;
assign n_5222 = ~n_5220 & ~n_5221;
assign n_5223 =  n_5219 &  n_5222;
assign n_5224 = ~x_2678 &  n_4400;
assign n_5225 = ~x_2674 &  n_4408;
assign n_5226 = ~n_5224 & ~n_5225;
assign n_5227 = ~x_2671 &  n_4410;
assign n_5228 = ~x_2672 &  n_4403;
assign n_5229 = ~n_5227 & ~n_5228;
assign n_5230 =  n_5226 &  n_5229;
assign n_5231 =  n_5223 &  n_5230;
assign n_5232 = ~x_2682 &  n_4397;
assign n_5233 = ~x_2683 &  n_4389;
assign n_5234 = ~n_5232 & ~n_5233;
assign n_5235 = ~x_2670 &  n_4395;
assign n_5236 = ~x_2676 &  n_4413;
assign n_5237 = ~n_5235 & ~n_5236;
assign n_5238 =  n_5234 &  n_5237;
assign n_5239 = ~x_2681 &  n_4419;
assign n_5240 = ~x_2679 &  n_4379;
assign n_5241 = ~n_5239 & ~n_5240;
assign n_5242 = ~x_2677 &  n_4383;
assign n_5243 = ~x_2684 &  n_4415;
assign n_5244 = ~n_5242 & ~n_5243;
assign n_5245 =  n_5241 &  n_5244;
assign n_5246 =  n_5238 &  n_5245;
assign n_5247 =  n_5231 &  n_5246;
assign n_5248 =  x_1523 & ~n_5247;
assign n_5249 = ~x_1523 &  n_5247;
assign n_5250 = ~n_5248 & ~n_5249;
assign n_5251 = ~x_2659 &  n_4421;
assign n_5252 = ~x_2660 &  n_4413;
assign n_5253 = ~n_5251 & ~n_5252;
assign n_5254 = ~x_2653 &  n_4387;
assign n_5255 = ~x_2668 &  n_4415;
assign n_5256 = ~n_5254 & ~n_5255;
assign n_5257 =  n_5253 &  n_5256;
assign n_5258 = ~x_2657 &  n_4424;
assign n_5259 = ~x_2667 &  n_4389;
assign n_5260 = ~n_5258 & ~n_5259;
assign n_5261 = ~x_2666 &  n_4397;
assign n_5262 = ~x_2661 &  n_4383;
assign n_5263 = ~n_5261 & ~n_5262;
assign n_5264 =  n_5260 &  n_5263;
assign n_5265 =  n_5257 &  n_5264;
assign n_5266 = ~x_2658 &  n_4408;
assign n_5267 = ~x_2662 &  n_4400;
assign n_5268 = ~n_5266 & ~n_5267;
assign n_5269 = ~x_2655 &  n_4410;
assign n_5270 = ~x_2656 &  n_4403;
assign n_5271 = ~n_5269 & ~n_5270;
assign n_5272 =  n_5268 &  n_5271;
assign n_5273 = ~x_2664 &  n_4426;
assign n_5274 = ~x_2654 &  n_4395;
assign n_5275 = ~n_5273 & ~n_5274;
assign n_5276 = ~x_2663 &  n_4379;
assign n_5277 = ~x_2665 &  n_4419;
assign n_5278 = ~n_5276 & ~n_5277;
assign n_5279 =  n_5275 &  n_5278;
assign n_5280 =  n_5272 &  n_5279;
assign n_5281 =  n_5265 &  n_5280;
assign n_5282 =  x_1524 & ~n_5281;
assign n_5283 = ~x_1524 &  n_5281;
assign n_5284 = ~n_5282 & ~n_5283;
assign n_5285 = ~x_2645 &  n_4383;
assign n_5286 = ~x_2640 &  n_4403;
assign n_5287 = ~n_5285 & ~n_5286;
assign n_5288 = ~x_2637 &  n_4387;
assign n_5289 = ~x_2642 &  n_4408;
assign n_5290 = ~n_5288 & ~n_5289;
assign n_5291 =  n_5287 &  n_5290;
assign n_5292 = ~x_2643 &  n_4421;
assign n_5293 = ~x_2639 &  n_4410;
assign n_5294 = ~n_5292 & ~n_5293;
assign n_5295 = ~x_2649 &  n_4419;
assign n_5296 = ~x_2651 &  n_4389;
assign n_5297 = ~n_5295 & ~n_5296;
assign n_5298 =  n_5294 &  n_5297;
assign n_5299 =  n_5291 &  n_5298;
assign n_5300 = ~x_2647 &  n_4379;
assign n_5301 = ~x_2650 &  n_4397;
assign n_5302 = ~n_5300 & ~n_5301;
assign n_5303 = ~x_2648 &  n_4426;
assign n_5304 = ~x_2641 &  n_4424;
assign n_5305 = ~n_5303 & ~n_5304;
assign n_5306 =  n_5302 &  n_5305;
assign n_5307 = ~x_2652 &  n_4415;
assign n_5308 = ~x_2638 &  n_4395;
assign n_5309 = ~n_5307 & ~n_5308;
assign n_5310 = ~x_2644 &  n_4413;
assign n_5311 = ~x_2646 &  n_4400;
assign n_5312 = ~n_5310 & ~n_5311;
assign n_5313 =  n_5309 &  n_5312;
assign n_5314 =  n_5306 &  n_5313;
assign n_5315 =  n_5299 &  n_5314;
assign n_5316 =  x_1525 & ~n_5315;
assign n_5317 = ~x_1525 &  n_5315;
assign n_5318 = ~n_5316 & ~n_5317;
assign n_5319 = ~x_2622 &  n_4395;
assign n_5320 = ~x_2628 &  n_4413;
assign n_5321 = ~n_5319 & ~n_5320;
assign n_5322 = ~x_2621 &  n_4387;
assign n_5323 = ~x_2631 &  n_4379;
assign n_5324 = ~n_5322 & ~n_5323;
assign n_5325 =  n_5321 &  n_5324;
assign n_5326 = ~x_2627 &  n_4421;
assign n_5327 = ~x_2633 &  n_4419;
assign n_5328 = ~n_5326 & ~n_5327;
assign n_5329 = ~x_2630 &  n_4400;
assign n_5330 = ~x_2624 &  n_4403;
assign n_5331 = ~n_5329 & ~n_5330;
assign n_5332 =  n_5328 &  n_5331;
assign n_5333 =  n_5325 &  n_5332;
assign n_5334 = ~x_2634 &  n_4397;
assign n_5335 = ~x_2626 &  n_4408;
assign n_5336 = ~n_5334 & ~n_5335;
assign n_5337 = ~x_2625 &  n_4424;
assign n_5338 = ~x_2623 &  n_4410;
assign n_5339 = ~n_5337 & ~n_5338;
assign n_5340 =  n_5336 &  n_5339;
assign n_5341 = ~x_2629 &  n_4383;
assign n_5342 = ~x_2635 &  n_4389;
assign n_5343 = ~n_5341 & ~n_5342;
assign n_5344 = ~x_2636 &  n_4415;
assign n_5345 = ~x_2632 &  n_4426;
assign n_5346 = ~n_5344 & ~n_5345;
assign n_5347 =  n_5343 &  n_5346;
assign n_5348 =  n_5340 &  n_5347;
assign n_5349 =  n_5333 &  n_5348;
assign n_5350 =  x_1526 & ~n_5349;
assign n_5351 = ~x_1526 &  n_5349;
assign n_5352 = ~n_5350 & ~n_5351;
assign n_5353 = ~x_2615 &  n_4379;
assign n_5354 = ~x_2608 &  n_4403;
assign n_5355 = ~n_5353 & ~n_5354;
assign n_5356 = ~x_2605 &  n_4387;
assign n_5357 = ~x_2609 &  n_4424;
assign n_5358 = ~n_5356 & ~n_5357;
assign n_5359 =  n_5355 &  n_5358;
assign n_5360 = ~x_2617 &  n_4419;
assign n_5361 = ~x_2614 &  n_4400;
assign n_5362 = ~n_5360 & ~n_5361;
assign n_5363 = ~x_2611 &  n_4421;
assign n_5364 = ~x_2612 &  n_4413;
assign n_5365 = ~n_5363 & ~n_5364;
assign n_5366 =  n_5362 &  n_5365;
assign n_5367 =  n_5359 &  n_5366;
assign n_5368 = ~x_2618 &  n_4397;
assign n_5369 = ~x_2607 &  n_4410;
assign n_5370 = ~n_5368 & ~n_5369;
assign n_5371 = ~x_2610 &  n_4408;
assign n_5372 = ~x_2620 &  n_4415;
assign n_5373 = ~n_5371 & ~n_5372;
assign n_5374 =  n_5370 &  n_5373;
assign n_5375 = ~x_2616 &  n_4426;
assign n_5376 = ~x_2619 &  n_4389;
assign n_5377 = ~n_5375 & ~n_5376;
assign n_5378 = ~x_2606 &  n_4395;
assign n_5379 = ~x_2613 &  n_4383;
assign n_5380 = ~n_5378 & ~n_5379;
assign n_5381 =  n_5377 &  n_5380;
assign n_5382 =  n_5374 &  n_5381;
assign n_5383 =  n_5367 &  n_5382;
assign n_5384 =  x_1527 & ~n_5383;
assign n_5385 = ~x_2589 &  n_4387;
assign n_5386 = ~x_2594 &  n_4408;
assign n_5387 = ~n_5385 & ~n_5386;
assign n_5388 = ~x_2596 &  n_4413;
assign n_5389 = ~x_2603 &  n_4389;
assign n_5390 = ~n_5388 & ~n_5389;
assign n_5391 =  n_5387 &  n_5390;
assign n_5392 = ~x_2600 &  n_4426;
assign n_5393 = ~x_2599 &  n_4379;
assign n_5394 = ~n_5392 & ~n_5393;
assign n_5395 = ~x_2593 &  n_4424;
assign n_5396 = ~x_2592 &  n_4403;
assign n_5397 = ~n_5395 & ~n_5396;
assign n_5398 =  n_5394 &  n_5397;
assign n_5399 =  n_5391 &  n_5398;
assign n_5400 = ~x_2604 &  n_4415;
assign n_5401 = ~x_2602 &  n_4397;
assign n_5402 = ~n_5400 & ~n_5401;
assign n_5403 = ~x_2597 &  n_4383;
assign n_5404 = ~x_2601 &  n_4419;
assign n_5405 = ~n_5403 & ~n_5404;
assign n_5406 =  n_5402 &  n_5405;
assign n_5407 = ~x_2595 &  n_4421;
assign n_5408 = ~x_2598 &  n_4400;
assign n_5409 = ~n_5407 & ~n_5408;
assign n_5410 = ~x_2591 &  n_4410;
assign n_5411 = ~x_2590 &  n_4395;
assign n_5412 = ~n_5410 & ~n_5411;
assign n_5413 =  n_5409 &  n_5412;
assign n_5414 =  n_5406 &  n_5413;
assign n_5415 =  n_5399 &  n_5414;
assign n_5416 =  x_1528 & ~n_5415;
assign n_5417 = ~x_1528 &  n_5415;
assign n_5418 = ~x_2559 &  n_4410;
assign n_5419 = ~x_1530 & ~n_5418;
assign n_5420 = ~x_2569 &  n_4419;
assign n_5421 = ~x_2570 &  n_4397;
assign n_5422 = ~n_5420 & ~n_5421;
assign n_5423 = ~x_2557 &  n_4387;
assign n_5424 = ~x_2572 &  n_4415;
assign n_5425 = ~n_5423 & ~n_5424;
assign n_5426 =  n_5422 &  n_5425;
assign n_5427 =  n_5419 &  n_5426;
assign n_5428 = ~x_2563 &  n_4421;
assign n_5429 = ~x_2566 &  n_4400;
assign n_5430 = ~x_2561 &  n_4424;
assign n_5431 = ~n_5429 & ~n_5430;
assign n_5432 = ~n_5428 &  n_5431;
assign n_5433 = ~x_2564 &  n_4413;
assign n_5434 = ~x_2558 &  n_4395;
assign n_5435 = ~n_5433 & ~n_5434;
assign n_5436 = ~x_2560 &  n_4403;
assign n_5437 = ~x_2571 &  n_4389;
assign n_5438 = ~n_5436 & ~n_5437;
assign n_5439 =  n_5435 &  n_5438;
assign n_5440 = ~x_2567 &  n_4379;
assign n_5441 = ~x_2568 &  n_4426;
assign n_5442 = ~n_5440 & ~n_5441;
assign n_5443 = ~x_2565 &  n_4383;
assign n_5444 = ~x_2562 &  n_4408;
assign n_5445 = ~n_5443 & ~n_5444;
assign n_5446 =  n_5442 &  n_5445;
assign n_5447 =  n_5439 &  n_5446;
assign n_5448 =  n_5432 &  n_5447;
assign n_5449 =  n_5427 &  n_5448;
assign n_5450 = ~x_1529 &  n_5449;
assign n_5451 = ~x_2573 &  n_4387;
assign n_5452 = ~x_2575 &  n_4410;
assign n_5453 = ~n_5451 & ~n_5452;
assign n_5454 = ~x_2587 &  n_4389;
assign n_5455 = ~x_2581 &  n_4383;
assign n_5456 = ~n_5454 & ~n_5455;
assign n_5457 =  n_5453 &  n_5456;
assign n_5458 = ~x_2582 &  n_4400;
assign n_5459 = ~x_2578 &  n_4408;
assign n_5460 = ~n_5458 & ~n_5459;
assign n_5461 = ~x_2576 &  n_4403;
assign n_5462 = ~x_2588 &  n_4415;
assign n_5463 = ~n_5461 & ~n_5462;
assign n_5464 =  n_5460 &  n_5463;
assign n_5465 =  n_5457 &  n_5464;
assign n_5466 = ~x_2586 &  n_4397;
assign n_5467 = ~x_2574 &  n_4395;
assign n_5468 = ~n_5466 & ~n_5467;
assign n_5469 = ~x_2580 &  n_4413;
assign n_5470 = ~x_2585 &  n_4419;
assign n_5471 = ~n_5469 & ~n_5470;
assign n_5472 =  n_5468 &  n_5471;
assign n_5473 = ~x_2583 &  n_4379;
assign n_5474 = ~x_2579 &  n_4421;
assign n_5475 = ~n_5473 & ~n_5474;
assign n_5476 = ~x_2577 &  n_4424;
assign n_5477 = ~x_2584 &  n_4426;
assign n_5478 = ~n_5476 & ~n_5477;
assign n_5479 =  n_5475 &  n_5478;
assign n_5480 =  n_5472 &  n_5479;
assign n_5481 =  n_5465 &  n_5480;
assign n_5482 = ~n_5450 & ~n_5481;
assign n_5483 =  x_1529 & ~n_5449;
assign n_5484 = ~n_5482 & ~n_5483;
assign n_5485 = ~n_5417 & ~n_5484;
assign n_5486 = ~n_5416 & ~n_5485;
assign n_5487 = ~x_1527 &  n_5383;
assign n_5488 = ~n_5384 & ~n_5487;
assign n_5489 = ~n_5486 &  n_5488;
assign n_5490 = ~n_5384 & ~n_5489;
assign n_5491 =  n_5352 & ~n_5490;
assign n_5492 = ~n_5350 & ~n_5491;
assign n_5493 =  n_5318 & ~n_5492;
assign n_5494 = ~n_5316 & ~n_5493;
assign n_5495 =  n_5284 & ~n_5494;
assign n_5496 = ~n_5282 & ~n_5495;
assign n_5497 =  n_5250 & ~n_5496;
assign n_5498 = ~n_5248 & ~n_5497;
assign n_5499 =  n_5216 & ~n_5498;
assign n_5500 = ~n_5214 & ~n_5499;
assign n_5501 =  n_5182 & ~n_5500;
assign n_5502 = ~n_5180 & ~n_5501;
assign n_5503 =  n_5148 & ~n_5502;
assign n_5504 = ~n_5146 & ~n_5503;
assign n_5505 =  n_5114 & ~n_5504;
assign n_5506 = ~n_5112 & ~n_5505;
assign n_5507 =  n_5080 & ~n_5506;
assign n_5508 = ~n_5078 & ~n_5507;
assign n_5509 =  n_5046 & ~n_5508;
assign n_5510 = ~n_5044 & ~n_5509;
assign n_5511 =  n_5012 & ~n_5510;
assign n_5512 = ~n_5010 & ~n_5511;
assign n_5513 =  n_4978 & ~n_5512;
assign n_5514 = ~n_4976 & ~n_5513;
assign n_5515 =  n_4944 & ~n_5514;
assign n_5516 = ~n_4942 & ~n_5515;
assign n_5517 =  n_4910 & ~n_5516;
assign n_5518 = ~n_4908 & ~n_5517;
assign n_5519 =  n_4876 & ~n_5518;
assign n_5520 = ~n_4874 & ~n_5519;
assign n_5521 =  n_4842 & ~n_5520;
assign n_5522 = ~n_4840 & ~n_5521;
assign n_5523 =  n_4808 & ~n_5522;
assign n_5524 = ~n_4806 & ~n_5523;
assign n_5525 =  n_4774 & ~n_5524;
assign n_5526 = ~n_4772 & ~n_5525;
assign n_5527 =  n_4740 & ~n_5526;
assign n_5528 = ~n_4738 & ~n_5527;
assign n_5529 =  n_4706 & ~n_5528;
assign n_5530 = ~n_4704 & ~n_5529;
assign n_5531 =  n_4672 & ~n_5530;
assign n_5532 = ~n_4670 & ~n_5531;
assign n_5533 =  n_4638 & ~n_5532;
assign n_5534 = ~n_4636 & ~n_5533;
assign n_5535 =  n_4604 & ~n_5534;
assign n_5536 = ~n_4602 & ~n_5535;
assign n_5537 =  n_4570 & ~n_5536;
assign n_5538 = ~n_4568 & ~n_5537;
assign n_5539 =  n_4536 & ~n_5538;
assign n_5540 = ~n_4534 & ~n_5539;
assign n_5541 =  n_4502 & ~n_5540;
assign n_5542 = ~n_4500 & ~n_5541;
assign n_5543 =  n_4468 & ~n_5542;
assign n_5544 = ~n_4466 & ~n_5543;
assign n_5545 =  n_4434 & ~n_5544;
assign n_5546 = ~n_4434 &  n_5544;
assign n_5547 = ~n_4375 & ~n_5546;
assign n_5548 = ~n_5545 &  n_5547;
assign n_5549 = ~n_4376 & ~n_5548;
assign n_5550 =  x_1561 &  n_4375;
assign n_5551 = ~n_4468 &  n_5542;
assign n_5552 = ~n_4375 & ~n_5543;
assign n_5553 = ~n_5551 &  n_5552;
assign n_5554 = ~n_5550 & ~n_5553;
assign n_5555 =  x_1500 &  n_4375;
assign n_5556 = ~n_4502 &  n_5540;
assign n_5557 = ~n_4375 & ~n_5556;
assign n_5558 = ~n_5541 &  n_5557;
assign n_5559 = ~n_5555 & ~n_5558;
assign n_5560 =  x_1554 &  n_4375;
assign n_5561 = ~n_4536 &  n_5538;
assign n_5562 = ~n_4375 & ~n_5539;
assign n_5563 = ~n_5561 &  n_5562;
assign n_5564 = ~n_5560 & ~n_5563;
assign n_5565 =  x_1531 &  n_4375;
assign n_5566 = ~n_4570 &  n_5536;
assign n_5567 = ~n_4375 & ~n_5537;
assign n_5568 = ~n_5566 &  n_5567;
assign n_5569 = ~n_5565 & ~n_5568;
assign n_5570 =  x_1532 &  n_4375;
assign n_5571 = ~n_4604 &  n_5534;
assign n_5572 = ~n_4375 & ~n_5535;
assign n_5573 = ~n_5571 &  n_5572;
assign n_5574 = ~n_5570 & ~n_5573;
assign n_5575 =  x_1553 &  n_4375;
assign n_5576 = ~n_4638 &  n_5532;
assign n_5577 = ~n_4375 & ~n_5533;
assign n_5578 = ~n_5576 &  n_5577;
assign n_5579 = ~n_5575 & ~n_5578;
assign n_5580 =  x_1552 &  n_4375;
assign n_5581 = ~n_4672 &  n_5530;
assign n_5582 = ~n_4375 & ~n_5531;
assign n_5583 = ~n_5581 &  n_5582;
assign n_5584 = ~n_5580 & ~n_5583;
assign n_5585 =  x_1533 &  n_4375;
assign n_5586 = ~n_4706 &  n_5528;
assign n_5587 = ~n_4375 & ~n_5529;
assign n_5588 = ~n_5586 &  n_5587;
assign n_5589 = ~n_5585 & ~n_5588;
assign n_5590 =  x_1536 &  n_4375;
assign n_5591 = ~n_4740 &  n_5526;
assign n_5592 = ~n_4375 & ~n_5527;
assign n_5593 = ~n_5591 &  n_5592;
assign n_5594 = ~n_5590 & ~n_5593;
assign n_5595 =  x_1550 &  n_4375;
assign n_5596 = ~n_4774 &  n_5524;
assign n_5597 = ~n_4375 & ~n_5525;
assign n_5598 = ~n_5596 &  n_5597;
assign n_5599 = ~n_5595 & ~n_5598;
assign n_5600 =  x_1551 &  n_4375;
assign n_5601 = ~n_4808 &  n_5522;
assign n_5602 = ~n_4375 & ~n_5523;
assign n_5603 = ~n_5601 &  n_5602;
assign n_5604 = ~n_5600 & ~n_5603;
assign n_5605 =  x_1535 &  n_4375;
assign n_5606 = ~n_4842 &  n_5520;
assign n_5607 = ~n_4375 & ~n_5521;
assign n_5608 = ~n_5606 &  n_5607;
assign n_5609 = ~n_5605 & ~n_5608;
assign n_5610 =  x_1537 &  n_4375;
assign n_5611 = ~n_4876 &  n_5518;
assign n_5612 = ~n_4375 & ~n_5519;
assign n_5613 = ~n_5611 &  n_5612;
assign n_5614 = ~n_5610 & ~n_5613;
assign n_5615 =  x_1534 &  n_4375;
assign n_5616 = ~n_4910 &  n_5516;
assign n_5617 = ~n_4375 & ~n_5517;
assign n_5618 = ~n_5616 &  n_5617;
assign n_5619 = ~n_5615 & ~n_5618;
assign n_5620 =  x_1560 &  n_4375;
assign n_5621 = ~n_4944 &  n_5514;
assign n_5622 = ~n_4375 & ~n_5515;
assign n_5623 = ~n_5621 &  n_5622;
assign n_5624 = ~n_5620 & ~n_5623;
assign n_5625 =  x_1545 &  n_4375;
assign n_5626 = ~n_4978 &  n_5512;
assign n_5627 = ~n_4375 & ~n_5513;
assign n_5628 = ~n_5626 &  n_5627;
assign n_5629 = ~n_5625 & ~n_5628;
assign n_5630 =  x_1546 &  n_4375;
assign n_5631 = ~n_5012 &  n_5510;
assign n_5632 = ~n_4375 & ~n_5511;
assign n_5633 = ~n_5631 &  n_5632;
assign n_5634 = ~n_5630 & ~n_5633;
assign n_5635 =  x_1540 &  n_4375;
assign n_5636 = ~n_5046 &  n_5508;
assign n_5637 = ~n_4375 & ~n_5509;
assign n_5638 = ~n_5636 &  n_5637;
assign n_5639 = ~n_5635 & ~n_5638;
assign n_5640 =  x_1547 &  n_4375;
assign n_5641 = ~n_5080 &  n_5506;
assign n_5642 = ~n_4375 & ~n_5507;
assign n_5643 = ~n_5641 &  n_5642;
assign n_5644 = ~n_5640 & ~n_5643;
assign n_5645 =  x_1549 &  n_4375;
assign n_5646 = ~n_5114 &  n_5504;
assign n_5647 = ~n_4375 & ~n_5505;
assign n_5648 = ~n_5646 &  n_5647;
assign n_5649 = ~n_5645 & ~n_5648;
assign n_5650 =  x_1541 &  n_4375;
assign n_5651 = ~n_5148 &  n_5502;
assign n_5652 = ~n_4375 & ~n_5503;
assign n_5653 = ~n_5651 &  n_5652;
assign n_5654 = ~n_5650 & ~n_5653;
assign n_5655 =  x_1544 &  n_4375;
assign n_5656 = ~n_5182 &  n_5500;
assign n_5657 = ~n_4375 & ~n_5501;
assign n_5658 = ~n_5656 &  n_5657;
assign n_5659 = ~n_5655 & ~n_5658;
assign n_5660 =  x_1539 &  n_4375;
assign n_5661 = ~n_5216 &  n_5498;
assign n_5662 = ~n_4375 & ~n_5499;
assign n_5663 = ~n_5661 &  n_5662;
assign n_5664 = ~n_5660 & ~n_5663;
assign n_5665 =  x_1538 &  n_4375;
assign n_5666 = ~n_5250 &  n_5496;
assign n_5667 = ~n_4375 & ~n_5497;
assign n_5668 = ~n_5666 &  n_5667;
assign n_5669 = ~n_5665 & ~n_5668;
assign n_5670 =  x_1543 &  n_4375;
assign n_5671 = ~n_5284 &  n_5494;
assign n_5672 = ~n_4375 & ~n_5495;
assign n_5673 = ~n_5671 &  n_5672;
assign n_5674 = ~n_5670 & ~n_5673;
assign n_5675 =  x_1542 &  n_4375;
assign n_5676 = ~n_5318 &  n_5492;
assign n_5677 = ~n_4375 & ~n_5493;
assign n_5678 = ~n_5676 &  n_5677;
assign n_5679 = ~n_5675 & ~n_5678;
assign n_5680 =  x_1556 &  n_4375;
assign n_5681 = ~n_5352 &  n_5490;
assign n_5682 = ~n_4375 & ~n_5491;
assign n_5683 = ~n_5681 &  n_5682;
assign n_5684 = ~n_5680 & ~n_5683;
assign n_5685 =  x_1548 &  n_4375;
assign n_5686 = ~n_5416 & ~n_5417;
assign n_5687 = ~n_5484 &  n_5686;
assign n_5688 =  n_5484 & ~n_5686;
assign n_5689 = ~n_4375 & ~n_5688;
assign n_5690 = ~n_5687 &  n_5689;
assign n_5691 = ~n_5685 & ~n_5690;
assign n_5692 =  x_1555 &  n_4375;
assign n_5693 =  n_5486 & ~n_5488;
assign n_5694 = ~n_4375 & ~n_5489;
assign n_5695 = ~n_5693 &  n_5694;
assign n_5696 = ~n_5692 & ~n_5695;
assign n_5697 =  n_5691 &  n_5696;
assign n_5698 =  n_5684 &  n_5697;
assign n_5699 =  n_5679 &  n_5698;
assign n_5700 =  n_5674 &  n_5699;
assign n_5701 =  n_5669 &  n_5700;
assign n_5702 =  n_5664 &  n_5701;
assign n_5703 =  n_5659 &  n_5702;
assign n_5704 =  n_5654 &  n_5703;
assign n_5705 =  n_5649 &  n_5704;
assign n_5706 =  n_5644 &  n_5705;
assign n_5707 =  n_5639 &  n_5706;
assign n_5708 =  n_5634 &  n_5707;
assign n_5709 =  n_5629 &  n_5708;
assign n_5710 =  n_5624 &  n_5709;
assign n_5711 =  n_5619 &  n_5710;
assign n_5712 =  n_5614 &  n_5711;
assign n_5713 =  n_5609 &  n_5712;
assign n_5714 =  n_5604 &  n_5713;
assign n_5715 =  n_5599 &  n_5714;
assign n_5716 =  n_5594 &  n_5715;
assign n_5717 =  n_5589 &  n_5716;
assign n_5718 =  n_5584 &  n_5717;
assign n_5719 =  n_5579 &  n_5718;
assign n_5720 =  n_5574 &  n_5719;
assign n_5721 =  n_5569 &  n_5720;
assign n_5722 =  n_5564 &  n_5721;
assign n_5723 =  n_5559 &  n_5722;
assign n_5724 =  n_5554 &  n_5723;
assign n_5725 =  n_5549 &  n_5724;
assign n_5726 =  x_1466 &  n_1522;
assign n_5727 = ~x_1467 & ~n_1525;
assign n_5728 = ~n_5726 &  n_5727;
assign n_5729 = ~n_4374 & ~n_5728;
assign n_5730 = ~n_5725 &  n_5729;
assign n_5731 = ~n_3617 & ~n_3634;
assign n_5732 = ~x_2421 & ~x_2422;
assign n_5733 = ~x_2423 & ~x_2424;
assign n_5734 =  n_5732 &  n_5733;
assign n_5735 = ~x_2417 & ~x_2418;
assign n_5736 = ~x_2419 & ~x_2420;
assign n_5737 =  n_5735 &  n_5736;
assign n_5738 =  n_5734 &  n_5737;
assign n_5739 = ~x_2429 & ~x_2430;
assign n_5740 = ~x_2431 & ~x_2432;
assign n_5741 =  n_5739 &  n_5740;
assign n_5742 = ~x_2425 & ~x_2426;
assign n_5743 = ~x_2427 & ~x_2428;
assign n_5744 =  n_5742 &  n_5743;
assign n_5745 =  n_5741 &  n_5744;
assign n_5746 =  n_5738 &  n_5745;
assign n_5747 = ~x_2405 & ~x_2406;
assign n_5748 = ~x_2407 & ~x_2408;
assign n_5749 =  n_5747 &  n_5748;
assign n_5750 = ~x_2403 & ~x_2404;
assign n_5751 =  n_3660 &  n_5750;
assign n_5752 =  n_5749 &  n_5751;
assign n_5753 = ~x_2413 & ~x_2414;
assign n_5754 = ~x_2415 & ~x_2416;
assign n_5755 =  n_5753 &  n_5754;
assign n_5756 = ~x_2409 & ~x_2410;
assign n_5757 = ~x_2411 & ~x_2412;
assign n_5758 =  n_5756 &  n_5757;
assign n_5759 =  n_5755 &  n_5758;
assign n_5760 =  n_5752 &  n_5759;
assign n_5761 =  n_5746 &  n_5760;
assign n_5762 =  n_3645 & ~n_5761;
assign n_5763 = ~x_2388 & ~x_2389;
assign n_5764 = ~x_2390 & ~x_2391;
assign n_5765 =  n_5763 &  n_5764;
assign n_5766 = ~x_2384 & ~x_2385;
assign n_5767 = ~x_2386 & ~x_2387;
assign n_5768 =  n_5766 &  n_5767;
assign n_5769 =  n_5765 &  n_5768;
assign n_5770 = ~x_2396 & ~x_2397;
assign n_5771 = ~x_2398 &  n_5770;
assign n_5772 = ~x_2392 & ~x_2393;
assign n_5773 = ~x_2394 & ~x_2395;
assign n_5774 =  n_5772 &  n_5773;
assign n_5775 =  n_5771 &  n_5774;
assign n_5776 =  n_5769 &  n_5775;
assign n_5777 = ~x_2372 & ~x_2373;
assign n_5778 = ~x_2374 & ~x_2375;
assign n_5779 =  n_5777 &  n_5778;
assign n_5780 = ~x_2368 & ~x_2369;
assign n_5781 = ~x_2370 & ~x_2371;
assign n_5782 =  n_5780 &  n_5781;
assign n_5783 =  n_5779 &  n_5782;
assign n_5784 = ~x_2380 & ~x_2381;
assign n_5785 = ~x_2382 & ~x_2383;
assign n_5786 =  n_5784 &  n_5785;
assign n_5787 = ~x_2376 & ~x_2377;
assign n_5788 = ~x_2378 & ~x_2379;
assign n_5789 =  n_5787 &  n_5788;
assign n_5790 =  n_5786 &  n_5789;
assign n_5791 =  n_5783 &  n_5790;
assign n_5792 =  n_5776 &  n_5791;
assign n_5793 =  n_3642 & ~n_5792;
assign n_5794 =  n_3656 & ~n_5793;
assign n_5795 = ~n_5762 &  n_5794;
assign n_5796 = ~n_5731 & ~n_5795;
assign n_5797 =  n_3263 &  n_3634;
assign n_5798 = ~n_3559 &  n_3616;
assign n_5799 = ~n_3571 & ~n_5798;
assign n_5800 = ~n_3573 & ~n_5799;
assign n_5801 =  n_3579 & ~n_5800;
assign n_5802 = ~n_3554 &  n_3574;
assign n_5803 = ~x_2436 & ~n_5802;
assign n_5804 =  n_5798 & ~n_5803;
assign n_5805 =  x_2436 &  n_3561;
assign n_5806 = ~n_3591 &  n_5805;
assign n_5807 = ~n_3586 &  n_5806;
assign n_5808 = ~n_3579 & ~n_5807;
assign n_5809 = ~n_5804 &  n_5808;
assign n_5810 = ~n_3626 & ~n_5809;
assign n_5811 = ~n_5801 &  n_5810;
assign n_5812 =  n_3598 &  n_3611;
assign n_5813 =  n_5811 &  n_5812;
assign n_5814 = ~n_4317 & ~n_4328;
assign n_5815 = ~n_4304 & ~n_4315;
assign n_5816 =  n_5814 &  n_5815;
assign n_5817 = ~i_1 & ~i_2;
assign n_5818 =  x_295 & ~n_5817;
assign n_5819 =  i_5 &  x_295;
assign n_5820 = ~i_6 &  n_5819;
assign n_5821 = ~n_4351 & ~n_5820;
assign n_5822 =  n_5818 &  n_5821;
assign n_5823 =  n_5822 & ~n_4355;
assign n_5824 =  i_3 &  x_295;
assign n_5825 = ~i_4 &  n_5824;
assign n_5826 = ~n_5825 &  n_4354;
assign n_5827 = ~n_5825 &  n_5821;
assign n_5828 = ~n_5826 & ~n_5827;
assign n_5829 = ~n_5823 &  n_5828;
assign n_5830 = ~n_1525 & ~n_5829;
assign n_5831 =  n_4349 & ~n_5829;
assign n_5832 = ~n_1522 & ~n_5831;
assign n_5833 =  x_2484 &  n_5832;
assign n_5834 =  x_2457 & ~n_5833;
assign n_5835 =  n_5830 & ~n_5834;
assign n_5836 = ~i_143 & ~x_2475;
assign n_5837 =  i_143 &  x_2475;
assign n_5838 = ~n_5836 & ~n_5837;
assign n_5839 =  i_145 & ~x_2474;
assign n_5840 = ~i_145 &  x_2474;
assign n_5841 = ~n_5839 & ~n_5840;
assign n_5842 = ~n_5838 &  n_5841;
assign n_5843 =  x_2476 & ~n_4323;
assign n_5844 = ~x_2476 &  n_4323;
assign n_5845 = ~n_5843 & ~n_5844;
assign n_5846 =  n_5842 &  n_5845;
assign n_5847 = ~x_2477 & ~n_4326;
assign n_5848 =  x_2477 &  n_4326;
assign n_5849 = ~n_5847 & ~n_5848;
assign n_5850 =  n_5816 & ~n_5849;
assign n_5851 =  n_5846 &  n_5850;
assign n_5852 =  x_2478 &  n_5851;
assign n_5853 = ~i_143 & ~x_2481;
assign n_5854 =  i_143 &  x_2481;
assign n_5855 = ~n_5853 & ~n_5854;
assign n_5856 =  i_145 & ~x_2480;
assign n_5857 = ~i_145 &  x_2480;
assign n_5858 = ~n_5856 & ~n_5857;
assign n_5859 = ~n_5855 &  n_5858;
assign n_5860 =  x_2482 & ~n_4326;
assign n_5861 = ~x_2482 &  n_4326;
assign n_5862 = ~n_5860 & ~n_5861;
assign n_5863 =  n_5859 &  n_5862;
assign n_5864 = ~x_2479 & ~n_4323;
assign n_5865 =  x_2479 &  n_4323;
assign n_5866 = ~n_5864 & ~n_5865;
assign n_5867 =  n_5816 & ~n_5866;
assign n_5868 =  n_5863 &  n_5867;
assign n_5869 =  x_2483 &  n_5868;
assign n_5870 = ~n_5852 & ~n_5869;
assign n_5871 = ~i_143 & ~x_2470;
assign n_5872 =  i_143 &  x_2470;
assign n_5873 = ~n_5871 & ~n_5872;
assign n_5874 =  i_145 & ~x_2469;
assign n_5875 = ~i_145 &  x_2469;
assign n_5876 = ~n_5874 & ~n_5875;
assign n_5877 = ~n_5873 &  n_5876;
assign n_5878 =  x_2471 & ~n_4323;
assign n_5879 = ~x_2471 &  n_4323;
assign n_5880 = ~n_5878 & ~n_5879;
assign n_5881 =  n_5877 &  n_5880;
assign n_5882 = ~x_2472 & ~n_4326;
assign n_5883 =  x_2472 &  n_4326;
assign n_5884 = ~n_5882 & ~n_5883;
assign n_5885 =  n_5816 & ~n_5884;
assign n_5886 =  n_5881 &  n_5885;
assign n_5887 =  x_2473 &  n_5886;
assign n_5888 = ~i_145 & ~x_2460;
assign n_5889 =  i_145 &  x_2460;
assign n_5890 = ~n_5888 & ~n_5889;
assign n_5891 =  i_143 & ~x_2459;
assign n_5892 = ~i_143 &  x_2459;
assign n_5893 = ~n_5891 & ~n_5892;
assign n_5894 = ~n_5890 &  n_5893;
assign n_5895 =  x_2461 & ~n_4326;
assign n_5896 = ~x_2461 &  n_4326;
assign n_5897 = ~n_5895 & ~n_5896;
assign n_5898 =  n_5894 &  n_5897;
assign n_5899 = ~x_2462 & ~n_4323;
assign n_5900 =  x_2462 &  n_4323;
assign n_5901 = ~n_5899 & ~n_5900;
assign n_5902 =  n_5816 & ~n_5901;
assign n_5903 =  n_5898 &  n_5902;
assign n_5904 =  x_2463 &  n_5903;
assign n_5905 = ~i_145 & ~x_2464;
assign n_5906 =  i_145 &  x_2464;
assign n_5907 = ~n_5905 & ~n_5906;
assign n_5908 =  i_143 & ~x_2466;
assign n_5909 = ~i_143 &  x_2466;
assign n_5910 = ~n_5908 & ~n_5909;
assign n_5911 = ~n_5907 &  n_5910;
assign n_5912 =  x_2465 & ~n_4323;
assign n_5913 = ~x_2465 &  n_4323;
assign n_5914 = ~n_5912 & ~n_5913;
assign n_5915 =  n_5911 &  n_5914;
assign n_5916 = ~x_2467 & ~n_4326;
assign n_5917 =  x_2467 &  n_4326;
assign n_5918 = ~n_5916 & ~n_5917;
assign n_5919 =  n_5816 & ~n_5918;
assign n_5920 =  n_5915 &  n_5919;
assign n_5921 =  x_2468 &  n_5920;
assign n_5922 = ~n_5904 & ~n_5921;
assign n_5923 = ~n_5887 &  n_5922;
assign n_5924 =  n_5870 &  n_5923;
assign n_5925 =  n_5835 &  n_5924;
assign n_5926 =  n_5816 &  n_5925;
assign n_5927 = ~x_2487 & ~x_2488;
assign n_5928 =  x_2486 & ~n_5927;
assign n_5929 =  n_5926 &  n_5928;
assign n_5930 = ~n_1525 &  n_4356;
assign n_5931 =  n_4349 &  n_4356;
assign n_5932 = ~n_1522 & ~n_5931;
assign n_5933 =  x_2485 &  n_5932;
assign n_5934 =  x_2458 & ~n_5933;
assign n_5935 =  n_5930 & ~n_5934;
assign n_5936 = ~n_5924 & ~n_5935;
assign n_5937 =  n_5835 &  n_5936;
assign n_5938 = ~i_2 & ~n_5821;
assign n_5939 =  n_4349 & ~n_5938;
assign n_5940 =  n_5823 & ~n_5939;
assign n_5941 =  n_4349 &  n_5818;
assign n_5942 =  n_5826 &  n_5941;
assign n_5943 =  x_2528 & ~n_5942;
assign n_5944 = ~n_5825 &  n_5822;
assign n_5945 =  n_5939 &  n_5944;
assign n_5946 =  x_2534 & ~n_5945;
assign n_5947 = ~n_5943 & ~n_5946;
assign n_5948 = ~n_5823 & ~n_5947;
assign n_5949 = ~n_4349 & ~n_4354;
assign n_5950 = ~n_5827 &  n_5949;
assign n_5951 = ~x_1731 & ~n_5950;
assign n_5952 = ~n_5948 &  n_5951;
assign n_5953 = ~n_5940 & ~n_5952;
assign n_5954 = ~x_1773 & ~n_4328;
assign n_5955 =  x_1773 &  n_4328;
assign n_5956 = ~n_5954 & ~n_5955;
assign n_5957 = ~x_1777 & ~n_4315;
assign n_5958 =  x_1777 &  n_4315;
assign n_5959 = ~n_5957 & ~n_5958;
assign n_5960 = ~i_143 &  x_1772;
assign n_5961 =  i_143 & ~x_1772;
assign n_5962 = ~n_5960 & ~n_5961;
assign n_5963 = ~i_145 &  x_1774;
assign n_5964 =  i_145 & ~x_1774;
assign n_5965 = ~n_5963 & ~n_5964;
assign n_5966 =  n_5962 &  n_5965;
assign n_5967 = ~n_5959 &  n_5966;
assign n_5968 = ~n_5956 &  n_5967;
assign n_5969 =  x_1776 & ~n_4323;
assign n_5970 = ~x_1775 &  n_4304;
assign n_5971 = ~n_5969 & ~n_5970;
assign n_5972 =  x_1775 & ~n_4304;
assign n_5973 = ~x_1776 &  n_4323;
assign n_5974 = ~n_5972 & ~n_5973;
assign n_5975 =  n_5971 &  n_5974;
assign n_5976 = ~x_1779 &  n_4317;
assign n_5977 =  x_1778 & ~n_4326;
assign n_5978 = ~n_5976 & ~n_5977;
assign n_5979 = ~x_1778 &  n_4326;
assign n_5980 =  x_1779 & ~n_4317;
assign n_5981 = ~n_5979 & ~n_5980;
assign n_5982 =  n_5978 &  n_5981;
assign n_5983 =  n_5975 &  n_5982;
assign n_5984 =  n_5968 &  n_5983;
assign n_5985 =  x_1467 &  n_1739;
assign n_5986 = ~n_5984 &  n_5985;
assign n_5987 = ~n_4349 &  n_5826;
assign n_5988 =  n_5818 &  n_5987;
assign n_5989 =  x_2529 &  n_5988;
assign n_5990 = ~n_5986 & ~n_5989;
assign n_5991 =  x_2435 &  n_3578;
assign n_5992 =  x_2452 & ~n_5991;
assign n_5993 =  x_1497 &  n_5992;
assign n_5994 =  x_1720 &  n_5992;
assign n_5995 = ~x_1496 &  n_5992;
assign n_5996 = ~n_5994 & ~n_5995;
assign n_5997 = ~x_1498 & ~x_2451;
assign n_5998 =  n_5996 &  n_5997;
assign n_5999 =  n_5993 & ~n_5998;
assign n_6000 = ~x_3157 &  n_5940;
assign n_6001 = ~n_5999 & ~n_6000;
assign n_6002 =  n_5990 &  n_6001;
assign n_6003 = ~i_7 & ~n_5824;
assign n_6004 =  n_4357 &  n_6003;
assign n_6005 =  n_4348 &  n_6004;
assign n_6006 =  n_6005 &  n_5822;
assign n_6007 =  x_2535 &  n_6006;
assign n_6008 =  n_4370 & ~n_5728;
assign n_6009 =  x_2544 &  n_6008;
assign n_6010 = ~x_2434 &  n_3570;
assign n_6011 =  x_2450 & ~x_3156;
assign n_6012 = ~n_6010 &  n_6011;
assign n_6013 = ~n_3571 & ~n_6012;
assign n_6014 = ~n_6009 & ~n_6013;
assign n_6015 = ~n_6007 &  n_6014;
assign n_6016 =  x_1754 & ~x_3156;
assign n_6017 = ~n_3555 &  n_6016;
assign n_6018 =  n_3570 &  n_6017;
assign n_6019 =  i_145 &  n_4323;
assign n_6020 = ~n_4326 & ~n_6019;
assign n_6021 =  n_5816 & ~n_6020;
assign n_6022 =  x_1729 & ~x_3073;
assign n_6023 =  x_3074 & ~x_3075;
assign n_6024 = ~n_6022 &  n_6023;
assign n_6025 = ~x_3236 & ~n_6024;
assign n_6026 =  n_1328 & ~n_6025;
assign n_6027 = ~n_6021 & ~n_6026;
assign n_6028 = ~n_6018 &  n_6027;
assign n_6029 =  x_1726 & ~x_3070;
assign n_6030 =  x_3071 & ~n_6029;
assign n_6031 = ~n_3676 & ~n_3679;
assign n_6032 = ~x_3072 &  n_6031;
assign n_6033 =  n_6030 &  n_6032;
assign n_6034 = ~x_3069 &  n_3685;
assign n_6035 =  n_6034 &  n_6030;
assign n_6036 = ~n_6033 & ~n_6035;
assign n_6037 =  x_226 &  n_1739;
assign n_6038 =  x_2524 & ~x_2526;
assign n_6039 = ~x_2527 &  n_6038;
assign n_6040 =  n_6037 & ~n_6039;
assign n_6041 = ~x_2434 &  x_3234;
assign n_6042 = ~x_2454 & ~x_2455;
assign n_6043 =  x_2456 & ~n_6042;
assign n_6044 = ~n_6041 & ~n_6043;
assign n_6045 =  n_3563 & ~n_6044;
assign n_6046 = ~n_6040 & ~n_6045;
assign n_6047 =  n_6036 &  n_6046;
assign n_6048 =  n_6028 &  n_6047;
assign n_6049 = ~x_2540 &  n_1739;
assign n_6050 = ~i_14 & ~i_222;
assign n_6051 =  x_295 & ~n_6050;
assign n_6052 =  i_221 &  x_295;
assign n_6053 =  n_6050 &  n_6052;
assign n_6054 = ~x_2541 &  n_6053;
assign n_6055 = ~n_6051 & ~n_6054;
assign n_6056 =  n_6049 &  n_6055;
assign n_6057 =  x_2542 &  n_6056;
assign n_6058 =  x_1498 &  n_5992;
assign n_6059 =  x_2451 &  n_6058;
assign n_6060 = ~n_5996 &  n_6059;
assign n_6061 = ~n_6057 & ~n_6060;
assign n_6062 =  n_6048 &  n_6061;
assign n_6063 = ~x_227 &  n_3673;
assign n_6064 = ~n_6022 &  n_6063;
assign n_6065 =  x_3074 &  n_6064;
assign n_6066 = ~x_2433 & ~n_3563;
assign n_6067 = ~i_218 &  n_3565;
assign n_6068 = ~x_1754 & ~n_3569;
assign n_6069 =  n_6067 & ~n_6068;
assign n_6070 = ~n_6066 &  n_6069;
assign n_6071 =  x_3155 &  n_3591;
assign n_6072 = ~n_6070 &  n_6071;
assign n_6073 = ~n_1325 &  n_6022;
assign n_6074 = ~n_6063 &  n_6073;
assign n_6075 = ~x_3074 &  n_6074;
assign n_6076 = ~n_6072 & ~n_6075;
assign n_6077 = ~n_6065 &  n_6076;
assign n_6078 =  x_2542 & ~x_2543;
assign n_6079 =  n_1525 &  n_6078;
assign n_6080 =  n_6055 &  n_6079;
assign n_6081 =  x_3239 &  n_3673;
assign n_6082 = ~x_3238 & ~n_6081;
assign n_6083 =  x_3237 &  n_6067;
assign n_6084 =  x_3235 &  n_1739;
assign n_6085 = ~n_6083 & ~n_6084;
assign n_6086 =  n_6082 &  n_6085;
assign n_6087 = ~n_6080 &  n_6086;
assign n_6088 = ~n_6049 &  n_6054;
assign n_6089 = ~x_2542 &  n_6088;
assign n_6090 = ~n_3676 &  n_6029;
assign n_6091 = ~n_6034 &  n_6090;
assign n_6092 = ~x_3071 &  n_6091;
assign n_6093 = ~n_6089 & ~n_6092;
assign n_6094 =  n_6087 &  n_6093;
assign n_6095 =  n_6077 &  n_6094;
assign n_6096 =  n_6062 &  n_6095;
assign n_6097 =  n_6015 &  n_6096;
assign n_6098 =  n_6002 &  n_6097;
assign n_6099 = ~n_5953 &  n_6098;
assign n_6100 = ~n_5937 &  n_6099;
assign n_6101 = ~n_5929 &  n_6100;
assign n_6102 = ~n_5813 &  n_6101;
assign n_6103 = ~n_5797 &  n_6102;
assign n_6104 = ~n_5796 &  n_6103;
assign n_6105 = ~n_5730 &  n_6104;
assign n_6106 =  x_3230 & ~n_6105;
assign n_6107 = ~x_3230 &  n_6105;
assign n_6108 = ~n_6106 & ~n_6107;
assign n_6109 =  x_1562 &  x_1736;
assign n_6110 = ~x_451 & ~n_6109;
assign n_6111 =  x_1732 & ~n_6110;
assign n_6112 = ~x_1562 & ~x_1736;
assign n_6113 =  i_80 &  x_295;
assign n_6114 =  i_79 & ~x_1732;
assign n_6115 = ~n_6113 &  n_6114;
assign n_6116 = ~n_4350 & ~n_5819;
assign n_6117 =  n_6115 &  n_6116;
assign n_6118 = ~n_4349 &  n_6117;
assign n_6119 = ~i_3 &  n_1739;
assign n_6120 =  n_6118 &  n_6119;
assign n_6121 = ~x_1733 & ~n_6120;
assign n_6122 = ~i_1 &  n_1739;
assign n_6123 =  n_6122 &  n_5824;
assign n_6124 =  n_6118 &  n_6123;
assign n_6125 = ~x_1735 & ~n_6124;
assign n_6126 =  i_79 &  n_1739;
assign n_6127 = ~n_6113 &  n_6126;
assign n_6128 =  n_6127 &  n_5988;
assign n_6129 = ~x_1732 & ~n_6128;
assign n_6130 =  n_6125 & ~n_6129;
assign n_6131 = ~n_4357 &  n_5987;
assign n_6132 = ~n_6006 & ~n_6131;
assign n_6133 =  n_6127 & ~n_6132;
assign n_6134 = ~x_1732 & ~n_6133;
assign n_6135 =  n_6130 & ~n_6134;
assign n_6136 = ~n_6121 &  n_6135;
assign n_6137 = ~n_6112 &  n_6136;
assign n_6138 = ~n_6111 & ~n_6137;
assign n_6139 =  x_3229 &  n_6138;
assign n_6140 = ~x_3229 & ~n_6138;
assign n_6141 = ~n_6139 & ~n_6140;
assign n_6142 =  n_1321 &  n_4291;
assign n_6143 = ~n_1220 & ~n_6142;
assign n_6144 =  x_230 &  x_1470;
assign n_6145 =  n_1714 & ~n_6144;
assign n_6146 = ~n_6143 & ~n_6145;
assign n_6147 = ~x_230 & ~x_1139;
assign n_6148 = ~x_1139 &  n_1126;
assign n_6149 = ~x_2358 &  n_447;
assign n_6150 = ~x_2360 &  n_449;
assign n_6151 = ~n_6149 & ~n_6150;
assign n_6152 = ~x_2364 &  n_441;
assign n_6153 = ~x_2362 &  n_444;
assign n_6154 = ~n_6152 & ~n_6153;
assign n_6155 =  n_6151 &  n_6154;
assign n_6156 = ~x_2365 &  n_460;
assign n_6157 = ~x_2363 &  n_468;
assign n_6158 = ~n_6156 & ~n_6157;
assign n_6159 = ~x_2359 &  n_463;
assign n_6160 = ~x_2361 &  n_466;
assign n_6161 = ~n_6159 & ~n_6160;
assign n_6162 =  n_6158 &  n_6161;
assign n_6163 =  n_6155 &  n_6162;
assign n_6164 =  x_231 &  n_6163;
assign n_6165 = ~n_6148 & ~n_6164;
assign n_6166 = ~x_1470 & ~n_6165;
assign n_6167 = ~n_6147 & ~n_6166;
assign n_6168 =  n_1713 & ~n_6167;
assign n_6169 =  x_1201 & ~n_436;
assign n_6170 =  n_436 &  n_6163;
assign n_6171 = ~n_6169 & ~n_6170;
assign n_6172 =  n_1321 & ~n_6171;
assign n_6173 = ~n_6168 & ~n_6172;
assign n_6174 = ~n_6146 & ~n_6173;
assign n_6175 =  x_3228 &  n_6146;
assign n_6176 = ~n_6174 & ~n_6175;
assign n_6177 =  x_3228 & ~n_6176;
assign n_6178 = ~x_3228 &  n_6176;
assign n_6179 = ~n_6177 & ~n_6178;
assign n_6180 = ~x_230 & ~x_1138;
assign n_6181 = ~x_1138 &  n_1126;
assign n_6182 = ~x_2356 &  n_441;
assign n_6183 = ~x_2354 &  n_444;
assign n_6184 = ~n_6182 & ~n_6183;
assign n_6185 = ~x_2352 &  n_449;
assign n_6186 = ~x_2350 &  n_447;
assign n_6187 = ~n_6185 & ~n_6186;
assign n_6188 =  n_6184 &  n_6187;
assign n_6189 = ~x_2357 &  n_460;
assign n_6190 = ~x_2353 &  n_466;
assign n_6191 = ~n_6189 & ~n_6190;
assign n_6192 = ~x_2351 &  n_463;
assign n_6193 = ~x_2355 &  n_468;
assign n_6194 = ~n_6192 & ~n_6193;
assign n_6195 =  n_6191 &  n_6194;
assign n_6196 =  n_6188 &  n_6195;
assign n_6197 =  x_231 &  n_6196;
assign n_6198 = ~n_6181 & ~n_6197;
assign n_6199 = ~x_1470 & ~n_6198;
assign n_6200 = ~n_6180 & ~n_6199;
assign n_6201 =  n_1713 & ~n_6200;
assign n_6202 =  x_1200 & ~n_436;
assign n_6203 =  n_436 &  n_6196;
assign n_6204 = ~n_6202 & ~n_6203;
assign n_6205 =  n_1321 & ~n_6204;
assign n_6206 = ~n_6201 & ~n_6205;
assign n_6207 = ~n_6146 & ~n_6206;
assign n_6208 =  x_3227 &  n_6146;
assign n_6209 = ~n_6207 & ~n_6208;
assign n_6210 =  x_3227 & ~n_6209;
assign n_6211 = ~x_3227 &  n_6209;
assign n_6212 = ~n_6210 & ~n_6211;
assign n_6213 = ~x_230 & ~x_1137;
assign n_6214 = ~x_1137 &  n_1126;
assign n_6215 = ~x_2344 &  n_449;
assign n_6216 = ~x_2342 &  n_447;
assign n_6217 = ~n_6215 & ~n_6216;
assign n_6218 = ~x_2348 &  n_441;
assign n_6219 = ~x_2346 &  n_444;
assign n_6220 = ~n_6218 & ~n_6219;
assign n_6221 =  n_6217 &  n_6220;
assign n_6222 = ~x_2345 &  n_466;
assign n_6223 = ~x_2347 &  n_468;
assign n_6224 = ~n_6222 & ~n_6223;
assign n_6225 = ~x_2343 &  n_463;
assign n_6226 = ~x_2349 &  n_460;
assign n_6227 = ~n_6225 & ~n_6226;
assign n_6228 =  n_6224 &  n_6227;
assign n_6229 =  n_6221 &  n_6228;
assign n_6230 =  x_231 &  n_6229;
assign n_6231 = ~n_6214 & ~n_6230;
assign n_6232 = ~x_1470 & ~n_6231;
assign n_6233 = ~n_6213 & ~n_6232;
assign n_6234 =  n_1713 & ~n_6233;
assign n_6235 =  x_1199 & ~n_436;
assign n_6236 =  n_436 &  n_6229;
assign n_6237 = ~n_6235 & ~n_6236;
assign n_6238 =  n_1321 & ~n_6237;
assign n_6239 = ~n_6234 & ~n_6238;
assign n_6240 = ~n_6146 & ~n_6239;
assign n_6241 =  x_3226 &  n_6146;
assign n_6242 = ~n_6240 & ~n_6241;
assign n_6243 =  x_3226 & ~n_6242;
assign n_6244 = ~x_3226 &  n_6242;
assign n_6245 = ~n_6243 & ~n_6244;
assign n_6246 = ~x_230 & ~x_1136;
assign n_6247 = ~x_1136 &  n_1126;
assign n_6248 = ~x_2334 &  n_447;
assign n_6249 = ~x_2336 &  n_449;
assign n_6250 = ~n_6248 & ~n_6249;
assign n_6251 = ~x_2338 &  n_444;
assign n_6252 = ~x_2340 &  n_441;
assign n_6253 = ~n_6251 & ~n_6252;
assign n_6254 =  n_6250 &  n_6253;
assign n_6255 = ~x_2339 &  n_468;
assign n_6256 = ~x_2341 &  n_460;
assign n_6257 = ~n_6255 & ~n_6256;
assign n_6258 = ~x_2335 &  n_463;
assign n_6259 = ~x_2337 &  n_466;
assign n_6260 = ~n_6258 & ~n_6259;
assign n_6261 =  n_6257 &  n_6260;
assign n_6262 =  n_6254 &  n_6261;
assign n_6263 =  x_231 &  n_6262;
assign n_6264 = ~n_6247 & ~n_6263;
assign n_6265 = ~x_1470 & ~n_6264;
assign n_6266 = ~n_6246 & ~n_6265;
assign n_6267 =  n_1713 & ~n_6266;
assign n_6268 =  x_1198 & ~n_436;
assign n_6269 =  n_436 &  n_6262;
assign n_6270 = ~n_6268 & ~n_6269;
assign n_6271 =  n_1321 & ~n_6270;
assign n_6272 = ~n_6267 & ~n_6271;
assign n_6273 = ~n_6146 & ~n_6272;
assign n_6274 =  x_3225 &  n_6146;
assign n_6275 = ~n_6273 & ~n_6274;
assign n_6276 =  x_3225 & ~n_6275;
assign n_6277 = ~x_3225 &  n_6275;
assign n_6278 = ~n_6276 & ~n_6277;
assign n_6279 = ~x_230 & ~x_1135;
assign n_6280 = ~x_1135 &  n_1126;
assign n_6281 = ~x_2328 &  n_449;
assign n_6282 = ~x_2330 &  n_444;
assign n_6283 = ~n_6281 & ~n_6282;
assign n_6284 = ~x_2332 &  n_441;
assign n_6285 = ~x_2326 &  n_447;
assign n_6286 = ~n_6284 & ~n_6285;
assign n_6287 =  n_6283 &  n_6286;
assign n_6288 = ~x_2331 &  n_468;
assign n_6289 = ~x_2329 &  n_466;
assign n_6290 = ~n_6288 & ~n_6289;
assign n_6291 = ~x_2327 &  n_463;
assign n_6292 = ~x_2333 &  n_460;
assign n_6293 = ~n_6291 & ~n_6292;
assign n_6294 =  n_6290 &  n_6293;
assign n_6295 =  n_6287 &  n_6294;
assign n_6296 =  x_231 &  n_6295;
assign n_6297 = ~n_6280 & ~n_6296;
assign n_6298 = ~x_1470 & ~n_6297;
assign n_6299 = ~n_6279 & ~n_6298;
assign n_6300 =  n_1713 & ~n_6299;
assign n_6301 =  x_1197 & ~n_436;
assign n_6302 =  n_436 &  n_6295;
assign n_6303 = ~n_6301 & ~n_6302;
assign n_6304 =  n_1321 & ~n_6303;
assign n_6305 = ~n_6300 & ~n_6304;
assign n_6306 = ~n_6146 & ~n_6305;
assign n_6307 =  x_3224 &  n_6146;
assign n_6308 = ~n_6306 & ~n_6307;
assign n_6309 =  x_3224 & ~n_6308;
assign n_6310 = ~x_3224 &  n_6308;
assign n_6311 = ~n_6309 & ~n_6310;
assign n_6312 = ~x_230 & ~x_1134;
assign n_6313 = ~x_1134 &  n_1126;
assign n_6314 = ~x_2318 &  n_447;
assign n_6315 = ~x_2320 &  n_449;
assign n_6316 = ~n_6314 & ~n_6315;
assign n_6317 = ~x_2324 &  n_441;
assign n_6318 = ~x_2322 &  n_444;
assign n_6319 = ~n_6317 & ~n_6318;
assign n_6320 =  n_6316 &  n_6319;
assign n_6321 = ~x_2321 &  n_466;
assign n_6322 = ~x_2323 &  n_468;
assign n_6323 = ~n_6321 & ~n_6322;
assign n_6324 = ~x_2325 &  n_460;
assign n_6325 = ~x_2319 &  n_463;
assign n_6326 = ~n_6324 & ~n_6325;
assign n_6327 =  n_6323 &  n_6326;
assign n_6328 =  n_6320 &  n_6327;
assign n_6329 =  x_231 &  n_6328;
assign n_6330 = ~n_6313 & ~n_6329;
assign n_6331 = ~x_1470 & ~n_6330;
assign n_6332 = ~n_6312 & ~n_6331;
assign n_6333 =  n_1713 & ~n_6332;
assign n_6334 =  x_1196 & ~n_436;
assign n_6335 =  n_436 &  n_6328;
assign n_6336 = ~n_6334 & ~n_6335;
assign n_6337 =  n_1321 & ~n_6336;
assign n_6338 = ~n_6333 & ~n_6337;
assign n_6339 = ~n_6146 & ~n_6338;
assign n_6340 =  x_3223 &  n_6146;
assign n_6341 = ~n_6339 & ~n_6340;
assign n_6342 =  x_3223 & ~n_6341;
assign n_6343 = ~x_3223 &  n_6341;
assign n_6344 = ~n_6342 & ~n_6343;
assign n_6345 = ~x_230 & ~x_1133;
assign n_6346 = ~x_1133 &  n_1126;
assign n_6347 = ~x_2310 &  n_447;
assign n_6348 = ~x_2312 &  n_449;
assign n_6349 = ~n_6347 & ~n_6348;
assign n_6350 = ~x_2316 &  n_441;
assign n_6351 = ~x_2314 &  n_444;
assign n_6352 = ~n_6350 & ~n_6351;
assign n_6353 =  n_6349 &  n_6352;
assign n_6354 = ~x_2317 &  n_460;
assign n_6355 = ~x_2315 &  n_468;
assign n_6356 = ~n_6354 & ~n_6355;
assign n_6357 = ~x_2311 &  n_463;
assign n_6358 = ~x_2313 &  n_466;
assign n_6359 = ~n_6357 & ~n_6358;
assign n_6360 =  n_6356 &  n_6359;
assign n_6361 =  n_6353 &  n_6360;
assign n_6362 =  x_231 &  n_6361;
assign n_6363 = ~n_6346 & ~n_6362;
assign n_6364 = ~x_1470 & ~n_6363;
assign n_6365 = ~n_6345 & ~n_6364;
assign n_6366 =  n_1713 & ~n_6365;
assign n_6367 =  x_1195 & ~n_436;
assign n_6368 =  n_436 &  n_6361;
assign n_6369 = ~n_6367 & ~n_6368;
assign n_6370 =  n_1321 & ~n_6369;
assign n_6371 = ~n_6366 & ~n_6370;
assign n_6372 = ~n_6146 & ~n_6371;
assign n_6373 =  x_3222 &  n_6146;
assign n_6374 = ~n_6372 & ~n_6373;
assign n_6375 =  x_3222 & ~n_6374;
assign n_6376 = ~x_3222 &  n_6374;
assign n_6377 = ~n_6375 & ~n_6376;
assign n_6378 = ~x_230 & ~x_1132;
assign n_6379 = ~x_1132 &  n_1126;
assign n_6380 = ~x_2304 &  n_449;
assign n_6381 = ~x_2306 &  n_444;
assign n_6382 = ~n_6380 & ~n_6381;
assign n_6383 = ~x_2308 &  n_441;
assign n_6384 = ~x_2302 &  n_447;
assign n_6385 = ~n_6383 & ~n_6384;
assign n_6386 =  n_6382 &  n_6385;
assign n_6387 = ~x_2307 &  n_468;
assign n_6388 = ~x_2305 &  n_466;
assign n_6389 = ~n_6387 & ~n_6388;
assign n_6390 = ~x_2303 &  n_463;
assign n_6391 = ~x_2309 &  n_460;
assign n_6392 = ~n_6390 & ~n_6391;
assign n_6393 =  n_6389 &  n_6392;
assign n_6394 =  n_6386 &  n_6393;
assign n_6395 =  x_231 &  n_6394;
assign n_6396 = ~n_6379 & ~n_6395;
assign n_6397 = ~x_1470 & ~n_6396;
assign n_6398 = ~n_6378 & ~n_6397;
assign n_6399 =  n_1713 & ~n_6398;
assign n_6400 =  x_1194 & ~n_436;
assign n_6401 =  n_436 &  n_6394;
assign n_6402 = ~n_6400 & ~n_6401;
assign n_6403 =  n_1321 & ~n_6402;
assign n_6404 = ~n_6399 & ~n_6403;
assign n_6405 =  x_3221 &  n_6404;
assign n_6406 = ~x_3221 & ~n_6404;
assign n_6407 = ~n_6405 & ~n_6406;
assign n_6408 =  n_6146 & ~n_4181;
assign n_6409 =  x_3220 & ~n_6408;
assign n_6410 = ~x_3220 &  n_6408;
assign n_6411 = ~n_6409 & ~n_6410;
assign n_6412 = ~x_230 & ~x_1131;
assign n_6413 = ~x_1131 &  n_1126;
assign n_6414 = ~x_2294 &  n_447;
assign n_6415 = ~x_2296 &  n_449;
assign n_6416 = ~n_6414 & ~n_6415;
assign n_6417 = ~x_2298 &  n_444;
assign n_6418 = ~x_2300 &  n_441;
assign n_6419 = ~n_6417 & ~n_6418;
assign n_6420 =  n_6416 &  n_6419;
assign n_6421 = ~x_2299 &  n_468;
assign n_6422 = ~x_2295 &  n_463;
assign n_6423 = ~n_6421 & ~n_6422;
assign n_6424 = ~x_2301 &  n_460;
assign n_6425 = ~x_2297 &  n_466;
assign n_6426 = ~n_6424 & ~n_6425;
assign n_6427 =  n_6423 &  n_6426;
assign n_6428 =  n_6420 &  n_6427;
assign n_6429 =  x_231 &  n_6428;
assign n_6430 = ~n_6413 & ~n_6429;
assign n_6431 = ~x_1470 & ~n_6430;
assign n_6432 = ~n_6412 & ~n_6431;
assign n_6433 =  n_1713 & ~n_6432;
assign n_6434 =  x_1193 & ~n_436;
assign n_6435 =  n_436 &  n_6428;
assign n_6436 = ~n_6434 & ~n_6435;
assign n_6437 =  n_1321 & ~n_6436;
assign n_6438 = ~n_6433 & ~n_6437;
assign n_6439 = ~n_6146 & ~n_6438;
assign n_6440 =  x_3219 &  n_6146;
assign n_6441 = ~n_6439 & ~n_6440;
assign n_6442 =  x_3219 & ~n_6441;
assign n_6443 = ~x_3219 &  n_6441;
assign n_6444 = ~n_6442 & ~n_6443;
assign n_6445 = ~x_230 & ~x_1130;
assign n_6446 = ~x_1130 &  n_1126;
assign n_6447 = ~x_2292 &  n_441;
assign n_6448 = ~x_2286 &  n_447;
assign n_6449 = ~n_6447 & ~n_6448;
assign n_6450 = ~x_2288 &  n_449;
assign n_6451 = ~x_2290 &  n_444;
assign n_6452 = ~n_6450 & ~n_6451;
assign n_6453 =  n_6449 &  n_6452;
assign n_6454 = ~x_2291 &  n_468;
assign n_6455 = ~x_2293 &  n_460;
assign n_6456 = ~n_6454 & ~n_6455;
assign n_6457 = ~x_2287 &  n_463;
assign n_6458 = ~x_2289 &  n_466;
assign n_6459 = ~n_6457 & ~n_6458;
assign n_6460 =  n_6456 &  n_6459;
assign n_6461 =  n_6453 &  n_6460;
assign n_6462 =  x_231 &  n_6461;
assign n_6463 = ~n_6446 & ~n_6462;
assign n_6464 = ~x_1470 & ~n_6463;
assign n_6465 = ~n_6445 & ~n_6464;
assign n_6466 =  n_1713 & ~n_6465;
assign n_6467 =  x_1192 & ~n_436;
assign n_6468 =  n_436 &  n_6461;
assign n_6469 = ~n_6467 & ~n_6468;
assign n_6470 =  n_1321 & ~n_6469;
assign n_6471 = ~n_6466 & ~n_6470;
assign n_6472 = ~n_6146 & ~n_6471;
assign n_6473 =  x_3218 &  n_6146;
assign n_6474 = ~n_6472 & ~n_6473;
assign n_6475 =  x_3218 & ~n_6474;
assign n_6476 = ~x_3218 &  n_6474;
assign n_6477 = ~n_6475 & ~n_6476;
assign n_6478 = ~x_230 & ~x_1129;
assign n_6479 = ~x_1129 &  n_1126;
assign n_6480 = ~x_2278 &  n_447;
assign n_6481 = ~x_2284 &  n_441;
assign n_6482 = ~n_6480 & ~n_6481;
assign n_6483 = ~x_2282 &  n_444;
assign n_6484 = ~x_2280 &  n_449;
assign n_6485 = ~n_6483 & ~n_6484;
assign n_6486 =  n_6482 &  n_6485;
assign n_6487 = ~x_2283 &  n_468;
assign n_6488 = ~x_2281 &  n_466;
assign n_6489 = ~n_6487 & ~n_6488;
assign n_6490 = ~x_2285 &  n_460;
assign n_6491 = ~x_2279 &  n_463;
assign n_6492 = ~n_6490 & ~n_6491;
assign n_6493 =  n_6489 &  n_6492;
assign n_6494 =  n_6486 &  n_6493;
assign n_6495 =  x_231 &  n_6494;
assign n_6496 = ~n_6479 & ~n_6495;
assign n_6497 = ~x_1470 & ~n_6496;
assign n_6498 = ~n_6478 & ~n_6497;
assign n_6499 =  n_1713 & ~n_6498;
assign n_6500 =  x_1191 & ~n_436;
assign n_6501 =  n_436 &  n_6494;
assign n_6502 = ~n_6500 & ~n_6501;
assign n_6503 =  n_1321 & ~n_6502;
assign n_6504 = ~n_6499 & ~n_6503;
assign n_6505 = ~n_6146 & ~n_6504;
assign n_6506 =  x_3217 &  n_6146;
assign n_6507 = ~n_6505 & ~n_6506;
assign n_6508 =  x_3217 & ~n_6507;
assign n_6509 = ~x_3217 &  n_6507;
assign n_6510 = ~n_6508 & ~n_6509;
assign n_6511 = ~x_230 & ~x_1128;
assign n_6512 = ~x_1128 &  n_1126;
assign n_6513 = ~x_2276 &  n_441;
assign n_6514 = ~x_2270 &  n_447;
assign n_6515 = ~n_6513 & ~n_6514;
assign n_6516 = ~x_2272 &  n_449;
assign n_6517 = ~x_2274 &  n_444;
assign n_6518 = ~n_6516 & ~n_6517;
assign n_6519 =  n_6515 &  n_6518;
assign n_6520 = ~x_2275 &  n_468;
assign n_6521 = ~x_2273 &  n_466;
assign n_6522 = ~n_6520 & ~n_6521;
assign n_6523 = ~x_2271 &  n_463;
assign n_6524 = ~x_2277 &  n_460;
assign n_6525 = ~n_6523 & ~n_6524;
assign n_6526 =  n_6522 &  n_6525;
assign n_6527 =  n_6519 &  n_6526;
assign n_6528 =  x_231 &  n_6527;
assign n_6529 = ~n_6512 & ~n_6528;
assign n_6530 = ~x_1470 & ~n_6529;
assign n_6531 = ~n_6511 & ~n_6530;
assign n_6532 =  n_1713 & ~n_6531;
assign n_6533 =  x_1190 & ~n_436;
assign n_6534 =  n_436 &  n_6527;
assign n_6535 = ~n_6533 & ~n_6534;
assign n_6536 =  n_1321 & ~n_6535;
assign n_6537 = ~n_6532 & ~n_6536;
assign n_6538 = ~n_6146 & ~n_6537;
assign n_6539 =  x_3216 &  n_6146;
assign n_6540 = ~n_6538 & ~n_6539;
assign n_6541 =  x_3216 & ~n_6540;
assign n_6542 = ~x_3216 &  n_6540;
assign n_6543 = ~n_6541 & ~n_6542;
assign n_6544 = ~x_230 & ~x_1127;
assign n_6545 = ~x_1127 &  n_1126;
assign n_6546 = ~x_2262 &  n_447;
assign n_6547 = ~x_2268 &  n_441;
assign n_6548 = ~n_6546 & ~n_6547;
assign n_6549 = ~x_2266 &  n_444;
assign n_6550 = ~x_2264 &  n_449;
assign n_6551 = ~n_6549 & ~n_6550;
assign n_6552 =  n_6548 &  n_6551;
assign n_6553 = ~x_2269 &  n_460;
assign n_6554 = ~x_2265 &  n_466;
assign n_6555 = ~n_6553 & ~n_6554;
assign n_6556 = ~x_2267 &  n_468;
assign n_6557 = ~x_2263 &  n_463;
assign n_6558 = ~n_6556 & ~n_6557;
assign n_6559 =  n_6555 &  n_6558;
assign n_6560 =  n_6552 &  n_6559;
assign n_6561 =  x_231 &  n_6560;
assign n_6562 = ~n_6545 & ~n_6561;
assign n_6563 = ~x_1470 & ~n_6562;
assign n_6564 = ~n_6544 & ~n_6563;
assign n_6565 =  n_1713 & ~n_6564;
assign n_6566 =  x_1189 & ~n_436;
assign n_6567 =  n_436 &  n_6560;
assign n_6568 = ~n_6566 & ~n_6567;
assign n_6569 =  n_1321 & ~n_6568;
assign n_6570 = ~n_6565 & ~n_6569;
assign n_6571 = ~n_6146 & ~n_6570;
assign n_6572 =  x_3215 &  n_6146;
assign n_6573 = ~n_6571 & ~n_6572;
assign n_6574 =  x_3215 & ~n_6573;
assign n_6575 = ~x_3215 &  n_6573;
assign n_6576 = ~n_6574 & ~n_6575;
assign n_6577 = ~x_230 & ~x_1126;
assign n_6578 = ~x_1126 &  n_1126;
assign n_6579 = ~x_2254 &  n_447;
assign n_6580 = ~x_2260 &  n_441;
assign n_6581 = ~n_6579 & ~n_6580;
assign n_6582 = ~x_2258 &  n_444;
assign n_6583 = ~x_2256 &  n_449;
assign n_6584 = ~n_6582 & ~n_6583;
assign n_6585 =  n_6581 &  n_6584;
assign n_6586 = ~x_2255 &  n_463;
assign n_6587 = ~x_2257 &  n_466;
assign n_6588 = ~n_6586 & ~n_6587;
assign n_6589 = ~x_2259 &  n_468;
assign n_6590 = ~x_2261 &  n_460;
assign n_6591 = ~n_6589 & ~n_6590;
assign n_6592 =  n_6588 &  n_6591;
assign n_6593 =  n_6585 &  n_6592;
assign n_6594 =  x_231 &  n_6593;
assign n_6595 = ~n_6578 & ~n_6594;
assign n_6596 = ~x_1470 & ~n_6595;
assign n_6597 = ~n_6577 & ~n_6596;
assign n_6598 =  n_1713 & ~n_6597;
assign n_6599 =  x_1188 & ~n_436;
assign n_6600 =  n_436 &  n_6593;
assign n_6601 = ~n_6599 & ~n_6600;
assign n_6602 =  n_1321 & ~n_6601;
assign n_6603 = ~n_6598 & ~n_6602;
assign n_6604 = ~n_6146 & ~n_6603;
assign n_6605 =  x_3214 &  n_6146;
assign n_6606 = ~n_6604 & ~n_6605;
assign n_6607 =  x_3214 & ~n_6606;
assign n_6608 = ~x_3214 &  n_6606;
assign n_6609 = ~n_6607 & ~n_6608;
assign n_6610 = ~x_230 & ~x_1125;
assign n_6611 = ~x_1125 &  n_1126;
assign n_6612 = ~x_2246 &  n_447;
assign n_6613 = ~x_2252 &  n_441;
assign n_6614 = ~n_6612 & ~n_6613;
assign n_6615 = ~x_2248 &  n_449;
assign n_6616 = ~x_2250 &  n_444;
assign n_6617 = ~n_6615 & ~n_6616;
assign n_6618 =  n_6614 &  n_6617;
assign n_6619 = ~x_2249 &  n_466;
assign n_6620 = ~x_2253 &  n_460;
assign n_6621 = ~n_6619 & ~n_6620;
assign n_6622 = ~x_2251 &  n_468;
assign n_6623 = ~x_2247 &  n_463;
assign n_6624 = ~n_6622 & ~n_6623;
assign n_6625 =  n_6621 &  n_6624;
assign n_6626 =  n_6618 &  n_6625;
assign n_6627 =  x_231 &  n_6626;
assign n_6628 = ~n_6611 & ~n_6627;
assign n_6629 = ~x_1470 & ~n_6628;
assign n_6630 = ~n_6610 & ~n_6629;
assign n_6631 =  n_1713 & ~n_6630;
assign n_6632 =  x_1187 & ~n_436;
assign n_6633 =  n_436 &  n_6626;
assign n_6634 = ~n_6632 & ~n_6633;
assign n_6635 =  n_1321 & ~n_6634;
assign n_6636 = ~n_6631 & ~n_6635;
assign n_6637 = ~n_6146 & ~n_6636;
assign n_6638 =  x_3213 &  n_6146;
assign n_6639 = ~n_6637 & ~n_6638;
assign n_6640 =  x_3213 & ~n_6639;
assign n_6641 = ~x_3213 &  n_6639;
assign n_6642 = ~n_6640 & ~n_6641;
assign n_6643 =  x_1186 & ~n_436;
assign n_6644 = ~x_2238 &  n_447;
assign n_6645 = ~x_2242 &  n_444;
assign n_6646 = ~n_6644 & ~n_6645;
assign n_6647 = ~x_2240 &  n_449;
assign n_6648 = ~x_2244 &  n_441;
assign n_6649 = ~n_6647 & ~n_6648;
assign n_6650 =  n_6646 &  n_6649;
assign n_6651 = ~x_2239 &  n_463;
assign n_6652 = ~x_2241 &  n_466;
assign n_6653 = ~n_6651 & ~n_6652;
assign n_6654 = ~x_2243 &  n_468;
assign n_6655 = ~x_2245 &  n_460;
assign n_6656 = ~n_6654 & ~n_6655;
assign n_6657 =  n_6653 &  n_6656;
assign n_6658 =  n_6650 &  n_6657;
assign n_6659 =  n_436 &  n_6658;
assign n_6660 = ~n_6643 & ~n_6659;
assign n_6661 =  n_1321 & ~n_6660;
assign n_6662 = ~x_230 & ~x_1124;
assign n_6663 = ~x_1124 &  n_1126;
assign n_6664 =  x_231 &  n_6658;
assign n_6665 = ~n_6663 & ~n_6664;
assign n_6666 = ~x_1470 & ~n_6665;
assign n_6667 = ~n_6662 & ~n_6666;
assign n_6668 =  n_1713 & ~n_6667;
assign n_6669 = ~n_6661 & ~n_6668;
assign n_6670 =  x_3212 &  n_6669;
assign n_6671 = ~x_3212 & ~n_6669;
assign n_6672 = ~n_6670 & ~n_6671;
assign n_6673 =  n_6146 & ~n_4072;
assign n_6674 =  x_3211 & ~n_6673;
assign n_6675 = ~x_3211 &  n_6673;
assign n_6676 = ~n_6674 & ~n_6675;
assign n_6677 = ~x_230 & ~x_1123;
assign n_6678 = ~x_1123 &  n_1126;
assign n_6679 = ~x_2236 &  n_441;
assign n_6680 = ~x_2232 &  n_449;
assign n_6681 = ~n_6679 & ~n_6680;
assign n_6682 = ~x_2234 &  n_444;
assign n_6683 = ~x_2230 &  n_447;
assign n_6684 = ~n_6682 & ~n_6683;
assign n_6685 =  n_6681 &  n_6684;
assign n_6686 = ~x_2231 &  n_463;
assign n_6687 = ~x_2237 &  n_460;
assign n_6688 = ~n_6686 & ~n_6687;
assign n_6689 = ~x_2233 &  n_466;
assign n_6690 = ~x_2235 &  n_468;
assign n_6691 = ~n_6689 & ~n_6690;
assign n_6692 =  n_6688 &  n_6691;
assign n_6693 =  n_6685 &  n_6692;
assign n_6694 =  x_231 &  n_6693;
assign n_6695 = ~n_6678 & ~n_6694;
assign n_6696 = ~x_1470 & ~n_6695;
assign n_6697 = ~n_6677 & ~n_6696;
assign n_6698 =  n_1713 & ~n_6697;
assign n_6699 =  x_1185 & ~n_436;
assign n_6700 =  n_436 &  n_6693;
assign n_6701 = ~n_6699 & ~n_6700;
assign n_6702 =  n_1321 & ~n_6701;
assign n_6703 = ~n_6698 & ~n_6702;
assign n_6704 = ~n_6146 & ~n_6703;
assign n_6705 =  x_3210 &  n_6146;
assign n_6706 = ~n_6704 & ~n_6705;
assign n_6707 =  x_3210 & ~n_6706;
assign n_6708 = ~x_3210 &  n_6706;
assign n_6709 = ~n_6707 & ~n_6708;
assign n_6710 = ~x_230 & ~x_1122;
assign n_6711 = ~x_1122 &  n_1126;
assign n_6712 = ~x_2228 &  n_441;
assign n_6713 = ~x_2224 &  n_449;
assign n_6714 = ~n_6712 & ~n_6713;
assign n_6715 = ~x_2226 &  n_444;
assign n_6716 = ~x_2222 &  n_447;
assign n_6717 = ~n_6715 & ~n_6716;
assign n_6718 =  n_6714 &  n_6717;
assign n_6719 = ~x_2227 &  n_468;
assign n_6720 = ~x_2229 &  n_460;
assign n_6721 = ~n_6719 & ~n_6720;
assign n_6722 = ~x_2225 &  n_466;
assign n_6723 = ~x_2223 &  n_463;
assign n_6724 = ~n_6722 & ~n_6723;
assign n_6725 =  n_6721 &  n_6724;
assign n_6726 =  n_6718 &  n_6725;
assign n_6727 =  x_231 &  n_6726;
assign n_6728 = ~n_6711 & ~n_6727;
assign n_6729 = ~x_1470 & ~n_6728;
assign n_6730 = ~n_6710 & ~n_6729;
assign n_6731 =  n_1713 & ~n_6730;
assign n_6732 =  x_1184 & ~n_436;
assign n_6733 =  n_436 &  n_6726;
assign n_6734 = ~n_6732 & ~n_6733;
assign n_6735 =  n_1321 & ~n_6734;
assign n_6736 = ~n_6731 & ~n_6735;
assign n_6737 = ~n_6146 & ~n_6736;
assign n_6738 =  x_3209 &  n_6146;
assign n_6739 = ~n_6737 & ~n_6738;
assign n_6740 =  x_3209 & ~n_6739;
assign n_6741 = ~x_3209 &  n_6739;
assign n_6742 = ~n_6740 & ~n_6741;
assign n_6743 = ~x_230 & ~x_1121;
assign n_6744 = ~x_1121 &  n_1126;
assign n_6745 = ~x_2220 &  n_441;
assign n_6746 = ~x_2216 &  n_449;
assign n_6747 = ~n_6745 & ~n_6746;
assign n_6748 = ~x_2218 &  n_444;
assign n_6749 = ~x_2214 &  n_447;
assign n_6750 = ~n_6748 & ~n_6749;
assign n_6751 =  n_6747 &  n_6750;
assign n_6752 = ~x_2219 &  n_468;
assign n_6753 = ~x_2221 &  n_460;
assign n_6754 = ~n_6752 & ~n_6753;
assign n_6755 = ~x_2215 &  n_463;
assign n_6756 = ~x_2217 &  n_466;
assign n_6757 = ~n_6755 & ~n_6756;
assign n_6758 =  n_6754 &  n_6757;
assign n_6759 =  n_6751 &  n_6758;
assign n_6760 =  x_231 &  n_6759;
assign n_6761 = ~n_6744 & ~n_6760;
assign n_6762 = ~x_1470 & ~n_6761;
assign n_6763 = ~n_6743 & ~n_6762;
assign n_6764 =  n_1713 & ~n_6763;
assign n_6765 =  x_1183 & ~n_436;
assign n_6766 =  n_436 &  n_6759;
assign n_6767 = ~n_6765 & ~n_6766;
assign n_6768 =  n_1321 & ~n_6767;
assign n_6769 = ~n_6764 & ~n_6768;
assign n_6770 = ~n_6146 & ~n_6769;
assign n_6771 =  x_3208 &  n_6146;
assign n_6772 = ~n_6770 & ~n_6771;
assign n_6773 =  x_3208 & ~n_6772;
assign n_6774 = ~x_3208 &  n_6772;
assign n_6775 = ~n_6773 & ~n_6774;
assign n_6776 = ~x_230 & ~x_1120;
assign n_6777 = ~x_1120 &  n_1126;
assign n_6778 = ~x_2210 &  n_444;
assign n_6779 = ~x_2208 &  n_449;
assign n_6780 = ~n_6778 & ~n_6779;
assign n_6781 = ~x_2212 &  n_441;
assign n_6782 = ~x_2206 &  n_447;
assign n_6783 = ~n_6781 & ~n_6782;
assign n_6784 =  n_6780 &  n_6783;
assign n_6785 = ~x_2209 &  n_466;
assign n_6786 = ~x_2211 &  n_468;
assign n_6787 = ~n_6785 & ~n_6786;
assign n_6788 = ~x_2213 &  n_460;
assign n_6789 = ~x_2207 &  n_463;
assign n_6790 = ~n_6788 & ~n_6789;
assign n_6791 =  n_6787 &  n_6790;
assign n_6792 =  n_6784 &  n_6791;
assign n_6793 =  x_231 &  n_6792;
assign n_6794 = ~n_6777 & ~n_6793;
assign n_6795 = ~x_1470 & ~n_6794;
assign n_6796 = ~n_6776 & ~n_6795;
assign n_6797 =  n_1713 & ~n_6796;
assign n_6798 =  x_1182 & ~n_436;
assign n_6799 =  n_436 &  n_6792;
assign n_6800 = ~n_6798 & ~n_6799;
assign n_6801 =  n_1321 & ~n_6800;
assign n_6802 = ~n_6797 & ~n_6801;
assign n_6803 = ~n_6146 & ~n_6802;
assign n_6804 =  x_3207 &  n_6146;
assign n_6805 = ~n_6803 & ~n_6804;
assign n_6806 =  x_3207 & ~n_6805;
assign n_6807 = ~x_3207 &  n_6805;
assign n_6808 = ~n_6806 & ~n_6807;
assign n_6809 = ~x_230 & ~x_1119;
assign n_6810 = ~x_1119 &  n_1126;
assign n_6811 = ~x_2200 &  n_449;
assign n_6812 = ~x_2202 &  n_444;
assign n_6813 = ~n_6811 & ~n_6812;
assign n_6814 = ~x_2204 &  n_441;
assign n_6815 = ~x_2198 &  n_447;
assign n_6816 = ~n_6814 & ~n_6815;
assign n_6817 =  n_6813 &  n_6816;
assign n_6818 = ~x_2203 &  n_468;
assign n_6819 = ~x_2205 &  n_460;
assign n_6820 = ~n_6818 & ~n_6819;
assign n_6821 = ~x_2199 &  n_463;
assign n_6822 = ~x_2201 &  n_466;
assign n_6823 = ~n_6821 & ~n_6822;
assign n_6824 =  n_6820 &  n_6823;
assign n_6825 =  n_6817 &  n_6824;
assign n_6826 =  x_231 &  n_6825;
assign n_6827 = ~n_6810 & ~n_6826;
assign n_6828 = ~x_1470 & ~n_6827;
assign n_6829 = ~n_6809 & ~n_6828;
assign n_6830 =  n_1713 & ~n_6829;
assign n_6831 =  x_1181 & ~n_436;
assign n_6832 =  n_436 &  n_6825;
assign n_6833 = ~n_6831 & ~n_6832;
assign n_6834 =  n_1321 & ~n_6833;
assign n_6835 = ~n_6830 & ~n_6834;
assign n_6836 = ~n_6146 & ~n_6835;
assign n_6837 =  x_3206 &  n_6146;
assign n_6838 = ~n_6836 & ~n_6837;
assign n_6839 =  x_3206 & ~n_6838;
assign n_6840 = ~x_3206 &  n_6838;
assign n_6841 = ~n_6839 & ~n_6840;
assign n_6842 = ~x_230 & ~x_1118;
assign n_6843 = ~x_1118 &  n_1126;
assign n_6844 = ~x_2196 &  n_441;
assign n_6845 = ~x_2192 &  n_449;
assign n_6846 = ~n_6844 & ~n_6845;
assign n_6847 = ~x_2194 &  n_444;
assign n_6848 = ~x_2190 &  n_447;
assign n_6849 = ~n_6847 & ~n_6848;
assign n_6850 =  n_6846 &  n_6849;
assign n_6851 = ~x_2191 &  n_463;
assign n_6852 = ~x_2195 &  n_468;
assign n_6853 = ~n_6851 & ~n_6852;
assign n_6854 = ~x_2193 &  n_466;
assign n_6855 = ~x_2197 &  n_460;
assign n_6856 = ~n_6854 & ~n_6855;
assign n_6857 =  n_6853 &  n_6856;
assign n_6858 =  n_6850 &  n_6857;
assign n_6859 =  x_231 &  n_6858;
assign n_6860 = ~n_6843 & ~n_6859;
assign n_6861 = ~x_1470 & ~n_6860;
assign n_6862 = ~n_6842 & ~n_6861;
assign n_6863 =  n_1713 & ~n_6862;
assign n_6864 =  x_1180 & ~n_436;
assign n_6865 =  n_436 &  n_6858;
assign n_6866 = ~n_6864 & ~n_6865;
assign n_6867 =  n_1321 & ~n_6866;
assign n_6868 = ~n_6863 & ~n_6867;
assign n_6869 = ~n_6146 & ~n_6868;
assign n_6870 =  x_3205 &  n_6146;
assign n_6871 = ~n_6869 & ~n_6870;
assign n_6872 =  x_3205 & ~n_6871;
assign n_6873 = ~x_3205 &  n_6871;
assign n_6874 = ~n_6872 & ~n_6873;
assign n_6875 = ~x_230 & ~x_1117;
assign n_6876 = ~x_1117 &  n_1126;
assign n_6877 = ~x_2188 &  n_441;
assign n_6878 = ~x_2184 &  n_449;
assign n_6879 = ~n_6877 & ~n_6878;
assign n_6880 = ~x_2186 &  n_444;
assign n_6881 = ~x_2182 &  n_447;
assign n_6882 = ~n_6880 & ~n_6881;
assign n_6883 =  n_6879 &  n_6882;
assign n_6884 = ~x_2187 &  n_468;
assign n_6885 = ~x_2189 &  n_460;
assign n_6886 = ~n_6884 & ~n_6885;
assign n_6887 = ~x_2185 &  n_466;
assign n_6888 = ~x_2183 &  n_463;
assign n_6889 = ~n_6887 & ~n_6888;
assign n_6890 =  n_6886 &  n_6889;
assign n_6891 =  n_6883 &  n_6890;
assign n_6892 =  x_231 &  n_6891;
assign n_6893 = ~n_6876 & ~n_6892;
assign n_6894 = ~x_1470 & ~n_6893;
assign n_6895 = ~n_6875 & ~n_6894;
assign n_6896 =  n_1713 & ~n_6895;
assign n_6897 =  x_1179 & ~n_436;
assign n_6898 =  n_436 &  n_6891;
assign n_6899 = ~n_6897 & ~n_6898;
assign n_6900 =  n_1321 & ~n_6899;
assign n_6901 = ~n_6896 & ~n_6900;
assign n_6902 = ~n_6146 & ~n_6901;
assign n_6903 =  x_3204 &  n_6146;
assign n_6904 = ~n_6902 & ~n_6903;
assign n_6905 =  x_3204 & ~n_6904;
assign n_6906 = ~x_3204 &  n_6904;
assign n_6907 = ~n_6905 & ~n_6906;
assign n_6908 = ~x_230 & ~x_1116;
assign n_6909 = ~x_1116 &  n_1126;
assign n_6910 = ~x_2174 &  n_447;
assign n_6911 = ~x_2180 &  n_441;
assign n_6912 = ~n_6910 & ~n_6911;
assign n_6913 = ~x_2178 &  n_444;
assign n_6914 = ~x_2176 &  n_449;
assign n_6915 = ~n_6913 & ~n_6914;
assign n_6916 =  n_6912 &  n_6915;
assign n_6917 = ~x_2179 &  n_468;
assign n_6918 = ~x_2177 &  n_466;
assign n_6919 = ~n_6917 & ~n_6918;
assign n_6920 = ~x_2181 &  n_460;
assign n_6921 = ~x_2175 &  n_463;
assign n_6922 = ~n_6920 & ~n_6921;
assign n_6923 =  n_6919 &  n_6922;
assign n_6924 =  n_6916 &  n_6923;
assign n_6925 =  x_231 &  n_6924;
assign n_6926 = ~n_6909 & ~n_6925;
assign n_6927 = ~x_1470 & ~n_6926;
assign n_6928 = ~n_6908 & ~n_6927;
assign n_6929 =  n_1713 & ~n_6928;
assign n_6930 =  x_1178 & ~n_436;
assign n_6931 =  n_436 &  n_6924;
assign n_6932 = ~n_6930 & ~n_6931;
assign n_6933 =  n_1321 & ~n_6932;
assign n_6934 = ~n_6929 & ~n_6933;
assign n_6935 =  x_3203 &  n_6934;
assign n_6936 = ~x_3203 & ~n_6934;
assign n_6937 = ~n_6935 & ~n_6936;
assign n_6938 =  n_6146 & ~n_4192;
assign n_6939 =  x_3202 & ~n_6938;
assign n_6940 = ~x_3202 &  n_6938;
assign n_6941 = ~n_6939 & ~n_6940;
assign n_6942 = ~x_230 & ~x_1115;
assign n_6943 = ~x_1115 &  n_1126;
assign n_6944 = ~x_2166 &  n_447;
assign n_6945 = ~x_2168 &  n_449;
assign n_6946 = ~n_6944 & ~n_6945;
assign n_6947 = ~x_2172 &  n_441;
assign n_6948 = ~x_2170 &  n_444;
assign n_6949 = ~n_6947 & ~n_6948;
assign n_6950 =  n_6946 &  n_6949;
assign n_6951 = ~x_2169 &  n_466;
assign n_6952 = ~x_2171 &  n_468;
assign n_6953 = ~n_6951 & ~n_6952;
assign n_6954 = ~x_2173 &  n_460;
assign n_6955 = ~x_2167 &  n_463;
assign n_6956 = ~n_6954 & ~n_6955;
assign n_6957 =  n_6953 &  n_6956;
assign n_6958 =  n_6950 &  n_6957;
assign n_6959 =  x_231 &  n_6958;
assign n_6960 = ~n_6943 & ~n_6959;
assign n_6961 = ~x_1470 & ~n_6960;
assign n_6962 = ~n_6942 & ~n_6961;
assign n_6963 =  n_1713 & ~n_6962;
assign n_6964 =  x_1177 & ~n_436;
assign n_6965 =  n_436 &  n_6958;
assign n_6966 = ~n_6964 & ~n_6965;
assign n_6967 =  n_1321 & ~n_6966;
assign n_6968 = ~n_6963 & ~n_6967;
assign n_6969 = ~n_6146 & ~n_6968;
assign n_6970 =  x_3201 &  n_6146;
assign n_6971 = ~n_6969 & ~n_6970;
assign n_6972 =  x_3201 & ~n_6971;
assign n_6973 = ~x_3201 &  n_6971;
assign n_6974 = ~n_6972 & ~n_6973;
assign n_6975 = ~x_230 & ~x_1114;
assign n_6976 = ~x_1114 &  n_1126;
assign n_6977 = ~x_2158 &  n_447;
assign n_6978 = ~x_2164 &  n_441;
assign n_6979 = ~n_6977 & ~n_6978;
assign n_6980 = ~x_2160 &  n_449;
assign n_6981 = ~x_2162 &  n_444;
assign n_6982 = ~n_6980 & ~n_6981;
assign n_6983 =  n_6979 &  n_6982;
assign n_6984 = ~x_2165 &  n_460;
assign n_6985 = ~x_2159 &  n_463;
assign n_6986 = ~n_6984 & ~n_6985;
assign n_6987 = ~x_2161 &  n_466;
assign n_6988 = ~x_2163 &  n_468;
assign n_6989 = ~n_6987 & ~n_6988;
assign n_6990 =  n_6986 &  n_6989;
assign n_6991 =  n_6983 &  n_6990;
assign n_6992 =  x_231 &  n_6991;
assign n_6993 = ~n_6976 & ~n_6992;
assign n_6994 = ~x_1470 & ~n_6993;
assign n_6995 = ~n_6975 & ~n_6994;
assign n_6996 =  n_1713 & ~n_6995;
assign n_6997 =  x_1176 & ~n_436;
assign n_6998 =  n_436 &  n_6991;
assign n_6999 = ~n_6997 & ~n_6998;
assign n_7000 =  n_1321 & ~n_6999;
assign n_7001 = ~n_6996 & ~n_7000;
assign n_7002 = ~n_6146 & ~n_7001;
assign n_7003 =  x_3200 &  n_6146;
assign n_7004 = ~n_7002 & ~n_7003;
assign n_7005 =  x_3200 & ~n_7004;
assign n_7006 = ~x_3200 &  n_7004;
assign n_7007 = ~n_7005 & ~n_7006;
assign n_7008 = ~x_230 & ~x_1113;
assign n_7009 = ~x_1113 &  n_1126;
assign n_7010 = ~x_2156 &  n_441;
assign n_7011 = ~x_2154 &  n_444;
assign n_7012 = ~n_7010 & ~n_7011;
assign n_7013 = ~x_2152 &  n_449;
assign n_7014 = ~x_2150 &  n_447;
assign n_7015 = ~n_7013 & ~n_7014;
assign n_7016 =  n_7012 &  n_7015;
assign n_7017 = ~x_2157 &  n_460;
assign n_7018 = ~x_2153 &  n_466;
assign n_7019 = ~n_7017 & ~n_7018;
assign n_7020 = ~x_2151 &  n_463;
assign n_7021 = ~x_2155 &  n_468;
assign n_7022 = ~n_7020 & ~n_7021;
assign n_7023 =  n_7019 &  n_7022;
assign n_7024 =  n_7016 &  n_7023;
assign n_7025 =  x_231 &  n_7024;
assign n_7026 = ~n_7009 & ~n_7025;
assign n_7027 = ~x_1470 & ~n_7026;
assign n_7028 = ~n_7008 & ~n_7027;
assign n_7029 =  n_1713 & ~n_7028;
assign n_7030 =  x_1175 & ~n_436;
assign n_7031 =  n_436 &  n_7024;
assign n_7032 = ~n_7030 & ~n_7031;
assign n_7033 =  n_1321 & ~n_7032;
assign n_7034 = ~n_7029 & ~n_7033;
assign n_7035 = ~n_6146 & ~n_7034;
assign n_7036 =  x_3199 &  n_6146;
assign n_7037 = ~n_7035 & ~n_7036;
assign n_7038 =  x_3199 & ~n_7037;
assign n_7039 = ~x_3199 &  n_7037;
assign n_7040 = ~n_7038 & ~n_7039;
assign n_7041 = ~x_230 & ~x_1112;
assign n_7042 = ~x_1112 &  n_1126;
assign n_7043 = ~x_2142 &  n_447;
assign n_7044 = ~x_2146 &  n_444;
assign n_7045 = ~n_7043 & ~n_7044;
assign n_7046 = ~x_2148 &  n_441;
assign n_7047 = ~x_2144 &  n_449;
assign n_7048 = ~n_7046 & ~n_7047;
assign n_7049 =  n_7045 &  n_7048;
assign n_7050 = ~x_2143 &  n_463;
assign n_7051 = ~x_2147 &  n_468;
assign n_7052 = ~n_7050 & ~n_7051;
assign n_7053 = ~x_2145 &  n_466;
assign n_7054 = ~x_2149 &  n_460;
assign n_7055 = ~n_7053 & ~n_7054;
assign n_7056 =  n_7052 &  n_7055;
assign n_7057 =  n_7049 &  n_7056;
assign n_7058 =  x_231 &  n_7057;
assign n_7059 = ~n_7042 & ~n_7058;
assign n_7060 = ~x_1470 & ~n_7059;
assign n_7061 = ~n_7041 & ~n_7060;
assign n_7062 =  n_1713 & ~n_7061;
assign n_7063 =  x_1174 & ~n_436;
assign n_7064 =  n_436 &  n_7057;
assign n_7065 = ~n_7063 & ~n_7064;
assign n_7066 =  n_1321 & ~n_7065;
assign n_7067 = ~n_7062 & ~n_7066;
assign n_7068 = ~n_6146 & ~n_7067;
assign n_7069 =  x_3198 &  n_6146;
assign n_7070 = ~n_7068 & ~n_7069;
assign n_7071 =  x_3198 & ~n_7070;
assign n_7072 = ~x_3198 &  n_7070;
assign n_7073 = ~n_7071 & ~n_7072;
assign n_7074 = ~x_230 & ~x_1111;
assign n_7075 = ~x_1111 &  n_1126;
assign n_7076 = ~x_2138 &  n_444;
assign n_7077 = ~x_2140 &  n_441;
assign n_7078 = ~n_7076 & ~n_7077;
assign n_7079 = ~x_2134 &  n_447;
assign n_7080 = ~x_2136 &  n_449;
assign n_7081 = ~n_7079 & ~n_7080;
assign n_7082 =  n_7078 &  n_7081;
assign n_7083 = ~x_2135 &  n_463;
assign n_7084 = ~x_2137 &  n_466;
assign n_7085 = ~n_7083 & ~n_7084;
assign n_7086 = ~x_2141 &  n_460;
assign n_7087 = ~x_2139 &  n_468;
assign n_7088 = ~n_7086 & ~n_7087;
assign n_7089 =  n_7085 &  n_7088;
assign n_7090 =  n_7082 &  n_7089;
assign n_7091 =  x_231 &  n_7090;
assign n_7092 = ~n_7075 & ~n_7091;
assign n_7093 = ~x_1470 & ~n_7092;
assign n_7094 = ~n_7074 & ~n_7093;
assign n_7095 =  n_1713 & ~n_7094;
assign n_7096 =  x_1173 & ~n_436;
assign n_7097 =  n_436 &  n_7090;
assign n_7098 = ~n_7096 & ~n_7097;
assign n_7099 =  n_1321 & ~n_7098;
assign n_7100 = ~n_7095 & ~n_7099;
assign n_7101 = ~n_6146 & ~n_7100;
assign n_7102 =  x_3197 &  n_6146;
assign n_7103 = ~n_7101 & ~n_7102;
assign n_7104 =  x_3197 & ~n_7103;
assign n_7105 = ~x_3197 &  n_7103;
assign n_7106 = ~n_7104 & ~n_7105;
assign n_7107 = ~x_230 & ~x_1110;
assign n_7108 = ~x_1110 &  n_1126;
assign n_7109 = ~x_2132 &  n_441;
assign n_7110 = ~x_2130 &  n_444;
assign n_7111 = ~n_7109 & ~n_7110;
assign n_7112 = ~x_2128 &  n_449;
assign n_7113 = ~x_2126 &  n_447;
assign n_7114 = ~n_7112 & ~n_7113;
assign n_7115 =  n_7111 &  n_7114;
assign n_7116 = ~x_2129 &  n_466;
assign n_7117 = ~x_2127 &  n_463;
assign n_7118 = ~n_7116 & ~n_7117;
assign n_7119 = ~x_2131 &  n_468;
assign n_7120 = ~x_2133 &  n_460;
assign n_7121 = ~n_7119 & ~n_7120;
assign n_7122 =  n_7118 &  n_7121;
assign n_7123 =  n_7115 &  n_7122;
assign n_7124 =  x_231 &  n_7123;
assign n_7125 = ~n_7108 & ~n_7124;
assign n_7126 = ~x_1470 & ~n_7125;
assign n_7127 = ~n_7107 & ~n_7126;
assign n_7128 =  n_1713 & ~n_7127;
assign n_7129 =  x_1172 & ~n_436;
assign n_7130 =  n_436 &  n_7123;
assign n_7131 = ~n_7129 & ~n_7130;
assign n_7132 =  n_1321 & ~n_7131;
assign n_7133 = ~n_7128 & ~n_7132;
assign n_7134 = ~n_6146 & ~n_7133;
assign n_7135 =  x_3196 &  n_6146;
assign n_7136 = ~n_7134 & ~n_7135;
assign n_7137 =  x_3196 & ~n_7136;
assign n_7138 = ~x_3196 &  n_7136;
assign n_7139 = ~n_7137 & ~n_7138;
assign n_7140 = ~x_230 & ~x_1109;
assign n_7141 = ~x_1109 &  n_1126;
assign n_7142 = ~x_2118 &  n_447;
assign n_7143 = ~x_2124 &  n_441;
assign n_7144 = ~n_7142 & ~n_7143;
assign n_7145 = ~x_2122 &  n_444;
assign n_7146 = ~x_2120 &  n_449;
assign n_7147 = ~n_7145 & ~n_7146;
assign n_7148 =  n_7144 &  n_7147;
assign n_7149 = ~x_2125 &  n_460;
assign n_7150 = ~x_2123 &  n_468;
assign n_7151 = ~n_7149 & ~n_7150;
assign n_7152 = ~x_2119 &  n_463;
assign n_7153 = ~x_2121 &  n_466;
assign n_7154 = ~n_7152 & ~n_7153;
assign n_7155 =  n_7151 &  n_7154;
assign n_7156 =  n_7148 &  n_7155;
assign n_7157 =  x_231 &  n_7156;
assign n_7158 = ~n_7141 & ~n_7157;
assign n_7159 = ~x_1470 & ~n_7158;
assign n_7160 = ~n_7140 & ~n_7159;
assign n_7161 =  n_1713 & ~n_7160;
assign n_7162 =  x_1171 & ~n_436;
assign n_7163 =  n_436 &  n_7156;
assign n_7164 = ~n_7162 & ~n_7163;
assign n_7165 =  n_1321 & ~n_7164;
assign n_7166 = ~n_7161 & ~n_7165;
assign n_7167 = ~n_6146 & ~n_7166;
assign n_7168 =  x_3195 &  n_6146;
assign n_7169 = ~n_7167 & ~n_7168;
assign n_7170 =  x_3195 & ~n_7169;
assign n_7171 = ~x_3195 &  n_7169;
assign n_7172 = ~n_7170 & ~n_7171;
assign n_7173 =  x_1170 & ~n_436;
assign n_7174 = ~x_2116 &  n_441;
assign n_7175 = ~x_2112 &  n_449;
assign n_7176 = ~n_7174 & ~n_7175;
assign n_7177 = ~x_2114 &  n_444;
assign n_7178 = ~x_2110 &  n_447;
assign n_7179 = ~n_7177 & ~n_7178;
assign n_7180 =  n_7176 &  n_7179;
assign n_7181 = ~x_2115 &  n_468;
assign n_7182 = ~x_2117 &  n_460;
assign n_7183 = ~n_7181 & ~n_7182;
assign n_7184 = ~x_2111 &  n_463;
assign n_7185 = ~x_2113 &  n_466;
assign n_7186 = ~n_7184 & ~n_7185;
assign n_7187 =  n_7183 &  n_7186;
assign n_7188 =  n_7180 &  n_7187;
assign n_7189 =  n_436 &  n_7188;
assign n_7190 = ~n_7173 & ~n_7189;
assign n_7191 =  n_1321 & ~n_7190;
assign n_7192 = ~x_230 & ~x_1108;
assign n_7193 = ~x_1108 &  n_1126;
assign n_7194 =  x_231 &  n_7188;
assign n_7195 = ~n_7193 & ~n_7194;
assign n_7196 = ~x_1470 & ~n_7195;
assign n_7197 = ~n_7192 & ~n_7196;
assign n_7198 =  n_1713 & ~n_7197;
assign n_7199 = ~n_7191 & ~n_7198;
assign n_7200 =  x_3194 &  n_7199;
assign n_7201 = ~x_3194 & ~n_7199;
assign n_7202 = ~n_7200 & ~n_7201;
assign n_7203 =  n_6146 & ~n_4068;
assign n_7204 =  x_3193 & ~n_7203;
assign n_7205 = ~x_3193 &  n_7203;
assign n_7206 = ~n_7204 & ~n_7205;
assign n_7207 = ~x_230 & ~x_1107;
assign n_7208 = ~x_1107 &  n_1126;
assign n_7209 = ~x_2102 &  n_447;
assign n_7210 = ~x_2106 &  n_444;
assign n_7211 = ~n_7209 & ~n_7210;
assign n_7212 = ~x_2104 &  n_449;
assign n_7213 = ~x_2108 &  n_441;
assign n_7214 = ~n_7212 & ~n_7213;
assign n_7215 =  n_7211 &  n_7214;
assign n_7216 = ~x_2103 &  n_463;
assign n_7217 = ~x_2105 &  n_466;
assign n_7218 = ~n_7216 & ~n_7217;
assign n_7219 = ~x_2107 &  n_468;
assign n_7220 = ~x_2109 &  n_460;
assign n_7221 = ~n_7219 & ~n_7220;
assign n_7222 =  n_7218 &  n_7221;
assign n_7223 =  n_7215 &  n_7222;
assign n_7224 =  x_231 &  n_7223;
assign n_7225 = ~n_7208 & ~n_7224;
assign n_7226 = ~x_1470 & ~n_7225;
assign n_7227 = ~n_7207 & ~n_7226;
assign n_7228 =  n_1713 & ~n_7227;
assign n_7229 =  x_1169 & ~n_436;
assign n_7230 =  n_436 &  n_7223;
assign n_7231 = ~n_7229 & ~n_7230;
assign n_7232 =  n_1321 & ~n_7231;
assign n_7233 = ~n_7228 & ~n_7232;
assign n_7234 = ~n_6146 & ~n_7233;
assign n_7235 =  x_3192 &  n_6146;
assign n_7236 = ~n_7234 & ~n_7235;
assign n_7237 =  x_3192 & ~n_7236;
assign n_7238 = ~x_3192 &  n_7236;
assign n_7239 = ~n_7237 & ~n_7238;
assign n_7240 = ~x_230 & ~x_1106;
assign n_7241 = ~x_1106 &  n_1126;
assign n_7242 = ~x_2094 &  n_447;
assign n_7243 = ~x_2098 &  n_444;
assign n_7244 = ~n_7242 & ~n_7243;
assign n_7245 = ~x_2096 &  n_449;
assign n_7246 = ~x_2100 &  n_441;
assign n_7247 = ~n_7245 & ~n_7246;
assign n_7248 =  n_7244 &  n_7247;
assign n_7249 = ~x_2095 &  n_463;
assign n_7250 = ~x_2101 &  n_460;
assign n_7251 = ~n_7249 & ~n_7250;
assign n_7252 = ~x_2097 &  n_466;
assign n_7253 = ~x_2099 &  n_468;
assign n_7254 = ~n_7252 & ~n_7253;
assign n_7255 =  n_7251 &  n_7254;
assign n_7256 =  n_7248 &  n_7255;
assign n_7257 =  x_231 &  n_7256;
assign n_7258 = ~n_7241 & ~n_7257;
assign n_7259 = ~x_1470 & ~n_7258;
assign n_7260 = ~n_7240 & ~n_7259;
assign n_7261 =  n_1713 & ~n_7260;
assign n_7262 =  x_1168 & ~n_436;
assign n_7263 =  n_436 &  n_7256;
assign n_7264 = ~n_7262 & ~n_7263;
assign n_7265 =  n_1321 & ~n_7264;
assign n_7266 = ~n_7261 & ~n_7265;
assign n_7267 = ~n_6146 & ~n_7266;
assign n_7268 =  x_3191 &  n_6146;
assign n_7269 = ~n_7267 & ~n_7268;
assign n_7270 =  x_3191 & ~n_7269;
assign n_7271 = ~x_3191 &  n_7269;
assign n_7272 = ~n_7270 & ~n_7271;
assign n_7273 = ~x_230 & ~x_1105;
assign n_7274 = ~x_1105 &  n_1126;
assign n_7275 = ~x_2088 &  n_449;
assign n_7276 = ~x_2090 &  n_444;
assign n_7277 = ~n_7275 & ~n_7276;
assign n_7278 = ~x_2092 &  n_441;
assign n_7279 = ~x_2086 &  n_447;
assign n_7280 = ~n_7278 & ~n_7279;
assign n_7281 =  n_7277 &  n_7280;
assign n_7282 = ~x_2091 &  n_468;
assign n_7283 = ~x_2093 &  n_460;
assign n_7284 = ~n_7282 & ~n_7283;
assign n_7285 = ~x_2087 &  n_463;
assign n_7286 = ~x_2089 &  n_466;
assign n_7287 = ~n_7285 & ~n_7286;
assign n_7288 =  n_7284 &  n_7287;
assign n_7289 =  n_7281 &  n_7288;
assign n_7290 =  x_231 &  n_7289;
assign n_7291 = ~n_7274 & ~n_7290;
assign n_7292 = ~x_1470 & ~n_7291;
assign n_7293 = ~n_7273 & ~n_7292;
assign n_7294 =  n_1713 & ~n_7293;
assign n_7295 =  x_1167 & ~n_436;
assign n_7296 =  n_436 &  n_7289;
assign n_7297 = ~n_7295 & ~n_7296;
assign n_7298 =  n_1321 & ~n_7297;
assign n_7299 = ~n_7294 & ~n_7298;
assign n_7300 = ~n_6146 & ~n_7299;
assign n_7301 =  x_3190 &  n_6146;
assign n_7302 = ~n_7300 & ~n_7301;
assign n_7303 =  x_3190 & ~n_7302;
assign n_7304 = ~x_3190 &  n_7302;
assign n_7305 = ~n_7303 & ~n_7304;
assign n_7306 = ~x_230 & ~x_1104;
assign n_7307 = ~x_1104 &  n_1126;
assign n_7308 = ~x_2078 &  n_447;
assign n_7309 = ~x_2080 &  n_449;
assign n_7310 = ~n_7308 & ~n_7309;
assign n_7311 = ~x_2084 &  n_441;
assign n_7312 = ~x_2082 &  n_444;
assign n_7313 = ~n_7311 & ~n_7312;
assign n_7314 =  n_7310 &  n_7313;
assign n_7315 = ~x_2081 &  n_466;
assign n_7316 = ~x_2083 &  n_468;
assign n_7317 = ~n_7315 & ~n_7316;
assign n_7318 = ~x_2085 &  n_460;
assign n_7319 = ~x_2079 &  n_463;
assign n_7320 = ~n_7318 & ~n_7319;
assign n_7321 =  n_7317 &  n_7320;
assign n_7322 =  n_7314 &  n_7321;
assign n_7323 =  x_231 &  n_7322;
assign n_7324 = ~n_7307 & ~n_7323;
assign n_7325 = ~x_1470 & ~n_7324;
assign n_7326 = ~n_7306 & ~n_7325;
assign n_7327 =  n_1713 & ~n_7326;
assign n_7328 =  x_1166 & ~n_436;
assign n_7329 =  n_436 &  n_7322;
assign n_7330 = ~n_7328 & ~n_7329;
assign n_7331 =  n_1321 & ~n_7330;
assign n_7332 = ~n_7327 & ~n_7331;
assign n_7333 = ~n_6146 & ~n_7332;
assign n_7334 =  x_3189 &  n_6146;
assign n_7335 = ~n_7333 & ~n_7334;
assign n_7336 =  x_3189 & ~n_7335;
assign n_7337 = ~x_3189 &  n_7335;
assign n_7338 = ~n_7336 & ~n_7337;
assign n_7339 = ~x_230 & ~x_1103;
assign n_7340 = ~x_1103 &  n_1126;
assign n_7341 = ~x_2074 &  n_444;
assign n_7342 = ~x_2076 &  n_441;
assign n_7343 = ~n_7341 & ~n_7342;
assign n_7344 = ~x_2072 &  n_449;
assign n_7345 = ~x_2070 &  n_447;
assign n_7346 = ~n_7344 & ~n_7345;
assign n_7347 =  n_7343 &  n_7346;
assign n_7348 = ~x_2075 &  n_468;
assign n_7349 = ~x_2077 &  n_460;
assign n_7350 = ~n_7348 & ~n_7349;
assign n_7351 = ~x_2073 &  n_466;
assign n_7352 = ~x_2071 &  n_463;
assign n_7353 = ~n_7351 & ~n_7352;
assign n_7354 =  n_7350 &  n_7353;
assign n_7355 =  n_7347 &  n_7354;
assign n_7356 =  x_231 &  n_7355;
assign n_7357 = ~n_7340 & ~n_7356;
assign n_7358 = ~x_1470 & ~n_7357;
assign n_7359 = ~n_7339 & ~n_7358;
assign n_7360 =  n_1713 & ~n_7359;
assign n_7361 =  x_1165 & ~n_436;
assign n_7362 =  n_436 &  n_7355;
assign n_7363 = ~n_7361 & ~n_7362;
assign n_7364 =  n_1321 & ~n_7363;
assign n_7365 = ~n_7360 & ~n_7364;
assign n_7366 = ~n_6146 & ~n_7365;
assign n_7367 =  x_3188 &  n_6146;
assign n_7368 = ~n_7366 & ~n_7367;
assign n_7369 =  x_3188 & ~n_7368;
assign n_7370 = ~x_3188 &  n_7368;
assign n_7371 = ~n_7369 & ~n_7370;
assign n_7372 = ~x_230 & ~x_1102;
assign n_7373 = ~x_1102 &  n_1126;
assign n_7374 = ~x_2062 &  n_447;
assign n_7375 = ~x_2066 &  n_444;
assign n_7376 = ~n_7374 & ~n_7375;
assign n_7377 = ~x_2068 &  n_441;
assign n_7378 = ~x_2064 &  n_449;
assign n_7379 = ~n_7377 & ~n_7378;
assign n_7380 =  n_7376 &  n_7379;
assign n_7381 = ~x_2063 &  n_463;
assign n_7382 = ~x_2067 &  n_468;
assign n_7383 = ~n_7381 & ~n_7382;
assign n_7384 = ~x_2065 &  n_466;
assign n_7385 = ~x_2069 &  n_460;
assign n_7386 = ~n_7384 & ~n_7385;
assign n_7387 =  n_7383 &  n_7386;
assign n_7388 =  n_7380 &  n_7387;
assign n_7389 =  x_231 &  n_7388;
assign n_7390 = ~n_7373 & ~n_7389;
assign n_7391 = ~x_1470 & ~n_7390;
assign n_7392 = ~n_7372 & ~n_7391;
assign n_7393 =  n_1713 & ~n_7392;
assign n_7394 =  x_1164 & ~n_436;
assign n_7395 =  n_436 &  n_7388;
assign n_7396 = ~n_7394 & ~n_7395;
assign n_7397 =  n_1321 & ~n_7396;
assign n_7398 = ~n_7393 & ~n_7397;
assign n_7399 = ~n_6146 & ~n_7398;
assign n_7400 =  x_3187 &  n_6146;
assign n_7401 = ~n_7399 & ~n_7400;
assign n_7402 =  x_3187 & ~n_7401;
assign n_7403 = ~x_3187 &  n_7401;
assign n_7404 = ~n_7402 & ~n_7403;
assign n_7405 = ~x_230 & ~x_1101;
assign n_7406 = ~x_1101 &  n_1126;
assign n_7407 = ~x_2054 &  n_447;
assign n_7408 = ~x_2060 &  n_441;
assign n_7409 = ~n_7407 & ~n_7408;
assign n_7410 = ~x_2056 &  n_449;
assign n_7411 = ~x_2058 &  n_444;
assign n_7412 = ~n_7410 & ~n_7411;
assign n_7413 =  n_7409 &  n_7412;
assign n_7414 = ~x_2055 &  n_463;
assign n_7415 = ~x_2061 &  n_460;
assign n_7416 = ~n_7414 & ~n_7415;
assign n_7417 = ~x_2059 &  n_468;
assign n_7418 = ~x_2057 &  n_466;
assign n_7419 = ~n_7417 & ~n_7418;
assign n_7420 =  n_7416 &  n_7419;
assign n_7421 =  n_7413 &  n_7420;
assign n_7422 =  x_231 &  n_7421;
assign n_7423 = ~n_7406 & ~n_7422;
assign n_7424 = ~x_1470 & ~n_7423;
assign n_7425 = ~n_7405 & ~n_7424;
assign n_7426 =  n_1713 & ~n_7425;
assign n_7427 =  x_1163 & ~n_436;
assign n_7428 =  n_436 &  n_7421;
assign n_7429 = ~n_7427 & ~n_7428;
assign n_7430 =  n_1321 & ~n_7429;
assign n_7431 = ~n_7426 & ~n_7430;
assign n_7432 = ~n_6146 & ~n_7431;
assign n_7433 =  x_3186 &  n_6146;
assign n_7434 = ~n_7432 & ~n_7433;
assign n_7435 =  x_3186 & ~n_7434;
assign n_7436 = ~x_3186 &  n_7434;
assign n_7437 = ~n_7435 & ~n_7436;
assign n_7438 = ~x_230 & ~x_1100;
assign n_7439 = ~x_1100 &  n_1126;
assign n_7440 = ~x_2052 &  n_441;
assign n_7441 = ~x_2048 &  n_449;
assign n_7442 = ~n_7440 & ~n_7441;
assign n_7443 = ~x_2050 &  n_444;
assign n_7444 = ~x_2046 &  n_447;
assign n_7445 = ~n_7443 & ~n_7444;
assign n_7446 =  n_7442 &  n_7445;
assign n_7447 = ~x_2051 &  n_468;
assign n_7448 = ~x_2053 &  n_460;
assign n_7449 = ~n_7447 & ~n_7448;
assign n_7450 = ~x_2047 &  n_463;
assign n_7451 = ~x_2049 &  n_466;
assign n_7452 = ~n_7450 & ~n_7451;
assign n_7453 =  n_7449 &  n_7452;
assign n_7454 =  n_7446 &  n_7453;
assign n_7455 =  x_231 &  n_7454;
assign n_7456 = ~n_7439 & ~n_7455;
assign n_7457 = ~x_1470 & ~n_7456;
assign n_7458 = ~n_7438 & ~n_7457;
assign n_7459 =  n_1713 & ~n_7458;
assign n_7460 =  x_1162 & ~n_436;
assign n_7461 =  n_436 &  n_7454;
assign n_7462 = ~n_7460 & ~n_7461;
assign n_7463 =  n_1321 & ~n_7462;
assign n_7464 = ~n_7459 & ~n_7463;
assign n_7465 =  x_3185 &  n_7464;
assign n_7466 = ~x_3185 & ~n_7464;
assign n_7467 = ~n_7465 & ~n_7466;
assign n_7468 =  n_6146 & ~n_4178;
assign n_7469 =  x_3184 & ~n_7468;
assign n_7470 = ~x_3184 &  n_7468;
assign n_7471 = ~n_7469 & ~n_7470;
assign n_7472 = ~x_230 & ~x_1099;
assign n_7473 = ~x_1099 &  n_1126;
assign n_7474 = ~x_2038 &  n_447;
assign n_7475 = ~x_2040 &  n_449;
assign n_7476 = ~n_7474 & ~n_7475;
assign n_7477 = ~x_2042 &  n_444;
assign n_7478 = ~x_2044 &  n_441;
assign n_7479 = ~n_7477 & ~n_7478;
assign n_7480 =  n_7476 &  n_7479;
assign n_7481 = ~x_2043 &  n_468;
assign n_7482 = ~x_2045 &  n_460;
assign n_7483 = ~n_7481 & ~n_7482;
assign n_7484 = ~x_2039 &  n_463;
assign n_7485 = ~x_2041 &  n_466;
assign n_7486 = ~n_7484 & ~n_7485;
assign n_7487 =  n_7483 &  n_7486;
assign n_7488 =  n_7480 &  n_7487;
assign n_7489 =  x_231 &  n_7488;
assign n_7490 = ~n_7473 & ~n_7489;
assign n_7491 = ~x_1470 & ~n_7490;
assign n_7492 = ~n_7472 & ~n_7491;
assign n_7493 =  n_1713 & ~n_7492;
assign n_7494 =  x_1161 & ~n_436;
assign n_7495 =  n_436 &  n_7488;
assign n_7496 = ~n_7494 & ~n_7495;
assign n_7497 =  n_1321 & ~n_7496;
assign n_7498 = ~n_7493 & ~n_7497;
assign n_7499 = ~n_6146 & ~n_7498;
assign n_7500 =  x_3183 &  n_6146;
assign n_7501 = ~n_7499 & ~n_7500;
assign n_7502 =  x_3183 & ~n_7501;
assign n_7503 = ~x_3183 &  n_7501;
assign n_7504 = ~n_7502 & ~n_7503;
assign n_7505 = ~x_230 & ~x_1098;
assign n_7506 = ~x_1098 &  n_1126;
assign n_7507 = ~x_2030 &  n_447;
assign n_7508 = ~x_2034 &  n_444;
assign n_7509 = ~n_7507 & ~n_7508;
assign n_7510 = ~x_2036 &  n_441;
assign n_7511 = ~x_2032 &  n_449;
assign n_7512 = ~n_7510 & ~n_7511;
assign n_7513 =  n_7509 &  n_7512;
assign n_7514 = ~x_2031 &  n_463;
assign n_7515 = ~x_2035 &  n_468;
assign n_7516 = ~n_7514 & ~n_7515;
assign n_7517 = ~x_2033 &  n_466;
assign n_7518 = ~x_2037 &  n_460;
assign n_7519 = ~n_7517 & ~n_7518;
assign n_7520 =  n_7516 &  n_7519;
assign n_7521 =  n_7513 &  n_7520;
assign n_7522 =  x_231 &  n_7521;
assign n_7523 = ~n_7506 & ~n_7522;
assign n_7524 = ~x_1470 & ~n_7523;
assign n_7525 = ~n_7505 & ~n_7524;
assign n_7526 =  n_1713 & ~n_7525;
assign n_7527 =  x_1160 & ~n_436;
assign n_7528 =  n_436 &  n_7521;
assign n_7529 = ~n_7527 & ~n_7528;
assign n_7530 =  n_1321 & ~n_7529;
assign n_7531 = ~n_7526 & ~n_7530;
assign n_7532 = ~n_6146 & ~n_7531;
assign n_7533 =  x_3182 &  n_6146;
assign n_7534 = ~n_7532 & ~n_7533;
assign n_7535 =  x_3182 & ~n_7534;
assign n_7536 = ~x_3182 &  n_7534;
assign n_7537 = ~n_7535 & ~n_7536;
assign n_7538 = ~x_230 & ~x_1097;
assign n_7539 = ~x_1097 &  n_1126;
assign n_7540 = ~x_2022 &  n_447;
assign n_7541 = ~x_2028 &  n_441;
assign n_7542 = ~n_7540 & ~n_7541;
assign n_7543 = ~x_2026 &  n_444;
assign n_7544 = ~x_2024 &  n_449;
assign n_7545 = ~n_7543 & ~n_7544;
assign n_7546 =  n_7542 &  n_7545;
assign n_7547 = ~x_2023 &  n_463;
assign n_7548 = ~x_2025 &  n_466;
assign n_7549 = ~n_7547 & ~n_7548;
assign n_7550 = ~x_2027 &  n_468;
assign n_7551 = ~x_2029 &  n_460;
assign n_7552 = ~n_7550 & ~n_7551;
assign n_7553 =  n_7549 &  n_7552;
assign n_7554 =  n_7546 &  n_7553;
assign n_7555 =  x_231 &  n_7554;
assign n_7556 = ~n_7539 & ~n_7555;
assign n_7557 = ~x_1470 & ~n_7556;
assign n_7558 = ~n_7538 & ~n_7557;
assign n_7559 =  n_1713 & ~n_7558;
assign n_7560 =  x_1159 & ~n_436;
assign n_7561 =  n_436 &  n_7554;
assign n_7562 = ~n_7560 & ~n_7561;
assign n_7563 =  n_1321 & ~n_7562;
assign n_7564 = ~n_7559 & ~n_7563;
assign n_7565 = ~n_6146 & ~n_7564;
assign n_7566 =  x_3181 &  n_6146;
assign n_7567 = ~n_7565 & ~n_7566;
assign n_7568 =  x_3181 & ~n_7567;
assign n_7569 = ~x_3181 &  n_7567;
assign n_7570 = ~n_7568 & ~n_7569;
assign n_7571 = ~x_230 & ~x_1096;
assign n_7572 = ~x_1096 &  n_1126;
assign n_7573 = ~x_2020 &  n_441;
assign n_7574 = ~x_2016 &  n_449;
assign n_7575 = ~n_7573 & ~n_7574;
assign n_7576 = ~x_2018 &  n_444;
assign n_7577 = ~x_2014 &  n_447;
assign n_7578 = ~n_7576 & ~n_7577;
assign n_7579 =  n_7575 &  n_7578;
assign n_7580 = ~x_2019 &  n_468;
assign n_7581 = ~x_2021 &  n_460;
assign n_7582 = ~n_7580 & ~n_7581;
assign n_7583 = ~x_2015 &  n_463;
assign n_7584 = ~x_2017 &  n_466;
assign n_7585 = ~n_7583 & ~n_7584;
assign n_7586 =  n_7582 &  n_7585;
assign n_7587 =  n_7579 &  n_7586;
assign n_7588 =  x_231 &  n_7587;
assign n_7589 = ~n_7572 & ~n_7588;
assign n_7590 = ~x_1470 & ~n_7589;
assign n_7591 = ~n_7571 & ~n_7590;
assign n_7592 =  n_1713 & ~n_7591;
assign n_7593 =  x_1158 & ~n_436;
assign n_7594 =  n_436 &  n_7587;
assign n_7595 = ~n_7593 & ~n_7594;
assign n_7596 =  n_1321 & ~n_7595;
assign n_7597 = ~n_7592 & ~n_7596;
assign n_7598 = ~n_6146 & ~n_7597;
assign n_7599 =  x_3180 &  n_6146;
assign n_7600 = ~n_7598 & ~n_7599;
assign n_7601 =  x_3180 & ~n_7600;
assign n_7602 = ~x_3180 &  n_7600;
assign n_7603 = ~n_7601 & ~n_7602;
assign n_7604 = ~x_230 & ~x_1095;
assign n_7605 = ~x_1095 &  n_1126;
assign n_7606 = ~x_2010 &  n_444;
assign n_7607 = ~x_2008 &  n_449;
assign n_7608 = ~n_7606 & ~n_7607;
assign n_7609 = ~x_2012 &  n_441;
assign n_7610 = ~x_2006 &  n_447;
assign n_7611 = ~n_7609 & ~n_7610;
assign n_7612 =  n_7608 &  n_7611;
assign n_7613 = ~x_2011 &  n_468;
assign n_7614 = ~x_2009 &  n_466;
assign n_7615 = ~n_7613 & ~n_7614;
assign n_7616 = ~x_2007 &  n_463;
assign n_7617 = ~x_2013 &  n_460;
assign n_7618 = ~n_7616 & ~n_7617;
assign n_7619 =  n_7615 &  n_7618;
assign n_7620 =  n_7612 &  n_7619;
assign n_7621 =  x_231 &  n_7620;
assign n_7622 = ~n_7605 & ~n_7621;
assign n_7623 = ~x_1470 & ~n_7622;
assign n_7624 = ~n_7604 & ~n_7623;
assign n_7625 =  n_1713 & ~n_7624;
assign n_7626 =  x_1157 & ~n_436;
assign n_7627 =  n_436 &  n_7620;
assign n_7628 = ~n_7626 & ~n_7627;
assign n_7629 =  n_1321 & ~n_7628;
assign n_7630 = ~n_7625 & ~n_7629;
assign n_7631 = ~n_6146 & ~n_7630;
assign n_7632 =  x_3179 &  n_6146;
assign n_7633 = ~n_7631 & ~n_7632;
assign n_7634 =  x_3179 & ~n_7633;
assign n_7635 = ~x_3179 &  n_7633;
assign n_7636 = ~n_7634 & ~n_7635;
assign n_7637 = ~x_230 & ~x_1094;
assign n_7638 = ~x_1094 &  n_1126;
assign n_7639 = ~x_2002 &  n_444;
assign n_7640 = ~x_2004 &  n_441;
assign n_7641 = ~n_7639 & ~n_7640;
assign n_7642 = ~x_2000 &  n_449;
assign n_7643 = ~x_1998 &  n_447;
assign n_7644 = ~n_7642 & ~n_7643;
assign n_7645 =  n_7641 &  n_7644;
assign n_7646 = ~x_1999 &  n_463;
assign n_7647 = ~x_2003 &  n_468;
assign n_7648 = ~n_7646 & ~n_7647;
assign n_7649 = ~x_2005 &  n_460;
assign n_7650 = ~x_2001 &  n_466;
assign n_7651 = ~n_7649 & ~n_7650;
assign n_7652 =  n_7648 &  n_7651;
assign n_7653 =  n_7645 &  n_7652;
assign n_7654 =  x_231 &  n_7653;
assign n_7655 = ~n_7638 & ~n_7654;
assign n_7656 = ~x_1470 & ~n_7655;
assign n_7657 = ~n_7637 & ~n_7656;
assign n_7658 =  n_1713 & ~n_7657;
assign n_7659 =  x_1156 & ~n_436;
assign n_7660 =  n_436 &  n_7653;
assign n_7661 = ~n_7659 & ~n_7660;
assign n_7662 =  n_1321 & ~n_7661;
assign n_7663 = ~n_7658 & ~n_7662;
assign n_7664 = ~n_6146 & ~n_7663;
assign n_7665 =  x_3178 &  n_6146;
assign n_7666 = ~n_7664 & ~n_7665;
assign n_7667 =  x_3178 & ~n_7666;
assign n_7668 = ~x_3178 &  n_7666;
assign n_7669 = ~n_7667 & ~n_7668;
assign n_7670 = ~x_230 & ~x_1093;
assign n_7671 = ~x_1093 &  n_1126;
assign n_7672 = ~x_1992 &  n_449;
assign n_7673 = ~x_1996 &  n_441;
assign n_7674 = ~n_7672 & ~n_7673;
assign n_7675 = ~x_1990 &  n_447;
assign n_7676 = ~x_1994 &  n_444;
assign n_7677 = ~n_7675 & ~n_7676;
assign n_7678 =  n_7674 &  n_7677;
assign n_7679 = ~x_1991 &  n_463;
assign n_7680 = ~x_1993 &  n_466;
assign n_7681 = ~n_7679 & ~n_7680;
assign n_7682 = ~x_1995 &  n_468;
assign n_7683 = ~x_1997 &  n_460;
assign n_7684 = ~n_7682 & ~n_7683;
assign n_7685 =  n_7681 &  n_7684;
assign n_7686 =  n_7678 &  n_7685;
assign n_7687 =  x_231 &  n_7686;
assign n_7688 = ~n_7671 & ~n_7687;
assign n_7689 = ~x_1470 & ~n_7688;
assign n_7690 = ~n_7670 & ~n_7689;
assign n_7691 =  n_1713 & ~n_7690;
assign n_7692 =  x_1155 & ~n_436;
assign n_7693 =  n_436 &  n_7686;
assign n_7694 = ~n_7692 & ~n_7693;
assign n_7695 =  n_1321 & ~n_7694;
assign n_7696 = ~n_7691 & ~n_7695;
assign n_7697 = ~n_6146 & ~n_7696;
assign n_7698 =  x_3177 &  n_6146;
assign n_7699 = ~n_7697 & ~n_7698;
assign n_7700 =  x_3177 & ~n_7699;
assign n_7701 = ~x_3177 &  n_7699;
assign n_7702 = ~n_7700 & ~n_7701;
assign n_7703 =  x_1154 & ~n_436;
assign n_7704 = ~x_1982 &  n_447;
assign n_7705 = ~x_1988 &  n_441;
assign n_7706 = ~n_7704 & ~n_7705;
assign n_7707 = ~x_1984 &  n_449;
assign n_7708 = ~x_1986 &  n_444;
assign n_7709 = ~n_7707 & ~n_7708;
assign n_7710 =  n_7706 &  n_7709;
assign n_7711 = ~x_1985 &  n_466;
assign n_7712 = ~x_1983 &  n_463;
assign n_7713 = ~n_7711 & ~n_7712;
assign n_7714 = ~x_1989 &  n_460;
assign n_7715 = ~x_1987 &  n_468;
assign n_7716 = ~n_7714 & ~n_7715;
assign n_7717 =  n_7713 &  n_7716;
assign n_7718 =  n_7710 &  n_7717;
assign n_7719 =  n_436 &  n_7718;
assign n_7720 = ~n_7703 & ~n_7719;
assign n_7721 =  n_1321 & ~n_7720;
assign n_7722 = ~x_230 & ~x_1092;
assign n_7723 = ~x_1092 &  n_1126;
assign n_7724 =  x_231 &  n_7718;
assign n_7725 = ~n_7723 & ~n_7724;
assign n_7726 = ~x_1470 & ~n_7725;
assign n_7727 = ~n_7722 & ~n_7726;
assign n_7728 =  n_1713 & ~n_7727;
assign n_7729 = ~n_7721 & ~n_7728;
assign n_7730 =  x_3176 &  n_7729;
assign n_7731 = ~x_3176 & ~n_7729;
assign n_7732 = ~n_7730 & ~n_7731;
assign n_7733 =  n_6146 & ~n_4197;
assign n_7734 =  x_3175 & ~n_7733;
assign n_7735 = ~x_3175 &  n_7733;
assign n_7736 = ~n_7734 & ~n_7735;
assign n_7737 = ~x_230 & ~x_1091;
assign n_7738 = ~x_1091 &  n_1126;
assign n_7739 = ~x_1974 &  n_447;
assign n_7740 = ~x_1980 &  n_441;
assign n_7741 = ~n_7739 & ~n_7740;
assign n_7742 = ~x_1976 &  n_449;
assign n_7743 = ~x_1978 &  n_444;
assign n_7744 = ~n_7742 & ~n_7743;
assign n_7745 =  n_7741 &  n_7744;
assign n_7746 = ~x_1977 &  n_466;
assign n_7747 = ~x_1981 &  n_460;
assign n_7748 = ~n_7746 & ~n_7747;
assign n_7749 = ~x_1979 &  n_468;
assign n_7750 = ~x_1975 &  n_463;
assign n_7751 = ~n_7749 & ~n_7750;
assign n_7752 =  n_7748 &  n_7751;
assign n_7753 =  n_7745 &  n_7752;
assign n_7754 =  x_231 &  n_7753;
assign n_7755 = ~n_7738 & ~n_7754;
assign n_7756 = ~x_1470 & ~n_7755;
assign n_7757 = ~n_7737 & ~n_7756;
assign n_7758 =  n_1713 & ~n_7757;
assign n_7759 =  x_1153 & ~n_436;
assign n_7760 =  n_436 &  n_7753;
assign n_7761 = ~n_7759 & ~n_7760;
assign n_7762 =  n_1321 & ~n_7761;
assign n_7763 = ~n_7758 & ~n_7762;
assign n_7764 = ~n_6146 & ~n_7763;
assign n_7765 =  x_3174 &  n_6146;
assign n_7766 = ~n_7764 & ~n_7765;
assign n_7767 =  x_3174 & ~n_7766;
assign n_7768 = ~x_3174 &  n_7766;
assign n_7769 = ~n_7767 & ~n_7768;
assign n_7770 = ~x_230 & ~x_1090;
assign n_7771 = ~x_1090 &  n_1126;
assign n_7772 = ~x_1966 &  n_447;
assign n_7773 = ~x_1972 &  n_441;
assign n_7774 = ~n_7772 & ~n_7773;
assign n_7775 = ~x_1968 &  n_449;
assign n_7776 = ~x_1970 &  n_444;
assign n_7777 = ~n_7775 & ~n_7776;
assign n_7778 =  n_7774 &  n_7777;
assign n_7779 = ~x_1967 &  n_463;
assign n_7780 = ~x_1973 &  n_460;
assign n_7781 = ~n_7779 & ~n_7780;
assign n_7782 = ~x_1971 &  n_468;
assign n_7783 = ~x_1969 &  n_466;
assign n_7784 = ~n_7782 & ~n_7783;
assign n_7785 =  n_7781 &  n_7784;
assign n_7786 =  n_7778 &  n_7785;
assign n_7787 =  x_231 &  n_7786;
assign n_7788 = ~n_7771 & ~n_7787;
assign n_7789 = ~x_1470 & ~n_7788;
assign n_7790 = ~n_7770 & ~n_7789;
assign n_7791 =  n_1713 & ~n_7790;
assign n_7792 =  x_1152 & ~n_436;
assign n_7793 =  n_436 &  n_7786;
assign n_7794 = ~n_7792 & ~n_7793;
assign n_7795 =  n_1321 & ~n_7794;
assign n_7796 = ~n_7791 & ~n_7795;
assign n_7797 = ~n_6146 & ~n_7796;
assign n_7798 =  x_3173 &  n_6146;
assign n_7799 = ~n_7797 & ~n_7798;
assign n_7800 =  x_3173 & ~n_7799;
assign n_7801 = ~x_3173 &  n_7799;
assign n_7802 = ~n_7800 & ~n_7801;
assign n_7803 = ~x_230 & ~x_1089;
assign n_7804 = ~x_1089 &  n_1126;
assign n_7805 = ~x_1958 &  n_447;
assign n_7806 = ~x_1964 &  n_441;
assign n_7807 = ~n_7805 & ~n_7806;
assign n_7808 = ~x_1962 &  n_444;
assign n_7809 = ~x_1960 &  n_449;
assign n_7810 = ~n_7808 & ~n_7809;
assign n_7811 =  n_7807 &  n_7810;
assign n_7812 = ~x_1965 &  n_460;
assign n_7813 = ~x_1961 &  n_466;
assign n_7814 = ~n_7812 & ~n_7813;
assign n_7815 = ~x_1963 &  n_468;
assign n_7816 = ~x_1959 &  n_463;
assign n_7817 = ~n_7815 & ~n_7816;
assign n_7818 =  n_7814 &  n_7817;
assign n_7819 =  n_7811 &  n_7818;
assign n_7820 =  x_231 &  n_7819;
assign n_7821 = ~n_7804 & ~n_7820;
assign n_7822 = ~x_1470 & ~n_7821;
assign n_7823 = ~n_7803 & ~n_7822;
assign n_7824 =  n_1713 & ~n_7823;
assign n_7825 =  x_1151 & ~n_436;
assign n_7826 =  n_436 &  n_7819;
assign n_7827 = ~n_7825 & ~n_7826;
assign n_7828 =  n_1321 & ~n_7827;
assign n_7829 = ~n_7824 & ~n_7828;
assign n_7830 = ~n_6146 & ~n_7829;
assign n_7831 =  x_3172 &  n_6146;
assign n_7832 = ~n_7830 & ~n_7831;
assign n_7833 =  x_3172 & ~n_7832;
assign n_7834 = ~x_3172 &  n_7832;
assign n_7835 = ~n_7833 & ~n_7834;
assign n_7836 = ~x_230 & ~x_1088;
assign n_7837 = ~x_1088 &  n_1126;
assign n_7838 = ~x_1950 &  n_447;
assign n_7839 = ~x_1952 &  n_449;
assign n_7840 = ~n_7838 & ~n_7839;
assign n_7841 = ~x_1956 &  n_441;
assign n_7842 = ~x_1954 &  n_444;
assign n_7843 = ~n_7841 & ~n_7842;
assign n_7844 =  n_7840 &  n_7843;
assign n_7845 = ~x_1953 &  n_466;
assign n_7846 = ~x_1951 &  n_463;
assign n_7847 = ~n_7845 & ~n_7846;
assign n_7848 = ~x_1957 &  n_460;
assign n_7849 = ~x_1955 &  n_468;
assign n_7850 = ~n_7848 & ~n_7849;
assign n_7851 =  n_7847 &  n_7850;
assign n_7852 =  n_7844 &  n_7851;
assign n_7853 =  x_231 &  n_7852;
assign n_7854 = ~n_7837 & ~n_7853;
assign n_7855 = ~x_1470 & ~n_7854;
assign n_7856 = ~n_7836 & ~n_7855;
assign n_7857 =  n_1713 & ~n_7856;
assign n_7858 =  x_1150 & ~n_436;
assign n_7859 =  n_436 &  n_7852;
assign n_7860 = ~n_7858 & ~n_7859;
assign n_7861 =  n_1321 & ~n_7860;
assign n_7862 = ~n_7857 & ~n_7861;
assign n_7863 = ~n_6146 & ~n_7862;
assign n_7864 =  x_3171 &  n_6146;
assign n_7865 = ~n_7863 & ~n_7864;
assign n_7866 =  x_3171 & ~n_7865;
assign n_7867 = ~x_3171 &  n_7865;
assign n_7868 = ~n_7866 & ~n_7867;
assign n_7869 = ~x_230 & ~x_1087;
assign n_7870 = ~x_1087 &  n_1126;
assign n_7871 = ~x_1942 &  n_447;
assign n_7872 = ~x_1946 &  n_444;
assign n_7873 = ~n_7871 & ~n_7872;
assign n_7874 = ~x_1944 &  n_449;
assign n_7875 = ~x_1948 &  n_441;
assign n_7876 = ~n_7874 & ~n_7875;
assign n_7877 =  n_7873 &  n_7876;
assign n_7878 = ~x_1945 &  n_466;
assign n_7879 = ~x_1947 &  n_468;
assign n_7880 = ~n_7878 & ~n_7879;
assign n_7881 = ~x_1949 &  n_460;
assign n_7882 = ~x_1943 &  n_463;
assign n_7883 = ~n_7881 & ~n_7882;
assign n_7884 =  n_7880 &  n_7883;
assign n_7885 =  n_7877 &  n_7884;
assign n_7886 =  x_231 &  n_7885;
assign n_7887 = ~n_7870 & ~n_7886;
assign n_7888 = ~x_1470 & ~n_7887;
assign n_7889 = ~n_7869 & ~n_7888;
assign n_7890 =  n_1713 & ~n_7889;
assign n_7891 =  x_1149 & ~n_436;
assign n_7892 =  n_436 &  n_7885;
assign n_7893 = ~n_7891 & ~n_7892;
assign n_7894 =  n_1321 & ~n_7893;
assign n_7895 = ~n_7890 & ~n_7894;
assign n_7896 = ~n_6146 & ~n_7895;
assign n_7897 =  x_3170 &  n_6146;
assign n_7898 = ~n_7896 & ~n_7897;
assign n_7899 =  x_3170 & ~n_7898;
assign n_7900 = ~x_3170 &  n_7898;
assign n_7901 = ~n_7899 & ~n_7900;
assign n_7902 = ~x_230 & ~x_1086;
assign n_7903 = ~x_1086 &  n_1126;
assign n_7904 = ~x_1940 &  n_441;
assign n_7905 = ~x_1936 &  n_449;
assign n_7906 = ~n_7904 & ~n_7905;
assign n_7907 = ~x_1938 &  n_444;
assign n_7908 = ~x_1934 &  n_447;
assign n_7909 = ~n_7907 & ~n_7908;
assign n_7910 =  n_7906 &  n_7909;
assign n_7911 = ~x_1935 &  n_463;
assign n_7912 = ~x_1939 &  n_468;
assign n_7913 = ~n_7911 & ~n_7912;
assign n_7914 = ~x_1937 &  n_466;
assign n_7915 = ~x_1941 &  n_460;
assign n_7916 = ~n_7914 & ~n_7915;
assign n_7917 =  n_7913 &  n_7916;
assign n_7918 =  n_7910 &  n_7917;
assign n_7919 =  x_231 &  n_7918;
assign n_7920 = ~n_7903 & ~n_7919;
assign n_7921 = ~x_1470 & ~n_7920;
assign n_7922 = ~n_7902 & ~n_7921;
assign n_7923 =  n_1713 & ~n_7922;
assign n_7924 =  x_1148 & ~n_436;
assign n_7925 =  n_436 &  n_7918;
assign n_7926 = ~n_7924 & ~n_7925;
assign n_7927 =  n_1321 & ~n_7926;
assign n_7928 = ~n_7923 & ~n_7927;
assign n_7929 = ~n_6146 & ~n_7928;
assign n_7930 =  x_3169 &  n_6146;
assign n_7931 = ~n_7929 & ~n_7930;
assign n_7932 =  x_3169 & ~n_7931;
assign n_7933 = ~x_3169 &  n_7931;
assign n_7934 = ~n_7932 & ~n_7933;
assign n_7935 = ~x_230 & ~x_1085;
assign n_7936 = ~x_1085 &  n_1126;
assign n_7937 = ~x_1928 &  n_449;
assign n_7938 = ~x_1932 &  n_441;
assign n_7939 = ~n_7937 & ~n_7938;
assign n_7940 = ~x_1926 &  n_447;
assign n_7941 = ~x_1930 &  n_444;
assign n_7942 = ~n_7940 & ~n_7941;
assign n_7943 =  n_7939 &  n_7942;
assign n_7944 = ~x_1927 &  n_463;
assign n_7945 = ~x_1929 &  n_466;
assign n_7946 = ~n_7944 & ~n_7945;
assign n_7947 = ~x_1931 &  n_468;
assign n_7948 = ~x_1933 &  n_460;
assign n_7949 = ~n_7947 & ~n_7948;
assign n_7950 =  n_7946 &  n_7949;
assign n_7951 =  n_7943 &  n_7950;
assign n_7952 =  x_231 &  n_7951;
assign n_7953 = ~n_7936 & ~n_7952;
assign n_7954 = ~x_1470 & ~n_7953;
assign n_7955 = ~n_7935 & ~n_7954;
assign n_7956 =  n_1713 & ~n_7955;
assign n_7957 =  x_1147 & ~n_436;
assign n_7958 =  n_436 &  n_7951;
assign n_7959 = ~n_7957 & ~n_7958;
assign n_7960 =  n_1321 & ~n_7959;
assign n_7961 = ~n_7956 & ~n_7960;
assign n_7962 = ~n_6146 & ~n_7961;
assign n_7963 =  x_3168 &  n_6146;
assign n_7964 = ~n_7962 & ~n_7963;
assign n_7965 =  x_3168 & ~n_7964;
assign n_7966 = ~x_3168 &  n_7964;
assign n_7967 = ~n_7965 & ~n_7966;
assign n_7968 = ~x_230 & ~x_1084;
assign n_7969 = ~x_1084 &  n_1126;
assign n_7970 = ~x_1924 &  n_441;
assign n_7971 = ~x_1920 &  n_449;
assign n_7972 = ~n_7970 & ~n_7971;
assign n_7973 = ~x_1922 &  n_444;
assign n_7974 = ~x_1918 &  n_447;
assign n_7975 = ~n_7973 & ~n_7974;
assign n_7976 =  n_7972 &  n_7975;
assign n_7977 = ~x_1919 &  n_463;
assign n_7978 = ~x_1923 &  n_468;
assign n_7979 = ~n_7977 & ~n_7978;
assign n_7980 = ~x_1921 &  n_466;
assign n_7981 = ~x_1925 &  n_460;
assign n_7982 = ~n_7980 & ~n_7981;
assign n_7983 =  n_7979 &  n_7982;
assign n_7984 =  n_7976 &  n_7983;
assign n_7985 =  x_231 &  n_7984;
assign n_7986 = ~n_7969 & ~n_7985;
assign n_7987 = ~x_1470 & ~n_7986;
assign n_7988 = ~n_7968 & ~n_7987;
assign n_7989 =  n_1713 & ~n_7988;
assign n_7990 =  x_1146 & ~n_436;
assign n_7991 =  n_436 &  n_7984;
assign n_7992 = ~n_7990 & ~n_7991;
assign n_7993 =  n_1321 & ~n_7992;
assign n_7994 = ~n_7989 & ~n_7993;
assign n_7995 =  x_3167 &  n_7994;
assign n_7996 = ~x_3167 & ~n_7994;
assign n_7997 = ~n_7995 & ~n_7996;
assign n_7998 =  n_6146 & ~n_4189;
assign n_7999 =  x_3166 & ~n_7998;
assign n_8000 = ~x_3166 &  n_7998;
assign n_8001 = ~n_7999 & ~n_8000;
assign n_8002 = ~x_230 & ~x_1075;
assign n_8003 = ~x_1075 &  n_1126;
assign n_8004 = ~x_1915 &  n_441;
assign n_8005 = ~x_1913 &  n_444;
assign n_8006 = ~n_8004 & ~n_8005;
assign n_8007 = ~x_1911 &  n_449;
assign n_8008 = ~x_1909 &  n_447;
assign n_8009 = ~n_8007 & ~n_8008;
assign n_8010 =  n_8006 &  n_8009;
assign n_8011 = ~x_1914 &  n_468;
assign n_8012 = ~x_1916 &  n_460;
assign n_8013 = ~n_8011 & ~n_8012;
assign n_8014 = ~x_1910 &  n_463;
assign n_8015 = ~x_1912 &  n_466;
assign n_8016 = ~n_8014 & ~n_8015;
assign n_8017 =  n_8013 &  n_8016;
assign n_8018 =  n_8010 &  n_8017;
assign n_8019 =  x_231 &  n_8018;
assign n_8020 = ~n_8003 & ~n_8019;
assign n_8021 = ~x_1470 & ~n_8020;
assign n_8022 = ~n_8002 & ~n_8021;
assign n_8023 =  n_1713 & ~n_8022;
assign n_8024 =  x_1145 & ~n_436;
assign n_8025 =  n_436 &  n_8018;
assign n_8026 = ~n_8024 & ~n_8025;
assign n_8027 =  n_1321 & ~n_8026;
assign n_8028 = ~n_8023 & ~n_8027;
assign n_8029 = ~n_6146 & ~n_8028;
assign n_8030 =  x_3165 &  n_6146;
assign n_8031 = ~n_8029 & ~n_8030;
assign n_8032 =  x_3165 & ~n_8031;
assign n_8033 = ~x_3165 &  n_8031;
assign n_8034 = ~n_8032 & ~n_8033;
assign n_8035 = ~x_230 & ~x_1066;
assign n_8036 = ~x_1066 &  n_1126;
assign n_8037 = ~x_1900 &  n_447;
assign n_8038 = ~x_1902 &  n_449;
assign n_8039 = ~n_8037 & ~n_8038;
assign n_8040 = ~x_1906 &  n_441;
assign n_8041 = ~x_1904 &  n_444;
assign n_8042 = ~n_8040 & ~n_8041;
assign n_8043 =  n_8039 &  n_8042;
assign n_8044 = ~x_1901 &  n_463;
assign n_8045 = ~x_1903 &  n_466;
assign n_8046 = ~n_8044 & ~n_8045;
assign n_8047 = ~x_1905 &  n_468;
assign n_8048 = ~x_1907 &  n_460;
assign n_8049 = ~n_8047 & ~n_8048;
assign n_8050 =  n_8046 &  n_8049;
assign n_8051 =  n_8043 &  n_8050;
assign n_8052 =  x_231 &  n_8051;
assign n_8053 = ~n_8036 & ~n_8052;
assign n_8054 = ~x_1470 & ~n_8053;
assign n_8055 = ~n_8035 & ~n_8054;
assign n_8056 =  n_1713 & ~n_8055;
assign n_8057 =  x_1144 & ~n_436;
assign n_8058 =  n_436 &  n_8051;
assign n_8059 = ~n_8057 & ~n_8058;
assign n_8060 =  n_1321 & ~n_8059;
assign n_8061 = ~n_8056 & ~n_8060;
assign n_8062 = ~n_6146 & ~n_8061;
assign n_8063 =  x_3164 &  n_6146;
assign n_8064 = ~n_8062 & ~n_8063;
assign n_8065 =  x_3164 & ~n_8064;
assign n_8066 = ~x_3164 &  n_8064;
assign n_8067 = ~n_8065 & ~n_8066;
assign n_8068 = ~x_230 & ~x_1057;
assign n_8069 = ~x_1057 &  n_1126;
assign n_8070 = ~x_1891 &  n_447;
assign n_8071 = ~x_1897 &  n_441;
assign n_8072 = ~n_8070 & ~n_8071;
assign n_8073 = ~x_1893 &  n_449;
assign n_8074 = ~x_1895 &  n_444;
assign n_8075 = ~n_8073 & ~n_8074;
assign n_8076 =  n_8072 &  n_8075;
assign n_8077 = ~x_1892 &  n_463;
assign n_8078 = ~x_1898 &  n_460;
assign n_8079 = ~n_8077 & ~n_8078;
assign n_8080 = ~x_1896 &  n_468;
assign n_8081 = ~x_1894 &  n_466;
assign n_8082 = ~n_8080 & ~n_8081;
assign n_8083 =  n_8079 &  n_8082;
assign n_8084 =  n_8076 &  n_8083;
assign n_8085 =  x_231 &  n_8084;
assign n_8086 = ~n_8069 & ~n_8085;
assign n_8087 = ~x_1470 & ~n_8086;
assign n_8088 = ~n_8068 & ~n_8087;
assign n_8089 =  n_1713 & ~n_8088;
assign n_8090 =  x_1143 & ~n_436;
assign n_8091 =  n_436 &  n_8084;
assign n_8092 = ~n_8090 & ~n_8091;
assign n_8093 =  n_1321 & ~n_8092;
assign n_8094 = ~n_8089 & ~n_8093;
assign n_8095 = ~n_6146 & ~n_8094;
assign n_8096 =  x_3163 &  n_6146;
assign n_8097 = ~n_8095 & ~n_8096;
assign n_8098 =  x_3163 & ~n_8097;
assign n_8099 = ~x_3163 &  n_8097;
assign n_8100 = ~n_8098 & ~n_8099;
assign n_8101 = ~x_230 & ~x_1048;
assign n_8102 = ~x_1048 &  n_1126;
assign n_8103 = ~x_1888 &  n_441;
assign n_8104 = ~x_1882 &  n_447;
assign n_8105 = ~n_8103 & ~n_8104;
assign n_8106 = ~x_1884 &  n_449;
assign n_8107 = ~x_1886 &  n_444;
assign n_8108 = ~n_8106 & ~n_8107;
assign n_8109 =  n_8105 &  n_8108;
assign n_8110 = ~x_1887 &  n_468;
assign n_8111 = ~x_1889 &  n_460;
assign n_8112 = ~n_8110 & ~n_8111;
assign n_8113 = ~x_1883 &  n_463;
assign n_8114 = ~x_1885 &  n_466;
assign n_8115 = ~n_8113 & ~n_8114;
assign n_8116 =  n_8112 &  n_8115;
assign n_8117 =  n_8109 &  n_8116;
assign n_8118 =  x_231 &  n_8117;
assign n_8119 = ~n_8102 & ~n_8118;
assign n_8120 = ~x_1470 & ~n_8119;
assign n_8121 = ~n_8101 & ~n_8120;
assign n_8122 =  n_1713 & ~n_8121;
assign n_8123 =  x_1142 & ~n_436;
assign n_8124 =  n_436 &  n_8117;
assign n_8125 = ~n_8123 & ~n_8124;
assign n_8126 =  n_1321 & ~n_8125;
assign n_8127 = ~n_8122 & ~n_8126;
assign n_8128 = ~n_6146 & ~n_8127;
assign n_8129 =  x_3162 &  n_6146;
assign n_8130 = ~n_8128 & ~n_8129;
assign n_8131 =  x_3162 & ~n_8130;
assign n_8132 = ~x_3162 &  n_8130;
assign n_8133 = ~n_8131 & ~n_8132;
assign n_8134 = ~x_230 & ~x_1039;
assign n_8135 = ~x_1039 &  n_1126;
assign n_8136 = ~x_1877 &  n_444;
assign n_8137 = ~x_1879 &  n_441;
assign n_8138 = ~n_8136 & ~n_8137;
assign n_8139 = ~x_1873 &  n_447;
assign n_8140 = ~x_1875 &  n_449;
assign n_8141 = ~n_8139 & ~n_8140;
assign n_8142 =  n_8138 &  n_8141;
assign n_8143 = ~x_1874 &  n_463;
assign n_8144 = ~x_1876 &  n_466;
assign n_8145 = ~n_8143 & ~n_8144;
assign n_8146 = ~x_1880 &  n_460;
assign n_8147 = ~x_1878 &  n_468;
assign n_8148 = ~n_8146 & ~n_8147;
assign n_8149 =  n_8145 &  n_8148;
assign n_8150 =  n_8142 &  n_8149;
assign n_8151 =  x_231 &  n_8150;
assign n_8152 = ~n_8135 & ~n_8151;
assign n_8153 = ~x_1470 & ~n_8152;
assign n_8154 = ~n_8134 & ~n_8153;
assign n_8155 =  n_1713 & ~n_8154;
assign n_8156 =  x_1141 & ~n_436;
assign n_8157 =  n_436 &  n_8150;
assign n_8158 = ~n_8156 & ~n_8157;
assign n_8159 =  n_1321 & ~n_8158;
assign n_8160 = ~n_8155 & ~n_8159;
assign n_8161 = ~n_6146 & ~n_8160;
assign n_8162 =  x_3161 &  n_6146;
assign n_8163 = ~n_8161 & ~n_8162;
assign n_8164 =  x_3161 & ~n_8163;
assign n_8165 = ~x_3161 &  n_8163;
assign n_8166 = ~n_8164 & ~n_8165;
assign n_8167 = ~x_230 & ~x_1030;
assign n_8168 = ~x_1030 &  n_1126;
assign n_8169 = ~x_1864 &  n_447;
assign n_8170 = ~x_1866 &  n_449;
assign n_8171 = ~n_8169 & ~n_8170;
assign n_8172 = ~x_1870 &  n_441;
assign n_8173 = ~x_1868 &  n_444;
assign n_8174 = ~n_8172 & ~n_8173;
assign n_8175 =  n_8171 &  n_8174;
assign n_8176 = ~x_1867 &  n_466;
assign n_8177 = ~x_1869 &  n_468;
assign n_8178 = ~n_8176 & ~n_8177;
assign n_8179 = ~x_1871 &  n_460;
assign n_8180 = ~x_1865 &  n_463;
assign n_8181 = ~n_8179 & ~n_8180;
assign n_8182 =  n_8178 &  n_8181;
assign n_8183 =  n_8175 &  n_8182;
assign n_8184 =  x_231 &  n_8183;
assign n_8185 = ~n_8168 & ~n_8184;
assign n_8186 = ~x_1470 & ~n_8185;
assign n_8187 = ~n_8167 & ~n_8186;
assign n_8188 =  n_1713 & ~n_8187;
assign n_8189 =  x_1140 & ~n_436;
assign n_8190 =  n_436 &  n_8183;
assign n_8191 = ~n_8189 & ~n_8190;
assign n_8192 =  n_1321 & ~n_8191;
assign n_8193 = ~n_8188 & ~n_8192;
assign n_8194 = ~n_6146 & ~n_8193;
assign n_8195 =  x_3160 &  n_6146;
assign n_8196 = ~n_8194 & ~n_8195;
assign n_8197 =  x_3160 & ~n_8196;
assign n_8198 = ~x_3160 &  n_8196;
assign n_8199 = ~n_8197 & ~n_8198;
assign n_8200 =  x_3159 &  n_6146;
assign n_8201 = ~x_3159 & ~n_6146;
assign n_8202 = ~n_8200 & ~n_8201;
assign n_8203 =  x_3158 &  n_6143;
assign n_8204 = ~x_3158 & ~n_6143;
assign n_8205 = ~n_8203 & ~n_8204;
assign n_8206 = ~n_6005 & ~n_5940;
assign n_8207 =  x_3157 & ~n_8206;
assign n_8208 = ~x_3157 &  n_8206;
assign n_8209 = ~n_8207 & ~n_8208;
assign n_8210 =  n_3617 & ~n_3670;
assign n_8211 =  x_3156 &  n_8210;
assign n_8212 = ~x_3156 & ~n_8210;
assign n_8213 = ~n_8211 & ~n_8212;
assign n_8214 =  n_6067 &  n_3633;
assign n_8215 =  x_3155 &  n_8214;
assign n_8216 = ~x_3155 & ~n_8214;
assign n_8217 = ~n_8215 & ~n_8216;
assign n_8218 = ~x_3154 & ~n_3702;
assign n_8219 = ~n_3699 & ~n_8218;
assign n_8220 =  x_3154 &  n_8219;
assign n_8221 = ~x_3154 & ~n_8219;
assign n_8222 = ~n_8220 & ~n_8221;
assign n_8223 = ~n_3701 &  n_3699;
assign n_8224 = ~n_3706 & ~n_8223;
assign n_8225 =  x_3153 &  n_8224;
assign n_8226 = ~x_3153 & ~n_8224;
assign n_8227 = ~n_8225 & ~n_8226;
assign n_8228 =  x_3152 & ~n_4341;
assign n_8229 =  i_143 &  n_4341;
assign n_8230 = ~n_8228 & ~n_8229;
assign n_8231 =  x_3152 & ~n_8230;
assign n_8232 = ~x_3152 &  n_8230;
assign n_8233 = ~n_8231 & ~n_8232;
assign n_8234 =  x_3151 & ~n_4341;
assign n_8235 =  n_4323 &  n_4341;
assign n_8236 = ~n_8234 & ~n_8235;
assign n_8237 =  x_3151 & ~n_8236;
assign n_8238 = ~x_3151 &  n_8236;
assign n_8239 = ~n_8237 & ~n_8238;
assign n_8240 =  x_3150 & ~n_4341;
assign n_8241 =  i_145 &  n_4341;
assign n_8242 = ~n_8240 & ~n_8241;
assign n_8243 =  x_3150 & ~n_8242;
assign n_8244 = ~x_3150 &  n_8242;
assign n_8245 = ~n_8243 & ~n_8244;
assign n_8246 =  x_3149 & ~n_4341;
assign n_8247 =  n_4304 &  n_4341;
assign n_8248 = ~n_8246 & ~n_8247;
assign n_8249 =  x_3149 & ~n_8248;
assign n_8250 = ~x_3149 &  n_8248;
assign n_8251 = ~n_8249 & ~n_8250;
assign n_8252 =  x_3148 & ~n_4341;
assign n_8253 =  n_4317 &  n_4341;
assign n_8254 = ~n_8252 & ~n_8253;
assign n_8255 =  x_3148 & ~n_8254;
assign n_8256 = ~x_3148 &  n_8254;
assign n_8257 = ~n_8255 & ~n_8256;
assign n_8258 =  x_3147 & ~n_4341;
assign n_8259 =  n_4328 &  n_4341;
assign n_8260 = ~n_8258 & ~n_8259;
assign n_8261 =  x_3147 & ~n_8260;
assign n_8262 = ~x_3147 &  n_8260;
assign n_8263 = ~n_8261 & ~n_8262;
assign n_8264 =  x_3146 & ~n_4341;
assign n_8265 =  n_4315 &  n_4341;
assign n_8266 = ~n_8264 & ~n_8265;
assign n_8267 =  x_3146 & ~n_8266;
assign n_8268 = ~x_3146 &  n_8266;
assign n_8269 = ~n_8267 & ~n_8268;
assign n_8270 =  x_3145 & ~n_4341;
assign n_8271 =  n_4326 &  n_4341;
assign n_8272 = ~n_8270 & ~n_8271;
assign n_8273 =  x_3145 & ~n_8272;
assign n_8274 = ~x_3145 &  n_8272;
assign n_8275 = ~n_8273 & ~n_8274;
assign n_8276 =  x_3144 &  n_4303;
assign n_8277 = ~x_3144 & ~n_4303;
assign n_8278 = ~n_8276 & ~n_8277;
assign n_8279 =  x_3143 &  n_4349;
assign n_8280 =  n_4360 &  n_8279;
assign n_8281 = ~n_4362 & ~n_8280;
assign n_8282 =  x_3143 & ~n_8281;
assign n_8283 = ~x_3143 &  n_8281;
assign n_8284 = ~n_8282 & ~n_8283;
assign n_8285 = ~x_3141 &  n_4361;
assign n_8286 = ~x_3142 & ~n_8285;
assign n_8287 =  x_3142 & ~n_8286;
assign n_8288 = ~x_3142 &  n_8286;
assign n_8289 = ~n_8287 & ~n_8288;
assign n_8290 = ~x_3141 &  n_4349;
assign n_8291 = ~n_8290 &  n_4360;
assign n_8292 =  x_3141 &  n_8291;
assign n_8293 = ~x_3141 & ~n_8291;
assign n_8294 = ~n_8292 & ~n_8293;
assign n_8295 =  x_3140 &  n_4294;
assign n_8296 = ~x_3140 & ~n_4294;
assign n_8297 = ~n_8295 & ~n_8296;
assign n_8298 =  x_3139 & ~n_3763;
assign n_8299 = ~x_3139 &  n_3763;
assign n_8300 = ~n_8298 & ~n_8299;
assign n_8301 =  x_3138 & ~n_3766;
assign n_8302 = ~x_3138 &  n_3766;
assign n_8303 = ~n_8301 & ~n_8302;
assign n_8304 =  x_3137 & ~n_3771;
assign n_8305 = ~x_3137 &  n_3771;
assign n_8306 = ~n_8304 & ~n_8305;
assign n_8307 =  x_3136 & ~n_3776;
assign n_8308 = ~x_3136 &  n_3776;
assign n_8309 = ~n_8307 & ~n_8308;
assign n_8310 =  x_3135 & ~n_3781;
assign n_8311 = ~x_3135 &  n_3781;
assign n_8312 = ~n_8310 & ~n_8311;
assign n_8313 =  x_3134 & ~n_3786;
assign n_8314 = ~x_3134 &  n_3786;
assign n_8315 = ~n_8313 & ~n_8314;
assign n_8316 =  x_3133 & ~n_3791;
assign n_8317 = ~x_3133 &  n_3791;
assign n_8318 = ~n_8316 & ~n_8317;
assign n_8319 =  x_3132 & ~n_3796;
assign n_8320 = ~x_3132 &  n_3796;
assign n_8321 = ~n_8319 & ~n_8320;
assign n_8322 =  x_3131 & ~n_3801;
assign n_8323 = ~x_3131 &  n_3801;
assign n_8324 = ~n_8322 & ~n_8323;
assign n_8325 =  x_3130 & ~n_3806;
assign n_8326 = ~x_3130 &  n_3806;
assign n_8327 = ~n_8325 & ~n_8326;
assign n_8328 =  x_3129 & ~n_3811;
assign n_8329 = ~x_3129 &  n_3811;
assign n_8330 = ~n_8328 & ~n_8329;
assign n_8331 =  x_3128 & ~n_3816;
assign n_8332 = ~x_3128 &  n_3816;
assign n_8333 = ~n_8331 & ~n_8332;
assign n_8334 =  x_3127 & ~n_3821;
assign n_8335 = ~x_3127 &  n_3821;
assign n_8336 = ~n_8334 & ~n_8335;
assign n_8337 =  x_3126 & ~n_3826;
assign n_8338 = ~x_3126 &  n_3826;
assign n_8339 = ~n_8337 & ~n_8338;
assign n_8340 =  x_3125 & ~n_3831;
assign n_8341 = ~x_3125 &  n_3831;
assign n_8342 = ~n_8340 & ~n_8341;
assign n_8343 =  x_3124 & ~n_3836;
assign n_8344 = ~x_3124 &  n_3836;
assign n_8345 = ~n_8343 & ~n_8344;
assign n_8346 =  x_3123 & ~n_3841;
assign n_8347 = ~x_3123 &  n_3841;
assign n_8348 = ~n_8346 & ~n_8347;
assign n_8349 =  x_3122 & ~n_3846;
assign n_8350 = ~x_3122 &  n_3846;
assign n_8351 = ~n_8349 & ~n_8350;
assign n_8352 =  x_3121 & ~n_3851;
assign n_8353 = ~x_3121 &  n_3851;
assign n_8354 = ~n_8352 & ~n_8353;
assign n_8355 =  x_3120 & ~n_3856;
assign n_8356 = ~x_3120 &  n_3856;
assign n_8357 = ~n_8355 & ~n_8356;
assign n_8358 =  x_3119 & ~n_3861;
assign n_8359 = ~x_3119 &  n_3861;
assign n_8360 = ~n_8358 & ~n_8359;
assign n_8361 =  x_3118 & ~n_3866;
assign n_8362 = ~x_3118 &  n_3866;
assign n_8363 = ~n_8361 & ~n_8362;
assign n_8364 =  x_3117 & ~n_3871;
assign n_8365 = ~x_3117 &  n_3871;
assign n_8366 = ~n_8364 & ~n_8365;
assign n_8367 =  x_3116 & ~n_3876;
assign n_8368 = ~x_3116 &  n_3876;
assign n_8369 = ~n_8367 & ~n_8368;
assign n_8370 =  x_3115 & ~n_3881;
assign n_8371 = ~x_3115 &  n_3881;
assign n_8372 = ~n_8370 & ~n_8371;
assign n_8373 =  x_3114 & ~n_3886;
assign n_8374 = ~x_3114 &  n_3886;
assign n_8375 = ~n_8373 & ~n_8374;
assign n_8376 =  x_3113 & ~n_3891;
assign n_8377 = ~x_3113 &  n_3891;
assign n_8378 = ~n_8376 & ~n_8377;
assign n_8379 =  x_3112 & ~n_3896;
assign n_8380 = ~x_3112 &  n_3896;
assign n_8381 = ~n_8379 & ~n_8380;
assign n_8382 =  x_3111 & ~n_3901;
assign n_8383 = ~x_3111 &  n_3901;
assign n_8384 = ~n_8382 & ~n_8383;
assign n_8385 =  x_3110 & ~n_3906;
assign n_8386 = ~x_3110 &  n_3906;
assign n_8387 = ~n_8385 & ~n_8386;
assign n_8388 =  x_3109 & ~n_3911;
assign n_8389 = ~x_3109 &  n_3911;
assign n_8390 = ~n_8388 & ~n_8389;
assign n_8391 =  x_3108 & ~n_1325;
assign n_8392 = ~x_3108 & ~n_3673;
assign n_8393 = ~n_8391 & ~n_8392;
assign n_8394 =  x_3108 &  n_8393;
assign n_8395 = ~x_3108 & ~n_8393;
assign n_8396 = ~n_8394 & ~n_8395;
assign n_8397 = ~x_3107 & ~n_6063;
assign n_8398 =  x_3107 & ~n_8397;
assign n_8399 = ~x_3107 &  n_8397;
assign n_8400 = ~n_8398 & ~n_8399;
assign n_8401 =  n_1508 & ~n_1493;
assign n_8402 = ~n_1487 &  n_8401;
assign n_8403 = ~n_1481 &  n_8402;
assign n_8404 = ~n_1475 &  n_8403;
assign n_8405 = ~n_1469 &  n_8404;
assign n_8406 = ~n_1463 &  n_8405;
assign n_8407 = ~n_1457 &  n_8406;
assign n_8408 = ~n_1451 &  n_8407;
assign n_8409 = ~n_1445 &  n_8408;
assign n_8410 = ~n_1439 &  n_8409;
assign n_8411 = ~n_1433 &  n_8410;
assign n_8412 = ~n_1427 &  n_8411;
assign n_8413 = ~n_1421 &  n_8412;
assign n_8414 = ~n_1415 &  n_8413;
assign n_8415 = ~n_1409 &  n_8414;
assign n_8416 = ~n_1403 &  n_8415;
assign n_8417 = ~n_1397 &  n_8416;
assign n_8418 = ~n_1391 &  n_8417;
assign n_8419 = ~n_1385 &  n_8418;
assign n_8420 = ~n_1379 &  n_8419;
assign n_8421 = ~n_1373 &  n_8420;
assign n_8422 = ~n_1367 &  n_8421;
assign n_8423 = ~n_1361 &  n_8422;
assign n_8424 = ~n_1355 &  n_8423;
assign n_8425 = ~n_1349 &  n_8424;
assign n_8426 = ~n_1343 &  n_8425;
assign n_8427 = ~n_1337 &  n_8426;
assign n_8428 = ~n_1331 &  n_8427;
assign n_8429 = ~n_8428 &  n_3527;
assign n_8430 =  n_8428 & ~n_3527;
assign n_8431 = ~n_8429 & ~n_8430;
assign n_8432 =  x_3106 & ~n_8431;
assign n_8433 = ~x_3106 &  n_8431;
assign n_8434 = ~n_8432 & ~n_8433;
assign n_8435 =  x_3105 & ~n_3527;
assign n_8436 = ~x_3105 &  n_3527;
assign n_8437 = ~n_8435 & ~n_8436;
assign n_8438 =  n_1331 & ~n_8427;
assign n_8439 = ~n_8438 & ~n_8428;
assign n_8440 =  x_3104 & ~n_8439;
assign n_8441 = ~x_3104 &  n_8439;
assign n_8442 = ~n_8440 & ~n_8441;
assign n_8443 =  n_1337 & ~n_8426;
assign n_8444 = ~n_8443 & ~n_8427;
assign n_8445 =  x_3103 & ~n_8444;
assign n_8446 = ~x_3103 &  n_8444;
assign n_8447 = ~n_8445 & ~n_8446;
assign n_8448 =  n_1343 & ~n_8425;
assign n_8449 = ~n_8448 & ~n_8426;
assign n_8450 =  x_3102 & ~n_8449;
assign n_8451 = ~x_3102 &  n_8449;
assign n_8452 = ~n_8450 & ~n_8451;
assign n_8453 =  n_1349 & ~n_8424;
assign n_8454 = ~n_8453 & ~n_8425;
assign n_8455 =  x_3101 & ~n_8454;
assign n_8456 = ~x_3101 &  n_8454;
assign n_8457 = ~n_8455 & ~n_8456;
assign n_8458 =  n_1355 & ~n_8423;
assign n_8459 = ~n_8458 & ~n_8424;
assign n_8460 =  x_3100 & ~n_8459;
assign n_8461 = ~x_3100 &  n_8459;
assign n_8462 = ~n_8460 & ~n_8461;
assign n_8463 =  n_1361 & ~n_8422;
assign n_8464 = ~n_8463 & ~n_8423;
assign n_8465 =  x_3099 & ~n_8464;
assign n_8466 = ~x_3099 &  n_8464;
assign n_8467 = ~n_8465 & ~n_8466;
assign n_8468 =  n_1367 & ~n_8421;
assign n_8469 = ~n_8468 & ~n_8422;
assign n_8470 =  x_3098 & ~n_8469;
assign n_8471 = ~x_3098 &  n_8469;
assign n_8472 = ~n_8470 & ~n_8471;
assign n_8473 =  n_1373 & ~n_8420;
assign n_8474 = ~n_8473 & ~n_8421;
assign n_8475 =  x_3097 & ~n_8474;
assign n_8476 = ~x_3097 &  n_8474;
assign n_8477 = ~n_8475 & ~n_8476;
assign n_8478 =  n_1379 & ~n_8419;
assign n_8479 = ~n_8478 & ~n_8420;
assign n_8480 =  x_3096 & ~n_8479;
assign n_8481 = ~x_3096 &  n_8479;
assign n_8482 = ~n_8480 & ~n_8481;
assign n_8483 =  n_1385 & ~n_8418;
assign n_8484 = ~n_8483 & ~n_8419;
assign n_8485 =  x_3095 & ~n_8484;
assign n_8486 = ~x_3095 &  n_8484;
assign n_8487 = ~n_8485 & ~n_8486;
assign n_8488 =  n_1391 & ~n_8417;
assign n_8489 = ~n_8488 & ~n_8418;
assign n_8490 =  x_3094 & ~n_8489;
assign n_8491 = ~x_3094 &  n_8489;
assign n_8492 = ~n_8490 & ~n_8491;
assign n_8493 =  n_1397 & ~n_8416;
assign n_8494 = ~n_8493 & ~n_8417;
assign n_8495 =  x_3093 & ~n_8494;
assign n_8496 = ~x_3093 &  n_8494;
assign n_8497 = ~n_8495 & ~n_8496;
assign n_8498 =  n_1403 & ~n_8415;
assign n_8499 = ~n_8498 & ~n_8416;
assign n_8500 =  x_3092 & ~n_8499;
assign n_8501 = ~x_3092 &  n_8499;
assign n_8502 = ~n_8500 & ~n_8501;
assign n_8503 =  n_1409 & ~n_8414;
assign n_8504 = ~n_8503 & ~n_8415;
assign n_8505 =  x_3091 & ~n_8504;
assign n_8506 = ~x_3091 &  n_8504;
assign n_8507 = ~n_8505 & ~n_8506;
assign n_8508 =  n_1415 & ~n_8413;
assign n_8509 = ~n_8508 & ~n_8414;
assign n_8510 =  x_3090 & ~n_8509;
assign n_8511 = ~x_3090 &  n_8509;
assign n_8512 = ~n_8510 & ~n_8511;
assign n_8513 =  n_1421 & ~n_8412;
assign n_8514 = ~n_8513 & ~n_8413;
assign n_8515 =  x_3089 & ~n_8514;
assign n_8516 = ~x_3089 &  n_8514;
assign n_8517 = ~n_8515 & ~n_8516;
assign n_8518 =  n_1427 & ~n_8411;
assign n_8519 = ~n_8518 & ~n_8412;
assign n_8520 =  x_3088 & ~n_8519;
assign n_8521 = ~x_3088 &  n_8519;
assign n_8522 = ~n_8520 & ~n_8521;
assign n_8523 =  n_1433 & ~n_8410;
assign n_8524 = ~n_8523 & ~n_8411;
assign n_8525 =  x_3087 & ~n_8524;
assign n_8526 = ~x_3087 &  n_8524;
assign n_8527 = ~n_8525 & ~n_8526;
assign n_8528 =  n_1439 & ~n_8409;
assign n_8529 = ~n_8528 & ~n_8410;
assign n_8530 =  x_3086 & ~n_8529;
assign n_8531 = ~x_3086 &  n_8529;
assign n_8532 = ~n_8530 & ~n_8531;
assign n_8533 =  n_1445 & ~n_8408;
assign n_8534 = ~n_8533 & ~n_8409;
assign n_8535 =  x_3085 & ~n_8534;
assign n_8536 = ~x_3085 &  n_8534;
assign n_8537 = ~n_8535 & ~n_8536;
assign n_8538 =  n_1451 & ~n_8407;
assign n_8539 = ~n_8538 & ~n_8408;
assign n_8540 =  x_3084 & ~n_8539;
assign n_8541 = ~x_3084 &  n_8539;
assign n_8542 = ~n_8540 & ~n_8541;
assign n_8543 =  n_1457 & ~n_8406;
assign n_8544 = ~n_8543 & ~n_8407;
assign n_8545 =  x_3083 & ~n_8544;
assign n_8546 = ~x_3083 &  n_8544;
assign n_8547 = ~n_8545 & ~n_8546;
assign n_8548 =  n_1463 & ~n_8405;
assign n_8549 = ~n_8548 & ~n_8406;
assign n_8550 =  x_3082 & ~n_8549;
assign n_8551 = ~x_3082 &  n_8549;
assign n_8552 = ~n_8550 & ~n_8551;
assign n_8553 =  n_1469 & ~n_8404;
assign n_8554 = ~n_8553 & ~n_8405;
assign n_8555 =  x_3081 & ~n_8554;
assign n_8556 = ~x_3081 &  n_8554;
assign n_8557 = ~n_8555 & ~n_8556;
assign n_8558 =  n_1475 & ~n_8403;
assign n_8559 = ~n_8558 & ~n_8404;
assign n_8560 =  x_3080 & ~n_8559;
assign n_8561 = ~x_3080 &  n_8559;
assign n_8562 = ~n_8560 & ~n_8561;
assign n_8563 =  n_1481 & ~n_8402;
assign n_8564 = ~n_8563 & ~n_8403;
assign n_8565 =  x_3079 & ~n_8564;
assign n_8566 = ~x_3079 &  n_8564;
assign n_8567 = ~n_8565 & ~n_8566;
assign n_8568 =  n_1487 & ~n_8401;
assign n_8569 = ~n_8568 & ~n_8402;
assign n_8570 =  x_3078 & ~n_8569;
assign n_8571 = ~x_3078 &  n_8569;
assign n_8572 = ~n_8570 & ~n_8571;
assign n_8573 = ~n_1508 &  n_1493;
assign n_8574 = ~n_8573 & ~n_8401;
assign n_8575 =  x_3077 & ~n_8574;
assign n_8576 = ~x_3077 &  n_8574;
assign n_8577 = ~n_8575 & ~n_8576;
assign n_8578 = ~n_1502 &  n_1505;
assign n_8579 = ~n_1506 & ~n_8578;
assign n_8580 =  x_3076 &  n_8579;
assign n_8581 = ~x_3076 & ~n_8579;
assign n_8582 = ~n_8580 & ~n_8581;
assign n_8583 =  x_3074 &  n_1328;
assign n_8584 = ~x_3075 & ~n_8583;
assign n_8585 = ~n_6073 & ~n_8584;
assign n_8586 =  x_3075 &  n_8585;
assign n_8587 = ~x_3075 & ~n_8585;
assign n_8588 = ~n_8586 & ~n_8587;
assign n_8589 =  x_3074 & ~n_6074;
assign n_8590 = ~n_6064 & ~n_8589;
assign n_8591 =  x_3074 & ~n_8590;
assign n_8592 = ~x_3074 &  n_8590;
assign n_8593 = ~n_8591 & ~n_8592;
assign n_8594 =  x_1729 & ~n_1325;
assign n_8595 =  x_3073 &  n_1325;
assign n_8596 = ~n_8594 & ~n_8595;
assign n_8597 =  x_3073 & ~n_8596;
assign n_8598 = ~x_3073 &  n_8596;
assign n_8599 = ~n_8597 & ~n_8598;
assign n_8600 =  x_3072 & ~n_6090;
assign n_8601 = ~n_8600 & ~n_6033;
assign n_8602 =  x_3072 & ~n_8601;
assign n_8603 = ~x_3072 &  n_8601;
assign n_8604 = ~n_8602 & ~n_8603;
assign n_8605 = ~n_6029 &  n_6034;
assign n_8606 =  x_3071 & ~n_6091;
assign n_8607 = ~n_8605 & ~n_8606;
assign n_8608 =  x_3071 & ~n_8607;
assign n_8609 = ~x_3071 &  n_8607;
assign n_8610 = ~n_8608 & ~n_8609;
assign n_8611 =  x_1726 & ~n_3676;
assign n_8612 =  x_3070 &  n_3676;
assign n_8613 = ~n_8611 & ~n_8612;
assign n_8614 =  x_3070 & ~n_8613;
assign n_8615 = ~x_3070 &  n_8613;
assign n_8616 = ~n_8614 & ~n_8615;
assign n_8617 = ~x_3069 &  n_3676;
assign n_8618 = ~n_6031 & ~n_8617;
assign n_8619 =  x_3069 &  n_8618;
assign n_8620 = ~x_3069 & ~n_8618;
assign n_8621 = ~n_8619 & ~n_8620;
assign n_8622 = ~x_2544 &  n_6008;
assign n_8623 = ~n_4374 &  n_5728;
assign n_8624 =  n_4370 &  n_8623;
assign n_8625 = ~n_8622 & ~n_8624;
assign n_8626 = ~x_2553 & ~n_8625;
assign n_8627 =  x_2554 &  n_8626;
assign n_8628 =  x_2555 &  x_2556;
assign n_8629 =  n_8627 &  n_8628;
assign n_8630 =  x_3068 & ~n_8629;
assign n_8631 =  x_1559 &  n_8629;
assign n_8632 = ~n_8630 & ~n_8631;
assign n_8633 =  x_3068 & ~n_8632;
assign n_8634 = ~x_3068 &  n_8632;
assign n_8635 = ~n_8633 & ~n_8634;
assign n_8636 =  x_2553 & ~n_8625;
assign n_8637 = ~x_2554 &  n_8628;
assign n_8638 =  n_8636 &  n_8637;
assign n_8639 =  x_3067 & ~n_8638;
assign n_8640 =  x_1559 &  n_8638;
assign n_8641 = ~n_8639 & ~n_8640;
assign n_8642 =  x_3067 & ~n_8641;
assign n_8643 = ~x_3067 &  n_8641;
assign n_8644 = ~n_8642 & ~n_8643;
assign n_8645 =  n_8626 &  n_8637;
assign n_8646 =  x_3066 & ~n_8645;
assign n_8647 =  x_1559 &  n_8645;
assign n_8648 = ~n_8646 & ~n_8647;
assign n_8649 =  x_3066 & ~n_8648;
assign n_8650 = ~x_3066 &  n_8648;
assign n_8651 = ~n_8649 & ~n_8650;
assign n_8652 =  x_2554 &  n_8636;
assign n_8653 = ~x_2555 &  x_2556;
assign n_8654 =  n_8652 &  n_8653;
assign n_8655 =  x_3065 & ~n_8654;
assign n_8656 =  x_1559 &  n_8654;
assign n_8657 = ~n_8655 & ~n_8656;
assign n_8658 =  x_3065 & ~n_8657;
assign n_8659 = ~x_3065 &  n_8657;
assign n_8660 = ~n_8658 & ~n_8659;
assign n_8661 =  n_8627 &  n_8653;
assign n_8662 =  x_3064 & ~n_8661;
assign n_8663 =  x_1559 &  n_8661;
assign n_8664 = ~n_8662 & ~n_8663;
assign n_8665 =  x_3064 & ~n_8664;
assign n_8666 = ~x_3064 &  n_8664;
assign n_8667 = ~n_8665 & ~n_8666;
assign n_8668 = ~x_2554 &  n_8653;
assign n_8669 =  n_8636 &  n_8668;
assign n_8670 =  x_3063 & ~n_8669;
assign n_8671 =  x_1559 &  n_8669;
assign n_8672 = ~n_8670 & ~n_8671;
assign n_8673 =  x_3063 & ~n_8672;
assign n_8674 = ~x_3063 &  n_8672;
assign n_8675 = ~n_8673 & ~n_8674;
assign n_8676 =  n_8626 &  n_8668;
assign n_8677 =  x_3062 & ~n_8676;
assign n_8678 =  x_1559 &  n_8676;
assign n_8679 = ~n_8677 & ~n_8678;
assign n_8680 =  x_3062 & ~n_8679;
assign n_8681 = ~x_3062 &  n_8679;
assign n_8682 = ~n_8680 & ~n_8681;
assign n_8683 =  x_2555 & ~x_2556;
assign n_8684 =  n_8652 &  n_8683;
assign n_8685 =  x_3061 & ~n_8684;
assign n_8686 =  x_1559 &  n_8684;
assign n_8687 = ~n_8685 & ~n_8686;
assign n_8688 =  x_3061 & ~n_8687;
assign n_8689 = ~x_3061 &  n_8687;
assign n_8690 = ~n_8688 & ~n_8689;
assign n_8691 =  n_8683 &  n_8627;
assign n_8692 =  x_3060 & ~n_8691;
assign n_8693 =  x_1559 &  n_8691;
assign n_8694 = ~n_8692 & ~n_8693;
assign n_8695 =  x_3060 & ~n_8694;
assign n_8696 = ~x_3060 &  n_8694;
assign n_8697 = ~n_8695 & ~n_8696;
assign n_8698 = ~x_2554 &  n_8683;
assign n_8699 =  n_8636 &  n_8698;
assign n_8700 =  x_3059 & ~n_8699;
assign n_8701 =  x_1559 &  n_8699;
assign n_8702 = ~n_8700 & ~n_8701;
assign n_8703 =  x_3059 & ~n_8702;
assign n_8704 = ~x_3059 &  n_8702;
assign n_8705 = ~n_8703 & ~n_8704;
assign n_8706 =  n_8626 &  n_8698;
assign n_8707 =  x_3058 & ~n_8706;
assign n_8708 =  x_1559 &  n_8706;
assign n_8709 = ~n_8707 & ~n_8708;
assign n_8710 =  x_3058 & ~n_8709;
assign n_8711 = ~x_3058 &  n_8709;
assign n_8712 = ~n_8710 & ~n_8711;
assign n_8713 = ~x_2555 & ~x_2556;
assign n_8714 =  n_8652 &  n_8713;
assign n_8715 =  x_3057 & ~n_8714;
assign n_8716 =  x_1559 &  n_8714;
assign n_8717 = ~n_8715 & ~n_8716;
assign n_8718 =  x_3057 & ~n_8717;
assign n_8719 = ~x_3057 &  n_8717;
assign n_8720 = ~n_8718 & ~n_8719;
assign n_8721 =  n_8713 &  n_8627;
assign n_8722 =  x_3056 & ~n_8721;
assign n_8723 =  x_1559 &  n_8721;
assign n_8724 = ~n_8722 & ~n_8723;
assign n_8725 =  x_3056 & ~n_8724;
assign n_8726 = ~x_3056 &  n_8724;
assign n_8727 = ~n_8725 & ~n_8726;
assign n_8728 = ~x_2554 &  n_8713;
assign n_8729 =  n_8636 &  n_8728;
assign n_8730 =  x_3055 & ~n_8729;
assign n_8731 =  x_1559 &  n_8729;
assign n_8732 = ~n_8730 & ~n_8731;
assign n_8733 =  x_3055 & ~n_8732;
assign n_8734 = ~x_3055 &  n_8732;
assign n_8735 = ~n_8733 & ~n_8734;
assign n_8736 =  n_8626 &  n_8728;
assign n_8737 =  x_3054 & ~n_8736;
assign n_8738 =  x_1559 &  n_8736;
assign n_8739 = ~n_8737 & ~n_8738;
assign n_8740 =  x_3054 & ~n_8739;
assign n_8741 = ~x_3054 &  n_8739;
assign n_8742 = ~n_8740 & ~n_8741;
assign n_8743 =  x_2555 &  n_8652;
assign n_8744 =  x_2556 &  n_8743;
assign n_8745 =  x_3053 & ~n_8744;
assign n_8746 =  x_1559 &  n_8744;
assign n_8747 = ~n_8745 & ~n_8746;
assign n_8748 =  x_3053 & ~n_8747;
assign n_8749 = ~x_3053 &  n_8747;
assign n_8750 = ~n_8748 & ~n_8749;
assign n_8751 =  x_3052 & ~n_8629;
assign n_8752 =  x_1558 &  n_8629;
assign n_8753 = ~n_8751 & ~n_8752;
assign n_8754 =  x_3052 & ~n_8753;
assign n_8755 = ~x_3052 &  n_8753;
assign n_8756 = ~n_8754 & ~n_8755;
assign n_8757 =  x_3051 & ~n_8638;
assign n_8758 =  x_1558 &  n_8638;
assign n_8759 = ~n_8757 & ~n_8758;
assign n_8760 =  x_3051 & ~n_8759;
assign n_8761 = ~x_3051 &  n_8759;
assign n_8762 = ~n_8760 & ~n_8761;
assign n_8763 =  x_3050 & ~n_8645;
assign n_8764 =  x_1558 &  n_8645;
assign n_8765 = ~n_8763 & ~n_8764;
assign n_8766 =  x_3050 & ~n_8765;
assign n_8767 = ~x_3050 &  n_8765;
assign n_8768 = ~n_8766 & ~n_8767;
assign n_8769 =  x_3049 & ~n_8654;
assign n_8770 =  x_1558 &  n_8654;
assign n_8771 = ~n_8769 & ~n_8770;
assign n_8772 =  x_3049 & ~n_8771;
assign n_8773 = ~x_3049 &  n_8771;
assign n_8774 = ~n_8772 & ~n_8773;
assign n_8775 =  x_3048 & ~n_8661;
assign n_8776 =  x_1558 &  n_8661;
assign n_8777 = ~n_8775 & ~n_8776;
assign n_8778 =  x_3048 & ~n_8777;
assign n_8779 = ~x_3048 &  n_8777;
assign n_8780 = ~n_8778 & ~n_8779;
assign n_8781 =  x_3047 & ~n_8669;
assign n_8782 =  x_1558 &  n_8669;
assign n_8783 = ~n_8781 & ~n_8782;
assign n_8784 =  x_3047 & ~n_8783;
assign n_8785 = ~x_3047 &  n_8783;
assign n_8786 = ~n_8784 & ~n_8785;
assign n_8787 =  x_3046 & ~n_8676;
assign n_8788 =  x_1558 &  n_8676;
assign n_8789 = ~n_8787 & ~n_8788;
assign n_8790 =  x_3046 & ~n_8789;
assign n_8791 = ~x_3046 &  n_8789;
assign n_8792 = ~n_8790 & ~n_8791;
assign n_8793 =  x_3045 & ~n_8684;
assign n_8794 =  x_1558 &  n_8684;
assign n_8795 = ~n_8793 & ~n_8794;
assign n_8796 =  x_3045 & ~n_8795;
assign n_8797 = ~x_3045 &  n_8795;
assign n_8798 = ~n_8796 & ~n_8797;
assign n_8799 =  x_3044 & ~n_8691;
assign n_8800 =  x_1558 &  n_8691;
assign n_8801 = ~n_8799 & ~n_8800;
assign n_8802 =  x_3044 & ~n_8801;
assign n_8803 = ~x_3044 &  n_8801;
assign n_8804 = ~n_8802 & ~n_8803;
assign n_8805 =  x_3043 & ~n_8699;
assign n_8806 =  x_1558 &  n_8699;
assign n_8807 = ~n_8805 & ~n_8806;
assign n_8808 =  x_3043 & ~n_8807;
assign n_8809 = ~x_3043 &  n_8807;
assign n_8810 = ~n_8808 & ~n_8809;
assign n_8811 =  x_3042 & ~n_8706;
assign n_8812 =  x_1558 &  n_8706;
assign n_8813 = ~n_8811 & ~n_8812;
assign n_8814 =  x_3042 & ~n_8813;
assign n_8815 = ~x_3042 &  n_8813;
assign n_8816 = ~n_8814 & ~n_8815;
assign n_8817 =  x_3041 & ~n_8714;
assign n_8818 =  x_1558 &  n_8714;
assign n_8819 = ~n_8817 & ~n_8818;
assign n_8820 =  x_3041 & ~n_8819;
assign n_8821 = ~x_3041 &  n_8819;
assign n_8822 = ~n_8820 & ~n_8821;
assign n_8823 =  x_3040 & ~n_8721;
assign n_8824 =  x_1558 &  n_8721;
assign n_8825 = ~n_8823 & ~n_8824;
assign n_8826 =  x_3040 & ~n_8825;
assign n_8827 = ~x_3040 &  n_8825;
assign n_8828 = ~n_8826 & ~n_8827;
assign n_8829 =  x_3039 & ~n_8729;
assign n_8830 =  x_1558 &  n_8729;
assign n_8831 = ~n_8829 & ~n_8830;
assign n_8832 =  x_3039 & ~n_8831;
assign n_8833 = ~x_3039 &  n_8831;
assign n_8834 = ~n_8832 & ~n_8833;
assign n_8835 =  x_3038 & ~n_8736;
assign n_8836 =  x_1558 &  n_8736;
assign n_8837 = ~n_8835 & ~n_8836;
assign n_8838 =  x_3038 & ~n_8837;
assign n_8839 = ~x_3038 &  n_8837;
assign n_8840 = ~n_8838 & ~n_8839;
assign n_8841 =  x_3037 & ~n_8744;
assign n_8842 =  x_1558 &  n_8744;
assign n_8843 = ~n_8841 & ~n_8842;
assign n_8844 =  x_3037 & ~n_8843;
assign n_8845 = ~x_3037 &  n_8843;
assign n_8846 = ~n_8844 & ~n_8845;
assign n_8847 =  x_3036 & ~n_8629;
assign n_8848 =  x_1501 &  n_8629;
assign n_8849 = ~n_8847 & ~n_8848;
assign n_8850 =  x_3036 & ~n_8849;
assign n_8851 = ~x_3036 &  n_8849;
assign n_8852 = ~n_8850 & ~n_8851;
assign n_8853 =  x_3035 & ~n_8638;
assign n_8854 =  x_1501 &  n_8638;
assign n_8855 = ~n_8853 & ~n_8854;
assign n_8856 =  x_3035 & ~n_8855;
assign n_8857 = ~x_3035 &  n_8855;
assign n_8858 = ~n_8856 & ~n_8857;
assign n_8859 =  x_3034 & ~n_8645;
assign n_8860 =  x_1501 &  n_8645;
assign n_8861 = ~n_8859 & ~n_8860;
assign n_8862 =  x_3034 & ~n_8861;
assign n_8863 = ~x_3034 &  n_8861;
assign n_8864 = ~n_8862 & ~n_8863;
assign n_8865 =  x_3033 & ~n_8654;
assign n_8866 =  x_1501 &  n_8654;
assign n_8867 = ~n_8865 & ~n_8866;
assign n_8868 =  x_3033 & ~n_8867;
assign n_8869 = ~x_3033 &  n_8867;
assign n_8870 = ~n_8868 & ~n_8869;
assign n_8871 =  x_3032 & ~n_8661;
assign n_8872 =  x_1501 &  n_8661;
assign n_8873 = ~n_8871 & ~n_8872;
assign n_8874 =  x_3032 & ~n_8873;
assign n_8875 = ~x_3032 &  n_8873;
assign n_8876 = ~n_8874 & ~n_8875;
assign n_8877 =  x_3031 & ~n_8669;
assign n_8878 =  x_1501 &  n_8669;
assign n_8879 = ~n_8877 & ~n_8878;
assign n_8880 =  x_3031 & ~n_8879;
assign n_8881 = ~x_3031 &  n_8879;
assign n_8882 = ~n_8880 & ~n_8881;
assign n_8883 =  x_3030 & ~n_8676;
assign n_8884 =  x_1501 &  n_8676;
assign n_8885 = ~n_8883 & ~n_8884;
assign n_8886 =  x_3030 & ~n_8885;
assign n_8887 = ~x_3030 &  n_8885;
assign n_8888 = ~n_8886 & ~n_8887;
assign n_8889 =  x_3029 & ~n_8684;
assign n_8890 =  x_1501 &  n_8684;
assign n_8891 = ~n_8889 & ~n_8890;
assign n_8892 =  x_3029 & ~n_8891;
assign n_8893 = ~x_3029 &  n_8891;
assign n_8894 = ~n_8892 & ~n_8893;
assign n_8895 =  x_3028 & ~n_8691;
assign n_8896 =  x_1501 &  n_8691;
assign n_8897 = ~n_8895 & ~n_8896;
assign n_8898 =  x_3028 & ~n_8897;
assign n_8899 = ~x_3028 &  n_8897;
assign n_8900 = ~n_8898 & ~n_8899;
assign n_8901 =  x_3027 & ~n_8699;
assign n_8902 =  x_1501 &  n_8699;
assign n_8903 = ~n_8901 & ~n_8902;
assign n_8904 =  x_3027 & ~n_8903;
assign n_8905 = ~x_3027 &  n_8903;
assign n_8906 = ~n_8904 & ~n_8905;
assign n_8907 =  x_3026 & ~n_8706;
assign n_8908 =  x_1501 &  n_8706;
assign n_8909 = ~n_8907 & ~n_8908;
assign n_8910 =  x_3026 & ~n_8909;
assign n_8911 = ~x_3026 &  n_8909;
assign n_8912 = ~n_8910 & ~n_8911;
assign n_8913 =  x_3025 & ~n_8714;
assign n_8914 =  x_1501 &  n_8714;
assign n_8915 = ~n_8913 & ~n_8914;
assign n_8916 =  x_3025 & ~n_8915;
assign n_8917 = ~x_3025 &  n_8915;
assign n_8918 = ~n_8916 & ~n_8917;
assign n_8919 =  x_3024 & ~n_8721;
assign n_8920 =  x_1501 &  n_8721;
assign n_8921 = ~n_8919 & ~n_8920;
assign n_8922 =  x_3024 & ~n_8921;
assign n_8923 = ~x_3024 &  n_8921;
assign n_8924 = ~n_8922 & ~n_8923;
assign n_8925 =  x_3023 & ~n_8729;
assign n_8926 =  x_1501 &  n_8729;
assign n_8927 = ~n_8925 & ~n_8926;
assign n_8928 =  x_3023 & ~n_8927;
assign n_8929 = ~x_3023 &  n_8927;
assign n_8930 = ~n_8928 & ~n_8929;
assign n_8931 =  x_3022 & ~n_8736;
assign n_8932 =  x_1501 &  n_8736;
assign n_8933 = ~n_8931 & ~n_8932;
assign n_8934 =  x_3022 & ~n_8933;
assign n_8935 = ~x_3022 &  n_8933;
assign n_8936 = ~n_8934 & ~n_8935;
assign n_8937 =  x_3021 & ~n_8744;
assign n_8938 =  x_1501 &  n_8744;
assign n_8939 = ~n_8937 & ~n_8938;
assign n_8940 =  x_3021 & ~n_8939;
assign n_8941 = ~x_3021 &  n_8939;
assign n_8942 = ~n_8940 & ~n_8941;
assign n_8943 =  x_3020 & ~n_8629;
assign n_8944 =  x_1502 &  n_8629;
assign n_8945 = ~n_8943 & ~n_8944;
assign n_8946 =  x_3020 & ~n_8945;
assign n_8947 = ~x_3020 &  n_8945;
assign n_8948 = ~n_8946 & ~n_8947;
assign n_8949 =  x_3019 & ~n_8638;
assign n_8950 =  x_1502 &  n_8638;
assign n_8951 = ~n_8949 & ~n_8950;
assign n_8952 =  x_3019 & ~n_8951;
assign n_8953 = ~x_3019 &  n_8951;
assign n_8954 = ~n_8952 & ~n_8953;
assign n_8955 =  x_3018 & ~n_8645;
assign n_8956 =  x_1502 &  n_8645;
assign n_8957 = ~n_8955 & ~n_8956;
assign n_8958 =  x_3018 & ~n_8957;
assign n_8959 = ~x_3018 &  n_8957;
assign n_8960 = ~n_8958 & ~n_8959;
assign n_8961 =  x_3017 & ~n_8654;
assign n_8962 =  x_1502 &  n_8654;
assign n_8963 = ~n_8961 & ~n_8962;
assign n_8964 =  x_3017 & ~n_8963;
assign n_8965 = ~x_3017 &  n_8963;
assign n_8966 = ~n_8964 & ~n_8965;
assign n_8967 =  x_3016 & ~n_8661;
assign n_8968 =  x_1502 &  n_8661;
assign n_8969 = ~n_8967 & ~n_8968;
assign n_8970 =  x_3016 & ~n_8969;
assign n_8971 = ~x_3016 &  n_8969;
assign n_8972 = ~n_8970 & ~n_8971;
assign n_8973 =  x_3015 & ~n_8669;
assign n_8974 =  x_1502 &  n_8669;
assign n_8975 = ~n_8973 & ~n_8974;
assign n_8976 =  x_3015 & ~n_8975;
assign n_8977 = ~x_3015 &  n_8975;
assign n_8978 = ~n_8976 & ~n_8977;
assign n_8979 =  x_3014 & ~n_8676;
assign n_8980 =  x_1502 &  n_8676;
assign n_8981 = ~n_8979 & ~n_8980;
assign n_8982 =  x_3014 & ~n_8981;
assign n_8983 = ~x_3014 &  n_8981;
assign n_8984 = ~n_8982 & ~n_8983;
assign n_8985 =  x_3013 & ~n_8684;
assign n_8986 =  x_1502 &  n_8684;
assign n_8987 = ~n_8985 & ~n_8986;
assign n_8988 =  x_3013 & ~n_8987;
assign n_8989 = ~x_3013 &  n_8987;
assign n_8990 = ~n_8988 & ~n_8989;
assign n_8991 =  x_3012 & ~n_8691;
assign n_8992 =  x_1502 &  n_8691;
assign n_8993 = ~n_8991 & ~n_8992;
assign n_8994 =  x_3012 & ~n_8993;
assign n_8995 = ~x_3012 &  n_8993;
assign n_8996 = ~n_8994 & ~n_8995;
assign n_8997 =  x_3011 & ~n_8699;
assign n_8998 =  x_1502 &  n_8699;
assign n_8999 = ~n_8997 & ~n_8998;
assign n_9000 =  x_3011 & ~n_8999;
assign n_9001 = ~x_3011 &  n_8999;
assign n_9002 = ~n_9000 & ~n_9001;
assign n_9003 =  x_3010 & ~n_8706;
assign n_9004 =  x_1502 &  n_8706;
assign n_9005 = ~n_9003 & ~n_9004;
assign n_9006 =  x_3010 & ~n_9005;
assign n_9007 = ~x_3010 &  n_9005;
assign n_9008 = ~n_9006 & ~n_9007;
assign n_9009 =  x_3009 & ~n_8714;
assign n_9010 =  x_1502 &  n_8714;
assign n_9011 = ~n_9009 & ~n_9010;
assign n_9012 =  x_3009 & ~n_9011;
assign n_9013 = ~x_3009 &  n_9011;
assign n_9014 = ~n_9012 & ~n_9013;
assign n_9015 =  x_3008 & ~n_8721;
assign n_9016 =  x_1502 &  n_8721;
assign n_9017 = ~n_9015 & ~n_9016;
assign n_9018 =  x_3008 & ~n_9017;
assign n_9019 = ~x_3008 &  n_9017;
assign n_9020 = ~n_9018 & ~n_9019;
assign n_9021 =  x_3007 & ~n_8729;
assign n_9022 =  x_1502 &  n_8729;
assign n_9023 = ~n_9021 & ~n_9022;
assign n_9024 =  x_3007 & ~n_9023;
assign n_9025 = ~x_3007 &  n_9023;
assign n_9026 = ~n_9024 & ~n_9025;
assign n_9027 =  x_3006 & ~n_8736;
assign n_9028 =  x_1502 &  n_8736;
assign n_9029 = ~n_9027 & ~n_9028;
assign n_9030 =  x_3006 & ~n_9029;
assign n_9031 = ~x_3006 &  n_9029;
assign n_9032 = ~n_9030 & ~n_9031;
assign n_9033 =  x_3005 & ~n_8744;
assign n_9034 =  x_1502 &  n_8744;
assign n_9035 = ~n_9033 & ~n_9034;
assign n_9036 =  x_3005 & ~n_9035;
assign n_9037 = ~x_3005 &  n_9035;
assign n_9038 = ~n_9036 & ~n_9037;
assign n_9039 =  x_3004 & ~n_8629;
assign n_9040 =  x_1503 &  n_8629;
assign n_9041 = ~n_9039 & ~n_9040;
assign n_9042 =  x_3004 & ~n_9041;
assign n_9043 = ~x_3004 &  n_9041;
assign n_9044 = ~n_9042 & ~n_9043;
assign n_9045 =  x_3003 & ~n_8638;
assign n_9046 =  x_1503 &  n_8638;
assign n_9047 = ~n_9045 & ~n_9046;
assign n_9048 =  x_3003 & ~n_9047;
assign n_9049 = ~x_3003 &  n_9047;
assign n_9050 = ~n_9048 & ~n_9049;
assign n_9051 =  x_3002 & ~n_8645;
assign n_9052 =  x_1503 &  n_8645;
assign n_9053 = ~n_9051 & ~n_9052;
assign n_9054 =  x_3002 & ~n_9053;
assign n_9055 = ~x_3002 &  n_9053;
assign n_9056 = ~n_9054 & ~n_9055;
assign n_9057 =  x_3001 & ~n_8654;
assign n_9058 =  x_1503 &  n_8654;
assign n_9059 = ~n_9057 & ~n_9058;
assign n_9060 =  x_3001 & ~n_9059;
assign n_9061 = ~x_3001 &  n_9059;
assign n_9062 = ~n_9060 & ~n_9061;
assign n_9063 =  x_3000 & ~n_8661;
assign n_9064 =  x_1503 &  n_8661;
assign n_9065 = ~n_9063 & ~n_9064;
assign n_9066 =  x_3000 & ~n_9065;
assign n_9067 = ~x_3000 &  n_9065;
assign n_9068 = ~n_9066 & ~n_9067;
assign n_9069 =  x_2999 & ~n_8669;
assign n_9070 =  x_1503 &  n_8669;
assign n_9071 = ~n_9069 & ~n_9070;
assign n_9072 =  x_2999 & ~n_9071;
assign n_9073 = ~x_2999 &  n_9071;
assign n_9074 = ~n_9072 & ~n_9073;
assign n_9075 =  x_2998 & ~n_8676;
assign n_9076 =  x_1503 &  n_8676;
assign n_9077 = ~n_9075 & ~n_9076;
assign n_9078 =  x_2998 & ~n_9077;
assign n_9079 = ~x_2998 &  n_9077;
assign n_9080 = ~n_9078 & ~n_9079;
assign n_9081 =  x_2997 & ~n_8684;
assign n_9082 =  x_1503 &  n_8684;
assign n_9083 = ~n_9081 & ~n_9082;
assign n_9084 =  x_2997 & ~n_9083;
assign n_9085 = ~x_2997 &  n_9083;
assign n_9086 = ~n_9084 & ~n_9085;
assign n_9087 =  x_2996 & ~n_8691;
assign n_9088 =  x_1503 &  n_8691;
assign n_9089 = ~n_9087 & ~n_9088;
assign n_9090 =  x_2996 & ~n_9089;
assign n_9091 = ~x_2996 &  n_9089;
assign n_9092 = ~n_9090 & ~n_9091;
assign n_9093 =  x_2995 & ~n_8699;
assign n_9094 =  x_1503 &  n_8699;
assign n_9095 = ~n_9093 & ~n_9094;
assign n_9096 =  x_2995 & ~n_9095;
assign n_9097 = ~x_2995 &  n_9095;
assign n_9098 = ~n_9096 & ~n_9097;
assign n_9099 =  x_2994 & ~n_8706;
assign n_9100 =  x_1503 &  n_8706;
assign n_9101 = ~n_9099 & ~n_9100;
assign n_9102 =  x_2994 & ~n_9101;
assign n_9103 = ~x_2994 &  n_9101;
assign n_9104 = ~n_9102 & ~n_9103;
assign n_9105 =  x_2993 & ~n_8714;
assign n_9106 =  x_1503 &  n_8714;
assign n_9107 = ~n_9105 & ~n_9106;
assign n_9108 =  x_2993 & ~n_9107;
assign n_9109 = ~x_2993 &  n_9107;
assign n_9110 = ~n_9108 & ~n_9109;
assign n_9111 =  x_2992 & ~n_8721;
assign n_9112 =  x_1503 &  n_8721;
assign n_9113 = ~n_9111 & ~n_9112;
assign n_9114 =  x_2992 & ~n_9113;
assign n_9115 = ~x_2992 &  n_9113;
assign n_9116 = ~n_9114 & ~n_9115;
assign n_9117 =  x_2991 & ~n_8729;
assign n_9118 =  x_1503 &  n_8729;
assign n_9119 = ~n_9117 & ~n_9118;
assign n_9120 =  x_2991 & ~n_9119;
assign n_9121 = ~x_2991 &  n_9119;
assign n_9122 = ~n_9120 & ~n_9121;
assign n_9123 =  x_2990 & ~n_8736;
assign n_9124 =  x_1503 &  n_8736;
assign n_9125 = ~n_9123 & ~n_9124;
assign n_9126 =  x_2990 & ~n_9125;
assign n_9127 = ~x_2990 &  n_9125;
assign n_9128 = ~n_9126 & ~n_9127;
assign n_9129 =  x_2989 & ~n_8744;
assign n_9130 =  x_1503 &  n_8744;
assign n_9131 = ~n_9129 & ~n_9130;
assign n_9132 =  x_2989 & ~n_9131;
assign n_9133 = ~x_2989 &  n_9131;
assign n_9134 = ~n_9132 & ~n_9133;
assign n_9135 =  x_2988 & ~n_8629;
assign n_9136 =  x_1504 &  n_8629;
assign n_9137 = ~n_9135 & ~n_9136;
assign n_9138 =  x_2988 & ~n_9137;
assign n_9139 = ~x_2988 &  n_9137;
assign n_9140 = ~n_9138 & ~n_9139;
assign n_9141 =  x_2987 & ~n_8638;
assign n_9142 =  x_1504 &  n_8638;
assign n_9143 = ~n_9141 & ~n_9142;
assign n_9144 =  x_2987 & ~n_9143;
assign n_9145 = ~x_2987 &  n_9143;
assign n_9146 = ~n_9144 & ~n_9145;
assign n_9147 =  x_2986 & ~n_8645;
assign n_9148 =  x_1504 &  n_8645;
assign n_9149 = ~n_9147 & ~n_9148;
assign n_9150 =  x_2986 & ~n_9149;
assign n_9151 = ~x_2986 &  n_9149;
assign n_9152 = ~n_9150 & ~n_9151;
assign n_9153 =  x_2985 & ~n_8654;
assign n_9154 =  x_1504 &  n_8654;
assign n_9155 = ~n_9153 & ~n_9154;
assign n_9156 =  x_2985 & ~n_9155;
assign n_9157 = ~x_2985 &  n_9155;
assign n_9158 = ~n_9156 & ~n_9157;
assign n_9159 =  x_2984 & ~n_8661;
assign n_9160 =  x_1504 &  n_8661;
assign n_9161 = ~n_9159 & ~n_9160;
assign n_9162 =  x_2984 & ~n_9161;
assign n_9163 = ~x_2984 &  n_9161;
assign n_9164 = ~n_9162 & ~n_9163;
assign n_9165 =  x_2983 & ~n_8669;
assign n_9166 =  x_1504 &  n_8669;
assign n_9167 = ~n_9165 & ~n_9166;
assign n_9168 =  x_2983 & ~n_9167;
assign n_9169 = ~x_2983 &  n_9167;
assign n_9170 = ~n_9168 & ~n_9169;
assign n_9171 =  x_2982 & ~n_8676;
assign n_9172 =  x_1504 &  n_8676;
assign n_9173 = ~n_9171 & ~n_9172;
assign n_9174 =  x_2982 & ~n_9173;
assign n_9175 = ~x_2982 &  n_9173;
assign n_9176 = ~n_9174 & ~n_9175;
assign n_9177 =  x_2981 & ~n_8684;
assign n_9178 =  x_1504 &  n_8684;
assign n_9179 = ~n_9177 & ~n_9178;
assign n_9180 =  x_2981 & ~n_9179;
assign n_9181 = ~x_2981 &  n_9179;
assign n_9182 = ~n_9180 & ~n_9181;
assign n_9183 =  x_2980 & ~n_8691;
assign n_9184 =  x_1504 &  n_8691;
assign n_9185 = ~n_9183 & ~n_9184;
assign n_9186 =  x_2980 & ~n_9185;
assign n_9187 = ~x_2980 &  n_9185;
assign n_9188 = ~n_9186 & ~n_9187;
assign n_9189 =  x_2979 & ~n_8699;
assign n_9190 =  x_1504 &  n_8699;
assign n_9191 = ~n_9189 & ~n_9190;
assign n_9192 =  x_2979 & ~n_9191;
assign n_9193 = ~x_2979 &  n_9191;
assign n_9194 = ~n_9192 & ~n_9193;
assign n_9195 =  x_2978 & ~n_8706;
assign n_9196 =  x_1504 &  n_8706;
assign n_9197 = ~n_9195 & ~n_9196;
assign n_9198 =  x_2978 & ~n_9197;
assign n_9199 = ~x_2978 &  n_9197;
assign n_9200 = ~n_9198 & ~n_9199;
assign n_9201 =  x_2977 & ~n_8714;
assign n_9202 =  x_1504 &  n_8714;
assign n_9203 = ~n_9201 & ~n_9202;
assign n_9204 =  x_2977 & ~n_9203;
assign n_9205 = ~x_2977 &  n_9203;
assign n_9206 = ~n_9204 & ~n_9205;
assign n_9207 =  x_2976 & ~n_8721;
assign n_9208 =  x_1504 &  n_8721;
assign n_9209 = ~n_9207 & ~n_9208;
assign n_9210 =  x_2976 & ~n_9209;
assign n_9211 = ~x_2976 &  n_9209;
assign n_9212 = ~n_9210 & ~n_9211;
assign n_9213 =  x_2975 & ~n_8729;
assign n_9214 =  x_1504 &  n_8729;
assign n_9215 = ~n_9213 & ~n_9214;
assign n_9216 =  x_2975 & ~n_9215;
assign n_9217 = ~x_2975 &  n_9215;
assign n_9218 = ~n_9216 & ~n_9217;
assign n_9219 =  x_2974 & ~n_8736;
assign n_9220 =  x_1504 &  n_8736;
assign n_9221 = ~n_9219 & ~n_9220;
assign n_9222 =  x_2974 & ~n_9221;
assign n_9223 = ~x_2974 &  n_9221;
assign n_9224 = ~n_9222 & ~n_9223;
assign n_9225 =  x_2973 & ~n_8744;
assign n_9226 =  x_1504 &  n_8744;
assign n_9227 = ~n_9225 & ~n_9226;
assign n_9228 =  x_2973 & ~n_9227;
assign n_9229 = ~x_2973 &  n_9227;
assign n_9230 = ~n_9228 & ~n_9229;
assign n_9231 =  x_2972 & ~n_8629;
assign n_9232 =  x_1505 &  n_8629;
assign n_9233 = ~n_9231 & ~n_9232;
assign n_9234 =  x_2972 & ~n_9233;
assign n_9235 = ~x_2972 &  n_9233;
assign n_9236 = ~n_9234 & ~n_9235;
assign n_9237 =  x_2971 & ~n_8638;
assign n_9238 =  x_1505 &  n_8638;
assign n_9239 = ~n_9237 & ~n_9238;
assign n_9240 =  x_2971 & ~n_9239;
assign n_9241 = ~x_2971 &  n_9239;
assign n_9242 = ~n_9240 & ~n_9241;
assign n_9243 =  x_2970 & ~n_8645;
assign n_9244 =  x_1505 &  n_8645;
assign n_9245 = ~n_9243 & ~n_9244;
assign n_9246 =  x_2970 & ~n_9245;
assign n_9247 = ~x_2970 &  n_9245;
assign n_9248 = ~n_9246 & ~n_9247;
assign n_9249 =  x_2969 & ~n_8654;
assign n_9250 =  x_1505 &  n_8654;
assign n_9251 = ~n_9249 & ~n_9250;
assign n_9252 =  x_2969 & ~n_9251;
assign n_9253 = ~x_2969 &  n_9251;
assign n_9254 = ~n_9252 & ~n_9253;
assign n_9255 =  x_2968 & ~n_8661;
assign n_9256 =  x_1505 &  n_8661;
assign n_9257 = ~n_9255 & ~n_9256;
assign n_9258 =  x_2968 & ~n_9257;
assign n_9259 = ~x_2968 &  n_9257;
assign n_9260 = ~n_9258 & ~n_9259;
assign n_9261 =  x_2967 & ~n_8669;
assign n_9262 =  x_1505 &  n_8669;
assign n_9263 = ~n_9261 & ~n_9262;
assign n_9264 =  x_2967 & ~n_9263;
assign n_9265 = ~x_2967 &  n_9263;
assign n_9266 = ~n_9264 & ~n_9265;
assign n_9267 =  x_2966 & ~n_8676;
assign n_9268 =  x_1505 &  n_8676;
assign n_9269 = ~n_9267 & ~n_9268;
assign n_9270 =  x_2966 & ~n_9269;
assign n_9271 = ~x_2966 &  n_9269;
assign n_9272 = ~n_9270 & ~n_9271;
assign n_9273 =  x_2965 & ~n_8684;
assign n_9274 =  x_1505 &  n_8684;
assign n_9275 = ~n_9273 & ~n_9274;
assign n_9276 =  x_2965 & ~n_9275;
assign n_9277 = ~x_2965 &  n_9275;
assign n_9278 = ~n_9276 & ~n_9277;
assign n_9279 =  x_2964 & ~n_8691;
assign n_9280 =  x_1505 &  n_8691;
assign n_9281 = ~n_9279 & ~n_9280;
assign n_9282 =  x_2964 & ~n_9281;
assign n_9283 = ~x_2964 &  n_9281;
assign n_9284 = ~n_9282 & ~n_9283;
assign n_9285 =  x_2963 & ~n_8699;
assign n_9286 =  x_1505 &  n_8699;
assign n_9287 = ~n_9285 & ~n_9286;
assign n_9288 =  x_2963 & ~n_9287;
assign n_9289 = ~x_2963 &  n_9287;
assign n_9290 = ~n_9288 & ~n_9289;
assign n_9291 =  x_2962 & ~n_8706;
assign n_9292 =  x_1505 &  n_8706;
assign n_9293 = ~n_9291 & ~n_9292;
assign n_9294 =  x_2962 & ~n_9293;
assign n_9295 = ~x_2962 &  n_9293;
assign n_9296 = ~n_9294 & ~n_9295;
assign n_9297 =  x_2961 & ~n_8714;
assign n_9298 =  x_1505 &  n_8714;
assign n_9299 = ~n_9297 & ~n_9298;
assign n_9300 =  x_2961 & ~n_9299;
assign n_9301 = ~x_2961 &  n_9299;
assign n_9302 = ~n_9300 & ~n_9301;
assign n_9303 =  x_2960 & ~n_8721;
assign n_9304 =  x_1505 &  n_8721;
assign n_9305 = ~n_9303 & ~n_9304;
assign n_9306 =  x_2960 & ~n_9305;
assign n_9307 = ~x_2960 &  n_9305;
assign n_9308 = ~n_9306 & ~n_9307;
assign n_9309 =  x_2959 & ~n_8729;
assign n_9310 =  x_1505 &  n_8729;
assign n_9311 = ~n_9309 & ~n_9310;
assign n_9312 =  x_2959 & ~n_9311;
assign n_9313 = ~x_2959 &  n_9311;
assign n_9314 = ~n_9312 & ~n_9313;
assign n_9315 =  x_2958 & ~n_8736;
assign n_9316 =  x_1505 &  n_8736;
assign n_9317 = ~n_9315 & ~n_9316;
assign n_9318 =  x_2958 & ~n_9317;
assign n_9319 = ~x_2958 &  n_9317;
assign n_9320 = ~n_9318 & ~n_9319;
assign n_9321 =  x_2957 & ~n_8744;
assign n_9322 =  x_1505 &  n_8744;
assign n_9323 = ~n_9321 & ~n_9322;
assign n_9324 =  x_2957 & ~n_9323;
assign n_9325 = ~x_2957 &  n_9323;
assign n_9326 = ~n_9324 & ~n_9325;
assign n_9327 =  x_2956 & ~n_8629;
assign n_9328 =  x_1506 &  n_8629;
assign n_9329 = ~n_9327 & ~n_9328;
assign n_9330 =  x_2956 & ~n_9329;
assign n_9331 = ~x_2956 &  n_9329;
assign n_9332 = ~n_9330 & ~n_9331;
assign n_9333 =  x_2955 & ~n_8638;
assign n_9334 =  x_1506 &  n_8638;
assign n_9335 = ~n_9333 & ~n_9334;
assign n_9336 =  x_2955 & ~n_9335;
assign n_9337 = ~x_2955 &  n_9335;
assign n_9338 = ~n_9336 & ~n_9337;
assign n_9339 =  x_2954 & ~n_8645;
assign n_9340 =  x_1506 &  n_8645;
assign n_9341 = ~n_9339 & ~n_9340;
assign n_9342 =  x_2954 & ~n_9341;
assign n_9343 = ~x_2954 &  n_9341;
assign n_9344 = ~n_9342 & ~n_9343;
assign n_9345 =  x_2953 & ~n_8654;
assign n_9346 =  x_1506 &  n_8654;
assign n_9347 = ~n_9345 & ~n_9346;
assign n_9348 =  x_2953 & ~n_9347;
assign n_9349 = ~x_2953 &  n_9347;
assign n_9350 = ~n_9348 & ~n_9349;
assign n_9351 =  x_2952 & ~n_8661;
assign n_9352 =  x_1506 &  n_8661;
assign n_9353 = ~n_9351 & ~n_9352;
assign n_9354 =  x_2952 & ~n_9353;
assign n_9355 = ~x_2952 &  n_9353;
assign n_9356 = ~n_9354 & ~n_9355;
assign n_9357 =  x_2951 & ~n_8669;
assign n_9358 =  x_1506 &  n_8669;
assign n_9359 = ~n_9357 & ~n_9358;
assign n_9360 =  x_2951 & ~n_9359;
assign n_9361 = ~x_2951 &  n_9359;
assign n_9362 = ~n_9360 & ~n_9361;
assign n_9363 =  x_2950 & ~n_8676;
assign n_9364 =  x_1506 &  n_8676;
assign n_9365 = ~n_9363 & ~n_9364;
assign n_9366 =  x_2950 & ~n_9365;
assign n_9367 = ~x_2950 &  n_9365;
assign n_9368 = ~n_9366 & ~n_9367;
assign n_9369 =  x_2949 & ~n_8684;
assign n_9370 =  x_1506 &  n_8684;
assign n_9371 = ~n_9369 & ~n_9370;
assign n_9372 =  x_2949 & ~n_9371;
assign n_9373 = ~x_2949 &  n_9371;
assign n_9374 = ~n_9372 & ~n_9373;
assign n_9375 =  x_2948 & ~n_8691;
assign n_9376 =  x_1506 &  n_8691;
assign n_9377 = ~n_9375 & ~n_9376;
assign n_9378 =  x_2948 & ~n_9377;
assign n_9379 = ~x_2948 &  n_9377;
assign n_9380 = ~n_9378 & ~n_9379;
assign n_9381 =  x_2947 & ~n_8699;
assign n_9382 =  x_1506 &  n_8699;
assign n_9383 = ~n_9381 & ~n_9382;
assign n_9384 =  x_2947 & ~n_9383;
assign n_9385 = ~x_2947 &  n_9383;
assign n_9386 = ~n_9384 & ~n_9385;
assign n_9387 =  x_2946 & ~n_8706;
assign n_9388 =  x_1506 &  n_8706;
assign n_9389 = ~n_9387 & ~n_9388;
assign n_9390 =  x_2946 & ~n_9389;
assign n_9391 = ~x_2946 &  n_9389;
assign n_9392 = ~n_9390 & ~n_9391;
assign n_9393 =  x_2945 & ~n_8714;
assign n_9394 =  x_1506 &  n_8714;
assign n_9395 = ~n_9393 & ~n_9394;
assign n_9396 =  x_2945 & ~n_9395;
assign n_9397 = ~x_2945 &  n_9395;
assign n_9398 = ~n_9396 & ~n_9397;
assign n_9399 =  x_2944 & ~n_8721;
assign n_9400 =  x_1506 &  n_8721;
assign n_9401 = ~n_9399 & ~n_9400;
assign n_9402 =  x_2944 & ~n_9401;
assign n_9403 = ~x_2944 &  n_9401;
assign n_9404 = ~n_9402 & ~n_9403;
assign n_9405 =  x_2943 & ~n_8729;
assign n_9406 =  x_1506 &  n_8729;
assign n_9407 = ~n_9405 & ~n_9406;
assign n_9408 =  x_2943 & ~n_9407;
assign n_9409 = ~x_2943 &  n_9407;
assign n_9410 = ~n_9408 & ~n_9409;
assign n_9411 =  x_2942 & ~n_8736;
assign n_9412 =  x_1506 &  n_8736;
assign n_9413 = ~n_9411 & ~n_9412;
assign n_9414 =  x_2942 & ~n_9413;
assign n_9415 = ~x_2942 &  n_9413;
assign n_9416 = ~n_9414 & ~n_9415;
assign n_9417 =  x_2941 & ~n_8744;
assign n_9418 =  x_1506 &  n_8744;
assign n_9419 = ~n_9417 & ~n_9418;
assign n_9420 =  x_2941 & ~n_9419;
assign n_9421 = ~x_2941 &  n_9419;
assign n_9422 = ~n_9420 & ~n_9421;
assign n_9423 =  x_2940 & ~n_8629;
assign n_9424 =  x_1507 &  n_8629;
assign n_9425 = ~n_9423 & ~n_9424;
assign n_9426 =  x_2940 & ~n_9425;
assign n_9427 = ~x_2940 &  n_9425;
assign n_9428 = ~n_9426 & ~n_9427;
assign n_9429 =  x_2939 & ~n_8638;
assign n_9430 =  x_1507 &  n_8638;
assign n_9431 = ~n_9429 & ~n_9430;
assign n_9432 =  x_2939 & ~n_9431;
assign n_9433 = ~x_2939 &  n_9431;
assign n_9434 = ~n_9432 & ~n_9433;
assign n_9435 =  x_2938 & ~n_8645;
assign n_9436 =  x_1507 &  n_8645;
assign n_9437 = ~n_9435 & ~n_9436;
assign n_9438 =  x_2938 & ~n_9437;
assign n_9439 = ~x_2938 &  n_9437;
assign n_9440 = ~n_9438 & ~n_9439;
assign n_9441 =  x_2937 & ~n_8654;
assign n_9442 =  x_1507 &  n_8654;
assign n_9443 = ~n_9441 & ~n_9442;
assign n_9444 =  x_2937 & ~n_9443;
assign n_9445 = ~x_2937 &  n_9443;
assign n_9446 = ~n_9444 & ~n_9445;
assign n_9447 =  x_2936 & ~n_8661;
assign n_9448 =  x_1507 &  n_8661;
assign n_9449 = ~n_9447 & ~n_9448;
assign n_9450 =  x_2936 & ~n_9449;
assign n_9451 = ~x_2936 &  n_9449;
assign n_9452 = ~n_9450 & ~n_9451;
assign n_9453 =  x_2935 & ~n_8669;
assign n_9454 =  x_1507 &  n_8669;
assign n_9455 = ~n_9453 & ~n_9454;
assign n_9456 =  x_2935 & ~n_9455;
assign n_9457 = ~x_2935 &  n_9455;
assign n_9458 = ~n_9456 & ~n_9457;
assign n_9459 =  x_2934 & ~n_8676;
assign n_9460 =  x_1507 &  n_8676;
assign n_9461 = ~n_9459 & ~n_9460;
assign n_9462 =  x_2934 & ~n_9461;
assign n_9463 = ~x_2934 &  n_9461;
assign n_9464 = ~n_9462 & ~n_9463;
assign n_9465 =  x_2933 & ~n_8684;
assign n_9466 =  x_1507 &  n_8684;
assign n_9467 = ~n_9465 & ~n_9466;
assign n_9468 =  x_2933 & ~n_9467;
assign n_9469 = ~x_2933 &  n_9467;
assign n_9470 = ~n_9468 & ~n_9469;
assign n_9471 =  x_2932 & ~n_8691;
assign n_9472 =  x_1507 &  n_8691;
assign n_9473 = ~n_9471 & ~n_9472;
assign n_9474 =  x_2932 & ~n_9473;
assign n_9475 = ~x_2932 &  n_9473;
assign n_9476 = ~n_9474 & ~n_9475;
assign n_9477 =  x_2931 & ~n_8699;
assign n_9478 =  x_1507 &  n_8699;
assign n_9479 = ~n_9477 & ~n_9478;
assign n_9480 =  x_2931 & ~n_9479;
assign n_9481 = ~x_2931 &  n_9479;
assign n_9482 = ~n_9480 & ~n_9481;
assign n_9483 =  x_2930 & ~n_8706;
assign n_9484 =  x_1507 &  n_8706;
assign n_9485 = ~n_9483 & ~n_9484;
assign n_9486 =  x_2930 & ~n_9485;
assign n_9487 = ~x_2930 &  n_9485;
assign n_9488 = ~n_9486 & ~n_9487;
assign n_9489 =  x_2929 & ~n_8714;
assign n_9490 =  x_1507 &  n_8714;
assign n_9491 = ~n_9489 & ~n_9490;
assign n_9492 =  x_2929 & ~n_9491;
assign n_9493 = ~x_2929 &  n_9491;
assign n_9494 = ~n_9492 & ~n_9493;
assign n_9495 =  x_2928 & ~n_8721;
assign n_9496 =  x_1507 &  n_8721;
assign n_9497 = ~n_9495 & ~n_9496;
assign n_9498 =  x_2928 & ~n_9497;
assign n_9499 = ~x_2928 &  n_9497;
assign n_9500 = ~n_9498 & ~n_9499;
assign n_9501 =  x_2927 & ~n_8729;
assign n_9502 =  x_1507 &  n_8729;
assign n_9503 = ~n_9501 & ~n_9502;
assign n_9504 =  x_2927 & ~n_9503;
assign n_9505 = ~x_2927 &  n_9503;
assign n_9506 = ~n_9504 & ~n_9505;
assign n_9507 =  x_2926 & ~n_8736;
assign n_9508 =  x_1507 &  n_8736;
assign n_9509 = ~n_9507 & ~n_9508;
assign n_9510 =  x_2926 & ~n_9509;
assign n_9511 = ~x_2926 &  n_9509;
assign n_9512 = ~n_9510 & ~n_9511;
assign n_9513 =  x_2925 & ~n_8744;
assign n_9514 =  x_1507 &  n_8744;
assign n_9515 = ~n_9513 & ~n_9514;
assign n_9516 =  x_2925 & ~n_9515;
assign n_9517 = ~x_2925 &  n_9515;
assign n_9518 = ~n_9516 & ~n_9517;
assign n_9519 =  x_2924 & ~n_8629;
assign n_9520 =  x_1508 &  n_8629;
assign n_9521 = ~n_9519 & ~n_9520;
assign n_9522 =  x_2924 & ~n_9521;
assign n_9523 = ~x_2924 &  n_9521;
assign n_9524 = ~n_9522 & ~n_9523;
assign n_9525 =  x_2923 & ~n_8638;
assign n_9526 =  x_1508 &  n_8638;
assign n_9527 = ~n_9525 & ~n_9526;
assign n_9528 =  x_2923 & ~n_9527;
assign n_9529 = ~x_2923 &  n_9527;
assign n_9530 = ~n_9528 & ~n_9529;
assign n_9531 =  x_2922 & ~n_8645;
assign n_9532 =  x_1508 &  n_8645;
assign n_9533 = ~n_9531 & ~n_9532;
assign n_9534 =  x_2922 & ~n_9533;
assign n_9535 = ~x_2922 &  n_9533;
assign n_9536 = ~n_9534 & ~n_9535;
assign n_9537 =  x_2921 & ~n_8654;
assign n_9538 =  x_1508 &  n_8654;
assign n_9539 = ~n_9537 & ~n_9538;
assign n_9540 =  x_2921 & ~n_9539;
assign n_9541 = ~x_2921 &  n_9539;
assign n_9542 = ~n_9540 & ~n_9541;
assign n_9543 =  x_2920 & ~n_8661;
assign n_9544 =  x_1508 &  n_8661;
assign n_9545 = ~n_9543 & ~n_9544;
assign n_9546 =  x_2920 & ~n_9545;
assign n_9547 = ~x_2920 &  n_9545;
assign n_9548 = ~n_9546 & ~n_9547;
assign n_9549 =  x_2919 & ~n_8669;
assign n_9550 =  x_1508 &  n_8669;
assign n_9551 = ~n_9549 & ~n_9550;
assign n_9552 =  x_2919 & ~n_9551;
assign n_9553 = ~x_2919 &  n_9551;
assign n_9554 = ~n_9552 & ~n_9553;
assign n_9555 =  x_2918 & ~n_8676;
assign n_9556 =  x_1508 &  n_8676;
assign n_9557 = ~n_9555 & ~n_9556;
assign n_9558 =  x_2918 & ~n_9557;
assign n_9559 = ~x_2918 &  n_9557;
assign n_9560 = ~n_9558 & ~n_9559;
assign n_9561 =  x_2917 & ~n_8684;
assign n_9562 =  x_1508 &  n_8684;
assign n_9563 = ~n_9561 & ~n_9562;
assign n_9564 =  x_2917 & ~n_9563;
assign n_9565 = ~x_2917 &  n_9563;
assign n_9566 = ~n_9564 & ~n_9565;
assign n_9567 =  x_2916 & ~n_8691;
assign n_9568 =  x_1508 &  n_8691;
assign n_9569 = ~n_9567 & ~n_9568;
assign n_9570 =  x_2916 & ~n_9569;
assign n_9571 = ~x_2916 &  n_9569;
assign n_9572 = ~n_9570 & ~n_9571;
assign n_9573 =  x_2915 & ~n_8699;
assign n_9574 =  x_1508 &  n_8699;
assign n_9575 = ~n_9573 & ~n_9574;
assign n_9576 =  x_2915 & ~n_9575;
assign n_9577 = ~x_2915 &  n_9575;
assign n_9578 = ~n_9576 & ~n_9577;
assign n_9579 =  x_2914 & ~n_8706;
assign n_9580 =  x_1508 &  n_8706;
assign n_9581 = ~n_9579 & ~n_9580;
assign n_9582 =  x_2914 & ~n_9581;
assign n_9583 = ~x_2914 &  n_9581;
assign n_9584 = ~n_9582 & ~n_9583;
assign n_9585 =  x_2913 & ~n_8714;
assign n_9586 =  x_1508 &  n_8714;
assign n_9587 = ~n_9585 & ~n_9586;
assign n_9588 =  x_2913 & ~n_9587;
assign n_9589 = ~x_2913 &  n_9587;
assign n_9590 = ~n_9588 & ~n_9589;
assign n_9591 =  x_2912 & ~n_8721;
assign n_9592 =  x_1508 &  n_8721;
assign n_9593 = ~n_9591 & ~n_9592;
assign n_9594 =  x_2912 & ~n_9593;
assign n_9595 = ~x_2912 &  n_9593;
assign n_9596 = ~n_9594 & ~n_9595;
assign n_9597 =  x_2911 & ~n_8729;
assign n_9598 =  x_1508 &  n_8729;
assign n_9599 = ~n_9597 & ~n_9598;
assign n_9600 =  x_2911 & ~n_9599;
assign n_9601 = ~x_2911 &  n_9599;
assign n_9602 = ~n_9600 & ~n_9601;
assign n_9603 =  x_2910 & ~n_8736;
assign n_9604 =  x_1508 &  n_8736;
assign n_9605 = ~n_9603 & ~n_9604;
assign n_9606 =  x_2910 & ~n_9605;
assign n_9607 = ~x_2910 &  n_9605;
assign n_9608 = ~n_9606 & ~n_9607;
assign n_9609 =  x_2909 & ~n_8744;
assign n_9610 =  x_1508 &  n_8744;
assign n_9611 = ~n_9609 & ~n_9610;
assign n_9612 =  x_2909 & ~n_9611;
assign n_9613 = ~x_2909 &  n_9611;
assign n_9614 = ~n_9612 & ~n_9613;
assign n_9615 =  x_2908 & ~n_8629;
assign n_9616 =  x_1509 &  n_8629;
assign n_9617 = ~n_9615 & ~n_9616;
assign n_9618 =  x_2908 & ~n_9617;
assign n_9619 = ~x_2908 &  n_9617;
assign n_9620 = ~n_9618 & ~n_9619;
assign n_9621 =  x_2907 & ~n_8638;
assign n_9622 =  x_1509 &  n_8638;
assign n_9623 = ~n_9621 & ~n_9622;
assign n_9624 =  x_2907 & ~n_9623;
assign n_9625 = ~x_2907 &  n_9623;
assign n_9626 = ~n_9624 & ~n_9625;
assign n_9627 =  x_2906 & ~n_8645;
assign n_9628 =  x_1509 &  n_8645;
assign n_9629 = ~n_9627 & ~n_9628;
assign n_9630 =  x_2906 & ~n_9629;
assign n_9631 = ~x_2906 &  n_9629;
assign n_9632 = ~n_9630 & ~n_9631;
assign n_9633 =  x_2905 & ~n_8654;
assign n_9634 =  x_1509 &  n_8654;
assign n_9635 = ~n_9633 & ~n_9634;
assign n_9636 =  x_2905 & ~n_9635;
assign n_9637 = ~x_2905 &  n_9635;
assign n_9638 = ~n_9636 & ~n_9637;
assign n_9639 =  x_2904 & ~n_8661;
assign n_9640 =  x_1509 &  n_8661;
assign n_9641 = ~n_9639 & ~n_9640;
assign n_9642 =  x_2904 & ~n_9641;
assign n_9643 = ~x_2904 &  n_9641;
assign n_9644 = ~n_9642 & ~n_9643;
assign n_9645 =  x_2903 & ~n_8669;
assign n_9646 =  x_1509 &  n_8669;
assign n_9647 = ~n_9645 & ~n_9646;
assign n_9648 =  x_2903 & ~n_9647;
assign n_9649 = ~x_2903 &  n_9647;
assign n_9650 = ~n_9648 & ~n_9649;
assign n_9651 =  x_2902 & ~n_8676;
assign n_9652 =  x_1509 &  n_8676;
assign n_9653 = ~n_9651 & ~n_9652;
assign n_9654 =  x_2902 & ~n_9653;
assign n_9655 = ~x_2902 &  n_9653;
assign n_9656 = ~n_9654 & ~n_9655;
assign n_9657 =  x_2901 & ~n_8684;
assign n_9658 =  x_1509 &  n_8684;
assign n_9659 = ~n_9657 & ~n_9658;
assign n_9660 =  x_2901 & ~n_9659;
assign n_9661 = ~x_2901 &  n_9659;
assign n_9662 = ~n_9660 & ~n_9661;
assign n_9663 =  x_2900 & ~n_8691;
assign n_9664 =  x_1509 &  n_8691;
assign n_9665 = ~n_9663 & ~n_9664;
assign n_9666 =  x_2900 & ~n_9665;
assign n_9667 = ~x_2900 &  n_9665;
assign n_9668 = ~n_9666 & ~n_9667;
assign n_9669 =  x_2899 & ~n_8699;
assign n_9670 =  x_1509 &  n_8699;
assign n_9671 = ~n_9669 & ~n_9670;
assign n_9672 =  x_2899 & ~n_9671;
assign n_9673 = ~x_2899 &  n_9671;
assign n_9674 = ~n_9672 & ~n_9673;
assign n_9675 =  x_2898 & ~n_8706;
assign n_9676 =  x_1509 &  n_8706;
assign n_9677 = ~n_9675 & ~n_9676;
assign n_9678 =  x_2898 & ~n_9677;
assign n_9679 = ~x_2898 &  n_9677;
assign n_9680 = ~n_9678 & ~n_9679;
assign n_9681 =  x_2897 & ~n_8714;
assign n_9682 =  x_1509 &  n_8714;
assign n_9683 = ~n_9681 & ~n_9682;
assign n_9684 =  x_2897 & ~n_9683;
assign n_9685 = ~x_2897 &  n_9683;
assign n_9686 = ~n_9684 & ~n_9685;
assign n_9687 =  x_2896 & ~n_8721;
assign n_9688 =  x_1509 &  n_8721;
assign n_9689 = ~n_9687 & ~n_9688;
assign n_9690 =  x_2896 & ~n_9689;
assign n_9691 = ~x_2896 &  n_9689;
assign n_9692 = ~n_9690 & ~n_9691;
assign n_9693 =  x_2895 & ~n_8729;
assign n_9694 =  x_1509 &  n_8729;
assign n_9695 = ~n_9693 & ~n_9694;
assign n_9696 =  x_2895 & ~n_9695;
assign n_9697 = ~x_2895 &  n_9695;
assign n_9698 = ~n_9696 & ~n_9697;
assign n_9699 =  x_2894 & ~n_8736;
assign n_9700 =  x_1509 &  n_8736;
assign n_9701 = ~n_9699 & ~n_9700;
assign n_9702 =  x_2894 & ~n_9701;
assign n_9703 = ~x_2894 &  n_9701;
assign n_9704 = ~n_9702 & ~n_9703;
assign n_9705 =  x_2893 & ~n_8744;
assign n_9706 =  x_1509 &  n_8744;
assign n_9707 = ~n_9705 & ~n_9706;
assign n_9708 =  x_2893 & ~n_9707;
assign n_9709 = ~x_2893 &  n_9707;
assign n_9710 = ~n_9708 & ~n_9709;
assign n_9711 =  x_2892 & ~n_8629;
assign n_9712 =  x_1510 &  n_8629;
assign n_9713 = ~n_9711 & ~n_9712;
assign n_9714 =  x_2892 & ~n_9713;
assign n_9715 = ~x_2892 &  n_9713;
assign n_9716 = ~n_9714 & ~n_9715;
assign n_9717 =  x_2891 & ~n_8638;
assign n_9718 =  x_1510 &  n_8638;
assign n_9719 = ~n_9717 & ~n_9718;
assign n_9720 =  x_2891 & ~n_9719;
assign n_9721 = ~x_2891 &  n_9719;
assign n_9722 = ~n_9720 & ~n_9721;
assign n_9723 =  x_2890 & ~n_8645;
assign n_9724 =  x_1510 &  n_8645;
assign n_9725 = ~n_9723 & ~n_9724;
assign n_9726 =  x_2890 & ~n_9725;
assign n_9727 = ~x_2890 &  n_9725;
assign n_9728 = ~n_9726 & ~n_9727;
assign n_9729 =  x_2889 & ~n_8654;
assign n_9730 =  x_1510 &  n_8654;
assign n_9731 = ~n_9729 & ~n_9730;
assign n_9732 =  x_2889 & ~n_9731;
assign n_9733 = ~x_2889 &  n_9731;
assign n_9734 = ~n_9732 & ~n_9733;
assign n_9735 =  x_2888 & ~n_8661;
assign n_9736 =  x_1510 &  n_8661;
assign n_9737 = ~n_9735 & ~n_9736;
assign n_9738 =  x_2888 & ~n_9737;
assign n_9739 = ~x_2888 &  n_9737;
assign n_9740 = ~n_9738 & ~n_9739;
assign n_9741 =  x_2887 & ~n_8669;
assign n_9742 =  x_1510 &  n_8669;
assign n_9743 = ~n_9741 & ~n_9742;
assign n_9744 =  x_2887 & ~n_9743;
assign n_9745 = ~x_2887 &  n_9743;
assign n_9746 = ~n_9744 & ~n_9745;
assign n_9747 =  x_2886 & ~n_8676;
assign n_9748 =  x_1510 &  n_8676;
assign n_9749 = ~n_9747 & ~n_9748;
assign n_9750 =  x_2886 & ~n_9749;
assign n_9751 = ~x_2886 &  n_9749;
assign n_9752 = ~n_9750 & ~n_9751;
assign n_9753 =  x_2885 & ~n_8684;
assign n_9754 =  x_1510 &  n_8684;
assign n_9755 = ~n_9753 & ~n_9754;
assign n_9756 =  x_2885 & ~n_9755;
assign n_9757 = ~x_2885 &  n_9755;
assign n_9758 = ~n_9756 & ~n_9757;
assign n_9759 =  x_2884 & ~n_8691;
assign n_9760 =  x_1510 &  n_8691;
assign n_9761 = ~n_9759 & ~n_9760;
assign n_9762 =  x_2884 & ~n_9761;
assign n_9763 = ~x_2884 &  n_9761;
assign n_9764 = ~n_9762 & ~n_9763;
assign n_9765 =  x_2883 & ~n_8699;
assign n_9766 =  x_1510 &  n_8699;
assign n_9767 = ~n_9765 & ~n_9766;
assign n_9768 =  x_2883 & ~n_9767;
assign n_9769 = ~x_2883 &  n_9767;
assign n_9770 = ~n_9768 & ~n_9769;
assign n_9771 =  x_2882 & ~n_8706;
assign n_9772 =  x_1510 &  n_8706;
assign n_9773 = ~n_9771 & ~n_9772;
assign n_9774 =  x_2882 & ~n_9773;
assign n_9775 = ~x_2882 &  n_9773;
assign n_9776 = ~n_9774 & ~n_9775;
assign n_9777 =  x_2881 & ~n_8714;
assign n_9778 =  x_1510 &  n_8714;
assign n_9779 = ~n_9777 & ~n_9778;
assign n_9780 =  x_2881 & ~n_9779;
assign n_9781 = ~x_2881 &  n_9779;
assign n_9782 = ~n_9780 & ~n_9781;
assign n_9783 =  x_2880 & ~n_8721;
assign n_9784 =  x_1510 &  n_8721;
assign n_9785 = ~n_9783 & ~n_9784;
assign n_9786 =  x_2880 & ~n_9785;
assign n_9787 = ~x_2880 &  n_9785;
assign n_9788 = ~n_9786 & ~n_9787;
assign n_9789 =  x_2879 & ~n_8729;
assign n_9790 =  x_1510 &  n_8729;
assign n_9791 = ~n_9789 & ~n_9790;
assign n_9792 =  x_2879 & ~n_9791;
assign n_9793 = ~x_2879 &  n_9791;
assign n_9794 = ~n_9792 & ~n_9793;
assign n_9795 =  x_2878 & ~n_8736;
assign n_9796 =  x_1510 &  n_8736;
assign n_9797 = ~n_9795 & ~n_9796;
assign n_9798 =  x_2878 & ~n_9797;
assign n_9799 = ~x_2878 &  n_9797;
assign n_9800 = ~n_9798 & ~n_9799;
assign n_9801 =  x_2877 & ~n_8744;
assign n_9802 =  x_1510 &  n_8744;
assign n_9803 = ~n_9801 & ~n_9802;
assign n_9804 =  x_2877 & ~n_9803;
assign n_9805 = ~x_2877 &  n_9803;
assign n_9806 = ~n_9804 & ~n_9805;
assign n_9807 =  x_2876 & ~n_8629;
assign n_9808 =  x_1511 &  n_8629;
assign n_9809 = ~n_9807 & ~n_9808;
assign n_9810 =  x_2876 & ~n_9809;
assign n_9811 = ~x_2876 &  n_9809;
assign n_9812 = ~n_9810 & ~n_9811;
assign n_9813 =  x_2875 & ~n_8638;
assign n_9814 =  x_1511 &  n_8638;
assign n_9815 = ~n_9813 & ~n_9814;
assign n_9816 =  x_2875 & ~n_9815;
assign n_9817 = ~x_2875 &  n_9815;
assign n_9818 = ~n_9816 & ~n_9817;
assign n_9819 =  x_2874 & ~n_8645;
assign n_9820 =  x_1511 &  n_8645;
assign n_9821 = ~n_9819 & ~n_9820;
assign n_9822 =  x_2874 & ~n_9821;
assign n_9823 = ~x_2874 &  n_9821;
assign n_9824 = ~n_9822 & ~n_9823;
assign n_9825 =  x_2873 & ~n_8654;
assign n_9826 =  x_1511 &  n_8654;
assign n_9827 = ~n_9825 & ~n_9826;
assign n_9828 =  x_2873 & ~n_9827;
assign n_9829 = ~x_2873 &  n_9827;
assign n_9830 = ~n_9828 & ~n_9829;
assign n_9831 =  x_2872 & ~n_8661;
assign n_9832 =  x_1511 &  n_8661;
assign n_9833 = ~n_9831 & ~n_9832;
assign n_9834 =  x_2872 & ~n_9833;
assign n_9835 = ~x_2872 &  n_9833;
assign n_9836 = ~n_9834 & ~n_9835;
assign n_9837 =  x_2871 & ~n_8669;
assign n_9838 =  x_1511 &  n_8669;
assign n_9839 = ~n_9837 & ~n_9838;
assign n_9840 =  x_2871 & ~n_9839;
assign n_9841 = ~x_2871 &  n_9839;
assign n_9842 = ~n_9840 & ~n_9841;
assign n_9843 =  x_2870 & ~n_8676;
assign n_9844 =  x_1511 &  n_8676;
assign n_9845 = ~n_9843 & ~n_9844;
assign n_9846 =  x_2870 & ~n_9845;
assign n_9847 = ~x_2870 &  n_9845;
assign n_9848 = ~n_9846 & ~n_9847;
assign n_9849 =  x_2869 & ~n_8684;
assign n_9850 =  x_1511 &  n_8684;
assign n_9851 = ~n_9849 & ~n_9850;
assign n_9852 =  x_2869 & ~n_9851;
assign n_9853 = ~x_2869 &  n_9851;
assign n_9854 = ~n_9852 & ~n_9853;
assign n_9855 =  x_2868 & ~n_8691;
assign n_9856 =  x_1511 &  n_8691;
assign n_9857 = ~n_9855 & ~n_9856;
assign n_9858 =  x_2868 & ~n_9857;
assign n_9859 = ~x_2868 &  n_9857;
assign n_9860 = ~n_9858 & ~n_9859;
assign n_9861 =  x_2867 & ~n_8699;
assign n_9862 =  x_1511 &  n_8699;
assign n_9863 = ~n_9861 & ~n_9862;
assign n_9864 =  x_2867 & ~n_9863;
assign n_9865 = ~x_2867 &  n_9863;
assign n_9866 = ~n_9864 & ~n_9865;
assign n_9867 =  x_2866 & ~n_8706;
assign n_9868 =  x_1511 &  n_8706;
assign n_9869 = ~n_9867 & ~n_9868;
assign n_9870 =  x_2866 & ~n_9869;
assign n_9871 = ~x_2866 &  n_9869;
assign n_9872 = ~n_9870 & ~n_9871;
assign n_9873 =  x_2865 & ~n_8714;
assign n_9874 =  x_1511 &  n_8714;
assign n_9875 = ~n_9873 & ~n_9874;
assign n_9876 =  x_2865 & ~n_9875;
assign n_9877 = ~x_2865 &  n_9875;
assign n_9878 = ~n_9876 & ~n_9877;
assign n_9879 =  x_2864 & ~n_8721;
assign n_9880 =  x_1511 &  n_8721;
assign n_9881 = ~n_9879 & ~n_9880;
assign n_9882 =  x_2864 & ~n_9881;
assign n_9883 = ~x_2864 &  n_9881;
assign n_9884 = ~n_9882 & ~n_9883;
assign n_9885 =  x_2863 & ~n_8729;
assign n_9886 =  x_1511 &  n_8729;
assign n_9887 = ~n_9885 & ~n_9886;
assign n_9888 =  x_2863 & ~n_9887;
assign n_9889 = ~x_2863 &  n_9887;
assign n_9890 = ~n_9888 & ~n_9889;
assign n_9891 =  x_2862 & ~n_8736;
assign n_9892 =  x_1511 &  n_8736;
assign n_9893 = ~n_9891 & ~n_9892;
assign n_9894 =  x_2862 & ~n_9893;
assign n_9895 = ~x_2862 &  n_9893;
assign n_9896 = ~n_9894 & ~n_9895;
assign n_9897 =  x_2861 & ~n_8744;
assign n_9898 =  x_1511 &  n_8744;
assign n_9899 = ~n_9897 & ~n_9898;
assign n_9900 =  x_2861 & ~n_9899;
assign n_9901 = ~x_2861 &  n_9899;
assign n_9902 = ~n_9900 & ~n_9901;
assign n_9903 =  x_2860 & ~n_8629;
assign n_9904 =  x_1512 &  n_8629;
assign n_9905 = ~n_9903 & ~n_9904;
assign n_9906 =  x_2860 & ~n_9905;
assign n_9907 = ~x_2860 &  n_9905;
assign n_9908 = ~n_9906 & ~n_9907;
assign n_9909 =  x_2859 & ~n_8638;
assign n_9910 =  x_1512 &  n_8638;
assign n_9911 = ~n_9909 & ~n_9910;
assign n_9912 =  x_2859 & ~n_9911;
assign n_9913 = ~x_2859 &  n_9911;
assign n_9914 = ~n_9912 & ~n_9913;
assign n_9915 =  x_2858 & ~n_8645;
assign n_9916 =  x_1512 &  n_8645;
assign n_9917 = ~n_9915 & ~n_9916;
assign n_9918 =  x_2858 & ~n_9917;
assign n_9919 = ~x_2858 &  n_9917;
assign n_9920 = ~n_9918 & ~n_9919;
assign n_9921 =  x_2857 & ~n_8654;
assign n_9922 =  x_1512 &  n_8654;
assign n_9923 = ~n_9921 & ~n_9922;
assign n_9924 =  x_2857 & ~n_9923;
assign n_9925 = ~x_2857 &  n_9923;
assign n_9926 = ~n_9924 & ~n_9925;
assign n_9927 =  x_2856 & ~n_8661;
assign n_9928 =  x_1512 &  n_8661;
assign n_9929 = ~n_9927 & ~n_9928;
assign n_9930 =  x_2856 & ~n_9929;
assign n_9931 = ~x_2856 &  n_9929;
assign n_9932 = ~n_9930 & ~n_9931;
assign n_9933 =  x_2855 & ~n_8669;
assign n_9934 =  x_1512 &  n_8669;
assign n_9935 = ~n_9933 & ~n_9934;
assign n_9936 =  x_2855 & ~n_9935;
assign n_9937 = ~x_2855 &  n_9935;
assign n_9938 = ~n_9936 & ~n_9937;
assign n_9939 =  x_2854 & ~n_8676;
assign n_9940 =  x_1512 &  n_8676;
assign n_9941 = ~n_9939 & ~n_9940;
assign n_9942 =  x_2854 & ~n_9941;
assign n_9943 = ~x_2854 &  n_9941;
assign n_9944 = ~n_9942 & ~n_9943;
assign n_9945 =  x_2853 & ~n_8684;
assign n_9946 =  x_1512 &  n_8684;
assign n_9947 = ~n_9945 & ~n_9946;
assign n_9948 =  x_2853 & ~n_9947;
assign n_9949 = ~x_2853 &  n_9947;
assign n_9950 = ~n_9948 & ~n_9949;
assign n_9951 =  x_2852 & ~n_8691;
assign n_9952 =  x_1512 &  n_8691;
assign n_9953 = ~n_9951 & ~n_9952;
assign n_9954 =  x_2852 & ~n_9953;
assign n_9955 = ~x_2852 &  n_9953;
assign n_9956 = ~n_9954 & ~n_9955;
assign n_9957 =  x_2851 & ~n_8699;
assign n_9958 =  x_1512 &  n_8699;
assign n_9959 = ~n_9957 & ~n_9958;
assign n_9960 =  x_2851 & ~n_9959;
assign n_9961 = ~x_2851 &  n_9959;
assign n_9962 = ~n_9960 & ~n_9961;
assign n_9963 =  x_2850 & ~n_8706;
assign n_9964 =  x_1512 &  n_8706;
assign n_9965 = ~n_9963 & ~n_9964;
assign n_9966 =  x_2850 & ~n_9965;
assign n_9967 = ~x_2850 &  n_9965;
assign n_9968 = ~n_9966 & ~n_9967;
assign n_9969 =  x_2849 & ~n_8714;
assign n_9970 =  x_1512 &  n_8714;
assign n_9971 = ~n_9969 & ~n_9970;
assign n_9972 =  x_2849 & ~n_9971;
assign n_9973 = ~x_2849 &  n_9971;
assign n_9974 = ~n_9972 & ~n_9973;
assign n_9975 =  x_2848 & ~n_8721;
assign n_9976 =  x_1512 &  n_8721;
assign n_9977 = ~n_9975 & ~n_9976;
assign n_9978 =  x_2848 & ~n_9977;
assign n_9979 = ~x_2848 &  n_9977;
assign n_9980 = ~n_9978 & ~n_9979;
assign n_9981 =  x_2847 & ~n_8729;
assign n_9982 =  x_1512 &  n_8729;
assign n_9983 = ~n_9981 & ~n_9982;
assign n_9984 =  x_2847 & ~n_9983;
assign n_9985 = ~x_2847 &  n_9983;
assign n_9986 = ~n_9984 & ~n_9985;
assign n_9987 =  x_2846 & ~n_8736;
assign n_9988 =  x_1512 &  n_8736;
assign n_9989 = ~n_9987 & ~n_9988;
assign n_9990 =  x_2846 & ~n_9989;
assign n_9991 = ~x_2846 &  n_9989;
assign n_9992 = ~n_9990 & ~n_9991;
assign n_9993 =  x_2845 & ~n_8744;
assign n_9994 =  x_1512 &  n_8744;
assign n_9995 = ~n_9993 & ~n_9994;
assign n_9996 =  x_2845 & ~n_9995;
assign n_9997 = ~x_2845 &  n_9995;
assign n_9998 = ~n_9996 & ~n_9997;
assign n_9999 =  x_2844 & ~n_8629;
assign n_10000 =  x_1513 &  n_8629;
assign n_10001 = ~n_9999 & ~n_10000;
assign n_10002 =  x_2844 & ~n_10001;
assign n_10003 = ~x_2844 &  n_10001;
assign n_10004 = ~n_10002 & ~n_10003;
assign n_10005 =  x_2843 & ~n_8638;
assign n_10006 =  x_1513 &  n_8638;
assign n_10007 = ~n_10005 & ~n_10006;
assign n_10008 =  x_2843 & ~n_10007;
assign n_10009 = ~x_2843 &  n_10007;
assign n_10010 = ~n_10008 & ~n_10009;
assign n_10011 =  x_2842 & ~n_8645;
assign n_10012 =  x_1513 &  n_8645;
assign n_10013 = ~n_10011 & ~n_10012;
assign n_10014 =  x_2842 & ~n_10013;
assign n_10015 = ~x_2842 &  n_10013;
assign n_10016 = ~n_10014 & ~n_10015;
assign n_10017 =  x_2841 & ~n_8654;
assign n_10018 =  x_1513 &  n_8654;
assign n_10019 = ~n_10017 & ~n_10018;
assign n_10020 =  x_2841 & ~n_10019;
assign n_10021 = ~x_2841 &  n_10019;
assign n_10022 = ~n_10020 & ~n_10021;
assign n_10023 =  x_2840 & ~n_8661;
assign n_10024 =  x_1513 &  n_8661;
assign n_10025 = ~n_10023 & ~n_10024;
assign n_10026 =  x_2840 & ~n_10025;
assign n_10027 = ~x_2840 &  n_10025;
assign n_10028 = ~n_10026 & ~n_10027;
assign n_10029 =  x_2839 & ~n_8669;
assign n_10030 =  x_1513 &  n_8669;
assign n_10031 = ~n_10029 & ~n_10030;
assign n_10032 =  x_2839 & ~n_10031;
assign n_10033 = ~x_2839 &  n_10031;
assign n_10034 = ~n_10032 & ~n_10033;
assign n_10035 =  x_2838 & ~n_8676;
assign n_10036 =  x_1513 &  n_8676;
assign n_10037 = ~n_10035 & ~n_10036;
assign n_10038 =  x_2838 & ~n_10037;
assign n_10039 = ~x_2838 &  n_10037;
assign n_10040 = ~n_10038 & ~n_10039;
assign n_10041 =  x_2837 & ~n_8684;
assign n_10042 =  x_1513 &  n_8684;
assign n_10043 = ~n_10041 & ~n_10042;
assign n_10044 =  x_2837 & ~n_10043;
assign n_10045 = ~x_2837 &  n_10043;
assign n_10046 = ~n_10044 & ~n_10045;
assign n_10047 =  x_2836 & ~n_8691;
assign n_10048 =  x_1513 &  n_8691;
assign n_10049 = ~n_10047 & ~n_10048;
assign n_10050 =  x_2836 & ~n_10049;
assign n_10051 = ~x_2836 &  n_10049;
assign n_10052 = ~n_10050 & ~n_10051;
assign n_10053 =  x_2835 & ~n_8699;
assign n_10054 =  x_1513 &  n_8699;
assign n_10055 = ~n_10053 & ~n_10054;
assign n_10056 =  x_2835 & ~n_10055;
assign n_10057 = ~x_2835 &  n_10055;
assign n_10058 = ~n_10056 & ~n_10057;
assign n_10059 =  x_2834 & ~n_8706;
assign n_10060 =  x_1513 &  n_8706;
assign n_10061 = ~n_10059 & ~n_10060;
assign n_10062 =  x_2834 & ~n_10061;
assign n_10063 = ~x_2834 &  n_10061;
assign n_10064 = ~n_10062 & ~n_10063;
assign n_10065 =  x_2833 & ~n_8714;
assign n_10066 =  x_1513 &  n_8714;
assign n_10067 = ~n_10065 & ~n_10066;
assign n_10068 =  x_2833 & ~n_10067;
assign n_10069 = ~x_2833 &  n_10067;
assign n_10070 = ~n_10068 & ~n_10069;
assign n_10071 =  x_2832 & ~n_8721;
assign n_10072 =  x_1513 &  n_8721;
assign n_10073 = ~n_10071 & ~n_10072;
assign n_10074 =  x_2832 & ~n_10073;
assign n_10075 = ~x_2832 &  n_10073;
assign n_10076 = ~n_10074 & ~n_10075;
assign n_10077 =  x_2831 & ~n_8729;
assign n_10078 =  x_1513 &  n_8729;
assign n_10079 = ~n_10077 & ~n_10078;
assign n_10080 =  x_2831 & ~n_10079;
assign n_10081 = ~x_2831 &  n_10079;
assign n_10082 = ~n_10080 & ~n_10081;
assign n_10083 =  x_2830 & ~n_8736;
assign n_10084 =  x_1513 &  n_8736;
assign n_10085 = ~n_10083 & ~n_10084;
assign n_10086 =  x_2830 & ~n_10085;
assign n_10087 = ~x_2830 &  n_10085;
assign n_10088 = ~n_10086 & ~n_10087;
assign n_10089 =  x_2829 & ~n_8744;
assign n_10090 =  x_1513 &  n_8744;
assign n_10091 = ~n_10089 & ~n_10090;
assign n_10092 =  x_2829 & ~n_10091;
assign n_10093 = ~x_2829 &  n_10091;
assign n_10094 = ~n_10092 & ~n_10093;
assign n_10095 =  x_2828 & ~n_8629;
assign n_10096 =  x_1514 &  n_8629;
assign n_10097 = ~n_10095 & ~n_10096;
assign n_10098 =  x_2828 & ~n_10097;
assign n_10099 = ~x_2828 &  n_10097;
assign n_10100 = ~n_10098 & ~n_10099;
assign n_10101 =  x_2827 & ~n_8638;
assign n_10102 =  x_1514 &  n_8638;
assign n_10103 = ~n_10101 & ~n_10102;
assign n_10104 =  x_2827 & ~n_10103;
assign n_10105 = ~x_2827 &  n_10103;
assign n_10106 = ~n_10104 & ~n_10105;
assign n_10107 =  x_2826 & ~n_8645;
assign n_10108 =  x_1514 &  n_8645;
assign n_10109 = ~n_10107 & ~n_10108;
assign n_10110 =  x_2826 & ~n_10109;
assign n_10111 = ~x_2826 &  n_10109;
assign n_10112 = ~n_10110 & ~n_10111;
assign n_10113 =  x_2825 & ~n_8654;
assign n_10114 =  x_1514 &  n_8654;
assign n_10115 = ~n_10113 & ~n_10114;
assign n_10116 =  x_2825 & ~n_10115;
assign n_10117 = ~x_2825 &  n_10115;
assign n_10118 = ~n_10116 & ~n_10117;
assign n_10119 =  x_2824 & ~n_8661;
assign n_10120 =  x_1514 &  n_8661;
assign n_10121 = ~n_10119 & ~n_10120;
assign n_10122 =  x_2824 & ~n_10121;
assign n_10123 = ~x_2824 &  n_10121;
assign n_10124 = ~n_10122 & ~n_10123;
assign n_10125 =  x_2823 & ~n_8669;
assign n_10126 =  x_1514 &  n_8669;
assign n_10127 = ~n_10125 & ~n_10126;
assign n_10128 =  x_2823 & ~n_10127;
assign n_10129 = ~x_2823 &  n_10127;
assign n_10130 = ~n_10128 & ~n_10129;
assign n_10131 =  x_2822 & ~n_8676;
assign n_10132 =  x_1514 &  n_8676;
assign n_10133 = ~n_10131 & ~n_10132;
assign n_10134 =  x_2822 & ~n_10133;
assign n_10135 = ~x_2822 &  n_10133;
assign n_10136 = ~n_10134 & ~n_10135;
assign n_10137 =  x_2821 & ~n_8684;
assign n_10138 =  x_1514 &  n_8684;
assign n_10139 = ~n_10137 & ~n_10138;
assign n_10140 =  x_2821 & ~n_10139;
assign n_10141 = ~x_2821 &  n_10139;
assign n_10142 = ~n_10140 & ~n_10141;
assign n_10143 =  x_2820 & ~n_8691;
assign n_10144 =  x_1514 &  n_8691;
assign n_10145 = ~n_10143 & ~n_10144;
assign n_10146 =  x_2820 & ~n_10145;
assign n_10147 = ~x_2820 &  n_10145;
assign n_10148 = ~n_10146 & ~n_10147;
assign n_10149 =  x_2819 & ~n_8699;
assign n_10150 =  x_1514 &  n_8699;
assign n_10151 = ~n_10149 & ~n_10150;
assign n_10152 =  x_2819 & ~n_10151;
assign n_10153 = ~x_2819 &  n_10151;
assign n_10154 = ~n_10152 & ~n_10153;
assign n_10155 =  x_2818 & ~n_8706;
assign n_10156 =  x_1514 &  n_8706;
assign n_10157 = ~n_10155 & ~n_10156;
assign n_10158 =  x_2818 & ~n_10157;
assign n_10159 = ~x_2818 &  n_10157;
assign n_10160 = ~n_10158 & ~n_10159;
assign n_10161 =  x_2817 & ~n_8714;
assign n_10162 =  x_1514 &  n_8714;
assign n_10163 = ~n_10161 & ~n_10162;
assign n_10164 =  x_2817 & ~n_10163;
assign n_10165 = ~x_2817 &  n_10163;
assign n_10166 = ~n_10164 & ~n_10165;
assign n_10167 =  x_2816 & ~n_8721;
assign n_10168 =  x_1514 &  n_8721;
assign n_10169 = ~n_10167 & ~n_10168;
assign n_10170 =  x_2816 & ~n_10169;
assign n_10171 = ~x_2816 &  n_10169;
assign n_10172 = ~n_10170 & ~n_10171;
assign n_10173 =  x_2815 & ~n_8729;
assign n_10174 =  x_1514 &  n_8729;
assign n_10175 = ~n_10173 & ~n_10174;
assign n_10176 =  x_2815 & ~n_10175;
assign n_10177 = ~x_2815 &  n_10175;
assign n_10178 = ~n_10176 & ~n_10177;
assign n_10179 =  x_2814 & ~n_8736;
assign n_10180 =  x_1514 &  n_8736;
assign n_10181 = ~n_10179 & ~n_10180;
assign n_10182 =  x_2814 & ~n_10181;
assign n_10183 = ~x_2814 &  n_10181;
assign n_10184 = ~n_10182 & ~n_10183;
assign n_10185 =  x_2813 & ~n_8744;
assign n_10186 =  x_1514 &  n_8744;
assign n_10187 = ~n_10185 & ~n_10186;
assign n_10188 =  x_2813 & ~n_10187;
assign n_10189 = ~x_2813 &  n_10187;
assign n_10190 = ~n_10188 & ~n_10189;
assign n_10191 =  x_2812 & ~n_8629;
assign n_10192 =  x_1515 &  n_8629;
assign n_10193 = ~n_10191 & ~n_10192;
assign n_10194 =  x_2812 & ~n_10193;
assign n_10195 = ~x_2812 &  n_10193;
assign n_10196 = ~n_10194 & ~n_10195;
assign n_10197 =  x_2811 & ~n_8638;
assign n_10198 =  x_1515 &  n_8638;
assign n_10199 = ~n_10197 & ~n_10198;
assign n_10200 =  x_2811 & ~n_10199;
assign n_10201 = ~x_2811 &  n_10199;
assign n_10202 = ~n_10200 & ~n_10201;
assign n_10203 =  x_2810 & ~n_8645;
assign n_10204 =  x_1515 &  n_8645;
assign n_10205 = ~n_10203 & ~n_10204;
assign n_10206 =  x_2810 & ~n_10205;
assign n_10207 = ~x_2810 &  n_10205;
assign n_10208 = ~n_10206 & ~n_10207;
assign n_10209 =  x_2809 & ~n_8654;
assign n_10210 =  x_1515 &  n_8654;
assign n_10211 = ~n_10209 & ~n_10210;
assign n_10212 =  x_2809 & ~n_10211;
assign n_10213 = ~x_2809 &  n_10211;
assign n_10214 = ~n_10212 & ~n_10213;
assign n_10215 =  x_2808 & ~n_8661;
assign n_10216 =  x_1515 &  n_8661;
assign n_10217 = ~n_10215 & ~n_10216;
assign n_10218 =  x_2808 & ~n_10217;
assign n_10219 = ~x_2808 &  n_10217;
assign n_10220 = ~n_10218 & ~n_10219;
assign n_10221 =  x_2807 & ~n_8669;
assign n_10222 =  x_1515 &  n_8669;
assign n_10223 = ~n_10221 & ~n_10222;
assign n_10224 =  x_2807 & ~n_10223;
assign n_10225 = ~x_2807 &  n_10223;
assign n_10226 = ~n_10224 & ~n_10225;
assign n_10227 =  x_2806 & ~n_8676;
assign n_10228 =  x_1515 &  n_8676;
assign n_10229 = ~n_10227 & ~n_10228;
assign n_10230 =  x_2806 & ~n_10229;
assign n_10231 = ~x_2806 &  n_10229;
assign n_10232 = ~n_10230 & ~n_10231;
assign n_10233 =  x_2805 & ~n_8684;
assign n_10234 =  x_1515 &  n_8684;
assign n_10235 = ~n_10233 & ~n_10234;
assign n_10236 =  x_2805 & ~n_10235;
assign n_10237 = ~x_2805 &  n_10235;
assign n_10238 = ~n_10236 & ~n_10237;
assign n_10239 =  x_2804 & ~n_8691;
assign n_10240 =  x_1515 &  n_8691;
assign n_10241 = ~n_10239 & ~n_10240;
assign n_10242 =  x_2804 & ~n_10241;
assign n_10243 = ~x_2804 &  n_10241;
assign n_10244 = ~n_10242 & ~n_10243;
assign n_10245 =  x_2803 & ~n_8699;
assign n_10246 =  x_1515 &  n_8699;
assign n_10247 = ~n_10245 & ~n_10246;
assign n_10248 =  x_2803 & ~n_10247;
assign n_10249 = ~x_2803 &  n_10247;
assign n_10250 = ~n_10248 & ~n_10249;
assign n_10251 =  x_2802 & ~n_8706;
assign n_10252 =  x_1515 &  n_8706;
assign n_10253 = ~n_10251 & ~n_10252;
assign n_10254 =  x_2802 & ~n_10253;
assign n_10255 = ~x_2802 &  n_10253;
assign n_10256 = ~n_10254 & ~n_10255;
assign n_10257 =  x_2801 & ~n_8714;
assign n_10258 =  x_1515 &  n_8714;
assign n_10259 = ~n_10257 & ~n_10258;
assign n_10260 =  x_2801 & ~n_10259;
assign n_10261 = ~x_2801 &  n_10259;
assign n_10262 = ~n_10260 & ~n_10261;
assign n_10263 =  x_2800 & ~n_8721;
assign n_10264 =  x_1515 &  n_8721;
assign n_10265 = ~n_10263 & ~n_10264;
assign n_10266 =  x_2800 & ~n_10265;
assign n_10267 = ~x_2800 &  n_10265;
assign n_10268 = ~n_10266 & ~n_10267;
assign n_10269 =  x_2799 & ~n_8729;
assign n_10270 =  x_1515 &  n_8729;
assign n_10271 = ~n_10269 & ~n_10270;
assign n_10272 =  x_2799 & ~n_10271;
assign n_10273 = ~x_2799 &  n_10271;
assign n_10274 = ~n_10272 & ~n_10273;
assign n_10275 =  x_2798 & ~n_8736;
assign n_10276 =  x_1515 &  n_8736;
assign n_10277 = ~n_10275 & ~n_10276;
assign n_10278 =  x_2798 & ~n_10277;
assign n_10279 = ~x_2798 &  n_10277;
assign n_10280 = ~n_10278 & ~n_10279;
assign n_10281 =  x_2797 & ~n_8744;
assign n_10282 =  x_1515 &  n_8744;
assign n_10283 = ~n_10281 & ~n_10282;
assign n_10284 =  x_2797 & ~n_10283;
assign n_10285 = ~x_2797 &  n_10283;
assign n_10286 = ~n_10284 & ~n_10285;
assign n_10287 =  x_2796 & ~n_8629;
assign n_10288 =  x_1516 &  n_8629;
assign n_10289 = ~n_10287 & ~n_10288;
assign n_10290 =  x_2796 & ~n_10289;
assign n_10291 = ~x_2796 &  n_10289;
assign n_10292 = ~n_10290 & ~n_10291;
assign n_10293 =  x_2795 & ~n_8638;
assign n_10294 =  x_1516 &  n_8638;
assign n_10295 = ~n_10293 & ~n_10294;
assign n_10296 =  x_2795 & ~n_10295;
assign n_10297 = ~x_2795 &  n_10295;
assign n_10298 = ~n_10296 & ~n_10297;
assign n_10299 =  x_2794 & ~n_8645;
assign n_10300 =  x_1516 &  n_8645;
assign n_10301 = ~n_10299 & ~n_10300;
assign n_10302 =  x_2794 & ~n_10301;
assign n_10303 = ~x_2794 &  n_10301;
assign n_10304 = ~n_10302 & ~n_10303;
assign n_10305 =  x_2793 & ~n_8654;
assign n_10306 =  x_1516 &  n_8654;
assign n_10307 = ~n_10305 & ~n_10306;
assign n_10308 =  x_2793 & ~n_10307;
assign n_10309 = ~x_2793 &  n_10307;
assign n_10310 = ~n_10308 & ~n_10309;
assign n_10311 =  x_2792 & ~n_8661;
assign n_10312 =  x_1516 &  n_8661;
assign n_10313 = ~n_10311 & ~n_10312;
assign n_10314 =  x_2792 & ~n_10313;
assign n_10315 = ~x_2792 &  n_10313;
assign n_10316 = ~n_10314 & ~n_10315;
assign n_10317 =  x_2791 & ~n_8669;
assign n_10318 =  x_1516 &  n_8669;
assign n_10319 = ~n_10317 & ~n_10318;
assign n_10320 =  x_2791 & ~n_10319;
assign n_10321 = ~x_2791 &  n_10319;
assign n_10322 = ~n_10320 & ~n_10321;
assign n_10323 =  x_2790 & ~n_8676;
assign n_10324 =  x_1516 &  n_8676;
assign n_10325 = ~n_10323 & ~n_10324;
assign n_10326 =  x_2790 & ~n_10325;
assign n_10327 = ~x_2790 &  n_10325;
assign n_10328 = ~n_10326 & ~n_10327;
assign n_10329 =  x_2789 & ~n_8684;
assign n_10330 =  x_1516 &  n_8684;
assign n_10331 = ~n_10329 & ~n_10330;
assign n_10332 =  x_2789 & ~n_10331;
assign n_10333 = ~x_2789 &  n_10331;
assign n_10334 = ~n_10332 & ~n_10333;
assign n_10335 =  x_2788 & ~n_8691;
assign n_10336 =  x_1516 &  n_8691;
assign n_10337 = ~n_10335 & ~n_10336;
assign n_10338 =  x_2788 & ~n_10337;
assign n_10339 = ~x_2788 &  n_10337;
assign n_10340 = ~n_10338 & ~n_10339;
assign n_10341 =  x_2787 & ~n_8699;
assign n_10342 =  x_1516 &  n_8699;
assign n_10343 = ~n_10341 & ~n_10342;
assign n_10344 =  x_2787 & ~n_10343;
assign n_10345 = ~x_2787 &  n_10343;
assign n_10346 = ~n_10344 & ~n_10345;
assign n_10347 =  x_2786 & ~n_8706;
assign n_10348 =  x_1516 &  n_8706;
assign n_10349 = ~n_10347 & ~n_10348;
assign n_10350 =  x_2786 & ~n_10349;
assign n_10351 = ~x_2786 &  n_10349;
assign n_10352 = ~n_10350 & ~n_10351;
assign n_10353 =  x_2785 & ~n_8714;
assign n_10354 =  x_1516 &  n_8714;
assign n_10355 = ~n_10353 & ~n_10354;
assign n_10356 =  x_2785 & ~n_10355;
assign n_10357 = ~x_2785 &  n_10355;
assign n_10358 = ~n_10356 & ~n_10357;
assign n_10359 =  x_2784 & ~n_8721;
assign n_10360 =  x_1516 &  n_8721;
assign n_10361 = ~n_10359 & ~n_10360;
assign n_10362 =  x_2784 & ~n_10361;
assign n_10363 = ~x_2784 &  n_10361;
assign n_10364 = ~n_10362 & ~n_10363;
assign n_10365 =  x_2783 & ~n_8729;
assign n_10366 =  x_1516 &  n_8729;
assign n_10367 = ~n_10365 & ~n_10366;
assign n_10368 =  x_2783 & ~n_10367;
assign n_10369 = ~x_2783 &  n_10367;
assign n_10370 = ~n_10368 & ~n_10369;
assign n_10371 =  x_2782 & ~n_8736;
assign n_10372 =  x_1516 &  n_8736;
assign n_10373 = ~n_10371 & ~n_10372;
assign n_10374 =  x_2782 & ~n_10373;
assign n_10375 = ~x_2782 &  n_10373;
assign n_10376 = ~n_10374 & ~n_10375;
assign n_10377 =  x_2781 & ~n_8744;
assign n_10378 =  x_1516 &  n_8744;
assign n_10379 = ~n_10377 & ~n_10378;
assign n_10380 =  x_2781 & ~n_10379;
assign n_10381 = ~x_2781 &  n_10379;
assign n_10382 = ~n_10380 & ~n_10381;
assign n_10383 =  x_2780 & ~n_8629;
assign n_10384 =  x_1517 &  n_8629;
assign n_10385 = ~n_10383 & ~n_10384;
assign n_10386 =  x_2780 & ~n_10385;
assign n_10387 = ~x_2780 &  n_10385;
assign n_10388 = ~n_10386 & ~n_10387;
assign n_10389 =  x_2779 & ~n_8638;
assign n_10390 =  x_1517 &  n_8638;
assign n_10391 = ~n_10389 & ~n_10390;
assign n_10392 =  x_2779 & ~n_10391;
assign n_10393 = ~x_2779 &  n_10391;
assign n_10394 = ~n_10392 & ~n_10393;
assign n_10395 =  x_2778 & ~n_8645;
assign n_10396 =  x_1517 &  n_8645;
assign n_10397 = ~n_10395 & ~n_10396;
assign n_10398 =  x_2778 & ~n_10397;
assign n_10399 = ~x_2778 &  n_10397;
assign n_10400 = ~n_10398 & ~n_10399;
assign n_10401 =  x_2777 & ~n_8654;
assign n_10402 =  x_1517 &  n_8654;
assign n_10403 = ~n_10401 & ~n_10402;
assign n_10404 =  x_2777 & ~n_10403;
assign n_10405 = ~x_2777 &  n_10403;
assign n_10406 = ~n_10404 & ~n_10405;
assign n_10407 =  x_2776 & ~n_8661;
assign n_10408 =  x_1517 &  n_8661;
assign n_10409 = ~n_10407 & ~n_10408;
assign n_10410 =  x_2776 & ~n_10409;
assign n_10411 = ~x_2776 &  n_10409;
assign n_10412 = ~n_10410 & ~n_10411;
assign n_10413 =  x_2775 & ~n_8669;
assign n_10414 =  x_1517 &  n_8669;
assign n_10415 = ~n_10413 & ~n_10414;
assign n_10416 =  x_2775 & ~n_10415;
assign n_10417 = ~x_2775 &  n_10415;
assign n_10418 = ~n_10416 & ~n_10417;
assign n_10419 =  x_2774 & ~n_8676;
assign n_10420 =  x_1517 &  n_8676;
assign n_10421 = ~n_10419 & ~n_10420;
assign n_10422 =  x_2774 & ~n_10421;
assign n_10423 = ~x_2774 &  n_10421;
assign n_10424 = ~n_10422 & ~n_10423;
assign n_10425 =  x_2773 & ~n_8684;
assign n_10426 =  x_1517 &  n_8684;
assign n_10427 = ~n_10425 & ~n_10426;
assign n_10428 =  x_2773 & ~n_10427;
assign n_10429 = ~x_2773 &  n_10427;
assign n_10430 = ~n_10428 & ~n_10429;
assign n_10431 =  x_2772 & ~n_8691;
assign n_10432 =  x_1517 &  n_8691;
assign n_10433 = ~n_10431 & ~n_10432;
assign n_10434 =  x_2772 & ~n_10433;
assign n_10435 = ~x_2772 &  n_10433;
assign n_10436 = ~n_10434 & ~n_10435;
assign n_10437 =  x_2771 & ~n_8699;
assign n_10438 =  x_1517 &  n_8699;
assign n_10439 = ~n_10437 & ~n_10438;
assign n_10440 =  x_2771 & ~n_10439;
assign n_10441 = ~x_2771 &  n_10439;
assign n_10442 = ~n_10440 & ~n_10441;
assign n_10443 =  x_2770 & ~n_8706;
assign n_10444 =  x_1517 &  n_8706;
assign n_10445 = ~n_10443 & ~n_10444;
assign n_10446 =  x_2770 & ~n_10445;
assign n_10447 = ~x_2770 &  n_10445;
assign n_10448 = ~n_10446 & ~n_10447;
assign n_10449 =  x_2769 & ~n_8714;
assign n_10450 =  x_1517 &  n_8714;
assign n_10451 = ~n_10449 & ~n_10450;
assign n_10452 =  x_2769 & ~n_10451;
assign n_10453 = ~x_2769 &  n_10451;
assign n_10454 = ~n_10452 & ~n_10453;
assign n_10455 =  x_2768 & ~n_8721;
assign n_10456 =  x_1517 &  n_8721;
assign n_10457 = ~n_10455 & ~n_10456;
assign n_10458 =  x_2768 & ~n_10457;
assign n_10459 = ~x_2768 &  n_10457;
assign n_10460 = ~n_10458 & ~n_10459;
assign n_10461 =  x_2767 & ~n_8729;
assign n_10462 =  x_1517 &  n_8729;
assign n_10463 = ~n_10461 & ~n_10462;
assign n_10464 =  x_2767 & ~n_10463;
assign n_10465 = ~x_2767 &  n_10463;
assign n_10466 = ~n_10464 & ~n_10465;
assign n_10467 =  x_2766 & ~n_8736;
assign n_10468 =  x_1517 &  n_8736;
assign n_10469 = ~n_10467 & ~n_10468;
assign n_10470 =  x_2766 & ~n_10469;
assign n_10471 = ~x_2766 &  n_10469;
assign n_10472 = ~n_10470 & ~n_10471;
assign n_10473 =  x_2765 & ~n_8744;
assign n_10474 =  x_1517 &  n_8744;
assign n_10475 = ~n_10473 & ~n_10474;
assign n_10476 =  x_2765 & ~n_10475;
assign n_10477 = ~x_2765 &  n_10475;
assign n_10478 = ~n_10476 & ~n_10477;
assign n_10479 =  x_2764 & ~n_8629;
assign n_10480 =  x_1518 &  n_8629;
assign n_10481 = ~n_10479 & ~n_10480;
assign n_10482 =  x_2764 & ~n_10481;
assign n_10483 = ~x_2764 &  n_10481;
assign n_10484 = ~n_10482 & ~n_10483;
assign n_10485 =  x_2763 & ~n_8638;
assign n_10486 =  x_1518 &  n_8638;
assign n_10487 = ~n_10485 & ~n_10486;
assign n_10488 =  x_2763 & ~n_10487;
assign n_10489 = ~x_2763 &  n_10487;
assign n_10490 = ~n_10488 & ~n_10489;
assign n_10491 =  x_2762 & ~n_8645;
assign n_10492 =  x_1518 &  n_8645;
assign n_10493 = ~n_10491 & ~n_10492;
assign n_10494 =  x_2762 & ~n_10493;
assign n_10495 = ~x_2762 &  n_10493;
assign n_10496 = ~n_10494 & ~n_10495;
assign n_10497 =  x_2761 & ~n_8654;
assign n_10498 =  x_1518 &  n_8654;
assign n_10499 = ~n_10497 & ~n_10498;
assign n_10500 =  x_2761 & ~n_10499;
assign n_10501 = ~x_2761 &  n_10499;
assign n_10502 = ~n_10500 & ~n_10501;
assign n_10503 =  x_2760 & ~n_8661;
assign n_10504 =  x_1518 &  n_8661;
assign n_10505 = ~n_10503 & ~n_10504;
assign n_10506 =  x_2760 & ~n_10505;
assign n_10507 = ~x_2760 &  n_10505;
assign n_10508 = ~n_10506 & ~n_10507;
assign n_10509 =  x_2759 & ~n_8669;
assign n_10510 =  x_1518 &  n_8669;
assign n_10511 = ~n_10509 & ~n_10510;
assign n_10512 =  x_2759 & ~n_10511;
assign n_10513 = ~x_2759 &  n_10511;
assign n_10514 = ~n_10512 & ~n_10513;
assign n_10515 =  x_2758 & ~n_8676;
assign n_10516 =  x_1518 &  n_8676;
assign n_10517 = ~n_10515 & ~n_10516;
assign n_10518 =  x_2758 & ~n_10517;
assign n_10519 = ~x_2758 &  n_10517;
assign n_10520 = ~n_10518 & ~n_10519;
assign n_10521 =  x_2757 & ~n_8684;
assign n_10522 =  x_1518 &  n_8684;
assign n_10523 = ~n_10521 & ~n_10522;
assign n_10524 =  x_2757 & ~n_10523;
assign n_10525 = ~x_2757 &  n_10523;
assign n_10526 = ~n_10524 & ~n_10525;
assign n_10527 =  x_2756 & ~n_8691;
assign n_10528 =  x_1518 &  n_8691;
assign n_10529 = ~n_10527 & ~n_10528;
assign n_10530 =  x_2756 & ~n_10529;
assign n_10531 = ~x_2756 &  n_10529;
assign n_10532 = ~n_10530 & ~n_10531;
assign n_10533 =  x_2755 & ~n_8699;
assign n_10534 =  x_1518 &  n_8699;
assign n_10535 = ~n_10533 & ~n_10534;
assign n_10536 =  x_2755 & ~n_10535;
assign n_10537 = ~x_2755 &  n_10535;
assign n_10538 = ~n_10536 & ~n_10537;
assign n_10539 =  x_2754 & ~n_8706;
assign n_10540 =  x_1518 &  n_8706;
assign n_10541 = ~n_10539 & ~n_10540;
assign n_10542 =  x_2754 & ~n_10541;
assign n_10543 = ~x_2754 &  n_10541;
assign n_10544 = ~n_10542 & ~n_10543;
assign n_10545 =  x_2753 & ~n_8714;
assign n_10546 =  x_1518 &  n_8714;
assign n_10547 = ~n_10545 & ~n_10546;
assign n_10548 =  x_2753 & ~n_10547;
assign n_10549 = ~x_2753 &  n_10547;
assign n_10550 = ~n_10548 & ~n_10549;
assign n_10551 =  x_2752 & ~n_8721;
assign n_10552 =  x_1518 &  n_8721;
assign n_10553 = ~n_10551 & ~n_10552;
assign n_10554 =  x_2752 & ~n_10553;
assign n_10555 = ~x_2752 &  n_10553;
assign n_10556 = ~n_10554 & ~n_10555;
assign n_10557 =  x_2751 & ~n_8729;
assign n_10558 =  x_1518 &  n_8729;
assign n_10559 = ~n_10557 & ~n_10558;
assign n_10560 =  x_2751 & ~n_10559;
assign n_10561 = ~x_2751 &  n_10559;
assign n_10562 = ~n_10560 & ~n_10561;
assign n_10563 =  x_2750 & ~n_8736;
assign n_10564 =  x_1518 &  n_8736;
assign n_10565 = ~n_10563 & ~n_10564;
assign n_10566 =  x_2750 & ~n_10565;
assign n_10567 = ~x_2750 &  n_10565;
assign n_10568 = ~n_10566 & ~n_10567;
assign n_10569 =  x_2749 & ~n_8744;
assign n_10570 =  x_1518 &  n_8744;
assign n_10571 = ~n_10569 & ~n_10570;
assign n_10572 =  x_2749 & ~n_10571;
assign n_10573 = ~x_2749 &  n_10571;
assign n_10574 = ~n_10572 & ~n_10573;
assign n_10575 =  x_2748 & ~n_8629;
assign n_10576 =  x_1519 &  n_8629;
assign n_10577 = ~n_10575 & ~n_10576;
assign n_10578 =  x_2748 & ~n_10577;
assign n_10579 = ~x_2748 &  n_10577;
assign n_10580 = ~n_10578 & ~n_10579;
assign n_10581 =  x_2747 & ~n_8638;
assign n_10582 =  x_1519 &  n_8638;
assign n_10583 = ~n_10581 & ~n_10582;
assign n_10584 =  x_2747 & ~n_10583;
assign n_10585 = ~x_2747 &  n_10583;
assign n_10586 = ~n_10584 & ~n_10585;
assign n_10587 =  x_2746 & ~n_8645;
assign n_10588 =  x_1519 &  n_8645;
assign n_10589 = ~n_10587 & ~n_10588;
assign n_10590 =  x_2746 & ~n_10589;
assign n_10591 = ~x_2746 &  n_10589;
assign n_10592 = ~n_10590 & ~n_10591;
assign n_10593 =  x_2745 & ~n_8654;
assign n_10594 =  x_1519 &  n_8654;
assign n_10595 = ~n_10593 & ~n_10594;
assign n_10596 =  x_2745 & ~n_10595;
assign n_10597 = ~x_2745 &  n_10595;
assign n_10598 = ~n_10596 & ~n_10597;
assign n_10599 =  x_2744 & ~n_8661;
assign n_10600 =  x_1519 &  n_8661;
assign n_10601 = ~n_10599 & ~n_10600;
assign n_10602 =  x_2744 & ~n_10601;
assign n_10603 = ~x_2744 &  n_10601;
assign n_10604 = ~n_10602 & ~n_10603;
assign n_10605 =  x_2743 & ~n_8669;
assign n_10606 =  x_1519 &  n_8669;
assign n_10607 = ~n_10605 & ~n_10606;
assign n_10608 =  x_2743 & ~n_10607;
assign n_10609 = ~x_2743 &  n_10607;
assign n_10610 = ~n_10608 & ~n_10609;
assign n_10611 =  x_2742 & ~n_8676;
assign n_10612 =  x_1519 &  n_8676;
assign n_10613 = ~n_10611 & ~n_10612;
assign n_10614 =  x_2742 & ~n_10613;
assign n_10615 = ~x_2742 &  n_10613;
assign n_10616 = ~n_10614 & ~n_10615;
assign n_10617 =  x_2741 & ~n_8684;
assign n_10618 =  x_1519 &  n_8684;
assign n_10619 = ~n_10617 & ~n_10618;
assign n_10620 =  x_2741 & ~n_10619;
assign n_10621 = ~x_2741 &  n_10619;
assign n_10622 = ~n_10620 & ~n_10621;
assign n_10623 =  x_2740 & ~n_8691;
assign n_10624 =  x_1519 &  n_8691;
assign n_10625 = ~n_10623 & ~n_10624;
assign n_10626 =  x_2740 & ~n_10625;
assign n_10627 = ~x_2740 &  n_10625;
assign n_10628 = ~n_10626 & ~n_10627;
assign n_10629 =  x_2739 & ~n_8699;
assign n_10630 =  x_1519 &  n_8699;
assign n_10631 = ~n_10629 & ~n_10630;
assign n_10632 =  x_2739 & ~n_10631;
assign n_10633 = ~x_2739 &  n_10631;
assign n_10634 = ~n_10632 & ~n_10633;
assign n_10635 =  x_2738 & ~n_8706;
assign n_10636 =  x_1519 &  n_8706;
assign n_10637 = ~n_10635 & ~n_10636;
assign n_10638 =  x_2738 & ~n_10637;
assign n_10639 = ~x_2738 &  n_10637;
assign n_10640 = ~n_10638 & ~n_10639;
assign n_10641 =  x_2737 & ~n_8714;
assign n_10642 =  x_1519 &  n_8714;
assign n_10643 = ~n_10641 & ~n_10642;
assign n_10644 =  x_2737 & ~n_10643;
assign n_10645 = ~x_2737 &  n_10643;
assign n_10646 = ~n_10644 & ~n_10645;
assign n_10647 =  x_2736 & ~n_8721;
assign n_10648 =  x_1519 &  n_8721;
assign n_10649 = ~n_10647 & ~n_10648;
assign n_10650 =  x_2736 & ~n_10649;
assign n_10651 = ~x_2736 &  n_10649;
assign n_10652 = ~n_10650 & ~n_10651;
assign n_10653 =  x_2735 & ~n_8729;
assign n_10654 =  x_1519 &  n_8729;
assign n_10655 = ~n_10653 & ~n_10654;
assign n_10656 =  x_2735 & ~n_10655;
assign n_10657 = ~x_2735 &  n_10655;
assign n_10658 = ~n_10656 & ~n_10657;
assign n_10659 =  x_2734 & ~n_8736;
assign n_10660 =  x_1519 &  n_8736;
assign n_10661 = ~n_10659 & ~n_10660;
assign n_10662 =  x_2734 & ~n_10661;
assign n_10663 = ~x_2734 &  n_10661;
assign n_10664 = ~n_10662 & ~n_10663;
assign n_10665 =  x_2733 & ~n_8744;
assign n_10666 =  x_1519 &  n_8744;
assign n_10667 = ~n_10665 & ~n_10666;
assign n_10668 =  x_2733 & ~n_10667;
assign n_10669 = ~x_2733 &  n_10667;
assign n_10670 = ~n_10668 & ~n_10669;
assign n_10671 =  x_2732 & ~n_8629;
assign n_10672 =  x_1520 &  n_8629;
assign n_10673 = ~n_10671 & ~n_10672;
assign n_10674 =  x_2732 & ~n_10673;
assign n_10675 = ~x_2732 &  n_10673;
assign n_10676 = ~n_10674 & ~n_10675;
assign n_10677 =  x_2731 & ~n_8638;
assign n_10678 =  x_1520 &  n_8638;
assign n_10679 = ~n_10677 & ~n_10678;
assign n_10680 =  x_2731 & ~n_10679;
assign n_10681 = ~x_2731 &  n_10679;
assign n_10682 = ~n_10680 & ~n_10681;
assign n_10683 =  x_2730 & ~n_8645;
assign n_10684 =  x_1520 &  n_8645;
assign n_10685 = ~n_10683 & ~n_10684;
assign n_10686 =  x_2730 & ~n_10685;
assign n_10687 = ~x_2730 &  n_10685;
assign n_10688 = ~n_10686 & ~n_10687;
assign n_10689 =  x_2729 & ~n_8654;
assign n_10690 =  x_1520 &  n_8654;
assign n_10691 = ~n_10689 & ~n_10690;
assign n_10692 =  x_2729 & ~n_10691;
assign n_10693 = ~x_2729 &  n_10691;
assign n_10694 = ~n_10692 & ~n_10693;
assign n_10695 =  x_2728 & ~n_8661;
assign n_10696 =  x_1520 &  n_8661;
assign n_10697 = ~n_10695 & ~n_10696;
assign n_10698 =  x_2728 & ~n_10697;
assign n_10699 = ~x_2728 &  n_10697;
assign n_10700 = ~n_10698 & ~n_10699;
assign n_10701 =  x_2727 & ~n_8669;
assign n_10702 =  x_1520 &  n_8669;
assign n_10703 = ~n_10701 & ~n_10702;
assign n_10704 =  x_2727 & ~n_10703;
assign n_10705 = ~x_2727 &  n_10703;
assign n_10706 = ~n_10704 & ~n_10705;
assign n_10707 =  x_2726 & ~n_8676;
assign n_10708 =  x_1520 &  n_8676;
assign n_10709 = ~n_10707 & ~n_10708;
assign n_10710 =  x_2726 & ~n_10709;
assign n_10711 = ~x_2726 &  n_10709;
assign n_10712 = ~n_10710 & ~n_10711;
assign n_10713 =  x_2725 & ~n_8684;
assign n_10714 =  x_1520 &  n_8684;
assign n_10715 = ~n_10713 & ~n_10714;
assign n_10716 =  x_2725 & ~n_10715;
assign n_10717 = ~x_2725 &  n_10715;
assign n_10718 = ~n_10716 & ~n_10717;
assign n_10719 =  x_2724 & ~n_8691;
assign n_10720 =  x_1520 &  n_8691;
assign n_10721 = ~n_10719 & ~n_10720;
assign n_10722 =  x_2724 & ~n_10721;
assign n_10723 = ~x_2724 &  n_10721;
assign n_10724 = ~n_10722 & ~n_10723;
assign n_10725 =  x_2723 & ~n_8699;
assign n_10726 =  x_1520 &  n_8699;
assign n_10727 = ~n_10725 & ~n_10726;
assign n_10728 =  x_2723 & ~n_10727;
assign n_10729 = ~x_2723 &  n_10727;
assign n_10730 = ~n_10728 & ~n_10729;
assign n_10731 =  x_2722 & ~n_8706;
assign n_10732 =  x_1520 &  n_8706;
assign n_10733 = ~n_10731 & ~n_10732;
assign n_10734 =  x_2722 & ~n_10733;
assign n_10735 = ~x_2722 &  n_10733;
assign n_10736 = ~n_10734 & ~n_10735;
assign n_10737 =  x_2721 & ~n_8714;
assign n_10738 =  x_1520 &  n_8714;
assign n_10739 = ~n_10737 & ~n_10738;
assign n_10740 =  x_2721 & ~n_10739;
assign n_10741 = ~x_2721 &  n_10739;
assign n_10742 = ~n_10740 & ~n_10741;
assign n_10743 =  x_2720 & ~n_8721;
assign n_10744 =  x_1520 &  n_8721;
assign n_10745 = ~n_10743 & ~n_10744;
assign n_10746 =  x_2720 & ~n_10745;
assign n_10747 = ~x_2720 &  n_10745;
assign n_10748 = ~n_10746 & ~n_10747;
assign n_10749 =  x_2719 & ~n_8729;
assign n_10750 =  x_1520 &  n_8729;
assign n_10751 = ~n_10749 & ~n_10750;
assign n_10752 =  x_2719 & ~n_10751;
assign n_10753 = ~x_2719 &  n_10751;
assign n_10754 = ~n_10752 & ~n_10753;
assign n_10755 =  x_2718 & ~n_8736;
assign n_10756 =  x_1520 &  n_8736;
assign n_10757 = ~n_10755 & ~n_10756;
assign n_10758 =  x_2718 & ~n_10757;
assign n_10759 = ~x_2718 &  n_10757;
assign n_10760 = ~n_10758 & ~n_10759;
assign n_10761 =  x_2717 & ~n_8744;
assign n_10762 =  x_1520 &  n_8744;
assign n_10763 = ~n_10761 & ~n_10762;
assign n_10764 =  x_2717 & ~n_10763;
assign n_10765 = ~x_2717 &  n_10763;
assign n_10766 = ~n_10764 & ~n_10765;
assign n_10767 =  x_2716 & ~n_8629;
assign n_10768 =  x_1521 &  n_8629;
assign n_10769 = ~n_10767 & ~n_10768;
assign n_10770 =  x_2716 & ~n_10769;
assign n_10771 = ~x_2716 &  n_10769;
assign n_10772 = ~n_10770 & ~n_10771;
assign n_10773 =  x_2715 & ~n_8638;
assign n_10774 =  x_1521 &  n_8638;
assign n_10775 = ~n_10773 & ~n_10774;
assign n_10776 =  x_2715 & ~n_10775;
assign n_10777 = ~x_2715 &  n_10775;
assign n_10778 = ~n_10776 & ~n_10777;
assign n_10779 =  x_2714 & ~n_8645;
assign n_10780 =  x_1521 &  n_8645;
assign n_10781 = ~n_10779 & ~n_10780;
assign n_10782 =  x_2714 & ~n_10781;
assign n_10783 = ~x_2714 &  n_10781;
assign n_10784 = ~n_10782 & ~n_10783;
assign n_10785 =  x_2713 & ~n_8654;
assign n_10786 =  x_1521 &  n_8654;
assign n_10787 = ~n_10785 & ~n_10786;
assign n_10788 =  x_2713 & ~n_10787;
assign n_10789 = ~x_2713 &  n_10787;
assign n_10790 = ~n_10788 & ~n_10789;
assign n_10791 =  x_2712 & ~n_8661;
assign n_10792 =  x_1521 &  n_8661;
assign n_10793 = ~n_10791 & ~n_10792;
assign n_10794 =  x_2712 & ~n_10793;
assign n_10795 = ~x_2712 &  n_10793;
assign n_10796 = ~n_10794 & ~n_10795;
assign n_10797 =  x_2711 & ~n_8669;
assign n_10798 =  x_1521 &  n_8669;
assign n_10799 = ~n_10797 & ~n_10798;
assign n_10800 =  x_2711 & ~n_10799;
assign n_10801 = ~x_2711 &  n_10799;
assign n_10802 = ~n_10800 & ~n_10801;
assign n_10803 =  x_2710 & ~n_8676;
assign n_10804 =  x_1521 &  n_8676;
assign n_10805 = ~n_10803 & ~n_10804;
assign n_10806 =  x_2710 & ~n_10805;
assign n_10807 = ~x_2710 &  n_10805;
assign n_10808 = ~n_10806 & ~n_10807;
assign n_10809 =  x_2709 & ~n_8684;
assign n_10810 =  x_1521 &  n_8684;
assign n_10811 = ~n_10809 & ~n_10810;
assign n_10812 =  x_2709 & ~n_10811;
assign n_10813 = ~x_2709 &  n_10811;
assign n_10814 = ~n_10812 & ~n_10813;
assign n_10815 =  x_2708 & ~n_8691;
assign n_10816 =  x_1521 &  n_8691;
assign n_10817 = ~n_10815 & ~n_10816;
assign n_10818 =  x_2708 & ~n_10817;
assign n_10819 = ~x_2708 &  n_10817;
assign n_10820 = ~n_10818 & ~n_10819;
assign n_10821 =  x_2707 & ~n_8699;
assign n_10822 =  x_1521 &  n_8699;
assign n_10823 = ~n_10821 & ~n_10822;
assign n_10824 =  x_2707 & ~n_10823;
assign n_10825 = ~x_2707 &  n_10823;
assign n_10826 = ~n_10824 & ~n_10825;
assign n_10827 =  x_2706 & ~n_8706;
assign n_10828 =  x_1521 &  n_8706;
assign n_10829 = ~n_10827 & ~n_10828;
assign n_10830 =  x_2706 & ~n_10829;
assign n_10831 = ~x_2706 &  n_10829;
assign n_10832 = ~n_10830 & ~n_10831;
assign n_10833 =  x_2705 & ~n_8714;
assign n_10834 =  x_1521 &  n_8714;
assign n_10835 = ~n_10833 & ~n_10834;
assign n_10836 =  x_2705 & ~n_10835;
assign n_10837 = ~x_2705 &  n_10835;
assign n_10838 = ~n_10836 & ~n_10837;
assign n_10839 =  x_2704 & ~n_8721;
assign n_10840 =  x_1521 &  n_8721;
assign n_10841 = ~n_10839 & ~n_10840;
assign n_10842 =  x_2704 & ~n_10841;
assign n_10843 = ~x_2704 &  n_10841;
assign n_10844 = ~n_10842 & ~n_10843;
assign n_10845 =  x_2703 & ~n_8729;
assign n_10846 =  x_1521 &  n_8729;
assign n_10847 = ~n_10845 & ~n_10846;
assign n_10848 =  x_2703 & ~n_10847;
assign n_10849 = ~x_2703 &  n_10847;
assign n_10850 = ~n_10848 & ~n_10849;
assign n_10851 =  x_2702 & ~n_8736;
assign n_10852 =  x_1521 &  n_8736;
assign n_10853 = ~n_10851 & ~n_10852;
assign n_10854 =  x_2702 & ~n_10853;
assign n_10855 = ~x_2702 &  n_10853;
assign n_10856 = ~n_10854 & ~n_10855;
assign n_10857 =  x_2701 & ~n_8744;
assign n_10858 =  x_1521 &  n_8744;
assign n_10859 = ~n_10857 & ~n_10858;
assign n_10860 =  x_2701 & ~n_10859;
assign n_10861 = ~x_2701 &  n_10859;
assign n_10862 = ~n_10860 & ~n_10861;
assign n_10863 =  x_2700 & ~n_8629;
assign n_10864 =  x_1522 &  n_8629;
assign n_10865 = ~n_10863 & ~n_10864;
assign n_10866 =  x_2700 & ~n_10865;
assign n_10867 = ~x_2700 &  n_10865;
assign n_10868 = ~n_10866 & ~n_10867;
assign n_10869 =  x_2699 & ~n_8638;
assign n_10870 =  x_1522 &  n_8638;
assign n_10871 = ~n_10869 & ~n_10870;
assign n_10872 =  x_2699 & ~n_10871;
assign n_10873 = ~x_2699 &  n_10871;
assign n_10874 = ~n_10872 & ~n_10873;
assign n_10875 =  x_2698 & ~n_8645;
assign n_10876 =  x_1522 &  n_8645;
assign n_10877 = ~n_10875 & ~n_10876;
assign n_10878 =  x_2698 & ~n_10877;
assign n_10879 = ~x_2698 &  n_10877;
assign n_10880 = ~n_10878 & ~n_10879;
assign n_10881 =  x_2697 & ~n_8654;
assign n_10882 =  x_1522 &  n_8654;
assign n_10883 = ~n_10881 & ~n_10882;
assign n_10884 =  x_2697 & ~n_10883;
assign n_10885 = ~x_2697 &  n_10883;
assign n_10886 = ~n_10884 & ~n_10885;
assign n_10887 =  x_2696 & ~n_8661;
assign n_10888 =  x_1522 &  n_8661;
assign n_10889 = ~n_10887 & ~n_10888;
assign n_10890 =  x_2696 & ~n_10889;
assign n_10891 = ~x_2696 &  n_10889;
assign n_10892 = ~n_10890 & ~n_10891;
assign n_10893 =  x_2695 & ~n_8669;
assign n_10894 =  x_1522 &  n_8669;
assign n_10895 = ~n_10893 & ~n_10894;
assign n_10896 =  x_2695 & ~n_10895;
assign n_10897 = ~x_2695 &  n_10895;
assign n_10898 = ~n_10896 & ~n_10897;
assign n_10899 =  x_2694 & ~n_8676;
assign n_10900 =  x_1522 &  n_8676;
assign n_10901 = ~n_10899 & ~n_10900;
assign n_10902 =  x_2694 & ~n_10901;
assign n_10903 = ~x_2694 &  n_10901;
assign n_10904 = ~n_10902 & ~n_10903;
assign n_10905 =  x_2693 & ~n_8684;
assign n_10906 =  x_1522 &  n_8684;
assign n_10907 = ~n_10905 & ~n_10906;
assign n_10908 =  x_2693 & ~n_10907;
assign n_10909 = ~x_2693 &  n_10907;
assign n_10910 = ~n_10908 & ~n_10909;
assign n_10911 =  x_2692 & ~n_8691;
assign n_10912 =  x_1522 &  n_8691;
assign n_10913 = ~n_10911 & ~n_10912;
assign n_10914 =  x_2692 & ~n_10913;
assign n_10915 = ~x_2692 &  n_10913;
assign n_10916 = ~n_10914 & ~n_10915;
assign n_10917 =  x_2691 & ~n_8699;
assign n_10918 =  x_1522 &  n_8699;
assign n_10919 = ~n_10917 & ~n_10918;
assign n_10920 =  x_2691 & ~n_10919;
assign n_10921 = ~x_2691 &  n_10919;
assign n_10922 = ~n_10920 & ~n_10921;
assign n_10923 =  x_2690 & ~n_8706;
assign n_10924 =  x_1522 &  n_8706;
assign n_10925 = ~n_10923 & ~n_10924;
assign n_10926 =  x_2690 & ~n_10925;
assign n_10927 = ~x_2690 &  n_10925;
assign n_10928 = ~n_10926 & ~n_10927;
assign n_10929 =  x_2689 & ~n_8714;
assign n_10930 =  x_1522 &  n_8714;
assign n_10931 = ~n_10929 & ~n_10930;
assign n_10932 =  x_2689 & ~n_10931;
assign n_10933 = ~x_2689 &  n_10931;
assign n_10934 = ~n_10932 & ~n_10933;
assign n_10935 =  x_2688 & ~n_8721;
assign n_10936 =  x_1522 &  n_8721;
assign n_10937 = ~n_10935 & ~n_10936;
assign n_10938 =  x_2688 & ~n_10937;
assign n_10939 = ~x_2688 &  n_10937;
assign n_10940 = ~n_10938 & ~n_10939;
assign n_10941 =  x_2687 & ~n_8729;
assign n_10942 =  x_1522 &  n_8729;
assign n_10943 = ~n_10941 & ~n_10942;
assign n_10944 =  x_2687 & ~n_10943;
assign n_10945 = ~x_2687 &  n_10943;
assign n_10946 = ~n_10944 & ~n_10945;
assign n_10947 =  x_2686 & ~n_8736;
assign n_10948 =  x_1522 &  n_8736;
assign n_10949 = ~n_10947 & ~n_10948;
assign n_10950 =  x_2686 & ~n_10949;
assign n_10951 = ~x_2686 &  n_10949;
assign n_10952 = ~n_10950 & ~n_10951;
assign n_10953 =  x_2685 & ~n_8744;
assign n_10954 =  x_1522 &  n_8744;
assign n_10955 = ~n_10953 & ~n_10954;
assign n_10956 =  x_2685 & ~n_10955;
assign n_10957 = ~x_2685 &  n_10955;
assign n_10958 = ~n_10956 & ~n_10957;
assign n_10959 =  x_2684 & ~n_8629;
assign n_10960 =  x_1523 &  n_8629;
assign n_10961 = ~n_10959 & ~n_10960;
assign n_10962 =  x_2684 & ~n_10961;
assign n_10963 = ~x_2684 &  n_10961;
assign n_10964 = ~n_10962 & ~n_10963;
assign n_10965 =  x_2683 & ~n_8638;
assign n_10966 =  x_1523 &  n_8638;
assign n_10967 = ~n_10965 & ~n_10966;
assign n_10968 =  x_2683 & ~n_10967;
assign n_10969 = ~x_2683 &  n_10967;
assign n_10970 = ~n_10968 & ~n_10969;
assign n_10971 =  x_2682 & ~n_8645;
assign n_10972 =  x_1523 &  n_8645;
assign n_10973 = ~n_10971 & ~n_10972;
assign n_10974 =  x_2682 & ~n_10973;
assign n_10975 = ~x_2682 &  n_10973;
assign n_10976 = ~n_10974 & ~n_10975;
assign n_10977 =  x_2681 & ~n_8654;
assign n_10978 =  x_1523 &  n_8654;
assign n_10979 = ~n_10977 & ~n_10978;
assign n_10980 =  x_2681 & ~n_10979;
assign n_10981 = ~x_2681 &  n_10979;
assign n_10982 = ~n_10980 & ~n_10981;
assign n_10983 =  x_2680 & ~n_8661;
assign n_10984 =  x_1523 &  n_8661;
assign n_10985 = ~n_10983 & ~n_10984;
assign n_10986 =  x_2680 & ~n_10985;
assign n_10987 = ~x_2680 &  n_10985;
assign n_10988 = ~n_10986 & ~n_10987;
assign n_10989 =  x_2679 & ~n_8669;
assign n_10990 =  x_1523 &  n_8669;
assign n_10991 = ~n_10989 & ~n_10990;
assign n_10992 =  x_2679 & ~n_10991;
assign n_10993 = ~x_2679 &  n_10991;
assign n_10994 = ~n_10992 & ~n_10993;
assign n_10995 =  x_2678 & ~n_8676;
assign n_10996 =  x_1523 &  n_8676;
assign n_10997 = ~n_10995 & ~n_10996;
assign n_10998 =  x_2678 & ~n_10997;
assign n_10999 = ~x_2678 &  n_10997;
assign n_11000 = ~n_10998 & ~n_10999;
assign n_11001 =  x_2677 & ~n_8684;
assign n_11002 =  x_1523 &  n_8684;
assign n_11003 = ~n_11001 & ~n_11002;
assign n_11004 =  x_2677 & ~n_11003;
assign n_11005 = ~x_2677 &  n_11003;
assign n_11006 = ~n_11004 & ~n_11005;
assign n_11007 =  x_2676 & ~n_8691;
assign n_11008 =  x_1523 &  n_8691;
assign n_11009 = ~n_11007 & ~n_11008;
assign n_11010 =  x_2676 & ~n_11009;
assign n_11011 = ~x_2676 &  n_11009;
assign n_11012 = ~n_11010 & ~n_11011;
assign n_11013 =  x_2675 & ~n_8699;
assign n_11014 =  x_1523 &  n_8699;
assign n_11015 = ~n_11013 & ~n_11014;
assign n_11016 =  x_2675 & ~n_11015;
assign n_11017 = ~x_2675 &  n_11015;
assign n_11018 = ~n_11016 & ~n_11017;
assign n_11019 =  x_2674 & ~n_8706;
assign n_11020 =  x_1523 &  n_8706;
assign n_11021 = ~n_11019 & ~n_11020;
assign n_11022 =  x_2674 & ~n_11021;
assign n_11023 = ~x_2674 &  n_11021;
assign n_11024 = ~n_11022 & ~n_11023;
assign n_11025 =  x_2673 & ~n_8714;
assign n_11026 =  x_1523 &  n_8714;
assign n_11027 = ~n_11025 & ~n_11026;
assign n_11028 =  x_2673 & ~n_11027;
assign n_11029 = ~x_2673 &  n_11027;
assign n_11030 = ~n_11028 & ~n_11029;
assign n_11031 =  x_2672 & ~n_8721;
assign n_11032 =  x_1523 &  n_8721;
assign n_11033 = ~n_11031 & ~n_11032;
assign n_11034 =  x_2672 & ~n_11033;
assign n_11035 = ~x_2672 &  n_11033;
assign n_11036 = ~n_11034 & ~n_11035;
assign n_11037 =  x_2671 & ~n_8729;
assign n_11038 =  x_1523 &  n_8729;
assign n_11039 = ~n_11037 & ~n_11038;
assign n_11040 =  x_2671 & ~n_11039;
assign n_11041 = ~x_2671 &  n_11039;
assign n_11042 = ~n_11040 & ~n_11041;
assign n_11043 =  x_2670 & ~n_8736;
assign n_11044 =  x_1523 &  n_8736;
assign n_11045 = ~n_11043 & ~n_11044;
assign n_11046 =  x_2670 & ~n_11045;
assign n_11047 = ~x_2670 &  n_11045;
assign n_11048 = ~n_11046 & ~n_11047;
assign n_11049 =  x_2669 & ~n_8744;
assign n_11050 =  x_1523 &  n_8744;
assign n_11051 = ~n_11049 & ~n_11050;
assign n_11052 =  x_2669 & ~n_11051;
assign n_11053 = ~x_2669 &  n_11051;
assign n_11054 = ~n_11052 & ~n_11053;
assign n_11055 =  x_2668 & ~n_8629;
assign n_11056 =  x_1524 &  n_8629;
assign n_11057 = ~n_11055 & ~n_11056;
assign n_11058 =  x_2668 & ~n_11057;
assign n_11059 = ~x_2668 &  n_11057;
assign n_11060 = ~n_11058 & ~n_11059;
assign n_11061 =  x_2667 & ~n_8638;
assign n_11062 =  x_1524 &  n_8638;
assign n_11063 = ~n_11061 & ~n_11062;
assign n_11064 =  x_2667 & ~n_11063;
assign n_11065 = ~x_2667 &  n_11063;
assign n_11066 = ~n_11064 & ~n_11065;
assign n_11067 =  x_2666 & ~n_8645;
assign n_11068 =  x_1524 &  n_8645;
assign n_11069 = ~n_11067 & ~n_11068;
assign n_11070 =  x_2666 & ~n_11069;
assign n_11071 = ~x_2666 &  n_11069;
assign n_11072 = ~n_11070 & ~n_11071;
assign n_11073 =  x_2665 & ~n_8654;
assign n_11074 =  x_1524 &  n_8654;
assign n_11075 = ~n_11073 & ~n_11074;
assign n_11076 =  x_2665 & ~n_11075;
assign n_11077 = ~x_2665 &  n_11075;
assign n_11078 = ~n_11076 & ~n_11077;
assign n_11079 =  x_2664 & ~n_8661;
assign n_11080 =  x_1524 &  n_8661;
assign n_11081 = ~n_11079 & ~n_11080;
assign n_11082 =  x_2664 & ~n_11081;
assign n_11083 = ~x_2664 &  n_11081;
assign n_11084 = ~n_11082 & ~n_11083;
assign n_11085 =  x_2663 & ~n_8669;
assign n_11086 =  x_1524 &  n_8669;
assign n_11087 = ~n_11085 & ~n_11086;
assign n_11088 =  x_2663 & ~n_11087;
assign n_11089 = ~x_2663 &  n_11087;
assign n_11090 = ~n_11088 & ~n_11089;
assign n_11091 =  x_2662 & ~n_8676;
assign n_11092 =  x_1524 &  n_8676;
assign n_11093 = ~n_11091 & ~n_11092;
assign n_11094 =  x_2662 & ~n_11093;
assign n_11095 = ~x_2662 &  n_11093;
assign n_11096 = ~n_11094 & ~n_11095;
assign n_11097 =  x_2661 & ~n_8684;
assign n_11098 =  x_1524 &  n_8684;
assign n_11099 = ~n_11097 & ~n_11098;
assign n_11100 =  x_2661 & ~n_11099;
assign n_11101 = ~x_2661 &  n_11099;
assign n_11102 = ~n_11100 & ~n_11101;
assign n_11103 =  x_2660 & ~n_8691;
assign n_11104 =  x_1524 &  n_8691;
assign n_11105 = ~n_11103 & ~n_11104;
assign n_11106 =  x_2660 & ~n_11105;
assign n_11107 = ~x_2660 &  n_11105;
assign n_11108 = ~n_11106 & ~n_11107;
assign n_11109 =  x_2659 & ~n_8699;
assign n_11110 =  x_1524 &  n_8699;
assign n_11111 = ~n_11109 & ~n_11110;
assign n_11112 =  x_2659 & ~n_11111;
assign n_11113 = ~x_2659 &  n_11111;
assign n_11114 = ~n_11112 & ~n_11113;
assign n_11115 =  x_2658 & ~n_8706;
assign n_11116 =  x_1524 &  n_8706;
assign n_11117 = ~n_11115 & ~n_11116;
assign n_11118 =  x_2658 & ~n_11117;
assign n_11119 = ~x_2658 &  n_11117;
assign n_11120 = ~n_11118 & ~n_11119;
assign n_11121 =  x_2657 & ~n_8714;
assign n_11122 =  x_1524 &  n_8714;
assign n_11123 = ~n_11121 & ~n_11122;
assign n_11124 =  x_2657 & ~n_11123;
assign n_11125 = ~x_2657 &  n_11123;
assign n_11126 = ~n_11124 & ~n_11125;
assign n_11127 =  x_2656 & ~n_8721;
assign n_11128 =  x_1524 &  n_8721;
assign n_11129 = ~n_11127 & ~n_11128;
assign n_11130 =  x_2656 & ~n_11129;
assign n_11131 = ~x_2656 &  n_11129;
assign n_11132 = ~n_11130 & ~n_11131;
assign n_11133 =  x_2655 & ~n_8729;
assign n_11134 =  x_1524 &  n_8729;
assign n_11135 = ~n_11133 & ~n_11134;
assign n_11136 =  x_2655 & ~n_11135;
assign n_11137 = ~x_2655 &  n_11135;
assign n_11138 = ~n_11136 & ~n_11137;
assign n_11139 =  x_2654 & ~n_8736;
assign n_11140 =  x_1524 &  n_8736;
assign n_11141 = ~n_11139 & ~n_11140;
assign n_11142 =  x_2654 & ~n_11141;
assign n_11143 = ~x_2654 &  n_11141;
assign n_11144 = ~n_11142 & ~n_11143;
assign n_11145 =  x_2653 & ~n_8744;
assign n_11146 =  x_1524 &  n_8744;
assign n_11147 = ~n_11145 & ~n_11146;
assign n_11148 =  x_2653 & ~n_11147;
assign n_11149 = ~x_2653 &  n_11147;
assign n_11150 = ~n_11148 & ~n_11149;
assign n_11151 =  x_2652 & ~n_8629;
assign n_11152 =  x_1525 &  n_8629;
assign n_11153 = ~n_11151 & ~n_11152;
assign n_11154 =  x_2652 & ~n_11153;
assign n_11155 = ~x_2652 &  n_11153;
assign n_11156 = ~n_11154 & ~n_11155;
assign n_11157 =  x_2651 & ~n_8638;
assign n_11158 =  x_1525 &  n_8638;
assign n_11159 = ~n_11157 & ~n_11158;
assign n_11160 =  x_2651 & ~n_11159;
assign n_11161 = ~x_2651 &  n_11159;
assign n_11162 = ~n_11160 & ~n_11161;
assign n_11163 =  x_2650 & ~n_8645;
assign n_11164 =  x_1525 &  n_8645;
assign n_11165 = ~n_11163 & ~n_11164;
assign n_11166 =  x_2650 & ~n_11165;
assign n_11167 = ~x_2650 &  n_11165;
assign n_11168 = ~n_11166 & ~n_11167;
assign n_11169 =  x_2649 & ~n_8654;
assign n_11170 =  x_1525 &  n_8654;
assign n_11171 = ~n_11169 & ~n_11170;
assign n_11172 =  x_2649 & ~n_11171;
assign n_11173 = ~x_2649 &  n_11171;
assign n_11174 = ~n_11172 & ~n_11173;
assign n_11175 =  x_2648 & ~n_8661;
assign n_11176 =  x_1525 &  n_8661;
assign n_11177 = ~n_11175 & ~n_11176;
assign n_11178 =  x_2648 & ~n_11177;
assign n_11179 = ~x_2648 &  n_11177;
assign n_11180 = ~n_11178 & ~n_11179;
assign n_11181 =  x_2647 & ~n_8669;
assign n_11182 =  x_1525 &  n_8669;
assign n_11183 = ~n_11181 & ~n_11182;
assign n_11184 =  x_2647 & ~n_11183;
assign n_11185 = ~x_2647 &  n_11183;
assign n_11186 = ~n_11184 & ~n_11185;
assign n_11187 =  x_2646 & ~n_8676;
assign n_11188 =  x_1525 &  n_8676;
assign n_11189 = ~n_11187 & ~n_11188;
assign n_11190 =  x_2646 & ~n_11189;
assign n_11191 = ~x_2646 &  n_11189;
assign n_11192 = ~n_11190 & ~n_11191;
assign n_11193 =  x_2645 & ~n_8684;
assign n_11194 =  x_1525 &  n_8684;
assign n_11195 = ~n_11193 & ~n_11194;
assign n_11196 =  x_2645 & ~n_11195;
assign n_11197 = ~x_2645 &  n_11195;
assign n_11198 = ~n_11196 & ~n_11197;
assign n_11199 =  x_2644 & ~n_8691;
assign n_11200 =  x_1525 &  n_8691;
assign n_11201 = ~n_11199 & ~n_11200;
assign n_11202 =  x_2644 & ~n_11201;
assign n_11203 = ~x_2644 &  n_11201;
assign n_11204 = ~n_11202 & ~n_11203;
assign n_11205 =  x_2643 & ~n_8699;
assign n_11206 =  x_1525 &  n_8699;
assign n_11207 = ~n_11205 & ~n_11206;
assign n_11208 =  x_2643 & ~n_11207;
assign n_11209 = ~x_2643 &  n_11207;
assign n_11210 = ~n_11208 & ~n_11209;
assign n_11211 =  x_2642 & ~n_8706;
assign n_11212 =  x_1525 &  n_8706;
assign n_11213 = ~n_11211 & ~n_11212;
assign n_11214 =  x_2642 & ~n_11213;
assign n_11215 = ~x_2642 &  n_11213;
assign n_11216 = ~n_11214 & ~n_11215;
assign n_11217 =  x_2641 & ~n_8714;
assign n_11218 =  x_1525 &  n_8714;
assign n_11219 = ~n_11217 & ~n_11218;
assign n_11220 =  x_2641 & ~n_11219;
assign n_11221 = ~x_2641 &  n_11219;
assign n_11222 = ~n_11220 & ~n_11221;
assign n_11223 =  x_2640 & ~n_8721;
assign n_11224 =  x_1525 &  n_8721;
assign n_11225 = ~n_11223 & ~n_11224;
assign n_11226 =  x_2640 & ~n_11225;
assign n_11227 = ~x_2640 &  n_11225;
assign n_11228 = ~n_11226 & ~n_11227;
assign n_11229 =  x_2639 & ~n_8729;
assign n_11230 =  x_1525 &  n_8729;
assign n_11231 = ~n_11229 & ~n_11230;
assign n_11232 =  x_2639 & ~n_11231;
assign n_11233 = ~x_2639 &  n_11231;
assign n_11234 = ~n_11232 & ~n_11233;
assign n_11235 =  x_2638 & ~n_8736;
assign n_11236 =  x_1525 &  n_8736;
assign n_11237 = ~n_11235 & ~n_11236;
assign n_11238 =  x_2638 & ~n_11237;
assign n_11239 = ~x_2638 &  n_11237;
assign n_11240 = ~n_11238 & ~n_11239;
assign n_11241 =  x_2637 & ~n_8744;
assign n_11242 =  x_1525 &  n_8744;
assign n_11243 = ~n_11241 & ~n_11242;
assign n_11244 =  x_2637 & ~n_11243;
assign n_11245 = ~x_2637 &  n_11243;
assign n_11246 = ~n_11244 & ~n_11245;
assign n_11247 =  x_2636 & ~n_8629;
assign n_11248 =  x_1526 &  n_8629;
assign n_11249 = ~n_11247 & ~n_11248;
assign n_11250 =  x_2636 & ~n_11249;
assign n_11251 = ~x_2636 &  n_11249;
assign n_11252 = ~n_11250 & ~n_11251;
assign n_11253 =  x_2635 & ~n_8638;
assign n_11254 =  x_1526 &  n_8638;
assign n_11255 = ~n_11253 & ~n_11254;
assign n_11256 =  x_2635 & ~n_11255;
assign n_11257 = ~x_2635 &  n_11255;
assign n_11258 = ~n_11256 & ~n_11257;
assign n_11259 =  x_2634 & ~n_8645;
assign n_11260 =  x_1526 &  n_8645;
assign n_11261 = ~n_11259 & ~n_11260;
assign n_11262 =  x_2634 & ~n_11261;
assign n_11263 = ~x_2634 &  n_11261;
assign n_11264 = ~n_11262 & ~n_11263;
assign n_11265 =  x_2633 & ~n_8654;
assign n_11266 =  x_1526 &  n_8654;
assign n_11267 = ~n_11265 & ~n_11266;
assign n_11268 =  x_2633 & ~n_11267;
assign n_11269 = ~x_2633 &  n_11267;
assign n_11270 = ~n_11268 & ~n_11269;
assign n_11271 =  x_2632 & ~n_8661;
assign n_11272 =  x_1526 &  n_8661;
assign n_11273 = ~n_11271 & ~n_11272;
assign n_11274 =  x_2632 & ~n_11273;
assign n_11275 = ~x_2632 &  n_11273;
assign n_11276 = ~n_11274 & ~n_11275;
assign n_11277 =  x_2631 & ~n_8669;
assign n_11278 =  x_1526 &  n_8669;
assign n_11279 = ~n_11277 & ~n_11278;
assign n_11280 =  x_2631 & ~n_11279;
assign n_11281 = ~x_2631 &  n_11279;
assign n_11282 = ~n_11280 & ~n_11281;
assign n_11283 =  x_2630 & ~n_8676;
assign n_11284 =  x_1526 &  n_8676;
assign n_11285 = ~n_11283 & ~n_11284;
assign n_11286 =  x_2630 & ~n_11285;
assign n_11287 = ~x_2630 &  n_11285;
assign n_11288 = ~n_11286 & ~n_11287;
assign n_11289 =  x_2629 & ~n_8684;
assign n_11290 =  x_1526 &  n_8684;
assign n_11291 = ~n_11289 & ~n_11290;
assign n_11292 =  x_2629 & ~n_11291;
assign n_11293 = ~x_2629 &  n_11291;
assign n_11294 = ~n_11292 & ~n_11293;
assign n_11295 =  x_2628 & ~n_8691;
assign n_11296 =  x_1526 &  n_8691;
assign n_11297 = ~n_11295 & ~n_11296;
assign n_11298 =  x_2628 & ~n_11297;
assign n_11299 = ~x_2628 &  n_11297;
assign n_11300 = ~n_11298 & ~n_11299;
assign n_11301 =  x_2627 & ~n_8699;
assign n_11302 =  x_1526 &  n_8699;
assign n_11303 = ~n_11301 & ~n_11302;
assign n_11304 =  x_2627 & ~n_11303;
assign n_11305 = ~x_2627 &  n_11303;
assign n_11306 = ~n_11304 & ~n_11305;
assign n_11307 =  x_2626 & ~n_8706;
assign n_11308 =  x_1526 &  n_8706;
assign n_11309 = ~n_11307 & ~n_11308;
assign n_11310 =  x_2626 & ~n_11309;
assign n_11311 = ~x_2626 &  n_11309;
assign n_11312 = ~n_11310 & ~n_11311;
assign n_11313 =  x_2625 & ~n_8714;
assign n_11314 =  x_1526 &  n_8714;
assign n_11315 = ~n_11313 & ~n_11314;
assign n_11316 =  x_2625 & ~n_11315;
assign n_11317 = ~x_2625 &  n_11315;
assign n_11318 = ~n_11316 & ~n_11317;
assign n_11319 =  x_2624 & ~n_8721;
assign n_11320 =  x_1526 &  n_8721;
assign n_11321 = ~n_11319 & ~n_11320;
assign n_11322 =  x_2624 & ~n_11321;
assign n_11323 = ~x_2624 &  n_11321;
assign n_11324 = ~n_11322 & ~n_11323;
assign n_11325 =  x_2623 & ~n_8729;
assign n_11326 =  x_1526 &  n_8729;
assign n_11327 = ~n_11325 & ~n_11326;
assign n_11328 =  x_2623 & ~n_11327;
assign n_11329 = ~x_2623 &  n_11327;
assign n_11330 = ~n_11328 & ~n_11329;
assign n_11331 =  x_2622 & ~n_8736;
assign n_11332 =  x_1526 &  n_8736;
assign n_11333 = ~n_11331 & ~n_11332;
assign n_11334 =  x_2622 & ~n_11333;
assign n_11335 = ~x_2622 &  n_11333;
assign n_11336 = ~n_11334 & ~n_11335;
assign n_11337 =  x_2621 & ~n_8744;
assign n_11338 =  x_1526 &  n_8744;
assign n_11339 = ~n_11337 & ~n_11338;
assign n_11340 =  x_2621 & ~n_11339;
assign n_11341 = ~x_2621 &  n_11339;
assign n_11342 = ~n_11340 & ~n_11341;
assign n_11343 =  x_2620 & ~n_8629;
assign n_11344 =  x_1527 &  n_8629;
assign n_11345 = ~n_11343 & ~n_11344;
assign n_11346 =  x_2620 & ~n_11345;
assign n_11347 = ~x_2620 &  n_11345;
assign n_11348 = ~n_11346 & ~n_11347;
assign n_11349 =  x_2619 & ~n_8638;
assign n_11350 =  x_1527 &  n_8638;
assign n_11351 = ~n_11349 & ~n_11350;
assign n_11352 =  x_2619 & ~n_11351;
assign n_11353 = ~x_2619 &  n_11351;
assign n_11354 = ~n_11352 & ~n_11353;
assign n_11355 =  x_2618 & ~n_8645;
assign n_11356 =  x_1527 &  n_8645;
assign n_11357 = ~n_11355 & ~n_11356;
assign n_11358 =  x_2618 & ~n_11357;
assign n_11359 = ~x_2618 &  n_11357;
assign n_11360 = ~n_11358 & ~n_11359;
assign n_11361 =  x_2617 & ~n_8654;
assign n_11362 =  x_1527 &  n_8654;
assign n_11363 = ~n_11361 & ~n_11362;
assign n_11364 =  x_2617 & ~n_11363;
assign n_11365 = ~x_2617 &  n_11363;
assign n_11366 = ~n_11364 & ~n_11365;
assign n_11367 =  x_2616 & ~n_8661;
assign n_11368 =  x_1527 &  n_8661;
assign n_11369 = ~n_11367 & ~n_11368;
assign n_11370 =  x_2616 & ~n_11369;
assign n_11371 = ~x_2616 &  n_11369;
assign n_11372 = ~n_11370 & ~n_11371;
assign n_11373 =  x_2615 & ~n_8669;
assign n_11374 =  x_1527 &  n_8669;
assign n_11375 = ~n_11373 & ~n_11374;
assign n_11376 =  x_2615 & ~n_11375;
assign n_11377 = ~x_2615 &  n_11375;
assign n_11378 = ~n_11376 & ~n_11377;
assign n_11379 =  x_2614 & ~n_8676;
assign n_11380 =  x_1527 &  n_8676;
assign n_11381 = ~n_11379 & ~n_11380;
assign n_11382 =  x_2614 & ~n_11381;
assign n_11383 = ~x_2614 &  n_11381;
assign n_11384 = ~n_11382 & ~n_11383;
assign n_11385 =  x_2613 & ~n_8684;
assign n_11386 =  x_1527 &  n_8684;
assign n_11387 = ~n_11385 & ~n_11386;
assign n_11388 =  x_2613 & ~n_11387;
assign n_11389 = ~x_2613 &  n_11387;
assign n_11390 = ~n_11388 & ~n_11389;
assign n_11391 =  x_2612 & ~n_8691;
assign n_11392 =  x_1527 &  n_8691;
assign n_11393 = ~n_11391 & ~n_11392;
assign n_11394 =  x_2612 & ~n_11393;
assign n_11395 = ~x_2612 &  n_11393;
assign n_11396 = ~n_11394 & ~n_11395;
assign n_11397 =  x_2611 & ~n_8699;
assign n_11398 =  x_1527 &  n_8699;
assign n_11399 = ~n_11397 & ~n_11398;
assign n_11400 =  x_2611 & ~n_11399;
assign n_11401 = ~x_2611 &  n_11399;
assign n_11402 = ~n_11400 & ~n_11401;
assign n_11403 =  x_2610 & ~n_8706;
assign n_11404 =  x_1527 &  n_8706;
assign n_11405 = ~n_11403 & ~n_11404;
assign n_11406 =  x_2610 & ~n_11405;
assign n_11407 = ~x_2610 &  n_11405;
assign n_11408 = ~n_11406 & ~n_11407;
assign n_11409 =  x_2609 & ~n_8714;
assign n_11410 =  x_1527 &  n_8714;
assign n_11411 = ~n_11409 & ~n_11410;
assign n_11412 =  x_2609 & ~n_11411;
assign n_11413 = ~x_2609 &  n_11411;
assign n_11414 = ~n_11412 & ~n_11413;
assign n_11415 =  x_2608 & ~n_8721;
assign n_11416 =  x_1527 &  n_8721;
assign n_11417 = ~n_11415 & ~n_11416;
assign n_11418 =  x_2608 & ~n_11417;
assign n_11419 = ~x_2608 &  n_11417;
assign n_11420 = ~n_11418 & ~n_11419;
assign n_11421 =  x_2607 & ~n_8729;
assign n_11422 =  x_1527 &  n_8729;
assign n_11423 = ~n_11421 & ~n_11422;
assign n_11424 =  x_2607 & ~n_11423;
assign n_11425 = ~x_2607 &  n_11423;
assign n_11426 = ~n_11424 & ~n_11425;
assign n_11427 =  x_2606 & ~n_8736;
assign n_11428 =  x_1527 &  n_8736;
assign n_11429 = ~n_11427 & ~n_11428;
assign n_11430 =  x_2606 & ~n_11429;
assign n_11431 = ~x_2606 &  n_11429;
assign n_11432 = ~n_11430 & ~n_11431;
assign n_11433 =  x_2605 & ~n_8744;
assign n_11434 =  x_1527 &  n_8744;
assign n_11435 = ~n_11433 & ~n_11434;
assign n_11436 =  x_2605 & ~n_11435;
assign n_11437 = ~x_2605 &  n_11435;
assign n_11438 = ~n_11436 & ~n_11437;
assign n_11439 =  x_2604 & ~n_8629;
assign n_11440 =  x_1528 &  n_8629;
assign n_11441 = ~n_11439 & ~n_11440;
assign n_11442 =  x_2604 & ~n_11441;
assign n_11443 = ~x_2604 &  n_11441;
assign n_11444 = ~n_11442 & ~n_11443;
assign n_11445 =  x_2603 & ~n_8638;
assign n_11446 =  x_1528 &  n_8638;
assign n_11447 = ~n_11445 & ~n_11446;
assign n_11448 =  x_2603 & ~n_11447;
assign n_11449 = ~x_2603 &  n_11447;
assign n_11450 = ~n_11448 & ~n_11449;
assign n_11451 =  x_2602 & ~n_8645;
assign n_11452 =  x_1528 &  n_8645;
assign n_11453 = ~n_11451 & ~n_11452;
assign n_11454 =  x_2602 & ~n_11453;
assign n_11455 = ~x_2602 &  n_11453;
assign n_11456 = ~n_11454 & ~n_11455;
assign n_11457 =  x_2601 & ~n_8654;
assign n_11458 =  x_1528 &  n_8654;
assign n_11459 = ~n_11457 & ~n_11458;
assign n_11460 =  x_2601 & ~n_11459;
assign n_11461 = ~x_2601 &  n_11459;
assign n_11462 = ~n_11460 & ~n_11461;
assign n_11463 =  x_2600 & ~n_8661;
assign n_11464 =  x_1528 &  n_8661;
assign n_11465 = ~n_11463 & ~n_11464;
assign n_11466 =  x_2600 & ~n_11465;
assign n_11467 = ~x_2600 &  n_11465;
assign n_11468 = ~n_11466 & ~n_11467;
assign n_11469 =  x_2599 & ~n_8669;
assign n_11470 =  x_1528 &  n_8669;
assign n_11471 = ~n_11469 & ~n_11470;
assign n_11472 =  x_2599 & ~n_11471;
assign n_11473 = ~x_2599 &  n_11471;
assign n_11474 = ~n_11472 & ~n_11473;
assign n_11475 =  x_2598 & ~n_8676;
assign n_11476 =  x_1528 &  n_8676;
assign n_11477 = ~n_11475 & ~n_11476;
assign n_11478 =  x_2598 & ~n_11477;
assign n_11479 = ~x_2598 &  n_11477;
assign n_11480 = ~n_11478 & ~n_11479;
assign n_11481 =  x_2597 & ~n_8684;
assign n_11482 =  x_1528 &  n_8684;
assign n_11483 = ~n_11481 & ~n_11482;
assign n_11484 =  x_2597 & ~n_11483;
assign n_11485 = ~x_2597 &  n_11483;
assign n_11486 = ~n_11484 & ~n_11485;
assign n_11487 =  x_2596 & ~n_8691;
assign n_11488 =  x_1528 &  n_8691;
assign n_11489 = ~n_11487 & ~n_11488;
assign n_11490 =  x_2596 & ~n_11489;
assign n_11491 = ~x_2596 &  n_11489;
assign n_11492 = ~n_11490 & ~n_11491;
assign n_11493 =  x_2595 & ~n_8699;
assign n_11494 =  x_1528 &  n_8699;
assign n_11495 = ~n_11493 & ~n_11494;
assign n_11496 =  x_2595 & ~n_11495;
assign n_11497 = ~x_2595 &  n_11495;
assign n_11498 = ~n_11496 & ~n_11497;
assign n_11499 =  x_2594 & ~n_8706;
assign n_11500 =  x_1528 &  n_8706;
assign n_11501 = ~n_11499 & ~n_11500;
assign n_11502 =  x_2594 & ~n_11501;
assign n_11503 = ~x_2594 &  n_11501;
assign n_11504 = ~n_11502 & ~n_11503;
assign n_11505 =  x_2593 & ~n_8714;
assign n_11506 =  x_1528 &  n_8714;
assign n_11507 = ~n_11505 & ~n_11506;
assign n_11508 =  x_2593 & ~n_11507;
assign n_11509 = ~x_2593 &  n_11507;
assign n_11510 = ~n_11508 & ~n_11509;
assign n_11511 =  x_2592 & ~n_8721;
assign n_11512 =  x_1528 &  n_8721;
assign n_11513 = ~n_11511 & ~n_11512;
assign n_11514 =  x_2592 & ~n_11513;
assign n_11515 = ~x_2592 &  n_11513;
assign n_11516 = ~n_11514 & ~n_11515;
assign n_11517 =  x_2591 & ~n_8729;
assign n_11518 =  x_1528 &  n_8729;
assign n_11519 = ~n_11517 & ~n_11518;
assign n_11520 =  x_2591 & ~n_11519;
assign n_11521 = ~x_2591 &  n_11519;
assign n_11522 = ~n_11520 & ~n_11521;
assign n_11523 =  x_2590 & ~n_8736;
assign n_11524 =  x_1528 &  n_8736;
assign n_11525 = ~n_11523 & ~n_11524;
assign n_11526 =  x_2590 & ~n_11525;
assign n_11527 = ~x_2590 &  n_11525;
assign n_11528 = ~n_11526 & ~n_11527;
assign n_11529 =  x_2589 & ~n_8744;
assign n_11530 =  x_1528 &  n_8744;
assign n_11531 = ~n_11529 & ~n_11530;
assign n_11532 =  x_2589 & ~n_11531;
assign n_11533 = ~x_2589 &  n_11531;
assign n_11534 = ~n_11532 & ~n_11533;
assign n_11535 =  x_2588 & ~n_8629;
assign n_11536 =  x_1529 &  n_8629;
assign n_11537 = ~n_11535 & ~n_11536;
assign n_11538 =  x_2588 & ~n_11537;
assign n_11539 = ~x_2588 &  n_11537;
assign n_11540 = ~n_11538 & ~n_11539;
assign n_11541 =  x_2587 & ~n_8638;
assign n_11542 =  x_1529 &  n_8638;
assign n_11543 = ~n_11541 & ~n_11542;
assign n_11544 =  x_2587 & ~n_11543;
assign n_11545 = ~x_2587 &  n_11543;
assign n_11546 = ~n_11544 & ~n_11545;
assign n_11547 =  x_2586 & ~n_8645;
assign n_11548 =  x_1529 &  n_8645;
assign n_11549 = ~n_11547 & ~n_11548;
assign n_11550 =  x_2586 & ~n_11549;
assign n_11551 = ~x_2586 &  n_11549;
assign n_11552 = ~n_11550 & ~n_11551;
assign n_11553 =  x_2585 & ~n_8654;
assign n_11554 =  x_1529 &  n_8654;
assign n_11555 = ~n_11553 & ~n_11554;
assign n_11556 =  x_2585 & ~n_11555;
assign n_11557 = ~x_2585 &  n_11555;
assign n_11558 = ~n_11556 & ~n_11557;
assign n_11559 =  x_2584 & ~n_8661;
assign n_11560 =  x_1529 &  n_8661;
assign n_11561 = ~n_11559 & ~n_11560;
assign n_11562 =  x_2584 & ~n_11561;
assign n_11563 = ~x_2584 &  n_11561;
assign n_11564 = ~n_11562 & ~n_11563;
assign n_11565 =  x_2583 & ~n_8669;
assign n_11566 =  x_1529 &  n_8669;
assign n_11567 = ~n_11565 & ~n_11566;
assign n_11568 =  x_2583 & ~n_11567;
assign n_11569 = ~x_2583 &  n_11567;
assign n_11570 = ~n_11568 & ~n_11569;
assign n_11571 =  x_2582 & ~n_8676;
assign n_11572 =  x_1529 &  n_8676;
assign n_11573 = ~n_11571 & ~n_11572;
assign n_11574 =  x_2582 & ~n_11573;
assign n_11575 = ~x_2582 &  n_11573;
assign n_11576 = ~n_11574 & ~n_11575;
assign n_11577 =  x_2581 & ~n_8684;
assign n_11578 =  x_1529 &  n_8684;
assign n_11579 = ~n_11577 & ~n_11578;
assign n_11580 =  x_2581 & ~n_11579;
assign n_11581 = ~x_2581 &  n_11579;
assign n_11582 = ~n_11580 & ~n_11581;
assign n_11583 =  x_2580 & ~n_8691;
assign n_11584 =  x_1529 &  n_8691;
assign n_11585 = ~n_11583 & ~n_11584;
assign n_11586 =  x_2580 & ~n_11585;
assign n_11587 = ~x_2580 &  n_11585;
assign n_11588 = ~n_11586 & ~n_11587;
assign n_11589 =  x_2579 & ~n_8699;
assign n_11590 =  x_1529 &  n_8699;
assign n_11591 = ~n_11589 & ~n_11590;
assign n_11592 =  x_2579 & ~n_11591;
assign n_11593 = ~x_2579 &  n_11591;
assign n_11594 = ~n_11592 & ~n_11593;
assign n_11595 =  x_2578 & ~n_8706;
assign n_11596 =  x_1529 &  n_8706;
assign n_11597 = ~n_11595 & ~n_11596;
assign n_11598 =  x_2578 & ~n_11597;
assign n_11599 = ~x_2578 &  n_11597;
assign n_11600 = ~n_11598 & ~n_11599;
assign n_11601 =  x_2577 & ~n_8714;
assign n_11602 =  x_1529 &  n_8714;
assign n_11603 = ~n_11601 & ~n_11602;
assign n_11604 =  x_2577 & ~n_11603;
assign n_11605 = ~x_2577 &  n_11603;
assign n_11606 = ~n_11604 & ~n_11605;
assign n_11607 =  x_2576 & ~n_8721;
assign n_11608 =  x_1529 &  n_8721;
assign n_11609 = ~n_11607 & ~n_11608;
assign n_11610 =  x_2576 & ~n_11609;
assign n_11611 = ~x_2576 &  n_11609;
assign n_11612 = ~n_11610 & ~n_11611;
assign n_11613 =  x_2575 & ~n_8729;
assign n_11614 =  x_1529 &  n_8729;
assign n_11615 = ~n_11613 & ~n_11614;
assign n_11616 =  x_2575 & ~n_11615;
assign n_11617 = ~x_2575 &  n_11615;
assign n_11618 = ~n_11616 & ~n_11617;
assign n_11619 =  x_2574 & ~n_8736;
assign n_11620 =  x_1529 &  n_8736;
assign n_11621 = ~n_11619 & ~n_11620;
assign n_11622 =  x_2574 & ~n_11621;
assign n_11623 = ~x_2574 &  n_11621;
assign n_11624 = ~n_11622 & ~n_11623;
assign n_11625 =  x_2573 & ~n_8744;
assign n_11626 =  x_1529 &  n_8744;
assign n_11627 = ~n_11625 & ~n_11626;
assign n_11628 =  x_2573 & ~n_11627;
assign n_11629 = ~x_2573 &  n_11627;
assign n_11630 = ~n_11628 & ~n_11629;
assign n_11631 =  x_2572 & ~n_8629;
assign n_11632 =  x_1530 &  n_8629;
assign n_11633 = ~n_11631 & ~n_11632;
assign n_11634 =  x_2572 & ~n_11633;
assign n_11635 = ~x_2572 &  n_11633;
assign n_11636 = ~n_11634 & ~n_11635;
assign n_11637 =  x_2571 & ~n_8638;
assign n_11638 =  x_1530 &  n_8638;
assign n_11639 = ~n_11637 & ~n_11638;
assign n_11640 =  x_2571 & ~n_11639;
assign n_11641 = ~x_2571 &  n_11639;
assign n_11642 = ~n_11640 & ~n_11641;
assign n_11643 =  x_2570 & ~n_8645;
assign n_11644 =  x_1530 &  n_8645;
assign n_11645 = ~n_11643 & ~n_11644;
assign n_11646 =  x_2570 & ~n_11645;
assign n_11647 = ~x_2570 &  n_11645;
assign n_11648 = ~n_11646 & ~n_11647;
assign n_11649 =  x_2569 & ~n_8654;
assign n_11650 =  x_1530 &  n_8654;
assign n_11651 = ~n_11649 & ~n_11650;
assign n_11652 =  x_2569 & ~n_11651;
assign n_11653 = ~x_2569 &  n_11651;
assign n_11654 = ~n_11652 & ~n_11653;
assign n_11655 =  x_2568 & ~n_8661;
assign n_11656 =  x_1530 &  n_8661;
assign n_11657 = ~n_11655 & ~n_11656;
assign n_11658 =  x_2568 & ~n_11657;
assign n_11659 = ~x_2568 &  n_11657;
assign n_11660 = ~n_11658 & ~n_11659;
assign n_11661 =  x_2567 & ~n_8669;
assign n_11662 =  x_1530 &  n_8669;
assign n_11663 = ~n_11661 & ~n_11662;
assign n_11664 =  x_2567 & ~n_11663;
assign n_11665 = ~x_2567 &  n_11663;
assign n_11666 = ~n_11664 & ~n_11665;
assign n_11667 =  x_2566 & ~n_8676;
assign n_11668 =  x_1530 &  n_8676;
assign n_11669 = ~n_11667 & ~n_11668;
assign n_11670 =  x_2566 & ~n_11669;
assign n_11671 = ~x_2566 &  n_11669;
assign n_11672 = ~n_11670 & ~n_11671;
assign n_11673 =  x_2565 & ~n_8684;
assign n_11674 =  x_1530 &  n_8684;
assign n_11675 = ~n_11673 & ~n_11674;
assign n_11676 =  x_2565 & ~n_11675;
assign n_11677 = ~x_2565 &  n_11675;
assign n_11678 = ~n_11676 & ~n_11677;
assign n_11679 =  x_2564 & ~n_8691;
assign n_11680 =  x_1530 &  n_8691;
assign n_11681 = ~n_11679 & ~n_11680;
assign n_11682 =  x_2564 & ~n_11681;
assign n_11683 = ~x_2564 &  n_11681;
assign n_11684 = ~n_11682 & ~n_11683;
assign n_11685 =  x_2563 & ~n_8699;
assign n_11686 =  x_1530 &  n_8699;
assign n_11687 = ~n_11685 & ~n_11686;
assign n_11688 =  x_2563 & ~n_11687;
assign n_11689 = ~x_2563 &  n_11687;
assign n_11690 = ~n_11688 & ~n_11689;
assign n_11691 =  x_2562 & ~n_8706;
assign n_11692 =  x_1530 &  n_8706;
assign n_11693 = ~n_11691 & ~n_11692;
assign n_11694 =  x_2562 & ~n_11693;
assign n_11695 = ~x_2562 &  n_11693;
assign n_11696 = ~n_11694 & ~n_11695;
assign n_11697 =  x_2561 & ~n_8714;
assign n_11698 =  x_1530 &  n_8714;
assign n_11699 = ~n_11697 & ~n_11698;
assign n_11700 =  x_2561 & ~n_11699;
assign n_11701 = ~x_2561 &  n_11699;
assign n_11702 = ~n_11700 & ~n_11701;
assign n_11703 =  x_2560 & ~n_8721;
assign n_11704 =  x_1530 &  n_8721;
assign n_11705 = ~n_11703 & ~n_11704;
assign n_11706 =  x_2560 & ~n_11705;
assign n_11707 = ~x_2560 &  n_11705;
assign n_11708 = ~n_11706 & ~n_11707;
assign n_11709 =  x_2559 & ~n_8729;
assign n_11710 =  x_1530 &  n_8729;
assign n_11711 = ~n_11709 & ~n_11710;
assign n_11712 =  x_2559 & ~n_11711;
assign n_11713 = ~x_2559 &  n_11711;
assign n_11714 = ~n_11712 & ~n_11713;
assign n_11715 =  x_2558 & ~n_8736;
assign n_11716 =  x_1530 &  n_8736;
assign n_11717 = ~n_11715 & ~n_11716;
assign n_11718 =  x_2558 & ~n_11717;
assign n_11719 = ~x_2558 &  n_11717;
assign n_11720 = ~n_11718 & ~n_11719;
assign n_11721 =  x_2557 & ~n_8744;
assign n_11722 =  x_1530 &  n_8744;
assign n_11723 = ~n_11721 & ~n_11722;
assign n_11724 =  x_2557 & ~n_11723;
assign n_11725 = ~x_2557 &  n_11723;
assign n_11726 = ~n_11724 & ~n_11725;
assign n_11727 =  x_2556 & ~n_8743;
assign n_11728 = ~n_11727 & ~n_8684;
assign n_11729 =  x_2556 & ~n_11728;
assign n_11730 = ~x_2556 &  n_11728;
assign n_11731 = ~n_11729 & ~n_11730;
assign n_11732 = ~x_2555 & ~n_8652;
assign n_11733 = ~n_11732 & ~n_8743;
assign n_11734 =  x_2555 &  n_11733;
assign n_11735 = ~x_2555 & ~n_11733;
assign n_11736 = ~n_11734 & ~n_11735;
assign n_11737 = ~x_2554 & ~n_8636;
assign n_11738 = ~n_11737 & ~n_8652;
assign n_11739 =  x_2554 &  n_11738;
assign n_11740 = ~x_2554 & ~n_11738;
assign n_11741 = ~n_11739 & ~n_11740;
assign n_11742 = ~x_2553 &  n_8625;
assign n_11743 = ~n_8636 & ~n_11742;
assign n_11744 =  x_2553 &  n_11743;
assign n_11745 = ~x_2553 & ~n_11743;
assign n_11746 = ~n_11744 & ~n_11745;
assign n_11747 =  x_2549 &  n_8623;
assign n_11748 =  x_2550 &  n_11747;
assign n_11749 =  x_2551 &  n_11748;
assign n_11750 =  x_2552 & ~n_11749;
assign n_11751 =  n_4383 &  n_8623;
assign n_11752 = ~n_11750 & ~n_11751;
assign n_11753 =  x_2552 & ~n_11752;
assign n_11754 = ~x_2552 &  n_11752;
assign n_11755 = ~n_11753 & ~n_11754;
assign n_11756 = ~x_2551 & ~n_11748;
assign n_11757 = ~n_11756 & ~n_11749;
assign n_11758 =  x_2551 &  n_11757;
assign n_11759 = ~x_2551 & ~n_11757;
assign n_11760 = ~n_11758 & ~n_11759;
assign n_11761 = ~x_2550 & ~n_11747;
assign n_11762 = ~n_11761 & ~n_11748;
assign n_11763 =  x_2550 &  n_11762;
assign n_11764 = ~x_2550 & ~n_11762;
assign n_11765 = ~n_11763 & ~n_11764;
assign n_11766 = ~x_2549 & ~n_8623;
assign n_11767 = ~n_11766 & ~n_11747;
assign n_11768 =  x_2549 &  n_11767;
assign n_11769 = ~x_2549 & ~n_11767;
assign n_11770 = ~n_11768 & ~n_11769;
assign n_11771 = ~n_4370 &  n_5728;
assign n_11772 = ~n_4374 &  n_11771;
assign n_11773 = ~n_11772 & ~n_8622;
assign n_11774 = ~x_2548 &  n_11773;
assign n_11775 =  x_2547 &  x_2548;
assign n_11776 = ~n_4371 & ~n_11775;
assign n_11777 =  n_11771 & ~n_11776;
assign n_11778 = ~n_11771 &  n_11776;
assign n_11779 = ~n_11777 & ~n_11778;
assign n_11780 = ~n_11773 &  n_11779;
assign n_11781 = ~n_11774 & ~n_11780;
assign n_11782 =  x_2548 &  n_11781;
assign n_11783 = ~x_2548 & ~n_11781;
assign n_11784 = ~n_11782 & ~n_11783;
assign n_11785 =  x_2547 & ~n_11773;
assign n_11786 = ~x_2547 &  n_11773;
assign n_11787 = ~n_11785 & ~n_11786;
assign n_11788 =  x_2547 &  n_11787;
assign n_11789 = ~x_2547 & ~n_11787;
assign n_11790 = ~n_11788 & ~n_11789;
assign n_11791 = ~n_11771 & ~n_11775;
assign n_11792 = ~n_4371 &  n_11771;
assign n_11793 = ~n_11791 & ~n_11792;
assign n_11794 = ~n_11773 &  n_11793;
assign n_11795 =  x_2546 &  n_11794;
assign n_11796 = ~x_2546 & ~n_11794;
assign n_11797 = ~n_11795 & ~n_11796;
assign n_11798 =  x_2546 &  n_11797;
assign n_11799 = ~x_2546 & ~n_11797;
assign n_11800 = ~n_11798 & ~n_11799;
assign n_11801 = ~n_11772 & ~n_11795;
assign n_11802 = ~n_4372 &  n_11771;
assign n_11803 = ~n_11801 & ~n_11802;
assign n_11804 = ~x_2545 &  n_11803;
assign n_11805 =  x_2545 & ~n_11803;
assign n_11806 = ~n_11804 & ~n_11805;
assign n_11807 =  x_2545 & ~n_11806;
assign n_11808 = ~x_2545 &  n_11806;
assign n_11809 = ~n_11807 & ~n_11808;
assign n_11810 = ~x_2545 & ~n_11771;
assign n_11811 = ~n_4373 &  n_11771;
assign n_11812 = ~n_11810 & ~n_11811;
assign n_11813 = ~n_11801 &  n_11812;
assign n_11814 =  x_2544 & ~n_11813;
assign n_11815 = ~x_2544 &  n_11813;
assign n_11816 = ~n_11814 & ~n_11815;
assign n_11817 =  x_2544 & ~n_11816;
assign n_11818 = ~x_2544 &  n_11816;
assign n_11819 = ~n_11817 & ~n_11818;
assign n_11820 =  x_2543 & ~n_6054;
assign n_11821 = ~n_11820 & ~n_6080;
assign n_11822 =  x_2543 & ~n_11821;
assign n_11823 = ~x_2543 &  n_11821;
assign n_11824 = ~n_11822 & ~n_11823;
assign n_11825 =  x_2542 & ~n_6088;
assign n_11826 = ~n_6056 & ~n_11825;
assign n_11827 =  x_2542 & ~n_11826;
assign n_11828 = ~x_2542 &  n_11826;
assign n_11829 = ~n_11827 & ~n_11828;
assign n_11830 =  x_2541 &  n_6051;
assign n_11831 = ~n_11830 & ~n_6053;
assign n_11832 =  x_2541 & ~n_11831;
assign n_11833 = ~x_2541 &  n_11831;
assign n_11834 = ~n_11832 & ~n_11833;
assign n_11835 =  x_2540 &  n_6051;
assign n_11836 =  n_1524 &  n_6050;
assign n_11837 = ~n_11835 & ~n_11836;
assign n_11838 =  x_2540 & ~n_11837;
assign n_11839 = ~x_2540 &  n_11837;
assign n_11840 = ~n_11838 & ~n_11839;
assign n_11841 = ~x_2535 &  n_6006;
assign n_11842 = ~x_2538 & ~x_2539;
assign n_11843 = ~x_2537 &  n_11842;
assign n_11844 = ~x_2535 & ~x_2536;
assign n_11845 =  n_11843 &  n_11844;
assign n_11846 =  n_5940 & ~n_11845;
assign n_11847 = ~n_11841 & ~n_11846;
assign n_11848 = ~x_2539 &  n_11847;
assign n_11849 =  x_2538 &  x_2539;
assign n_11850 = ~n_11849 & ~n_11842;
assign n_11851 =  n_5940 & ~n_11850;
assign n_11852 = ~n_5940 &  n_11850;
assign n_11853 = ~n_11851 & ~n_11852;
assign n_11854 = ~n_11847 &  n_11853;
assign n_11855 = ~n_11848 & ~n_11854;
assign n_11856 =  x_2539 &  n_11855;
assign n_11857 = ~x_2539 & ~n_11855;
assign n_11858 = ~n_11856 & ~n_11857;
assign n_11859 = ~x_2538 & ~n_11847;
assign n_11860 =  x_2538 &  n_11847;
assign n_11861 = ~n_11859 & ~n_11860;
assign n_11862 =  x_2538 & ~n_11861;
assign n_11863 = ~x_2538 &  n_11861;
assign n_11864 = ~n_11862 & ~n_11863;
assign n_11865 = ~n_5940 &  n_11849;
assign n_11866 =  n_5940 &  n_11842;
assign n_11867 = ~n_11865 & ~n_11866;
assign n_11868 = ~n_11847 & ~n_11867;
assign n_11869 =  x_2537 &  n_11868;
assign n_11870 = ~x_2537 & ~n_11868;
assign n_11871 = ~n_11869 & ~n_11870;
assign n_11872 =  x_2537 &  n_11871;
assign n_11873 = ~x_2537 & ~n_11871;
assign n_11874 = ~n_11872 & ~n_11873;
assign n_11875 =  x_2537 &  n_11865;
assign n_11876 =  n_5940 &  n_11843;
assign n_11877 = ~n_11875 & ~n_11876;
assign n_11878 = ~n_11847 & ~n_11877;
assign n_11879 = ~x_2536 &  n_11878;
assign n_11880 =  x_2536 & ~n_11878;
assign n_11881 = ~n_11879 & ~n_11880;
assign n_11882 =  x_2536 & ~n_11881;
assign n_11883 = ~x_2536 &  n_11881;
assign n_11884 = ~n_11882 & ~n_11883;
assign n_11885 =  x_2536 & ~n_11875;
assign n_11886 = ~x_2536 & ~n_11876;
assign n_11887 = ~n_11886 & ~n_11847;
assign n_11888 = ~n_11885 &  n_11887;
assign n_11889 =  x_2535 &  n_11888;
assign n_11890 = ~x_2535 & ~n_11888;
assign n_11891 = ~n_11889 & ~n_11890;
assign n_11892 =  x_2535 &  n_11891;
assign n_11893 = ~x_2535 & ~n_11891;
assign n_11894 = ~n_11892 & ~n_11893;
assign n_11895 =  x_2534 & ~n_5940;
assign n_11896 = ~n_6006 & ~n_11895;
assign n_11897 =  x_2534 & ~n_11896;
assign n_11898 = ~x_2534 &  n_11896;
assign n_11899 = ~n_11897 & ~n_11898;
assign n_11900 = ~x_2529 &  n_5988;
assign n_11901 = ~x_2532 & ~x_2533;
assign n_11902 = ~x_2531 &  n_11901;
assign n_11903 = ~x_2529 & ~x_2530;
assign n_11904 =  n_11902 &  n_11903;
assign n_11905 =  n_5940 & ~n_11904;
assign n_11906 = ~n_11900 & ~n_11905;
assign n_11907 = ~x_2533 &  n_11906;
assign n_11908 =  x_2532 &  x_2533;
assign n_11909 = ~n_11908 & ~n_11901;
assign n_11910 =  n_5940 & ~n_11909;
assign n_11911 = ~n_5940 &  n_11909;
assign n_11912 = ~n_11910 & ~n_11911;
assign n_11913 = ~n_11906 &  n_11912;
assign n_11914 = ~n_11907 & ~n_11913;
assign n_11915 =  x_2533 &  n_11914;
assign n_11916 = ~x_2533 & ~n_11914;
assign n_11917 = ~n_11915 & ~n_11916;
assign n_11918 = ~x_2532 & ~n_11906;
assign n_11919 =  x_2532 &  n_11906;
assign n_11920 = ~n_11918 & ~n_11919;
assign n_11921 =  x_2532 & ~n_11920;
assign n_11922 = ~x_2532 &  n_11920;
assign n_11923 = ~n_11921 & ~n_11922;
assign n_11924 = ~n_5940 &  n_11908;
assign n_11925 =  n_5940 &  n_11901;
assign n_11926 = ~n_11924 & ~n_11925;
assign n_11927 = ~n_11906 & ~n_11926;
assign n_11928 =  x_2531 &  n_11927;
assign n_11929 = ~x_2531 & ~n_11927;
assign n_11930 = ~n_11928 & ~n_11929;
assign n_11931 =  x_2531 &  n_11930;
assign n_11932 = ~x_2531 & ~n_11930;
assign n_11933 = ~n_11931 & ~n_11932;
assign n_11934 =  x_2531 &  n_11924;
assign n_11935 =  n_5940 &  n_11902;
assign n_11936 = ~n_11934 & ~n_11935;
assign n_11937 = ~n_11906 & ~n_11936;
assign n_11938 = ~x_2530 &  n_11937;
assign n_11939 =  x_2530 & ~n_11937;
assign n_11940 = ~n_11938 & ~n_11939;
assign n_11941 =  x_2530 & ~n_11940;
assign n_11942 = ~x_2530 &  n_11940;
assign n_11943 = ~n_11941 & ~n_11942;
assign n_11944 =  x_2530 & ~n_11934;
assign n_11945 = ~x_2530 & ~n_11935;
assign n_11946 = ~n_11945 & ~n_11906;
assign n_11947 = ~n_11944 &  n_11946;
assign n_11948 =  x_2529 &  n_11947;
assign n_11949 = ~x_2529 & ~n_11947;
assign n_11950 = ~n_11948 & ~n_11949;
assign n_11951 =  x_2529 &  n_11950;
assign n_11952 = ~x_2529 & ~n_11950;
assign n_11953 = ~n_11951 & ~n_11952;
assign n_11954 =  x_2528 & ~n_5940;
assign n_11955 = ~n_5988 & ~n_11954;
assign n_11956 =  x_2528 & ~n_11955;
assign n_11957 = ~x_2528 &  n_11955;
assign n_11958 = ~n_11956 & ~n_11957;
assign n_11959 =  x_2526 &  n_6037;
assign n_11960 =  x_2527 &  n_1522;
assign n_11961 = ~n_11959 & ~n_11960;
assign n_11962 =  x_2527 & ~n_11961;
assign n_11963 = ~x_2527 &  n_11961;
assign n_11964 = ~n_11962 & ~n_11963;
assign n_11965 =  x_2525 &  n_6037;
assign n_11966 =  x_2526 &  n_1522;
assign n_11967 = ~n_11965 & ~n_11966;
assign n_11968 =  x_2526 & ~n_11967;
assign n_11969 = ~x_2526 &  n_11967;
assign n_11970 = ~n_11968 & ~n_11969;
assign n_11971 =  x_2525 &  n_1522;
assign n_11972 = ~n_6037 & ~n_11971;
assign n_11973 =  x_2525 & ~n_11972;
assign n_11974 = ~x_2525 &  n_11972;
assign n_11975 = ~n_11973 & ~n_11974;
assign n_11976 = ~x_226 &  n_1739;
assign n_11977 = ~x_2524 & ~n_11976;
assign n_11978 =  x_2524 & ~n_11977;
assign n_11979 = ~x_2524 &  n_11977;
assign n_11980 = ~n_11978 & ~n_11979;
assign n_11981 =  n_1708 & ~n_1702;
assign n_11982 = ~n_1696 &  n_11981;
assign n_11983 = ~n_1690 &  n_11982;
assign n_11984 = ~n_1684 &  n_11983;
assign n_11985 = ~n_1678 &  n_11984;
assign n_11986 = ~n_1672 &  n_11985;
assign n_11987 = ~n_1666 &  n_11986;
assign n_11988 = ~n_1660 &  n_11987;
assign n_11989 = ~n_1654 &  n_11988;
assign n_11990 = ~n_1648 &  n_11989;
assign n_11991 = ~n_1642 &  n_11990;
assign n_11992 = ~n_1636 &  n_11991;
assign n_11993 = ~n_1630 &  n_11992;
assign n_11994 = ~n_1624 &  n_11993;
assign n_11995 = ~n_1618 &  n_11994;
assign n_11996 = ~n_1612 &  n_11995;
assign n_11997 = ~n_1606 &  n_11996;
assign n_11998 = ~n_1600 &  n_11997;
assign n_11999 = ~n_1594 &  n_11998;
assign n_12000 = ~n_1588 &  n_11999;
assign n_12001 = ~n_1582 &  n_12000;
assign n_12002 = ~n_1576 &  n_12001;
assign n_12003 = ~n_1570 &  n_12002;
assign n_12004 = ~n_1564 &  n_12003;
assign n_12005 = ~n_1558 &  n_12004;
assign n_12006 = ~n_1552 &  n_12005;
assign n_12007 = ~n_1546 &  n_12006;
assign n_12008 = ~n_1540 &  n_12007;
assign n_12009 = ~n_1534 &  n_12008;
assign n_12010 = ~n_1528 &  n_12009;
assign n_12011 = ~n_12010 &  n_3948;
assign n_12012 =  n_12010 & ~n_3948;
assign n_12013 = ~n_12011 & ~n_12012;
assign n_12014 =  x_2523 & ~n_12013;
assign n_12015 = ~x_2523 &  n_12013;
assign n_12016 = ~n_12014 & ~n_12015;
assign n_12017 =  x_2522 & ~n_3948;
assign n_12018 = ~x_2522 &  n_3948;
assign n_12019 = ~n_12017 & ~n_12018;
assign n_12020 =  n_1528 & ~n_12009;
assign n_12021 = ~n_12020 & ~n_12010;
assign n_12022 =  x_2521 & ~n_12021;
assign n_12023 = ~x_2521 &  n_12021;
assign n_12024 = ~n_12022 & ~n_12023;
assign n_12025 =  n_1534 & ~n_12008;
assign n_12026 = ~n_12025 & ~n_12009;
assign n_12027 =  x_2520 & ~n_12026;
assign n_12028 = ~x_2520 &  n_12026;
assign n_12029 = ~n_12027 & ~n_12028;
assign n_12030 =  n_1540 & ~n_12007;
assign n_12031 = ~n_12030 & ~n_12008;
assign n_12032 =  x_2519 & ~n_12031;
assign n_12033 = ~x_2519 &  n_12031;
assign n_12034 = ~n_12032 & ~n_12033;
assign n_12035 =  n_1546 & ~n_12006;
assign n_12036 = ~n_12035 & ~n_12007;
assign n_12037 =  x_2518 & ~n_12036;
assign n_12038 = ~x_2518 &  n_12036;
assign n_12039 = ~n_12037 & ~n_12038;
assign n_12040 =  n_1552 & ~n_12005;
assign n_12041 = ~n_12040 & ~n_12006;
assign n_12042 =  x_2517 & ~n_12041;
assign n_12043 = ~x_2517 &  n_12041;
assign n_12044 = ~n_12042 & ~n_12043;
assign n_12045 =  n_1558 & ~n_12004;
assign n_12046 = ~n_12045 & ~n_12005;
assign n_12047 =  x_2516 & ~n_12046;
assign n_12048 = ~x_2516 &  n_12046;
assign n_12049 = ~n_12047 & ~n_12048;
assign n_12050 =  n_1564 & ~n_12003;
assign n_12051 = ~n_12050 & ~n_12004;
assign n_12052 =  x_2515 & ~n_12051;
assign n_12053 = ~x_2515 &  n_12051;
assign n_12054 = ~n_12052 & ~n_12053;
assign n_12055 =  n_1570 & ~n_12002;
assign n_12056 = ~n_12055 & ~n_12003;
assign n_12057 =  x_2514 & ~n_12056;
assign n_12058 = ~x_2514 &  n_12056;
assign n_12059 = ~n_12057 & ~n_12058;
assign n_12060 =  n_1576 & ~n_12001;
assign n_12061 = ~n_12060 & ~n_12002;
assign n_12062 =  x_2513 & ~n_12061;
assign n_12063 = ~x_2513 &  n_12061;
assign n_12064 = ~n_12062 & ~n_12063;
assign n_12065 =  n_1582 & ~n_12000;
assign n_12066 = ~n_12065 & ~n_12001;
assign n_12067 =  x_2512 & ~n_12066;
assign n_12068 = ~x_2512 &  n_12066;
assign n_12069 = ~n_12067 & ~n_12068;
assign n_12070 =  n_1588 & ~n_11999;
assign n_12071 = ~n_12070 & ~n_12000;
assign n_12072 =  x_2511 & ~n_12071;
assign n_12073 = ~x_2511 &  n_12071;
assign n_12074 = ~n_12072 & ~n_12073;
assign n_12075 =  n_1594 & ~n_11998;
assign n_12076 = ~n_12075 & ~n_11999;
assign n_12077 =  x_2510 & ~n_12076;
assign n_12078 = ~x_2510 &  n_12076;
assign n_12079 = ~n_12077 & ~n_12078;
assign n_12080 =  n_1600 & ~n_11997;
assign n_12081 = ~n_12080 & ~n_11998;
assign n_12082 =  x_2509 & ~n_12081;
assign n_12083 = ~x_2509 &  n_12081;
assign n_12084 = ~n_12082 & ~n_12083;
assign n_12085 =  n_1606 & ~n_11996;
assign n_12086 = ~n_12085 & ~n_11997;
assign n_12087 =  x_2508 & ~n_12086;
assign n_12088 = ~x_2508 &  n_12086;
assign n_12089 = ~n_12087 & ~n_12088;
assign n_12090 =  n_1612 & ~n_11995;
assign n_12091 = ~n_12090 & ~n_11996;
assign n_12092 =  x_2507 & ~n_12091;
assign n_12093 = ~x_2507 &  n_12091;
assign n_12094 = ~n_12092 & ~n_12093;
assign n_12095 =  n_1618 & ~n_11994;
assign n_12096 = ~n_12095 & ~n_11995;
assign n_12097 =  x_2506 & ~n_12096;
assign n_12098 = ~x_2506 &  n_12096;
assign n_12099 = ~n_12097 & ~n_12098;
assign n_12100 =  n_1624 & ~n_11993;
assign n_12101 = ~n_12100 & ~n_11994;
assign n_12102 =  x_2505 & ~n_12101;
assign n_12103 = ~x_2505 &  n_12101;
assign n_12104 = ~n_12102 & ~n_12103;
assign n_12105 =  n_1630 & ~n_11992;
assign n_12106 = ~n_12105 & ~n_11993;
assign n_12107 =  x_2504 & ~n_12106;
assign n_12108 = ~x_2504 &  n_12106;
assign n_12109 = ~n_12107 & ~n_12108;
assign n_12110 =  n_1636 & ~n_11991;
assign n_12111 = ~n_12110 & ~n_11992;
assign n_12112 =  x_2503 & ~n_12111;
assign n_12113 = ~x_2503 &  n_12111;
assign n_12114 = ~n_12112 & ~n_12113;
assign n_12115 =  n_1642 & ~n_11990;
assign n_12116 = ~n_12115 & ~n_11991;
assign n_12117 =  x_2502 & ~n_12116;
assign n_12118 = ~x_2502 &  n_12116;
assign n_12119 = ~n_12117 & ~n_12118;
assign n_12120 =  n_1648 & ~n_11989;
assign n_12121 = ~n_12120 & ~n_11990;
assign n_12122 =  x_2501 & ~n_12121;
assign n_12123 = ~x_2501 &  n_12121;
assign n_12124 = ~n_12122 & ~n_12123;
assign n_12125 =  n_1654 & ~n_11988;
assign n_12126 = ~n_12125 & ~n_11989;
assign n_12127 =  x_2500 & ~n_12126;
assign n_12128 = ~x_2500 &  n_12126;
assign n_12129 = ~n_12127 & ~n_12128;
assign n_12130 =  n_1660 & ~n_11987;
assign n_12131 = ~n_12130 & ~n_11988;
assign n_12132 =  x_2499 & ~n_12131;
assign n_12133 = ~x_2499 &  n_12131;
assign n_12134 = ~n_12132 & ~n_12133;
assign n_12135 =  n_1666 & ~n_11986;
assign n_12136 = ~n_11987 & ~n_12135;
assign n_12137 =  x_2498 & ~n_12136;
assign n_12138 = ~x_2498 &  n_12136;
assign n_12139 = ~n_12137 & ~n_12138;
assign n_12140 =  n_1672 & ~n_11985;
assign n_12141 = ~n_12140 & ~n_11986;
assign n_12142 =  x_2497 & ~n_12141;
assign n_12143 = ~x_2497 &  n_12141;
assign n_12144 = ~n_12142 & ~n_12143;
assign n_12145 =  n_1678 & ~n_11984;
assign n_12146 = ~n_12145 & ~n_11985;
assign n_12147 =  x_2496 & ~n_12146;
assign n_12148 = ~x_2496 &  n_12146;
assign n_12149 = ~n_12147 & ~n_12148;
assign n_12150 =  n_1684 & ~n_11983;
assign n_12151 = ~n_12150 & ~n_11984;
assign n_12152 =  x_2495 & ~n_12151;
assign n_12153 = ~x_2495 &  n_12151;
assign n_12154 = ~n_12152 & ~n_12153;
assign n_12155 =  n_1690 & ~n_11982;
assign n_12156 = ~n_12155 & ~n_11983;
assign n_12157 =  x_2494 & ~n_12156;
assign n_12158 = ~x_2494 &  n_12156;
assign n_12159 = ~n_12157 & ~n_12158;
assign n_12160 =  n_1696 & ~n_11981;
assign n_12161 = ~n_12160 & ~n_11982;
assign n_12162 =  x_2493 & ~n_12161;
assign n_12163 = ~x_2493 &  n_12161;
assign n_12164 = ~n_12162 & ~n_12163;
assign n_12165 = ~n_11981 & ~n_3959;
assign n_12166 =  x_2492 &  n_12165;
assign n_12167 = ~x_2492 & ~n_12165;
assign n_12168 = ~n_12166 & ~n_12167;
assign n_12169 = ~n_5924 &  n_5935;
assign n_12170 = ~n_5835 &  n_12169;
assign n_12171 = ~n_5935 & ~n_5928;
assign n_12172 =  n_5925 &  n_12171;
assign n_12173 = ~n_12170 & ~n_12172;
assign n_12174 =  n_5926 & ~n_12173;
assign n_12175 = ~x_2473 & ~x_2489;
assign n_12176 =  n_12174 & ~n_12175;
assign n_12177 =  x_2490 &  x_2491;
assign n_12178 = ~x_2483 & ~n_12177;
assign n_12179 =  x_2490 & ~x_2491;
assign n_12180 = ~x_2478 & ~n_12179;
assign n_12181 = ~x_2489 & ~x_2490;
assign n_12182 =  x_2491 &  n_12181;
assign n_12183 = ~x_2468 & ~n_12182;
assign n_12184 =  x_2463 &  x_2491;
assign n_12185 = ~n_12183 & ~n_12184;
assign n_12186 = ~n_12180 & ~n_12185;
assign n_12187 = ~n_12178 & ~n_12186;
assign n_12188 =  n_12176 & ~n_12187;
assign n_12189 =  n_5816 & ~n_12173;
assign n_12190 =  x_2491 & ~n_12189;
assign n_12191 = ~n_5852 &  n_5921;
assign n_12192 = ~n_5869 & ~n_12191;
assign n_12193 = ~n_5887 & ~n_12192;
assign n_12194 =  n_12189 &  n_12193;
assign n_12195 = ~n_12190 & ~n_12194;
assign n_12196 = ~n_12188 &  n_12195;
assign n_12197 =  x_2491 & ~n_12196;
assign n_12198 = ~x_2491 &  n_12196;
assign n_12199 = ~n_12197 & ~n_12198;
assign n_12200 = ~n_12180 & ~n_12178;
assign n_12201 =  x_2463 &  x_2468;
assign n_12202 =  x_2490 &  n_12201;
assign n_12203 =  n_12200 & ~n_12202;
assign n_12204 =  n_12176 & ~n_12203;
assign n_12205 =  x_2490 & ~n_12189;
assign n_12206 = ~n_5870 & ~n_5887;
assign n_12207 =  n_12189 &  n_12206;
assign n_12208 = ~n_12205 & ~n_12207;
assign n_12209 = ~n_12204 &  n_12208;
assign n_12210 =  x_2490 & ~n_12209;
assign n_12211 = ~x_2490 &  n_12209;
assign n_12212 = ~n_12210 & ~n_12211;
assign n_12213 = ~x_2491 &  n_12181;
assign n_12214 = ~x_2463 & ~n_12213;
assign n_12215 =  n_12200 & ~n_12183;
assign n_12216 = ~n_12214 &  n_12215;
assign n_12217 =  n_5925 &  n_12216;
assign n_12218 =  n_12189 & ~n_12217;
assign n_12219 =  x_2489 & ~n_12218;
assign n_12220 =  n_5925 &  n_12175;
assign n_12221 = ~n_5887 & ~n_12220;
assign n_12222 =  n_12189 & ~n_12221;
assign n_12223 = ~n_12219 & ~n_12222;
assign n_12224 =  x_2489 & ~n_12223;
assign n_12225 = ~x_2489 &  n_12223;
assign n_12226 = ~n_12224 & ~n_12225;
assign n_12227 = ~x_2488 & ~n_12189;
assign n_12228 =  x_2487 &  x_2488;
assign n_12229 = ~n_5927 & ~n_12228;
assign n_12230 =  n_12170 & ~n_12229;
assign n_12231 = ~n_12170 &  n_12229;
assign n_12232 = ~n_12230 & ~n_12231;
assign n_12233 =  n_12189 &  n_12232;
assign n_12234 = ~n_12227 & ~n_12233;
assign n_12235 =  x_2488 &  n_12234;
assign n_12236 = ~x_2488 & ~n_12234;
assign n_12237 = ~n_12235 & ~n_12236;
assign n_12238 =  x_2487 & ~n_12189;
assign n_12239 = ~x_2487 &  n_12189;
assign n_12240 = ~n_12238 & ~n_12239;
assign n_12241 =  x_2487 & ~n_12240;
assign n_12242 = ~x_2487 &  n_12240;
assign n_12243 = ~n_12241 & ~n_12242;
assign n_12244 = ~n_12170 & ~n_12228;
assign n_12245 =  n_12170 & ~n_5927;
assign n_12246 = ~n_12244 & ~n_12245;
assign n_12247 =  n_12189 &  n_12246;
assign n_12248 = ~x_2486 &  n_12247;
assign n_12249 =  x_2486 & ~n_12247;
assign n_12250 = ~n_12248 & ~n_12249;
assign n_12251 =  x_2486 & ~n_12250;
assign n_12252 = ~x_2486 &  n_12250;
assign n_12253 = ~n_12251 & ~n_12252;
assign n_12254 =  n_5930 & ~n_5932;
assign n_12255 =  x_2485 &  n_12254;
assign n_12256 = ~x_2485 & ~n_12254;
assign n_12257 = ~n_12255 & ~n_12256;
assign n_12258 =  n_5830 & ~n_5832;
assign n_12259 =  x_2484 &  n_12258;
assign n_12260 = ~x_2484 & ~n_12258;
assign n_12261 = ~n_12259 & ~n_12260;
assign n_12262 =  n_12174 &  n_12177;
assign n_12263 = ~n_5926 & ~n_12173;
assign n_12264 =  n_5868 &  n_12263;
assign n_12265 =  x_2483 & ~n_12264;
assign n_12266 = ~n_12262 & ~n_12265;
assign n_12267 =  x_2483 & ~n_12266;
assign n_12268 = ~x_2483 &  n_12266;
assign n_12269 = ~n_12267 & ~n_12268;
assign n_12270 =  x_2482 & ~n_12262;
assign n_12271 =  n_4326 &  n_12262;
assign n_12272 = ~n_12270 & ~n_12271;
assign n_12273 =  x_2482 & ~n_12272;
assign n_12274 = ~x_2482 &  n_12272;
assign n_12275 = ~n_12273 & ~n_12274;
assign n_12276 =  x_2481 & ~n_12262;
assign n_12277 =  i_143 &  n_12262;
assign n_12278 = ~n_12276 & ~n_12277;
assign n_12279 =  x_2481 & ~n_12278;
assign n_12280 = ~x_2481 &  n_12278;
assign n_12281 = ~n_12279 & ~n_12280;
assign n_12282 =  x_2480 & ~n_12262;
assign n_12283 =  i_145 &  n_12262;
assign n_12284 = ~n_12282 & ~n_12283;
assign n_12285 =  x_2480 & ~n_12284;
assign n_12286 = ~x_2480 &  n_12284;
assign n_12287 = ~n_12285 & ~n_12286;
assign n_12288 =  x_2479 & ~n_12262;
assign n_12289 =  n_4323 &  n_12262;
assign n_12290 = ~n_12288 & ~n_12289;
assign n_12291 =  x_2479 & ~n_12290;
assign n_12292 = ~x_2479 &  n_12290;
assign n_12293 = ~n_12291 & ~n_12292;
assign n_12294 =  n_12174 &  n_12179;
assign n_12295 =  n_5851 &  n_12263;
assign n_12296 =  x_2478 & ~n_12295;
assign n_12297 = ~n_12294 & ~n_12296;
assign n_12298 =  x_2478 & ~n_12297;
assign n_12299 = ~x_2478 &  n_12297;
assign n_12300 = ~n_12298 & ~n_12299;
assign n_12301 =  x_2477 & ~n_12294;
assign n_12302 =  n_4326 &  n_12294;
assign n_12303 = ~n_12301 & ~n_12302;
assign n_12304 =  x_2477 & ~n_12303;
assign n_12305 = ~x_2477 &  n_12303;
assign n_12306 = ~n_12304 & ~n_12305;
assign n_12307 =  x_2476 & ~n_12294;
assign n_12308 =  n_4323 &  n_12294;
assign n_12309 = ~n_12307 & ~n_12308;
assign n_12310 =  x_2476 & ~n_12309;
assign n_12311 = ~x_2476 &  n_12309;
assign n_12312 = ~n_12310 & ~n_12311;
assign n_12313 =  x_2475 & ~n_12294;
assign n_12314 =  i_143 &  n_12294;
assign n_12315 = ~n_12313 & ~n_12314;
assign n_12316 =  x_2475 & ~n_12315;
assign n_12317 = ~x_2475 &  n_12315;
assign n_12318 = ~n_12316 & ~n_12317;
assign n_12319 =  x_2474 & ~n_12294;
assign n_12320 =  i_145 &  n_12294;
assign n_12321 = ~n_12319 & ~n_12320;
assign n_12322 =  x_2474 & ~n_12321;
assign n_12323 = ~x_2474 &  n_12321;
assign n_12324 = ~n_12322 & ~n_12323;
assign n_12325 =  n_5886 & ~n_12173;
assign n_12326 =  x_2473 & ~n_12325;
assign n_12327 = ~n_12176 & ~n_12326;
assign n_12328 =  x_2473 & ~n_12327;
assign n_12329 = ~x_2473 &  n_12327;
assign n_12330 = ~n_12328 & ~n_12329;
assign n_12331 =  x_2489 &  n_12174;
assign n_12332 =  x_2472 & ~n_12331;
assign n_12333 =  n_4326 &  n_12331;
assign n_12334 = ~n_12332 & ~n_12333;
assign n_12335 =  x_2472 & ~n_12334;
assign n_12336 = ~x_2472 &  n_12334;
assign n_12337 = ~n_12335 & ~n_12336;
assign n_12338 =  x_2471 & ~n_12331;
assign n_12339 =  n_4323 &  n_12331;
assign n_12340 = ~n_12338 & ~n_12339;
assign n_12341 =  x_2471 & ~n_12340;
assign n_12342 = ~x_2471 &  n_12340;
assign n_12343 = ~n_12341 & ~n_12342;
assign n_12344 =  x_2470 & ~n_12331;
assign n_12345 =  i_143 &  n_12331;
assign n_12346 = ~n_12344 & ~n_12345;
assign n_12347 =  x_2470 & ~n_12346;
assign n_12348 = ~x_2470 &  n_12346;
assign n_12349 = ~n_12347 & ~n_12348;
assign n_12350 =  x_2469 & ~n_12331;
assign n_12351 =  i_145 &  n_12331;
assign n_12352 = ~n_12350 & ~n_12351;
assign n_12353 =  x_2469 & ~n_12352;
assign n_12354 = ~x_2469 &  n_12352;
assign n_12355 = ~n_12353 & ~n_12354;
assign n_12356 =  n_12174 &  n_12182;
assign n_12357 =  n_5920 &  n_12263;
assign n_12358 =  x_2468 & ~n_12357;
assign n_12359 = ~n_12356 & ~n_12358;
assign n_12360 =  x_2468 & ~n_12359;
assign n_12361 = ~x_2468 &  n_12359;
assign n_12362 = ~n_12360 & ~n_12361;
assign n_12363 =  x_2467 & ~n_12356;
assign n_12364 =  n_4326 &  n_12356;
assign n_12365 = ~n_12363 & ~n_12364;
assign n_12366 =  x_2467 & ~n_12365;
assign n_12367 = ~x_2467 &  n_12365;
assign n_12368 = ~n_12366 & ~n_12367;
assign n_12369 =  x_2466 & ~n_12356;
assign n_12370 =  i_143 &  n_12356;
assign n_12371 = ~n_12369 & ~n_12370;
assign n_12372 =  x_2466 & ~n_12371;
assign n_12373 = ~x_2466 &  n_12371;
assign n_12374 = ~n_12372 & ~n_12373;
assign n_12375 =  x_2465 & ~n_12356;
assign n_12376 =  n_4323 &  n_12356;
assign n_12377 = ~n_12375 & ~n_12376;
assign n_12378 =  x_2465 & ~n_12377;
assign n_12379 = ~x_2465 &  n_12377;
assign n_12380 = ~n_12378 & ~n_12379;
assign n_12381 =  x_2464 & ~n_12356;
assign n_12382 =  i_145 &  n_12356;
assign n_12383 = ~n_12381 & ~n_12382;
assign n_12384 =  x_2464 & ~n_12383;
assign n_12385 = ~x_2464 &  n_12383;
assign n_12386 = ~n_12384 & ~n_12385;
assign n_12387 =  n_12213 &  n_12174;
assign n_12388 =  n_5903 &  n_12263;
assign n_12389 =  x_2463 & ~n_12388;
assign n_12390 = ~n_12387 & ~n_12389;
assign n_12391 =  x_2463 & ~n_12390;
assign n_12392 = ~x_2463 &  n_12390;
assign n_12393 = ~n_12391 & ~n_12392;
assign n_12394 =  x_2462 & ~n_12387;
assign n_12395 =  n_4323 &  n_12387;
assign n_12396 = ~n_12394 & ~n_12395;
assign n_12397 =  x_2462 & ~n_12396;
assign n_12398 = ~x_2462 &  n_12396;
assign n_12399 = ~n_12397 & ~n_12398;
assign n_12400 =  x_2461 & ~n_12387;
assign n_12401 =  n_4326 &  n_12387;
assign n_12402 = ~n_12400 & ~n_12401;
assign n_12403 =  x_2461 & ~n_12402;
assign n_12404 = ~x_2461 &  n_12402;
assign n_12405 = ~n_12403 & ~n_12404;
assign n_12406 =  x_2460 & ~n_12387;
assign n_12407 =  i_145 &  n_12387;
assign n_12408 = ~n_12406 & ~n_12407;
assign n_12409 =  x_2460 & ~n_12408;
assign n_12410 = ~x_2460 &  n_12408;
assign n_12411 = ~n_12409 & ~n_12410;
assign n_12412 =  x_2459 & ~n_12387;
assign n_12413 =  i_143 &  n_12387;
assign n_12414 = ~n_12412 & ~n_12413;
assign n_12415 =  x_2459 & ~n_12414;
assign n_12416 = ~x_2459 &  n_12414;
assign n_12417 = ~n_12415 & ~n_12416;
assign n_12418 =  x_2458 &  n_5930;
assign n_12419 = ~x_2458 & ~n_5930;
assign n_12420 = ~n_12418 & ~n_12419;
assign n_12421 =  x_2457 &  n_5830;
assign n_12422 = ~x_2457 & ~n_5830;
assign n_12423 = ~n_12421 & ~n_12422;
assign n_12424 = ~x_2442 &  n_3559;
assign n_12425 =  n_3570 & ~n_12424;
assign n_12426 = ~x_2440 &  n_12425;
assign n_12427 =  x_2454 &  x_2455;
assign n_12428 =  n_12426 &  n_12427;
assign n_12429 = ~x_2456 & ~n_12428;
assign n_12430 =  n_12426 & ~n_12427;
assign n_12431 = ~n_3563 & ~n_12425;
assign n_12432 = ~x_2440 &  n_12431;
assign n_12433 =  x_2456 & ~n_12432;
assign n_12434 = ~n_12430 &  n_12433;
assign n_12435 = ~n_12429 & ~n_12434;
assign n_12436 =  x_2456 &  n_12435;
assign n_12437 = ~x_2456 & ~n_12435;
assign n_12438 = ~n_12436 & ~n_12437;
assign n_12439 =  x_2455 &  n_12432;
assign n_12440 = ~n_6042 &  n_12430;
assign n_12441 = ~n_12439 & ~n_12440;
assign n_12442 =  x_2455 & ~n_12441;
assign n_12443 = ~x_2455 &  n_12441;
assign n_12444 = ~n_12442 & ~n_12443;
assign n_12445 =  x_2454 &  n_12431;
assign n_12446 = ~x_2454 &  n_12425;
assign n_12447 = ~x_2440 & ~n_12446;
assign n_12448 = ~n_12445 &  n_12447;
assign n_12449 =  x_2454 & ~n_12448;
assign n_12450 = ~x_2454 &  n_12448;
assign n_12451 = ~n_12449 & ~n_12450;
assign n_12452 = ~x_1495 &  n_5992;
assign n_12453 =  x_2453 &  n_12452;
assign n_12454 = ~n_12453 &  n_5995;
assign n_12455 =  x_2453 &  n_12454;
assign n_12456 = ~x_2453 & ~n_12454;
assign n_12457 = ~n_12455 & ~n_12456;
assign n_12458 = ~n_12453 & ~n_5994;
assign n_12459 = ~x_1498 &  n_12458;
assign n_12460 =  n_5993 & ~n_12459;
assign n_12461 = ~n_3612 & ~n_12460;
assign n_12462 =  x_2452 &  n_12461;
assign n_12463 = ~x_2452 & ~n_12461;
assign n_12464 = ~n_12462 & ~n_12463;
assign n_12465 =  n_3563 &  n_6067;
assign n_12466 = ~x_2451 & ~n_12465;
assign n_12467 =  x_1761 & ~n_12466;
assign n_12468 = ~x_1768 &  x_2451;
assign n_12469 = ~n_3570 &  n_12468;
assign n_12470 = ~n_12467 & ~n_12469;
assign n_12471 =  x_2451 & ~n_12470;
assign n_12472 = ~x_2451 &  n_12470;
assign n_12473 = ~n_12471 & ~n_12472;
assign n_12474 =  x_2450 & ~n_3626;
assign n_12475 = ~n_3612 &  n_12474;
assign n_12476 = ~n_3634 & ~n_12475;
assign n_12477 =  x_2450 & ~n_12476;
assign n_12478 = ~x_2450 &  n_12476;
assign n_12479 = ~n_12477 & ~n_12478;
assign n_12480 =  x_2449 & ~n_3714;
assign n_12481 = ~x_2449 &  n_3714;
assign n_12482 = ~n_12480 & ~n_12481;
assign n_12483 = ~x_2448 & ~n_3634;
assign n_12484 =  x_2448 & ~n_12483;
assign n_12485 = ~x_2448 &  n_12483;
assign n_12486 = ~n_12484 & ~n_12485;
assign n_12487 = ~x_2447 & ~n_3634;
assign n_12488 = ~n_12487 & ~n_3716;
assign n_12489 =  x_2447 &  n_12488;
assign n_12490 = ~x_2447 & ~n_12488;
assign n_12491 = ~n_12489 & ~n_12490;
assign n_12492 =  x_2446 & ~n_3665;
assign n_12493 = ~x_2446 &  n_3665;
assign n_12494 = ~n_12492 & ~n_12493;
assign n_12495 =  x_2445 & ~n_3658;
assign n_12496 = ~x_2445 &  n_3658;
assign n_12497 = ~n_12495 & ~n_12496;
assign n_12498 =  x_2444 & ~n_3650;
assign n_12499 = ~x_2444 &  n_3650;
assign n_12500 = ~n_12498 & ~n_12499;
assign n_12501 =  x_2443 & ~n_3640;
assign n_12502 = ~x_2443 &  n_3640;
assign n_12503 = ~n_12501 & ~n_12502;
assign n_12504 =  x_2442 & ~n_3670;
assign n_12505 = ~x_2442 &  n_3670;
assign n_12506 = ~n_12504 & ~n_12505;
assign n_12507 =  x_2441 &  n_5811;
assign n_12508 = ~x_2441 & ~n_5811;
assign n_12509 = ~n_12507 & ~n_12508;
assign n_12510 = ~x_1765 & ~x_1766;
assign n_12511 =  x_309 & ~x_1489;
assign n_12512 =  x_310 &  n_12511;
assign n_12513 =  n_12510 &  n_12512;
assign n_12514 = ~x_1755 & ~x_1757;
assign n_12515 = ~x_1756 &  n_12514;
assign n_12516 =  x_1487 & ~n_12515;
assign n_12517 = ~x_1488 & ~n_12516;
assign n_12518 = ~x_1765 & ~n_12517;
assign n_12519 =  x_1762 &  n_12465;
assign n_12520 = ~n_12518 &  n_12519;
assign n_12521 = ~n_12513 & ~n_12520;
assign n_12522 =  x_1767 & ~n_12521;
assign n_12523 =  x_1756 &  x_1759;
assign n_12524 =  n_12511 &  n_12523;
assign n_12525 = ~n_12513 &  n_12524;
assign n_12526 =  x_1756 &  n_12514;
assign n_12527 = ~n_12525 & ~n_12526;
assign n_12528 = ~n_12522 &  n_12527;
assign n_12529 = ~x_310 &  n_12511;
assign n_12530 =  n_12510 &  n_12529;
assign n_12531 = ~x_1765 &  x_1766;
assign n_12532 = ~x_1489 &  n_12531;
assign n_12533 =  n_3644 & ~n_12532;
assign n_12534 =  n_6067 &  n_12533;
assign n_12535 = ~n_12530 & ~n_12534;
assign n_12536 =  x_1760 & ~n_12535;
assign n_12537 = ~x_1490 &  n_3256;
assign n_12538 =  n_12514 &  n_12537;
assign n_12539 = ~n_3718 & ~n_12538;
assign n_12540 = ~x_1756 & ~n_12539;
assign n_12541 = ~n_12536 & ~n_12540;
assign n_12542 =  n_12528 &  n_12541;
assign n_12543 =  x_1755 &  n_12542;
assign n_12544 = ~n_12524 & ~n_3719;
assign n_12545 = ~x_310 & ~n_12544;
assign n_12546 = ~x_1760 & ~x_1767;
assign n_12547 = ~n_12545 &  n_12546;
assign n_12548 = ~n_12542 & ~n_12547;
assign n_12549 = ~n_12543 & ~n_12548;
assign n_12550 =  x_1756 &  n_12528;
assign n_12551 =  x_1762 & ~n_12517;
assign n_12552 = ~n_12513 &  n_12551;
assign n_12553 =  x_1767 &  n_12552;
assign n_12554 =  x_1765 &  n_12529;
assign n_12555 =  n_6067 &  n_12554;
assign n_12556 =  x_1760 &  n_12555;
assign n_12557 =  n_12526 &  n_3636;
assign n_12558 =  n_12514 & ~n_12557;
assign n_12559 =  n_12523 & ~n_12529;
assign n_12560 =  x_310 &  x_1758;
assign n_12561 = ~n_12559 & ~n_12560;
assign n_12562 = ~n_12558 &  n_12561;
assign n_12563 = ~n_12556 &  n_12562;
assign n_12564 = ~n_12553 &  n_12563;
assign n_12565 = ~n_12542 & ~n_12564;
assign n_12566 = ~n_12550 & ~n_12565;
assign n_12567 =  x_1767 & ~n_12552;
assign n_12568 = ~x_1760 & ~n_12559;
assign n_12569 = ~n_12555 & ~n_12568;
assign n_12570 =  x_1758 & ~n_3644;
assign n_12571 = ~n_12557 & ~n_12570;
assign n_12572 = ~n_12569 &  n_12571;
assign n_12573 = ~n_12567 &  n_12572;
assign n_12574 = ~n_12542 & ~n_12573;
assign n_12575 =  x_1757 &  n_12542;
assign n_12576 = ~n_12574 & ~n_12575;
assign n_12577 =  n_12566 & ~n_12576;
assign n_12578 =  n_12549 &  n_12577;
assign n_12579 =  n_3636 &  n_12578;
assign n_12580 = ~n_12549 &  n_12576;
assign n_12581 =  n_12566 &  n_12580;
assign n_12582 = ~x_310 &  n_12581;
assign n_12583 = ~n_12566 & ~n_12576;
assign n_12584 =  x_310 &  n_12583;
assign n_12585 =  x_1768 &  n_12517;
assign n_12586 =  n_12584 &  n_12585;
assign n_12587 = ~n_12582 & ~n_12586;
assign n_12588 =  x_1489 & ~n_12587;
assign n_12589 = ~n_12517 &  n_12529;
assign n_12590 =  x_1760 &  n_12531;
assign n_12591 =  n_12589 &  n_12590;
assign n_12592 =  x_1765 & ~x_1766;
assign n_12593 =  n_12512 &  n_12592;
assign n_12594 = ~n_12530 & ~n_12593;
assign n_12595 =  n_6067 &  n_12523;
assign n_12596 = ~n_12594 &  n_12595;
assign n_12597 =  x_1767 &  n_12593;
assign n_12598 =  x_1761 & ~n_12597;
assign n_12599 = ~n_12596 &  n_12598;
assign n_12600 = ~n_12591 &  n_12599;
assign n_12601 = ~n_12588 &  n_12600;
assign n_12602 = ~n_12579 & ~n_12601;
assign n_12603 = ~x_1761 & ~n_12602;
assign n_12604 =  x_2440 &  n_12603;
assign n_12605 = ~x_2440 & ~n_12603;
assign n_12606 = ~n_12604 & ~n_12605;
assign n_12607 =  x_2439 &  n_3634;
assign n_12608 = ~x_2439 & ~n_3634;
assign n_12609 = ~n_12607 & ~n_12608;
assign n_12610 =  x_2438 &  n_3612;
assign n_12611 = ~x_2438 & ~n_3612;
assign n_12612 = ~n_12610 & ~n_12611;
assign n_12613 =  x_2437 &  n_3633;
assign n_12614 = ~x_2437 & ~n_3633;
assign n_12615 = ~n_12613 & ~n_12614;
assign n_12616 =  x_2436 &  n_3611;
assign n_12617 = ~x_2436 & ~n_3611;
assign n_12618 = ~n_12616 & ~n_12617;
assign n_12619 =  x_2435 &  n_3599;
assign n_12620 = ~x_2435 & ~n_3599;
assign n_12621 = ~n_12619 & ~n_12620;
assign n_12622 =  x_2434 & ~n_3570;
assign n_12623 = ~n_6010 & ~n_12622;
assign n_12624 =  x_2433 &  n_3569;
assign n_12625 = ~x_2433 & ~n_3569;
assign n_12626 = ~n_12624 & ~n_12625;
assign n_12627 = ~n_6067 &  n_12530;
assign n_12628 = ~n_12581 &  n_12627;
assign n_12629 = ~n_12578 & ~n_12628;
assign n_12630 = ~x_312 &  x_454;
assign n_12631 = ~x_312 &  x_456;
assign n_12632 = ~x_482 & ~x_483;
assign n_12633 = ~x_484 & ~x_485;
assign n_12634 =  n_12632 &  n_12633;
assign n_12635 = ~x_478 & ~x_479;
assign n_12636 = ~x_480 & ~x_481;
assign n_12637 =  n_12635 &  n_12636;
assign n_12638 = ~x_474 & ~x_475;
assign n_12639 = ~x_476 & ~x_477;
assign n_12640 =  n_12638 &  n_12639;
assign n_12641 =  n_12637 &  n_12640;
assign n_12642 =  n_12634 &  n_12641;
assign n_12643 = ~x_462 & ~x_463;
assign n_12644 = ~x_464 & ~x_465;
assign n_12645 =  n_12643 &  n_12644;
assign n_12646 = ~x_458 & ~x_459;
assign n_12647 = ~x_460 & ~x_461;
assign n_12648 =  n_12646 &  n_12647;
assign n_12649 =  n_12645 &  n_12648;
assign n_12650 = ~x_470 & ~x_471;
assign n_12651 = ~x_472 & ~x_473;
assign n_12652 =  n_12650 &  n_12651;
assign n_12653 = ~x_466 & ~x_467;
assign n_12654 = ~x_468 & ~x_469;
assign n_12655 =  n_12653 &  n_12654;
assign n_12656 =  n_12652 &  n_12655;
assign n_12657 =  n_12649 &  n_12656;
assign n_12658 =  n_12642 &  n_12657;
assign n_12659 = ~x_457 &  n_12658;
assign n_12660 =  n_12631 &  n_12659;
assign n_12661 = ~x_455 &  n_12660;
assign n_12662 =  n_12630 &  n_12661;
assign n_12663 = ~x_873 &  n_12662;
assign n_12664 =  x_455 &  n_12660;
assign n_12665 = ~n_12630 &  n_12664;
assign n_12666 = ~x_879 &  n_12665;
assign n_12667 = ~n_12663 & ~n_12666;
assign n_12668 =  n_12630 &  n_12664;
assign n_12669 = ~x_876 &  n_12668;
assign n_12670 = ~n_12630 &  n_12661;
assign n_12671 = ~x_875 &  n_12670;
assign n_12672 = ~n_12669 & ~n_12671;
assign n_12673 =  n_12667 &  n_12672;
assign n_12674 = ~x_456 &  x_457;
assign n_12675 =  n_12658 &  n_12674;
assign n_12676 = ~x_455 &  n_12675;
assign n_12677 = ~n_12630 &  n_12676;
assign n_12678 = ~x_869 &  n_12677;
assign n_12679 = ~x_312 &  x_455;
assign n_12680 =  n_12679 &  n_12675;
assign n_12681 = ~x_454 &  n_12680;
assign n_12682 = ~x_880 &  n_12681;
assign n_12683 = ~n_12678 & ~n_12682;
assign n_12684 =  n_12630 &  n_12676;
assign n_12685 = ~x_871 &  n_12684;
assign n_12686 =  x_454 &  n_12680;
assign n_12687 = ~x_870 &  n_12686;
assign n_12688 = ~n_12685 & ~n_12687;
assign n_12689 =  n_12683 &  n_12688;
assign n_12690 = ~n_12631 &  n_12659;
assign n_12691 =  n_12679 &  n_12690;
assign n_12692 =  x_454 &  n_12691;
assign n_12693 = ~x_872 &  n_12692;
assign n_12694 = ~n_12679 &  n_12690;
assign n_12695 = ~n_12630 &  n_12694;
assign n_12696 = ~x_878 &  n_12695;
assign n_12697 = ~n_12693 & ~n_12696;
assign n_12698 = ~x_454 &  n_12691;
assign n_12699 = ~x_874 &  n_12698;
assign n_12700 =  n_12630 &  n_12694;
assign n_12701 = ~x_877 &  n_12700;
assign n_12702 = ~n_12699 & ~n_12701;
assign n_12703 =  n_12697 &  n_12702;
assign n_12704 =  n_12689 &  n_12703;
assign n_12705 =  n_12673 &  n_12704;
assign n_12706 =  n_12629 &  n_12705;
assign n_12707 = ~x_1759 & ~n_12581;
assign n_12708 = ~n_12579 &  n_12707;
assign n_12709 =  x_2398 &  n_12578;
assign n_12710 = ~n_12708 & ~n_12709;
assign n_12711 = ~n_12706 &  n_12710;
assign n_12712 = ~x_2432 &  n_12708;
assign n_12713 = ~n_12711 & ~n_12712;
assign n_12714 =  x_2432 &  n_12713;
assign n_12715 = ~x_2432 & ~n_12713;
assign n_12716 = ~n_12714 & ~n_12715;
assign n_12717 = ~x_866 &  n_12698;
assign n_12718 = ~x_857 &  n_12665;
assign n_12719 = ~n_12717 & ~n_12718;
assign n_12720 = ~x_861 &  n_12662;
assign n_12721 = ~x_865 &  n_12692;
assign n_12722 = ~n_12720 & ~n_12721;
assign n_12723 =  n_12719 &  n_12722;
assign n_12724 = ~x_859 &  n_12677;
assign n_12725 = ~x_863 &  n_12684;
assign n_12726 = ~n_12724 & ~n_12725;
assign n_12727 = ~x_867 &  n_12681;
assign n_12728 = ~x_858 &  n_12686;
assign n_12729 = ~n_12727 & ~n_12728;
assign n_12730 =  n_12726 &  n_12729;
assign n_12731 = ~x_864 &  n_12700;
assign n_12732 = ~x_860 &  n_12668;
assign n_12733 = ~n_12731 & ~n_12732;
assign n_12734 = ~x_868 &  n_12670;
assign n_12735 = ~x_862 &  n_12695;
assign n_12736 = ~n_12734 & ~n_12735;
assign n_12737 =  n_12733 &  n_12736;
assign n_12738 =  n_12730 &  n_12737;
assign n_12739 =  n_12723 &  n_12738;
assign n_12740 =  n_12629 &  n_12739;
assign n_12741 =  x_2397 &  n_12578;
assign n_12742 = ~n_12708 & ~n_12741;
assign n_12743 = ~n_12740 &  n_12742;
assign n_12744 = ~x_2431 &  n_12708;
assign n_12745 = ~n_12743 & ~n_12744;
assign n_12746 =  x_2431 &  n_12745;
assign n_12747 = ~x_2431 & ~n_12745;
assign n_12748 = ~n_12746 & ~n_12747;
assign n_12749 = ~x_848 &  n_12665;
assign n_12750 = ~x_854 &  n_12670;
assign n_12751 = ~n_12749 & ~n_12750;
assign n_12752 = ~x_847 &  n_12695;
assign n_12753 = ~x_853 &  n_12700;
assign n_12754 = ~n_12752 & ~n_12753;
assign n_12755 =  n_12751 &  n_12754;
assign n_12756 = ~x_856 &  n_12686;
assign n_12757 = ~x_855 &  n_12677;
assign n_12758 = ~n_12756 & ~n_12757;
assign n_12759 = ~x_849 &  n_12684;
assign n_12760 = ~x_850 &  n_12681;
assign n_12761 = ~n_12759 & ~n_12760;
assign n_12762 =  n_12758 &  n_12761;
assign n_12763 = ~x_846 &  n_12662;
assign n_12764 = ~x_852 &  n_12668;
assign n_12765 = ~n_12763 & ~n_12764;
assign n_12766 = ~x_851 &  n_12698;
assign n_12767 = ~x_845 &  n_12692;
assign n_12768 = ~n_12766 & ~n_12767;
assign n_12769 =  n_12765 &  n_12768;
assign n_12770 =  n_12762 &  n_12769;
assign n_12771 =  n_12755 &  n_12770;
assign n_12772 =  n_12629 &  n_12771;
assign n_12773 =  x_2396 &  n_12578;
assign n_12774 = ~n_12708 & ~n_12773;
assign n_12775 = ~n_12772 &  n_12774;
assign n_12776 = ~x_2430 &  n_12708;
assign n_12777 = ~n_12775 & ~n_12776;
assign n_12778 =  x_2430 &  n_12777;
assign n_12779 = ~x_2430 & ~n_12777;
assign n_12780 = ~n_12778 & ~n_12779;
assign n_12781 = ~x_843 &  n_12695;
assign n_12782 = ~x_841 &  n_12665;
assign n_12783 = ~n_12781 & ~n_12782;
assign n_12784 = ~x_835 &  n_12670;
assign n_12785 = ~x_836 &  n_12700;
assign n_12786 = ~n_12784 & ~n_12785;
assign n_12787 =  n_12783 &  n_12786;
assign n_12788 = ~x_833 &  n_12684;
assign n_12789 = ~x_844 &  n_12677;
assign n_12790 = ~n_12788 & ~n_12789;
assign n_12791 = ~x_838 &  n_12681;
assign n_12792 = ~x_839 &  n_12686;
assign n_12793 = ~n_12791 & ~n_12792;
assign n_12794 =  n_12790 &  n_12793;
assign n_12795 = ~x_842 &  n_12668;
assign n_12796 = ~x_840 &  n_12698;
assign n_12797 = ~n_12795 & ~n_12796;
assign n_12798 = ~x_834 &  n_12662;
assign n_12799 = ~x_837 &  n_12692;
assign n_12800 = ~n_12798 & ~n_12799;
assign n_12801 =  n_12797 &  n_12800;
assign n_12802 =  n_12794 &  n_12801;
assign n_12803 =  n_12787 &  n_12802;
assign n_12804 =  n_12629 &  n_12803;
assign n_12805 =  x_2395 &  n_12578;
assign n_12806 = ~n_12708 & ~n_12805;
assign n_12807 = ~n_12804 &  n_12806;
assign n_12808 = ~x_2429 &  n_12708;
assign n_12809 = ~n_12807 & ~n_12808;
assign n_12810 =  x_2429 &  n_12809;
assign n_12811 = ~x_2429 & ~n_12809;
assign n_12812 = ~n_12810 & ~n_12811;
assign n_12813 = ~x_828 &  n_12692;
assign n_12814 = ~x_829 &  n_12700;
assign n_12815 = ~n_12813 & ~n_12814;
assign n_12816 = ~x_821 &  n_12695;
assign n_12817 = ~x_832 &  n_12668;
assign n_12818 = ~n_12816 & ~n_12817;
assign n_12819 =  n_12815 &  n_12818;
assign n_12820 = ~x_826 &  n_12677;
assign n_12821 = ~x_823 &  n_12681;
assign n_12822 = ~n_12820 & ~n_12821;
assign n_12823 = ~x_822 &  n_12686;
assign n_12824 = ~x_830 &  n_12684;
assign n_12825 = ~n_12823 & ~n_12824;
assign n_12826 =  n_12822 &  n_12825;
assign n_12827 = ~x_825 &  n_12665;
assign n_12828 = ~x_827 &  n_12698;
assign n_12829 = ~n_12827 & ~n_12828;
assign n_12830 = ~x_831 &  n_12670;
assign n_12831 = ~x_824 &  n_12662;
assign n_12832 = ~n_12830 & ~n_12831;
assign n_12833 =  n_12829 &  n_12832;
assign n_12834 =  n_12826 &  n_12833;
assign n_12835 =  n_12819 &  n_12834;
assign n_12836 =  n_12629 &  n_12835;
assign n_12837 =  x_2394 &  n_12578;
assign n_12838 = ~n_12708 & ~n_12837;
assign n_12839 = ~n_12836 &  n_12838;
assign n_12840 = ~x_2428 &  n_12708;
assign n_12841 = ~n_12839 & ~n_12840;
assign n_12842 =  x_2428 &  n_12841;
assign n_12843 = ~x_2428 & ~n_12841;
assign n_12844 = ~n_12842 & ~n_12843;
assign n_12845 = ~x_820 &  n_12665;
assign n_12846 = ~x_814 &  n_12662;
assign n_12847 = ~n_12845 & ~n_12846;
assign n_12848 = ~x_813 &  n_12692;
assign n_12849 = ~x_815 &  n_12698;
assign n_12850 = ~n_12848 & ~n_12849;
assign n_12851 =  n_12847 &  n_12850;
assign n_12852 = ~x_816 &  n_12677;
assign n_12853 = ~x_809 &  n_12684;
assign n_12854 = ~n_12852 & ~n_12853;
assign n_12855 = ~x_818 &  n_12686;
assign n_12856 = ~x_817 &  n_12681;
assign n_12857 = ~n_12855 & ~n_12856;
assign n_12858 =  n_12854 &  n_12857;
assign n_12859 = ~x_810 &  n_12700;
assign n_12860 = ~x_812 &  n_12695;
assign n_12861 = ~n_12859 & ~n_12860;
assign n_12862 = ~x_819 &  n_12670;
assign n_12863 = ~x_811 &  n_12668;
assign n_12864 = ~n_12862 & ~n_12863;
assign n_12865 =  n_12861 &  n_12864;
assign n_12866 =  n_12858 &  n_12865;
assign n_12867 =  n_12851 &  n_12866;
assign n_12868 =  n_12629 &  n_12867;
assign n_12869 =  x_2393 &  n_12578;
assign n_12870 = ~n_12708 & ~n_12869;
assign n_12871 = ~n_12868 &  n_12870;
assign n_12872 = ~x_2427 &  n_12708;
assign n_12873 = ~n_12871 & ~n_12872;
assign n_12874 =  x_2427 &  n_12873;
assign n_12875 = ~x_2427 & ~n_12873;
assign n_12876 = ~n_12874 & ~n_12875;
assign n_12877 = ~x_808 &  n_12670;
assign n_12878 = ~x_802 &  n_12662;
assign n_12879 = ~n_12877 & ~n_12878;
assign n_12880 = ~x_801 &  n_12665;
assign n_12881 = ~x_803 &  n_12700;
assign n_12882 = ~n_12880 & ~n_12881;
assign n_12883 =  n_12879 &  n_12882;
assign n_12884 = ~x_804 &  n_12677;
assign n_12885 = ~x_797 &  n_12681;
assign n_12886 = ~n_12884 & ~n_12885;
assign n_12887 = ~x_806 &  n_12686;
assign n_12888 = ~x_805 &  n_12684;
assign n_12889 = ~n_12887 & ~n_12888;
assign n_12890 =  n_12886 &  n_12889;
assign n_12891 = ~x_798 &  n_12668;
assign n_12892 = ~x_800 &  n_12698;
assign n_12893 = ~n_12891 & ~n_12892;
assign n_12894 = ~x_807 &  n_12695;
assign n_12895 = ~x_799 &  n_12692;
assign n_12896 = ~n_12894 & ~n_12895;
assign n_12897 =  n_12893 &  n_12896;
assign n_12898 =  n_12890 &  n_12897;
assign n_12899 =  n_12883 &  n_12898;
assign n_12900 =  n_12629 &  n_12899;
assign n_12901 =  x_2392 &  n_12578;
assign n_12902 = ~n_12708 & ~n_12901;
assign n_12903 = ~n_12900 &  n_12902;
assign n_12904 = ~x_2426 &  n_12708;
assign n_12905 = ~n_12903 & ~n_12904;
assign n_12906 =  x_2426 &  n_12905;
assign n_12907 = ~x_2426 & ~n_12905;
assign n_12908 = ~n_12906 & ~n_12907;
assign n_12909 = ~x_793 &  n_12692;
assign n_12910 = ~x_788 &  n_12698;
assign n_12911 = ~n_12909 & ~n_12910;
assign n_12912 = ~x_785 &  n_12668;
assign n_12913 = ~x_789 &  n_12662;
assign n_12914 = ~n_12912 & ~n_12913;
assign n_12915 =  n_12911 &  n_12914;
assign n_12916 = ~x_791 &  n_12686;
assign n_12917 = ~x_786 &  n_12677;
assign n_12918 = ~n_12916 & ~n_12917;
assign n_12919 = ~x_796 &  n_12684;
assign n_12920 = ~x_795 &  n_12681;
assign n_12921 = ~n_12919 & ~n_12920;
assign n_12922 =  n_12918 &  n_12921;
assign n_12923 = ~x_787 &  n_12700;
assign n_12924 = ~x_792 &  n_12665;
assign n_12925 = ~n_12923 & ~n_12924;
assign n_12926 = ~x_794 &  n_12670;
assign n_12927 = ~x_790 &  n_12695;
assign n_12928 = ~n_12926 & ~n_12927;
assign n_12929 =  n_12925 &  n_12928;
assign n_12930 =  n_12922 &  n_12929;
assign n_12931 =  n_12915 &  n_12930;
assign n_12932 =  n_12629 &  n_12931;
assign n_12933 =  x_2391 &  n_12578;
assign n_12934 = ~n_12708 & ~n_12933;
assign n_12935 = ~n_12932 &  n_12934;
assign n_12936 = ~x_2425 &  n_12708;
assign n_12937 = ~n_12935 & ~n_12936;
assign n_12938 =  x_2425 &  n_12937;
assign n_12939 = ~x_2425 & ~n_12937;
assign n_12940 = ~n_12938 & ~n_12939;
assign n_12941 = ~x_777 &  n_12662;
assign n_12942 = ~x_783 &  n_12665;
assign n_12943 = ~n_12941 & ~n_12942;
assign n_12944 = ~x_780 &  n_12700;
assign n_12945 = ~x_779 &  n_12670;
assign n_12946 = ~n_12944 & ~n_12945;
assign n_12947 =  n_12943 &  n_12946;
assign n_12948 = ~x_773 &  n_12677;
assign n_12949 = ~x_784 &  n_12681;
assign n_12950 = ~n_12948 & ~n_12949;
assign n_12951 = ~x_775 &  n_12684;
assign n_12952 = ~x_774 &  n_12686;
assign n_12953 = ~n_12951 & ~n_12952;
assign n_12954 =  n_12950 &  n_12953;
assign n_12955 = ~x_776 &  n_12692;
assign n_12956 = ~x_782 &  n_12668;
assign n_12957 = ~n_12955 & ~n_12956;
assign n_12958 = ~x_778 &  n_12698;
assign n_12959 = ~x_781 &  n_12695;
assign n_12960 = ~n_12958 & ~n_12959;
assign n_12961 =  n_12957 &  n_12960;
assign n_12962 =  n_12954 &  n_12961;
assign n_12963 =  n_12947 &  n_12962;
assign n_12964 =  n_12629 &  n_12963;
assign n_12965 =  x_2390 &  n_12578;
assign n_12966 = ~n_12708 & ~n_12965;
assign n_12967 = ~n_12964 &  n_12966;
assign n_12968 = ~x_2424 &  n_12708;
assign n_12969 = ~n_12967 & ~n_12968;
assign n_12970 =  x_2424 &  n_12969;
assign n_12971 = ~x_2424 & ~n_12969;
assign n_12972 = ~n_12970 & ~n_12971;
assign n_12973 = ~x_770 &  n_12692;
assign n_12974 = ~x_761 &  n_12700;
assign n_12975 = ~n_12973 & ~n_12974;
assign n_12976 = ~x_765 &  n_12662;
assign n_12977 = ~x_769 &  n_12695;
assign n_12978 = ~n_12976 & ~n_12977;
assign n_12979 =  n_12975 &  n_12978;
assign n_12980 = ~x_763 &  n_12684;
assign n_12981 = ~x_767 &  n_12681;
assign n_12982 = ~n_12980 & ~n_12981;
assign n_12983 = ~x_771 &  n_12677;
assign n_12984 = ~x_762 &  n_12686;
assign n_12985 = ~n_12983 & ~n_12984;
assign n_12986 =  n_12982 &  n_12985;
assign n_12987 = ~x_768 &  n_12670;
assign n_12988 = ~x_764 &  n_12668;
assign n_12989 = ~n_12987 & ~n_12988;
assign n_12990 = ~x_772 &  n_12698;
assign n_12991 = ~x_766 &  n_12665;
assign n_12992 = ~n_12990 & ~n_12991;
assign n_12993 =  n_12989 &  n_12992;
assign n_12994 =  n_12986 &  n_12993;
assign n_12995 =  n_12979 &  n_12994;
assign n_12996 =  n_12629 &  n_12995;
assign n_12997 =  x_2389 &  n_12578;
assign n_12998 = ~n_12708 & ~n_12997;
assign n_12999 = ~n_12996 &  n_12998;
assign n_13000 = ~x_2423 &  n_12708;
assign n_13001 = ~n_12999 & ~n_13000;
assign n_13002 =  x_2423 &  n_13001;
assign n_13003 = ~x_2423 & ~n_13001;
assign n_13004 = ~n_13002 & ~n_13003;
assign n_13005 = ~x_759 &  n_12665;
assign n_13006 = ~x_752 &  n_12700;
assign n_13007 = ~n_13005 & ~n_13006;
assign n_13008 = ~x_753 &  n_12668;
assign n_13009 = ~x_757 &  n_12692;
assign n_13010 = ~n_13008 & ~n_13009;
assign n_13011 =  n_13007 &  n_13010;
assign n_13012 = ~x_754 &  n_12677;
assign n_13013 = ~x_755 &  n_12681;
assign n_13014 = ~n_13012 & ~n_13013;
assign n_13015 = ~x_749 &  n_12686;
assign n_13016 = ~x_758 &  n_12684;
assign n_13017 = ~n_13015 & ~n_13016;
assign n_13018 =  n_13014 &  n_13017;
assign n_13019 = ~x_756 &  n_12695;
assign n_13020 = ~x_751 &  n_12662;
assign n_13021 = ~n_13019 & ~n_13020;
assign n_13022 = ~x_760 &  n_12670;
assign n_13023 = ~x_750 &  n_12698;
assign n_13024 = ~n_13022 & ~n_13023;
assign n_13025 =  n_13021 &  n_13024;
assign n_13026 =  n_13018 &  n_13025;
assign n_13027 =  n_13011 &  n_13026;
assign n_13028 =  n_12629 &  n_13027;
assign n_13029 =  x_2388 &  n_12578;
assign n_13030 = ~n_12708 & ~n_13029;
assign n_13031 = ~n_13028 &  n_13030;
assign n_13032 = ~x_2422 &  n_12708;
assign n_13033 = ~n_13031 & ~n_13032;
assign n_13034 =  x_2422 &  n_13033;
assign n_13035 = ~x_2422 & ~n_13033;
assign n_13036 = ~n_13034 & ~n_13035;
assign n_13037 = ~x_746 &  n_12670;
assign n_13038 = ~x_737 &  n_12692;
assign n_13039 = ~n_13037 & ~n_13038;
assign n_13040 = ~x_741 &  n_12665;
assign n_13041 = ~x_745 &  n_12698;
assign n_13042 = ~n_13040 & ~n_13041;
assign n_13043 =  n_13039 &  n_13042;
assign n_13044 = ~x_739 &  n_12677;
assign n_13045 = ~x_744 &  n_12686;
assign n_13046 = ~n_13044 & ~n_13045;
assign n_13047 = ~x_748 &  n_12681;
assign n_13048 = ~x_738 &  n_12684;
assign n_13049 = ~n_13047 & ~n_13048;
assign n_13050 =  n_13046 &  n_13049;
assign n_13051 = ~x_747 &  n_12695;
assign n_13052 = ~x_740 &  n_12662;
assign n_13053 = ~n_13051 & ~n_13052;
assign n_13054 = ~x_743 &  n_12668;
assign n_13055 = ~x_742 &  n_12700;
assign n_13056 = ~n_13054 & ~n_13055;
assign n_13057 =  n_13053 &  n_13056;
assign n_13058 =  n_13050 &  n_13057;
assign n_13059 =  n_13043 &  n_13058;
assign n_13060 =  n_12629 &  n_13059;
assign n_13061 =  x_2387 &  n_12578;
assign n_13062 = ~n_12708 & ~n_13061;
assign n_13063 = ~n_13060 &  n_13062;
assign n_13064 = ~x_2421 &  n_12708;
assign n_13065 = ~n_13063 & ~n_13064;
assign n_13066 =  x_2421 &  n_13065;
assign n_13067 = ~x_2421 & ~n_13065;
assign n_13068 = ~n_13066 & ~n_13067;
assign n_13069 = ~x_725 &  n_12692;
assign n_13070 = ~x_728 &  n_12670;
assign n_13071 = ~n_13069 & ~n_13070;
assign n_13072 = ~x_726 &  n_12665;
assign n_13073 = ~x_733 &  n_12698;
assign n_13074 = ~n_13072 & ~n_13073;
assign n_13075 =  n_13071 &  n_13074;
assign n_13076 = ~x_730 &  n_12681;
assign n_13077 = ~x_729 &  n_12686;
assign n_13078 = ~n_13076 & ~n_13077;
assign n_13079 = ~x_731 &  n_12684;
assign n_13080 = ~x_734 &  n_12677;
assign n_13081 = ~n_13079 & ~n_13080;
assign n_13082 =  n_13078 &  n_13081;
assign n_13083 = ~x_736 &  n_12695;
assign n_13084 = ~x_732 &  n_12662;
assign n_13085 = ~n_13083 & ~n_13084;
assign n_13086 = ~x_735 &  n_12700;
assign n_13087 = ~x_727 &  n_12668;
assign n_13088 = ~n_13086 & ~n_13087;
assign n_13089 =  n_13085 &  n_13088;
assign n_13090 =  n_13082 &  n_13089;
assign n_13091 =  n_13075 &  n_13090;
assign n_13092 =  n_12629 &  n_13091;
assign n_13093 =  x_2386 &  n_12578;
assign n_13094 = ~n_12708 & ~n_13093;
assign n_13095 = ~n_13092 &  n_13094;
assign n_13096 = ~x_2420 &  n_12708;
assign n_13097 = ~n_13095 & ~n_13096;
assign n_13098 =  x_2420 &  n_13097;
assign n_13099 = ~x_2420 & ~n_13097;
assign n_13100 = ~n_13098 & ~n_13099;
assign n_13101 = ~x_722 &  n_12670;
assign n_13102 = ~x_713 &  n_12700;
assign n_13103 = ~n_13101 & ~n_13102;
assign n_13104 = ~x_717 &  n_12692;
assign n_13105 = ~x_721 &  n_12695;
assign n_13106 = ~n_13104 & ~n_13105;
assign n_13107 =  n_13103 &  n_13106;
assign n_13108 = ~x_715 &  n_12686;
assign n_13109 = ~x_720 &  n_12684;
assign n_13110 = ~n_13108 & ~n_13109;
assign n_13111 = ~x_724 &  n_12677;
assign n_13112 = ~x_714 &  n_12681;
assign n_13113 = ~n_13111 & ~n_13112;
assign n_13114 =  n_13110 &  n_13113;
assign n_13115 = ~x_723 &  n_12698;
assign n_13116 = ~x_716 &  n_12668;
assign n_13117 = ~n_13115 & ~n_13116;
assign n_13118 = ~x_719 &  n_12665;
assign n_13119 = ~x_718 &  n_12662;
assign n_13120 = ~n_13118 & ~n_13119;
assign n_13121 =  n_13117 &  n_13120;
assign n_13122 =  n_13114 &  n_13121;
assign n_13123 =  n_13107 &  n_13122;
assign n_13124 =  n_12629 &  n_13123;
assign n_13125 =  x_2385 &  n_12578;
assign n_13126 = ~n_12708 & ~n_13125;
assign n_13127 = ~n_13124 &  n_13126;
assign n_13128 = ~x_2419 &  n_12708;
assign n_13129 = ~n_13127 & ~n_13128;
assign n_13130 =  x_2419 &  n_13129;
assign n_13131 = ~x_2419 & ~n_13129;
assign n_13132 = ~n_13130 & ~n_13131;
assign n_13133 = ~x_711 &  n_12692;
assign n_13134 = ~x_701 &  n_12700;
assign n_13135 = ~n_13133 & ~n_13134;
assign n_13136 = ~x_705 &  n_12698;
assign n_13137 = ~x_710 &  n_12670;
assign n_13138 = ~n_13136 & ~n_13137;
assign n_13139 =  n_13135 &  n_13138;
assign n_13140 = ~x_703 &  n_12684;
assign n_13141 = ~x_709 &  n_12677;
assign n_13142 = ~n_13140 & ~n_13141;
assign n_13143 = ~x_712 &  n_12686;
assign n_13144 = ~x_702 &  n_12681;
assign n_13145 = ~n_13143 & ~n_13144;
assign n_13146 =  n_13142 &  n_13145;
assign n_13147 = ~x_708 &  n_12668;
assign n_13148 = ~x_704 &  n_12662;
assign n_13149 = ~n_13147 & ~n_13148;
assign n_13150 = ~x_707 &  n_12665;
assign n_13151 = ~x_706 &  n_12695;
assign n_13152 = ~n_13150 & ~n_13151;
assign n_13153 =  n_13149 &  n_13152;
assign n_13154 =  n_13146 &  n_13153;
assign n_13155 =  n_13139 &  n_13154;
assign n_13156 =  n_12629 &  n_13155;
assign n_13157 =  x_2384 &  n_12578;
assign n_13158 = ~n_12708 & ~n_13157;
assign n_13159 = ~n_13156 &  n_13158;
assign n_13160 = ~x_2418 &  n_12708;
assign n_13161 = ~n_13159 & ~n_13160;
assign n_13162 =  x_2418 &  n_13161;
assign n_13163 = ~x_2418 & ~n_13161;
assign n_13164 = ~n_13162 & ~n_13163;
assign n_13165 = ~x_693 &  n_12668;
assign n_13166 = ~x_697 &  n_12700;
assign n_13167 = ~n_13165 & ~n_13166;
assign n_13168 = ~x_691 &  n_12692;
assign n_13169 = ~x_695 &  n_12670;
assign n_13170 = ~n_13168 & ~n_13169;
assign n_13171 =  n_13167 &  n_13170;
assign n_13172 = ~x_689 &  n_12681;
assign n_13173 = ~x_700 &  n_12677;
assign n_13174 = ~n_13172 & ~n_13173;
assign n_13175 = ~x_699 &  n_12684;
assign n_13176 = ~x_690 &  n_12686;
assign n_13177 = ~n_13175 & ~n_13176;
assign n_13178 =  n_13174 &  n_13177;
assign n_13179 = ~x_698 &  n_12665;
assign n_13180 = ~x_696 &  n_12698;
assign n_13181 = ~n_13179 & ~n_13180;
assign n_13182 = ~x_694 &  n_12662;
assign n_13183 = ~x_692 &  n_12695;
assign n_13184 = ~n_13182 & ~n_13183;
assign n_13185 =  n_13181 &  n_13184;
assign n_13186 =  n_13178 &  n_13185;
assign n_13187 =  n_13171 &  n_13186;
assign n_13188 =  n_12629 &  n_13187;
assign n_13189 =  x_2383 &  n_12578;
assign n_13190 = ~n_12708 & ~n_13189;
assign n_13191 = ~n_13188 &  n_13190;
assign n_13192 = ~x_2417 &  n_12708;
assign n_13193 = ~n_13191 & ~n_13192;
assign n_13194 =  x_2417 &  n_13193;
assign n_13195 = ~x_2417 & ~n_13193;
assign n_13196 = ~n_13194 & ~n_13195;
assign n_13197 = ~x_685 &  n_12668;
assign n_13198 = ~x_680 &  n_12670;
assign n_13199 = ~n_13197 & ~n_13198;
assign n_13200 = ~x_677 &  n_12700;
assign n_13201 = ~x_681 &  n_12662;
assign n_13202 = ~n_13200 & ~n_13201;
assign n_13203 =  n_13199 &  n_13202;
assign n_13204 = ~x_683 &  n_12686;
assign n_13205 = ~x_678 &  n_12684;
assign n_13206 = ~n_13204 & ~n_13205;
assign n_13207 = ~x_688 &  n_12681;
assign n_13208 = ~x_687 &  n_12677;
assign n_13209 = ~n_13207 & ~n_13208;
assign n_13210 =  n_13206 &  n_13209;
assign n_13211 = ~x_679 &  n_12665;
assign n_13212 = ~x_684 &  n_12695;
assign n_13213 = ~n_13211 & ~n_13212;
assign n_13214 = ~x_686 &  n_12692;
assign n_13215 = ~x_682 &  n_12698;
assign n_13216 = ~n_13214 & ~n_13215;
assign n_13217 =  n_13213 &  n_13216;
assign n_13218 =  n_13210 &  n_13217;
assign n_13219 =  n_13203 &  n_13218;
assign n_13220 =  n_12629 &  n_13219;
assign n_13221 =  x_2382 &  n_12578;
assign n_13222 = ~n_12708 & ~n_13221;
assign n_13223 = ~n_13220 &  n_13222;
assign n_13224 = ~x_2416 &  n_12708;
assign n_13225 = ~n_13223 & ~n_13224;
assign n_13226 =  x_2416 &  n_13225;
assign n_13227 = ~x_2416 & ~n_13225;
assign n_13228 = ~n_13226 & ~n_13227;
assign n_13229 = ~x_669 &  n_12698;
assign n_13230 = ~x_673 &  n_12700;
assign n_13231 = ~n_13229 & ~n_13230;
assign n_13232 = ~x_671 &  n_12670;
assign n_13233 = ~x_672 &  n_12695;
assign n_13234 = ~n_13232 & ~n_13233;
assign n_13235 =  n_13231 &  n_13234;
assign n_13236 = ~x_665 &  n_12684;
assign n_13237 = ~x_676 &  n_12681;
assign n_13238 = ~n_13236 & ~n_13237;
assign n_13239 = ~x_675 &  n_12677;
assign n_13240 = ~x_667 &  n_12686;
assign n_13241 = ~n_13239 & ~n_13240;
assign n_13242 =  n_13238 &  n_13241;
assign n_13243 = ~x_674 &  n_12665;
assign n_13244 = ~x_670 &  n_12692;
assign n_13245 = ~n_13243 & ~n_13244;
assign n_13246 = ~x_666 &  n_12662;
assign n_13247 = ~x_668 &  n_12668;
assign n_13248 = ~n_13246 & ~n_13247;
assign n_13249 =  n_13245 &  n_13248;
assign n_13250 =  n_13242 &  n_13249;
assign n_13251 =  n_13235 &  n_13250;
assign n_13252 =  n_12629 &  n_13251;
assign n_13253 =  x_2381 &  n_12578;
assign n_13254 = ~n_12708 & ~n_13253;
assign n_13255 = ~n_13252 &  n_13254;
assign n_13256 = ~x_2415 &  n_12708;
assign n_13257 = ~n_13255 & ~n_13256;
assign n_13258 =  x_2415 &  n_13257;
assign n_13259 = ~x_2415 & ~n_13257;
assign n_13260 = ~n_13258 & ~n_13259;
assign n_13261 = ~x_660 &  n_12662;
assign n_13262 = ~x_661 &  n_12700;
assign n_13263 = ~n_13261 & ~n_13262;
assign n_13264 = ~x_653 &  n_12698;
assign n_13265 = ~x_664 &  n_12670;
assign n_13266 = ~n_13264 & ~n_13265;
assign n_13267 =  n_13263 &  n_13266;
assign n_13268 = ~x_658 &  n_12686;
assign n_13269 = ~x_655 &  n_12684;
assign n_13270 = ~n_13268 & ~n_13269;
assign n_13271 = ~x_654 &  n_12681;
assign n_13272 = ~x_662 &  n_12677;
assign n_13273 = ~n_13271 & ~n_13272;
assign n_13274 =  n_13270 &  n_13273;
assign n_13275 = ~x_657 &  n_12695;
assign n_13276 = ~x_659 &  n_12692;
assign n_13277 = ~n_13275 & ~n_13276;
assign n_13278 = ~x_663 &  n_12668;
assign n_13279 = ~x_656 &  n_12665;
assign n_13280 = ~n_13278 & ~n_13279;
assign n_13281 =  n_13277 &  n_13280;
assign n_13282 =  n_13274 &  n_13281;
assign n_13283 =  n_13267 &  n_13282;
assign n_13284 =  n_12629 &  n_13283;
assign n_13285 =  x_2380 &  n_12578;
assign n_13286 = ~n_12708 & ~n_13285;
assign n_13287 = ~n_13284 &  n_13286;
assign n_13288 = ~x_2414 &  n_12708;
assign n_13289 = ~n_13287 & ~n_13288;
assign n_13290 =  x_2414 &  n_13289;
assign n_13291 = ~x_2414 & ~n_13289;
assign n_13292 = ~n_13290 & ~n_13291;
assign n_13293 = ~x_652 &  n_12700;
assign n_13294 = ~x_646 &  n_12665;
assign n_13295 = ~n_13293 & ~n_13294;
assign n_13296 = ~x_645 &  n_12698;
assign n_13297 = ~x_647 &  n_12692;
assign n_13298 = ~n_13296 & ~n_13297;
assign n_13299 =  n_13295 &  n_13298;
assign n_13300 = ~x_648 &  n_12684;
assign n_13301 = ~x_641 &  n_12686;
assign n_13302 = ~n_13300 & ~n_13301;
assign n_13303 = ~x_650 &  n_12677;
assign n_13304 = ~x_649 &  n_12681;
assign n_13305 = ~n_13303 & ~n_13304;
assign n_13306 =  n_13302 &  n_13305;
assign n_13307 = ~x_642 &  n_12668;
assign n_13308 = ~x_644 &  n_12695;
assign n_13309 = ~n_13307 & ~n_13308;
assign n_13310 = ~x_651 &  n_12670;
assign n_13311 = ~x_643 &  n_12662;
assign n_13312 = ~n_13310 & ~n_13311;
assign n_13313 =  n_13309 &  n_13312;
assign n_13314 =  n_13306 &  n_13313;
assign n_13315 =  n_13299 &  n_13314;
assign n_13316 =  n_12629 &  n_13315;
assign n_13317 =  x_2379 &  n_12578;
assign n_13318 = ~n_12708 & ~n_13317;
assign n_13319 = ~n_13316 &  n_13318;
assign n_13320 = ~x_2413 &  n_12708;
assign n_13321 = ~n_13319 & ~n_13320;
assign n_13322 =  x_2413 &  n_13321;
assign n_13323 = ~x_2413 & ~n_13321;
assign n_13324 = ~n_13322 & ~n_13323;
assign n_13325 = ~x_636 &  n_12700;
assign n_13326 = ~x_637 &  n_12692;
assign n_13327 = ~n_13325 & ~n_13326;
assign n_13328 = ~x_629 &  n_12698;
assign n_13329 = ~x_640 &  n_12695;
assign n_13330 = ~n_13328 & ~n_13329;
assign n_13331 =  n_13327 &  n_13330;
assign n_13332 = ~x_634 &  n_12677;
assign n_13333 = ~x_631 &  n_12684;
assign n_13334 = ~n_13332 & ~n_13333;
assign n_13335 = ~x_630 &  n_12681;
assign n_13336 = ~x_638 &  n_12686;
assign n_13337 = ~n_13335 & ~n_13336;
assign n_13338 =  n_13334 &  n_13337;
assign n_13339 = ~x_633 &  n_12665;
assign n_13340 = ~x_635 &  n_12670;
assign n_13341 = ~n_13339 & ~n_13340;
assign n_13342 = ~x_639 &  n_12662;
assign n_13343 = ~x_632 &  n_12668;
assign n_13344 = ~n_13342 & ~n_13343;
assign n_13345 =  n_13341 &  n_13344;
assign n_13346 =  n_13338 &  n_13345;
assign n_13347 =  n_13331 &  n_13346;
assign n_13348 =  n_12629 &  n_13347;
assign n_13349 =  x_2378 &  n_12578;
assign n_13350 = ~n_12708 & ~n_13349;
assign n_13351 = ~n_13348 &  n_13350;
assign n_13352 = ~x_2412 &  n_12708;
assign n_13353 = ~n_13351 & ~n_13352;
assign n_13354 =  x_2412 &  n_13353;
assign n_13355 = ~x_2412 & ~n_13353;
assign n_13356 = ~n_13354 & ~n_13355;
assign n_13357 = ~x_624 &  n_12662;
assign n_13358 = ~x_622 &  n_12668;
assign n_13359 = ~n_13357 & ~n_13358;
assign n_13360 = ~x_625 &  n_12695;
assign n_13361 = ~x_618 &  n_12670;
assign n_13362 = ~n_13360 & ~n_13361;
assign n_13363 =  n_13359 &  n_13362;
assign n_13364 = ~x_620 &  n_12686;
assign n_13365 = ~x_619 &  n_12681;
assign n_13366 = ~n_13364 & ~n_13365;
assign n_13367 = ~x_627 &  n_12684;
assign n_13368 = ~x_628 &  n_12677;
assign n_13369 = ~n_13367 & ~n_13368;
assign n_13370 =  n_13366 &  n_13369;
assign n_13371 = ~x_626 &  n_12700;
assign n_13372 = ~x_623 &  n_12665;
assign n_13373 = ~n_13371 & ~n_13372;
assign n_13374 = ~x_621 &  n_12692;
assign n_13375 = ~x_617 &  n_12698;
assign n_13376 = ~n_13374 & ~n_13375;
assign n_13377 =  n_13373 &  n_13376;
assign n_13378 =  n_13370 &  n_13377;
assign n_13379 =  n_13363 &  n_13378;
assign n_13380 =  n_12629 &  n_13379;
assign n_13381 =  x_2377 &  n_12578;
assign n_13382 = ~n_12708 & ~n_13381;
assign n_13383 = ~n_13380 &  n_13382;
assign n_13384 = ~x_2411 &  n_12708;
assign n_13385 = ~n_13383 & ~n_13384;
assign n_13386 =  x_2411 &  n_13385;
assign n_13387 = ~x_2411 & ~n_13385;
assign n_13388 = ~n_13386 & ~n_13387;
assign n_13389 = ~x_612 &  n_12668;
assign n_13390 = ~x_610 &  n_12662;
assign n_13391 = ~n_13389 & ~n_13390;
assign n_13392 = ~x_613 &  n_12665;
assign n_13393 = ~x_606 &  n_12695;
assign n_13394 = ~n_13392 & ~n_13393;
assign n_13395 =  n_13391 &  n_13394;
assign n_13396 = ~x_607 &  n_12681;
assign n_13397 = ~x_605 &  n_12686;
assign n_13398 = ~n_13396 & ~n_13397;
assign n_13399 = ~x_608 &  n_12677;
assign n_13400 = ~x_616 &  n_12684;
assign n_13401 = ~n_13399 & ~n_13400;
assign n_13402 =  n_13398 &  n_13401;
assign n_13403 = ~x_614 &  n_12692;
assign n_13404 = ~x_615 &  n_12670;
assign n_13405 = ~n_13403 & ~n_13404;
assign n_13406 = ~x_611 &  n_12698;
assign n_13407 = ~x_609 &  n_12700;
assign n_13408 = ~n_13406 & ~n_13407;
assign n_13409 =  n_13405 &  n_13408;
assign n_13410 =  n_13402 &  n_13409;
assign n_13411 =  n_13395 &  n_13410;
assign n_13412 =  n_12629 &  n_13411;
assign n_13413 =  x_2376 &  n_12578;
assign n_13414 = ~n_12708 & ~n_13413;
assign n_13415 = ~n_13412 &  n_13414;
assign n_13416 = ~x_2410 &  n_12708;
assign n_13417 = ~n_13415 & ~n_13416;
assign n_13418 =  x_2410 &  n_13417;
assign n_13419 = ~x_2410 & ~n_13417;
assign n_13420 = ~n_13418 & ~n_13419;
assign n_13421 = ~x_598 &  n_12700;
assign n_13422 = ~x_602 &  n_12662;
assign n_13423 = ~n_13421 & ~n_13422;
assign n_13424 = ~x_604 &  n_12698;
assign n_13425 = ~x_603 &  n_12665;
assign n_13426 = ~n_13424 & ~n_13425;
assign n_13427 =  n_13423 &  n_13426;
assign n_13428 = ~x_593 &  n_12684;
assign n_13429 = ~x_595 &  n_12677;
assign n_13430 = ~n_13428 & ~n_13429;
assign n_13431 = ~x_594 &  n_12681;
assign n_13432 = ~x_601 &  n_12686;
assign n_13433 = ~n_13431 & ~n_13432;
assign n_13434 =  n_13430 &  n_13433;
assign n_13435 = ~x_597 &  n_12692;
assign n_13436 = ~x_596 &  n_12670;
assign n_13437 = ~n_13435 & ~n_13436;
assign n_13438 = ~x_599 &  n_12668;
assign n_13439 = ~x_600 &  n_12695;
assign n_13440 = ~n_13438 & ~n_13439;
assign n_13441 =  n_13437 &  n_13440;
assign n_13442 =  n_13434 &  n_13441;
assign n_13443 =  n_13427 &  n_13442;
assign n_13444 =  n_12629 &  n_13443;
assign n_13445 =  x_2375 &  n_12578;
assign n_13446 = ~n_12708 & ~n_13445;
assign n_13447 = ~n_13444 &  n_13446;
assign n_13448 = ~x_2409 &  n_12708;
assign n_13449 = ~n_13447 & ~n_13448;
assign n_13450 =  x_2409 &  n_13449;
assign n_13451 = ~x_2409 & ~n_13449;
assign n_13452 = ~n_13450 & ~n_13451;
assign n_13453 = ~x_590 &  n_12662;
assign n_13454 = ~x_581 &  n_12668;
assign n_13455 = ~n_13453 & ~n_13454;
assign n_13456 = ~x_585 &  n_12670;
assign n_13457 = ~x_589 &  n_12698;
assign n_13458 = ~n_13456 & ~n_13457;
assign n_13459 =  n_13455 &  n_13458;
assign n_13460 = ~x_583 &  n_12686;
assign n_13461 = ~x_587 &  n_12681;
assign n_13462 = ~n_13460 & ~n_13461;
assign n_13463 = ~x_591 &  n_12677;
assign n_13464 = ~x_582 &  n_12684;
assign n_13465 = ~n_13463 & ~n_13464;
assign n_13466 =  n_13462 &  n_13465;
assign n_13467 = ~x_588 &  n_12692;
assign n_13468 = ~x_584 &  n_12695;
assign n_13469 = ~n_13467 & ~n_13468;
assign n_13470 = ~x_592 &  n_12700;
assign n_13471 = ~x_586 &  n_12665;
assign n_13472 = ~n_13470 & ~n_13471;
assign n_13473 =  n_13469 &  n_13472;
assign n_13474 =  n_13466 &  n_13473;
assign n_13475 =  n_13459 &  n_13474;
assign n_13476 =  n_12629 &  n_13475;
assign n_13477 =  x_2374 &  n_12578;
assign n_13478 = ~n_12708 & ~n_13477;
assign n_13479 = ~n_13476 &  n_13478;
assign n_13480 = ~x_2408 &  n_12708;
assign n_13481 = ~n_13479 & ~n_13480;
assign n_13482 =  x_2408 &  n_13481;
assign n_13483 = ~x_2408 & ~n_13481;
assign n_13484 = ~n_13482 & ~n_13483;
assign n_13485 = ~x_576 &  n_12700;
assign n_13486 = ~x_577 &  n_12692;
assign n_13487 = ~n_13485 & ~n_13486;
assign n_13488 = ~x_569 &  n_12698;
assign n_13489 = ~x_580 &  n_12695;
assign n_13490 = ~n_13488 & ~n_13489;
assign n_13491 =  n_13487 &  n_13490;
assign n_13492 = ~x_574 &  n_12677;
assign n_13493 = ~x_571 &  n_12684;
assign n_13494 = ~n_13492 & ~n_13493;
assign n_13495 = ~x_570 &  n_12681;
assign n_13496 = ~x_578 &  n_12686;
assign n_13497 = ~n_13495 & ~n_13496;
assign n_13498 =  n_13494 &  n_13497;
assign n_13499 = ~x_573 &  n_12665;
assign n_13500 = ~x_575 &  n_12670;
assign n_13501 = ~n_13499 & ~n_13500;
assign n_13502 = ~x_579 &  n_12662;
assign n_13503 = ~x_572 &  n_12668;
assign n_13504 = ~n_13502 & ~n_13503;
assign n_13505 =  n_13501 &  n_13504;
assign n_13506 =  n_13498 &  n_13505;
assign n_13507 =  n_13491 &  n_13506;
assign n_13508 =  n_12629 &  n_13507;
assign n_13509 =  x_2373 &  n_12578;
assign n_13510 = ~n_12708 & ~n_13509;
assign n_13511 = ~n_13508 &  n_13510;
assign n_13512 = ~x_2407 &  n_12708;
assign n_13513 = ~n_13511 & ~n_13512;
assign n_13514 =  x_2407 &  n_13513;
assign n_13515 = ~x_2407 & ~n_13513;
assign n_13516 = ~n_13514 & ~n_13515;
assign n_13517 = ~x_560 &  n_12700;
assign n_13518 = ~x_566 &  n_12662;
assign n_13519 = ~n_13517 & ~n_13518;
assign n_13520 = ~x_568 &  n_12692;
assign n_13521 = ~x_567 &  n_12668;
assign n_13522 = ~n_13520 & ~n_13521;
assign n_13523 =  n_13519 &  n_13522;
assign n_13524 = ~x_557 &  n_12686;
assign n_13525 = ~x_564 &  n_12681;
assign n_13526 = ~n_13524 & ~n_13525;
assign n_13527 = ~x_561 &  n_12677;
assign n_13528 = ~x_562 &  n_12684;
assign n_13529 = ~n_13527 & ~n_13528;
assign n_13530 =  n_13526 &  n_13529;
assign n_13531 = ~x_563 &  n_12665;
assign n_13532 = ~x_559 &  n_12695;
assign n_13533 = ~n_13531 & ~n_13532;
assign n_13534 = ~x_558 &  n_12698;
assign n_13535 = ~x_565 &  n_12670;
assign n_13536 = ~n_13534 & ~n_13535;
assign n_13537 =  n_13533 &  n_13536;
assign n_13538 =  n_13530 &  n_13537;
assign n_13539 =  n_13523 &  n_13538;
assign n_13540 =  n_12629 &  n_13539;
assign n_13541 =  x_2372 &  n_12578;
assign n_13542 = ~n_12708 & ~n_13541;
assign n_13543 = ~n_13540 &  n_13542;
assign n_13544 = ~x_2406 &  n_12708;
assign n_13545 = ~n_13543 & ~n_13544;
assign n_13546 =  x_2406 &  n_13545;
assign n_13547 = ~x_2406 & ~n_13545;
assign n_13548 = ~n_13546 & ~n_13547;
assign n_13549 = ~x_555 &  n_12692;
assign n_13550 = ~x_548 &  n_12700;
assign n_13551 = ~n_13549 & ~n_13550;
assign n_13552 = ~x_546 &  n_12698;
assign n_13553 = ~x_552 &  n_12670;
assign n_13554 = ~n_13552 & ~n_13553;
assign n_13555 =  n_13551 &  n_13554;
assign n_13556 = ~x_550 &  n_12684;
assign n_13557 = ~x_549 &  n_12686;
assign n_13558 = ~n_13556 & ~n_13557;
assign n_13559 = ~x_545 &  n_12677;
assign n_13560 = ~x_551 &  n_12681;
assign n_13561 = ~n_13559 & ~n_13560;
assign n_13562 =  n_13558 &  n_13561;
assign n_13563 = ~x_554 &  n_12668;
assign n_13564 = ~x_553 &  n_12662;
assign n_13565 = ~n_13563 & ~n_13564;
assign n_13566 = ~x_556 &  n_12665;
assign n_13567 = ~x_547 &  n_12695;
assign n_13568 = ~n_13566 & ~n_13567;
assign n_13569 =  n_13565 &  n_13568;
assign n_13570 =  n_13562 &  n_13569;
assign n_13571 =  n_13555 &  n_13570;
assign n_13572 =  n_12629 &  n_13571;
assign n_13573 =  x_2371 &  n_12578;
assign n_13574 = ~n_12708 & ~n_13573;
assign n_13575 = ~n_13572 &  n_13574;
assign n_13576 = ~x_2405 &  n_12708;
assign n_13577 = ~n_13575 & ~n_13576;
assign n_13578 =  x_2405 &  n_13577;
assign n_13579 = ~x_2405 & ~n_13577;
assign n_13580 = ~n_13578 & ~n_13579;
assign n_13581 = ~x_536 &  n_12698;
assign n_13582 = ~x_542 &  n_12700;
assign n_13583 = ~n_13581 & ~n_13582;
assign n_13584 = ~x_544 &  n_12670;
assign n_13585 = ~x_543 &  n_12695;
assign n_13586 = ~n_13584 & ~n_13585;
assign n_13587 =  n_13583 &  n_13586;
assign n_13588 = ~x_533 &  n_12677;
assign n_13589 = ~x_540 &  n_12681;
assign n_13590 = ~n_13588 & ~n_13589;
assign n_13591 = ~x_537 &  n_12684;
assign n_13592 = ~x_538 &  n_12686;
assign n_13593 = ~n_13591 & ~n_13592;
assign n_13594 =  n_13590 &  n_13593;
assign n_13595 = ~x_539 &  n_12665;
assign n_13596 = ~x_535 &  n_12668;
assign n_13597 = ~n_13595 & ~n_13596;
assign n_13598 = ~x_534 &  n_12692;
assign n_13599 = ~x_541 &  n_12662;
assign n_13600 = ~n_13598 & ~n_13599;
assign n_13601 =  n_13597 &  n_13600;
assign n_13602 =  n_13594 &  n_13601;
assign n_13603 =  n_13587 &  n_13602;
assign n_13604 =  n_12629 &  n_13603;
assign n_13605 =  x_2370 &  n_12578;
assign n_13606 = ~n_12708 & ~n_13605;
assign n_13607 = ~n_13604 &  n_13606;
assign n_13608 = ~x_2404 &  n_12708;
assign n_13609 = ~n_13607 & ~n_13608;
assign n_13610 =  x_2404 &  n_13609;
assign n_13611 = ~x_2404 & ~n_13609;
assign n_13612 = ~n_13610 & ~n_13611;
assign n_13613 = ~x_525 &  n_12698;
assign n_13614 = ~x_529 &  n_12692;
assign n_13615 = ~n_13613 & ~n_13614;
assign n_13616 = ~x_523 &  n_12695;
assign n_13617 = ~x_527 &  n_12670;
assign n_13618 = ~n_13616 & ~n_13617;
assign n_13619 =  n_13615 &  n_13618;
assign n_13620 = ~x_521 &  n_12681;
assign n_13621 = ~x_532 &  n_12686;
assign n_13622 = ~n_13620 & ~n_13621;
assign n_13623 = ~x_531 &  n_12677;
assign n_13624 = ~x_522 &  n_12684;
assign n_13625 = ~n_13623 & ~n_13624;
assign n_13626 =  n_13622 &  n_13625;
assign n_13627 = ~x_530 &  n_12668;
assign n_13628 = ~x_528 &  n_12665;
assign n_13629 = ~n_13627 & ~n_13628;
assign n_13630 = ~x_526 &  n_12700;
assign n_13631 = ~x_524 &  n_12662;
assign n_13632 = ~n_13630 & ~n_13631;
assign n_13633 =  n_13629 &  n_13632;
assign n_13634 =  n_13626 &  n_13633;
assign n_13635 =  n_13619 &  n_13634;
assign n_13636 =  n_12629 &  n_13635;
assign n_13637 =  x_2369 &  n_12578;
assign n_13638 = ~n_12708 & ~n_13637;
assign n_13639 = ~n_13636 &  n_13638;
assign n_13640 = ~x_2403 &  n_12708;
assign n_13641 = ~n_13639 & ~n_13640;
assign n_13642 =  x_2403 &  n_13641;
assign n_13643 = ~x_2403 & ~n_13641;
assign n_13644 = ~n_13642 & ~n_13643;
assign n_13645 = ~x_518 &  n_12700;
assign n_13646 = ~x_509 &  n_12698;
assign n_13647 = ~n_13645 & ~n_13646;
assign n_13648 = ~x_513 &  n_12695;
assign n_13649 = ~x_517 &  n_12670;
assign n_13650 = ~n_13648 & ~n_13649;
assign n_13651 =  n_13647 &  n_13650;
assign n_13652 = ~x_511 &  n_12677;
assign n_13653 = ~x_516 &  n_12686;
assign n_13654 = ~n_13652 & ~n_13653;
assign n_13655 = ~x_520 &  n_12681;
assign n_13656 = ~x_510 &  n_12684;
assign n_13657 = ~n_13655 & ~n_13656;
assign n_13658 =  n_13654 &  n_13657;
assign n_13659 = ~x_519 &  n_12692;
assign n_13660 = ~x_512 &  n_12662;
assign n_13661 = ~n_13659 & ~n_13660;
assign n_13662 = ~x_515 &  n_12668;
assign n_13663 = ~x_514 &  n_12665;
assign n_13664 = ~n_13662 & ~n_13663;
assign n_13665 =  n_13661 &  n_13664;
assign n_13666 =  n_13658 &  n_13665;
assign n_13667 =  n_13651 &  n_13666;
assign n_13668 =  n_12629 &  n_13667;
assign n_13669 =  x_2368 &  n_12578;
assign n_13670 = ~n_12708 & ~n_13669;
assign n_13671 = ~n_13668 &  n_13670;
assign n_13672 = ~x_2402 &  n_12708;
assign n_13673 = ~n_13671 & ~n_13672;
assign n_13674 =  x_2402 &  n_13673;
assign n_13675 = ~x_2402 & ~n_13673;
assign n_13676 = ~n_13674 & ~n_13675;
assign n_13677 = ~x_499 &  n_12670;
assign n_13678 = ~x_506 &  n_12695;
assign n_13679 = ~n_13677 & ~n_13678;
assign n_13680 = ~x_501 &  n_12665;
assign n_13681 = ~x_498 &  n_12698;
assign n_13682 = ~n_13680 & ~n_13681;
assign n_13683 =  n_13679 &  n_13682;
assign n_13684 = ~x_497 &  n_12684;
assign n_13685 = ~x_508 &  n_12681;
assign n_13686 = ~n_13684 & ~n_13685;
assign n_13687 = ~x_502 &  n_12677;
assign n_13688 = ~x_505 &  n_12686;
assign n_13689 = ~n_13687 & ~n_13688;
assign n_13690 =  n_13686 &  n_13689;
assign n_13691 = ~x_503 &  n_12692;
assign n_13692 = ~x_500 &  n_12668;
assign n_13693 = ~n_13691 & ~n_13692;
assign n_13694 = ~x_504 &  n_12662;
assign n_13695 = ~x_507 &  n_12700;
assign n_13696 = ~n_13694 & ~n_13695;
assign n_13697 =  n_13693 &  n_13696;
assign n_13698 =  n_13690 &  n_13697;
assign n_13699 =  n_13683 &  n_13698;
assign n_13700 =  n_12629 &  n_13699;
assign n_13701 =  x_2367 &  n_12578;
assign n_13702 = ~n_12708 & ~n_13701;
assign n_13703 = ~n_13700 &  n_13702;
assign n_13704 = ~x_2401 &  n_12708;
assign n_13705 = ~n_13703 & ~n_13704;
assign n_13706 =  x_2401 &  n_13705;
assign n_13707 = ~x_2401 & ~n_13705;
assign n_13708 = ~n_13706 & ~n_13707;
assign n_13709 = ~x_489 &  n_12662;
assign n_13710 = ~x_494 &  n_12692;
assign n_13711 = ~n_13709 & ~n_13710;
assign n_13712 = ~x_495 &  n_12668;
assign n_13713 = ~x_488 &  n_12695;
assign n_13714 = ~n_13712 & ~n_13713;
assign n_13715 =  n_13711 &  n_13714;
assign n_13716 = ~x_492 &  n_12677;
assign n_13717 = ~x_487 &  n_12681;
assign n_13718 = ~n_13716 & ~n_13717;
assign n_13719 = ~x_486 &  n_12686;
assign n_13720 = ~x_496 &  n_12684;
assign n_13721 = ~n_13719 & ~n_13720;
assign n_13722 =  n_13718 &  n_13721;
assign n_13723 = ~x_493 &  n_12665;
assign n_13724 = ~x_491 &  n_12670;
assign n_13725 = ~n_13723 & ~n_13724;
assign n_13726 = ~x_490 &  n_12698;
assign n_13727 = ~x_453 &  n_12700;
assign n_13728 = ~n_13726 & ~n_13727;
assign n_13729 =  n_13725 &  n_13728;
assign n_13730 =  n_13722 &  n_13729;
assign n_13731 =  n_13715 &  n_13730;
assign n_13732 =  n_12629 &  n_13731;
assign n_13733 = ~x_2366 &  n_12578;
assign n_13734 = ~n_13733 & ~n_12708;
assign n_13735 = ~n_13732 &  n_13734;
assign n_13736 =  x_2400 &  n_12708;
assign n_13737 = ~n_13735 & ~n_13736;
assign n_13738 =  x_2400 & ~n_13737;
assign n_13739 = ~x_2400 &  n_13737;
assign n_13740 = ~n_13738 & ~n_13739;
assign n_13741 =  n_12529 &  n_12578;
assign n_13742 =  x_1759 &  n_12592;
assign n_13743 =  n_12529 &  n_13742;
assign n_13744 =  x_2399 & ~n_13743;
assign n_13745 = ~n_13741 & ~n_13744;
assign n_13746 =  x_2399 & ~n_13745;
assign n_13747 = ~x_2399 &  n_13745;
assign n_13748 = ~n_13746 & ~n_13747;
assign n_13749 =  x_434 &  n_3307;
assign n_13750 =  x_2398 &  n_3308;
assign n_13751 = ~n_13749 & ~n_13750;
assign n_13752 =  x_2398 & ~n_13751;
assign n_13753 = ~x_2398 &  n_13751;
assign n_13754 = ~n_13752 & ~n_13753;
assign n_13755 =  x_433 &  n_3307;
assign n_13756 =  x_2397 &  n_3308;
assign n_13757 = ~n_13755 & ~n_13756;
assign n_13758 =  x_2397 & ~n_13757;
assign n_13759 = ~x_2397 &  n_13757;
assign n_13760 = ~n_13758 & ~n_13759;
assign n_13761 =  x_432 &  n_3307;
assign n_13762 =  x_2396 &  n_3308;
assign n_13763 = ~n_13761 & ~n_13762;
assign n_13764 =  x_2396 & ~n_13763;
assign n_13765 = ~x_2396 &  n_13763;
assign n_13766 = ~n_13764 & ~n_13765;
assign n_13767 =  x_431 &  n_3307;
assign n_13768 =  x_2395 &  n_3308;
assign n_13769 = ~n_13767 & ~n_13768;
assign n_13770 =  x_2395 & ~n_13769;
assign n_13771 = ~x_2395 &  n_13769;
assign n_13772 = ~n_13770 & ~n_13771;
assign n_13773 =  x_430 &  n_3307;
assign n_13774 =  x_2394 &  n_3308;
assign n_13775 = ~n_13773 & ~n_13774;
assign n_13776 =  x_2394 & ~n_13775;
assign n_13777 = ~x_2394 &  n_13775;
assign n_13778 = ~n_13776 & ~n_13777;
assign n_13779 =  x_429 &  n_3307;
assign n_13780 =  x_2393 &  n_3308;
assign n_13781 = ~n_13779 & ~n_13780;
assign n_13782 =  x_2393 & ~n_13781;
assign n_13783 = ~x_2393 &  n_13781;
assign n_13784 = ~n_13782 & ~n_13783;
assign n_13785 =  x_428 &  n_3307;
assign n_13786 =  x_2392 &  n_3308;
assign n_13787 = ~n_13785 & ~n_13786;
assign n_13788 =  x_2392 & ~n_13787;
assign n_13789 = ~x_2392 &  n_13787;
assign n_13790 = ~n_13788 & ~n_13789;
assign n_13791 =  x_427 &  n_3307;
assign n_13792 =  x_2391 &  n_3308;
assign n_13793 = ~n_13791 & ~n_13792;
assign n_13794 =  x_2391 & ~n_13793;
assign n_13795 = ~x_2391 &  n_13793;
assign n_13796 = ~n_13794 & ~n_13795;
assign n_13797 =  x_426 &  n_3307;
assign n_13798 =  x_2390 &  n_3308;
assign n_13799 = ~n_13797 & ~n_13798;
assign n_13800 =  x_2390 & ~n_13799;
assign n_13801 = ~x_2390 &  n_13799;
assign n_13802 = ~n_13800 & ~n_13801;
assign n_13803 =  x_425 &  n_3307;
assign n_13804 =  x_2389 &  n_3308;
assign n_13805 = ~n_13803 & ~n_13804;
assign n_13806 =  x_2389 & ~n_13805;
assign n_13807 = ~x_2389 &  n_13805;
assign n_13808 = ~n_13806 & ~n_13807;
assign n_13809 =  x_424 &  n_3307;
assign n_13810 =  x_2388 &  n_3308;
assign n_13811 = ~n_13809 & ~n_13810;
assign n_13812 =  x_2388 & ~n_13811;
assign n_13813 = ~x_2388 &  n_13811;
assign n_13814 = ~n_13812 & ~n_13813;
assign n_13815 =  x_423 &  n_3307;
assign n_13816 =  x_2387 &  n_3308;
assign n_13817 = ~n_13815 & ~n_13816;
assign n_13818 =  x_2387 & ~n_13817;
assign n_13819 = ~x_2387 &  n_13817;
assign n_13820 = ~n_13818 & ~n_13819;
assign n_13821 =  x_422 &  n_3307;
assign n_13822 =  x_2386 &  n_3308;
assign n_13823 = ~n_13821 & ~n_13822;
assign n_13824 =  x_2386 & ~n_13823;
assign n_13825 = ~x_2386 &  n_13823;
assign n_13826 = ~n_13824 & ~n_13825;
assign n_13827 =  x_421 &  n_3307;
assign n_13828 =  x_2385 &  n_3308;
assign n_13829 = ~n_13827 & ~n_13828;
assign n_13830 =  x_2385 & ~n_13829;
assign n_13831 = ~x_2385 &  n_13829;
assign n_13832 = ~n_13830 & ~n_13831;
assign n_13833 =  x_420 &  n_3307;
assign n_13834 =  x_2384 &  n_3308;
assign n_13835 = ~n_13833 & ~n_13834;
assign n_13836 =  x_2384 & ~n_13835;
assign n_13837 = ~x_2384 &  n_13835;
assign n_13838 = ~n_13836 & ~n_13837;
assign n_13839 =  x_419 &  n_3307;
assign n_13840 =  x_2383 &  n_3308;
assign n_13841 = ~n_13839 & ~n_13840;
assign n_13842 =  x_2383 & ~n_13841;
assign n_13843 = ~x_2383 &  n_13841;
assign n_13844 = ~n_13842 & ~n_13843;
assign n_13845 =  x_418 &  n_3307;
assign n_13846 =  x_2382 &  n_3308;
assign n_13847 = ~n_13845 & ~n_13846;
assign n_13848 =  x_2382 & ~n_13847;
assign n_13849 = ~x_2382 &  n_13847;
assign n_13850 = ~n_13848 & ~n_13849;
assign n_13851 =  x_417 &  n_3307;
assign n_13852 =  x_2381 &  n_3308;
assign n_13853 = ~n_13851 & ~n_13852;
assign n_13854 =  x_2381 & ~n_13853;
assign n_13855 = ~x_2381 &  n_13853;
assign n_13856 = ~n_13854 & ~n_13855;
assign n_13857 =  x_416 &  n_3307;
assign n_13858 =  x_2380 &  n_3308;
assign n_13859 = ~n_13857 & ~n_13858;
assign n_13860 =  x_2380 & ~n_13859;
assign n_13861 = ~x_2380 &  n_13859;
assign n_13862 = ~n_13860 & ~n_13861;
assign n_13863 =  x_415 &  n_3307;
assign n_13864 =  x_2379 &  n_3308;
assign n_13865 = ~n_13863 & ~n_13864;
assign n_13866 =  x_2379 & ~n_13865;
assign n_13867 = ~x_2379 &  n_13865;
assign n_13868 = ~n_13866 & ~n_13867;
assign n_13869 =  x_414 &  n_3307;
assign n_13870 =  x_2378 &  n_3308;
assign n_13871 = ~n_13869 & ~n_13870;
assign n_13872 =  x_2378 & ~n_13871;
assign n_13873 = ~x_2378 &  n_13871;
assign n_13874 = ~n_13872 & ~n_13873;
assign n_13875 =  x_413 &  n_3307;
assign n_13876 =  x_2377 &  n_3308;
assign n_13877 = ~n_13875 & ~n_13876;
assign n_13878 =  x_2377 & ~n_13877;
assign n_13879 = ~x_2377 &  n_13877;
assign n_13880 = ~n_13878 & ~n_13879;
assign n_13881 =  x_412 &  n_3307;
assign n_13882 =  x_2376 &  n_3308;
assign n_13883 = ~n_13881 & ~n_13882;
assign n_13884 =  x_2376 & ~n_13883;
assign n_13885 = ~x_2376 &  n_13883;
assign n_13886 = ~n_13884 & ~n_13885;
assign n_13887 =  x_411 &  n_3307;
assign n_13888 =  x_2375 &  n_3308;
assign n_13889 = ~n_13887 & ~n_13888;
assign n_13890 =  x_2375 & ~n_13889;
assign n_13891 = ~x_2375 &  n_13889;
assign n_13892 = ~n_13890 & ~n_13891;
assign n_13893 =  x_410 &  n_3307;
assign n_13894 =  x_2374 &  n_3308;
assign n_13895 = ~n_13893 & ~n_13894;
assign n_13896 =  x_2374 & ~n_13895;
assign n_13897 = ~x_2374 &  n_13895;
assign n_13898 = ~n_13896 & ~n_13897;
assign n_13899 =  x_409 &  n_3307;
assign n_13900 =  x_2373 &  n_3308;
assign n_13901 = ~n_13899 & ~n_13900;
assign n_13902 =  x_2373 & ~n_13901;
assign n_13903 = ~x_2373 &  n_13901;
assign n_13904 = ~n_13902 & ~n_13903;
assign n_13905 =  x_408 &  n_3307;
assign n_13906 =  x_2372 &  n_3308;
assign n_13907 = ~n_13905 & ~n_13906;
assign n_13908 =  x_2372 & ~n_13907;
assign n_13909 = ~x_2372 &  n_13907;
assign n_13910 = ~n_13908 & ~n_13909;
assign n_13911 =  x_407 &  n_3307;
assign n_13912 =  x_2371 &  n_3308;
assign n_13913 = ~n_13911 & ~n_13912;
assign n_13914 =  x_2371 & ~n_13913;
assign n_13915 = ~x_2371 &  n_13913;
assign n_13916 = ~n_13914 & ~n_13915;
assign n_13917 =  x_406 &  n_3307;
assign n_13918 =  x_2370 &  n_3308;
assign n_13919 = ~n_13917 & ~n_13918;
assign n_13920 =  x_2370 & ~n_13919;
assign n_13921 = ~x_2370 &  n_13919;
assign n_13922 = ~n_13920 & ~n_13921;
assign n_13923 =  x_405 &  n_3307;
assign n_13924 =  x_2369 &  n_3308;
assign n_13925 = ~n_13923 & ~n_13924;
assign n_13926 =  x_2369 & ~n_13925;
assign n_13927 = ~x_2369 &  n_13925;
assign n_13928 = ~n_13926 & ~n_13927;
assign n_13929 =  x_404 &  n_3307;
assign n_13930 =  x_2368 &  n_3308;
assign n_13931 = ~n_13929 & ~n_13930;
assign n_13932 =  x_2368 & ~n_13931;
assign n_13933 = ~x_2368 &  n_13931;
assign n_13934 = ~n_13932 & ~n_13933;
assign n_13935 =  x_403 &  n_3307;
assign n_13936 =  x_2367 &  n_3308;
assign n_13937 = ~n_13935 & ~n_13936;
assign n_13938 =  x_2367 & ~n_13937;
assign n_13939 = ~x_2367 &  n_13937;
assign n_13940 = ~n_13938 & ~n_13939;
assign n_13941 = ~x_402 &  n_3307;
assign n_13942 =  x_2366 &  n_3308;
assign n_13943 = ~n_13941 & ~n_13942;
assign n_13944 =  x_2366 & ~n_13943;
assign n_13945 = ~x_2366 &  n_13943;
assign n_13946 = ~n_13944 & ~n_13945;
assign n_13947 =  x_2365 & ~n_1761;
assign n_13948 =  i_216 &  n_1751;
assign n_13949 =  n_1761 &  n_13948;
assign n_13950 = ~n_13947 & ~n_13949;
assign n_13951 =  x_2365 & ~n_13950;
assign n_13952 = ~x_2365 &  n_13950;
assign n_13953 = ~n_13951 & ~n_13952;
assign n_13954 =  x_2364 & ~n_1770;
assign n_13955 =  n_1770 &  n_13948;
assign n_13956 = ~n_13954 & ~n_13955;
assign n_13957 =  x_2364 & ~n_13956;
assign n_13958 = ~x_2364 &  n_13956;
assign n_13959 = ~n_13957 & ~n_13958;
assign n_13960 =  x_2363 & ~n_1778;
assign n_13961 =  n_1778 &  n_13948;
assign n_13962 = ~n_13960 & ~n_13961;
assign n_13963 =  x_2363 & ~n_13962;
assign n_13964 = ~x_2363 &  n_13962;
assign n_13965 = ~n_13963 & ~n_13964;
assign n_13966 =  x_2362 & ~n_1785;
assign n_13967 =  n_1785 &  n_13948;
assign n_13968 = ~n_13966 & ~n_13967;
assign n_13969 =  x_2362 & ~n_13968;
assign n_13970 = ~x_2362 &  n_13968;
assign n_13971 = ~n_13969 & ~n_13970;
assign n_13972 =  x_2361 & ~n_1792;
assign n_13973 =  n_1792 &  n_13948;
assign n_13974 = ~n_13972 & ~n_13973;
assign n_13975 =  x_2361 & ~n_13974;
assign n_13976 = ~x_2361 &  n_13974;
assign n_13977 = ~n_13975 & ~n_13976;
assign n_13978 =  x_2360 & ~n_1799;
assign n_13979 =  n_1799 &  n_13948;
assign n_13980 = ~n_13978 & ~n_13979;
assign n_13981 =  x_2360 & ~n_13980;
assign n_13982 = ~x_2360 &  n_13980;
assign n_13983 = ~n_13981 & ~n_13982;
assign n_13984 =  x_2359 & ~n_1806;
assign n_13985 =  n_1806 &  n_13948;
assign n_13986 = ~n_13984 & ~n_13985;
assign n_13987 =  x_2359 & ~n_13986;
assign n_13988 = ~x_2359 &  n_13986;
assign n_13989 = ~n_13987 & ~n_13988;
assign n_13990 =  n_1750 & ~n_13948;
assign n_13991 = ~x_2358 & ~n_1750;
assign n_13992 = ~n_13990 & ~n_13991;
assign n_13993 =  x_2358 &  n_13992;
assign n_13994 = ~x_2358 & ~n_13992;
assign n_13995 = ~n_13993 & ~n_13994;
assign n_13996 =  x_2357 & ~n_1761;
assign n_13997 =  i_215 &  n_1751;
assign n_13998 =  n_1761 &  n_13997;
assign n_13999 = ~n_13996 & ~n_13998;
assign n_14000 =  x_2357 & ~n_13999;
assign n_14001 = ~x_2357 &  n_13999;
assign n_14002 = ~n_14000 & ~n_14001;
assign n_14003 =  x_2356 & ~n_1770;
assign n_14004 =  n_1770 &  n_13997;
assign n_14005 = ~n_14003 & ~n_14004;
assign n_14006 =  x_2356 & ~n_14005;
assign n_14007 = ~x_2356 &  n_14005;
assign n_14008 = ~n_14006 & ~n_14007;
assign n_14009 =  x_2355 & ~n_1778;
assign n_14010 =  n_1778 &  n_13997;
assign n_14011 = ~n_14009 & ~n_14010;
assign n_14012 =  x_2355 & ~n_14011;
assign n_14013 = ~x_2355 &  n_14011;
assign n_14014 = ~n_14012 & ~n_14013;
assign n_14015 =  x_2354 & ~n_1785;
assign n_14016 =  n_1785 &  n_13997;
assign n_14017 = ~n_14015 & ~n_14016;
assign n_14018 =  x_2354 & ~n_14017;
assign n_14019 = ~x_2354 &  n_14017;
assign n_14020 = ~n_14018 & ~n_14019;
assign n_14021 =  x_2353 & ~n_1792;
assign n_14022 =  n_1792 &  n_13997;
assign n_14023 = ~n_14021 & ~n_14022;
assign n_14024 =  x_2353 & ~n_14023;
assign n_14025 = ~x_2353 &  n_14023;
assign n_14026 = ~n_14024 & ~n_14025;
assign n_14027 =  x_2352 & ~n_1799;
assign n_14028 =  n_1799 &  n_13997;
assign n_14029 = ~n_14027 & ~n_14028;
assign n_14030 =  x_2352 & ~n_14029;
assign n_14031 = ~x_2352 &  n_14029;
assign n_14032 = ~n_14030 & ~n_14031;
assign n_14033 =  x_2351 & ~n_1806;
assign n_14034 =  n_1806 &  n_13997;
assign n_14035 = ~n_14033 & ~n_14034;
assign n_14036 =  x_2351 & ~n_14035;
assign n_14037 = ~x_2351 &  n_14035;
assign n_14038 = ~n_14036 & ~n_14037;
assign n_14039 =  n_1750 & ~n_13997;
assign n_14040 = ~x_2350 & ~n_1750;
assign n_14041 = ~n_14039 & ~n_14040;
assign n_14042 =  x_2350 &  n_14041;
assign n_14043 = ~x_2350 & ~n_14041;
assign n_14044 = ~n_14042 & ~n_14043;
assign n_14045 =  x_2349 & ~n_1761;
assign n_14046 =  i_214 &  n_1751;
assign n_14047 =  n_1761 &  n_14046;
assign n_14048 = ~n_14045 & ~n_14047;
assign n_14049 =  x_2349 & ~n_14048;
assign n_14050 = ~x_2349 &  n_14048;
assign n_14051 = ~n_14049 & ~n_14050;
assign n_14052 =  x_2348 & ~n_1770;
assign n_14053 =  n_1770 &  n_14046;
assign n_14054 = ~n_14052 & ~n_14053;
assign n_14055 =  x_2348 & ~n_14054;
assign n_14056 = ~x_2348 &  n_14054;
assign n_14057 = ~n_14055 & ~n_14056;
assign n_14058 =  x_2347 & ~n_1778;
assign n_14059 =  n_1778 &  n_14046;
assign n_14060 = ~n_14058 & ~n_14059;
assign n_14061 =  x_2347 & ~n_14060;
assign n_14062 = ~x_2347 &  n_14060;
assign n_14063 = ~n_14061 & ~n_14062;
assign n_14064 =  x_2346 & ~n_1785;
assign n_14065 =  n_1785 &  n_14046;
assign n_14066 = ~n_14064 & ~n_14065;
assign n_14067 =  x_2346 & ~n_14066;
assign n_14068 = ~x_2346 &  n_14066;
assign n_14069 = ~n_14067 & ~n_14068;
assign n_14070 =  x_2345 & ~n_1792;
assign n_14071 =  n_1792 &  n_14046;
assign n_14072 = ~n_14070 & ~n_14071;
assign n_14073 =  x_2345 & ~n_14072;
assign n_14074 = ~x_2345 &  n_14072;
assign n_14075 = ~n_14073 & ~n_14074;
assign n_14076 =  x_2344 & ~n_1799;
assign n_14077 =  n_1799 &  n_14046;
assign n_14078 = ~n_14076 & ~n_14077;
assign n_14079 =  x_2344 & ~n_14078;
assign n_14080 = ~x_2344 &  n_14078;
assign n_14081 = ~n_14079 & ~n_14080;
assign n_14082 =  x_2343 & ~n_1806;
assign n_14083 =  n_1806 &  n_14046;
assign n_14084 = ~n_14082 & ~n_14083;
assign n_14085 =  x_2343 & ~n_14084;
assign n_14086 = ~x_2343 &  n_14084;
assign n_14087 = ~n_14085 & ~n_14086;
assign n_14088 =  n_1750 & ~n_14046;
assign n_14089 = ~x_2342 & ~n_1750;
assign n_14090 = ~n_14088 & ~n_14089;
assign n_14091 =  x_2342 &  n_14090;
assign n_14092 = ~x_2342 & ~n_14090;
assign n_14093 = ~n_14091 & ~n_14092;
assign n_14094 =  x_2341 & ~n_1761;
assign n_14095 =  i_213 &  n_1751;
assign n_14096 =  n_1761 &  n_14095;
assign n_14097 = ~n_14094 & ~n_14096;
assign n_14098 =  x_2341 & ~n_14097;
assign n_14099 = ~x_2341 &  n_14097;
assign n_14100 = ~n_14098 & ~n_14099;
assign n_14101 =  x_2340 & ~n_1770;
assign n_14102 =  n_1770 &  n_14095;
assign n_14103 = ~n_14101 & ~n_14102;
assign n_14104 =  x_2340 & ~n_14103;
assign n_14105 = ~x_2340 &  n_14103;
assign n_14106 = ~n_14104 & ~n_14105;
assign n_14107 =  x_2339 & ~n_1778;
assign n_14108 =  n_1778 &  n_14095;
assign n_14109 = ~n_14107 & ~n_14108;
assign n_14110 =  x_2339 & ~n_14109;
assign n_14111 = ~x_2339 &  n_14109;
assign n_14112 = ~n_14110 & ~n_14111;
assign n_14113 =  x_2338 & ~n_1785;
assign n_14114 =  n_1785 &  n_14095;
assign n_14115 = ~n_14113 & ~n_14114;
assign n_14116 =  x_2338 & ~n_14115;
assign n_14117 = ~x_2338 &  n_14115;
assign n_14118 = ~n_14116 & ~n_14117;
assign n_14119 =  x_2337 & ~n_1792;
assign n_14120 =  n_1792 &  n_14095;
assign n_14121 = ~n_14119 & ~n_14120;
assign n_14122 =  x_2337 & ~n_14121;
assign n_14123 = ~x_2337 &  n_14121;
assign n_14124 = ~n_14122 & ~n_14123;
assign n_14125 =  x_2336 & ~n_1799;
assign n_14126 =  n_1799 &  n_14095;
assign n_14127 = ~n_14125 & ~n_14126;
assign n_14128 =  x_2336 & ~n_14127;
assign n_14129 = ~x_2336 &  n_14127;
assign n_14130 = ~n_14128 & ~n_14129;
assign n_14131 =  x_2335 & ~n_1806;
assign n_14132 =  n_1806 &  n_14095;
assign n_14133 = ~n_14131 & ~n_14132;
assign n_14134 =  x_2335 & ~n_14133;
assign n_14135 = ~x_2335 &  n_14133;
assign n_14136 = ~n_14134 & ~n_14135;
assign n_14137 =  n_1750 & ~n_14095;
assign n_14138 = ~x_2334 & ~n_1750;
assign n_14139 = ~n_14137 & ~n_14138;
assign n_14140 =  x_2334 &  n_14139;
assign n_14141 = ~x_2334 & ~n_14139;
assign n_14142 = ~n_14140 & ~n_14141;
assign n_14143 =  x_2333 & ~n_1761;
assign n_14144 =  i_212 &  n_1751;
assign n_14145 =  n_1761 &  n_14144;
assign n_14146 = ~n_14143 & ~n_14145;
assign n_14147 =  x_2333 & ~n_14146;
assign n_14148 = ~x_2333 &  n_14146;
assign n_14149 = ~n_14147 & ~n_14148;
assign n_14150 =  x_2332 & ~n_1770;
assign n_14151 =  n_1770 &  n_14144;
assign n_14152 = ~n_14150 & ~n_14151;
assign n_14153 =  x_2332 & ~n_14152;
assign n_14154 = ~x_2332 &  n_14152;
assign n_14155 = ~n_14153 & ~n_14154;
assign n_14156 =  x_2331 & ~n_1778;
assign n_14157 =  n_1778 &  n_14144;
assign n_14158 = ~n_14156 & ~n_14157;
assign n_14159 =  x_2331 & ~n_14158;
assign n_14160 = ~x_2331 &  n_14158;
assign n_14161 = ~n_14159 & ~n_14160;
assign n_14162 =  x_2330 & ~n_1785;
assign n_14163 =  n_1785 &  n_14144;
assign n_14164 = ~n_14162 & ~n_14163;
assign n_14165 =  x_2330 & ~n_14164;
assign n_14166 = ~x_2330 &  n_14164;
assign n_14167 = ~n_14165 & ~n_14166;
assign n_14168 =  x_2329 & ~n_1792;
assign n_14169 =  n_1792 &  n_14144;
assign n_14170 = ~n_14168 & ~n_14169;
assign n_14171 =  x_2329 & ~n_14170;
assign n_14172 = ~x_2329 &  n_14170;
assign n_14173 = ~n_14171 & ~n_14172;
assign n_14174 =  x_2328 & ~n_1799;
assign n_14175 =  n_1799 &  n_14144;
assign n_14176 = ~n_14174 & ~n_14175;
assign n_14177 =  x_2328 & ~n_14176;
assign n_14178 = ~x_2328 &  n_14176;
assign n_14179 = ~n_14177 & ~n_14178;
assign n_14180 =  x_2327 & ~n_1806;
assign n_14181 =  n_1806 &  n_14144;
assign n_14182 = ~n_14180 & ~n_14181;
assign n_14183 =  x_2327 & ~n_14182;
assign n_14184 = ~x_2327 &  n_14182;
assign n_14185 = ~n_14183 & ~n_14184;
assign n_14186 =  n_1750 & ~n_14144;
assign n_14187 = ~x_2326 & ~n_1750;
assign n_14188 = ~n_14186 & ~n_14187;
assign n_14189 =  x_2326 &  n_14188;
assign n_14190 = ~x_2326 & ~n_14188;
assign n_14191 = ~n_14189 & ~n_14190;
assign n_14192 =  x_2325 & ~n_1761;
assign n_14193 =  i_211 &  n_1751;
assign n_14194 =  n_1761 &  n_14193;
assign n_14195 = ~n_14192 & ~n_14194;
assign n_14196 =  x_2325 & ~n_14195;
assign n_14197 = ~x_2325 &  n_14195;
assign n_14198 = ~n_14196 & ~n_14197;
assign n_14199 =  x_2324 & ~n_1770;
assign n_14200 =  n_1770 &  n_14193;
assign n_14201 = ~n_14199 & ~n_14200;
assign n_14202 =  x_2324 & ~n_14201;
assign n_14203 = ~x_2324 &  n_14201;
assign n_14204 = ~n_14202 & ~n_14203;
assign n_14205 =  x_2323 & ~n_1778;
assign n_14206 =  n_1778 &  n_14193;
assign n_14207 = ~n_14205 & ~n_14206;
assign n_14208 =  x_2323 & ~n_14207;
assign n_14209 = ~x_2323 &  n_14207;
assign n_14210 = ~n_14208 & ~n_14209;
assign n_14211 =  x_2322 & ~n_1785;
assign n_14212 =  n_1785 &  n_14193;
assign n_14213 = ~n_14211 & ~n_14212;
assign n_14214 =  x_2322 & ~n_14213;
assign n_14215 = ~x_2322 &  n_14213;
assign n_14216 = ~n_14214 & ~n_14215;
assign n_14217 =  x_2321 & ~n_1792;
assign n_14218 =  n_1792 &  n_14193;
assign n_14219 = ~n_14217 & ~n_14218;
assign n_14220 =  x_2321 & ~n_14219;
assign n_14221 = ~x_2321 &  n_14219;
assign n_14222 = ~n_14220 & ~n_14221;
assign n_14223 =  x_2320 & ~n_1799;
assign n_14224 =  n_1799 &  n_14193;
assign n_14225 = ~n_14223 & ~n_14224;
assign n_14226 =  x_2320 & ~n_14225;
assign n_14227 = ~x_2320 &  n_14225;
assign n_14228 = ~n_14226 & ~n_14227;
assign n_14229 =  x_2319 & ~n_1806;
assign n_14230 =  n_1806 &  n_14193;
assign n_14231 = ~n_14229 & ~n_14230;
assign n_14232 =  x_2319 & ~n_14231;
assign n_14233 = ~x_2319 &  n_14231;
assign n_14234 = ~n_14232 & ~n_14233;
assign n_14235 =  n_1750 & ~n_14193;
assign n_14236 = ~x_2318 & ~n_1750;
assign n_14237 = ~n_14235 & ~n_14236;
assign n_14238 =  x_2318 &  n_14237;
assign n_14239 = ~x_2318 & ~n_14237;
assign n_14240 = ~n_14238 & ~n_14239;
assign n_14241 =  x_2317 & ~n_1761;
assign n_14242 =  i_210 &  n_1751;
assign n_14243 =  n_1761 &  n_14242;
assign n_14244 = ~n_14241 & ~n_14243;
assign n_14245 =  x_2317 & ~n_14244;
assign n_14246 = ~x_2317 &  n_14244;
assign n_14247 = ~n_14245 & ~n_14246;
assign n_14248 =  x_2316 & ~n_1770;
assign n_14249 =  n_1770 &  n_14242;
assign n_14250 = ~n_14248 & ~n_14249;
assign n_14251 =  x_2316 & ~n_14250;
assign n_14252 = ~x_2316 &  n_14250;
assign n_14253 = ~n_14251 & ~n_14252;
assign n_14254 =  x_2315 & ~n_1778;
assign n_14255 =  n_1778 &  n_14242;
assign n_14256 = ~n_14254 & ~n_14255;
assign n_14257 =  x_2315 & ~n_14256;
assign n_14258 = ~x_2315 &  n_14256;
assign n_14259 = ~n_14257 & ~n_14258;
assign n_14260 =  x_2314 & ~n_1785;
assign n_14261 =  n_1785 &  n_14242;
assign n_14262 = ~n_14260 & ~n_14261;
assign n_14263 =  x_2314 & ~n_14262;
assign n_14264 = ~x_2314 &  n_14262;
assign n_14265 = ~n_14263 & ~n_14264;
assign n_14266 =  x_2313 & ~n_1792;
assign n_14267 =  n_1792 &  n_14242;
assign n_14268 = ~n_14266 & ~n_14267;
assign n_14269 =  x_2313 & ~n_14268;
assign n_14270 = ~x_2313 &  n_14268;
assign n_14271 = ~n_14269 & ~n_14270;
assign n_14272 =  x_2312 & ~n_1799;
assign n_14273 =  n_1799 &  n_14242;
assign n_14274 = ~n_14272 & ~n_14273;
assign n_14275 =  x_2312 & ~n_14274;
assign n_14276 = ~x_2312 &  n_14274;
assign n_14277 = ~n_14275 & ~n_14276;
assign n_14278 =  x_2311 & ~n_1806;
assign n_14279 =  n_1806 &  n_14242;
assign n_14280 = ~n_14278 & ~n_14279;
assign n_14281 =  x_2311 & ~n_14280;
assign n_14282 = ~x_2311 &  n_14280;
assign n_14283 = ~n_14281 & ~n_14282;
assign n_14284 =  n_1750 & ~n_14242;
assign n_14285 = ~x_2310 & ~n_1750;
assign n_14286 = ~n_14284 & ~n_14285;
assign n_14287 =  x_2310 &  n_14286;
assign n_14288 = ~x_2310 & ~n_14286;
assign n_14289 = ~n_14287 & ~n_14288;
assign n_14290 =  x_2309 & ~n_1761;
assign n_14291 =  i_209 &  n_1751;
assign n_14292 =  n_1761 &  n_14291;
assign n_14293 = ~n_14290 & ~n_14292;
assign n_14294 =  x_2309 & ~n_14293;
assign n_14295 = ~x_2309 &  n_14293;
assign n_14296 = ~n_14294 & ~n_14295;
assign n_14297 =  x_2308 & ~n_1770;
assign n_14298 =  n_1770 &  n_14291;
assign n_14299 = ~n_14297 & ~n_14298;
assign n_14300 =  x_2308 & ~n_14299;
assign n_14301 = ~x_2308 &  n_14299;
assign n_14302 = ~n_14300 & ~n_14301;
assign n_14303 =  x_2307 & ~n_1778;
assign n_14304 =  n_1778 &  n_14291;
assign n_14305 = ~n_14303 & ~n_14304;
assign n_14306 =  x_2307 & ~n_14305;
assign n_14307 = ~x_2307 &  n_14305;
assign n_14308 = ~n_14306 & ~n_14307;
assign n_14309 =  x_2306 & ~n_1785;
assign n_14310 =  n_1785 &  n_14291;
assign n_14311 = ~n_14309 & ~n_14310;
assign n_14312 =  x_2306 & ~n_14311;
assign n_14313 = ~x_2306 &  n_14311;
assign n_14314 = ~n_14312 & ~n_14313;
assign n_14315 =  x_2305 & ~n_1792;
assign n_14316 =  n_1792 &  n_14291;
assign n_14317 = ~n_14315 & ~n_14316;
assign n_14318 =  x_2305 & ~n_14317;
assign n_14319 = ~x_2305 &  n_14317;
assign n_14320 = ~n_14318 & ~n_14319;
assign n_14321 =  x_2304 & ~n_1799;
assign n_14322 =  n_1799 &  n_14291;
assign n_14323 = ~n_14321 & ~n_14322;
assign n_14324 =  x_2304 & ~n_14323;
assign n_14325 = ~x_2304 &  n_14323;
assign n_14326 = ~n_14324 & ~n_14325;
assign n_14327 =  x_2303 & ~n_1806;
assign n_14328 =  n_1806 &  n_14291;
assign n_14329 = ~n_14327 & ~n_14328;
assign n_14330 =  x_2303 & ~n_14329;
assign n_14331 = ~x_2303 &  n_14329;
assign n_14332 = ~n_14330 & ~n_14331;
assign n_14333 =  n_1750 & ~n_14291;
assign n_14334 = ~x_2302 & ~n_1750;
assign n_14335 = ~n_14333 & ~n_14334;
assign n_14336 =  x_2302 &  n_14335;
assign n_14337 = ~x_2302 & ~n_14335;
assign n_14338 = ~n_14336 & ~n_14337;
assign n_14339 =  x_2301 & ~n_1761;
assign n_14340 =  i_208 &  n_1751;
assign n_14341 =  n_1761 &  n_14340;
assign n_14342 = ~n_14339 & ~n_14341;
assign n_14343 =  x_2301 & ~n_14342;
assign n_14344 = ~x_2301 &  n_14342;
assign n_14345 = ~n_14343 & ~n_14344;
assign n_14346 =  x_2300 & ~n_1770;
assign n_14347 =  n_1770 &  n_14340;
assign n_14348 = ~n_14346 & ~n_14347;
assign n_14349 =  x_2300 & ~n_14348;
assign n_14350 = ~x_2300 &  n_14348;
assign n_14351 = ~n_14349 & ~n_14350;
assign n_14352 =  x_2299 & ~n_1778;
assign n_14353 =  n_1778 &  n_14340;
assign n_14354 = ~n_14352 & ~n_14353;
assign n_14355 =  x_2299 & ~n_14354;
assign n_14356 = ~x_2299 &  n_14354;
assign n_14357 = ~n_14355 & ~n_14356;
assign n_14358 =  x_2298 & ~n_1785;
assign n_14359 =  n_1785 &  n_14340;
assign n_14360 = ~n_14358 & ~n_14359;
assign n_14361 =  x_2298 & ~n_14360;
assign n_14362 = ~x_2298 &  n_14360;
assign n_14363 = ~n_14361 & ~n_14362;
assign n_14364 =  x_2297 & ~n_1792;
assign n_14365 =  n_1792 &  n_14340;
assign n_14366 = ~n_14364 & ~n_14365;
assign n_14367 =  x_2297 & ~n_14366;
assign n_14368 = ~x_2297 &  n_14366;
assign n_14369 = ~n_14367 & ~n_14368;
assign n_14370 =  x_2296 & ~n_1799;
assign n_14371 =  n_1799 &  n_14340;
assign n_14372 = ~n_14370 & ~n_14371;
assign n_14373 =  x_2296 & ~n_14372;
assign n_14374 = ~x_2296 &  n_14372;
assign n_14375 = ~n_14373 & ~n_14374;
assign n_14376 =  x_2295 & ~n_1806;
assign n_14377 =  n_1806 &  n_14340;
assign n_14378 = ~n_14376 & ~n_14377;
assign n_14379 =  x_2295 & ~n_14378;
assign n_14380 = ~x_2295 &  n_14378;
assign n_14381 = ~n_14379 & ~n_14380;
assign n_14382 =  n_1750 & ~n_14340;
assign n_14383 = ~x_2294 & ~n_1750;
assign n_14384 = ~n_14382 & ~n_14383;
assign n_14385 =  x_2294 &  n_14384;
assign n_14386 = ~x_2294 & ~n_14384;
assign n_14387 = ~n_14385 & ~n_14386;
assign n_14388 =  x_2293 & ~n_1761;
assign n_14389 =  i_207 &  n_1751;
assign n_14390 =  n_1761 &  n_14389;
assign n_14391 = ~n_14388 & ~n_14390;
assign n_14392 =  x_2293 & ~n_14391;
assign n_14393 = ~x_2293 &  n_14391;
assign n_14394 = ~n_14392 & ~n_14393;
assign n_14395 =  x_2292 & ~n_1770;
assign n_14396 =  n_1770 &  n_14389;
assign n_14397 = ~n_14395 & ~n_14396;
assign n_14398 =  x_2292 & ~n_14397;
assign n_14399 = ~x_2292 &  n_14397;
assign n_14400 = ~n_14398 & ~n_14399;
assign n_14401 =  x_2291 & ~n_1778;
assign n_14402 =  n_1778 &  n_14389;
assign n_14403 = ~n_14401 & ~n_14402;
assign n_14404 =  x_2291 & ~n_14403;
assign n_14405 = ~x_2291 &  n_14403;
assign n_14406 = ~n_14404 & ~n_14405;
assign n_14407 =  x_2290 & ~n_1785;
assign n_14408 =  n_1785 &  n_14389;
assign n_14409 = ~n_14407 & ~n_14408;
assign n_14410 =  x_2290 & ~n_14409;
assign n_14411 = ~x_2290 &  n_14409;
assign n_14412 = ~n_14410 & ~n_14411;
assign n_14413 =  x_2289 & ~n_1792;
assign n_14414 =  n_1792 &  n_14389;
assign n_14415 = ~n_14413 & ~n_14414;
assign n_14416 =  x_2289 & ~n_14415;
assign n_14417 = ~x_2289 &  n_14415;
assign n_14418 = ~n_14416 & ~n_14417;
assign n_14419 =  x_2288 & ~n_1799;
assign n_14420 =  n_1799 &  n_14389;
assign n_14421 = ~n_14419 & ~n_14420;
assign n_14422 =  x_2288 & ~n_14421;
assign n_14423 = ~x_2288 &  n_14421;
assign n_14424 = ~n_14422 & ~n_14423;
assign n_14425 =  x_2287 & ~n_1806;
assign n_14426 =  n_1806 &  n_14389;
assign n_14427 = ~n_14425 & ~n_14426;
assign n_14428 =  x_2287 & ~n_14427;
assign n_14429 = ~x_2287 &  n_14427;
assign n_14430 = ~n_14428 & ~n_14429;
assign n_14431 =  n_1750 & ~n_14389;
assign n_14432 = ~x_2286 & ~n_1750;
assign n_14433 = ~n_14431 & ~n_14432;
assign n_14434 =  x_2286 &  n_14433;
assign n_14435 = ~x_2286 & ~n_14433;
assign n_14436 = ~n_14434 & ~n_14435;
assign n_14437 =  x_2285 & ~n_1761;
assign n_14438 =  i_206 &  n_1751;
assign n_14439 =  n_1761 &  n_14438;
assign n_14440 = ~n_14437 & ~n_14439;
assign n_14441 =  x_2285 & ~n_14440;
assign n_14442 = ~x_2285 &  n_14440;
assign n_14443 = ~n_14441 & ~n_14442;
assign n_14444 =  x_2284 & ~n_1770;
assign n_14445 =  n_1770 &  n_14438;
assign n_14446 = ~n_14444 & ~n_14445;
assign n_14447 =  x_2284 & ~n_14446;
assign n_14448 = ~x_2284 &  n_14446;
assign n_14449 = ~n_14447 & ~n_14448;
assign n_14450 =  x_2283 & ~n_1778;
assign n_14451 =  n_1778 &  n_14438;
assign n_14452 = ~n_14450 & ~n_14451;
assign n_14453 =  x_2283 & ~n_14452;
assign n_14454 = ~x_2283 &  n_14452;
assign n_14455 = ~n_14453 & ~n_14454;
assign n_14456 =  x_2282 & ~n_1785;
assign n_14457 =  n_1785 &  n_14438;
assign n_14458 = ~n_14456 & ~n_14457;
assign n_14459 =  x_2282 & ~n_14458;
assign n_14460 = ~x_2282 &  n_14458;
assign n_14461 = ~n_14459 & ~n_14460;
assign n_14462 =  x_2281 & ~n_1792;
assign n_14463 =  n_1792 &  n_14438;
assign n_14464 = ~n_14462 & ~n_14463;
assign n_14465 =  x_2281 & ~n_14464;
assign n_14466 = ~x_2281 &  n_14464;
assign n_14467 = ~n_14465 & ~n_14466;
assign n_14468 =  x_2280 & ~n_1799;
assign n_14469 =  n_1799 &  n_14438;
assign n_14470 = ~n_14468 & ~n_14469;
assign n_14471 =  x_2280 & ~n_14470;
assign n_14472 = ~x_2280 &  n_14470;
assign n_14473 = ~n_14471 & ~n_14472;
assign n_14474 =  x_2279 & ~n_1806;
assign n_14475 =  n_1806 &  n_14438;
assign n_14476 = ~n_14474 & ~n_14475;
assign n_14477 =  x_2279 & ~n_14476;
assign n_14478 = ~x_2279 &  n_14476;
assign n_14479 = ~n_14477 & ~n_14478;
assign n_14480 =  n_1750 & ~n_14438;
assign n_14481 = ~x_2278 & ~n_1750;
assign n_14482 = ~n_14480 & ~n_14481;
assign n_14483 =  x_2278 &  n_14482;
assign n_14484 = ~x_2278 & ~n_14482;
assign n_14485 = ~n_14483 & ~n_14484;
assign n_14486 =  x_2277 & ~n_1761;
assign n_14487 =  i_205 &  n_1751;
assign n_14488 =  n_1761 &  n_14487;
assign n_14489 = ~n_14486 & ~n_14488;
assign n_14490 =  x_2277 & ~n_14489;
assign n_14491 = ~x_2277 &  n_14489;
assign n_14492 = ~n_14490 & ~n_14491;
assign n_14493 =  x_2276 & ~n_1770;
assign n_14494 =  n_1770 &  n_14487;
assign n_14495 = ~n_14493 & ~n_14494;
assign n_14496 =  x_2276 & ~n_14495;
assign n_14497 = ~x_2276 &  n_14495;
assign n_14498 = ~n_14496 & ~n_14497;
assign n_14499 =  x_2275 & ~n_1778;
assign n_14500 =  n_1778 &  n_14487;
assign n_14501 = ~n_14499 & ~n_14500;
assign n_14502 =  x_2275 & ~n_14501;
assign n_14503 = ~x_2275 &  n_14501;
assign n_14504 = ~n_14502 & ~n_14503;
assign n_14505 =  x_2274 & ~n_1785;
assign n_14506 =  n_1785 &  n_14487;
assign n_14507 = ~n_14505 & ~n_14506;
assign n_14508 =  x_2274 & ~n_14507;
assign n_14509 = ~x_2274 &  n_14507;
assign n_14510 = ~n_14508 & ~n_14509;
assign n_14511 =  x_2273 & ~n_1792;
assign n_14512 =  n_1792 &  n_14487;
assign n_14513 = ~n_14511 & ~n_14512;
assign n_14514 =  x_2273 & ~n_14513;
assign n_14515 = ~x_2273 &  n_14513;
assign n_14516 = ~n_14514 & ~n_14515;
assign n_14517 =  x_2272 & ~n_1799;
assign n_14518 =  n_1799 &  n_14487;
assign n_14519 = ~n_14517 & ~n_14518;
assign n_14520 =  x_2272 & ~n_14519;
assign n_14521 = ~x_2272 &  n_14519;
assign n_14522 = ~n_14520 & ~n_14521;
assign n_14523 =  x_2271 & ~n_1806;
assign n_14524 =  n_1806 &  n_14487;
assign n_14525 = ~n_14523 & ~n_14524;
assign n_14526 =  x_2271 & ~n_14525;
assign n_14527 = ~x_2271 &  n_14525;
assign n_14528 = ~n_14526 & ~n_14527;
assign n_14529 =  n_1750 & ~n_14487;
assign n_14530 = ~x_2270 & ~n_1750;
assign n_14531 = ~n_14529 & ~n_14530;
assign n_14532 =  x_2270 &  n_14531;
assign n_14533 = ~x_2270 & ~n_14531;
assign n_14534 = ~n_14532 & ~n_14533;
assign n_14535 =  x_2269 & ~n_1761;
assign n_14536 =  i_204 &  n_1751;
assign n_14537 =  n_1761 &  n_14536;
assign n_14538 = ~n_14535 & ~n_14537;
assign n_14539 =  x_2269 & ~n_14538;
assign n_14540 = ~x_2269 &  n_14538;
assign n_14541 = ~n_14539 & ~n_14540;
assign n_14542 =  x_2268 & ~n_1770;
assign n_14543 =  n_1770 &  n_14536;
assign n_14544 = ~n_14542 & ~n_14543;
assign n_14545 =  x_2268 & ~n_14544;
assign n_14546 = ~x_2268 &  n_14544;
assign n_14547 = ~n_14545 & ~n_14546;
assign n_14548 =  x_2267 & ~n_1778;
assign n_14549 =  n_1778 &  n_14536;
assign n_14550 = ~n_14548 & ~n_14549;
assign n_14551 =  x_2267 & ~n_14550;
assign n_14552 = ~x_2267 &  n_14550;
assign n_14553 = ~n_14551 & ~n_14552;
assign n_14554 =  x_2266 & ~n_1785;
assign n_14555 =  n_1785 &  n_14536;
assign n_14556 = ~n_14554 & ~n_14555;
assign n_14557 =  x_2266 & ~n_14556;
assign n_14558 = ~x_2266 &  n_14556;
assign n_14559 = ~n_14557 & ~n_14558;
assign n_14560 =  x_2265 & ~n_1792;
assign n_14561 =  n_1792 &  n_14536;
assign n_14562 = ~n_14560 & ~n_14561;
assign n_14563 =  x_2265 & ~n_14562;
assign n_14564 = ~x_2265 &  n_14562;
assign n_14565 = ~n_14563 & ~n_14564;
assign n_14566 =  x_2264 & ~n_1799;
assign n_14567 =  n_1799 &  n_14536;
assign n_14568 = ~n_14566 & ~n_14567;
assign n_14569 =  x_2264 & ~n_14568;
assign n_14570 = ~x_2264 &  n_14568;
assign n_14571 = ~n_14569 & ~n_14570;
assign n_14572 =  x_2263 & ~n_1806;
assign n_14573 =  n_1806 &  n_14536;
assign n_14574 = ~n_14572 & ~n_14573;
assign n_14575 =  x_2263 & ~n_14574;
assign n_14576 = ~x_2263 &  n_14574;
assign n_14577 = ~n_14575 & ~n_14576;
assign n_14578 =  n_1750 & ~n_14536;
assign n_14579 = ~x_2262 & ~n_1750;
assign n_14580 = ~n_14578 & ~n_14579;
assign n_14581 =  x_2262 &  n_14580;
assign n_14582 = ~x_2262 & ~n_14580;
assign n_14583 = ~n_14581 & ~n_14582;
assign n_14584 =  x_2261 & ~n_1761;
assign n_14585 =  i_203 &  n_1751;
assign n_14586 =  n_1761 &  n_14585;
assign n_14587 = ~n_14584 & ~n_14586;
assign n_14588 =  x_2261 & ~n_14587;
assign n_14589 = ~x_2261 &  n_14587;
assign n_14590 = ~n_14588 & ~n_14589;
assign n_14591 =  x_2260 & ~n_1770;
assign n_14592 =  n_1770 &  n_14585;
assign n_14593 = ~n_14591 & ~n_14592;
assign n_14594 =  x_2260 & ~n_14593;
assign n_14595 = ~x_2260 &  n_14593;
assign n_14596 = ~n_14594 & ~n_14595;
assign n_14597 =  x_2259 & ~n_1778;
assign n_14598 =  n_1778 &  n_14585;
assign n_14599 = ~n_14597 & ~n_14598;
assign n_14600 =  x_2259 & ~n_14599;
assign n_14601 = ~x_2259 &  n_14599;
assign n_14602 = ~n_14600 & ~n_14601;
assign n_14603 =  x_2258 & ~n_1785;
assign n_14604 =  n_1785 &  n_14585;
assign n_14605 = ~n_14603 & ~n_14604;
assign n_14606 =  x_2258 & ~n_14605;
assign n_14607 = ~x_2258 &  n_14605;
assign n_14608 = ~n_14606 & ~n_14607;
assign n_14609 =  x_2257 & ~n_1792;
assign n_14610 =  n_1792 &  n_14585;
assign n_14611 = ~n_14609 & ~n_14610;
assign n_14612 =  x_2257 & ~n_14611;
assign n_14613 = ~x_2257 &  n_14611;
assign n_14614 = ~n_14612 & ~n_14613;
assign n_14615 =  x_2256 & ~n_1799;
assign n_14616 =  n_1799 &  n_14585;
assign n_14617 = ~n_14615 & ~n_14616;
assign n_14618 =  x_2256 & ~n_14617;
assign n_14619 = ~x_2256 &  n_14617;
assign n_14620 = ~n_14618 & ~n_14619;
assign n_14621 =  x_2255 & ~n_1806;
assign n_14622 =  n_1806 &  n_14585;
assign n_14623 = ~n_14621 & ~n_14622;
assign n_14624 =  x_2255 & ~n_14623;
assign n_14625 = ~x_2255 &  n_14623;
assign n_14626 = ~n_14624 & ~n_14625;
assign n_14627 =  n_1750 & ~n_14585;
assign n_14628 = ~x_2254 & ~n_1750;
assign n_14629 = ~n_14627 & ~n_14628;
assign n_14630 =  x_2254 &  n_14629;
assign n_14631 = ~x_2254 & ~n_14629;
assign n_14632 = ~n_14630 & ~n_14631;
assign n_14633 =  x_2253 & ~n_1761;
assign n_14634 =  i_202 &  n_1751;
assign n_14635 =  n_1761 &  n_14634;
assign n_14636 = ~n_14633 & ~n_14635;
assign n_14637 =  x_2253 & ~n_14636;
assign n_14638 = ~x_2253 &  n_14636;
assign n_14639 = ~n_14637 & ~n_14638;
assign n_14640 =  x_2252 & ~n_1770;
assign n_14641 =  n_1770 &  n_14634;
assign n_14642 = ~n_14640 & ~n_14641;
assign n_14643 =  x_2252 & ~n_14642;
assign n_14644 = ~x_2252 &  n_14642;
assign n_14645 = ~n_14643 & ~n_14644;
assign n_14646 =  x_2251 & ~n_1778;
assign n_14647 =  n_1778 &  n_14634;
assign n_14648 = ~n_14646 & ~n_14647;
assign n_14649 =  x_2251 & ~n_14648;
assign n_14650 = ~x_2251 &  n_14648;
assign n_14651 = ~n_14649 & ~n_14650;
assign n_14652 =  x_2250 & ~n_1785;
assign n_14653 =  n_1785 &  n_14634;
assign n_14654 = ~n_14652 & ~n_14653;
assign n_14655 =  x_2250 & ~n_14654;
assign n_14656 = ~x_2250 &  n_14654;
assign n_14657 = ~n_14655 & ~n_14656;
assign n_14658 =  x_2249 & ~n_1792;
assign n_14659 =  n_1792 &  n_14634;
assign n_14660 = ~n_14658 & ~n_14659;
assign n_14661 =  x_2249 & ~n_14660;
assign n_14662 = ~x_2249 &  n_14660;
assign n_14663 = ~n_14661 & ~n_14662;
assign n_14664 =  x_2248 & ~n_1799;
assign n_14665 =  n_1799 &  n_14634;
assign n_14666 = ~n_14664 & ~n_14665;
assign n_14667 =  x_2248 & ~n_14666;
assign n_14668 = ~x_2248 &  n_14666;
assign n_14669 = ~n_14667 & ~n_14668;
assign n_14670 =  x_2247 & ~n_1806;
assign n_14671 =  n_1806 &  n_14634;
assign n_14672 = ~n_14670 & ~n_14671;
assign n_14673 =  x_2247 & ~n_14672;
assign n_14674 = ~x_2247 &  n_14672;
assign n_14675 = ~n_14673 & ~n_14674;
assign n_14676 =  n_1750 & ~n_14634;
assign n_14677 = ~x_2246 & ~n_1750;
assign n_14678 = ~n_14676 & ~n_14677;
assign n_14679 =  x_2246 &  n_14678;
assign n_14680 = ~x_2246 & ~n_14678;
assign n_14681 = ~n_14679 & ~n_14680;
assign n_14682 =  x_2245 & ~n_1761;
assign n_14683 =  i_201 &  n_1751;
assign n_14684 =  n_1761 &  n_14683;
assign n_14685 = ~n_14682 & ~n_14684;
assign n_14686 =  x_2245 & ~n_14685;
assign n_14687 = ~x_2245 &  n_14685;
assign n_14688 = ~n_14686 & ~n_14687;
assign n_14689 =  x_2244 & ~n_1770;
assign n_14690 =  n_1770 &  n_14683;
assign n_14691 = ~n_14689 & ~n_14690;
assign n_14692 =  x_2244 & ~n_14691;
assign n_14693 = ~x_2244 &  n_14691;
assign n_14694 = ~n_14692 & ~n_14693;
assign n_14695 =  x_2243 & ~n_1778;
assign n_14696 =  n_1778 &  n_14683;
assign n_14697 = ~n_14695 & ~n_14696;
assign n_14698 =  x_2243 & ~n_14697;
assign n_14699 = ~x_2243 &  n_14697;
assign n_14700 = ~n_14698 & ~n_14699;
assign n_14701 =  x_2242 & ~n_1785;
assign n_14702 =  n_1785 &  n_14683;
assign n_14703 = ~n_14701 & ~n_14702;
assign n_14704 =  x_2242 & ~n_14703;
assign n_14705 = ~x_2242 &  n_14703;
assign n_14706 = ~n_14704 & ~n_14705;
assign n_14707 =  x_2241 & ~n_1792;
assign n_14708 =  n_1792 &  n_14683;
assign n_14709 = ~n_14707 & ~n_14708;
assign n_14710 =  x_2241 & ~n_14709;
assign n_14711 = ~x_2241 &  n_14709;
assign n_14712 = ~n_14710 & ~n_14711;
assign n_14713 =  x_2240 & ~n_1799;
assign n_14714 =  n_1799 &  n_14683;
assign n_14715 = ~n_14713 & ~n_14714;
assign n_14716 =  x_2240 & ~n_14715;
assign n_14717 = ~x_2240 &  n_14715;
assign n_14718 = ~n_14716 & ~n_14717;
assign n_14719 =  x_2239 & ~n_1806;
assign n_14720 =  n_1806 &  n_14683;
assign n_14721 = ~n_14719 & ~n_14720;
assign n_14722 =  x_2239 & ~n_14721;
assign n_14723 = ~x_2239 &  n_14721;
assign n_14724 = ~n_14722 & ~n_14723;
assign n_14725 =  n_1750 & ~n_14683;
assign n_14726 = ~x_2238 & ~n_1750;
assign n_14727 = ~n_14725 & ~n_14726;
assign n_14728 =  x_2238 &  n_14727;
assign n_14729 = ~x_2238 & ~n_14727;
assign n_14730 = ~n_14728 & ~n_14729;
assign n_14731 =  x_2237 & ~n_1761;
assign n_14732 =  i_200 &  n_1751;
assign n_14733 =  n_1761 &  n_14732;
assign n_14734 = ~n_14731 & ~n_14733;
assign n_14735 =  x_2237 & ~n_14734;
assign n_14736 = ~x_2237 &  n_14734;
assign n_14737 = ~n_14735 & ~n_14736;
assign n_14738 =  x_2236 & ~n_1770;
assign n_14739 =  n_1770 &  n_14732;
assign n_14740 = ~n_14738 & ~n_14739;
assign n_14741 =  x_2236 & ~n_14740;
assign n_14742 = ~x_2236 &  n_14740;
assign n_14743 = ~n_14741 & ~n_14742;
assign n_14744 =  x_2235 & ~n_1778;
assign n_14745 =  n_1778 &  n_14732;
assign n_14746 = ~n_14744 & ~n_14745;
assign n_14747 =  x_2235 & ~n_14746;
assign n_14748 = ~x_2235 &  n_14746;
assign n_14749 = ~n_14747 & ~n_14748;
assign n_14750 =  x_2234 & ~n_1785;
assign n_14751 =  n_1785 &  n_14732;
assign n_14752 = ~n_14750 & ~n_14751;
assign n_14753 =  x_2234 & ~n_14752;
assign n_14754 = ~x_2234 &  n_14752;
assign n_14755 = ~n_14753 & ~n_14754;
assign n_14756 =  x_2233 & ~n_1792;
assign n_14757 =  n_1792 &  n_14732;
assign n_14758 = ~n_14756 & ~n_14757;
assign n_14759 =  x_2233 & ~n_14758;
assign n_14760 = ~x_2233 &  n_14758;
assign n_14761 = ~n_14759 & ~n_14760;
assign n_14762 =  x_2232 & ~n_1799;
assign n_14763 =  n_1799 &  n_14732;
assign n_14764 = ~n_14762 & ~n_14763;
assign n_14765 =  x_2232 & ~n_14764;
assign n_14766 = ~x_2232 &  n_14764;
assign n_14767 = ~n_14765 & ~n_14766;
assign n_14768 =  x_2231 & ~n_1806;
assign n_14769 =  n_1806 &  n_14732;
assign n_14770 = ~n_14768 & ~n_14769;
assign n_14771 =  x_2231 & ~n_14770;
assign n_14772 = ~x_2231 &  n_14770;
assign n_14773 = ~n_14771 & ~n_14772;
assign n_14774 =  n_1750 & ~n_14732;
assign n_14775 = ~x_2230 & ~n_1750;
assign n_14776 = ~n_14774 & ~n_14775;
assign n_14777 =  x_2230 &  n_14776;
assign n_14778 = ~x_2230 & ~n_14776;
assign n_14779 = ~n_14777 & ~n_14778;
assign n_14780 =  x_2229 & ~n_1761;
assign n_14781 =  i_199 &  n_1751;
assign n_14782 =  n_1761 &  n_14781;
assign n_14783 = ~n_14780 & ~n_14782;
assign n_14784 =  x_2229 & ~n_14783;
assign n_14785 = ~x_2229 &  n_14783;
assign n_14786 = ~n_14784 & ~n_14785;
assign n_14787 =  x_2228 & ~n_1770;
assign n_14788 =  n_1770 &  n_14781;
assign n_14789 = ~n_14787 & ~n_14788;
assign n_14790 =  x_2228 & ~n_14789;
assign n_14791 = ~x_2228 &  n_14789;
assign n_14792 = ~n_14790 & ~n_14791;
assign n_14793 =  x_2227 & ~n_1778;
assign n_14794 =  n_1778 &  n_14781;
assign n_14795 = ~n_14793 & ~n_14794;
assign n_14796 =  x_2227 & ~n_14795;
assign n_14797 = ~x_2227 &  n_14795;
assign n_14798 = ~n_14796 & ~n_14797;
assign n_14799 =  x_2226 & ~n_1785;
assign n_14800 =  n_1785 &  n_14781;
assign n_14801 = ~n_14799 & ~n_14800;
assign n_14802 =  x_2226 & ~n_14801;
assign n_14803 = ~x_2226 &  n_14801;
assign n_14804 = ~n_14802 & ~n_14803;
assign n_14805 =  x_2225 & ~n_1792;
assign n_14806 =  n_1792 &  n_14781;
assign n_14807 = ~n_14805 & ~n_14806;
assign n_14808 =  x_2225 & ~n_14807;
assign n_14809 = ~x_2225 &  n_14807;
assign n_14810 = ~n_14808 & ~n_14809;
assign n_14811 =  x_2224 & ~n_1799;
assign n_14812 =  n_1799 &  n_14781;
assign n_14813 = ~n_14811 & ~n_14812;
assign n_14814 =  x_2224 & ~n_14813;
assign n_14815 = ~x_2224 &  n_14813;
assign n_14816 = ~n_14814 & ~n_14815;
assign n_14817 =  x_2223 & ~n_1806;
assign n_14818 =  n_1806 &  n_14781;
assign n_14819 = ~n_14817 & ~n_14818;
assign n_14820 =  x_2223 & ~n_14819;
assign n_14821 = ~x_2223 &  n_14819;
assign n_14822 = ~n_14820 & ~n_14821;
assign n_14823 =  n_1750 & ~n_14781;
assign n_14824 = ~x_2222 & ~n_1750;
assign n_14825 = ~n_14823 & ~n_14824;
assign n_14826 =  x_2222 &  n_14825;
assign n_14827 = ~x_2222 & ~n_14825;
assign n_14828 = ~n_14826 & ~n_14827;
assign n_14829 =  x_2221 & ~n_1761;
assign n_14830 =  i_198 &  n_1751;
assign n_14831 =  n_1761 &  n_14830;
assign n_14832 = ~n_14829 & ~n_14831;
assign n_14833 =  x_2221 & ~n_14832;
assign n_14834 = ~x_2221 &  n_14832;
assign n_14835 = ~n_14833 & ~n_14834;
assign n_14836 =  x_2220 & ~n_1770;
assign n_14837 =  n_1770 &  n_14830;
assign n_14838 = ~n_14836 & ~n_14837;
assign n_14839 =  x_2220 & ~n_14838;
assign n_14840 = ~x_2220 &  n_14838;
assign n_14841 = ~n_14839 & ~n_14840;
assign n_14842 =  x_2219 & ~n_1778;
assign n_14843 =  n_1778 &  n_14830;
assign n_14844 = ~n_14842 & ~n_14843;
assign n_14845 =  x_2219 & ~n_14844;
assign n_14846 = ~x_2219 &  n_14844;
assign n_14847 = ~n_14845 & ~n_14846;
assign n_14848 =  x_2218 & ~n_1785;
assign n_14849 =  n_1785 &  n_14830;
assign n_14850 = ~n_14848 & ~n_14849;
assign n_14851 =  x_2218 & ~n_14850;
assign n_14852 = ~x_2218 &  n_14850;
assign n_14853 = ~n_14851 & ~n_14852;
assign n_14854 =  x_2217 & ~n_1792;
assign n_14855 =  n_1792 &  n_14830;
assign n_14856 = ~n_14854 & ~n_14855;
assign n_14857 =  x_2217 & ~n_14856;
assign n_14858 = ~x_2217 &  n_14856;
assign n_14859 = ~n_14857 & ~n_14858;
assign n_14860 =  x_2216 & ~n_1799;
assign n_14861 =  n_1799 &  n_14830;
assign n_14862 = ~n_14860 & ~n_14861;
assign n_14863 =  x_2216 & ~n_14862;
assign n_14864 = ~x_2216 &  n_14862;
assign n_14865 = ~n_14863 & ~n_14864;
assign n_14866 =  x_2215 & ~n_1806;
assign n_14867 =  n_1806 &  n_14830;
assign n_14868 = ~n_14866 & ~n_14867;
assign n_14869 =  x_2215 & ~n_14868;
assign n_14870 = ~x_2215 &  n_14868;
assign n_14871 = ~n_14869 & ~n_14870;
assign n_14872 =  n_1750 & ~n_14830;
assign n_14873 = ~x_2214 & ~n_1750;
assign n_14874 = ~n_14872 & ~n_14873;
assign n_14875 =  x_2214 &  n_14874;
assign n_14876 = ~x_2214 & ~n_14874;
assign n_14877 = ~n_14875 & ~n_14876;
assign n_14878 =  x_2213 & ~n_1761;
assign n_14879 =  i_197 &  n_1751;
assign n_14880 =  n_1761 &  n_14879;
assign n_14881 = ~n_14878 & ~n_14880;
assign n_14882 =  x_2213 & ~n_14881;
assign n_14883 = ~x_2213 &  n_14881;
assign n_14884 = ~n_14882 & ~n_14883;
assign n_14885 =  x_2212 & ~n_1770;
assign n_14886 =  n_1770 &  n_14879;
assign n_14887 = ~n_14885 & ~n_14886;
assign n_14888 =  x_2212 & ~n_14887;
assign n_14889 = ~x_2212 &  n_14887;
assign n_14890 = ~n_14888 & ~n_14889;
assign n_14891 =  x_2211 & ~n_1778;
assign n_14892 =  n_1778 &  n_14879;
assign n_14893 = ~n_14891 & ~n_14892;
assign n_14894 =  x_2211 & ~n_14893;
assign n_14895 = ~x_2211 &  n_14893;
assign n_14896 = ~n_14894 & ~n_14895;
assign n_14897 =  x_2210 & ~n_1785;
assign n_14898 =  n_1785 &  n_14879;
assign n_14899 = ~n_14897 & ~n_14898;
assign n_14900 =  x_2210 & ~n_14899;
assign n_14901 = ~x_2210 &  n_14899;
assign n_14902 = ~n_14900 & ~n_14901;
assign n_14903 =  x_2209 & ~n_1792;
assign n_14904 =  n_1792 &  n_14879;
assign n_14905 = ~n_14903 & ~n_14904;
assign n_14906 =  x_2209 & ~n_14905;
assign n_14907 = ~x_2209 &  n_14905;
assign n_14908 = ~n_14906 & ~n_14907;
assign n_14909 =  x_2208 & ~n_1799;
assign n_14910 =  n_1799 &  n_14879;
assign n_14911 = ~n_14909 & ~n_14910;
assign n_14912 =  x_2208 & ~n_14911;
assign n_14913 = ~x_2208 &  n_14911;
assign n_14914 = ~n_14912 & ~n_14913;
assign n_14915 =  x_2207 & ~n_1806;
assign n_14916 =  n_1806 &  n_14879;
assign n_14917 = ~n_14915 & ~n_14916;
assign n_14918 =  x_2207 & ~n_14917;
assign n_14919 = ~x_2207 &  n_14917;
assign n_14920 = ~n_14918 & ~n_14919;
assign n_14921 =  n_1750 & ~n_14879;
assign n_14922 = ~x_2206 & ~n_1750;
assign n_14923 = ~n_14921 & ~n_14922;
assign n_14924 =  x_2206 &  n_14923;
assign n_14925 = ~x_2206 & ~n_14923;
assign n_14926 = ~n_14924 & ~n_14925;
assign n_14927 =  x_2205 & ~n_1761;
assign n_14928 =  i_196 &  n_1751;
assign n_14929 =  n_1761 &  n_14928;
assign n_14930 = ~n_14927 & ~n_14929;
assign n_14931 =  x_2205 & ~n_14930;
assign n_14932 = ~x_2205 &  n_14930;
assign n_14933 = ~n_14931 & ~n_14932;
assign n_14934 =  x_2204 & ~n_1770;
assign n_14935 =  n_1770 &  n_14928;
assign n_14936 = ~n_14934 & ~n_14935;
assign n_14937 =  x_2204 & ~n_14936;
assign n_14938 = ~x_2204 &  n_14936;
assign n_14939 = ~n_14937 & ~n_14938;
assign n_14940 =  x_2203 & ~n_1778;
assign n_14941 =  n_1778 &  n_14928;
assign n_14942 = ~n_14940 & ~n_14941;
assign n_14943 =  x_2203 & ~n_14942;
assign n_14944 = ~x_2203 &  n_14942;
assign n_14945 = ~n_14943 & ~n_14944;
assign n_14946 =  x_2202 & ~n_1785;
assign n_14947 =  n_1785 &  n_14928;
assign n_14948 = ~n_14946 & ~n_14947;
assign n_14949 =  x_2202 & ~n_14948;
assign n_14950 = ~x_2202 &  n_14948;
assign n_14951 = ~n_14949 & ~n_14950;
assign n_14952 =  x_2201 & ~n_1792;
assign n_14953 =  n_1792 &  n_14928;
assign n_14954 = ~n_14952 & ~n_14953;
assign n_14955 =  x_2201 & ~n_14954;
assign n_14956 = ~x_2201 &  n_14954;
assign n_14957 = ~n_14955 & ~n_14956;
assign n_14958 =  x_2200 & ~n_1799;
assign n_14959 =  n_1799 &  n_14928;
assign n_14960 = ~n_14958 & ~n_14959;
assign n_14961 =  x_2200 & ~n_14960;
assign n_14962 = ~x_2200 &  n_14960;
assign n_14963 = ~n_14961 & ~n_14962;
assign n_14964 =  x_2199 & ~n_1806;
assign n_14965 =  n_1806 &  n_14928;
assign n_14966 = ~n_14964 & ~n_14965;
assign n_14967 =  x_2199 & ~n_14966;
assign n_14968 = ~x_2199 &  n_14966;
assign n_14969 = ~n_14967 & ~n_14968;
assign n_14970 =  n_1750 & ~n_14928;
assign n_14971 = ~x_2198 & ~n_1750;
assign n_14972 = ~n_14970 & ~n_14971;
assign n_14973 =  x_2198 &  n_14972;
assign n_14974 = ~x_2198 & ~n_14972;
assign n_14975 = ~n_14973 & ~n_14974;
assign n_14976 =  x_2197 & ~n_1761;
assign n_14977 =  i_195 &  n_1751;
assign n_14978 =  n_1761 &  n_14977;
assign n_14979 = ~n_14976 & ~n_14978;
assign n_14980 =  x_2197 & ~n_14979;
assign n_14981 = ~x_2197 &  n_14979;
assign n_14982 = ~n_14980 & ~n_14981;
assign n_14983 =  x_2196 & ~n_1770;
assign n_14984 =  n_1770 &  n_14977;
assign n_14985 = ~n_14983 & ~n_14984;
assign n_14986 =  x_2196 & ~n_14985;
assign n_14987 = ~x_2196 &  n_14985;
assign n_14988 = ~n_14986 & ~n_14987;
assign n_14989 =  x_2195 & ~n_1778;
assign n_14990 =  n_1778 &  n_14977;
assign n_14991 = ~n_14989 & ~n_14990;
assign n_14992 =  x_2195 & ~n_14991;
assign n_14993 = ~x_2195 &  n_14991;
assign n_14994 = ~n_14992 & ~n_14993;
assign n_14995 =  x_2194 & ~n_1785;
assign n_14996 =  n_1785 &  n_14977;
assign n_14997 = ~n_14995 & ~n_14996;
assign n_14998 =  x_2194 & ~n_14997;
assign n_14999 = ~x_2194 &  n_14997;
assign n_15000 = ~n_14998 & ~n_14999;
assign n_15001 =  x_2193 & ~n_1792;
assign n_15002 =  n_1792 &  n_14977;
assign n_15003 = ~n_15001 & ~n_15002;
assign n_15004 =  x_2193 & ~n_15003;
assign n_15005 = ~x_2193 &  n_15003;
assign n_15006 = ~n_15004 & ~n_15005;
assign n_15007 =  x_2192 & ~n_1799;
assign n_15008 =  n_1799 &  n_14977;
assign n_15009 = ~n_15007 & ~n_15008;
assign n_15010 =  x_2192 & ~n_15009;
assign n_15011 = ~x_2192 &  n_15009;
assign n_15012 = ~n_15010 & ~n_15011;
assign n_15013 =  x_2191 & ~n_1806;
assign n_15014 =  n_1806 &  n_14977;
assign n_15015 = ~n_15013 & ~n_15014;
assign n_15016 =  x_2191 & ~n_15015;
assign n_15017 = ~x_2191 &  n_15015;
assign n_15018 = ~n_15016 & ~n_15017;
assign n_15019 =  n_1750 & ~n_14977;
assign n_15020 = ~x_2190 & ~n_1750;
assign n_15021 = ~n_15019 & ~n_15020;
assign n_15022 =  x_2190 &  n_15021;
assign n_15023 = ~x_2190 & ~n_15021;
assign n_15024 = ~n_15022 & ~n_15023;
assign n_15025 =  x_2189 & ~n_1761;
assign n_15026 =  i_194 &  n_1751;
assign n_15027 =  n_1761 &  n_15026;
assign n_15028 = ~n_15025 & ~n_15027;
assign n_15029 =  x_2189 & ~n_15028;
assign n_15030 = ~x_2189 &  n_15028;
assign n_15031 = ~n_15029 & ~n_15030;
assign n_15032 =  x_2188 & ~n_1770;
assign n_15033 =  n_1770 &  n_15026;
assign n_15034 = ~n_15032 & ~n_15033;
assign n_15035 =  x_2188 & ~n_15034;
assign n_15036 = ~x_2188 &  n_15034;
assign n_15037 = ~n_15035 & ~n_15036;
assign n_15038 =  x_2187 & ~n_1778;
assign n_15039 =  n_1778 &  n_15026;
assign n_15040 = ~n_15038 & ~n_15039;
assign n_15041 =  x_2187 & ~n_15040;
assign n_15042 = ~x_2187 &  n_15040;
assign n_15043 = ~n_15041 & ~n_15042;
assign n_15044 =  x_2186 & ~n_1785;
assign n_15045 =  n_1785 &  n_15026;
assign n_15046 = ~n_15044 & ~n_15045;
assign n_15047 =  x_2186 & ~n_15046;
assign n_15048 = ~x_2186 &  n_15046;
assign n_15049 = ~n_15047 & ~n_15048;
assign n_15050 =  x_2185 & ~n_1792;
assign n_15051 =  n_1792 &  n_15026;
assign n_15052 = ~n_15050 & ~n_15051;
assign n_15053 =  x_2185 & ~n_15052;
assign n_15054 = ~x_2185 &  n_15052;
assign n_15055 = ~n_15053 & ~n_15054;
assign n_15056 =  x_2184 & ~n_1799;
assign n_15057 =  n_1799 &  n_15026;
assign n_15058 = ~n_15056 & ~n_15057;
assign n_15059 =  x_2184 & ~n_15058;
assign n_15060 = ~x_2184 &  n_15058;
assign n_15061 = ~n_15059 & ~n_15060;
assign n_15062 =  x_2183 & ~n_1806;
assign n_15063 =  n_1806 &  n_15026;
assign n_15064 = ~n_15062 & ~n_15063;
assign n_15065 =  x_2183 & ~n_15064;
assign n_15066 = ~x_2183 &  n_15064;
assign n_15067 = ~n_15065 & ~n_15066;
assign n_15068 =  n_1750 & ~n_15026;
assign n_15069 = ~x_2182 & ~n_1750;
assign n_15070 = ~n_15068 & ~n_15069;
assign n_15071 =  x_2182 &  n_15070;
assign n_15072 = ~x_2182 & ~n_15070;
assign n_15073 = ~n_15071 & ~n_15072;
assign n_15074 =  x_2181 & ~n_1761;
assign n_15075 =  i_193 &  n_1751;
assign n_15076 =  n_1761 &  n_15075;
assign n_15077 = ~n_15074 & ~n_15076;
assign n_15078 =  x_2181 & ~n_15077;
assign n_15079 = ~x_2181 &  n_15077;
assign n_15080 = ~n_15078 & ~n_15079;
assign n_15081 =  x_2180 & ~n_1770;
assign n_15082 =  n_1770 &  n_15075;
assign n_15083 = ~n_15081 & ~n_15082;
assign n_15084 =  x_2180 & ~n_15083;
assign n_15085 = ~x_2180 &  n_15083;
assign n_15086 = ~n_15084 & ~n_15085;
assign n_15087 =  x_2179 & ~n_1778;
assign n_15088 =  n_1778 &  n_15075;
assign n_15089 = ~n_15087 & ~n_15088;
assign n_15090 =  x_2179 & ~n_15089;
assign n_15091 = ~x_2179 &  n_15089;
assign n_15092 = ~n_15090 & ~n_15091;
assign n_15093 =  x_2178 & ~n_1785;
assign n_15094 =  n_1785 &  n_15075;
assign n_15095 = ~n_15093 & ~n_15094;
assign n_15096 =  x_2178 & ~n_15095;
assign n_15097 = ~x_2178 &  n_15095;
assign n_15098 = ~n_15096 & ~n_15097;
assign n_15099 =  x_2177 & ~n_1792;
assign n_15100 =  n_1792 &  n_15075;
assign n_15101 = ~n_15099 & ~n_15100;
assign n_15102 =  x_2177 & ~n_15101;
assign n_15103 = ~x_2177 &  n_15101;
assign n_15104 = ~n_15102 & ~n_15103;
assign n_15105 =  x_2176 & ~n_1799;
assign n_15106 =  n_1799 &  n_15075;
assign n_15107 = ~n_15105 & ~n_15106;
assign n_15108 =  x_2176 & ~n_15107;
assign n_15109 = ~x_2176 &  n_15107;
assign n_15110 = ~n_15108 & ~n_15109;
assign n_15111 =  x_2175 & ~n_1806;
assign n_15112 =  n_1806 &  n_15075;
assign n_15113 = ~n_15111 & ~n_15112;
assign n_15114 =  x_2175 & ~n_15113;
assign n_15115 = ~x_2175 &  n_15113;
assign n_15116 = ~n_15114 & ~n_15115;
assign n_15117 =  n_1750 & ~n_15075;
assign n_15118 = ~x_2174 & ~n_1750;
assign n_15119 = ~n_15117 & ~n_15118;
assign n_15120 =  x_2174 &  n_15119;
assign n_15121 = ~x_2174 & ~n_15119;
assign n_15122 = ~n_15120 & ~n_15121;
assign n_15123 =  x_2173 & ~n_1761;
assign n_15124 =  i_192 &  n_1751;
assign n_15125 =  n_1761 &  n_15124;
assign n_15126 = ~n_15123 & ~n_15125;
assign n_15127 =  x_2173 & ~n_15126;
assign n_15128 = ~x_2173 &  n_15126;
assign n_15129 = ~n_15127 & ~n_15128;
assign n_15130 =  x_2172 & ~n_1770;
assign n_15131 =  n_1770 &  n_15124;
assign n_15132 = ~n_15130 & ~n_15131;
assign n_15133 =  x_2172 & ~n_15132;
assign n_15134 = ~x_2172 &  n_15132;
assign n_15135 = ~n_15133 & ~n_15134;
assign n_15136 =  x_2171 & ~n_1778;
assign n_15137 =  n_1778 &  n_15124;
assign n_15138 = ~n_15136 & ~n_15137;
assign n_15139 =  x_2171 & ~n_15138;
assign n_15140 = ~x_2171 &  n_15138;
assign n_15141 = ~n_15139 & ~n_15140;
assign n_15142 =  x_2170 & ~n_1785;
assign n_15143 =  n_1785 &  n_15124;
assign n_15144 = ~n_15142 & ~n_15143;
assign n_15145 =  x_2170 & ~n_15144;
assign n_15146 = ~x_2170 &  n_15144;
assign n_15147 = ~n_15145 & ~n_15146;
assign n_15148 =  x_2169 & ~n_1792;
assign n_15149 =  n_1792 &  n_15124;
assign n_15150 = ~n_15148 & ~n_15149;
assign n_15151 =  x_2169 & ~n_15150;
assign n_15152 = ~x_2169 &  n_15150;
assign n_15153 = ~n_15151 & ~n_15152;
assign n_15154 =  x_2168 & ~n_1799;
assign n_15155 =  n_1799 &  n_15124;
assign n_15156 = ~n_15154 & ~n_15155;
assign n_15157 =  x_2168 & ~n_15156;
assign n_15158 = ~x_2168 &  n_15156;
assign n_15159 = ~n_15157 & ~n_15158;
assign n_15160 =  x_2167 & ~n_1806;
assign n_15161 =  n_1806 &  n_15124;
assign n_15162 = ~n_15160 & ~n_15161;
assign n_15163 =  x_2167 & ~n_15162;
assign n_15164 = ~x_2167 &  n_15162;
assign n_15165 = ~n_15163 & ~n_15164;
assign n_15166 =  n_1750 & ~n_15124;
assign n_15167 = ~x_2166 & ~n_1750;
assign n_15168 = ~n_15166 & ~n_15167;
assign n_15169 =  x_2166 &  n_15168;
assign n_15170 = ~x_2166 & ~n_15168;
assign n_15171 = ~n_15169 & ~n_15170;
assign n_15172 =  x_2165 & ~n_1761;
assign n_15173 =  n_1761 &  n_1752;
assign n_15174 = ~n_15172 & ~n_15173;
assign n_15175 =  x_2165 & ~n_15174;
assign n_15176 = ~x_2165 &  n_15174;
assign n_15177 = ~n_15175 & ~n_15176;
assign n_15178 =  x_2164 & ~n_1770;
assign n_15179 =  n_1770 &  n_1752;
assign n_15180 = ~n_15178 & ~n_15179;
assign n_15181 =  x_2164 & ~n_15180;
assign n_15182 = ~x_2164 &  n_15180;
assign n_15183 = ~n_15181 & ~n_15182;
assign n_15184 =  x_2163 & ~n_1778;
assign n_15185 =  n_1778 &  n_1752;
assign n_15186 = ~n_15184 & ~n_15185;
assign n_15187 =  x_2163 & ~n_15186;
assign n_15188 = ~x_2163 &  n_15186;
assign n_15189 = ~n_15187 & ~n_15188;
assign n_15190 =  x_2162 & ~n_1785;
assign n_15191 =  n_1785 &  n_1752;
assign n_15192 = ~n_15190 & ~n_15191;
assign n_15193 =  x_2162 & ~n_15192;
assign n_15194 = ~x_2162 &  n_15192;
assign n_15195 = ~n_15193 & ~n_15194;
assign n_15196 =  x_2161 & ~n_1792;
assign n_15197 =  n_1792 &  n_1752;
assign n_15198 = ~n_15196 & ~n_15197;
assign n_15199 =  x_2161 & ~n_15198;
assign n_15200 = ~x_2161 &  n_15198;
assign n_15201 = ~n_15199 & ~n_15200;
assign n_15202 =  x_2160 & ~n_1799;
assign n_15203 =  n_1799 &  n_1752;
assign n_15204 = ~n_15202 & ~n_15203;
assign n_15205 =  x_2160 & ~n_15204;
assign n_15206 = ~x_2160 &  n_15204;
assign n_15207 = ~n_15205 & ~n_15206;
assign n_15208 =  x_2159 & ~n_1806;
assign n_15209 =  n_1806 &  n_1752;
assign n_15210 = ~n_15208 & ~n_15209;
assign n_15211 =  x_2159 & ~n_15210;
assign n_15212 = ~x_2159 &  n_15210;
assign n_15213 = ~n_15211 & ~n_15212;
assign n_15214 =  x_1883 & ~n_1806;
assign n_15215 =  n_1806 &  n_3481;
assign n_15216 = ~n_15214 & ~n_15215;
assign n_15217 =  x_1883 & ~n_15216;
assign n_15218 = ~x_1883 &  n_15216;
assign n_15219 = ~n_15217 & ~n_15218;
assign n_15220 =  n_1750 & ~n_3481;
assign n_15221 = ~x_1882 & ~n_1750;
assign n_15222 = ~n_15220 & ~n_15221;
assign n_15223 =  x_1882 &  n_15222;
assign n_15224 = ~x_1882 & ~n_15222;
assign n_15225 = ~n_15223 & ~n_15224;
assign n_15226 =  x_1881 &  n_3308;
assign n_15227 =  x_448 &  n_3307;
assign n_15228 = ~n_15226 & ~n_15227;
assign n_15229 =  x_1881 & ~n_15228;
assign n_15230 = ~x_1881 &  n_15228;
assign n_15231 = ~n_15229 & ~n_15230;
assign n_15232 =  x_1880 & ~n_1761;
assign n_15233 =  i_156 &  n_1751;
assign n_15234 =  n_1761 &  n_15233;
assign n_15235 = ~n_15232 & ~n_15234;
assign n_15236 =  x_1880 & ~n_15235;
assign n_15237 = ~x_1880 &  n_15235;
assign n_15238 = ~n_15236 & ~n_15237;
assign n_15239 =  x_1879 & ~n_1770;
assign n_15240 =  n_1770 &  n_15233;
assign n_15241 = ~n_15239 & ~n_15240;
assign n_15242 =  x_1879 & ~n_15241;
assign n_15243 = ~x_1879 &  n_15241;
assign n_15244 = ~n_15242 & ~n_15243;
assign n_15245 =  x_1878 & ~n_1778;
assign n_15246 =  n_1778 &  n_15233;
assign n_15247 = ~n_15245 & ~n_15246;
assign n_15248 =  x_1878 & ~n_15247;
assign n_15249 = ~x_1878 &  n_15247;
assign n_15250 = ~n_15248 & ~n_15249;
assign n_15251 =  x_1877 & ~n_1785;
assign n_15252 =  n_1785 &  n_15233;
assign n_15253 = ~n_15251 & ~n_15252;
assign n_15254 =  x_1877 & ~n_15253;
assign n_15255 = ~x_1877 &  n_15253;
assign n_15256 = ~n_15254 & ~n_15255;
assign n_15257 =  x_1876 & ~n_1792;
assign n_15258 =  n_1792 &  n_15233;
assign n_15259 = ~n_15257 & ~n_15258;
assign n_15260 =  x_1876 & ~n_15259;
assign n_15261 = ~x_1876 &  n_15259;
assign n_15262 = ~n_15260 & ~n_15261;
assign n_15263 =  x_1875 & ~n_1799;
assign n_15264 =  n_1799 &  n_15233;
assign n_15265 = ~n_15263 & ~n_15264;
assign n_15266 =  x_1875 & ~n_15265;
assign n_15267 = ~x_1875 &  n_15265;
assign n_15268 = ~n_15266 & ~n_15267;
assign n_15269 =  x_1874 & ~n_1806;
assign n_15270 =  n_1806 &  n_15233;
assign n_15271 = ~n_15269 & ~n_15270;
assign n_15272 =  x_1874 & ~n_15271;
assign n_15273 = ~x_1874 &  n_15271;
assign n_15274 = ~n_15272 & ~n_15273;
assign n_15275 =  n_1750 & ~n_15233;
assign n_15276 = ~x_1873 & ~n_1750;
assign n_15277 = ~n_15275 & ~n_15276;
assign n_15278 =  x_1873 &  n_15277;
assign n_15279 = ~x_1873 & ~n_15277;
assign n_15280 = ~n_15278 & ~n_15279;
assign n_15281 =  x_1872 &  n_3308;
assign n_15282 = ~x_444 &  n_3307;
assign n_15283 = ~n_15281 & ~n_15282;
assign n_15284 =  x_1872 & ~n_15283;
assign n_15285 = ~x_1872 &  n_15283;
assign n_15286 = ~n_15284 & ~n_15285;
assign n_15287 =  x_1871 & ~n_1761;
assign n_15288 =  i_155 &  n_1751;
assign n_15289 =  n_1761 &  n_15288;
assign n_15290 = ~n_15287 & ~n_15289;
assign n_15291 =  x_1871 & ~n_15290;
assign n_15292 = ~x_1871 &  n_15290;
assign n_15293 = ~n_15291 & ~n_15292;
assign n_15294 =  x_1870 & ~n_1770;
assign n_15295 =  n_1770 &  n_15288;
assign n_15296 = ~n_15294 & ~n_15295;
assign n_15297 =  x_1870 & ~n_15296;
assign n_15298 = ~x_1870 &  n_15296;
assign n_15299 = ~n_15297 & ~n_15298;
assign n_15300 =  x_1869 & ~n_1778;
assign n_15301 =  n_1778 &  n_15288;
assign n_15302 = ~n_15300 & ~n_15301;
assign n_15303 =  x_1869 & ~n_15302;
assign n_15304 = ~x_1869 &  n_15302;
assign n_15305 = ~n_15303 & ~n_15304;
assign n_15306 =  x_1868 & ~n_1785;
assign n_15307 =  n_1785 &  n_15288;
assign n_15308 = ~n_15306 & ~n_15307;
assign n_15309 =  x_1868 & ~n_15308;
assign n_15310 = ~x_1868 &  n_15308;
assign n_15311 = ~n_15309 & ~n_15310;
assign n_15312 =  x_1867 & ~n_1792;
assign n_15313 =  n_1792 &  n_15288;
assign n_15314 = ~n_15312 & ~n_15313;
assign n_15315 =  x_1867 & ~n_15314;
assign n_15316 = ~x_1867 &  n_15314;
assign n_15317 = ~n_15315 & ~n_15316;
assign n_15318 =  x_1866 & ~n_1799;
assign n_15319 =  n_1799 &  n_15288;
assign n_15320 = ~n_15318 & ~n_15319;
assign n_15321 =  x_1866 & ~n_15320;
assign n_15322 = ~x_1866 &  n_15320;
assign n_15323 = ~n_15321 & ~n_15322;
assign n_15324 =  x_1865 & ~n_1806;
assign n_15325 =  n_1806 &  n_15288;
assign n_15326 = ~n_15324 & ~n_15325;
assign n_15327 =  x_1865 & ~n_15326;
assign n_15328 = ~x_1865 &  n_15326;
assign n_15329 = ~n_15327 & ~n_15328;
assign n_15330 =  n_1750 & ~n_15288;
assign n_15331 = ~x_1864 & ~n_1750;
assign n_15332 = ~n_15330 & ~n_15331;
assign n_15333 =  x_1864 &  n_15332;
assign n_15334 = ~x_1864 & ~n_15332;
assign n_15335 = ~n_15333 & ~n_15334;
assign n_15336 =  x_1863 &  n_3308;
assign n_15337 =  x_447 &  n_3307;
assign n_15338 = ~n_15336 & ~n_15337;
assign n_15339 =  x_1863 & ~n_15338;
assign n_15340 = ~x_1863 &  n_15338;
assign n_15341 = ~n_15339 & ~n_15340;
assign n_15342 =  x_1862 &  n_3308;
assign n_15343 = ~x_443 &  n_3307;
assign n_15344 = ~n_15342 & ~n_15343;
assign n_15345 =  x_1862 & ~n_15344;
assign n_15346 = ~x_1862 &  n_15344;
assign n_15347 = ~n_15345 & ~n_15346;
assign n_15348 =  x_1861 & ~n_1761;
assign n_15349 =  i_154 &  n_1751;
assign n_15350 =  n_1761 &  n_15349;
assign n_15351 = ~n_15348 & ~n_15350;
assign n_15352 =  x_1861 & ~n_15351;
assign n_15353 = ~x_1861 &  n_15351;
assign n_15354 = ~n_15352 & ~n_15353;
assign n_15355 =  x_1860 & ~n_1770;
assign n_15356 =  n_1770 &  n_15349;
assign n_15357 = ~n_15355 & ~n_15356;
assign n_15358 =  x_1860 & ~n_15357;
assign n_15359 = ~x_1860 &  n_15357;
assign n_15360 = ~n_15358 & ~n_15359;
assign n_15361 =  x_1859 & ~n_1778;
assign n_15362 =  n_1778 &  n_15349;
assign n_15363 = ~n_15361 & ~n_15362;
assign n_15364 =  x_1859 & ~n_15363;
assign n_15365 = ~x_1859 &  n_15363;
assign n_15366 = ~n_15364 & ~n_15365;
assign n_15367 =  x_1858 & ~n_1785;
assign n_15368 =  n_1785 &  n_15349;
assign n_15369 = ~n_15367 & ~n_15368;
assign n_15370 =  x_1858 & ~n_15369;
assign n_15371 = ~x_1858 &  n_15369;
assign n_15372 = ~n_15370 & ~n_15371;
assign n_15373 =  x_1857 & ~n_1792;
assign n_15374 =  n_1792 &  n_15349;
assign n_15375 = ~n_15373 & ~n_15374;
assign n_15376 =  x_1857 & ~n_15375;
assign n_15377 = ~x_1857 &  n_15375;
assign n_15378 = ~n_15376 & ~n_15377;
assign n_15379 =  x_1856 & ~n_1799;
assign n_15380 =  n_1799 &  n_15349;
assign n_15381 = ~n_15379 & ~n_15380;
assign n_15382 =  x_1856 & ~n_15381;
assign n_15383 = ~x_1856 &  n_15381;
assign n_15384 = ~n_15382 & ~n_15383;
assign n_15385 =  x_1855 & ~n_1806;
assign n_15386 =  n_1806 &  n_15349;
assign n_15387 = ~n_15385 & ~n_15386;
assign n_15388 =  x_1855 & ~n_15387;
assign n_15389 = ~x_1855 &  n_15387;
assign n_15390 = ~n_15388 & ~n_15389;
assign n_15391 =  n_1750 & ~n_15349;
assign n_15392 = ~x_1854 & ~n_1750;
assign n_15393 = ~n_15391 & ~n_15392;
assign n_15394 =  x_1854 &  n_15393;
assign n_15395 = ~x_1854 & ~n_15393;
assign n_15396 = ~n_15394 & ~n_15395;
assign n_15397 =  x_1853 & ~n_1761;
assign n_15398 =  i_153 &  n_1751;
assign n_15399 =  n_1761 &  n_15398;
assign n_15400 = ~n_15397 & ~n_15399;
assign n_15401 =  x_1853 & ~n_15400;
assign n_15402 = ~x_1853 &  n_15400;
assign n_15403 = ~n_15401 & ~n_15402;
assign n_15404 =  x_1852 & ~n_1770;
assign n_15405 =  n_1770 &  n_15398;
assign n_15406 = ~n_15404 & ~n_15405;
assign n_15407 =  x_1852 & ~n_15406;
assign n_15408 = ~x_1852 &  n_15406;
assign n_15409 = ~n_15407 & ~n_15408;
assign n_15410 =  x_1851 & ~n_1778;
assign n_15411 =  n_1778 &  n_15398;
assign n_15412 = ~n_15410 & ~n_15411;
assign n_15413 =  x_1851 & ~n_15412;
assign n_15414 = ~x_1851 &  n_15412;
assign n_15415 = ~n_15413 & ~n_15414;
assign n_15416 =  x_1850 & ~n_1785;
assign n_15417 =  n_1785 &  n_15398;
assign n_15418 = ~n_15416 & ~n_15417;
assign n_15419 =  x_1850 & ~n_15418;
assign n_15420 = ~x_1850 &  n_15418;
assign n_15421 = ~n_15419 & ~n_15420;
assign n_15422 =  x_1849 & ~n_1792;
assign n_15423 =  n_1792 &  n_15398;
assign n_15424 = ~n_15422 & ~n_15423;
assign n_15425 =  x_1849 & ~n_15424;
assign n_15426 = ~x_1849 &  n_15424;
assign n_15427 = ~n_15425 & ~n_15426;
assign n_15428 =  x_1848 & ~n_1799;
assign n_15429 =  n_1799 &  n_15398;
assign n_15430 = ~n_15428 & ~n_15429;
assign n_15431 =  x_1848 & ~n_15430;
assign n_15432 = ~x_1848 &  n_15430;
assign n_15433 = ~n_15431 & ~n_15432;
assign n_15434 =  x_1847 & ~n_1806;
assign n_15435 =  n_1806 &  n_15398;
assign n_15436 = ~n_15434 & ~n_15435;
assign n_15437 =  x_1847 & ~n_15436;
assign n_15438 = ~x_1847 &  n_15436;
assign n_15439 = ~n_15437 & ~n_15438;
assign n_15440 =  n_1750 & ~n_15398;
assign n_15441 = ~x_1846 & ~n_1750;
assign n_15442 = ~n_15440 & ~n_15441;
assign n_15443 =  x_1846 &  n_15442;
assign n_15444 = ~x_1846 & ~n_15442;
assign n_15445 = ~n_15443 & ~n_15444;
assign n_15446 =  x_1845 & ~n_1739;
assign n_15447 =  i_142 &  n_1739;
assign n_15448 = ~n_15446 & ~n_15447;
assign n_15449 =  x_1845 & ~n_15448;
assign n_15450 = ~x_1845 &  n_15448;
assign n_15451 = ~n_15449 & ~n_15450;
assign n_15452 =  x_1844 & ~n_1739;
assign n_15453 =  i_140 &  n_1739;
assign n_15454 = ~n_15452 & ~n_15453;
assign n_15455 =  x_1844 & ~n_15454;
assign n_15456 = ~x_1844 &  n_15454;
assign n_15457 = ~n_15455 & ~n_15456;
assign n_15458 =  x_1843 & ~n_1739;
assign n_15459 =  i_138 &  n_1739;
assign n_15460 = ~n_15458 & ~n_15459;
assign n_15461 =  x_1843 & ~n_15460;
assign n_15462 = ~x_1843 &  n_15460;
assign n_15463 = ~n_15461 & ~n_15462;
assign n_15464 =  x_1842 & ~n_1739;
assign n_15465 =  i_136 &  n_1739;
assign n_15466 = ~n_15464 & ~n_15465;
assign n_15467 =  x_1842 & ~n_15466;
assign n_15468 = ~x_1842 &  n_15466;
assign n_15469 = ~n_15467 & ~n_15468;
assign n_15470 =  x_1841 & ~n_1739;
assign n_15471 =  i_134 &  n_1739;
assign n_15472 = ~n_15470 & ~n_15471;
assign n_15473 =  x_1841 & ~n_15472;
assign n_15474 = ~x_1841 &  n_15472;
assign n_15475 = ~n_15473 & ~n_15474;
assign n_15476 =  x_1840 & ~n_1739;
assign n_15477 =  i_132 &  n_1739;
assign n_15478 = ~n_15476 & ~n_15477;
assign n_15479 =  x_1840 & ~n_15478;
assign n_15480 = ~x_1840 &  n_15478;
assign n_15481 = ~n_15479 & ~n_15480;
assign n_15482 =  x_1839 & ~n_1739;
assign n_15483 =  i_130 &  n_1739;
assign n_15484 = ~n_15482 & ~n_15483;
assign n_15485 =  x_1839 & ~n_15484;
assign n_15486 = ~x_1839 &  n_15484;
assign n_15487 = ~n_15485 & ~n_15486;
assign n_15488 =  x_1838 & ~n_1739;
assign n_15489 =  i_128 &  n_1739;
assign n_15490 = ~n_15488 & ~n_15489;
assign n_15491 =  x_1838 & ~n_15490;
assign n_15492 = ~x_1838 &  n_15490;
assign n_15493 = ~n_15491 & ~n_15492;
assign n_15494 =  x_1837 & ~n_1739;
assign n_15495 =  i_126 &  n_1739;
assign n_15496 = ~n_15494 & ~n_15495;
assign n_15497 =  x_1837 & ~n_15496;
assign n_15498 = ~x_1837 &  n_15496;
assign n_15499 = ~n_15497 & ~n_15498;
assign n_15500 =  x_1836 & ~n_1739;
assign n_15501 =  i_124 &  n_1739;
assign n_15502 = ~n_15500 & ~n_15501;
assign n_15503 =  x_1836 & ~n_15502;
assign n_15504 = ~x_1836 &  n_15502;
assign n_15505 = ~n_15503 & ~n_15504;
assign n_15506 =  x_1835 & ~n_1739;
assign n_15507 =  i_122 &  n_1739;
assign n_15508 = ~n_15506 & ~n_15507;
assign n_15509 =  x_1835 & ~n_15508;
assign n_15510 = ~x_1835 &  n_15508;
assign n_15511 = ~n_15509 & ~n_15510;
assign n_15512 =  x_1834 & ~n_1739;
assign n_15513 =  i_120 &  n_1739;
assign n_15514 = ~n_15512 & ~n_15513;
assign n_15515 =  x_1834 & ~n_15514;
assign n_15516 = ~x_1834 &  n_15514;
assign n_15517 = ~n_15515 & ~n_15516;
assign n_15518 =  x_1833 & ~n_1739;
assign n_15519 =  i_118 &  n_1739;
assign n_15520 = ~n_15518 & ~n_15519;
assign n_15521 =  x_1833 & ~n_15520;
assign n_15522 = ~x_1833 &  n_15520;
assign n_15523 = ~n_15521 & ~n_15522;
assign n_15524 =  x_1832 & ~n_1739;
assign n_15525 =  i_116 &  n_1739;
assign n_15526 = ~n_15524 & ~n_15525;
assign n_15527 =  x_1832 & ~n_15526;
assign n_15528 = ~x_1832 &  n_15526;
assign n_15529 = ~n_15527 & ~n_15528;
assign n_15530 =  x_1831 & ~n_1739;
assign n_15531 =  i_114 &  n_1739;
assign n_15532 = ~n_15530 & ~n_15531;
assign n_15533 =  x_1831 & ~n_15532;
assign n_15534 = ~x_1831 &  n_15532;
assign n_15535 = ~n_15533 & ~n_15534;
assign n_15536 =  x_1830 & ~n_1739;
assign n_15537 =  i_112 &  n_1739;
assign n_15538 = ~n_15536 & ~n_15537;
assign n_15539 =  x_1830 & ~n_15538;
assign n_15540 = ~x_1830 &  n_15538;
assign n_15541 = ~n_15539 & ~n_15540;
assign n_15542 =  x_1829 & ~n_1739;
assign n_15543 =  i_110 &  n_1739;
assign n_15544 = ~n_15542 & ~n_15543;
assign n_15545 =  x_1829 & ~n_15544;
assign n_15546 = ~x_1829 &  n_15544;
assign n_15547 = ~n_15545 & ~n_15546;
assign n_15548 =  x_1828 & ~n_1739;
assign n_15549 =  i_108 &  n_1739;
assign n_15550 = ~n_15548 & ~n_15549;
assign n_15551 =  x_1828 & ~n_15550;
assign n_15552 = ~x_1828 &  n_15550;
assign n_15553 = ~n_15551 & ~n_15552;
assign n_15554 =  x_1827 & ~n_1739;
assign n_15555 =  i_106 &  n_1739;
assign n_15556 = ~n_15554 & ~n_15555;
assign n_15557 =  x_1827 & ~n_15556;
assign n_15558 = ~x_1827 &  n_15556;
assign n_15559 = ~n_15557 & ~n_15558;
assign n_15560 =  x_1826 & ~n_1739;
assign n_15561 =  i_104 &  n_1739;
assign n_15562 = ~n_15560 & ~n_15561;
assign n_15563 =  x_1826 & ~n_15562;
assign n_15564 = ~x_1826 &  n_15562;
assign n_15565 = ~n_15563 & ~n_15564;
assign n_15566 =  x_1825 & ~n_1739;
assign n_15567 =  i_102 &  n_1739;
assign n_15568 = ~n_15566 & ~n_15567;
assign n_15569 =  x_1825 & ~n_15568;
assign n_15570 = ~x_1825 &  n_15568;
assign n_15571 = ~n_15569 & ~n_15570;
assign n_15572 =  x_1824 & ~n_1739;
assign n_15573 =  i_100 &  n_1739;
assign n_15574 = ~n_15572 & ~n_15573;
assign n_15575 =  x_1824 & ~n_15574;
assign n_15576 = ~x_1824 &  n_15574;
assign n_15577 = ~n_15575 & ~n_15576;
assign n_15578 =  x_1823 & ~n_1739;
assign n_15579 =  i_98 &  n_1739;
assign n_15580 = ~n_15578 & ~n_15579;
assign n_15581 =  x_1823 & ~n_15580;
assign n_15582 = ~x_1823 &  n_15580;
assign n_15583 = ~n_15581 & ~n_15582;
assign n_15584 =  x_1822 & ~n_1739;
assign n_15585 =  i_96 &  n_1739;
assign n_15586 = ~n_15584 & ~n_15585;
assign n_15587 =  x_1822 & ~n_15586;
assign n_15588 = ~x_1822 &  n_15586;
assign n_15589 = ~n_15587 & ~n_15588;
assign n_15590 =  x_1821 & ~n_1739;
assign n_15591 =  i_94 &  n_1739;
assign n_15592 = ~n_15590 & ~n_15591;
assign n_15593 =  x_1821 & ~n_15592;
assign n_15594 = ~x_1821 &  n_15592;
assign n_15595 = ~n_15593 & ~n_15594;
assign n_15596 =  x_1820 & ~n_1739;
assign n_15597 =  i_92 &  n_1739;
assign n_15598 = ~n_15596 & ~n_15597;
assign n_15599 =  x_1820 & ~n_15598;
assign n_15600 = ~x_1820 &  n_15598;
assign n_15601 = ~n_15599 & ~n_15600;
assign n_15602 =  x_1819 & ~n_1739;
assign n_15603 =  i_90 &  n_1739;
assign n_15604 = ~n_15602 & ~n_15603;
assign n_15605 =  x_1819 & ~n_15604;
assign n_15606 = ~x_1819 &  n_15604;
assign n_15607 = ~n_15605 & ~n_15606;
assign n_15608 =  x_1818 & ~n_1739;
assign n_15609 =  i_88 &  n_1739;
assign n_15610 = ~n_15608 & ~n_15609;
assign n_15611 =  x_1818 & ~n_15610;
assign n_15612 = ~x_1818 &  n_15610;
assign n_15613 = ~n_15611 & ~n_15612;
assign n_15614 =  x_1817 & ~n_1739;
assign n_15615 =  i_86 &  n_1739;
assign n_15616 = ~n_15614 & ~n_15615;
assign n_15617 =  x_1817 & ~n_15616;
assign n_15618 = ~x_1817 &  n_15616;
assign n_15619 = ~n_15617 & ~n_15618;
assign n_15620 =  x_1816 & ~n_1739;
assign n_15621 =  i_84 &  n_1739;
assign n_15622 = ~n_15620 & ~n_15621;
assign n_15623 =  x_1816 & ~n_15622;
assign n_15624 = ~x_1816 &  n_15622;
assign n_15625 = ~n_15623 & ~n_15624;
assign n_15626 =  x_1815 & ~n_1739;
assign n_15627 =  i_82 &  n_1739;
assign n_15628 = ~n_15626 & ~n_15627;
assign n_15629 =  x_1815 & ~n_15628;
assign n_15630 = ~x_1815 &  n_15628;
assign n_15631 = ~n_15629 & ~n_15630;
assign n_15632 =  x_1814 & ~n_1739;
assign n_15633 =  i_80 &  n_1739;
assign n_15634 = ~n_15632 & ~n_15633;
assign n_15635 =  x_1814 & ~n_15634;
assign n_15636 = ~x_1814 &  n_15634;
assign n_15637 = ~n_15635 & ~n_15636;
assign n_15638 =  x_1813 & ~n_1739;
assign n_15639 = ~n_6126 & ~n_15638;
assign n_15640 =  x_1813 & ~n_15639;
assign n_15641 = ~x_1813 &  n_15639;
assign n_15642 = ~n_15640 & ~n_15641;
assign n_15643 =  x_1812 & ~n_1739;
assign n_15644 =  i_78 &  n_1739;
assign n_15645 = ~n_15643 & ~n_15644;
assign n_15646 =  x_1812 & ~n_15645;
assign n_15647 = ~x_1812 &  n_15645;
assign n_15648 = ~n_15646 & ~n_15647;
assign n_15649 =  x_1811 & ~n_1739;
assign n_15650 =  i_76 &  n_1739;
assign n_15651 = ~n_15649 & ~n_15650;
assign n_15652 =  x_1811 & ~n_15651;
assign n_15653 = ~x_1811 &  n_15651;
assign n_15654 = ~n_15652 & ~n_15653;
assign n_15655 =  x_1810 & ~n_1739;
assign n_15656 =  i_74 &  n_1739;
assign n_15657 = ~n_15655 & ~n_15656;
assign n_15658 =  x_1810 & ~n_15657;
assign n_15659 = ~x_1810 &  n_15657;
assign n_15660 = ~n_15658 & ~n_15659;
assign n_15661 =  x_1809 & ~n_1739;
assign n_15662 =  i_72 &  n_1739;
assign n_15663 = ~n_15661 & ~n_15662;
assign n_15664 =  x_1809 & ~n_15663;
assign n_15665 = ~x_1809 &  n_15663;
assign n_15666 = ~n_15664 & ~n_15665;
assign n_15667 =  x_1808 & ~n_1739;
assign n_15668 =  i_70 &  n_1739;
assign n_15669 = ~n_15667 & ~n_15668;
assign n_15670 =  x_1808 & ~n_15669;
assign n_15671 = ~x_1808 &  n_15669;
assign n_15672 = ~n_15670 & ~n_15671;
assign n_15673 =  x_1807 & ~n_1739;
assign n_15674 =  i_68 &  n_1739;
assign n_15675 = ~n_15673 & ~n_15674;
assign n_15676 =  x_1807 & ~n_15675;
assign n_15677 = ~x_1807 &  n_15675;
assign n_15678 = ~n_15676 & ~n_15677;
assign n_15679 =  x_1806 & ~n_1739;
assign n_15680 =  i_66 &  n_1739;
assign n_15681 = ~n_15679 & ~n_15680;
assign n_15682 =  x_1806 & ~n_15681;
assign n_15683 = ~x_1806 &  n_15681;
assign n_15684 = ~n_15682 & ~n_15683;
assign n_15685 =  x_1805 & ~n_1739;
assign n_15686 =  i_64 &  n_1739;
assign n_15687 = ~n_15685 & ~n_15686;
assign n_15688 =  x_1805 & ~n_15687;
assign n_15689 = ~x_1805 &  n_15687;
assign n_15690 = ~n_15688 & ~n_15689;
assign n_15691 =  x_1804 & ~n_1739;
assign n_15692 =  i_62 &  n_1739;
assign n_15693 = ~n_15691 & ~n_15692;
assign n_15694 =  x_1804 & ~n_15693;
assign n_15695 = ~x_1804 &  n_15693;
assign n_15696 = ~n_15694 & ~n_15695;
assign n_15697 =  x_1803 & ~n_1739;
assign n_15698 =  i_60 &  n_1739;
assign n_15699 = ~n_15697 & ~n_15698;
assign n_15700 =  x_1803 & ~n_15699;
assign n_15701 = ~x_1803 &  n_15699;
assign n_15702 = ~n_15700 & ~n_15701;
assign n_15703 =  x_1802 & ~n_1739;
assign n_15704 =  i_58 &  n_1739;
assign n_15705 = ~n_15703 & ~n_15704;
assign n_15706 =  x_1802 & ~n_15705;
assign n_15707 = ~x_1802 &  n_15705;
assign n_15708 = ~n_15706 & ~n_15707;
assign n_15709 =  x_1801 & ~n_1739;
assign n_15710 =  i_56 &  n_1739;
assign n_15711 = ~n_15709 & ~n_15710;
assign n_15712 =  x_1801 & ~n_15711;
assign n_15713 = ~x_1801 &  n_15711;
assign n_15714 = ~n_15712 & ~n_15713;
assign n_15715 =  x_1800 & ~n_1739;
assign n_15716 =  i_54 &  n_1739;
assign n_15717 = ~n_15715 & ~n_15716;
assign n_15718 =  x_1800 & ~n_15717;
assign n_15719 = ~x_1800 &  n_15717;
assign n_15720 = ~n_15718 & ~n_15719;
assign n_15721 =  x_1799 & ~n_1739;
assign n_15722 =  i_52 &  n_1739;
assign n_15723 = ~n_15721 & ~n_15722;
assign n_15724 =  x_1799 & ~n_15723;
assign n_15725 = ~x_1799 &  n_15723;
assign n_15726 = ~n_15724 & ~n_15725;
assign n_15727 =  x_1798 & ~n_1739;
assign n_15728 =  i_50 &  n_1739;
assign n_15729 = ~n_15727 & ~n_15728;
assign n_15730 =  x_1798 & ~n_15729;
assign n_15731 = ~x_1798 &  n_15729;
assign n_15732 = ~n_15730 & ~n_15731;
assign n_15733 =  x_1797 & ~n_1739;
assign n_15734 =  i_48 &  n_1739;
assign n_15735 = ~n_15733 & ~n_15734;
assign n_15736 =  x_1797 & ~n_15735;
assign n_15737 = ~x_1797 &  n_15735;
assign n_15738 = ~n_15736 & ~n_15737;
assign n_15739 =  x_1796 & ~n_1739;
assign n_15740 =  i_46 &  n_1739;
assign n_15741 = ~n_15739 & ~n_15740;
assign n_15742 =  x_1796 & ~n_15741;
assign n_15743 = ~x_1796 &  n_15741;
assign n_15744 = ~n_15742 & ~n_15743;
assign n_15745 =  x_1795 & ~n_1739;
assign n_15746 =  i_44 &  n_1739;
assign n_15747 = ~n_15745 & ~n_15746;
assign n_15748 =  x_1795 & ~n_15747;
assign n_15749 = ~x_1795 &  n_15747;
assign n_15750 = ~n_15748 & ~n_15749;
assign n_15751 =  x_1794 & ~n_1739;
assign n_15752 =  i_42 &  n_1739;
assign n_15753 = ~n_15751 & ~n_15752;
assign n_15754 =  x_1794 & ~n_15753;
assign n_15755 = ~x_1794 &  n_15753;
assign n_15756 = ~n_15754 & ~n_15755;
assign n_15757 =  x_1793 & ~n_1739;
assign n_15758 =  i_40 &  n_1739;
assign n_15759 = ~n_15757 & ~n_15758;
assign n_15760 =  x_1793 & ~n_15759;
assign n_15761 = ~x_1793 &  n_15759;
assign n_15762 = ~n_15760 & ~n_15761;
assign n_15763 =  x_1792 & ~n_1739;
assign n_15764 =  i_38 &  n_1739;
assign n_15765 = ~n_15763 & ~n_15764;
assign n_15766 =  x_1792 & ~n_15765;
assign n_15767 = ~x_1792 &  n_15765;
assign n_15768 = ~n_15766 & ~n_15767;
assign n_15769 =  x_1791 & ~n_1739;
assign n_15770 =  i_36 &  n_1739;
assign n_15771 = ~n_15769 & ~n_15770;
assign n_15772 =  x_1791 & ~n_15771;
assign n_15773 = ~x_1791 &  n_15771;
assign n_15774 = ~n_15772 & ~n_15773;
assign n_15775 =  x_1790 & ~n_1739;
assign n_15776 =  i_34 &  n_1739;
assign n_15777 = ~n_15775 & ~n_15776;
assign n_15778 =  x_1790 & ~n_15777;
assign n_15779 = ~x_1790 &  n_15777;
assign n_15780 = ~n_15778 & ~n_15779;
assign n_15781 =  x_1789 & ~n_1739;
assign n_15782 =  i_32 &  n_1739;
assign n_15783 = ~n_15781 & ~n_15782;
assign n_15784 =  x_1789 & ~n_15783;
assign n_15785 = ~x_1789 &  n_15783;
assign n_15786 = ~n_15784 & ~n_15785;
assign n_15787 =  x_1788 & ~n_1739;
assign n_15788 =  i_30 &  n_1739;
assign n_15789 = ~n_15787 & ~n_15788;
assign n_15790 =  x_1788 & ~n_15789;
assign n_15791 = ~x_1788 &  n_15789;
assign n_15792 = ~n_15790 & ~n_15791;
assign n_15793 =  x_1787 & ~n_1739;
assign n_15794 =  i_28 &  n_1739;
assign n_15795 = ~n_15793 & ~n_15794;
assign n_15796 =  x_1787 & ~n_15795;
assign n_15797 = ~x_1787 &  n_15795;
assign n_15798 = ~n_15796 & ~n_15797;
assign n_15799 =  x_1786 & ~n_1739;
assign n_15800 =  i_26 &  n_1739;
assign n_15801 = ~n_15799 & ~n_15800;
assign n_15802 =  x_1786 & ~n_15801;
assign n_15803 = ~x_1786 &  n_15801;
assign n_15804 = ~n_15802 & ~n_15803;
assign n_15805 =  x_1785 & ~n_1739;
assign n_15806 =  i_24 &  n_1739;
assign n_15807 = ~n_15805 & ~n_15806;
assign n_15808 =  x_1785 & ~n_15807;
assign n_15809 = ~x_1785 &  n_15807;
assign n_15810 = ~n_15808 & ~n_15809;
assign n_15811 =  x_1784 & ~n_1739;
assign n_15812 =  i_22 &  n_1739;
assign n_15813 = ~n_15811 & ~n_15812;
assign n_15814 =  x_1784 & ~n_15813;
assign n_15815 = ~x_1784 &  n_15813;
assign n_15816 = ~n_15814 & ~n_15815;
assign n_15817 =  x_1783 & ~n_1739;
assign n_15818 =  i_20 &  n_1739;
assign n_15819 = ~n_15817 & ~n_15818;
assign n_15820 =  x_1783 & ~n_15819;
assign n_15821 = ~x_1783 &  n_15819;
assign n_15822 = ~n_15820 & ~n_15821;
assign n_15823 =  x_1782 & ~n_1739;
assign n_15824 =  i_18 &  n_1739;
assign n_15825 = ~n_15823 & ~n_15824;
assign n_15826 =  x_1782 & ~n_15825;
assign n_15827 = ~x_1782 &  n_15825;
assign n_15828 = ~n_15826 & ~n_15827;
assign n_15829 =  x_1781 & ~n_1739;
assign n_15830 =  i_16 &  n_1739;
assign n_15831 = ~n_15829 & ~n_15830;
assign n_15832 =  x_1781 & ~n_15831;
assign n_15833 = ~x_1781 &  n_15831;
assign n_15834 = ~n_15832 & ~n_15833;
assign n_15835 =  x_1780 & ~n_1739;
assign n_15836 =  i_15 &  n_1739;
assign n_15837 = ~n_15835 & ~n_15836;
assign n_15838 =  x_1780 & ~n_15837;
assign n_15839 = ~x_1780 &  n_15837;
assign n_15840 = ~n_15838 & ~n_15839;
assign n_15841 =  x_1779 & ~n_1739;
assign n_15842 =  i_150 &  n_1739;
assign n_15843 = ~n_15841 & ~n_15842;
assign n_15844 =  x_1779 & ~n_15843;
assign n_15845 = ~x_1779 &  n_15843;
assign n_15846 = ~n_15844 & ~n_15845;
assign n_15847 =  x_1778 & ~n_1739;
assign n_15848 =  i_149 &  n_1739;
assign n_15849 = ~n_15847 & ~n_15848;
assign n_15850 =  x_1778 & ~n_15849;
assign n_15851 = ~x_1778 &  n_15849;
assign n_15852 = ~n_15850 & ~n_15851;
assign n_15853 =  x_1777 & ~n_1739;
assign n_15854 =  i_148 &  n_1739;
assign n_15855 = ~n_15853 & ~n_15854;
assign n_15856 =  x_1777 & ~n_15855;
assign n_15857 = ~x_1777 &  n_15855;
assign n_15858 = ~n_15856 & ~n_15857;
assign n_15859 =  x_1776 & ~n_1739;
assign n_15860 =  i_147 &  n_1739;
assign n_15861 = ~n_15859 & ~n_15860;
assign n_15862 =  x_1776 & ~n_15861;
assign n_15863 = ~x_1776 &  n_15861;
assign n_15864 = ~n_15862 & ~n_15863;
assign n_15865 =  x_1775 & ~n_1739;
assign n_15866 =  i_146 &  n_1739;
assign n_15867 = ~n_15865 & ~n_15866;
assign n_15868 =  x_1775 & ~n_15867;
assign n_15869 = ~x_1775 &  n_15867;
assign n_15870 = ~n_15868 & ~n_15869;
assign n_15871 =  x_1774 & ~n_1739;
assign n_15872 =  i_145 &  n_1739;
assign n_15873 = ~n_15871 & ~n_15872;
assign n_15874 =  x_1774 & ~n_15873;
assign n_15875 = ~x_1774 &  n_15873;
assign n_15876 = ~n_15874 & ~n_15875;
assign n_15877 =  x_1773 & ~n_1739;
assign n_15878 =  i_144 &  n_1739;
assign n_15879 = ~n_15877 & ~n_15878;
assign n_15880 =  x_1773 & ~n_15879;
assign n_15881 = ~x_1773 &  n_15879;
assign n_15882 = ~n_15880 & ~n_15881;
assign n_15883 =  x_1772 & ~n_1739;
assign n_15884 =  i_143 &  n_1739;
assign n_15885 = ~n_15883 & ~n_15884;
assign n_15886 =  x_1772 & ~n_15885;
assign n_15887 = ~x_1772 &  n_15885;
assign n_15888 = ~n_15886 & ~n_15887;
assign n_15889 = ~n_3263 &  n_3281;
assign n_15890 = ~x_1771 & ~n_15889;
assign n_15891 =  n_3294 & ~n_15890;
assign n_15892 = ~n_3246 &  n_3245;
assign n_15893 =  x_1761 &  n_3257;
assign n_15894 =  n_3253 &  n_15893;
assign n_15895 = ~n_15892 & ~n_15894;
assign n_15896 =  x_1768 & ~n_3294;
assign n_15897 = ~n_15895 &  n_15896;
assign n_15898 = ~n_15891 & ~n_15897;
assign n_15899 =  x_1771 & ~n_15898;
assign n_15900 = ~x_1771 &  n_15898;
assign n_15901 = ~n_15899 & ~n_15900;
assign n_15902 =  x_1759 &  n_12533;
assign n_15903 = ~n_12554 &  n_15902;
assign n_15904 = ~x_1770 & ~n_15902;
assign n_15905 = ~n_12581 &  n_15904;
assign n_15906 = ~n_15903 & ~n_15905;
assign n_15907 =  x_1770 &  n_15906;
assign n_15908 = ~x_1770 & ~n_15906;
assign n_15909 = ~n_15907 & ~n_15908;
assign n_15910 =  x_1763 &  n_3308;
assign n_15911 =  x_435 & ~n_15910;
assign n_15912 =  n_12532 &  n_12584;
assign n_15913 = ~n_12549 &  n_12577;
assign n_15914 =  x_1762 & ~n_15913;
assign n_15915 = ~n_15912 &  n_15914;
assign n_15916 = ~x_1489 & ~x_1765;
assign n_15917 =  n_1751 & ~n_15916;
assign n_15918 = ~n_3263 &  n_15917;
assign n_15919 =  n_12583 &  n_15918;
assign n_15920 = ~n_15915 & ~n_15919;
assign n_15921 = ~x_442 &  n_3307;
assign n_15922 = ~n_15910 & ~n_15921;
assign n_15923 =  n_15920 & ~n_15922;
assign n_15924 = ~n_15911 &  n_15923;
assign n_15925 =  x_1769 &  n_15924;
assign n_15926 = ~x_1769 & ~n_15924;
assign n_15927 = ~n_15925 & ~n_15926;
assign n_15928 =  n_12584 & ~n_15916;
assign n_15929 = ~x_1768 & ~n_12581;
assign n_15930 = ~n_15928 &  n_15929;
assign n_15931 =  n_12551 &  n_15912;
assign n_15932 = ~n_15913 & ~n_15931;
assign n_15933 = ~n_15930 &  n_15932;
assign n_15934 =  x_1768 &  n_15933;
assign n_15935 = ~x_1768 & ~n_15933;
assign n_15936 = ~n_15934 & ~n_15935;
assign n_15937 =  n_12549 &  n_12583;
assign n_15938 =  x_1767 &  n_15937;
assign n_15939 = ~x_1767 & ~n_15937;
assign n_15940 = ~n_15938 & ~n_15939;
assign n_15941 =  n_12512 &  n_12551;
assign n_15942 =  x_1770 &  n_12589;
assign n_15943 = ~n_15941 & ~n_15942;
assign n_15944 = ~n_12537 &  n_15943;
assign n_15945 = ~n_15913 &  n_15944;
assign n_15946 =  x_1766 &  n_15945;
assign n_15947 =  x_1491 &  n_12537;
assign n_15948 = ~n_12537 & ~n_15943;
assign n_15949 = ~x_1766 &  n_15948;
assign n_15950 = ~n_15947 & ~n_15949;
assign n_15951 = ~n_15946 &  n_15950;
assign n_15952 =  x_1766 & ~n_15951;
assign n_15953 = ~x_1766 &  n_15951;
assign n_15954 = ~n_15952 & ~n_15953;
assign n_15955 =  x_1765 &  n_15945;
assign n_15956 = ~n_12531 & ~n_12592;
assign n_15957 =  n_15948 &  n_15956;
assign n_15958 = ~n_15957 & ~n_15947;
assign n_15959 = ~n_15955 &  n_15958;
assign n_15960 =  x_1765 & ~n_15959;
assign n_15961 = ~x_1765 &  n_15959;
assign n_15962 = ~n_15960 & ~n_15961;
assign n_15963 =  n_6125 & ~n_6134;
assign n_15964 = ~n_6130 & ~n_15963;
assign n_15965 = ~n_15964 & ~n_6135;
assign n_15966 =  n_6121 & ~n_15965;
assign n_15967 = ~n_6109 & ~n_15966;
assign n_15968 =  n_6121 &  n_15964;
assign n_15969 = ~x_1600 & ~x_1601;
assign n_15970 = ~x_1598 & ~x_1599;
assign n_15971 =  n_15969 &  n_15970;
assign n_15972 = ~x_1734 &  n_15971;
assign n_15973 =  n_15968 &  n_15972;
assign n_15974 = ~n_15967 & ~n_15973;
assign n_15975 =  x_1764 & ~n_6137;
assign n_15976 = ~n_15966 &  n_15975;
assign n_15977 = ~n_15974 & ~n_15976;
assign n_15978 =  x_1764 & ~n_15977;
assign n_15979 = ~x_1764 &  n_15977;
assign n_15980 = ~n_15978 & ~n_15979;
assign n_15981 =  x_1763 & ~n_15922;
assign n_15982 = ~x_1763 &  n_15922;
assign n_15983 = ~n_15981 & ~n_15982;
assign n_15984 =  x_1762 & ~n_15920;
assign n_15985 = ~x_1762 &  n_15920;
assign n_15986 = ~n_15984 & ~n_15985;
assign n_15987 =  x_1761 & ~n_12602;
assign n_15988 = ~x_1761 &  n_12602;
assign n_15989 = ~n_15987 & ~n_15988;
assign n_15990 =  x_1760 &  n_12581;
assign n_15991 = ~x_1760 & ~n_12581;
assign n_15992 = ~n_15990 & ~n_15991;
assign n_15993 =  x_1759 &  n_12580;
assign n_15994 = ~x_1759 & ~n_12580;
assign n_15995 = ~n_15993 & ~n_15994;
assign n_15996 =  x_1758 &  n_12578;
assign n_15997 = ~x_1758 & ~n_12578;
assign n_15998 = ~n_15996 & ~n_15997;
assign n_15999 =  x_1757 & ~n_12576;
assign n_16000 = ~x_1757 &  n_12576;
assign n_16001 = ~n_15999 & ~n_16000;
assign n_16002 =  x_1756 & ~n_12566;
assign n_16003 = ~x_1756 &  n_12566;
assign n_16004 = ~n_16002 & ~n_16003;
assign n_16005 =  x_1755 & ~n_12549;
assign n_16006 = ~x_1755 &  n_12549;
assign n_16007 = ~n_16005 & ~n_16006;
assign n_16008 =  x_1754 &  n_3563;
assign n_16009 = ~x_1754 & ~n_3563;
assign n_16010 = ~n_16008 & ~n_16009;
assign n_16011 =  x_1753 &  n_15910;
assign n_16012 = ~x_1753 & ~n_15910;
assign n_16013 = ~n_16011 & ~n_16012;
assign n_16014 =  x_1752 &  n_3308;
assign n_16015 = ~x_438 &  n_3307;
assign n_16016 = ~n_16014 & ~n_16015;
assign n_16017 =  x_1752 & ~n_16016;
assign n_16018 = ~x_1752 &  n_16016;
assign n_16019 = ~n_16017 & ~n_16018;
assign n_16020 = ~x_441 &  n_3286;
assign n_16021 = ~x_435 & ~x_436;
assign n_16022 = ~x_437 & ~x_439;
assign n_16023 = ~x_440 &  n_16022;
assign n_16024 =  n_16021 &  n_16023;
assign n_16025 =  n_16020 &  n_16024;
assign n_16026 =  n_3306 & ~n_16025;
assign n_16027 =  x_1751 & ~n_16026;
assign n_16028 = ~x_1751 &  n_16026;
assign n_16029 = ~n_16027 & ~n_16028;
assign n_16030 =  n_3306 & ~n_16020;
assign n_16031 =  x_1750 &  n_16030;
assign n_16032 = ~x_1750 & ~n_16030;
assign n_16033 = ~n_16031 & ~n_16032;
assign n_16034 =  x_1749 &  n_3307;
assign n_16035 = ~x_1749 & ~n_3307;
assign n_16036 = ~n_16034 & ~n_16035;
assign n_16037 =  x_1748 & ~n_3306;
assign n_16038 = ~x_1748 &  n_3306;
assign n_16039 = ~n_16037 & ~n_16038;
assign n_16040 =  x_1747 &  n_3286;
assign n_16041 = ~x_1747 & ~n_3286;
assign n_16042 = ~n_16040 & ~n_16041;
assign n_16043 =  x_1746 &  n_3305;
assign n_16044 = ~x_1746 & ~n_3305;
assign n_16045 = ~n_16043 & ~n_16044;
assign n_16046 =  x_1745 &  n_3298;
assign n_16047 = ~x_1745 & ~n_3298;
assign n_16048 = ~n_16046 & ~n_16047;
assign n_16049 =  x_1744 & ~n_1739;
assign n_16050 =  i_2 &  n_1739;
assign n_16051 = ~n_16049 & ~n_16050;
assign n_16052 =  x_1744 & ~n_16051;
assign n_16053 = ~x_1744 &  n_16051;
assign n_16054 = ~n_16052 & ~n_16053;
assign n_16055 =  x_1743 & ~n_1739;
assign n_16056 =  i_4 &  n_1739;
assign n_16057 = ~n_16055 & ~n_16056;
assign n_16058 =  x_1743 & ~n_16057;
assign n_16059 = ~x_1743 &  n_16057;
assign n_16060 = ~n_16058 & ~n_16059;
assign n_16061 =  x_1742 & ~n_1739;
assign n_16062 =  i_8 &  n_1739;
assign n_16063 = ~n_16061 & ~n_16062;
assign n_16064 =  x_1742 & ~n_16063;
assign n_16065 = ~x_1742 &  n_16063;
assign n_16066 = ~n_16064 & ~n_16065;
assign n_16067 =  x_1741 & ~n_1739;
assign n_16068 = ~i_7 &  n_1739;
assign n_16069 = ~n_16067 & ~n_16068;
assign n_16070 =  x_1741 & ~n_16069;
assign n_16071 = ~x_1741 &  n_16069;
assign n_16072 = ~n_16070 & ~n_16071;
assign n_16073 =  x_1740 & ~n_1739;
assign n_16074 =  i_6 &  n_1739;
assign n_16075 = ~n_16073 & ~n_16074;
assign n_16076 =  x_1740 & ~n_16075;
assign n_16077 = ~x_1740 &  n_16075;
assign n_16078 = ~n_16076 & ~n_16077;
assign n_16079 =  x_1739 & ~n_1739;
assign n_16080 = ~i_5 &  n_1739;
assign n_16081 = ~n_16079 & ~n_16080;
assign n_16082 =  x_1739 & ~n_16081;
assign n_16083 = ~x_1739 &  n_16081;
assign n_16084 = ~n_16082 & ~n_16083;
assign n_16085 =  x_1738 & ~n_1739;
assign n_16086 = ~n_6119 & ~n_16085;
assign n_16087 =  x_1738 & ~n_16086;
assign n_16088 = ~x_1738 &  n_16086;
assign n_16089 = ~n_16087 & ~n_16088;
assign n_16090 =  x_1737 & ~n_1739;
assign n_16091 = ~n_6122 & ~n_16090;
assign n_16092 =  x_1737 & ~n_16091;
assign n_16093 = ~x_1737 &  n_16091;
assign n_16094 = ~n_16092 & ~n_16093;
assign n_16095 = ~x_1736 &  n_6136;
assign n_16096 =  x_1736 &  n_16095;
assign n_16097 = ~x_1736 & ~n_16095;
assign n_16098 = ~n_16096 & ~n_16097;
assign n_16099 =  n_6121 &  n_15963;
assign n_16100 = ~n_15964 & ~n_16099;
assign n_16101 = ~n_15966 & ~n_16100;
assign n_16102 = ~n_6109 & ~n_16099;
assign n_16103 = ~n_16101 &  n_16102;
assign n_16104 =  x_1735 & ~n_16103;
assign n_16105 = ~x_1735 &  n_16103;
assign n_16106 = ~n_16104 & ~n_16105;
assign n_16107 =  x_1734 &  n_16101;
assign n_16108 = ~x_1734 & ~n_16101;
assign n_16109 = ~n_16107 & ~n_16108;
assign n_16110 = ~n_6111 &  n_6130;
assign n_16111 = ~n_16099 &  n_16110;
assign n_16112 =  x_1733 &  n_16111;
assign n_16113 = ~x_1733 & ~n_16111;
assign n_16114 = ~n_16112 & ~n_16113;
assign n_16115 =  x_1732 & ~n_15968;
assign n_16116 = ~x_1732 &  n_15968;
assign n_16117 = ~n_16115 & ~n_16116;
assign n_16118 =  x_1731 &  n_6005;
assign n_16119 = ~x_1731 & ~n_6005;
assign n_16120 = ~n_16118 & ~n_16119;
assign n_16121 =  x_1730 &  n_6124;
assign n_16122 = ~x_1730 & ~n_6124;
assign n_16123 = ~n_16121 & ~n_16122;
assign n_16124 =  x_1729 & ~n_3673;
assign n_16125 = ~x_1723 & ~x_1724;
assign n_16126 = ~n_3679 & ~n_16125;
assign n_16127 =  n_3678 & ~n_16126;
assign n_16128 = ~x_308 &  n_3674;
assign n_16129 = ~x_1723 &  n_16128;
assign n_16130 = ~n_16127 & ~n_16129;
assign n_16131 =  n_3683 &  n_16130;
assign n_16132 =  n_16131 & ~n_4287;
assign n_16133 =  n_16124 & ~n_16132;
assign n_16134 =  x_1723 & ~x_1724;
assign n_16135 =  n_16128 &  n_16134;
assign n_16136 = ~n_4284 & ~n_16135;
assign n_16137 =  n_3696 & ~n_16136;
assign n_16138 = ~x_1727 &  n_3673;
assign n_16139 = ~x_1729 & ~n_16138;
assign n_16140 = ~n_16137 &  n_16139;
assign n_16141 = ~n_16133 & ~n_16140;
assign n_16142 = ~x_308 & ~n_4284;
assign n_16143 =  n_3678 &  n_16134;
assign n_16144 =  n_16142 & ~n_16143;
assign n_16145 =  n_4280 & ~n_16144;
assign n_16146 =  n_16132 &  n_16145;
assign n_16147 = ~n_16141 & ~n_16146;
assign n_16148 =  x_1729 & ~n_16147;
assign n_16149 = ~x_1729 &  n_16147;
assign n_16150 = ~n_16148 & ~n_16149;
assign n_16151 = ~n_3673 &  n_16132;
assign n_16152 = ~x_308 &  n_4287;
assign n_16153 =  n_3679 & ~n_16152;
assign n_16154 =  x_308 & ~n_4287;
assign n_16155 = ~n_3676 & ~n_16154;
assign n_16156 = ~n_16153 &  n_16155;
assign n_16157 =  x_308 &  x_1722;
assign n_16158 =  n_3685 &  n_16157;
assign n_16159 =  n_3673 & ~n_16158;
assign n_16160 = ~n_16156 &  n_16159;
assign n_16161 = ~x_1727 & ~n_16160;
assign n_16162 = ~n_16151 &  n_16161;
assign n_16163 = ~n_3674 & ~n_4282;
assign n_16164 = ~x_1724 & ~n_16163;
assign n_16165 = ~n_4284 & ~n_3685;
assign n_16166 =  n_3695 &  n_16165;
assign n_16167 = ~n_16164 &  n_16166;
assign n_16168 = ~n_4287 &  n_16167;
assign n_16169 =  n_3673 &  n_16152;
assign n_16170 =  n_1328 & ~n_16154;
assign n_16171 =  n_3685 & ~n_16170;
assign n_16172 = ~n_16169 &  n_16171;
assign n_16173 =  x_1726 & ~n_16172;
assign n_16174 =  x_308 &  x_1721;
assign n_16175 =  x_1726 &  n_16174;
assign n_16176 =  n_3673 &  n_16175;
assign n_16177 = ~n_16173 & ~n_16176;
assign n_16178 = ~n_16168 & ~n_16177;
assign n_16179 = ~n_4289 & ~n_3686;
assign n_16180 = ~n_16178 &  n_16179;
assign n_16181 = ~n_16162 &  n_16180;
assign n_16182 = ~x_1728 &  n_16181;
assign n_16183 =  x_308 &  x_1725;
assign n_16184 =  n_1328 &  n_6031;
assign n_16185 =  n_1328 &  n_3685;
assign n_16186 =  n_3673 &  n_6031;
assign n_16187 = ~n_16185 & ~n_16186;
assign n_16188 =  n_4287 & ~n_16187;
assign n_16189 = ~n_16184 & ~n_16188;
assign n_16190 = ~n_3677 & ~n_3691;
assign n_16191 =  n_3673 &  n_3685;
assign n_16192 = ~n_16190 &  n_16191;
assign n_16193 =  n_16189 & ~n_16192;
assign n_16194 =  n_16183 & ~n_16193;
assign n_16195 = ~n_16194 &  n_16181;
assign n_16196 = ~x_308 & ~n_3691;
assign n_16197 = ~n_3673 &  n_3691;
assign n_16198 = ~n_16196 & ~n_16197;
assign n_16199 = ~x_1726 &  n_3691;
assign n_16200 = ~n_16125 & ~n_16199;
assign n_16201 = ~n_16198 & ~n_16200;
assign n_16202 = ~n_4287 & ~n_3685;
assign n_16203 =  x_1727 &  n_16202;
assign n_16204 = ~n_16201 &  n_16203;
assign n_16205 =  x_1725 & ~n_16142;
assign n_16206 = ~n_16138 & ~n_16205;
assign n_16207 = ~n_16204 &  n_16206;
assign n_16208 = ~n_16195 &  n_16207;
assign n_16209 = ~n_16182 & ~n_16208;
assign n_16210 = ~x_1721 & ~n_16125;
assign n_16211 =  n_16202 &  n_16210;
assign n_16212 = ~n_16174 & ~n_16211;
assign n_16213 =  x_1729 & ~n_16212;
assign n_16214 = ~n_3688 & ~n_16213;
assign n_16215 = ~n_16209 &  n_16214;
assign n_16216 =  x_1728 & ~n_16215;
assign n_16217 = ~x_1728 &  n_16215;
assign n_16218 = ~n_16216 & ~n_16217;
assign n_16219 =  x_308 & ~n_3677;
assign n_16220 =  n_3677 &  n_3685;
assign n_16221 = ~n_16219 & ~n_16220;
assign n_16222 =  n_16125 &  n_16221;
assign n_16223 = ~n_4287 & ~n_16222;
assign n_16224 =  x_1728 & ~n_16223;
assign n_16225 = ~x_308 & ~x_1728;
assign n_16226 = ~n_3685 &  n_16225;
assign n_16227 = ~n_3673 & ~n_16226;
assign n_16228 = ~n_16224 &  n_16227;
assign n_16229 = ~n_16195 &  n_16228;
assign n_16230 = ~x_1727 & ~n_16229;
assign n_16231 = ~n_16125 &  n_16197;
assign n_16232 = ~x_1722 & ~x_1726;
assign n_16233 =  n_3685 & ~n_16232;
assign n_16234 = ~x_1722 & ~x_1728;
assign n_16235 =  x_308 & ~n_16234;
assign n_16236 =  x_1727 & ~n_16235;
assign n_16237 = ~n_16233 &  n_16236;
assign n_16238 = ~n_16231 &  n_16237;
assign n_16239 = ~n_16195 &  n_16238;
assign n_16240 = ~n_16230 & ~n_16239;
assign n_16241 =  x_1727 &  n_16240;
assign n_16242 = ~x_1727 & ~n_16240;
assign n_16243 = ~n_16241 & ~n_16242;
assign n_16244 = ~n_3685 & ~n_16168;
assign n_16245 =  x_1726 & ~n_16244;
assign n_16246 =  n_4282 &  n_16231;
assign n_16247 = ~n_16220 & ~n_16246;
assign n_16248 =  n_4280 & ~n_16247;
assign n_16249 =  n_3685 &  n_3686;
assign n_16250 =  x_1724 &  n_16129;
assign n_16251 = ~n_16220 & ~n_16250;
assign n_16252 =  x_1729 & ~n_16251;
assign n_16253 = ~n_16249 & ~n_16252;
assign n_16254 = ~n_3673 & ~n_16253;
assign n_16255 = ~n_16248 & ~n_16254;
assign n_16256 = ~n_16245 &  n_16255;
assign n_16257 =  x_1726 & ~n_16256;
assign n_16258 = ~x_1726 &  n_16256;
assign n_16259 = ~n_16257 & ~n_16258;
assign n_16260 =  x_1725 & ~n_4291;
assign n_16261 = ~x_1725 &  n_4291;
assign n_16262 = ~n_16260 & ~n_16261;
assign n_16263 =  n_16247 &  n_16144;
assign n_16264 =  x_308 & ~n_16184;
assign n_16265 =  n_16264 & ~n_16192;
assign n_16266 =  x_1725 & ~n_16265;
assign n_16267 = ~n_16263 &  n_16266;
assign n_16268 =  n_16124 & ~n_16131;
assign n_16269 =  n_16268 & ~n_16222;
assign n_16270 = ~x_308 &  n_1328;
assign n_16271 =  n_3685 & ~n_16270;
assign n_16272 =  x_1726 & ~n_16271;
assign n_16273 = ~n_16272 & ~n_16176;
assign n_16274 =  n_16166 & ~n_16135;
assign n_16275 = ~n_16273 & ~n_16274;
assign n_16276 =  x_1728 &  n_16138;
assign n_16277 = ~x_308 &  n_6031;
assign n_16278 = ~n_16277 & ~n_16158;
assign n_16279 =  n_16276 & ~n_16278;
assign n_16280 = ~n_16275 & ~n_16279;
assign n_16281 = ~n_16269 &  n_16280;
assign n_16282 = ~n_16267 &  n_16281;
assign n_16283 =  n_16276 & ~n_16277;
assign n_16284 = ~x_1726 & ~n_16264;
assign n_16285 = ~n_16272 & ~n_16284;
assign n_16286 =  n_4284 &  n_16285;
assign n_16287 = ~n_16283 & ~n_16286;
assign n_16288 = ~n_16282 & ~n_16287;
assign n_16289 =  x_1724 &  n_16282;
assign n_16290 = ~n_16288 & ~n_16289;
assign n_16291 =  x_1724 & ~n_16290;
assign n_16292 = ~x_1724 &  n_16290;
assign n_16293 = ~n_16291 & ~n_16292;
assign n_16294 =  n_16276 &  n_16220;
assign n_16295 =  n_3673 &  n_16199;
assign n_16296 = ~x_1729 & ~n_16295;
assign n_16297 =  n_16285 &  n_16296;
assign n_16298 = ~n_16294 & ~n_16297;
assign n_16299 = ~n_16298 & ~n_16282;
assign n_16300 =  x_1723 &  n_16282;
assign n_16301 = ~n_16299 & ~n_16300;
assign n_16302 =  x_1723 & ~n_16301;
assign n_16303 = ~x_1723 &  n_16301;
assign n_16304 = ~n_16302 & ~n_16303;
assign n_16305 =  n_4280 & ~n_4286;
assign n_16306 =  n_16276 &  n_16156;
assign n_16307 = ~n_16305 & ~n_16306;
assign n_16308 = ~n_16268 &  n_16307;
assign n_16309 =  n_16183 & ~n_16189;
assign n_16310 = ~n_16167 &  n_16173;
assign n_16311 = ~n_16309 & ~n_16310;
assign n_16312 =  n_16308 &  n_16311;
assign n_16313 =  x_1722 &  n_16312;
assign n_16314 = ~n_3673 &  n_16285;
assign n_16315 = ~n_16196 &  n_3696;
assign n_16316 = ~n_3691 & ~n_3685;
assign n_16317 = ~x_308 & ~x_1726;
assign n_16318 = ~n_16316 &  n_16317;
assign n_16319 = ~n_16315 & ~n_16318;
assign n_16320 =  x_1724 & ~n_16197;
assign n_16321 = ~n_16319 &  n_16320;
assign n_16322 = ~n_16314 & ~n_16321;
assign n_16323 = ~x_1729 & ~n_16322;
assign n_16324 =  x_1724 &  x_1729;
assign n_16325 = ~n_16221 &  n_16324;
assign n_16326 = ~n_16283 & ~n_16325;
assign n_16327 = ~n_16323 &  n_16326;
assign n_16328 = ~n_16312 & ~n_16327;
assign n_16329 = ~n_16313 & ~n_16328;
assign n_16330 =  x_1722 & ~n_16329;
assign n_16331 = ~x_1722 &  n_16329;
assign n_16332 = ~n_16330 & ~n_16331;
assign n_16333 =  x_1723 &  n_16198;
assign n_16334 = ~n_16333 &  n_16272;
assign n_16335 =  x_1723 & ~n_16316;
assign n_16336 = ~x_308 & ~n_16335;
assign n_16337 = ~n_3673 & ~n_16196;
assign n_16338 = ~x_1729 & ~n_16337;
assign n_16339 = ~n_16336 &  n_16338;
assign n_16340 = ~x_1726 & ~n_16339;
assign n_16341 = ~n_16334 & ~n_16340;
assign n_16342 = ~n_3685 &  n_16283;
assign n_16343 =  x_1723 &  n_16124;
assign n_16344 = ~n_16221 &  n_16343;
assign n_16345 = ~n_16342 & ~n_16344;
assign n_16346 = ~n_16341 &  n_16345;
assign n_16347 = ~n_16312 & ~n_16346;
assign n_16348 =  x_1721 &  n_16312;
assign n_16349 = ~n_16347 & ~n_16348;
assign n_16350 =  x_1721 & ~n_16349;
assign n_16351 = ~x_1721 &  n_16349;
assign n_16352 = ~n_16350 & ~n_16351;
assign n_16353 =  x_1720 &  n_12453;
assign n_16354 = ~n_16353 & ~n_12458;
assign n_16355 =  x_1720 &  n_16354;
assign n_16356 = ~x_1720 & ~n_16354;
assign n_16357 = ~n_16355 & ~n_16356;
assign n_16358 = ~x_1749 & ~n_3243;
assign n_16359 =  x_1719 &  n_16358;
assign n_16360 = ~x_1719 & ~n_16358;
assign n_16361 = ~n_16359 & ~n_16360;
assign n_16362 =  x_1761 &  n_12515;
assign n_16363 =  x_1718 &  n_16362;
assign n_16364 = ~x_1718 & ~n_16362;
assign n_16365 = ~n_16363 & ~n_16364;
assign n_16366 =  x_1725 &  x_1726;
assign n_16367 =  x_1729 & ~n_4368;
assign n_16368 = ~n_16366 & ~n_16367;
assign n_16369 =  x_1717 & ~n_16368;
assign n_16370 = ~x_1717 &  n_16368;
assign n_16371 = ~n_16369 & ~n_16370;
assign n_16372 =  x_1716 & ~n_1761;
assign n_16373 =  x_1917 &  n_1761;
assign n_16374 = ~n_16372 & ~n_16373;
assign n_16375 =  x_1716 & ~n_16374;
assign n_16376 = ~x_1716 &  n_16374;
assign n_16377 = ~n_16375 & ~n_16376;
assign n_16378 =  x_1715 & ~n_1770;
assign n_16379 =  x_1917 &  n_1770;
assign n_16380 = ~n_16378 & ~n_16379;
assign n_16381 =  x_1715 & ~n_16380;
assign n_16382 = ~x_1715 &  n_16380;
assign n_16383 = ~n_16381 & ~n_16382;
assign n_16384 =  x_1714 & ~n_1778;
assign n_16385 =  x_1917 &  n_1778;
assign n_16386 = ~n_16384 & ~n_16385;
assign n_16387 =  x_1714 & ~n_16386;
assign n_16388 = ~x_1714 &  n_16386;
assign n_16389 = ~n_16387 & ~n_16388;
assign n_16390 =  x_1713 & ~n_1785;
assign n_16391 =  x_1917 &  n_1785;
assign n_16392 = ~n_16390 & ~n_16391;
assign n_16393 =  x_1713 & ~n_16392;
assign n_16394 = ~x_1713 &  n_16392;
assign n_16395 = ~n_16393 & ~n_16394;
assign n_16396 =  x_1712 & ~n_1792;
assign n_16397 =  x_1917 &  n_1792;
assign n_16398 = ~n_16396 & ~n_16397;
assign n_16399 =  x_1712 & ~n_16398;
assign n_16400 = ~x_1712 &  n_16398;
assign n_16401 = ~n_16399 & ~n_16400;
assign n_16402 =  x_1711 & ~n_1799;
assign n_16403 =  x_1917 &  n_1799;
assign n_16404 = ~n_16402 & ~n_16403;
assign n_16405 =  x_1711 & ~n_16404;
assign n_16406 = ~x_1711 &  n_16404;
assign n_16407 = ~n_16405 & ~n_16406;
assign n_16408 =  x_1710 & ~n_1806;
assign n_16409 =  x_1917 &  n_1806;
assign n_16410 = ~n_16408 & ~n_16409;
assign n_16411 =  x_1710 & ~n_16410;
assign n_16412 = ~x_1710 &  n_16410;
assign n_16413 = ~n_16411 & ~n_16412;
assign n_16414 =  x_1709 & ~n_1750;
assign n_16415 =  x_1917 &  n_1750;
assign n_16416 = ~n_16414 & ~n_16415;
assign n_16417 =  x_1709 & ~n_16416;
assign n_16418 = ~x_1709 &  n_16416;
assign n_16419 = ~n_16417 & ~n_16418;
assign n_16420 =  x_1708 & ~n_1761;
assign n_16421 = ~x_1908 &  n_1761;
assign n_16422 = ~n_16420 & ~n_16421;
assign n_16423 =  x_1708 & ~n_16422;
assign n_16424 = ~x_1708 &  n_16422;
assign n_16425 = ~n_16423 & ~n_16424;
assign n_16426 =  x_1707 & ~n_1770;
assign n_16427 = ~x_1908 &  n_1770;
assign n_16428 = ~n_16426 & ~n_16427;
assign n_16429 =  x_1707 & ~n_16428;
assign n_16430 = ~x_1707 &  n_16428;
assign n_16431 = ~n_16429 & ~n_16430;
assign n_16432 =  x_1706 & ~n_1778;
assign n_16433 = ~x_1908 &  n_1778;
assign n_16434 = ~n_16432 & ~n_16433;
assign n_16435 =  x_1706 & ~n_16434;
assign n_16436 = ~x_1706 &  n_16434;
assign n_16437 = ~n_16435 & ~n_16436;
assign n_16438 =  x_1705 & ~n_1785;
assign n_16439 = ~x_1908 &  n_1785;
assign n_16440 = ~n_16438 & ~n_16439;
assign n_16441 =  x_1705 & ~n_16440;
assign n_16442 = ~x_1705 &  n_16440;
assign n_16443 = ~n_16441 & ~n_16442;
assign n_16444 =  x_1704 & ~n_1792;
assign n_16445 = ~x_1908 &  n_1792;
assign n_16446 = ~n_16444 & ~n_16445;
assign n_16447 =  x_1704 & ~n_16446;
assign n_16448 = ~x_1704 &  n_16446;
assign n_16449 = ~n_16447 & ~n_16448;
assign n_16450 =  x_1703 & ~n_1799;
assign n_16451 = ~x_1908 &  n_1799;
assign n_16452 = ~n_16450 & ~n_16451;
assign n_16453 =  x_1703 & ~n_16452;
assign n_16454 = ~x_1703 &  n_16452;
assign n_16455 = ~n_16453 & ~n_16454;
assign n_16456 =  x_1702 & ~n_1806;
assign n_16457 = ~x_1908 &  n_1806;
assign n_16458 = ~n_16456 & ~n_16457;
assign n_16459 =  x_1702 & ~n_16458;
assign n_16460 = ~x_1702 &  n_16458;
assign n_16461 = ~n_16459 & ~n_16460;
assign n_16462 =  x_1701 & ~n_1750;
assign n_16463 = ~x_1908 &  n_1750;
assign n_16464 = ~n_16462 & ~n_16463;
assign n_16465 =  x_1701 & ~n_16464;
assign n_16466 = ~x_1701 &  n_16464;
assign n_16467 = ~n_16465 & ~n_16466;
assign n_16468 =  x_1700 & ~n_1761;
assign n_16469 =  x_1899 &  n_1761;
assign n_16470 = ~n_16468 & ~n_16469;
assign n_16471 =  x_1700 & ~n_16470;
assign n_16472 = ~x_1700 &  n_16470;
assign n_16473 = ~n_16471 & ~n_16472;
assign n_16474 =  x_1699 & ~n_1770;
assign n_16475 =  x_1899 &  n_1770;
assign n_16476 = ~n_16474 & ~n_16475;
assign n_16477 =  x_1699 & ~n_16476;
assign n_16478 = ~x_1699 &  n_16476;
assign n_16479 = ~n_16477 & ~n_16478;
assign n_16480 =  x_1698 & ~n_1778;
assign n_16481 =  x_1899 &  n_1778;
assign n_16482 = ~n_16480 & ~n_16481;
assign n_16483 =  x_1698 & ~n_16482;
assign n_16484 = ~x_1698 &  n_16482;
assign n_16485 = ~n_16483 & ~n_16484;
assign n_16486 =  x_1697 & ~n_1785;
assign n_16487 =  x_1899 &  n_1785;
assign n_16488 = ~n_16486 & ~n_16487;
assign n_16489 =  x_1697 & ~n_16488;
assign n_16490 = ~x_1697 &  n_16488;
assign n_16491 = ~n_16489 & ~n_16490;
assign n_16492 =  x_1696 & ~n_1792;
assign n_16493 =  x_1899 &  n_1792;
assign n_16494 = ~n_16492 & ~n_16493;
assign n_16495 =  x_1696 & ~n_16494;
assign n_16496 = ~x_1696 &  n_16494;
assign n_16497 = ~n_16495 & ~n_16496;
assign n_16498 =  x_1695 & ~n_1799;
assign n_16499 =  x_1899 &  n_1799;
assign n_16500 = ~n_16498 & ~n_16499;
assign n_16501 =  x_1695 & ~n_16500;
assign n_16502 = ~x_1695 &  n_16500;
assign n_16503 = ~n_16501 & ~n_16502;
assign n_16504 =  x_1694 & ~n_1806;
assign n_16505 =  x_1899 &  n_1806;
assign n_16506 = ~n_16504 & ~n_16505;
assign n_16507 =  x_1694 & ~n_16506;
assign n_16508 = ~x_1694 &  n_16506;
assign n_16509 = ~n_16507 & ~n_16508;
assign n_16510 =  x_1693 & ~n_1750;
assign n_16511 =  x_1899 &  n_1750;
assign n_16512 = ~n_16510 & ~n_16511;
assign n_16513 =  x_1693 & ~n_16512;
assign n_16514 = ~x_1693 &  n_16512;
assign n_16515 = ~n_16513 & ~n_16514;
assign n_16516 =  x_1692 & ~n_1761;
assign n_16517 = ~x_1890 &  n_1761;
assign n_16518 = ~n_16516 & ~n_16517;
assign n_16519 =  x_1692 & ~n_16518;
assign n_16520 = ~x_1692 &  n_16518;
assign n_16521 = ~n_16519 & ~n_16520;
assign n_16522 =  x_1691 & ~n_1770;
assign n_16523 = ~x_1890 &  n_1770;
assign n_16524 = ~n_16522 & ~n_16523;
assign n_16525 =  x_1691 & ~n_16524;
assign n_16526 = ~x_1691 &  n_16524;
assign n_16527 = ~n_16525 & ~n_16526;
assign n_16528 =  x_1690 & ~n_1778;
assign n_16529 = ~x_1890 &  n_1778;
assign n_16530 = ~n_16528 & ~n_16529;
assign n_16531 =  x_1690 & ~n_16530;
assign n_16532 = ~x_1690 &  n_16530;
assign n_16533 = ~n_16531 & ~n_16532;
assign n_16534 =  x_1689 & ~n_1785;
assign n_16535 = ~x_1890 &  n_1785;
assign n_16536 = ~n_16534 & ~n_16535;
assign n_16537 =  x_1689 & ~n_16536;
assign n_16538 = ~x_1689 &  n_16536;
assign n_16539 = ~n_16537 & ~n_16538;
assign n_16540 =  x_1688 & ~n_1792;
assign n_16541 = ~x_1890 &  n_1792;
assign n_16542 = ~n_16540 & ~n_16541;
assign n_16543 =  x_1688 & ~n_16542;
assign n_16544 = ~x_1688 &  n_16542;
assign n_16545 = ~n_16543 & ~n_16544;
assign n_16546 =  x_1687 & ~n_1799;
assign n_16547 = ~x_1890 &  n_1799;
assign n_16548 = ~n_16546 & ~n_16547;
assign n_16549 =  x_1687 & ~n_16548;
assign n_16550 = ~x_1687 &  n_16548;
assign n_16551 = ~n_16549 & ~n_16550;
assign n_16552 =  x_1686 & ~n_1806;
assign n_16553 = ~x_1890 &  n_1806;
assign n_16554 = ~n_16552 & ~n_16553;
assign n_16555 =  x_1686 & ~n_16554;
assign n_16556 = ~x_1686 &  n_16554;
assign n_16557 = ~n_16555 & ~n_16556;
assign n_16558 =  x_1685 & ~n_1750;
assign n_16559 = ~x_1890 &  n_1750;
assign n_16560 = ~n_16558 & ~n_16559;
assign n_16561 =  x_1685 & ~n_16560;
assign n_16562 = ~x_1685 &  n_16560;
assign n_16563 = ~n_16561 & ~n_16562;
assign n_16564 =  x_1684 & ~n_1761;
assign n_16565 =  x_1881 &  n_1761;
assign n_16566 = ~n_16564 & ~n_16565;
assign n_16567 =  x_1684 & ~n_16566;
assign n_16568 = ~x_1684 &  n_16566;
assign n_16569 = ~n_16567 & ~n_16568;
assign n_16570 =  x_1683 & ~n_1770;
assign n_16571 =  x_1881 &  n_1770;
assign n_16572 = ~n_16570 & ~n_16571;
assign n_16573 =  x_1683 & ~n_16572;
assign n_16574 = ~x_1683 &  n_16572;
assign n_16575 = ~n_16573 & ~n_16574;
assign n_16576 =  x_1682 & ~n_1778;
assign n_16577 =  x_1881 &  n_1778;
assign n_16578 = ~n_16576 & ~n_16577;
assign n_16579 =  x_1682 & ~n_16578;
assign n_16580 = ~x_1682 &  n_16578;
assign n_16581 = ~n_16579 & ~n_16580;
assign n_16582 =  x_1681 & ~n_1785;
assign n_16583 =  x_1881 &  n_1785;
assign n_16584 = ~n_16582 & ~n_16583;
assign n_16585 =  x_1681 & ~n_16584;
assign n_16586 = ~x_1681 &  n_16584;
assign n_16587 = ~n_16585 & ~n_16586;
assign n_16588 =  x_1680 & ~n_1792;
assign n_16589 =  x_1881 &  n_1792;
assign n_16590 = ~n_16588 & ~n_16589;
assign n_16591 =  x_1680 & ~n_16590;
assign n_16592 = ~x_1680 &  n_16590;
assign n_16593 = ~n_16591 & ~n_16592;
assign n_16594 =  x_1679 & ~n_1799;
assign n_16595 =  x_1881 &  n_1799;
assign n_16596 = ~n_16594 & ~n_16595;
assign n_16597 =  x_1679 & ~n_16596;
assign n_16598 = ~x_1679 &  n_16596;
assign n_16599 = ~n_16597 & ~n_16598;
assign n_16600 =  x_1678 & ~n_1806;
assign n_16601 =  x_1881 &  n_1806;
assign n_16602 = ~n_16600 & ~n_16601;
assign n_16603 =  x_1678 & ~n_16602;
assign n_16604 = ~x_1678 &  n_16602;
assign n_16605 = ~n_16603 & ~n_16604;
assign n_16606 =  x_1677 & ~n_1750;
assign n_16607 =  x_1881 &  n_1750;
assign n_16608 = ~n_16606 & ~n_16607;
assign n_16609 =  x_1677 & ~n_16608;
assign n_16610 = ~x_1677 &  n_16608;
assign n_16611 = ~n_16609 & ~n_16610;
assign n_16612 =  x_1676 & ~n_1761;
assign n_16613 = ~x_1872 &  n_1761;
assign n_16614 = ~n_16612 & ~n_16613;
assign n_16615 =  x_1676 & ~n_16614;
assign n_16616 = ~x_1676 &  n_16614;
assign n_16617 = ~n_16615 & ~n_16616;
assign n_16618 =  x_1675 & ~n_1770;
assign n_16619 = ~x_1872 &  n_1770;
assign n_16620 = ~n_16618 & ~n_16619;
assign n_16621 =  x_1675 & ~n_16620;
assign n_16622 = ~x_1675 &  n_16620;
assign n_16623 = ~n_16621 & ~n_16622;
assign n_16624 =  x_1674 & ~n_1778;
assign n_16625 = ~x_1872 &  n_1778;
assign n_16626 = ~n_16624 & ~n_16625;
assign n_16627 =  x_1674 & ~n_16626;
assign n_16628 = ~x_1674 &  n_16626;
assign n_16629 = ~n_16627 & ~n_16628;
assign n_16630 =  x_1673 & ~n_1785;
assign n_16631 = ~x_1872 &  n_1785;
assign n_16632 = ~n_16630 & ~n_16631;
assign n_16633 =  x_1673 & ~n_16632;
assign n_16634 = ~x_1673 &  n_16632;
assign n_16635 = ~n_16633 & ~n_16634;
assign n_16636 =  x_1672 & ~n_1792;
assign n_16637 = ~x_1872 &  n_1792;
assign n_16638 = ~n_16636 & ~n_16637;
assign n_16639 =  x_1672 & ~n_16638;
assign n_16640 = ~x_1672 &  n_16638;
assign n_16641 = ~n_16639 & ~n_16640;
assign n_16642 =  x_1671 & ~n_1799;
assign n_16643 = ~x_1872 &  n_1799;
assign n_16644 = ~n_16642 & ~n_16643;
assign n_16645 =  x_1671 & ~n_16644;
assign n_16646 = ~x_1671 &  n_16644;
assign n_16647 = ~n_16645 & ~n_16646;
assign n_16648 =  x_1670 & ~n_1806;
assign n_16649 = ~x_1872 &  n_1806;
assign n_16650 = ~n_16648 & ~n_16649;
assign n_16651 =  x_1670 & ~n_16650;
assign n_16652 = ~x_1670 &  n_16650;
assign n_16653 = ~n_16651 & ~n_16652;
assign n_16654 =  x_1669 & ~n_1750;
assign n_16655 = ~x_1872 &  n_1750;
assign n_16656 = ~n_16654 & ~n_16655;
assign n_16657 =  x_1669 & ~n_16656;
assign n_16658 = ~x_1669 &  n_16656;
assign n_16659 = ~n_16657 & ~n_16658;
assign n_16660 =  x_1668 & ~n_1761;
assign n_16661 =  x_1863 &  n_1761;
assign n_16662 = ~n_16660 & ~n_16661;
assign n_16663 =  x_1668 & ~n_16662;
assign n_16664 = ~x_1668 &  n_16662;
assign n_16665 = ~n_16663 & ~n_16664;
assign n_16666 =  x_1667 & ~n_1770;
assign n_16667 =  x_1863 &  n_1770;
assign n_16668 = ~n_16666 & ~n_16667;
assign n_16669 =  x_1667 & ~n_16668;
assign n_16670 = ~x_1667 &  n_16668;
assign n_16671 = ~n_16669 & ~n_16670;
assign n_16672 =  x_1666 & ~n_1778;
assign n_16673 =  x_1863 &  n_1778;
assign n_16674 = ~n_16672 & ~n_16673;
assign n_16675 =  x_1666 & ~n_16674;
assign n_16676 = ~x_1666 &  n_16674;
assign n_16677 = ~n_16675 & ~n_16676;
assign n_16678 =  x_1665 & ~n_1785;
assign n_16679 =  x_1863 &  n_1785;
assign n_16680 = ~n_16678 & ~n_16679;
assign n_16681 =  x_1665 & ~n_16680;
assign n_16682 = ~x_1665 &  n_16680;
assign n_16683 = ~n_16681 & ~n_16682;
assign n_16684 =  x_1664 & ~n_1792;
assign n_16685 =  x_1863 &  n_1792;
assign n_16686 = ~n_16684 & ~n_16685;
assign n_16687 =  x_1664 & ~n_16686;
assign n_16688 = ~x_1664 &  n_16686;
assign n_16689 = ~n_16687 & ~n_16688;
assign n_16690 =  x_1663 & ~n_1799;
assign n_16691 =  x_1863 &  n_1799;
assign n_16692 = ~n_16690 & ~n_16691;
assign n_16693 =  x_1663 & ~n_16692;
assign n_16694 = ~x_1663 &  n_16692;
assign n_16695 = ~n_16693 & ~n_16694;
assign n_16696 =  x_1662 & ~n_1806;
assign n_16697 =  x_1863 &  n_1806;
assign n_16698 = ~n_16696 & ~n_16697;
assign n_16699 =  x_1662 & ~n_16698;
assign n_16700 = ~x_1662 &  n_16698;
assign n_16701 = ~n_16699 & ~n_16700;
assign n_16702 =  x_1661 & ~n_1750;
assign n_16703 =  x_1863 &  n_1750;
assign n_16704 = ~n_16702 & ~n_16703;
assign n_16705 =  x_1661 & ~n_16704;
assign n_16706 = ~x_1661 &  n_16704;
assign n_16707 = ~n_16705 & ~n_16706;
assign n_16708 =  x_1660 & ~n_1761;
assign n_16709 = ~x_1862 &  n_1761;
assign n_16710 = ~n_16708 & ~n_16709;
assign n_16711 =  x_1660 & ~n_16710;
assign n_16712 = ~x_1660 &  n_16710;
assign n_16713 = ~n_16711 & ~n_16712;
assign n_16714 =  x_1659 & ~n_1770;
assign n_16715 = ~x_1862 &  n_1770;
assign n_16716 = ~n_16714 & ~n_16715;
assign n_16717 =  x_1659 & ~n_16716;
assign n_16718 = ~x_1659 &  n_16716;
assign n_16719 = ~n_16717 & ~n_16718;
assign n_16720 =  x_1658 & ~n_1778;
assign n_16721 = ~x_1862 &  n_1778;
assign n_16722 = ~n_16720 & ~n_16721;
assign n_16723 =  x_1658 & ~n_16722;
assign n_16724 = ~x_1658 &  n_16722;
assign n_16725 = ~n_16723 & ~n_16724;
assign n_16726 =  x_1657 & ~n_1785;
assign n_16727 = ~x_1862 &  n_1785;
assign n_16728 = ~n_16726 & ~n_16727;
assign n_16729 =  x_1657 & ~n_16728;
assign n_16730 = ~x_1657 &  n_16728;
assign n_16731 = ~n_16729 & ~n_16730;
assign n_16732 =  x_1656 & ~n_1792;
assign n_16733 = ~x_1862 &  n_1792;
assign n_16734 = ~n_16732 & ~n_16733;
assign n_16735 =  x_1656 & ~n_16734;
assign n_16736 = ~x_1656 &  n_16734;
assign n_16737 = ~n_16735 & ~n_16736;
assign n_16738 =  x_1655 & ~n_1799;
assign n_16739 = ~x_1862 &  n_1799;
assign n_16740 = ~n_16738 & ~n_16739;
assign n_16741 =  x_1655 & ~n_16740;
assign n_16742 = ~x_1655 &  n_16740;
assign n_16743 = ~n_16741 & ~n_16742;
assign n_16744 =  x_1654 & ~n_1806;
assign n_16745 = ~x_1862 &  n_1806;
assign n_16746 = ~n_16744 & ~n_16745;
assign n_16747 =  x_1654 & ~n_16746;
assign n_16748 = ~x_1654 &  n_16746;
assign n_16749 = ~n_16747 & ~n_16748;
assign n_16750 =  x_1653 & ~n_1750;
assign n_16751 = ~x_1862 &  n_1750;
assign n_16752 = ~n_16750 & ~n_16751;
assign n_16753 =  x_1653 & ~n_16752;
assign n_16754 = ~x_1653 &  n_16752;
assign n_16755 = ~n_16753 & ~n_16754;
assign n_16756 =  x_1652 & ~n_1719;
assign n_16757 = ~x_1652 &  n_1719;
assign n_16758 = ~n_16756 & ~n_16757;
assign n_16759 = ~x_1562 &  x_1736;
assign n_16760 =  x_1651 & ~n_16759;
assign n_16761 =  x_1845 &  n_16759;
assign n_16762 = ~n_16760 & ~n_16761;
assign n_16763 =  x_1651 & ~n_16762;
assign n_16764 = ~x_1651 &  n_16762;
assign n_16765 = ~n_16763 & ~n_16764;
assign n_16766 =  x_1650 & ~n_16759;
assign n_16767 =  x_1844 &  n_16759;
assign n_16768 = ~n_16766 & ~n_16767;
assign n_16769 =  x_1650 & ~n_16768;
assign n_16770 = ~x_1650 &  n_16768;
assign n_16771 = ~n_16769 & ~n_16770;
assign n_16772 =  x_1649 & ~n_16759;
assign n_16773 =  x_1843 &  n_16759;
assign n_16774 = ~n_16772 & ~n_16773;
assign n_16775 =  x_1649 & ~n_16774;
assign n_16776 = ~x_1649 &  n_16774;
assign n_16777 = ~n_16775 & ~n_16776;
assign n_16778 =  x_1648 & ~n_16759;
assign n_16779 =  x_1842 &  n_16759;
assign n_16780 = ~n_16778 & ~n_16779;
assign n_16781 =  x_1648 & ~n_16780;
assign n_16782 = ~x_1648 &  n_16780;
assign n_16783 = ~n_16781 & ~n_16782;
assign n_16784 =  x_1647 & ~n_16759;
assign n_16785 =  x_1841 &  n_16759;
assign n_16786 = ~n_16784 & ~n_16785;
assign n_16787 =  x_1647 & ~n_16786;
assign n_16788 = ~x_1647 &  n_16786;
assign n_16789 = ~n_16787 & ~n_16788;
assign n_16790 =  x_1646 & ~n_16759;
assign n_16791 =  x_1840 &  n_16759;
assign n_16792 = ~n_16790 & ~n_16791;
assign n_16793 =  x_1646 & ~n_16792;
assign n_16794 = ~x_1646 &  n_16792;
assign n_16795 = ~n_16793 & ~n_16794;
assign n_16796 =  x_1645 & ~n_16759;
assign n_16797 =  x_1839 &  n_16759;
assign n_16798 = ~n_16796 & ~n_16797;
assign n_16799 =  x_1645 & ~n_16798;
assign n_16800 = ~x_1645 &  n_16798;
assign n_16801 = ~n_16799 & ~n_16800;
assign n_16802 =  x_1644 & ~n_16759;
assign n_16803 =  x_1838 &  n_16759;
assign n_16804 = ~n_16802 & ~n_16803;
assign n_16805 =  x_1644 & ~n_16804;
assign n_16806 = ~x_1644 &  n_16804;
assign n_16807 = ~n_16805 & ~n_16806;
assign n_16808 =  x_1643 & ~n_16759;
assign n_16809 =  x_1837 &  n_16759;
assign n_16810 = ~n_16808 & ~n_16809;
assign n_16811 =  x_1643 & ~n_16810;
assign n_16812 = ~x_1643 &  n_16810;
assign n_16813 = ~n_16811 & ~n_16812;
assign n_16814 =  x_1642 & ~n_16759;
assign n_16815 =  x_1836 &  n_16759;
assign n_16816 = ~n_16814 & ~n_16815;
assign n_16817 =  x_1642 & ~n_16816;
assign n_16818 = ~x_1642 &  n_16816;
assign n_16819 = ~n_16817 & ~n_16818;
assign n_16820 =  x_1641 & ~n_16759;
assign n_16821 =  x_1835 &  n_16759;
assign n_16822 = ~n_16820 & ~n_16821;
assign n_16823 =  x_1641 & ~n_16822;
assign n_16824 = ~x_1641 &  n_16822;
assign n_16825 = ~n_16823 & ~n_16824;
assign n_16826 =  x_1640 & ~n_16759;
assign n_16827 =  x_1834 &  n_16759;
assign n_16828 = ~n_16826 & ~n_16827;
assign n_16829 =  x_1640 & ~n_16828;
assign n_16830 = ~x_1640 &  n_16828;
assign n_16831 = ~n_16829 & ~n_16830;
assign n_16832 =  x_1639 & ~n_16759;
assign n_16833 =  x_1833 &  n_16759;
assign n_16834 = ~n_16832 & ~n_16833;
assign n_16835 =  x_1639 & ~n_16834;
assign n_16836 = ~x_1639 &  n_16834;
assign n_16837 = ~n_16835 & ~n_16836;
assign n_16838 =  x_1638 & ~n_16759;
assign n_16839 =  x_1832 &  n_16759;
assign n_16840 = ~n_16838 & ~n_16839;
assign n_16841 =  x_1638 & ~n_16840;
assign n_16842 = ~x_1638 &  n_16840;
assign n_16843 = ~n_16841 & ~n_16842;
assign n_16844 =  x_1637 & ~n_16759;
assign n_16845 =  x_1831 &  n_16759;
assign n_16846 = ~n_16844 & ~n_16845;
assign n_16847 =  x_1637 & ~n_16846;
assign n_16848 = ~x_1637 &  n_16846;
assign n_16849 = ~n_16847 & ~n_16848;
assign n_16850 =  x_1636 & ~n_16759;
assign n_16851 =  x_1830 &  n_16759;
assign n_16852 = ~n_16850 & ~n_16851;
assign n_16853 =  x_1636 & ~n_16852;
assign n_16854 = ~x_1636 &  n_16852;
assign n_16855 = ~n_16853 & ~n_16854;
assign n_16856 =  x_1635 & ~n_16759;
assign n_16857 =  x_1829 &  n_16759;
assign n_16858 = ~n_16856 & ~n_16857;
assign n_16859 =  x_1635 & ~n_16858;
assign n_16860 = ~x_1635 &  n_16858;
assign n_16861 = ~n_16859 & ~n_16860;
assign n_16862 =  x_1634 & ~n_16759;
assign n_16863 =  x_1828 &  n_16759;
assign n_16864 = ~n_16862 & ~n_16863;
assign n_16865 =  x_1634 & ~n_16864;
assign n_16866 = ~x_1634 &  n_16864;
assign n_16867 = ~n_16865 & ~n_16866;
assign n_16868 =  x_1633 & ~n_16759;
assign n_16869 =  x_1827 &  n_16759;
assign n_16870 = ~n_16868 & ~n_16869;
assign n_16871 =  x_1633 & ~n_16870;
assign n_16872 = ~x_1633 &  n_16870;
assign n_16873 = ~n_16871 & ~n_16872;
assign n_16874 =  x_1632 & ~n_16759;
assign n_16875 =  x_1826 &  n_16759;
assign n_16876 = ~n_16874 & ~n_16875;
assign n_16877 =  x_1632 & ~n_16876;
assign n_16878 = ~x_1632 &  n_16876;
assign n_16879 = ~n_16877 & ~n_16878;
assign n_16880 =  x_1631 & ~n_16759;
assign n_16881 =  x_1825 &  n_16759;
assign n_16882 = ~n_16880 & ~n_16881;
assign n_16883 =  x_1631 & ~n_16882;
assign n_16884 = ~x_1631 &  n_16882;
assign n_16885 = ~n_16883 & ~n_16884;
assign n_16886 =  x_1630 & ~n_16759;
assign n_16887 =  x_1824 &  n_16759;
assign n_16888 = ~n_16886 & ~n_16887;
assign n_16889 =  x_1630 & ~n_16888;
assign n_16890 = ~x_1630 &  n_16888;
assign n_16891 = ~n_16889 & ~n_16890;
assign n_16892 =  x_1629 & ~n_16759;
assign n_16893 =  x_1823 &  n_16759;
assign n_16894 = ~n_16892 & ~n_16893;
assign n_16895 =  x_1629 & ~n_16894;
assign n_16896 = ~x_1629 &  n_16894;
assign n_16897 = ~n_16895 & ~n_16896;
assign n_16898 =  x_1628 & ~n_16759;
assign n_16899 =  x_1822 &  n_16759;
assign n_16900 = ~n_16898 & ~n_16899;
assign n_16901 =  x_1628 & ~n_16900;
assign n_16902 = ~x_1628 &  n_16900;
assign n_16903 = ~n_16901 & ~n_16902;
assign n_16904 =  x_1627 & ~n_16759;
assign n_16905 =  x_1821 &  n_16759;
assign n_16906 = ~n_16904 & ~n_16905;
assign n_16907 =  x_1627 & ~n_16906;
assign n_16908 = ~x_1627 &  n_16906;
assign n_16909 = ~n_16907 & ~n_16908;
assign n_16910 =  x_1626 & ~n_16759;
assign n_16911 =  x_1820 &  n_16759;
assign n_16912 = ~n_16910 & ~n_16911;
assign n_16913 =  x_1626 & ~n_16912;
assign n_16914 = ~x_1626 &  n_16912;
assign n_16915 = ~n_16913 & ~n_16914;
assign n_16916 =  x_1625 & ~n_16759;
assign n_16917 =  x_1819 &  n_16759;
assign n_16918 = ~n_16916 & ~n_16917;
assign n_16919 =  x_1625 & ~n_16918;
assign n_16920 = ~x_1625 &  n_16918;
assign n_16921 = ~n_16919 & ~n_16920;
assign n_16922 =  x_1624 & ~n_16759;
assign n_16923 =  x_1818 &  n_16759;
assign n_16924 = ~n_16922 & ~n_16923;
assign n_16925 =  x_1624 & ~n_16924;
assign n_16926 = ~x_1624 &  n_16924;
assign n_16927 = ~n_16925 & ~n_16926;
assign n_16928 =  x_1623 & ~n_16759;
assign n_16929 =  x_1817 &  n_16759;
assign n_16930 = ~n_16928 & ~n_16929;
assign n_16931 =  x_1623 & ~n_16930;
assign n_16932 = ~x_1623 &  n_16930;
assign n_16933 = ~n_16931 & ~n_16932;
assign n_16934 =  x_1622 & ~n_16759;
assign n_16935 =  x_1816 &  n_16759;
assign n_16936 = ~n_16934 & ~n_16935;
assign n_16937 =  x_1622 & ~n_16936;
assign n_16938 = ~x_1622 &  n_16936;
assign n_16939 = ~n_16937 & ~n_16938;
assign n_16940 =  x_1621 & ~n_16759;
assign n_16941 =  x_1815 &  n_16759;
assign n_16942 = ~n_16940 & ~n_16941;
assign n_16943 =  x_1621 & ~n_16942;
assign n_16944 = ~x_1621 &  n_16942;
assign n_16945 = ~n_16943 & ~n_16944;
assign n_16946 =  x_1620 & ~n_16759;
assign n_16947 =  x_1814 &  n_16759;
assign n_16948 = ~n_16946 & ~n_16947;
assign n_16949 =  x_1620 & ~n_16948;
assign n_16950 = ~x_1620 &  n_16948;
assign n_16951 = ~n_16949 & ~n_16950;
assign n_16952 =  x_1619 & ~n_16759;
assign n_16953 =  x_1813 &  n_16759;
assign n_16954 = ~n_16952 & ~n_16953;
assign n_16955 =  x_1619 & ~n_16954;
assign n_16956 = ~x_1619 &  n_16954;
assign n_16957 = ~n_16955 & ~n_16956;
assign n_16958 =  x_1618 &  n_16759;
assign n_16959 = ~x_1618 & ~n_16759;
assign n_16960 = ~n_16958 & ~n_16959;
assign n_16961 =  x_1617 & ~n_1785;
assign n_16962 = ~x_1763 &  n_1785;
assign n_16963 = ~n_16961 & ~n_16962;
assign n_16964 =  x_1617 & ~n_16963;
assign n_16965 = ~x_1617 &  n_16963;
assign n_16966 = ~n_16964 & ~n_16965;
assign n_16967 =  x_1616 & ~n_1778;
assign n_16968 = ~x_1763 &  n_1778;
assign n_16969 = ~n_16967 & ~n_16968;
assign n_16970 =  x_1616 & ~n_16969;
assign n_16971 = ~x_1616 &  n_16969;
assign n_16972 = ~n_16970 & ~n_16971;
assign n_16973 =  x_1615 & ~n_1799;
assign n_16974 = ~x_1763 &  n_1799;
assign n_16975 = ~n_16973 & ~n_16974;
assign n_16976 =  x_1615 & ~n_16975;
assign n_16977 = ~x_1615 &  n_16975;
assign n_16978 = ~n_16976 & ~n_16977;
assign n_16979 =  x_1614 & ~n_1792;
assign n_16980 = ~x_1763 &  n_1792;
assign n_16981 = ~n_16979 & ~n_16980;
assign n_16982 =  x_1614 & ~n_16981;
assign n_16983 = ~x_1614 &  n_16981;
assign n_16984 = ~n_16982 & ~n_16983;
assign n_16985 =  x_1613 & ~n_1770;
assign n_16986 = ~x_1763 &  n_1770;
assign n_16987 = ~n_16985 & ~n_16986;
assign n_16988 =  x_1613 & ~n_16987;
assign n_16989 = ~x_1613 &  n_16987;
assign n_16990 = ~n_16988 & ~n_16989;
assign n_16991 =  x_1612 & ~n_1750;
assign n_16992 = ~x_1763 &  n_1750;
assign n_16993 = ~n_16991 & ~n_16992;
assign n_16994 =  x_1612 & ~n_16993;
assign n_16995 = ~x_1612 &  n_16993;
assign n_16996 = ~n_16994 & ~n_16995;
assign n_16997 =  x_1611 & ~n_1806;
assign n_16998 = ~x_1763 &  n_1806;
assign n_16999 = ~n_16997 & ~n_16998;
assign n_17000 =  x_1611 & ~n_16999;
assign n_17001 = ~x_1611 &  n_16999;
assign n_17002 = ~n_17000 & ~n_17001;
assign n_17003 =  x_1610 & ~n_1761;
assign n_17004 = ~x_1763 &  n_1761;
assign n_17005 = ~n_17003 & ~n_17004;
assign n_17006 =  x_1610 & ~n_17005;
assign n_17007 = ~x_1610 &  n_17005;
assign n_17008 = ~n_17006 & ~n_17007;
assign n_17009 =  x_1609 & ~n_1785;
assign n_17010 = ~x_1752 &  n_1785;
assign n_17011 = ~n_17009 & ~n_17010;
assign n_17012 =  x_1609 & ~n_17011;
assign n_17013 = ~x_1609 &  n_17011;
assign n_17014 = ~n_17012 & ~n_17013;
assign n_17015 =  x_1608 & ~n_1761;
assign n_17016 = ~x_1752 &  n_1761;
assign n_17017 = ~n_17015 & ~n_17016;
assign n_17018 =  x_1608 & ~n_17017;
assign n_17019 = ~x_1608 &  n_17017;
assign n_17020 = ~n_17018 & ~n_17019;
assign n_17021 =  x_1607 & ~n_1792;
assign n_17022 = ~x_1752 &  n_1792;
assign n_17023 = ~n_17021 & ~n_17022;
assign n_17024 =  x_1607 & ~n_17023;
assign n_17025 = ~x_1607 &  n_17023;
assign n_17026 = ~n_17024 & ~n_17025;
assign n_17027 =  x_1606 & ~n_1770;
assign n_17028 = ~x_1752 &  n_1770;
assign n_17029 = ~n_17027 & ~n_17028;
assign n_17030 =  x_1606 & ~n_17029;
assign n_17031 = ~x_1606 &  n_17029;
assign n_17032 = ~n_17030 & ~n_17031;
assign n_17033 =  x_1605 & ~n_1799;
assign n_17034 = ~x_1752 &  n_1799;
assign n_17035 = ~n_17033 & ~n_17034;
assign n_17036 =  x_1605 & ~n_17035;
assign n_17037 = ~x_1605 &  n_17035;
assign n_17038 = ~n_17036 & ~n_17037;
assign n_17039 =  x_1604 & ~n_1750;
assign n_17040 = ~x_1752 &  n_1750;
assign n_17041 = ~n_17039 & ~n_17040;
assign n_17042 =  x_1604 & ~n_17041;
assign n_17043 = ~x_1604 &  n_17041;
assign n_17044 = ~n_17042 & ~n_17043;
assign n_17045 =  x_1603 & ~n_1806;
assign n_17046 = ~x_1752 &  n_1806;
assign n_17047 = ~n_17045 & ~n_17046;
assign n_17048 =  x_1603 & ~n_17047;
assign n_17049 = ~x_1603 &  n_17047;
assign n_17050 = ~n_17048 & ~n_17049;
assign n_17051 =  x_1602 & ~n_1778;
assign n_17052 = ~x_1752 &  n_1778;
assign n_17053 = ~n_17051 & ~n_17052;
assign n_17054 =  x_1602 & ~n_17053;
assign n_17055 = ~x_1602 &  n_17053;
assign n_17056 = ~n_17054 & ~n_17055;
assign n_17057 =  x_1600 &  x_1601;
assign n_17058 = ~n_15969 & ~n_17057;
assign n_17059 = ~x_1747 &  n_3247;
assign n_17060 =  n_3274 &  n_17059;
assign n_17061 = ~x_1596 & ~n_3268;
assign n_17062 = ~n_3293 & ~n_17061;
assign n_17063 = ~n_17060 &  n_17062;
assign n_17064 = ~n_3267 & ~n_17063;
assign n_17065 =  x_1732 &  n_17064;
assign n_17066 = ~x_1598 &  n_17065;
assign n_17067 = ~x_1732 & ~n_17064;
assign n_17068 =  n_17067 & ~n_15971;
assign n_17069 = ~n_17066 & ~n_17068;
assign n_17070 = ~x_1600 &  n_17069;
assign n_17071 = ~n_17066 & ~n_17070;
assign n_17072 = ~n_17058 & ~n_17071;
assign n_17073 =  n_17058 &  n_17071;
assign n_17074 = ~n_17072 & ~n_17073;
assign n_17075 =  x_1601 &  n_17074;
assign n_17076 = ~x_1601 & ~n_17074;
assign n_17077 = ~n_17075 & ~n_17076;
assign n_17078 =  x_1600 & ~n_17069;
assign n_17079 = ~n_17078 & ~n_17070;
assign n_17080 =  x_1600 &  n_17079;
assign n_17081 = ~x_1600 & ~n_17079;
assign n_17082 = ~n_17080 & ~n_17081;
assign n_17083 =  n_15969 &  n_17067;
assign n_17084 =  n_17057 &  n_17065;
assign n_17085 = ~n_17083 & ~n_17084;
assign n_17086 = ~n_17069 & ~n_17085;
assign n_17087 = ~x_1599 &  n_17086;
assign n_17088 =  x_1599 & ~n_17086;
assign n_17089 = ~n_17087 & ~n_17088;
assign n_17090 =  x_1599 & ~n_17089;
assign n_17091 = ~x_1599 &  n_17089;
assign n_17092 = ~n_17090 & ~n_17091;
assign n_17093 =  x_1598 & ~n_17083;
assign n_17094 = ~x_1598 & ~n_17084;
assign n_17095 =  x_1599 & ~n_17094;
assign n_17096 = ~n_17093 & ~n_17095;
assign n_17097 =  x_1598 & ~n_17096;
assign n_17098 = ~x_1598 &  n_17096;
assign n_17099 = ~n_17097 & ~n_17098;
assign n_17100 = ~x_1597 & ~n_1715;
assign n_17101 =  n_1718 & ~n_17100;
assign n_17102 =  x_1597 &  n_17101;
assign n_17103 = ~x_1597 & ~n_17101;
assign n_17104 = ~n_17102 & ~n_17103;
assign n_17105 =  x_1596 & ~n_17064;
assign n_17106 = ~x_1596 &  n_17064;
assign n_17107 = ~n_17105 & ~n_17106;
assign n_17108 =  x_1596 &  n_3244;
assign n_17109 = ~n_3247 &  n_17108;
assign n_17110 = ~x_1594 & ~n_17109;
assign n_17111 =  x_1594 &  n_17109;
assign n_17112 = ~n_3266 & ~n_17111;
assign n_17113 = ~n_17110 &  n_17112;
assign n_17114 =  n_17113 &  n_17063;
assign n_17115 =  x_1595 &  n_17114;
assign n_17116 = ~x_1595 & ~n_17114;
assign n_17117 = ~n_17115 & ~n_17116;
assign n_17118 =  x_1594 &  n_17113;
assign n_17119 = ~x_1594 & ~n_17113;
assign n_17120 = ~n_17118 & ~n_17119;
assign n_17121 =  x_452 &  x_1593;
assign n_17122 =  n_17121 &  n_17111;
assign n_17123 = ~n_17121 & ~n_17111;
assign n_17124 = ~n_17122 & ~n_17123;
assign n_17125 =  x_1593 &  n_17124;
assign n_17126 = ~x_1593 & ~n_17124;
assign n_17127 = ~n_17125 & ~n_17126;
assign n_17128 =  x_1592 &  n_17122;
assign n_17129 =  x_452 &  x_1592;
assign n_17130 = ~n_17129 & ~n_17122;
assign n_17131 = ~n_17128 & ~n_17130;
assign n_17132 =  x_1592 &  n_17131;
assign n_17133 = ~x_1592 & ~n_17131;
assign n_17134 = ~n_17132 & ~n_17133;
assign n_17135 =  x_1563 &  n_17128;
assign n_17136 = ~x_1591 & ~n_17135;
assign n_17137 =  x_1591 &  n_17135;
assign n_17138 = ~n_3266 & ~n_17137;
assign n_17139 = ~n_17136 &  n_17138;
assign n_17140 =  x_1591 &  n_17139;
assign n_17141 = ~x_1591 & ~n_17139;
assign n_17142 = ~n_17140 & ~n_17141;
assign n_17143 = ~x_1590 & ~n_17137;
assign n_17144 =  x_1590 &  n_17137;
assign n_17145 = ~n_3266 & ~n_17144;
assign n_17146 = ~n_17143 &  n_17145;
assign n_17147 =  x_1590 &  n_17146;
assign n_17148 = ~x_1590 & ~n_17146;
assign n_17149 = ~n_17147 & ~n_17148;
assign n_17150 = ~x_1589 & ~n_17144;
assign n_17151 =  x_1589 &  n_17144;
assign n_17152 = ~n_3266 & ~n_17151;
assign n_17153 = ~n_17150 &  n_17152;
assign n_17154 =  x_1589 &  n_17153;
assign n_17155 = ~x_1589 & ~n_17153;
assign n_17156 = ~n_17154 & ~n_17155;
assign n_17157 = ~x_1588 & ~n_17151;
assign n_17158 =  x_1588 &  n_17151;
assign n_17159 = ~n_3266 & ~n_17158;
assign n_17160 = ~n_17157 &  n_17159;
assign n_17161 =  x_1588 &  n_17160;
assign n_17162 = ~x_1588 & ~n_17160;
assign n_17163 = ~n_17161 & ~n_17162;
assign n_17164 = ~x_1587 & ~n_17158;
assign n_17165 =  x_1587 &  n_17158;
assign n_17166 = ~n_3266 & ~n_17165;
assign n_17167 = ~n_17164 &  n_17166;
assign n_17168 =  x_1587 &  n_17167;
assign n_17169 = ~x_1587 & ~n_17167;
assign n_17170 = ~n_17168 & ~n_17169;
assign n_17171 = ~x_1586 & ~n_17165;
assign n_17172 =  x_1586 &  n_17165;
assign n_17173 = ~n_3266 & ~n_17172;
assign n_17174 = ~n_17171 &  n_17173;
assign n_17175 =  x_1586 &  n_17174;
assign n_17176 = ~x_1586 & ~n_17174;
assign n_17177 = ~n_17175 & ~n_17176;
assign n_17178 = ~x_1585 & ~n_17172;
assign n_17179 =  x_1585 &  n_17172;
assign n_17180 = ~n_3266 & ~n_17179;
assign n_17181 = ~n_17178 &  n_17180;
assign n_17182 =  x_1585 &  n_17181;
assign n_17183 = ~x_1585 & ~n_17181;
assign n_17184 = ~n_17182 & ~n_17183;
assign n_17185 = ~x_1584 & ~n_17179;
assign n_17186 =  x_1584 &  n_17179;
assign n_17187 = ~n_3266 & ~n_17186;
assign n_17188 = ~n_17185 &  n_17187;
assign n_17189 =  x_1584 &  n_17188;
assign n_17190 = ~x_1584 & ~n_17188;
assign n_17191 = ~n_17189 & ~n_17190;
assign n_17192 = ~x_1583 & ~n_17186;
assign n_17193 =  x_1583 &  n_17186;
assign n_17194 = ~n_3266 & ~n_17193;
assign n_17195 = ~n_17192 &  n_17194;
assign n_17196 =  x_1583 &  n_17195;
assign n_17197 = ~x_1583 & ~n_17195;
assign n_17198 = ~n_17196 & ~n_17197;
assign n_17199 = ~x_1582 & ~n_17193;
assign n_17200 =  x_1582 &  n_17193;
assign n_17201 = ~n_3266 & ~n_17200;
assign n_17202 = ~n_17199 &  n_17201;
assign n_17203 =  x_1582 &  n_17202;
assign n_17204 = ~x_1582 & ~n_17202;
assign n_17205 = ~n_17203 & ~n_17204;
assign n_17206 = ~x_1581 & ~n_17200;
assign n_17207 =  x_1581 &  n_17200;
assign n_17208 = ~n_3266 & ~n_17207;
assign n_17209 = ~n_17206 &  n_17208;
assign n_17210 =  x_1581 &  n_17209;
assign n_17211 = ~x_1581 & ~n_17209;
assign n_17212 = ~n_17210 & ~n_17211;
assign n_17213 = ~x_1580 & ~n_17207;
assign n_17214 =  x_1580 &  n_17207;
assign n_17215 = ~n_3266 & ~n_17214;
assign n_17216 = ~n_17213 &  n_17215;
assign n_17217 =  x_1580 &  n_17216;
assign n_17218 = ~x_1580 & ~n_17216;
assign n_17219 = ~n_17217 & ~n_17218;
assign n_17220 = ~x_1579 & ~n_17214;
assign n_17221 =  x_1579 &  n_17214;
assign n_17222 = ~n_3266 & ~n_17221;
assign n_17223 = ~n_17220 &  n_17222;
assign n_17224 =  x_1579 &  n_17223;
assign n_17225 = ~x_1579 & ~n_17223;
assign n_17226 = ~n_17224 & ~n_17225;
assign n_17227 = ~x_1578 & ~n_17221;
assign n_17228 =  x_1578 &  n_17221;
assign n_17229 = ~n_3266 & ~n_17228;
assign n_17230 = ~n_17227 &  n_17229;
assign n_17231 =  x_1578 &  n_17230;
assign n_17232 = ~x_1578 & ~n_17230;
assign n_17233 = ~n_17231 & ~n_17232;
assign n_17234 = ~x_1577 & ~n_17228;
assign n_17235 =  x_1577 &  n_17228;
assign n_17236 = ~n_3266 & ~n_17235;
assign n_17237 = ~n_17234 &  n_17236;
assign n_17238 =  x_1577 &  n_17237;
assign n_17239 = ~x_1577 & ~n_17237;
assign n_17240 = ~n_17238 & ~n_17239;
assign n_17241 = ~x_1576 & ~n_17235;
assign n_17242 =  x_1576 &  n_17235;
assign n_17243 = ~n_3266 & ~n_17242;
assign n_17244 = ~n_17241 &  n_17243;
assign n_17245 =  x_1576 &  n_17244;
assign n_17246 = ~x_1576 & ~n_17244;
assign n_17247 = ~n_17245 & ~n_17246;
assign n_17248 = ~x_1575 & ~n_17242;
assign n_17249 =  x_1575 &  n_17242;
assign n_17250 = ~n_3266 & ~n_17249;
assign n_17251 = ~n_17248 &  n_17250;
assign n_17252 =  x_1575 &  n_17251;
assign n_17253 = ~x_1575 & ~n_17251;
assign n_17254 = ~n_17252 & ~n_17253;
assign n_17255 = ~x_1574 & ~n_17249;
assign n_17256 =  x_1574 &  n_17249;
assign n_17257 = ~n_3266 & ~n_17256;
assign n_17258 = ~n_17255 &  n_17257;
assign n_17259 =  x_1574 &  n_17258;
assign n_17260 = ~x_1574 & ~n_17258;
assign n_17261 = ~n_17259 & ~n_17260;
assign n_17262 = ~x_1573 & ~n_17256;
assign n_17263 =  x_1573 &  n_17256;
assign n_17264 = ~n_3266 & ~n_17263;
assign n_17265 = ~n_17262 &  n_17264;
assign n_17266 =  x_1573 &  n_17265;
assign n_17267 = ~x_1573 & ~n_17265;
assign n_17268 = ~n_17266 & ~n_17267;
assign n_17269 = ~x_1572 & ~n_17263;
assign n_17270 =  x_1572 &  n_17263;
assign n_17271 = ~n_3266 & ~n_17270;
assign n_17272 = ~n_17269 &  n_17271;
assign n_17273 =  x_1572 &  n_17272;
assign n_17274 = ~x_1572 & ~n_17272;
assign n_17275 = ~n_17273 & ~n_17274;
assign n_17276 = ~x_1571 & ~n_17270;
assign n_17277 =  x_1571 &  n_17270;
assign n_17278 = ~n_3266 & ~n_17277;
assign n_17279 = ~n_17276 &  n_17278;
assign n_17280 =  x_1571 &  n_17279;
assign n_17281 = ~x_1571 & ~n_17279;
assign n_17282 = ~n_17280 & ~n_17281;
assign n_17283 = ~x_1570 & ~n_17277;
assign n_17284 =  x_1570 &  n_17277;
assign n_17285 = ~n_3266 & ~n_17284;
assign n_17286 = ~n_17283 &  n_17285;
assign n_17287 =  x_1570 &  n_17286;
assign n_17288 = ~x_1570 & ~n_17286;
assign n_17289 = ~n_17287 & ~n_17288;
assign n_17290 = ~x_1569 & ~n_17284;
assign n_17291 =  x_1569 &  n_17284;
assign n_17292 = ~n_3266 & ~n_17291;
assign n_17293 = ~n_17290 &  n_17292;
assign n_17294 =  x_1569 &  n_17293;
assign n_17295 = ~x_1569 & ~n_17293;
assign n_17296 = ~n_17294 & ~n_17295;
assign n_17297 = ~x_1568 & ~n_17291;
assign n_17298 =  x_1568 &  n_17291;
assign n_17299 = ~n_3266 & ~n_17298;
assign n_17300 = ~n_17297 &  n_17299;
assign n_17301 =  x_1568 &  n_17300;
assign n_17302 = ~x_1568 & ~n_17300;
assign n_17303 = ~n_17301 & ~n_17302;
assign n_17304 = ~x_1567 & ~n_17298;
assign n_17305 =  x_1567 &  n_17298;
assign n_17306 = ~n_3266 & ~n_17305;
assign n_17307 = ~n_17304 &  n_17306;
assign n_17308 =  x_1567 &  n_17307;
assign n_17309 = ~x_1567 & ~n_17307;
assign n_17310 = ~n_17308 & ~n_17309;
assign n_17311 = ~x_1566 & ~n_17305;
assign n_17312 =  x_1566 &  n_17305;
assign n_17313 = ~n_3266 & ~n_17312;
assign n_17314 = ~n_17311 &  n_17313;
assign n_17315 =  x_1566 &  n_17314;
assign n_17316 = ~x_1566 & ~n_17314;
assign n_17317 = ~n_17315 & ~n_17316;
assign n_17318 = ~x_1565 & ~n_17312;
assign n_17319 =  x_1565 &  n_17312;
assign n_17320 = ~n_3266 & ~n_17319;
assign n_17321 = ~n_17318 &  n_17320;
assign n_17322 =  x_1565 &  n_17321;
assign n_17323 = ~x_1565 & ~n_17321;
assign n_17324 = ~n_17322 & ~n_17323;
assign n_17325 =  x_1564 &  n_17319;
assign n_17326 = ~x_1564 & ~n_17319;
assign n_17327 = ~n_3266 & ~n_17326;
assign n_17328 = ~n_17325 &  n_17327;
assign n_17329 =  x_1564 &  n_17328;
assign n_17330 = ~x_1564 & ~n_17328;
assign n_17331 = ~n_17329 & ~n_17330;
assign n_17332 = ~x_1563 & ~n_17128;
assign n_17333 = ~n_3266 & ~n_17135;
assign n_17334 = ~n_17332 &  n_17333;
assign n_17335 =  x_1563 &  n_17334;
assign n_17336 = ~x_1563 & ~n_17334;
assign n_17337 = ~n_17335 & ~n_17336;
assign n_17338 = ~n_6109 & ~n_6112;
assign n_17339 =  x_1562 &  n_17338;
assign n_17340 = ~x_1562 & ~n_17338;
assign n_17341 = ~n_17339 & ~n_17340;
assign n_17342 =  x_1561 & ~n_5554;
assign n_17343 = ~x_1561 &  n_5554;
assign n_17344 = ~n_17342 & ~n_17343;
assign n_17345 =  x_1560 & ~n_5624;
assign n_17346 = ~x_1560 &  n_5624;
assign n_17347 = ~n_17345 & ~n_17346;
assign n_17348 =  x_1530 & ~n_4375;
assign n_17349 =  x_1529 &  n_17348;
assign n_17350 =  x_1528 &  n_17349;
assign n_17351 =  x_1527 &  n_17350;
assign n_17352 =  x_1526 &  n_17351;
assign n_17353 =  x_1525 &  n_17352;
assign n_17354 =  x_1524 &  n_17353;
assign n_17355 =  x_1523 &  n_17354;
assign n_17356 =  x_1522 &  n_17355;
assign n_17357 =  x_1521 &  n_17356;
assign n_17358 =  x_1520 &  n_17357;
assign n_17359 =  x_1519 &  n_17358;
assign n_17360 =  x_1518 &  n_17359;
assign n_17361 =  x_1517 &  n_17360;
assign n_17362 =  x_1516 &  n_17361;
assign n_17363 =  x_1515 &  n_17362;
assign n_17364 =  x_1514 &  n_17363;
assign n_17365 =  x_1513 &  n_17364;
assign n_17366 =  x_1512 &  n_17365;
assign n_17367 =  x_1511 &  n_17366;
assign n_17368 =  x_1510 &  n_17367;
assign n_17369 =  x_1509 &  n_17368;
assign n_17370 =  x_1508 &  n_17369;
assign n_17371 =  x_1507 &  n_17370;
assign n_17372 =  x_1506 &  n_17371;
assign n_17373 =  x_1505 &  n_17372;
assign n_17374 =  x_1504 &  n_17373;
assign n_17375 =  x_1503 &  n_17374;
assign n_17376 =  x_1502 &  n_17375;
assign n_17377 =  x_1501 &  n_17376;
assign n_17378 =  x_1558 &  n_17377;
assign n_17379 = ~x_1559 & ~n_17378;
assign n_17380 =  x_1559 &  n_17378;
assign n_17381 = ~n_17379 & ~n_17380;
assign n_17382 =  x_1559 &  n_17381;
assign n_17383 = ~x_1559 & ~n_17381;
assign n_17384 = ~n_17382 & ~n_17383;
assign n_17385 = ~x_1558 & ~n_17377;
assign n_17386 = ~n_17385 & ~n_17378;
assign n_17387 =  x_1558 &  n_17386;
assign n_17388 = ~x_1558 & ~n_17386;
assign n_17389 = ~n_17387 & ~n_17388;
assign n_17390 =  x_1557 & ~n_5549;
assign n_17391 = ~x_1557 &  n_5549;
assign n_17392 = ~n_17390 & ~n_17391;
assign n_17393 =  x_1556 & ~n_5684;
assign n_17394 = ~x_1556 &  n_5684;
assign n_17395 = ~n_17393 & ~n_17394;
assign n_17396 =  x_1555 & ~n_5696;
assign n_17397 = ~x_1555 &  n_5696;
assign n_17398 = ~n_17396 & ~n_17397;
assign n_17399 =  x_1554 & ~n_5564;
assign n_17400 = ~x_1554 &  n_5564;
assign n_17401 = ~n_17399 & ~n_17400;
assign n_17402 =  x_1553 & ~n_5579;
assign n_17403 = ~x_1553 &  n_5579;
assign n_17404 = ~n_17402 & ~n_17403;
assign n_17405 =  x_1552 & ~n_5584;
assign n_17406 = ~x_1552 &  n_5584;
assign n_17407 = ~n_17405 & ~n_17406;
assign n_17408 =  x_1551 & ~n_5604;
assign n_17409 = ~x_1551 &  n_5604;
assign n_17410 = ~n_17408 & ~n_17409;
assign n_17411 =  x_1550 & ~n_5599;
assign n_17412 = ~x_1550 &  n_5599;
assign n_17413 = ~n_17411 & ~n_17412;
assign n_17414 =  x_1549 & ~n_5649;
assign n_17415 = ~x_1549 &  n_5649;
assign n_17416 = ~n_17414 & ~n_17415;
assign n_17417 =  x_1548 & ~n_5691;
assign n_17418 = ~x_1548 &  n_5691;
assign n_17419 = ~n_17417 & ~n_17418;
assign n_17420 =  x_1547 & ~n_5644;
assign n_17421 = ~x_1547 &  n_5644;
assign n_17422 = ~n_17420 & ~n_17421;
assign n_17423 =  x_1546 & ~n_5634;
assign n_17424 = ~x_1546 &  n_5634;
assign n_17425 = ~n_17423 & ~n_17424;
assign n_17426 =  x_1545 & ~n_5629;
assign n_17427 = ~x_1545 &  n_5629;
assign n_17428 = ~n_17426 & ~n_17427;
assign n_17429 =  x_1544 & ~n_5659;
assign n_17430 = ~x_1544 &  n_5659;
assign n_17431 = ~n_17429 & ~n_17430;
assign n_17432 =  x_1543 & ~n_5674;
assign n_17433 = ~x_1543 &  n_5674;
assign n_17434 = ~n_17432 & ~n_17433;
assign n_17435 =  x_1542 & ~n_5679;
assign n_17436 = ~x_1542 &  n_5679;
assign n_17437 = ~n_17435 & ~n_17436;
assign n_17438 =  x_1541 & ~n_5654;
assign n_17439 = ~x_1541 &  n_5654;
assign n_17440 = ~n_17438 & ~n_17439;
assign n_17441 =  x_1540 & ~n_5639;
assign n_17442 = ~x_1540 &  n_5639;
assign n_17443 = ~n_17441 & ~n_17442;
assign n_17444 =  x_1539 & ~n_5664;
assign n_17445 = ~x_1539 &  n_5664;
assign n_17446 = ~n_17444 & ~n_17445;
assign n_17447 =  x_1538 & ~n_5669;
assign n_17448 = ~x_1538 &  n_5669;
assign n_17449 = ~n_17447 & ~n_17448;
assign n_17450 =  x_1537 & ~n_5614;
assign n_17451 = ~x_1537 &  n_5614;
assign n_17452 = ~n_17450 & ~n_17451;
assign n_17453 =  x_1536 & ~n_5594;
assign n_17454 = ~x_1536 &  n_5594;
assign n_17455 = ~n_17453 & ~n_17454;
assign n_17456 =  x_1535 & ~n_5609;
assign n_17457 = ~x_1535 &  n_5609;
assign n_17458 = ~n_17456 & ~n_17457;
assign n_17459 =  x_1534 & ~n_5619;
assign n_17460 = ~x_1534 &  n_5619;
assign n_17461 = ~n_17459 & ~n_17460;
assign n_17462 =  x_1533 & ~n_5589;
assign n_17463 = ~x_1533 &  n_5589;
assign n_17464 = ~n_17462 & ~n_17463;
assign n_17465 =  x_1532 & ~n_5574;
assign n_17466 = ~x_1532 &  n_5574;
assign n_17467 = ~n_17465 & ~n_17466;
assign n_17468 =  x_1531 & ~n_5569;
assign n_17469 = ~x_1531 &  n_5569;
assign n_17470 = ~n_17468 & ~n_17469;
assign n_17471 = ~x_1530 &  n_4375;
assign n_17472 = ~n_17348 & ~n_17471;
assign n_17473 =  x_1530 &  n_17472;
assign n_17474 = ~x_1530 & ~n_17472;
assign n_17475 = ~n_17473 & ~n_17474;
assign n_17476 = ~x_1529 & ~n_17348;
assign n_17477 = ~n_17349 & ~n_17476;
assign n_17478 =  x_1529 &  n_17477;
assign n_17479 = ~x_1529 & ~n_17477;
assign n_17480 = ~n_17478 & ~n_17479;
assign n_17481 = ~x_1528 & ~n_17349;
assign n_17482 = ~n_17350 & ~n_17481;
assign n_17483 =  x_1528 &  n_17482;
assign n_17484 = ~x_1528 & ~n_17482;
assign n_17485 = ~n_17483 & ~n_17484;
assign n_17486 = ~x_1527 & ~n_17350;
assign n_17487 = ~n_17351 & ~n_17486;
assign n_17488 =  x_1527 &  n_17487;
assign n_17489 = ~x_1527 & ~n_17487;
assign n_17490 = ~n_17488 & ~n_17489;
assign n_17491 = ~x_1526 & ~n_17351;
assign n_17492 = ~n_17352 & ~n_17491;
assign n_17493 =  x_1526 &  n_17492;
assign n_17494 = ~x_1526 & ~n_17492;
assign n_17495 = ~n_17493 & ~n_17494;
assign n_17496 = ~x_1525 & ~n_17352;
assign n_17497 = ~n_17353 & ~n_17496;
assign n_17498 =  x_1525 &  n_17497;
assign n_17499 = ~x_1525 & ~n_17497;
assign n_17500 = ~n_17498 & ~n_17499;
assign n_17501 = ~x_1524 & ~n_17353;
assign n_17502 = ~n_17354 & ~n_17501;
assign n_17503 =  x_1524 &  n_17502;
assign n_17504 = ~x_1524 & ~n_17502;
assign n_17505 = ~n_17503 & ~n_17504;
assign n_17506 = ~x_1523 & ~n_17354;
assign n_17507 = ~n_17355 & ~n_17506;
assign n_17508 =  x_1523 &  n_17507;
assign n_17509 = ~x_1523 & ~n_17507;
assign n_17510 = ~n_17508 & ~n_17509;
assign n_17511 = ~x_1522 & ~n_17355;
assign n_17512 = ~n_17356 & ~n_17511;
assign n_17513 =  x_1522 &  n_17512;
assign n_17514 = ~x_1522 & ~n_17512;
assign n_17515 = ~n_17513 & ~n_17514;
assign n_17516 = ~x_1521 & ~n_17356;
assign n_17517 = ~n_17357 & ~n_17516;
assign n_17518 =  x_1521 &  n_17517;
assign n_17519 = ~x_1521 & ~n_17517;
assign n_17520 = ~n_17518 & ~n_17519;
assign n_17521 = ~x_1520 & ~n_17357;
assign n_17522 = ~n_17358 & ~n_17521;
assign n_17523 =  x_1520 &  n_17522;
assign n_17524 = ~x_1520 & ~n_17522;
assign n_17525 = ~n_17523 & ~n_17524;
assign n_17526 = ~x_1519 & ~n_17358;
assign n_17527 = ~n_17359 & ~n_17526;
assign n_17528 =  x_1519 &  n_17527;
assign n_17529 = ~x_1519 & ~n_17527;
assign n_17530 = ~n_17528 & ~n_17529;
assign n_17531 = ~x_1518 & ~n_17359;
assign n_17532 = ~n_17360 & ~n_17531;
assign n_17533 =  x_1518 &  n_17532;
assign n_17534 = ~x_1518 & ~n_17532;
assign n_17535 = ~n_17533 & ~n_17534;
assign n_17536 = ~x_1517 & ~n_17360;
assign n_17537 = ~n_17361 & ~n_17536;
assign n_17538 =  x_1517 &  n_17537;
assign n_17539 = ~x_1517 & ~n_17537;
assign n_17540 = ~n_17538 & ~n_17539;
assign n_17541 = ~x_1516 & ~n_17361;
assign n_17542 = ~n_17362 & ~n_17541;
assign n_17543 =  x_1516 &  n_17542;
assign n_17544 = ~x_1516 & ~n_17542;
assign n_17545 = ~n_17543 & ~n_17544;
assign n_17546 = ~x_1515 & ~n_17362;
assign n_17547 = ~n_17363 & ~n_17546;
assign n_17548 =  x_1515 &  n_17547;
assign n_17549 = ~x_1515 & ~n_17547;
assign n_17550 = ~n_17548 & ~n_17549;
assign n_17551 = ~x_1514 & ~n_17363;
assign n_17552 = ~n_17364 & ~n_17551;
assign n_17553 =  x_1514 &  n_17552;
assign n_17554 = ~x_1514 & ~n_17552;
assign n_17555 = ~n_17553 & ~n_17554;
assign n_17556 = ~x_1513 & ~n_17364;
assign n_17557 = ~n_17365 & ~n_17556;
assign n_17558 =  x_1513 &  n_17557;
assign n_17559 = ~x_1513 & ~n_17557;
assign n_17560 = ~n_17558 & ~n_17559;
assign n_17561 = ~x_1512 & ~n_17365;
assign n_17562 = ~n_17366 & ~n_17561;
assign n_17563 =  x_1512 &  n_17562;
assign n_17564 = ~x_1512 & ~n_17562;
assign n_17565 = ~n_17563 & ~n_17564;
assign n_17566 = ~x_1511 & ~n_17366;
assign n_17567 = ~n_17367 & ~n_17566;
assign n_17568 =  x_1511 &  n_17567;
assign n_17569 = ~x_1511 & ~n_17567;
assign n_17570 = ~n_17568 & ~n_17569;
assign n_17571 = ~x_1510 & ~n_17367;
assign n_17572 = ~n_17368 & ~n_17571;
assign n_17573 =  x_1510 &  n_17572;
assign n_17574 = ~x_1510 & ~n_17572;
assign n_17575 = ~n_17573 & ~n_17574;
assign n_17576 = ~x_1509 & ~n_17368;
assign n_17577 = ~n_17369 & ~n_17576;
assign n_17578 =  x_1509 &  n_17577;
assign n_17579 = ~x_1509 & ~n_17577;
assign n_17580 = ~n_17578 & ~n_17579;
assign n_17581 = ~x_1508 & ~n_17369;
assign n_17582 = ~n_17370 & ~n_17581;
assign n_17583 =  x_1508 &  n_17582;
assign n_17584 = ~x_1508 & ~n_17582;
assign n_17585 = ~n_17583 & ~n_17584;
assign n_17586 = ~x_1507 & ~n_17370;
assign n_17587 = ~n_17371 & ~n_17586;
assign n_17588 =  x_1507 &  n_17587;
assign n_17589 = ~x_1507 & ~n_17587;
assign n_17590 = ~n_17588 & ~n_17589;
assign n_17591 = ~x_1506 & ~n_17371;
assign n_17592 = ~n_17372 & ~n_17591;
assign n_17593 =  x_1506 &  n_17592;
assign n_17594 = ~x_1506 & ~n_17592;
assign n_17595 = ~n_17593 & ~n_17594;
assign n_17596 = ~x_1505 & ~n_17372;
assign n_17597 = ~n_17373 & ~n_17596;
assign n_17598 =  x_1505 &  n_17597;
assign n_17599 = ~x_1505 & ~n_17597;
assign n_17600 = ~n_17598 & ~n_17599;
assign n_17601 = ~x_1504 & ~n_17373;
assign n_17602 = ~n_17374 & ~n_17601;
assign n_17603 =  x_1504 &  n_17602;
assign n_17604 = ~x_1504 & ~n_17602;
assign n_17605 = ~n_17603 & ~n_17604;
assign n_17606 = ~x_1503 & ~n_17374;
assign n_17607 = ~n_17375 & ~n_17606;
assign n_17608 =  x_1503 &  n_17607;
assign n_17609 = ~x_1503 & ~n_17607;
assign n_17610 = ~n_17608 & ~n_17609;
assign n_17611 = ~x_1502 & ~n_17375;
assign n_17612 = ~n_17376 & ~n_17611;
assign n_17613 =  x_1502 &  n_17612;
assign n_17614 = ~x_1502 & ~n_17612;
assign n_17615 = ~n_17613 & ~n_17614;
assign n_17616 = ~x_1501 & ~n_17376;
assign n_17617 = ~n_17616 & ~n_17377;
assign n_17618 =  x_1501 &  n_17617;
assign n_17619 = ~x_1501 & ~n_17617;
assign n_17620 = ~n_17618 & ~n_17619;
assign n_17621 =  x_1500 & ~n_5559;
assign n_17622 = ~x_1500 &  n_5559;
assign n_17623 = ~n_17621 & ~n_17622;
assign n_17624 =  x_1499 & ~n_4369;
assign n_17625 = ~x_1499 &  n_4369;
assign n_17626 = ~n_17624 & ~n_17625;
assign n_17627 =  n_6058 &  n_16353;
assign n_17628 = ~n_6058 & ~n_16353;
assign n_17629 = ~n_17627 & ~n_17628;
assign n_17630 =  x_1498 &  n_17629;
assign n_17631 = ~x_1498 & ~n_17629;
assign n_17632 = ~n_17630 & ~n_17631;
assign n_17633 = ~n_5993 & ~n_17627;
assign n_17634 =  x_1497 & ~n_17633;
assign n_17635 = ~x_1497 &  n_17633;
assign n_17636 = ~n_17634 & ~n_17635;
assign n_17637 =  x_1496 &  n_12453;
assign n_17638 = ~x_1496 & ~n_12453;
assign n_17639 = ~n_17637 & ~n_17638;
assign n_17640 =  x_1495 &  n_12452;
assign n_17641 = ~x_1495 & ~n_12452;
assign n_17642 = ~n_17640 & ~n_17641;
assign n_17643 =  x_1494 & ~n_1749;
assign n_17644 = ~n_1785 & ~n_17643;
assign n_17645 =  x_1494 & ~n_17644;
assign n_17646 = ~x_1494 &  n_17644;
assign n_17647 = ~n_17645 & ~n_17646;
assign n_17648 = ~x_1493 & ~n_1748;
assign n_17649 = ~n_1749 & ~n_17648;
assign n_17650 =  x_1493 &  n_17649;
assign n_17651 = ~x_1493 & ~n_17649;
assign n_17652 = ~n_17650 & ~n_17651;
assign n_17653 =  x_1492 & ~x_1771;
assign n_17654 = ~n_1759 & ~n_17653;
assign n_17655 =  x_1492 & ~n_17654;
assign n_17656 = ~x_1492 &  n_17654;
assign n_17657 = ~n_17655 & ~n_17656;
assign n_17658 = ~x_1752 &  n_3287;
assign n_17659 =  x_1491 & ~n_3267;
assign n_17660 = ~n_17658 & ~n_17659;
assign n_17661 =  x_1491 & ~n_17660;
assign n_17662 = ~x_1491 &  n_17660;
assign n_17663 = ~n_17661 & ~n_17662;
assign n_17664 = ~x_1490 & ~n_3240;
assign n_17665 = ~n_3241 & ~n_17664;
assign n_17666 =  x_1490 &  n_17665;
assign n_17667 = ~x_1490 & ~n_17665;
assign n_17668 = ~n_17666 & ~n_17667;
assign n_17669 = ~x_1746 & ~n_3293;
assign n_17670 =  x_1489 & ~n_17669;
assign n_17671 =  n_3243 &  n_3256;
assign n_17672 = ~n_17670 & ~n_17671;
assign n_17673 =  x_1489 & ~n_17672;
assign n_17674 = ~x_1489 &  n_17672;
assign n_17675 = ~n_17673 & ~n_17674;
assign n_17676 =  x_1758 &  n_12511;
assign n_17677 =  x_1488 &  n_17676;
assign n_17678 = ~x_1488 & ~n_17676;
assign n_17679 = ~n_17677 & ~n_17678;
assign n_17680 = ~x_1758 & ~n_12517;
assign n_17681 =  x_1487 &  n_17680;
assign n_17682 = ~x_1487 & ~n_17680;
assign n_17683 = ~n_17681 & ~n_17682;
assign n_17684 =  x_1486 &  n_17658;
assign n_17685 = ~x_1486 & ~n_17658;
assign n_17686 = ~n_17684 & ~n_17685;
assign n_17687 = ~x_1769 &  n_3244;
assign n_17688 = ~n_3243 &  n_17687;
assign n_17689 = ~x_1483 &  n_17688;
assign n_17690 = ~x_1484 &  n_17689;
assign n_17691 =  x_1485 & ~n_17690;
assign n_17692 =  n_17689 &  n_3246;
assign n_17693 =  x_1748 & ~n_17692;
assign n_17694 = ~n_17691 &  n_17693;
assign n_17695 = ~n_3266 & ~n_17694;
assign n_17696 =  x_1485 &  n_17695;
assign n_17697 = ~x_1485 & ~n_17695;
assign n_17698 = ~n_17696 & ~n_17697;
assign n_17699 =  x_1484 & ~n_17689;
assign n_17700 = ~n_17699 & ~n_17690;
assign n_17701 =  x_1748 & ~n_17700;
assign n_17702 =  x_1484 &  n_17701;
assign n_17703 = ~x_1484 & ~n_17701;
assign n_17704 = ~n_17702 & ~n_17703;
assign n_17705 =  x_1483 & ~n_17688;
assign n_17706 = ~n_17689 & ~n_17705;
assign n_17707 =  x_1748 & ~n_17706;
assign n_17708 =  x_1483 &  n_17707;
assign n_17709 = ~x_1483 & ~n_17707;
assign n_17710 = ~n_17708 & ~n_17709;
assign n_17711 = ~x_229 & ~n_510;
assign n_17712 =  n_1712 & ~n_17711;
assign n_17713 =  n_1713 & ~n_17712;
assign n_17714 =  x_1482 &  n_17713;
assign n_17715 = ~x_1482 & ~n_17713;
assign n_17716 = ~n_17714 & ~n_17715;
assign n_17717 =  n_1713 &  n_17711;
assign n_17718 =  x_1481 &  n_17717;
assign n_17719 = ~x_1481 & ~n_17717;
assign n_17720 = ~n_17718 & ~n_17719;
assign n_17721 =  x_1480 & ~n_1806;
assign n_17722 =  x_1750 &  n_1806;
assign n_17723 = ~n_17721 & ~n_17722;
assign n_17724 =  x_1480 & ~n_17723;
assign n_17725 = ~x_1480 &  n_17723;
assign n_17726 = ~n_17724 & ~n_17725;
assign n_17727 =  x_1479 & ~n_1799;
assign n_17728 =  x_1750 &  n_1799;
assign n_17729 = ~n_17727 & ~n_17728;
assign n_17730 =  x_1479 & ~n_17729;
assign n_17731 = ~x_1479 &  n_17729;
assign n_17732 = ~n_17730 & ~n_17731;
assign n_17733 =  x_1478 & ~n_1770;
assign n_17734 =  x_1750 &  n_1770;
assign n_17735 = ~n_17733 & ~n_17734;
assign n_17736 =  x_1478 & ~n_17735;
assign n_17737 = ~x_1478 &  n_17735;
assign n_17738 = ~n_17736 & ~n_17737;
assign n_17739 =  x_1477 & ~n_1778;
assign n_17740 =  x_1750 &  n_1778;
assign n_17741 = ~n_17739 & ~n_17740;
assign n_17742 =  x_1477 & ~n_17741;
assign n_17743 = ~x_1477 &  n_17741;
assign n_17744 = ~n_17742 & ~n_17743;
assign n_17745 =  x_1476 & ~n_1761;
assign n_17746 =  x_1750 &  n_1761;
assign n_17747 = ~n_17745 & ~n_17746;
assign n_17748 =  x_1476 & ~n_17747;
assign n_17749 = ~x_1476 &  n_17747;
assign n_17750 = ~n_17748 & ~n_17749;
assign n_17751 =  x_1475 & ~n_1750;
assign n_17752 =  x_1750 &  n_1750;
assign n_17753 = ~n_17751 & ~n_17752;
assign n_17754 =  x_1475 & ~n_17753;
assign n_17755 = ~x_1475 &  n_17753;
assign n_17756 = ~n_17754 & ~n_17755;
assign n_17757 =  x_1474 & ~n_1785;
assign n_17758 =  x_1750 &  n_1785;
assign n_17759 = ~n_17757 & ~n_17758;
assign n_17760 =  x_1474 & ~n_17759;
assign n_17761 = ~x_1474 &  n_17759;
assign n_17762 = ~n_17760 & ~n_17761;
assign n_17763 =  x_1473 & ~n_1792;
assign n_17764 =  x_1750 &  n_1792;
assign n_17765 = ~n_17763 & ~n_17764;
assign n_17766 =  x_1473 & ~n_17765;
assign n_17767 = ~x_1473 &  n_17765;
assign n_17768 = ~n_17766 & ~n_17767;
assign n_17769 =  x_1472 &  n_1717;
assign n_17770 = ~x_1472 & ~n_1717;
assign n_17771 = ~n_17769 & ~n_17770;
assign n_17772 =  x_1471 &  n_1723;
assign n_17773 = ~x_1471 & ~n_1723;
assign n_17774 = ~n_17772 & ~n_17773;
assign n_17775 = ~x_1470 & ~n_1716;
assign n_17776 = ~n_1723 & ~n_17775;
assign n_17777 =  x_1469 &  n_1715;
assign n_17778 = ~x_1469 & ~n_1715;
assign n_17779 = ~n_17777 & ~n_17778;
assign n_17780 =  x_1468 &  n_1713;
assign n_17781 = ~x_1468 & ~n_1713;
assign n_17782 = ~n_17780 & ~n_17781;
assign n_17783 = ~x_1467 & ~n_1739;
assign n_17784 = ~n_5985 & ~n_17783;
assign n_17785 = ~x_1466 & ~n_1522;
assign n_17786 = ~n_5726 & ~n_17785;
assign n_17787 = ~x_881 &  x_1732;
assign n_17788 = ~x_882 &  n_17787;
assign n_17789 = ~x_883 &  n_17788;
assign n_17790 =  x_1465 & ~n_17789;
assign n_17791 = ~x_1013 &  n_6109;
assign n_17792 = ~x_1012 & ~x_1562;
assign n_17793 =  x_1618 & ~x_1651;
assign n_17794 = ~n_17792 & ~n_17793;
assign n_17795 = ~n_17791 &  n_17794;
assign n_17796 = ~x_3229 & ~n_17795;
assign n_17797 = ~x_1812 &  x_3229;
assign n_17798 =  x_1732 & ~n_17797;
assign n_17799 = ~n_17796 &  n_17798;
assign n_17800 =  n_17789 &  n_17799;
assign n_17801 = ~n_17790 & ~n_17800;
assign n_17802 =  x_1465 & ~n_17801;
assign n_17803 = ~x_1465 &  n_17801;
assign n_17804 = ~n_17802 & ~n_17803;
assign n_17805 =  x_881 &  x_1732;
assign n_17806 = ~x_882 &  n_17805;
assign n_17807 = ~x_883 &  n_17806;
assign n_17808 =  x_1464 & ~n_17807;
assign n_17809 =  n_17807 &  n_17799;
assign n_17810 = ~n_17808 & ~n_17809;
assign n_17811 =  x_1464 & ~n_17810;
assign n_17812 = ~x_1464 &  n_17810;
assign n_17813 = ~n_17811 & ~n_17812;
assign n_17814 =  x_882 &  n_17787;
assign n_17815 = ~x_883 &  n_17814;
assign n_17816 =  x_1463 & ~n_17815;
assign n_17817 =  n_17815 &  n_17799;
assign n_17818 = ~n_17816 & ~n_17817;
assign n_17819 =  x_1463 & ~n_17818;
assign n_17820 = ~x_1463 &  n_17818;
assign n_17821 = ~n_17819 & ~n_17820;
assign n_17822 =  x_882 &  n_17805;
assign n_17823 = ~x_883 &  n_17822;
assign n_17824 =  x_1462 & ~n_17823;
assign n_17825 =  n_17823 &  n_17799;
assign n_17826 = ~n_17824 & ~n_17825;
assign n_17827 =  x_1462 & ~n_17826;
assign n_17828 = ~x_1462 &  n_17826;
assign n_17829 = ~n_17827 & ~n_17828;
assign n_17830 =  x_883 &  n_17788;
assign n_17831 =  x_1461 & ~n_17830;
assign n_17832 =  n_17830 &  n_17799;
assign n_17833 = ~n_17831 & ~n_17832;
assign n_17834 =  x_1461 & ~n_17833;
assign n_17835 = ~x_1461 &  n_17833;
assign n_17836 = ~n_17834 & ~n_17835;
assign n_17837 =  x_883 &  n_17806;
assign n_17838 =  x_1460 & ~n_17837;
assign n_17839 =  n_17837 &  n_17799;
assign n_17840 = ~n_17838 & ~n_17839;
assign n_17841 =  x_1460 & ~n_17840;
assign n_17842 = ~x_1460 &  n_17840;
assign n_17843 = ~n_17841 & ~n_17842;
assign n_17844 =  x_883 &  n_17814;
assign n_17845 =  x_1459 & ~n_17844;
assign n_17846 =  n_17844 &  n_17799;
assign n_17847 = ~n_17845 & ~n_17846;
assign n_17848 =  x_1459 & ~n_17847;
assign n_17849 = ~x_1459 &  n_17847;
assign n_17850 = ~n_17848 & ~n_17849;
assign n_17851 =  x_883 &  n_17822;
assign n_17852 =  x_1458 & ~n_17851;
assign n_17853 =  n_17851 &  n_17799;
assign n_17854 = ~n_17852 & ~n_17853;
assign n_17855 =  x_1458 & ~n_17854;
assign n_17856 = ~x_1458 &  n_17854;
assign n_17857 = ~n_17855 & ~n_17856;
assign n_17858 =  x_1457 & ~n_17789;
assign n_17859 = ~x_1011 &  n_6109;
assign n_17860 =  x_1618 & ~x_1650;
assign n_17861 = ~x_1010 & ~x_1562;
assign n_17862 = ~n_17860 & ~n_17861;
assign n_17863 = ~n_17859 &  n_17862;
assign n_17864 = ~x_3229 & ~n_17863;
assign n_17865 = ~x_1811 &  x_3229;
assign n_17866 =  x_1732 & ~n_17865;
assign n_17867 = ~n_17864 &  n_17866;
assign n_17868 =  n_17789 &  n_17867;
assign n_17869 = ~n_17858 & ~n_17868;
assign n_17870 =  x_1457 & ~n_17869;
assign n_17871 = ~x_1457 &  n_17869;
assign n_17872 = ~n_17870 & ~n_17871;
assign n_17873 =  x_1456 & ~n_17807;
assign n_17874 =  n_17807 &  n_17867;
assign n_17875 = ~n_17873 & ~n_17874;
assign n_17876 =  x_1456 & ~n_17875;
assign n_17877 = ~x_1456 &  n_17875;
assign n_17878 = ~n_17876 & ~n_17877;
assign n_17879 =  x_1455 & ~n_17815;
assign n_17880 =  n_17815 &  n_17867;
assign n_17881 = ~n_17879 & ~n_17880;
assign n_17882 =  x_1455 & ~n_17881;
assign n_17883 = ~x_1455 &  n_17881;
assign n_17884 = ~n_17882 & ~n_17883;
assign n_17885 =  x_1454 & ~n_17823;
assign n_17886 =  n_17823 &  n_17867;
assign n_17887 = ~n_17885 & ~n_17886;
assign n_17888 =  x_1454 & ~n_17887;
assign n_17889 = ~x_1454 &  n_17887;
assign n_17890 = ~n_17888 & ~n_17889;
assign n_17891 =  x_1453 & ~n_17830;
assign n_17892 =  n_17830 &  n_17867;
assign n_17893 = ~n_17891 & ~n_17892;
assign n_17894 =  x_1453 & ~n_17893;
assign n_17895 = ~x_1453 &  n_17893;
assign n_17896 = ~n_17894 & ~n_17895;
assign n_17897 =  x_1452 & ~n_17837;
assign n_17898 =  n_17837 &  n_17867;
assign n_17899 = ~n_17897 & ~n_17898;
assign n_17900 =  x_1452 & ~n_17899;
assign n_17901 = ~x_1452 &  n_17899;
assign n_17902 = ~n_17900 & ~n_17901;
assign n_17903 =  x_1451 & ~n_17844;
assign n_17904 =  n_17844 &  n_17867;
assign n_17905 = ~n_17903 & ~n_17904;
assign n_17906 =  x_1451 & ~n_17905;
assign n_17907 = ~x_1451 &  n_17905;
assign n_17908 = ~n_17906 & ~n_17907;
assign n_17909 =  x_1450 & ~n_17851;
assign n_17910 =  n_17851 &  n_17867;
assign n_17911 = ~n_17909 & ~n_17910;
assign n_17912 =  x_1450 & ~n_17911;
assign n_17913 = ~x_1450 &  n_17911;
assign n_17914 = ~n_17912 & ~n_17913;
assign n_17915 =  x_1449 & ~n_17789;
assign n_17916 = ~x_1009 &  n_6109;
assign n_17917 = ~x_1008 & ~x_1562;
assign n_17918 =  x_1618 & ~x_1649;
assign n_17919 = ~n_17917 & ~n_17918;
assign n_17920 = ~n_17916 &  n_17919;
assign n_17921 = ~x_3229 & ~n_17920;
assign n_17922 = ~x_1810 &  x_3229;
assign n_17923 =  x_1732 & ~n_17922;
assign n_17924 = ~n_17921 &  n_17923;
assign n_17925 =  n_17789 &  n_17924;
assign n_17926 = ~n_17915 & ~n_17925;
assign n_17927 =  x_1449 & ~n_17926;
assign n_17928 = ~x_1449 &  n_17926;
assign n_17929 = ~n_17927 & ~n_17928;
assign n_17930 =  x_1448 & ~n_17807;
assign n_17931 =  n_17807 &  n_17924;
assign n_17932 = ~n_17930 & ~n_17931;
assign n_17933 =  x_1448 & ~n_17932;
assign n_17934 = ~x_1448 &  n_17932;
assign n_17935 = ~n_17933 & ~n_17934;
assign n_17936 =  x_1447 & ~n_17815;
assign n_17937 =  n_17815 &  n_17924;
assign n_17938 = ~n_17936 & ~n_17937;
assign n_17939 =  x_1447 & ~n_17938;
assign n_17940 = ~x_1447 &  n_17938;
assign n_17941 = ~n_17939 & ~n_17940;
assign n_17942 =  x_1446 & ~n_17823;
assign n_17943 =  n_17823 &  n_17924;
assign n_17944 = ~n_17942 & ~n_17943;
assign n_17945 =  x_1446 & ~n_17944;
assign n_17946 = ~x_1446 &  n_17944;
assign n_17947 = ~n_17945 & ~n_17946;
assign n_17948 =  x_1445 & ~n_17830;
assign n_17949 =  n_17830 &  n_17924;
assign n_17950 = ~n_17948 & ~n_17949;
assign n_17951 =  x_1445 & ~n_17950;
assign n_17952 = ~x_1445 &  n_17950;
assign n_17953 = ~n_17951 & ~n_17952;
assign n_17954 =  x_1444 & ~n_17837;
assign n_17955 =  n_17837 &  n_17924;
assign n_17956 = ~n_17954 & ~n_17955;
assign n_17957 =  x_1444 & ~n_17956;
assign n_17958 = ~x_1444 &  n_17956;
assign n_17959 = ~n_17957 & ~n_17958;
assign n_17960 =  x_1443 & ~n_17844;
assign n_17961 =  n_17844 &  n_17924;
assign n_17962 = ~n_17960 & ~n_17961;
assign n_17963 =  x_1443 & ~n_17962;
assign n_17964 = ~x_1443 &  n_17962;
assign n_17965 = ~n_17963 & ~n_17964;
assign n_17966 =  x_1442 & ~n_17851;
assign n_17967 =  n_17851 &  n_17924;
assign n_17968 = ~n_17966 & ~n_17967;
assign n_17969 =  x_1442 & ~n_17968;
assign n_17970 = ~x_1442 &  n_17968;
assign n_17971 = ~n_17969 & ~n_17970;
assign n_17972 =  x_1441 & ~n_17789;
assign n_17973 = ~x_1007 &  n_6109;
assign n_17974 = ~x_1006 & ~x_1562;
assign n_17975 =  x_1618 & ~x_1648;
assign n_17976 = ~n_17974 & ~n_17975;
assign n_17977 = ~n_17973 &  n_17976;
assign n_17978 = ~x_3229 & ~n_17977;
assign n_17979 = ~x_1809 &  x_3229;
assign n_17980 =  x_1732 & ~n_17979;
assign n_17981 = ~n_17978 &  n_17980;
assign n_17982 =  n_17789 &  n_17981;
assign n_17983 = ~n_17972 & ~n_17982;
assign n_17984 =  x_1441 & ~n_17983;
assign n_17985 = ~x_1441 &  n_17983;
assign n_17986 = ~n_17984 & ~n_17985;
assign n_17987 =  x_1440 & ~n_17807;
assign n_17988 =  n_17807 &  n_17981;
assign n_17989 = ~n_17987 & ~n_17988;
assign n_17990 =  x_1440 & ~n_17989;
assign n_17991 = ~x_1440 &  n_17989;
assign n_17992 = ~n_17990 & ~n_17991;
assign n_17993 =  x_1439 & ~n_17815;
assign n_17994 =  n_17815 &  n_17981;
assign n_17995 = ~n_17993 & ~n_17994;
assign n_17996 =  x_1439 & ~n_17995;
assign n_17997 = ~x_1439 &  n_17995;
assign n_17998 = ~n_17996 & ~n_17997;
assign n_17999 =  x_1438 & ~n_17823;
assign n_18000 =  n_17823 &  n_17981;
assign n_18001 = ~n_17999 & ~n_18000;
assign n_18002 =  x_1438 & ~n_18001;
assign n_18003 = ~x_1438 &  n_18001;
assign n_18004 = ~n_18002 & ~n_18003;
assign n_18005 =  x_1437 & ~n_17830;
assign n_18006 =  n_17830 &  n_17981;
assign n_18007 = ~n_18005 & ~n_18006;
assign n_18008 =  x_1437 & ~n_18007;
assign n_18009 = ~x_1437 &  n_18007;
assign n_18010 = ~n_18008 & ~n_18009;
assign n_18011 =  x_1436 & ~n_17837;
assign n_18012 =  n_17837 &  n_17981;
assign n_18013 = ~n_18011 & ~n_18012;
assign n_18014 =  x_1436 & ~n_18013;
assign n_18015 = ~x_1436 &  n_18013;
assign n_18016 = ~n_18014 & ~n_18015;
assign n_18017 =  x_1435 & ~n_17844;
assign n_18018 =  n_17844 &  n_17981;
assign n_18019 = ~n_18017 & ~n_18018;
assign n_18020 =  x_1435 & ~n_18019;
assign n_18021 = ~x_1435 &  n_18019;
assign n_18022 = ~n_18020 & ~n_18021;
assign n_18023 =  x_1434 & ~n_17851;
assign n_18024 =  n_17851 &  n_17981;
assign n_18025 = ~n_18023 & ~n_18024;
assign n_18026 =  x_1434 & ~n_18025;
assign n_18027 = ~x_1434 &  n_18025;
assign n_18028 = ~n_18026 & ~n_18027;
assign n_18029 =  x_1433 & ~n_17789;
assign n_18030 = ~x_1005 &  n_6109;
assign n_18031 = ~x_1004 & ~x_1562;
assign n_18032 =  x_1618 & ~x_1647;
assign n_18033 = ~n_18031 & ~n_18032;
assign n_18034 = ~n_18030 &  n_18033;
assign n_18035 = ~x_3229 & ~n_18034;
assign n_18036 = ~x_1808 &  x_3229;
assign n_18037 =  x_1732 & ~n_18036;
assign n_18038 = ~n_18035 &  n_18037;
assign n_18039 =  n_17789 &  n_18038;
assign n_18040 = ~n_18029 & ~n_18039;
assign n_18041 =  x_1433 & ~n_18040;
assign n_18042 = ~x_1433 &  n_18040;
assign n_18043 = ~n_18041 & ~n_18042;
assign n_18044 =  x_1432 & ~n_17807;
assign n_18045 =  n_17807 &  n_18038;
assign n_18046 = ~n_18044 & ~n_18045;
assign n_18047 =  x_1432 & ~n_18046;
assign n_18048 = ~x_1432 &  n_18046;
assign n_18049 = ~n_18047 & ~n_18048;
assign n_18050 =  x_1431 & ~n_17815;
assign n_18051 =  n_17815 &  n_18038;
assign n_18052 = ~n_18050 & ~n_18051;
assign n_18053 =  x_1431 & ~n_18052;
assign n_18054 = ~x_1431 &  n_18052;
assign n_18055 = ~n_18053 & ~n_18054;
assign n_18056 =  x_1430 & ~n_17823;
assign n_18057 =  n_17823 &  n_18038;
assign n_18058 = ~n_18056 & ~n_18057;
assign n_18059 =  x_1430 & ~n_18058;
assign n_18060 = ~x_1430 &  n_18058;
assign n_18061 = ~n_18059 & ~n_18060;
assign n_18062 =  x_1429 & ~n_17830;
assign n_18063 =  n_17830 &  n_18038;
assign n_18064 = ~n_18062 & ~n_18063;
assign n_18065 =  x_1429 & ~n_18064;
assign n_18066 = ~x_1429 &  n_18064;
assign n_18067 = ~n_18065 & ~n_18066;
assign n_18068 =  x_1428 & ~n_17837;
assign n_18069 =  n_17837 &  n_18038;
assign n_18070 = ~n_18068 & ~n_18069;
assign n_18071 =  x_1428 & ~n_18070;
assign n_18072 = ~x_1428 &  n_18070;
assign n_18073 = ~n_18071 & ~n_18072;
assign n_18074 =  x_1427 & ~n_17844;
assign n_18075 =  n_17844 &  n_18038;
assign n_18076 = ~n_18074 & ~n_18075;
assign n_18077 =  x_1427 & ~n_18076;
assign n_18078 = ~x_1427 &  n_18076;
assign n_18079 = ~n_18077 & ~n_18078;
assign n_18080 =  x_1426 & ~n_17851;
assign n_18081 =  n_17851 &  n_18038;
assign n_18082 = ~n_18080 & ~n_18081;
assign n_18083 =  x_1426 & ~n_18082;
assign n_18084 = ~x_1426 &  n_18082;
assign n_18085 = ~n_18083 & ~n_18084;
assign n_18086 =  x_1425 & ~n_17789;
assign n_18087 = ~x_1003 &  n_6109;
assign n_18088 = ~x_1002 & ~x_1562;
assign n_18089 =  x_1618 & ~x_1646;
assign n_18090 = ~n_18088 & ~n_18089;
assign n_18091 = ~n_18087 &  n_18090;
assign n_18092 = ~x_3229 & ~n_18091;
assign n_18093 = ~x_1807 &  x_3229;
assign n_18094 =  x_1732 & ~n_18093;
assign n_18095 = ~n_18092 &  n_18094;
assign n_18096 =  n_17789 &  n_18095;
assign n_18097 = ~n_18086 & ~n_18096;
assign n_18098 =  x_1425 & ~n_18097;
assign n_18099 = ~x_1425 &  n_18097;
assign n_18100 = ~n_18098 & ~n_18099;
assign n_18101 =  x_1424 & ~n_17807;
assign n_18102 =  n_17807 &  n_18095;
assign n_18103 = ~n_18101 & ~n_18102;
assign n_18104 =  x_1424 & ~n_18103;
assign n_18105 = ~x_1424 &  n_18103;
assign n_18106 = ~n_18104 & ~n_18105;
assign n_18107 =  x_1423 & ~n_17815;
assign n_18108 =  n_17815 &  n_18095;
assign n_18109 = ~n_18107 & ~n_18108;
assign n_18110 =  x_1423 & ~n_18109;
assign n_18111 = ~x_1423 &  n_18109;
assign n_18112 = ~n_18110 & ~n_18111;
assign n_18113 =  x_1422 & ~n_17823;
assign n_18114 =  n_17823 &  n_18095;
assign n_18115 = ~n_18113 & ~n_18114;
assign n_18116 =  x_1422 & ~n_18115;
assign n_18117 = ~x_1422 &  n_18115;
assign n_18118 = ~n_18116 & ~n_18117;
assign n_18119 =  x_1421 & ~n_17830;
assign n_18120 =  n_17830 &  n_18095;
assign n_18121 = ~n_18119 & ~n_18120;
assign n_18122 =  x_1421 & ~n_18121;
assign n_18123 = ~x_1421 &  n_18121;
assign n_18124 = ~n_18122 & ~n_18123;
assign n_18125 =  x_1420 & ~n_17837;
assign n_18126 =  n_17837 &  n_18095;
assign n_18127 = ~n_18125 & ~n_18126;
assign n_18128 =  x_1420 & ~n_18127;
assign n_18129 = ~x_1420 &  n_18127;
assign n_18130 = ~n_18128 & ~n_18129;
assign n_18131 =  x_1419 & ~n_17844;
assign n_18132 =  n_17844 &  n_18095;
assign n_18133 = ~n_18131 & ~n_18132;
assign n_18134 =  x_1419 & ~n_18133;
assign n_18135 = ~x_1419 &  n_18133;
assign n_18136 = ~n_18134 & ~n_18135;
assign n_18137 =  x_1418 & ~n_17851;
assign n_18138 =  n_17851 &  n_18095;
assign n_18139 = ~n_18137 & ~n_18138;
assign n_18140 =  x_1418 & ~n_18139;
assign n_18141 = ~x_1418 &  n_18139;
assign n_18142 = ~n_18140 & ~n_18141;
assign n_18143 =  x_1417 & ~n_17789;
assign n_18144 = ~x_1001 &  n_6109;
assign n_18145 = ~x_1000 & ~x_1562;
assign n_18146 =  x_1618 & ~x_1645;
assign n_18147 = ~n_18145 & ~n_18146;
assign n_18148 = ~n_18144 &  n_18147;
assign n_18149 = ~x_3229 & ~n_18148;
assign n_18150 = ~x_1806 &  x_3229;
assign n_18151 =  x_1732 & ~n_18150;
assign n_18152 = ~n_18149 &  n_18151;
assign n_18153 =  n_17789 &  n_18152;
assign n_18154 = ~n_18143 & ~n_18153;
assign n_18155 =  x_1417 & ~n_18154;
assign n_18156 = ~x_1417 &  n_18154;
assign n_18157 = ~n_18155 & ~n_18156;
assign n_18158 =  x_1416 & ~n_17807;
assign n_18159 =  n_17807 &  n_18152;
assign n_18160 = ~n_18158 & ~n_18159;
assign n_18161 =  x_1416 & ~n_18160;
assign n_18162 = ~x_1416 &  n_18160;
assign n_18163 = ~n_18161 & ~n_18162;
assign n_18164 =  x_1415 & ~n_17815;
assign n_18165 =  n_17815 &  n_18152;
assign n_18166 = ~n_18164 & ~n_18165;
assign n_18167 =  x_1415 & ~n_18166;
assign n_18168 = ~x_1415 &  n_18166;
assign n_18169 = ~n_18167 & ~n_18168;
assign n_18170 =  x_1414 & ~n_17823;
assign n_18171 =  n_17823 &  n_18152;
assign n_18172 = ~n_18170 & ~n_18171;
assign n_18173 =  x_1414 & ~n_18172;
assign n_18174 = ~x_1414 &  n_18172;
assign n_18175 = ~n_18173 & ~n_18174;
assign n_18176 =  x_1413 & ~n_17830;
assign n_18177 =  n_17830 &  n_18152;
assign n_18178 = ~n_18176 & ~n_18177;
assign n_18179 =  x_1413 & ~n_18178;
assign n_18180 = ~x_1413 &  n_18178;
assign n_18181 = ~n_18179 & ~n_18180;
assign n_18182 =  x_1412 & ~n_17837;
assign n_18183 =  n_17837 &  n_18152;
assign n_18184 = ~n_18182 & ~n_18183;
assign n_18185 =  x_1412 & ~n_18184;
assign n_18186 = ~x_1412 &  n_18184;
assign n_18187 = ~n_18185 & ~n_18186;
assign n_18188 =  x_1411 & ~n_17844;
assign n_18189 =  n_17844 &  n_18152;
assign n_18190 = ~n_18188 & ~n_18189;
assign n_18191 =  x_1411 & ~n_18190;
assign n_18192 = ~x_1411 &  n_18190;
assign n_18193 = ~n_18191 & ~n_18192;
assign n_18194 =  x_1410 & ~n_17851;
assign n_18195 =  n_17851 &  n_18152;
assign n_18196 = ~n_18194 & ~n_18195;
assign n_18197 =  x_1410 & ~n_18196;
assign n_18198 = ~x_1410 &  n_18196;
assign n_18199 = ~n_18197 & ~n_18198;
assign n_18200 =  x_1409 & ~n_17789;
assign n_18201 = ~x_999 &  n_6109;
assign n_18202 =  x_1618 & ~x_1644;
assign n_18203 = ~x_998 & ~x_1562;
assign n_18204 = ~n_18202 & ~n_18203;
assign n_18205 = ~n_18201 &  n_18204;
assign n_18206 = ~x_3229 & ~n_18205;
assign n_18207 = ~x_1805 &  x_3229;
assign n_18208 =  x_1732 & ~n_18207;
assign n_18209 = ~n_18206 &  n_18208;
assign n_18210 =  n_17789 &  n_18209;
assign n_18211 = ~n_18200 & ~n_18210;
assign n_18212 =  x_1409 & ~n_18211;
assign n_18213 = ~x_1409 &  n_18211;
assign n_18214 = ~n_18212 & ~n_18213;
assign n_18215 =  x_1408 & ~n_17807;
assign n_18216 =  n_17807 &  n_18209;
assign n_18217 = ~n_18215 & ~n_18216;
assign n_18218 =  x_1408 & ~n_18217;
assign n_18219 = ~x_1408 &  n_18217;
assign n_18220 = ~n_18218 & ~n_18219;
assign n_18221 =  x_1407 & ~n_17815;
assign n_18222 =  n_17815 &  n_18209;
assign n_18223 = ~n_18221 & ~n_18222;
assign n_18224 =  x_1407 & ~n_18223;
assign n_18225 = ~x_1407 &  n_18223;
assign n_18226 = ~n_18224 & ~n_18225;
assign n_18227 =  x_1406 & ~n_17823;
assign n_18228 =  n_17823 &  n_18209;
assign n_18229 = ~n_18227 & ~n_18228;
assign n_18230 =  x_1406 & ~n_18229;
assign n_18231 = ~x_1406 &  n_18229;
assign n_18232 = ~n_18230 & ~n_18231;
assign n_18233 =  x_1405 & ~n_17830;
assign n_18234 =  n_17830 &  n_18209;
assign n_18235 = ~n_18233 & ~n_18234;
assign n_18236 =  x_1405 & ~n_18235;
assign n_18237 = ~x_1405 &  n_18235;
assign n_18238 = ~n_18236 & ~n_18237;
assign n_18239 =  x_1404 & ~n_17837;
assign n_18240 =  n_17837 &  n_18209;
assign n_18241 = ~n_18239 & ~n_18240;
assign n_18242 =  x_1404 & ~n_18241;
assign n_18243 = ~x_1404 &  n_18241;
assign n_18244 = ~n_18242 & ~n_18243;
assign n_18245 =  x_1403 & ~n_17844;
assign n_18246 =  n_17844 &  n_18209;
assign n_18247 = ~n_18245 & ~n_18246;
assign n_18248 =  x_1403 & ~n_18247;
assign n_18249 = ~x_1403 &  n_18247;
assign n_18250 = ~n_18248 & ~n_18249;
assign n_18251 =  x_1402 & ~n_17851;
assign n_18252 =  n_17851 &  n_18209;
assign n_18253 = ~n_18251 & ~n_18252;
assign n_18254 =  x_1402 & ~n_18253;
assign n_18255 = ~x_1402 &  n_18253;
assign n_18256 = ~n_18254 & ~n_18255;
assign n_18257 =  x_1401 & ~n_17789;
assign n_18258 = ~x_997 &  n_6109;
assign n_18259 =  x_1618 & ~x_1643;
assign n_18260 = ~x_996 & ~x_1562;
assign n_18261 = ~n_18259 & ~n_18260;
assign n_18262 = ~n_18258 &  n_18261;
assign n_18263 = ~x_3229 & ~n_18262;
assign n_18264 = ~x_1804 &  x_3229;
assign n_18265 =  x_1732 & ~n_18264;
assign n_18266 = ~n_18263 &  n_18265;
assign n_18267 =  n_17789 &  n_18266;
assign n_18268 = ~n_18257 & ~n_18267;
assign n_18269 =  x_1401 & ~n_18268;
assign n_18270 = ~x_1401 &  n_18268;
assign n_18271 = ~n_18269 & ~n_18270;
assign n_18272 =  x_1400 & ~n_17807;
assign n_18273 =  n_17807 &  n_18266;
assign n_18274 = ~n_18272 & ~n_18273;
assign n_18275 =  x_1400 & ~n_18274;
assign n_18276 = ~x_1400 &  n_18274;
assign n_18277 = ~n_18275 & ~n_18276;
assign n_18278 =  x_1399 & ~n_17815;
assign n_18279 =  n_17815 &  n_18266;
assign n_18280 = ~n_18278 & ~n_18279;
assign n_18281 =  x_1399 & ~n_18280;
assign n_18282 = ~x_1399 &  n_18280;
assign n_18283 = ~n_18281 & ~n_18282;
assign n_18284 =  x_1398 & ~n_17823;
assign n_18285 =  n_17823 &  n_18266;
assign n_18286 = ~n_18284 & ~n_18285;
assign n_18287 =  x_1398 & ~n_18286;
assign n_18288 = ~x_1398 &  n_18286;
assign n_18289 = ~n_18287 & ~n_18288;
assign n_18290 =  x_1397 & ~n_17830;
assign n_18291 =  n_17830 &  n_18266;
assign n_18292 = ~n_18290 & ~n_18291;
assign n_18293 =  x_1397 & ~n_18292;
assign n_18294 = ~x_1397 &  n_18292;
assign n_18295 = ~n_18293 & ~n_18294;
assign n_18296 =  x_1396 & ~n_17837;
assign n_18297 =  n_17837 &  n_18266;
assign n_18298 = ~n_18296 & ~n_18297;
assign n_18299 =  x_1396 & ~n_18298;
assign n_18300 = ~x_1396 &  n_18298;
assign n_18301 = ~n_18299 & ~n_18300;
assign n_18302 =  x_1395 & ~n_17844;
assign n_18303 =  n_17844 &  n_18266;
assign n_18304 = ~n_18302 & ~n_18303;
assign n_18305 =  x_1395 & ~n_18304;
assign n_18306 = ~x_1395 &  n_18304;
assign n_18307 = ~n_18305 & ~n_18306;
assign n_18308 =  x_1394 & ~n_17851;
assign n_18309 =  n_17851 &  n_18266;
assign n_18310 = ~n_18308 & ~n_18309;
assign n_18311 =  x_1394 & ~n_18310;
assign n_18312 = ~x_1394 &  n_18310;
assign n_18313 = ~n_18311 & ~n_18312;
assign n_18314 =  x_1393 & ~n_17789;
assign n_18315 = ~x_995 &  n_6109;
assign n_18316 =  x_1618 & ~x_1642;
assign n_18317 = ~x_994 & ~x_1562;
assign n_18318 = ~n_18316 & ~n_18317;
assign n_18319 = ~n_18315 &  n_18318;
assign n_18320 = ~x_3229 & ~n_18319;
assign n_18321 = ~x_1803 &  x_3229;
assign n_18322 =  x_1732 & ~n_18321;
assign n_18323 = ~n_18320 &  n_18322;
assign n_18324 =  n_17789 &  n_18323;
assign n_18325 = ~n_18314 & ~n_18324;
assign n_18326 =  x_1393 & ~n_18325;
assign n_18327 = ~x_1393 &  n_18325;
assign n_18328 = ~n_18326 & ~n_18327;
assign n_18329 =  x_1392 & ~n_17807;
assign n_18330 =  n_17807 &  n_18323;
assign n_18331 = ~n_18329 & ~n_18330;
assign n_18332 =  x_1392 & ~n_18331;
assign n_18333 = ~x_1392 &  n_18331;
assign n_18334 = ~n_18332 & ~n_18333;
assign n_18335 =  x_1391 & ~n_17815;
assign n_18336 =  n_17815 &  n_18323;
assign n_18337 = ~n_18335 & ~n_18336;
assign n_18338 =  x_1391 & ~n_18337;
assign n_18339 = ~x_1391 &  n_18337;
assign n_18340 = ~n_18338 & ~n_18339;
assign n_18341 =  x_1390 & ~n_17823;
assign n_18342 =  n_17823 &  n_18323;
assign n_18343 = ~n_18341 & ~n_18342;
assign n_18344 =  x_1390 & ~n_18343;
assign n_18345 = ~x_1390 &  n_18343;
assign n_18346 = ~n_18344 & ~n_18345;
assign n_18347 =  x_1389 & ~n_17830;
assign n_18348 =  n_17830 &  n_18323;
assign n_18349 = ~n_18347 & ~n_18348;
assign n_18350 =  x_1389 & ~n_18349;
assign n_18351 = ~x_1389 &  n_18349;
assign n_18352 = ~n_18350 & ~n_18351;
assign n_18353 =  x_1388 & ~n_17837;
assign n_18354 =  n_17837 &  n_18323;
assign n_18355 = ~n_18353 & ~n_18354;
assign n_18356 =  x_1388 & ~n_18355;
assign n_18357 = ~x_1388 &  n_18355;
assign n_18358 = ~n_18356 & ~n_18357;
assign n_18359 =  x_1387 & ~n_17844;
assign n_18360 =  n_17844 &  n_18323;
assign n_18361 = ~n_18359 & ~n_18360;
assign n_18362 =  x_1387 & ~n_18361;
assign n_18363 = ~x_1387 &  n_18361;
assign n_18364 = ~n_18362 & ~n_18363;
assign n_18365 =  x_1386 & ~n_17851;
assign n_18366 =  n_17851 &  n_18323;
assign n_18367 = ~n_18365 & ~n_18366;
assign n_18368 =  x_1386 & ~n_18367;
assign n_18369 = ~x_1386 &  n_18367;
assign n_18370 = ~n_18368 & ~n_18369;
assign n_18371 =  x_1385 & ~n_17789;
assign n_18372 = ~x_993 &  n_6109;
assign n_18373 = ~x_992 & ~x_1562;
assign n_18374 =  x_1618 & ~x_1641;
assign n_18375 = ~n_18373 & ~n_18374;
assign n_18376 = ~n_18372 &  n_18375;
assign n_18377 = ~x_3229 & ~n_18376;
assign n_18378 = ~x_1802 &  x_3229;
assign n_18379 =  x_1732 & ~n_18378;
assign n_18380 = ~n_18377 &  n_18379;
assign n_18381 =  n_17789 &  n_18380;
assign n_18382 = ~n_18371 & ~n_18381;
assign n_18383 =  x_1385 & ~n_18382;
assign n_18384 = ~x_1385 &  n_18382;
assign n_18385 = ~n_18383 & ~n_18384;
assign n_18386 =  x_1384 & ~n_17807;
assign n_18387 =  n_17807 &  n_18380;
assign n_18388 = ~n_18386 & ~n_18387;
assign n_18389 =  x_1384 & ~n_18388;
assign n_18390 = ~x_1384 &  n_18388;
assign n_18391 = ~n_18389 & ~n_18390;
assign n_18392 =  x_1383 & ~n_17815;
assign n_18393 =  n_17815 &  n_18380;
assign n_18394 = ~n_18392 & ~n_18393;
assign n_18395 =  x_1383 & ~n_18394;
assign n_18396 = ~x_1383 &  n_18394;
assign n_18397 = ~n_18395 & ~n_18396;
assign n_18398 =  x_1382 & ~n_17823;
assign n_18399 =  n_17823 &  n_18380;
assign n_18400 = ~n_18398 & ~n_18399;
assign n_18401 =  x_1382 & ~n_18400;
assign n_18402 = ~x_1382 &  n_18400;
assign n_18403 = ~n_18401 & ~n_18402;
assign n_18404 =  x_1381 & ~n_17830;
assign n_18405 =  n_17830 &  n_18380;
assign n_18406 = ~n_18404 & ~n_18405;
assign n_18407 =  x_1381 & ~n_18406;
assign n_18408 = ~x_1381 &  n_18406;
assign n_18409 = ~n_18407 & ~n_18408;
assign n_18410 =  x_1380 & ~n_17837;
assign n_18411 =  n_17837 &  n_18380;
assign n_18412 = ~n_18410 & ~n_18411;
assign n_18413 =  x_1380 & ~n_18412;
assign n_18414 = ~x_1380 &  n_18412;
assign n_18415 = ~n_18413 & ~n_18414;
assign n_18416 =  x_1379 & ~n_17844;
assign n_18417 =  n_17844 &  n_18380;
assign n_18418 = ~n_18416 & ~n_18417;
assign n_18419 =  x_1379 & ~n_18418;
assign n_18420 = ~x_1379 &  n_18418;
assign n_18421 = ~n_18419 & ~n_18420;
assign n_18422 =  x_1378 & ~n_17851;
assign n_18423 =  n_17851 &  n_18380;
assign n_18424 = ~n_18422 & ~n_18423;
assign n_18425 =  x_1378 & ~n_18424;
assign n_18426 = ~x_1378 &  n_18424;
assign n_18427 = ~n_18425 & ~n_18426;
assign n_18428 =  x_1377 & ~n_17789;
assign n_18429 = ~x_991 &  n_6109;
assign n_18430 = ~x_990 & ~x_1562;
assign n_18431 =  x_1618 & ~x_1640;
assign n_18432 = ~n_18430 & ~n_18431;
assign n_18433 = ~n_18429 &  n_18432;
assign n_18434 = ~x_3229 & ~n_18433;
assign n_18435 = ~x_1801 &  x_3229;
assign n_18436 =  x_1732 & ~n_18435;
assign n_18437 = ~n_18434 &  n_18436;
assign n_18438 =  n_17789 &  n_18437;
assign n_18439 = ~n_18428 & ~n_18438;
assign n_18440 =  x_1377 & ~n_18439;
assign n_18441 = ~x_1377 &  n_18439;
assign n_18442 = ~n_18440 & ~n_18441;
assign n_18443 =  x_1376 & ~n_17807;
assign n_18444 =  n_17807 &  n_18437;
assign n_18445 = ~n_18443 & ~n_18444;
assign n_18446 =  x_1376 & ~n_18445;
assign n_18447 = ~x_1376 &  n_18445;
assign n_18448 = ~n_18446 & ~n_18447;
assign n_18449 =  x_1375 & ~n_17815;
assign n_18450 =  n_17815 &  n_18437;
assign n_18451 = ~n_18449 & ~n_18450;
assign n_18452 =  x_1375 & ~n_18451;
assign n_18453 = ~x_1375 &  n_18451;
assign n_18454 = ~n_18452 & ~n_18453;
assign n_18455 =  x_1374 & ~n_17823;
assign n_18456 =  n_17823 &  n_18437;
assign n_18457 = ~n_18455 & ~n_18456;
assign n_18458 =  x_1374 & ~n_18457;
assign n_18459 = ~x_1374 &  n_18457;
assign n_18460 = ~n_18458 & ~n_18459;
assign n_18461 =  x_1373 & ~n_17830;
assign n_18462 =  n_17830 &  n_18437;
assign n_18463 = ~n_18461 & ~n_18462;
assign n_18464 =  x_1373 & ~n_18463;
assign n_18465 = ~x_1373 &  n_18463;
assign n_18466 = ~n_18464 & ~n_18465;
assign n_18467 =  x_1372 & ~n_17837;
assign n_18468 =  n_17837 &  n_18437;
assign n_18469 = ~n_18467 & ~n_18468;
assign n_18470 =  x_1372 & ~n_18469;
assign n_18471 = ~x_1372 &  n_18469;
assign n_18472 = ~n_18470 & ~n_18471;
assign n_18473 =  x_1371 & ~n_17844;
assign n_18474 =  n_17844 &  n_18437;
assign n_18475 = ~n_18473 & ~n_18474;
assign n_18476 =  x_1371 & ~n_18475;
assign n_18477 = ~x_1371 &  n_18475;
assign n_18478 = ~n_18476 & ~n_18477;
assign n_18479 =  x_1370 & ~n_17851;
assign n_18480 =  n_17851 &  n_18437;
assign n_18481 = ~n_18479 & ~n_18480;
assign n_18482 =  x_1370 & ~n_18481;
assign n_18483 = ~x_1370 &  n_18481;
assign n_18484 = ~n_18482 & ~n_18483;
assign n_18485 =  x_1369 & ~n_17789;
assign n_18486 = ~x_989 &  n_6109;
assign n_18487 = ~x_988 & ~x_1562;
assign n_18488 =  x_1618 & ~x_1639;
assign n_18489 = ~n_18487 & ~n_18488;
assign n_18490 = ~n_18486 &  n_18489;
assign n_18491 = ~x_3229 & ~n_18490;
assign n_18492 = ~x_1800 &  x_3229;
assign n_18493 =  x_1732 & ~n_18492;
assign n_18494 = ~n_18491 &  n_18493;
assign n_18495 =  n_17789 &  n_18494;
assign n_18496 = ~n_18485 & ~n_18495;
assign n_18497 =  x_1369 & ~n_18496;
assign n_18498 = ~x_1369 &  n_18496;
assign n_18499 = ~n_18497 & ~n_18498;
assign n_18500 =  x_1368 & ~n_17807;
assign n_18501 =  n_17807 &  n_18494;
assign n_18502 = ~n_18500 & ~n_18501;
assign n_18503 =  x_1368 & ~n_18502;
assign n_18504 = ~x_1368 &  n_18502;
assign n_18505 = ~n_18503 & ~n_18504;
assign n_18506 =  x_1367 & ~n_17815;
assign n_18507 =  n_17815 &  n_18494;
assign n_18508 = ~n_18506 & ~n_18507;
assign n_18509 =  x_1367 & ~n_18508;
assign n_18510 = ~x_1367 &  n_18508;
assign n_18511 = ~n_18509 & ~n_18510;
assign n_18512 =  x_1366 & ~n_17823;
assign n_18513 =  n_17823 &  n_18494;
assign n_18514 = ~n_18512 & ~n_18513;
assign n_18515 =  x_1366 & ~n_18514;
assign n_18516 = ~x_1366 &  n_18514;
assign n_18517 = ~n_18515 & ~n_18516;
assign n_18518 =  x_1365 & ~n_17830;
assign n_18519 =  n_17830 &  n_18494;
assign n_18520 = ~n_18518 & ~n_18519;
assign n_18521 =  x_1365 & ~n_18520;
assign n_18522 = ~x_1365 &  n_18520;
assign n_18523 = ~n_18521 & ~n_18522;
assign n_18524 =  x_1364 & ~n_17837;
assign n_18525 =  n_17837 &  n_18494;
assign n_18526 = ~n_18524 & ~n_18525;
assign n_18527 =  x_1364 & ~n_18526;
assign n_18528 = ~x_1364 &  n_18526;
assign n_18529 = ~n_18527 & ~n_18528;
assign n_18530 =  x_1363 & ~n_17844;
assign n_18531 =  n_17844 &  n_18494;
assign n_18532 = ~n_18530 & ~n_18531;
assign n_18533 =  x_1363 & ~n_18532;
assign n_18534 = ~x_1363 &  n_18532;
assign n_18535 = ~n_18533 & ~n_18534;
assign n_18536 =  x_1362 & ~n_17851;
assign n_18537 =  n_17851 &  n_18494;
assign n_18538 = ~n_18536 & ~n_18537;
assign n_18539 =  x_1362 & ~n_18538;
assign n_18540 = ~x_1362 &  n_18538;
assign n_18541 = ~n_18539 & ~n_18540;
assign n_18542 =  x_1361 & ~n_17789;
assign n_18543 = ~x_987 &  n_6109;
assign n_18544 = ~x_986 & ~x_1562;
assign n_18545 =  x_1618 & ~x_1638;
assign n_18546 = ~n_18544 & ~n_18545;
assign n_18547 = ~n_18543 &  n_18546;
assign n_18548 = ~x_3229 & ~n_18547;
assign n_18549 = ~x_1799 &  x_3229;
assign n_18550 =  x_1732 & ~n_18549;
assign n_18551 = ~n_18548 &  n_18550;
assign n_18552 =  n_17789 &  n_18551;
assign n_18553 = ~n_18542 & ~n_18552;
assign n_18554 =  x_1361 & ~n_18553;
assign n_18555 = ~x_1361 &  n_18553;
assign n_18556 = ~n_18554 & ~n_18555;
assign n_18557 =  x_1360 & ~n_17807;
assign n_18558 =  n_17807 &  n_18551;
assign n_18559 = ~n_18557 & ~n_18558;
assign n_18560 =  x_1360 & ~n_18559;
assign n_18561 = ~x_1360 &  n_18559;
assign n_18562 = ~n_18560 & ~n_18561;
assign n_18563 =  x_1359 & ~n_17815;
assign n_18564 =  n_17815 &  n_18551;
assign n_18565 = ~n_18563 & ~n_18564;
assign n_18566 =  x_1359 & ~n_18565;
assign n_18567 = ~x_1359 &  n_18565;
assign n_18568 = ~n_18566 & ~n_18567;
assign n_18569 =  x_1358 & ~n_17823;
assign n_18570 =  n_17823 &  n_18551;
assign n_18571 = ~n_18569 & ~n_18570;
assign n_18572 =  x_1358 & ~n_18571;
assign n_18573 = ~x_1358 &  n_18571;
assign n_18574 = ~n_18572 & ~n_18573;
assign n_18575 =  x_1357 & ~n_17830;
assign n_18576 =  n_17830 &  n_18551;
assign n_18577 = ~n_18575 & ~n_18576;
assign n_18578 =  x_1357 & ~n_18577;
assign n_18579 = ~x_1357 &  n_18577;
assign n_18580 = ~n_18578 & ~n_18579;
assign n_18581 =  x_1356 & ~n_17837;
assign n_18582 =  n_17837 &  n_18551;
assign n_18583 = ~n_18581 & ~n_18582;
assign n_18584 =  x_1356 & ~n_18583;
assign n_18585 = ~x_1356 &  n_18583;
assign n_18586 = ~n_18584 & ~n_18585;
assign n_18587 =  x_1355 & ~n_17844;
assign n_18588 =  n_17844 &  n_18551;
assign n_18589 = ~n_18587 & ~n_18588;
assign n_18590 =  x_1355 & ~n_18589;
assign n_18591 = ~x_1355 &  n_18589;
assign n_18592 = ~n_18590 & ~n_18591;
assign n_18593 =  x_1354 & ~n_17851;
assign n_18594 =  n_17851 &  n_18551;
assign n_18595 = ~n_18593 & ~n_18594;
assign n_18596 =  x_1354 & ~n_18595;
assign n_18597 = ~x_1354 &  n_18595;
assign n_18598 = ~n_18596 & ~n_18597;
assign n_18599 =  x_1353 & ~n_17789;
assign n_18600 = ~x_985 &  n_6109;
assign n_18601 = ~x_984 & ~x_1562;
assign n_18602 =  x_1618 & ~x_1637;
assign n_18603 = ~n_18601 & ~n_18602;
assign n_18604 = ~n_18600 &  n_18603;
assign n_18605 = ~x_3229 & ~n_18604;
assign n_18606 = ~x_1798 &  x_3229;
assign n_18607 =  x_1732 & ~n_18606;
assign n_18608 = ~n_18605 &  n_18607;
assign n_18609 =  n_17789 &  n_18608;
assign n_18610 = ~n_18599 & ~n_18609;
assign n_18611 =  x_1353 & ~n_18610;
assign n_18612 = ~x_1353 &  n_18610;
assign n_18613 = ~n_18611 & ~n_18612;
assign n_18614 =  x_1352 & ~n_17807;
assign n_18615 =  n_17807 &  n_18608;
assign n_18616 = ~n_18614 & ~n_18615;
assign n_18617 =  x_1352 & ~n_18616;
assign n_18618 = ~x_1352 &  n_18616;
assign n_18619 = ~n_18617 & ~n_18618;
assign n_18620 =  x_1351 & ~n_17815;
assign n_18621 =  n_17815 &  n_18608;
assign n_18622 = ~n_18620 & ~n_18621;
assign n_18623 =  x_1351 & ~n_18622;
assign n_18624 = ~x_1351 &  n_18622;
assign n_18625 = ~n_18623 & ~n_18624;
assign n_18626 =  x_1350 & ~n_17823;
assign n_18627 =  n_17823 &  n_18608;
assign n_18628 = ~n_18626 & ~n_18627;
assign n_18629 =  x_1350 & ~n_18628;
assign n_18630 = ~x_1350 &  n_18628;
assign n_18631 = ~n_18629 & ~n_18630;
assign n_18632 =  x_1349 & ~n_17830;
assign n_18633 =  n_17830 &  n_18608;
assign n_18634 = ~n_18632 & ~n_18633;
assign n_18635 =  x_1349 & ~n_18634;
assign n_18636 = ~x_1349 &  n_18634;
assign n_18637 = ~n_18635 & ~n_18636;
assign n_18638 =  x_1348 & ~n_17837;
assign n_18639 =  n_17837 &  n_18608;
assign n_18640 = ~n_18638 & ~n_18639;
assign n_18641 =  x_1348 & ~n_18640;
assign n_18642 = ~x_1348 &  n_18640;
assign n_18643 = ~n_18641 & ~n_18642;
assign n_18644 =  x_1347 & ~n_17844;
assign n_18645 =  n_17844 &  n_18608;
assign n_18646 = ~n_18644 & ~n_18645;
assign n_18647 =  x_1347 & ~n_18646;
assign n_18648 = ~x_1347 &  n_18646;
assign n_18649 = ~n_18647 & ~n_18648;
assign n_18650 =  x_1346 & ~n_17851;
assign n_18651 =  n_17851 &  n_18608;
assign n_18652 = ~n_18650 & ~n_18651;
assign n_18653 =  x_1346 & ~n_18652;
assign n_18654 = ~x_1346 &  n_18652;
assign n_18655 = ~n_18653 & ~n_18654;
assign n_18656 =  x_1345 & ~n_17789;
assign n_18657 = ~x_983 &  n_6109;
assign n_18658 =  x_1618 & ~x_1636;
assign n_18659 = ~x_982 & ~x_1562;
assign n_18660 = ~n_18658 & ~n_18659;
assign n_18661 = ~n_18657 &  n_18660;
assign n_18662 = ~x_3229 & ~n_18661;
assign n_18663 = ~x_1797 &  x_3229;
assign n_18664 =  x_1732 & ~n_18663;
assign n_18665 = ~n_18662 &  n_18664;
assign n_18666 =  n_17789 &  n_18665;
assign n_18667 = ~n_18656 & ~n_18666;
assign n_18668 =  x_1345 & ~n_18667;
assign n_18669 = ~x_1345 &  n_18667;
assign n_18670 = ~n_18668 & ~n_18669;
assign n_18671 =  x_1344 & ~n_17807;
assign n_18672 =  n_17807 &  n_18665;
assign n_18673 = ~n_18671 & ~n_18672;
assign n_18674 =  x_1344 & ~n_18673;
assign n_18675 = ~x_1344 &  n_18673;
assign n_18676 = ~n_18674 & ~n_18675;
assign n_18677 =  x_1343 & ~n_17815;
assign n_18678 =  n_17815 &  n_18665;
assign n_18679 = ~n_18677 & ~n_18678;
assign n_18680 =  x_1343 & ~n_18679;
assign n_18681 = ~x_1343 &  n_18679;
assign n_18682 = ~n_18680 & ~n_18681;
assign n_18683 =  x_1342 & ~n_17823;
assign n_18684 =  n_17823 &  n_18665;
assign n_18685 = ~n_18683 & ~n_18684;
assign n_18686 =  x_1342 & ~n_18685;
assign n_18687 = ~x_1342 &  n_18685;
assign n_18688 = ~n_18686 & ~n_18687;
assign n_18689 =  x_1341 & ~n_17830;
assign n_18690 =  n_17830 &  n_18665;
assign n_18691 = ~n_18689 & ~n_18690;
assign n_18692 =  x_1341 & ~n_18691;
assign n_18693 = ~x_1341 &  n_18691;
assign n_18694 = ~n_18692 & ~n_18693;
assign n_18695 =  x_1340 & ~n_17837;
assign n_18696 =  n_17837 &  n_18665;
assign n_18697 = ~n_18695 & ~n_18696;
assign n_18698 =  x_1340 & ~n_18697;
assign n_18699 = ~x_1340 &  n_18697;
assign n_18700 = ~n_18698 & ~n_18699;
assign n_18701 =  x_1339 & ~n_17844;
assign n_18702 =  n_17844 &  n_18665;
assign n_18703 = ~n_18701 & ~n_18702;
assign n_18704 =  x_1339 & ~n_18703;
assign n_18705 = ~x_1339 &  n_18703;
assign n_18706 = ~n_18704 & ~n_18705;
assign n_18707 =  x_1338 & ~n_17851;
assign n_18708 =  n_17851 &  n_18665;
assign n_18709 = ~n_18707 & ~n_18708;
assign n_18710 =  x_1338 & ~n_18709;
assign n_18711 = ~x_1338 &  n_18709;
assign n_18712 = ~n_18710 & ~n_18711;
assign n_18713 =  x_1337 & ~n_17789;
assign n_18714 = ~x_981 &  n_6109;
assign n_18715 = ~x_980 & ~x_1562;
assign n_18716 =  x_1618 & ~x_1635;
assign n_18717 = ~n_18715 & ~n_18716;
assign n_18718 = ~n_18714 &  n_18717;
assign n_18719 = ~x_3229 & ~n_18718;
assign n_18720 = ~x_1796 &  x_3229;
assign n_18721 =  x_1732 & ~n_18720;
assign n_18722 = ~n_18719 &  n_18721;
assign n_18723 =  n_17789 &  n_18722;
assign n_18724 = ~n_18713 & ~n_18723;
assign n_18725 =  x_1337 & ~n_18724;
assign n_18726 = ~x_1337 &  n_18724;
assign n_18727 = ~n_18725 & ~n_18726;
assign n_18728 =  x_1336 & ~n_17807;
assign n_18729 =  n_17807 &  n_18722;
assign n_18730 = ~n_18728 & ~n_18729;
assign n_18731 =  x_1336 & ~n_18730;
assign n_18732 = ~x_1336 &  n_18730;
assign n_18733 = ~n_18731 & ~n_18732;
assign n_18734 =  x_1335 & ~n_17815;
assign n_18735 =  n_17815 &  n_18722;
assign n_18736 = ~n_18734 & ~n_18735;
assign n_18737 =  x_1335 & ~n_18736;
assign n_18738 = ~x_1335 &  n_18736;
assign n_18739 = ~n_18737 & ~n_18738;
assign n_18740 =  x_1334 & ~n_17823;
assign n_18741 =  n_17823 &  n_18722;
assign n_18742 = ~n_18740 & ~n_18741;
assign n_18743 =  x_1334 & ~n_18742;
assign n_18744 = ~x_1334 &  n_18742;
assign n_18745 = ~n_18743 & ~n_18744;
assign n_18746 =  x_1333 & ~n_17830;
assign n_18747 =  n_17830 &  n_18722;
assign n_18748 = ~n_18746 & ~n_18747;
assign n_18749 =  x_1333 & ~n_18748;
assign n_18750 = ~x_1333 &  n_18748;
assign n_18751 = ~n_18749 & ~n_18750;
assign n_18752 =  x_1332 & ~n_17837;
assign n_18753 =  n_17837 &  n_18722;
assign n_18754 = ~n_18752 & ~n_18753;
assign n_18755 =  x_1332 & ~n_18754;
assign n_18756 = ~x_1332 &  n_18754;
assign n_18757 = ~n_18755 & ~n_18756;
assign n_18758 =  x_1331 & ~n_17844;
assign n_18759 =  n_17844 &  n_18722;
assign n_18760 = ~n_18758 & ~n_18759;
assign n_18761 =  x_1331 & ~n_18760;
assign n_18762 = ~x_1331 &  n_18760;
assign n_18763 = ~n_18761 & ~n_18762;
assign n_18764 =  x_1330 & ~n_17851;
assign n_18765 =  n_17851 &  n_18722;
assign n_18766 = ~n_18764 & ~n_18765;
assign n_18767 =  x_1330 & ~n_18766;
assign n_18768 = ~x_1330 &  n_18766;
assign n_18769 = ~n_18767 & ~n_18768;
assign n_18770 =  x_1329 & ~n_17789;
assign n_18771 = ~x_979 &  n_6109;
assign n_18772 =  x_1618 & ~x_1634;
assign n_18773 = ~x_978 & ~x_1562;
assign n_18774 = ~n_18772 & ~n_18773;
assign n_18775 = ~n_18771 &  n_18774;
assign n_18776 = ~x_3229 & ~n_18775;
assign n_18777 = ~x_1795 &  x_3229;
assign n_18778 =  x_1732 & ~n_18777;
assign n_18779 = ~n_18776 &  n_18778;
assign n_18780 =  n_17789 &  n_18779;
assign n_18781 = ~n_18770 & ~n_18780;
assign n_18782 =  x_1329 & ~n_18781;
assign n_18783 = ~x_1329 &  n_18781;
assign n_18784 = ~n_18782 & ~n_18783;
assign n_18785 =  x_1328 & ~n_17807;
assign n_18786 =  n_17807 &  n_18779;
assign n_18787 = ~n_18785 & ~n_18786;
assign n_18788 =  x_1328 & ~n_18787;
assign n_18789 = ~x_1328 &  n_18787;
assign n_18790 = ~n_18788 & ~n_18789;
assign n_18791 =  x_1327 & ~n_17815;
assign n_18792 =  n_17815 &  n_18779;
assign n_18793 = ~n_18791 & ~n_18792;
assign n_18794 =  x_1327 & ~n_18793;
assign n_18795 = ~x_1327 &  n_18793;
assign n_18796 = ~n_18794 & ~n_18795;
assign n_18797 =  x_1326 & ~n_17823;
assign n_18798 =  n_17823 &  n_18779;
assign n_18799 = ~n_18797 & ~n_18798;
assign n_18800 =  x_1326 & ~n_18799;
assign n_18801 = ~x_1326 &  n_18799;
assign n_18802 = ~n_18800 & ~n_18801;
assign n_18803 =  x_1325 & ~n_17830;
assign n_18804 =  n_17830 &  n_18779;
assign n_18805 = ~n_18803 & ~n_18804;
assign n_18806 =  x_1325 & ~n_18805;
assign n_18807 = ~x_1325 &  n_18805;
assign n_18808 = ~n_18806 & ~n_18807;
assign n_18809 =  x_1324 & ~n_17837;
assign n_18810 =  n_17837 &  n_18779;
assign n_18811 = ~n_18809 & ~n_18810;
assign n_18812 =  x_1324 & ~n_18811;
assign n_18813 = ~x_1324 &  n_18811;
assign n_18814 = ~n_18812 & ~n_18813;
assign n_18815 =  x_1323 & ~n_17844;
assign n_18816 =  n_17844 &  n_18779;
assign n_18817 = ~n_18815 & ~n_18816;
assign n_18818 =  x_1323 & ~n_18817;
assign n_18819 = ~x_1323 &  n_18817;
assign n_18820 = ~n_18818 & ~n_18819;
assign n_18821 =  x_1322 & ~n_17851;
assign n_18822 =  n_17851 &  n_18779;
assign n_18823 = ~n_18821 & ~n_18822;
assign n_18824 =  x_1322 & ~n_18823;
assign n_18825 = ~x_1322 &  n_18823;
assign n_18826 = ~n_18824 & ~n_18825;
assign n_18827 =  x_1321 & ~n_17789;
assign n_18828 = ~x_977 &  n_6109;
assign n_18829 = ~x_976 & ~x_1562;
assign n_18830 =  x_1618 & ~x_1633;
assign n_18831 = ~n_18829 & ~n_18830;
assign n_18832 = ~n_18828 &  n_18831;
assign n_18833 = ~x_3229 & ~n_18832;
assign n_18834 = ~x_1794 &  x_3229;
assign n_18835 =  x_1732 & ~n_18834;
assign n_18836 = ~n_18833 &  n_18835;
assign n_18837 =  n_17789 &  n_18836;
assign n_18838 = ~n_18827 & ~n_18837;
assign n_18839 =  x_1321 & ~n_18838;
assign n_18840 = ~x_1321 &  n_18838;
assign n_18841 = ~n_18839 & ~n_18840;
assign n_18842 =  x_1320 & ~n_17807;
assign n_18843 =  n_17807 &  n_18836;
assign n_18844 = ~n_18842 & ~n_18843;
assign n_18845 =  x_1320 & ~n_18844;
assign n_18846 = ~x_1320 &  n_18844;
assign n_18847 = ~n_18845 & ~n_18846;
assign n_18848 =  x_1319 & ~n_17815;
assign n_18849 =  n_17815 &  n_18836;
assign n_18850 = ~n_18848 & ~n_18849;
assign n_18851 =  x_1319 & ~n_18850;
assign n_18852 = ~x_1319 &  n_18850;
assign n_18853 = ~n_18851 & ~n_18852;
assign n_18854 =  x_1318 & ~n_17823;
assign n_18855 =  n_17823 &  n_18836;
assign n_18856 = ~n_18854 & ~n_18855;
assign n_18857 =  x_1318 & ~n_18856;
assign n_18858 = ~x_1318 &  n_18856;
assign n_18859 = ~n_18857 & ~n_18858;
assign n_18860 =  x_1317 & ~n_17830;
assign n_18861 =  n_17830 &  n_18836;
assign n_18862 = ~n_18860 & ~n_18861;
assign n_18863 =  x_1317 & ~n_18862;
assign n_18864 = ~x_1317 &  n_18862;
assign n_18865 = ~n_18863 & ~n_18864;
assign n_18866 =  x_1316 & ~n_17837;
assign n_18867 =  n_17837 &  n_18836;
assign n_18868 = ~n_18866 & ~n_18867;
assign n_18869 =  x_1316 & ~n_18868;
assign n_18870 = ~x_1316 &  n_18868;
assign n_18871 = ~n_18869 & ~n_18870;
assign n_18872 =  x_1315 & ~n_17844;
assign n_18873 =  n_17844 &  n_18836;
assign n_18874 = ~n_18872 & ~n_18873;
assign n_18875 =  x_1315 & ~n_18874;
assign n_18876 = ~x_1315 &  n_18874;
assign n_18877 = ~n_18875 & ~n_18876;
assign n_18878 =  x_1314 & ~n_17851;
assign n_18879 =  n_17851 &  n_18836;
assign n_18880 = ~n_18878 & ~n_18879;
assign n_18881 =  x_1314 & ~n_18880;
assign n_18882 = ~x_1314 &  n_18880;
assign n_18883 = ~n_18881 & ~n_18882;
assign n_18884 =  x_1313 & ~n_17789;
assign n_18885 = ~x_975 &  n_6109;
assign n_18886 = ~x_974 & ~x_1562;
assign n_18887 =  x_1618 & ~x_1632;
assign n_18888 = ~n_18886 & ~n_18887;
assign n_18889 = ~n_18885 &  n_18888;
assign n_18890 = ~x_3229 & ~n_18889;
assign n_18891 = ~x_1793 &  x_3229;
assign n_18892 =  x_1732 & ~n_18891;
assign n_18893 = ~n_18890 &  n_18892;
assign n_18894 =  n_17789 &  n_18893;
assign n_18895 = ~n_18884 & ~n_18894;
assign n_18896 =  x_1313 & ~n_18895;
assign n_18897 = ~x_1313 &  n_18895;
assign n_18898 = ~n_18896 & ~n_18897;
assign n_18899 =  x_1312 & ~n_17807;
assign n_18900 =  n_17807 &  n_18893;
assign n_18901 = ~n_18899 & ~n_18900;
assign n_18902 =  x_1312 & ~n_18901;
assign n_18903 = ~x_1312 &  n_18901;
assign n_18904 = ~n_18902 & ~n_18903;
assign n_18905 =  x_1311 & ~n_17815;
assign n_18906 =  n_17815 &  n_18893;
assign n_18907 = ~n_18905 & ~n_18906;
assign n_18908 =  x_1311 & ~n_18907;
assign n_18909 = ~x_1311 &  n_18907;
assign n_18910 = ~n_18908 & ~n_18909;
assign n_18911 =  x_1310 & ~n_17823;
assign n_18912 =  n_17823 &  n_18893;
assign n_18913 = ~n_18911 & ~n_18912;
assign n_18914 =  x_1310 & ~n_18913;
assign n_18915 = ~x_1310 &  n_18913;
assign n_18916 = ~n_18914 & ~n_18915;
assign n_18917 =  x_1309 & ~n_17830;
assign n_18918 =  n_17830 &  n_18893;
assign n_18919 = ~n_18917 & ~n_18918;
assign n_18920 =  x_1309 & ~n_18919;
assign n_18921 = ~x_1309 &  n_18919;
assign n_18922 = ~n_18920 & ~n_18921;
assign n_18923 =  x_1308 & ~n_17837;
assign n_18924 =  n_17837 &  n_18893;
assign n_18925 = ~n_18923 & ~n_18924;
assign n_18926 =  x_1308 & ~n_18925;
assign n_18927 = ~x_1308 &  n_18925;
assign n_18928 = ~n_18926 & ~n_18927;
assign n_18929 =  x_1307 & ~n_17844;
assign n_18930 =  n_17844 &  n_18893;
assign n_18931 = ~n_18929 & ~n_18930;
assign n_18932 =  x_1307 & ~n_18931;
assign n_18933 = ~x_1307 &  n_18931;
assign n_18934 = ~n_18932 & ~n_18933;
assign n_18935 =  x_1306 & ~n_17851;
assign n_18936 =  n_17851 &  n_18893;
assign n_18937 = ~n_18935 & ~n_18936;
assign n_18938 =  x_1306 & ~n_18937;
assign n_18939 = ~x_1306 &  n_18937;
assign n_18940 = ~n_18938 & ~n_18939;
assign n_18941 =  x_1305 & ~n_17789;
assign n_18942 = ~x_973 &  n_6109;
assign n_18943 = ~x_972 & ~x_1562;
assign n_18944 =  x_1618 & ~x_1631;
assign n_18945 = ~n_18943 & ~n_18944;
assign n_18946 = ~n_18942 &  n_18945;
assign n_18947 = ~x_3229 & ~n_18946;
assign n_18948 = ~x_1792 &  x_3229;
assign n_18949 =  x_1732 & ~n_18948;
assign n_18950 = ~n_18947 &  n_18949;
assign n_18951 =  n_17789 &  n_18950;
assign n_18952 = ~n_18941 & ~n_18951;
assign n_18953 =  x_1305 & ~n_18952;
assign n_18954 = ~x_1305 &  n_18952;
assign n_18955 = ~n_18953 & ~n_18954;
assign n_18956 =  x_1304 & ~n_17807;
assign n_18957 =  n_17807 &  n_18950;
assign n_18958 = ~n_18956 & ~n_18957;
assign n_18959 =  x_1304 & ~n_18958;
assign n_18960 = ~x_1304 &  n_18958;
assign n_18961 = ~n_18959 & ~n_18960;
assign n_18962 =  x_1303 & ~n_17815;
assign n_18963 =  n_17815 &  n_18950;
assign n_18964 = ~n_18962 & ~n_18963;
assign n_18965 =  x_1303 & ~n_18964;
assign n_18966 = ~x_1303 &  n_18964;
assign n_18967 = ~n_18965 & ~n_18966;
assign n_18968 =  x_1302 & ~n_17823;
assign n_18969 =  n_17823 &  n_18950;
assign n_18970 = ~n_18968 & ~n_18969;
assign n_18971 =  x_1302 & ~n_18970;
assign n_18972 = ~x_1302 &  n_18970;
assign n_18973 = ~n_18971 & ~n_18972;
assign n_18974 =  x_1301 & ~n_17830;
assign n_18975 =  n_17830 &  n_18950;
assign n_18976 = ~n_18974 & ~n_18975;
assign n_18977 =  x_1301 & ~n_18976;
assign n_18978 = ~x_1301 &  n_18976;
assign n_18979 = ~n_18977 & ~n_18978;
assign n_18980 =  x_1300 & ~n_17837;
assign n_18981 =  n_17837 &  n_18950;
assign n_18982 = ~n_18980 & ~n_18981;
assign n_18983 =  x_1300 & ~n_18982;
assign n_18984 = ~x_1300 &  n_18982;
assign n_18985 = ~n_18983 & ~n_18984;
assign n_18986 =  x_1299 & ~n_17844;
assign n_18987 =  n_17844 &  n_18950;
assign n_18988 = ~n_18986 & ~n_18987;
assign n_18989 =  x_1299 & ~n_18988;
assign n_18990 = ~x_1299 &  n_18988;
assign n_18991 = ~n_18989 & ~n_18990;
assign n_18992 =  x_1298 & ~n_17851;
assign n_18993 =  n_17851 &  n_18950;
assign n_18994 = ~n_18992 & ~n_18993;
assign n_18995 =  x_1298 & ~n_18994;
assign n_18996 = ~x_1298 &  n_18994;
assign n_18997 = ~n_18995 & ~n_18996;
assign n_18998 =  x_1297 & ~n_17789;
assign n_18999 = ~x_971 &  n_6109;
assign n_19000 = ~x_970 & ~x_1562;
assign n_19001 =  x_1618 & ~x_1630;
assign n_19002 = ~n_19000 & ~n_19001;
assign n_19003 = ~n_18999 &  n_19002;
assign n_19004 = ~x_3229 & ~n_19003;
assign n_19005 = ~x_1791 &  x_3229;
assign n_19006 =  x_1732 & ~n_19005;
assign n_19007 = ~n_19004 &  n_19006;
assign n_19008 =  n_17789 &  n_19007;
assign n_19009 = ~n_18998 & ~n_19008;
assign n_19010 =  x_1297 & ~n_19009;
assign n_19011 = ~x_1297 &  n_19009;
assign n_19012 = ~n_19010 & ~n_19011;
assign n_19013 =  x_1296 & ~n_17807;
assign n_19014 =  n_17807 &  n_19007;
assign n_19015 = ~n_19013 & ~n_19014;
assign n_19016 =  x_1296 & ~n_19015;
assign n_19017 = ~x_1296 &  n_19015;
assign n_19018 = ~n_19016 & ~n_19017;
assign n_19019 =  x_1295 & ~n_17815;
assign n_19020 =  n_17815 &  n_19007;
assign n_19021 = ~n_19019 & ~n_19020;
assign n_19022 =  x_1295 & ~n_19021;
assign n_19023 = ~x_1295 &  n_19021;
assign n_19024 = ~n_19022 & ~n_19023;
assign n_19025 =  x_1294 & ~n_17823;
assign n_19026 =  n_17823 &  n_19007;
assign n_19027 = ~n_19025 & ~n_19026;
assign n_19028 =  x_1294 & ~n_19027;
assign n_19029 = ~x_1294 &  n_19027;
assign n_19030 = ~n_19028 & ~n_19029;
assign n_19031 =  x_1293 & ~n_17830;
assign n_19032 =  n_17830 &  n_19007;
assign n_19033 = ~n_19031 & ~n_19032;
assign n_19034 =  x_1293 & ~n_19033;
assign n_19035 = ~x_1293 &  n_19033;
assign n_19036 = ~n_19034 & ~n_19035;
assign n_19037 =  x_1292 & ~n_17837;
assign n_19038 =  n_17837 &  n_19007;
assign n_19039 = ~n_19037 & ~n_19038;
assign n_19040 =  x_1292 & ~n_19039;
assign n_19041 = ~x_1292 &  n_19039;
assign n_19042 = ~n_19040 & ~n_19041;
assign n_19043 =  x_1291 & ~n_17844;
assign n_19044 =  n_17844 &  n_19007;
assign n_19045 = ~n_19043 & ~n_19044;
assign n_19046 =  x_1291 & ~n_19045;
assign n_19047 = ~x_1291 &  n_19045;
assign n_19048 = ~n_19046 & ~n_19047;
assign n_19049 =  x_1290 & ~n_17851;
assign n_19050 =  n_17851 &  n_19007;
assign n_19051 = ~n_19049 & ~n_19050;
assign n_19052 =  x_1290 & ~n_19051;
assign n_19053 = ~x_1290 &  n_19051;
assign n_19054 = ~n_19052 & ~n_19053;
assign n_19055 =  x_1289 & ~n_17789;
assign n_19056 = ~x_969 &  n_6109;
assign n_19057 = ~x_968 & ~x_1562;
assign n_19058 =  x_1618 & ~x_1629;
assign n_19059 = ~n_19057 & ~n_19058;
assign n_19060 = ~n_19056 &  n_19059;
assign n_19061 = ~x_3229 & ~n_19060;
assign n_19062 = ~x_1790 &  x_3229;
assign n_19063 =  x_1732 & ~n_19062;
assign n_19064 = ~n_19061 &  n_19063;
assign n_19065 =  n_17789 &  n_19064;
assign n_19066 = ~n_19055 & ~n_19065;
assign n_19067 =  x_1289 & ~n_19066;
assign n_19068 = ~x_1289 &  n_19066;
assign n_19069 = ~n_19067 & ~n_19068;
assign n_19070 =  x_1288 & ~n_17807;
assign n_19071 =  n_17807 &  n_19064;
assign n_19072 = ~n_19070 & ~n_19071;
assign n_19073 =  x_1288 & ~n_19072;
assign n_19074 = ~x_1288 &  n_19072;
assign n_19075 = ~n_19073 & ~n_19074;
assign n_19076 =  x_1287 & ~n_17815;
assign n_19077 =  n_17815 &  n_19064;
assign n_19078 = ~n_19076 & ~n_19077;
assign n_19079 =  x_1287 & ~n_19078;
assign n_19080 = ~x_1287 &  n_19078;
assign n_19081 = ~n_19079 & ~n_19080;
assign n_19082 =  x_1286 & ~n_17823;
assign n_19083 =  n_17823 &  n_19064;
assign n_19084 = ~n_19082 & ~n_19083;
assign n_19085 =  x_1286 & ~n_19084;
assign n_19086 = ~x_1286 &  n_19084;
assign n_19087 = ~n_19085 & ~n_19086;
assign n_19088 =  x_1285 & ~n_17830;
assign n_19089 =  n_17830 &  n_19064;
assign n_19090 = ~n_19088 & ~n_19089;
assign n_19091 =  x_1285 & ~n_19090;
assign n_19092 = ~x_1285 &  n_19090;
assign n_19093 = ~n_19091 & ~n_19092;
assign n_19094 =  x_1284 & ~n_17837;
assign n_19095 =  n_17837 &  n_19064;
assign n_19096 = ~n_19094 & ~n_19095;
assign n_19097 =  x_1284 & ~n_19096;
assign n_19098 = ~x_1284 &  n_19096;
assign n_19099 = ~n_19097 & ~n_19098;
assign n_19100 =  x_1283 & ~n_17844;
assign n_19101 =  n_17844 &  n_19064;
assign n_19102 = ~n_19100 & ~n_19101;
assign n_19103 =  x_1283 & ~n_19102;
assign n_19104 = ~x_1283 &  n_19102;
assign n_19105 = ~n_19103 & ~n_19104;
assign n_19106 =  x_1282 & ~n_17851;
assign n_19107 =  n_17851 &  n_19064;
assign n_19108 = ~n_19106 & ~n_19107;
assign n_19109 =  x_1282 & ~n_19108;
assign n_19110 = ~x_1282 &  n_19108;
assign n_19111 = ~n_19109 & ~n_19110;
assign n_19112 =  x_1281 & ~n_17789;
assign n_19113 = ~x_967 &  n_6109;
assign n_19114 =  x_1618 & ~x_1628;
assign n_19115 = ~x_966 & ~x_1562;
assign n_19116 = ~n_19114 & ~n_19115;
assign n_19117 = ~n_19113 &  n_19116;
assign n_19118 = ~x_3229 & ~n_19117;
assign n_19119 = ~x_1789 &  x_3229;
assign n_19120 =  x_1732 & ~n_19119;
assign n_19121 = ~n_19118 &  n_19120;
assign n_19122 =  n_17789 &  n_19121;
assign n_19123 = ~n_19112 & ~n_19122;
assign n_19124 =  x_1281 & ~n_19123;
assign n_19125 = ~x_1281 &  n_19123;
assign n_19126 = ~n_19124 & ~n_19125;
assign n_19127 =  x_1280 & ~n_17807;
assign n_19128 =  n_17807 &  n_19121;
assign n_19129 = ~n_19127 & ~n_19128;
assign n_19130 =  x_1280 & ~n_19129;
assign n_19131 = ~x_1280 &  n_19129;
assign n_19132 = ~n_19130 & ~n_19131;
assign n_19133 =  x_1279 & ~n_17815;
assign n_19134 =  n_17815 &  n_19121;
assign n_19135 = ~n_19133 & ~n_19134;
assign n_19136 =  x_1279 & ~n_19135;
assign n_19137 = ~x_1279 &  n_19135;
assign n_19138 = ~n_19136 & ~n_19137;
assign n_19139 =  x_1278 & ~n_17823;
assign n_19140 =  n_17823 &  n_19121;
assign n_19141 = ~n_19139 & ~n_19140;
assign n_19142 =  x_1278 & ~n_19141;
assign n_19143 = ~x_1278 &  n_19141;
assign n_19144 = ~n_19142 & ~n_19143;
assign n_19145 =  x_1277 & ~n_17830;
assign n_19146 =  n_17830 &  n_19121;
assign n_19147 = ~n_19145 & ~n_19146;
assign n_19148 =  x_1277 & ~n_19147;
assign n_19149 = ~x_1277 &  n_19147;
assign n_19150 = ~n_19148 & ~n_19149;
assign n_19151 =  x_1276 & ~n_17837;
assign n_19152 =  n_17837 &  n_19121;
assign n_19153 = ~n_19151 & ~n_19152;
assign n_19154 =  x_1276 & ~n_19153;
assign n_19155 = ~x_1276 &  n_19153;
assign n_19156 = ~n_19154 & ~n_19155;
assign n_19157 =  x_1275 & ~n_17844;
assign n_19158 =  n_17844 &  n_19121;
assign n_19159 = ~n_19157 & ~n_19158;
assign n_19160 =  x_1275 & ~n_19159;
assign n_19161 = ~x_1275 &  n_19159;
assign n_19162 = ~n_19160 & ~n_19161;
assign n_19163 =  x_1274 & ~n_17851;
assign n_19164 =  n_17851 &  n_19121;
assign n_19165 = ~n_19163 & ~n_19164;
assign n_19166 =  x_1274 & ~n_19165;
assign n_19167 = ~x_1274 &  n_19165;
assign n_19168 = ~n_19166 & ~n_19167;
assign n_19169 =  x_1273 & ~n_17789;
assign n_19170 = ~x_965 &  n_6109;
assign n_19171 =  x_1618 & ~x_1627;
assign n_19172 = ~x_964 & ~x_1562;
assign n_19173 = ~n_19171 & ~n_19172;
assign n_19174 = ~n_19170 &  n_19173;
assign n_19175 = ~x_3229 & ~n_19174;
assign n_19176 = ~x_1788 &  x_3229;
assign n_19177 =  x_1732 & ~n_19176;
assign n_19178 = ~n_19175 &  n_19177;
assign n_19179 =  n_17789 &  n_19178;
assign n_19180 = ~n_19169 & ~n_19179;
assign n_19181 =  x_1273 & ~n_19180;
assign n_19182 = ~x_1273 &  n_19180;
assign n_19183 = ~n_19181 & ~n_19182;
assign n_19184 =  x_1272 & ~n_17807;
assign n_19185 =  n_17807 &  n_19178;
assign n_19186 = ~n_19184 & ~n_19185;
assign n_19187 =  x_1272 & ~n_19186;
assign n_19188 = ~x_1272 &  n_19186;
assign n_19189 = ~n_19187 & ~n_19188;
assign n_19190 =  x_1271 & ~n_17815;
assign n_19191 =  n_17815 &  n_19178;
assign n_19192 = ~n_19190 & ~n_19191;
assign n_19193 =  x_1271 & ~n_19192;
assign n_19194 = ~x_1271 &  n_19192;
assign n_19195 = ~n_19193 & ~n_19194;
assign n_19196 =  x_1270 & ~n_17823;
assign n_19197 =  n_17823 &  n_19178;
assign n_19198 = ~n_19196 & ~n_19197;
assign n_19199 =  x_1270 & ~n_19198;
assign n_19200 = ~x_1270 &  n_19198;
assign n_19201 = ~n_19199 & ~n_19200;
assign n_19202 =  x_1269 & ~n_17830;
assign n_19203 =  n_17830 &  n_19178;
assign n_19204 = ~n_19202 & ~n_19203;
assign n_19205 =  x_1269 & ~n_19204;
assign n_19206 = ~x_1269 &  n_19204;
assign n_19207 = ~n_19205 & ~n_19206;
assign n_19208 =  x_1268 & ~n_17837;
assign n_19209 =  n_17837 &  n_19178;
assign n_19210 = ~n_19208 & ~n_19209;
assign n_19211 =  x_1268 & ~n_19210;
assign n_19212 = ~x_1268 &  n_19210;
assign n_19213 = ~n_19211 & ~n_19212;
assign n_19214 =  x_1267 & ~n_17844;
assign n_19215 =  n_17844 &  n_19178;
assign n_19216 = ~n_19214 & ~n_19215;
assign n_19217 =  x_1267 & ~n_19216;
assign n_19218 = ~x_1267 &  n_19216;
assign n_19219 = ~n_19217 & ~n_19218;
assign n_19220 =  x_1266 & ~n_17851;
assign n_19221 =  n_17851 &  n_19178;
assign n_19222 = ~n_19220 & ~n_19221;
assign n_19223 =  x_1266 & ~n_19222;
assign n_19224 = ~x_1266 &  n_19222;
assign n_19225 = ~n_19223 & ~n_19224;
assign n_19226 =  x_1265 & ~n_17789;
assign n_19227 = ~x_963 &  n_6109;
assign n_19228 =  x_1618 & ~x_1626;
assign n_19229 = ~x_962 & ~x_1562;
assign n_19230 = ~n_19228 & ~n_19229;
assign n_19231 = ~n_19227 &  n_19230;
assign n_19232 = ~x_3229 & ~n_19231;
assign n_19233 = ~x_1787 &  x_3229;
assign n_19234 =  x_1732 & ~n_19233;
assign n_19235 = ~n_19232 &  n_19234;
assign n_19236 =  n_17789 &  n_19235;
assign n_19237 = ~n_19226 & ~n_19236;
assign n_19238 =  x_1265 & ~n_19237;
assign n_19239 = ~x_1265 &  n_19237;
assign n_19240 = ~n_19238 & ~n_19239;
assign n_19241 =  x_1264 & ~n_17807;
assign n_19242 =  n_17807 &  n_19235;
assign n_19243 = ~n_19241 & ~n_19242;
assign n_19244 =  x_1264 & ~n_19243;
assign n_19245 = ~x_1264 &  n_19243;
assign n_19246 = ~n_19244 & ~n_19245;
assign n_19247 =  x_1263 & ~n_17815;
assign n_19248 =  n_17815 &  n_19235;
assign n_19249 = ~n_19247 & ~n_19248;
assign n_19250 =  x_1263 & ~n_19249;
assign n_19251 = ~x_1263 &  n_19249;
assign n_19252 = ~n_19250 & ~n_19251;
assign n_19253 =  x_1262 & ~n_17823;
assign n_19254 =  n_17823 &  n_19235;
assign n_19255 = ~n_19253 & ~n_19254;
assign n_19256 =  x_1262 & ~n_19255;
assign n_19257 = ~x_1262 &  n_19255;
assign n_19258 = ~n_19256 & ~n_19257;
assign n_19259 =  x_1261 & ~n_17830;
assign n_19260 =  n_17830 &  n_19235;
assign n_19261 = ~n_19259 & ~n_19260;
assign n_19262 =  x_1261 & ~n_19261;
assign n_19263 = ~x_1261 &  n_19261;
assign n_19264 = ~n_19262 & ~n_19263;
assign n_19265 =  x_1260 & ~n_17837;
assign n_19266 =  n_17837 &  n_19235;
assign n_19267 = ~n_19265 & ~n_19266;
assign n_19268 =  x_1260 & ~n_19267;
assign n_19269 = ~x_1260 &  n_19267;
assign n_19270 = ~n_19268 & ~n_19269;
assign n_19271 =  x_1259 & ~n_17844;
assign n_19272 =  n_17844 &  n_19235;
assign n_19273 = ~n_19271 & ~n_19272;
assign n_19274 =  x_1259 & ~n_19273;
assign n_19275 = ~x_1259 &  n_19273;
assign n_19276 = ~n_19274 & ~n_19275;
assign n_19277 =  x_1258 & ~n_17851;
assign n_19278 =  n_17851 &  n_19235;
assign n_19279 = ~n_19277 & ~n_19278;
assign n_19280 =  x_1258 & ~n_19279;
assign n_19281 = ~x_1258 &  n_19279;
assign n_19282 = ~n_19280 & ~n_19281;
assign n_19283 =  x_1257 & ~n_17789;
assign n_19284 = ~x_961 &  n_6109;
assign n_19285 = ~x_960 & ~x_1562;
assign n_19286 =  x_1618 & ~x_1625;
assign n_19287 = ~n_19285 & ~n_19286;
assign n_19288 = ~n_19284 &  n_19287;
assign n_19289 = ~x_3229 & ~n_19288;
assign n_19290 = ~x_1786 &  x_3229;
assign n_19291 =  x_1732 & ~n_19290;
assign n_19292 = ~n_19289 &  n_19291;
assign n_19293 =  n_17789 &  n_19292;
assign n_19294 = ~n_19283 & ~n_19293;
assign n_19295 =  x_1257 & ~n_19294;
assign n_19296 = ~x_1257 &  n_19294;
assign n_19297 = ~n_19295 & ~n_19296;
assign n_19298 =  x_1256 & ~n_17807;
assign n_19299 =  n_17807 &  n_19292;
assign n_19300 = ~n_19298 & ~n_19299;
assign n_19301 =  x_1256 & ~n_19300;
assign n_19302 = ~x_1256 &  n_19300;
assign n_19303 = ~n_19301 & ~n_19302;
assign n_19304 =  x_1255 & ~n_17815;
assign n_19305 =  n_17815 &  n_19292;
assign n_19306 = ~n_19304 & ~n_19305;
assign n_19307 =  x_1255 & ~n_19306;
assign n_19308 = ~x_1255 &  n_19306;
assign n_19309 = ~n_19307 & ~n_19308;
assign n_19310 =  x_1254 & ~n_17823;
assign n_19311 =  n_17823 &  n_19292;
assign n_19312 = ~n_19310 & ~n_19311;
assign n_19313 =  x_1254 & ~n_19312;
assign n_19314 = ~x_1254 &  n_19312;
assign n_19315 = ~n_19313 & ~n_19314;
assign n_19316 =  x_1253 & ~n_17830;
assign n_19317 =  n_17830 &  n_19292;
assign n_19318 = ~n_19316 & ~n_19317;
assign n_19319 =  x_1253 & ~n_19318;
assign n_19320 = ~x_1253 &  n_19318;
assign n_19321 = ~n_19319 & ~n_19320;
assign n_19322 =  x_1252 & ~n_17837;
assign n_19323 =  n_17837 &  n_19292;
assign n_19324 = ~n_19322 & ~n_19323;
assign n_19325 =  x_1252 & ~n_19324;
assign n_19326 = ~x_1252 &  n_19324;
assign n_19327 = ~n_19325 & ~n_19326;
assign n_19328 =  x_1251 & ~n_17844;
assign n_19329 =  n_17844 &  n_19292;
assign n_19330 = ~n_19328 & ~n_19329;
assign n_19331 =  x_1251 & ~n_19330;
assign n_19332 = ~x_1251 &  n_19330;
assign n_19333 = ~n_19331 & ~n_19332;
assign n_19334 =  x_1250 & ~n_17851;
assign n_19335 =  n_17851 &  n_19292;
assign n_19336 = ~n_19334 & ~n_19335;
assign n_19337 =  x_1250 & ~n_19336;
assign n_19338 = ~x_1250 &  n_19336;
assign n_19339 = ~n_19337 & ~n_19338;
assign n_19340 =  x_1249 & ~n_17789;
assign n_19341 = ~x_959 &  n_6109;
assign n_19342 = ~x_958 & ~x_1562;
assign n_19343 =  x_1618 & ~x_1624;
assign n_19344 = ~n_19342 & ~n_19343;
assign n_19345 = ~n_19341 &  n_19344;
assign n_19346 = ~x_3229 & ~n_19345;
assign n_19347 = ~x_1785 &  x_3229;
assign n_19348 =  x_1732 & ~n_19347;
assign n_19349 = ~n_19346 &  n_19348;
assign n_19350 =  n_17789 &  n_19349;
assign n_19351 = ~n_19340 & ~n_19350;
assign n_19352 =  x_1249 & ~n_19351;
assign n_19353 = ~x_1249 &  n_19351;
assign n_19354 = ~n_19352 & ~n_19353;
assign n_19355 =  x_1248 & ~n_17807;
assign n_19356 =  n_17807 &  n_19349;
assign n_19357 = ~n_19355 & ~n_19356;
assign n_19358 =  x_1248 & ~n_19357;
assign n_19359 = ~x_1248 &  n_19357;
assign n_19360 = ~n_19358 & ~n_19359;
assign n_19361 =  x_1247 & ~n_17815;
assign n_19362 =  n_17815 &  n_19349;
assign n_19363 = ~n_19361 & ~n_19362;
assign n_19364 =  x_1247 & ~n_19363;
assign n_19365 = ~x_1247 &  n_19363;
assign n_19366 = ~n_19364 & ~n_19365;
assign n_19367 =  x_1246 & ~n_17823;
assign n_19368 =  n_17823 &  n_19349;
assign n_19369 = ~n_19367 & ~n_19368;
assign n_19370 =  x_1246 & ~n_19369;
assign n_19371 = ~x_1246 &  n_19369;
assign n_19372 = ~n_19370 & ~n_19371;
assign n_19373 =  x_1245 & ~n_17830;
assign n_19374 =  n_17830 &  n_19349;
assign n_19375 = ~n_19373 & ~n_19374;
assign n_19376 =  x_1245 & ~n_19375;
assign n_19377 = ~x_1245 &  n_19375;
assign n_19378 = ~n_19376 & ~n_19377;
assign n_19379 =  x_1244 & ~n_17837;
assign n_19380 =  n_17837 &  n_19349;
assign n_19381 = ~n_19379 & ~n_19380;
assign n_19382 =  x_1244 & ~n_19381;
assign n_19383 = ~x_1244 &  n_19381;
assign n_19384 = ~n_19382 & ~n_19383;
assign n_19385 =  x_1243 & ~n_17844;
assign n_19386 =  n_17844 &  n_19349;
assign n_19387 = ~n_19385 & ~n_19386;
assign n_19388 =  x_1243 & ~n_19387;
assign n_19389 = ~x_1243 &  n_19387;
assign n_19390 = ~n_19388 & ~n_19389;
assign n_19391 =  x_1242 & ~n_17851;
assign n_19392 =  n_17851 &  n_19349;
assign n_19393 = ~n_19391 & ~n_19392;
assign n_19394 =  x_1242 & ~n_19393;
assign n_19395 = ~x_1242 &  n_19393;
assign n_19396 = ~n_19394 & ~n_19395;
assign n_19397 =  x_1241 & ~n_17789;
assign n_19398 = ~x_957 &  n_6109;
assign n_19399 = ~x_956 & ~x_1562;
assign n_19400 =  x_1618 & ~x_1623;
assign n_19401 = ~n_19399 & ~n_19400;
assign n_19402 = ~n_19398 &  n_19401;
assign n_19403 = ~x_3229 & ~n_19402;
assign n_19404 = ~x_1784 &  x_3229;
assign n_19405 =  x_1732 & ~n_19404;
assign n_19406 = ~n_19403 &  n_19405;
assign n_19407 =  n_17789 &  n_19406;
assign n_19408 = ~n_19397 & ~n_19407;
assign n_19409 =  x_1241 & ~n_19408;
assign n_19410 = ~x_1241 &  n_19408;
assign n_19411 = ~n_19409 & ~n_19410;
assign n_19412 =  x_1240 & ~n_17807;
assign n_19413 =  n_17807 &  n_19406;
assign n_19414 = ~n_19412 & ~n_19413;
assign n_19415 =  x_1240 & ~n_19414;
assign n_19416 = ~x_1240 &  n_19414;
assign n_19417 = ~n_19415 & ~n_19416;
assign n_19418 =  x_1239 & ~n_17815;
assign n_19419 =  n_17815 &  n_19406;
assign n_19420 = ~n_19418 & ~n_19419;
assign n_19421 =  x_1239 & ~n_19420;
assign n_19422 = ~x_1239 &  n_19420;
assign n_19423 = ~n_19421 & ~n_19422;
assign n_19424 =  x_1238 & ~n_17823;
assign n_19425 =  n_17823 &  n_19406;
assign n_19426 = ~n_19424 & ~n_19425;
assign n_19427 =  x_1238 & ~n_19426;
assign n_19428 = ~x_1238 &  n_19426;
assign n_19429 = ~n_19427 & ~n_19428;
assign n_19430 =  x_1237 & ~n_17830;
assign n_19431 =  n_17830 &  n_19406;
assign n_19432 = ~n_19430 & ~n_19431;
assign n_19433 =  x_1237 & ~n_19432;
assign n_19434 = ~x_1237 &  n_19432;
assign n_19435 = ~n_19433 & ~n_19434;
assign n_19436 =  x_1236 & ~n_17837;
assign n_19437 =  n_17837 &  n_19406;
assign n_19438 = ~n_19436 & ~n_19437;
assign n_19439 =  x_1236 & ~n_19438;
assign n_19440 = ~x_1236 &  n_19438;
assign n_19441 = ~n_19439 & ~n_19440;
assign n_19442 =  x_1235 & ~n_17844;
assign n_19443 =  n_17844 &  n_19406;
assign n_19444 = ~n_19442 & ~n_19443;
assign n_19445 =  x_1235 & ~n_19444;
assign n_19446 = ~x_1235 &  n_19444;
assign n_19447 = ~n_19445 & ~n_19446;
assign n_19448 =  x_1234 & ~n_17851;
assign n_19449 =  n_17851 &  n_19406;
assign n_19450 = ~n_19448 & ~n_19449;
assign n_19451 =  x_1234 & ~n_19450;
assign n_19452 = ~x_1234 &  n_19450;
assign n_19453 = ~n_19451 & ~n_19452;
assign n_19454 =  x_1233 & ~n_17789;
assign n_19455 = ~x_955 &  n_6109;
assign n_19456 = ~x_954 & ~x_1562;
assign n_19457 =  x_1618 & ~x_1622;
assign n_19458 = ~n_19456 & ~n_19457;
assign n_19459 = ~n_19455 &  n_19458;
assign n_19460 = ~x_3229 & ~n_19459;
assign n_19461 = ~x_1783 &  x_3229;
assign n_19462 =  x_1732 & ~n_19461;
assign n_19463 = ~n_19460 &  n_19462;
assign n_19464 =  n_17789 &  n_19463;
assign n_19465 = ~n_19454 & ~n_19464;
assign n_19466 =  x_1233 & ~n_19465;
assign n_19467 = ~x_1233 &  n_19465;
assign n_19468 = ~n_19466 & ~n_19467;
assign n_19469 =  x_1232 & ~n_17807;
assign n_19470 =  n_17807 &  n_19463;
assign n_19471 = ~n_19469 & ~n_19470;
assign n_19472 =  x_1232 & ~n_19471;
assign n_19473 = ~x_1232 &  n_19471;
assign n_19474 = ~n_19472 & ~n_19473;
assign n_19475 =  x_1231 & ~n_17815;
assign n_19476 =  n_17815 &  n_19463;
assign n_19477 = ~n_19475 & ~n_19476;
assign n_19478 =  x_1231 & ~n_19477;
assign n_19479 = ~x_1231 &  n_19477;
assign n_19480 = ~n_19478 & ~n_19479;
assign n_19481 =  x_1230 & ~n_17823;
assign n_19482 =  n_17823 &  n_19463;
assign n_19483 = ~n_19481 & ~n_19482;
assign n_19484 =  x_1230 & ~n_19483;
assign n_19485 = ~x_1230 &  n_19483;
assign n_19486 = ~n_19484 & ~n_19485;
assign n_19487 =  x_1229 & ~n_17830;
assign n_19488 =  n_17830 &  n_19463;
assign n_19489 = ~n_19487 & ~n_19488;
assign n_19490 =  x_1229 & ~n_19489;
assign n_19491 = ~x_1229 &  n_19489;
assign n_19492 = ~n_19490 & ~n_19491;
assign n_19493 =  x_1228 & ~n_17837;
assign n_19494 =  n_17837 &  n_19463;
assign n_19495 = ~n_19493 & ~n_19494;
assign n_19496 =  x_1228 & ~n_19495;
assign n_19497 = ~x_1228 &  n_19495;
assign n_19498 = ~n_19496 & ~n_19497;
assign n_19499 =  x_1227 & ~n_17844;
assign n_19500 =  n_17844 &  n_19463;
assign n_19501 = ~n_19499 & ~n_19500;
assign n_19502 =  x_1227 & ~n_19501;
assign n_19503 = ~x_1227 &  n_19501;
assign n_19504 = ~n_19502 & ~n_19503;
assign n_19505 =  x_1226 & ~n_17851;
assign n_19506 =  n_17851 &  n_19463;
assign n_19507 = ~n_19505 & ~n_19506;
assign n_19508 =  x_1226 & ~n_19507;
assign n_19509 = ~x_1226 &  n_19507;
assign n_19510 = ~n_19508 & ~n_19509;
assign n_19511 =  x_1225 & ~n_17789;
assign n_19512 = ~x_953 &  n_6109;
assign n_19513 = ~x_952 & ~x_1562;
assign n_19514 =  x_1618 & ~x_1621;
assign n_19515 = ~n_19513 & ~n_19514;
assign n_19516 = ~n_19512 &  n_19515;
assign n_19517 = ~x_3229 & ~n_19516;
assign n_19518 = ~x_1782 &  x_3229;
assign n_19519 =  x_1732 & ~n_19518;
assign n_19520 = ~n_19517 &  n_19519;
assign n_19521 =  n_17789 &  n_19520;
assign n_19522 = ~n_19511 & ~n_19521;
assign n_19523 =  x_1225 & ~n_19522;
assign n_19524 = ~x_1225 &  n_19522;
assign n_19525 = ~n_19523 & ~n_19524;
assign n_19526 =  x_1224 & ~n_17807;
assign n_19527 =  n_17807 &  n_19520;
assign n_19528 = ~n_19526 & ~n_19527;
assign n_19529 =  x_1224 & ~n_19528;
assign n_19530 = ~x_1224 &  n_19528;
assign n_19531 = ~n_19529 & ~n_19530;
assign n_19532 =  x_1223 & ~n_17815;
assign n_19533 =  n_17815 &  n_19520;
assign n_19534 = ~n_19532 & ~n_19533;
assign n_19535 =  x_1223 & ~n_19534;
assign n_19536 = ~x_1223 &  n_19534;
assign n_19537 = ~n_19535 & ~n_19536;
assign n_19538 =  x_1222 & ~n_17823;
assign n_19539 =  n_17823 &  n_19520;
assign n_19540 = ~n_19538 & ~n_19539;
assign n_19541 =  x_1222 & ~n_19540;
assign n_19542 = ~x_1222 &  n_19540;
assign n_19543 = ~n_19541 & ~n_19542;
assign n_19544 =  x_1221 & ~n_17830;
assign n_19545 =  n_17830 &  n_19520;
assign n_19546 = ~n_19544 & ~n_19545;
assign n_19547 =  x_1221 & ~n_19546;
assign n_19548 = ~x_1221 &  n_19546;
assign n_19549 = ~n_19547 & ~n_19548;
assign n_19550 =  x_1220 & ~n_17837;
assign n_19551 =  n_17837 &  n_19520;
assign n_19552 = ~n_19550 & ~n_19551;
assign n_19553 =  x_1220 & ~n_19552;
assign n_19554 = ~x_1220 &  n_19552;
assign n_19555 = ~n_19553 & ~n_19554;
assign n_19556 =  x_1219 & ~n_17844;
assign n_19557 =  n_17844 &  n_19520;
assign n_19558 = ~n_19556 & ~n_19557;
assign n_19559 =  x_1219 & ~n_19558;
assign n_19560 = ~x_1219 &  n_19558;
assign n_19561 = ~n_19559 & ~n_19560;
assign n_19562 =  x_1218 & ~n_17851;
assign n_19563 =  n_17851 &  n_19520;
assign n_19564 = ~n_19562 & ~n_19563;
assign n_19565 =  x_1218 & ~n_19564;
assign n_19566 = ~x_1218 &  n_19564;
assign n_19567 = ~n_19565 & ~n_19566;
assign n_19568 =  x_1217 & ~n_17789;
assign n_19569 = ~x_951 &  n_6109;
assign n_19570 =  x_1618 & ~x_1620;
assign n_19571 = ~x_950 & ~x_1562;
assign n_19572 = ~n_19570 & ~n_19571;
assign n_19573 = ~n_19569 &  n_19572;
assign n_19574 = ~x_3229 & ~n_19573;
assign n_19575 = ~x_1781 &  x_3229;
assign n_19576 =  x_1732 & ~n_19575;
assign n_19577 = ~n_19574 &  n_19576;
assign n_19578 =  n_17789 &  n_19577;
assign n_19579 = ~n_19568 & ~n_19578;
assign n_19580 =  x_1217 & ~n_19579;
assign n_19581 = ~x_1217 &  n_19579;
assign n_19582 = ~n_19580 & ~n_19581;
assign n_19583 =  x_1216 & ~n_17807;
assign n_19584 =  n_17807 &  n_19577;
assign n_19585 = ~n_19583 & ~n_19584;
assign n_19586 =  x_1216 & ~n_19585;
assign n_19587 = ~x_1216 &  n_19585;
assign n_19588 = ~n_19586 & ~n_19587;
assign n_19589 =  x_1215 & ~n_17815;
assign n_19590 =  n_17815 &  n_19577;
assign n_19591 = ~n_19589 & ~n_19590;
assign n_19592 =  x_1215 & ~n_19591;
assign n_19593 = ~x_1215 &  n_19591;
assign n_19594 = ~n_19592 & ~n_19593;
assign n_19595 =  x_1214 & ~n_17823;
assign n_19596 =  n_17823 &  n_19577;
assign n_19597 = ~n_19595 & ~n_19596;
assign n_19598 =  x_1214 & ~n_19597;
assign n_19599 = ~x_1214 &  n_19597;
assign n_19600 = ~n_19598 & ~n_19599;
assign n_19601 =  x_1213 & ~n_17830;
assign n_19602 =  n_17830 &  n_19577;
assign n_19603 = ~n_19601 & ~n_19602;
assign n_19604 =  x_1213 & ~n_19603;
assign n_19605 = ~x_1213 &  n_19603;
assign n_19606 = ~n_19604 & ~n_19605;
assign n_19607 =  x_1212 & ~n_17837;
assign n_19608 =  n_17837 &  n_19577;
assign n_19609 = ~n_19607 & ~n_19608;
assign n_19610 =  x_1212 & ~n_19609;
assign n_19611 = ~x_1212 &  n_19609;
assign n_19612 = ~n_19610 & ~n_19611;
assign n_19613 =  x_1211 & ~n_17844;
assign n_19614 =  n_17844 &  n_19577;
assign n_19615 = ~n_19613 & ~n_19614;
assign n_19616 =  x_1211 & ~n_19615;
assign n_19617 = ~x_1211 &  n_19615;
assign n_19618 = ~n_19616 & ~n_19617;
assign n_19619 =  x_1210 & ~n_17851;
assign n_19620 =  n_17851 &  n_19577;
assign n_19621 = ~n_19619 & ~n_19620;
assign n_19622 =  x_1210 & ~n_19621;
assign n_19623 = ~x_1210 &  n_19621;
assign n_19624 = ~n_19622 & ~n_19623;
assign n_19625 =  x_1209 & ~n_17789;
assign n_19626 = ~x_949 &  n_6109;
assign n_19627 = ~x_948 & ~x_1562;
assign n_19628 =  x_1618 & ~x_1619;
assign n_19629 = ~n_19627 & ~n_19628;
assign n_19630 = ~n_19626 &  n_19629;
assign n_19631 = ~x_3229 & ~n_19630;
assign n_19632 = ~x_1780 &  x_3229;
assign n_19633 =  x_1732 & ~n_19632;
assign n_19634 = ~n_19631 &  n_19633;
assign n_19635 =  n_17789 &  n_19634;
assign n_19636 = ~n_19625 & ~n_19635;
assign n_19637 =  x_1209 & ~n_19636;
assign n_19638 = ~x_1209 &  n_19636;
assign n_19639 = ~n_19637 & ~n_19638;
assign n_19640 =  x_1208 & ~n_17807;
assign n_19641 =  n_17807 &  n_19634;
assign n_19642 = ~n_19640 & ~n_19641;
assign n_19643 =  x_1208 & ~n_19642;
assign n_19644 = ~x_1208 &  n_19642;
assign n_19645 = ~n_19643 & ~n_19644;
assign n_19646 =  x_1207 & ~n_17815;
assign n_19647 =  n_17815 &  n_19634;
assign n_19648 = ~n_19646 & ~n_19647;
assign n_19649 =  x_1207 & ~n_19648;
assign n_19650 = ~x_1207 &  n_19648;
assign n_19651 = ~n_19649 & ~n_19650;
assign n_19652 =  x_1206 & ~n_17823;
assign n_19653 =  n_17823 &  n_19634;
assign n_19654 = ~n_19652 & ~n_19653;
assign n_19655 =  x_1206 & ~n_19654;
assign n_19656 = ~x_1206 &  n_19654;
assign n_19657 = ~n_19655 & ~n_19656;
assign n_19658 =  x_1205 & ~n_17830;
assign n_19659 =  n_17830 &  n_19634;
assign n_19660 = ~n_19658 & ~n_19659;
assign n_19661 =  x_1205 & ~n_19660;
assign n_19662 = ~x_1205 &  n_19660;
assign n_19663 = ~n_19661 & ~n_19662;
assign n_19664 =  x_1204 & ~n_17837;
assign n_19665 =  n_17837 &  n_19634;
assign n_19666 = ~n_19664 & ~n_19665;
assign n_19667 =  x_1204 & ~n_19666;
assign n_19668 = ~x_1204 &  n_19666;
assign n_19669 = ~n_19667 & ~n_19668;
assign n_19670 =  x_1203 & ~n_17844;
assign n_19671 =  n_17844 &  n_19634;
assign n_19672 = ~n_19670 & ~n_19671;
assign n_19673 =  x_1203 & ~n_19672;
assign n_19674 = ~x_1203 &  n_19672;
assign n_19675 = ~n_19673 & ~n_19674;
assign n_19676 =  x_1202 & ~n_17851;
assign n_19677 =  n_17851 &  n_19634;
assign n_19678 = ~n_19676 & ~n_19677;
assign n_19679 =  x_1202 & ~n_19678;
assign n_19680 = ~x_1202 &  n_19678;
assign n_19681 = ~n_19679 & ~n_19680;
assign n_19682 =  x_1201 & ~n_6171;
assign n_19683 = ~x_1201 &  n_6171;
assign n_19684 = ~n_19682 & ~n_19683;
assign n_19685 =  x_1200 & ~n_6204;
assign n_19686 = ~x_1200 &  n_6204;
assign n_19687 = ~n_19685 & ~n_19686;
assign n_19688 =  x_1199 & ~n_6237;
assign n_19689 = ~x_1199 &  n_6237;
assign n_19690 = ~n_19688 & ~n_19689;
assign n_19691 =  x_1198 & ~n_6270;
assign n_19692 = ~x_1198 &  n_6270;
assign n_19693 = ~n_19691 & ~n_19692;
assign n_19694 =  x_1197 & ~n_6303;
assign n_19695 = ~x_1197 &  n_6303;
assign n_19696 = ~n_19694 & ~n_19695;
assign n_19697 =  x_1196 & ~n_6336;
assign n_19698 = ~x_1196 &  n_6336;
assign n_19699 = ~n_19697 & ~n_19698;
assign n_19700 =  x_1195 & ~n_6369;
assign n_19701 = ~x_1195 &  n_6369;
assign n_19702 = ~n_19700 & ~n_19701;
assign n_19703 =  x_1194 & ~n_6402;
assign n_19704 = ~x_1194 &  n_6402;
assign n_19705 = ~n_19703 & ~n_19704;
assign n_19706 =  x_1193 & ~n_6436;
assign n_19707 = ~x_1193 &  n_6436;
assign n_19708 = ~n_19706 & ~n_19707;
assign n_19709 =  x_1192 & ~n_6469;
assign n_19710 = ~x_1192 &  n_6469;
assign n_19711 = ~n_19709 & ~n_19710;
assign n_19712 =  x_1191 & ~n_6502;
assign n_19713 = ~x_1191 &  n_6502;
assign n_19714 = ~n_19712 & ~n_19713;
assign n_19715 =  x_1190 & ~n_6535;
assign n_19716 = ~x_1190 &  n_6535;
assign n_19717 = ~n_19715 & ~n_19716;
assign n_19718 =  x_1189 & ~n_6568;
assign n_19719 = ~x_1189 &  n_6568;
assign n_19720 = ~n_19718 & ~n_19719;
assign n_19721 =  x_1188 & ~n_6601;
assign n_19722 = ~x_1188 &  n_6601;
assign n_19723 = ~n_19721 & ~n_19722;
assign n_19724 =  x_1187 & ~n_6634;
assign n_19725 = ~x_1187 &  n_6634;
assign n_19726 = ~n_19724 & ~n_19725;
assign n_19727 =  x_1186 & ~n_6660;
assign n_19728 = ~x_1186 &  n_6660;
assign n_19729 = ~n_19727 & ~n_19728;
assign n_19730 =  x_1185 & ~n_6701;
assign n_19731 = ~x_1185 &  n_6701;
assign n_19732 = ~n_19730 & ~n_19731;
assign n_19733 =  x_1184 & ~n_6734;
assign n_19734 = ~x_1184 &  n_6734;
assign n_19735 = ~n_19733 & ~n_19734;
assign n_19736 =  x_1183 & ~n_6767;
assign n_19737 = ~x_1183 &  n_6767;
assign n_19738 = ~n_19736 & ~n_19737;
assign n_19739 =  x_1182 & ~n_6800;
assign n_19740 = ~x_1182 &  n_6800;
assign n_19741 = ~n_19739 & ~n_19740;
assign n_19742 =  x_1181 & ~n_6833;
assign n_19743 = ~x_1181 &  n_6833;
assign n_19744 = ~n_19742 & ~n_19743;
assign n_19745 =  x_1180 & ~n_6866;
assign n_19746 = ~x_1180 &  n_6866;
assign n_19747 = ~n_19745 & ~n_19746;
assign n_19748 =  x_1179 & ~n_6899;
assign n_19749 = ~x_1179 &  n_6899;
assign n_19750 = ~n_19748 & ~n_19749;
assign n_19751 =  x_1178 & ~n_6932;
assign n_19752 = ~x_1178 &  n_6932;
assign n_19753 = ~n_19751 & ~n_19752;
assign n_19754 =  x_1177 & ~n_6966;
assign n_19755 = ~x_1177 &  n_6966;
assign n_19756 = ~n_19754 & ~n_19755;
assign n_19757 =  x_1176 & ~n_6999;
assign n_19758 = ~x_1176 &  n_6999;
assign n_19759 = ~n_19757 & ~n_19758;
assign n_19760 =  x_1175 & ~n_7032;
assign n_19761 = ~x_1175 &  n_7032;
assign n_19762 = ~n_19760 & ~n_19761;
assign n_19763 =  x_1174 & ~n_7065;
assign n_19764 = ~x_1174 &  n_7065;
assign n_19765 = ~n_19763 & ~n_19764;
assign n_19766 =  x_1173 & ~n_7098;
assign n_19767 = ~x_1173 &  n_7098;
assign n_19768 = ~n_19766 & ~n_19767;
assign n_19769 =  x_1172 & ~n_7131;
assign n_19770 = ~x_1172 &  n_7131;
assign n_19771 = ~n_19769 & ~n_19770;
assign n_19772 =  x_1171 & ~n_7164;
assign n_19773 = ~x_1171 &  n_7164;
assign n_19774 = ~n_19772 & ~n_19773;
assign n_19775 =  x_1170 & ~n_7190;
assign n_19776 = ~x_1170 &  n_7190;
assign n_19777 = ~n_19775 & ~n_19776;
assign n_19778 =  x_1169 & ~n_7231;
assign n_19779 = ~x_1169 &  n_7231;
assign n_19780 = ~n_19778 & ~n_19779;
assign n_19781 =  x_1168 & ~n_7264;
assign n_19782 = ~x_1168 &  n_7264;
assign n_19783 = ~n_19781 & ~n_19782;
assign n_19784 =  x_1167 & ~n_7297;
assign n_19785 = ~x_1167 &  n_7297;
assign n_19786 = ~n_19784 & ~n_19785;
assign n_19787 =  x_1166 & ~n_7330;
assign n_19788 = ~x_1166 &  n_7330;
assign n_19789 = ~n_19787 & ~n_19788;
assign n_19790 =  x_1165 & ~n_7363;
assign n_19791 = ~x_1165 &  n_7363;
assign n_19792 = ~n_19790 & ~n_19791;
assign n_19793 =  x_1164 & ~n_7396;
assign n_19794 = ~x_1164 &  n_7396;
assign n_19795 = ~n_19793 & ~n_19794;
assign n_19796 =  x_1163 & ~n_7429;
assign n_19797 = ~x_1163 &  n_7429;
assign n_19798 = ~n_19796 & ~n_19797;
assign n_19799 =  x_1162 & ~n_7462;
assign n_19800 = ~x_1162 &  n_7462;
assign n_19801 = ~n_19799 & ~n_19800;
assign n_19802 =  x_1161 & ~n_7496;
assign n_19803 = ~x_1161 &  n_7496;
assign n_19804 = ~n_19802 & ~n_19803;
assign n_19805 =  x_1160 & ~n_7529;
assign n_19806 = ~x_1160 &  n_7529;
assign n_19807 = ~n_19805 & ~n_19806;
assign n_19808 =  x_1159 & ~n_7562;
assign n_19809 = ~x_1159 &  n_7562;
assign n_19810 = ~n_19808 & ~n_19809;
assign n_19811 =  x_1158 & ~n_7595;
assign n_19812 = ~x_1158 &  n_7595;
assign n_19813 = ~n_19811 & ~n_19812;
assign n_19814 =  x_1157 & ~n_7628;
assign n_19815 = ~x_1157 &  n_7628;
assign n_19816 = ~n_19814 & ~n_19815;
assign n_19817 =  x_1156 & ~n_7661;
assign n_19818 = ~x_1156 &  n_7661;
assign n_19819 = ~n_19817 & ~n_19818;
assign n_19820 =  x_1155 & ~n_7694;
assign n_19821 = ~x_1155 &  n_7694;
assign n_19822 = ~n_19820 & ~n_19821;
assign n_19823 =  x_1154 & ~n_7720;
assign n_19824 = ~x_1154 &  n_7720;
assign n_19825 = ~n_19823 & ~n_19824;
assign n_19826 =  x_1153 & ~n_7761;
assign n_19827 = ~x_1153 &  n_7761;
assign n_19828 = ~n_19826 & ~n_19827;
assign n_19829 =  x_1152 & ~n_7794;
assign n_19830 = ~x_1152 &  n_7794;
assign n_19831 = ~n_19829 & ~n_19830;
assign n_19832 =  x_1151 & ~n_7827;
assign n_19833 = ~x_1151 &  n_7827;
assign n_19834 = ~n_19832 & ~n_19833;
assign n_19835 =  x_1150 & ~n_7860;
assign n_19836 = ~x_1150 &  n_7860;
assign n_19837 = ~n_19835 & ~n_19836;
assign n_19838 =  x_1149 & ~n_7893;
assign n_19839 = ~x_1149 &  n_7893;
assign n_19840 = ~n_19838 & ~n_19839;
assign n_19841 =  x_1148 & ~n_7926;
assign n_19842 = ~x_1148 &  n_7926;
assign n_19843 = ~n_19841 & ~n_19842;
assign n_19844 =  x_1147 & ~n_7959;
assign n_19845 = ~x_1147 &  n_7959;
assign n_19846 = ~n_19844 & ~n_19845;
assign n_19847 =  x_1146 & ~n_7992;
assign n_19848 = ~x_1146 &  n_7992;
assign n_19849 = ~n_19847 & ~n_19848;
assign n_19850 =  x_1145 & ~n_8026;
assign n_19851 = ~x_1145 &  n_8026;
assign n_19852 = ~n_19850 & ~n_19851;
assign n_19853 =  x_1144 & ~n_8059;
assign n_19854 = ~x_1144 &  n_8059;
assign n_19855 = ~n_19853 & ~n_19854;
assign n_19856 =  x_1143 & ~n_8092;
assign n_19857 = ~x_1143 &  n_8092;
assign n_19858 = ~n_19856 & ~n_19857;
assign n_19859 =  x_1142 & ~n_8125;
assign n_19860 = ~x_1142 &  n_8125;
assign n_19861 = ~n_19859 & ~n_19860;
assign n_19862 =  x_1141 & ~n_8158;
assign n_19863 = ~x_1141 &  n_8158;
assign n_19864 = ~n_19862 & ~n_19863;
assign n_19865 =  x_1140 & ~n_8191;
assign n_19866 = ~x_1140 &  n_8191;
assign n_19867 = ~n_19865 & ~n_19866;
assign n_19868 =  x_1139 &  n_6165;
assign n_19869 = ~x_1139 & ~n_6165;
assign n_19870 = ~n_19868 & ~n_19869;
assign n_19871 =  x_1138 &  n_6198;
assign n_19872 = ~x_1138 & ~n_6198;
assign n_19873 = ~n_19871 & ~n_19872;
assign n_19874 =  x_1137 &  n_6231;
assign n_19875 = ~x_1137 & ~n_6231;
assign n_19876 = ~n_19874 & ~n_19875;
assign n_19877 =  x_1136 &  n_6264;
assign n_19878 = ~x_1136 & ~n_6264;
assign n_19879 = ~n_19877 & ~n_19878;
assign n_19880 =  x_1135 &  n_6297;
assign n_19881 = ~x_1135 & ~n_6297;
assign n_19882 = ~n_19880 & ~n_19881;
assign n_19883 =  x_1134 &  n_6330;
assign n_19884 = ~x_1134 & ~n_6330;
assign n_19885 = ~n_19883 & ~n_19884;
assign n_19886 =  x_1133 &  n_6363;
assign n_19887 = ~x_1133 & ~n_6363;
assign n_19888 = ~n_19886 & ~n_19887;
assign n_19889 =  x_1132 &  n_6396;
assign n_19890 = ~x_1132 & ~n_6396;
assign n_19891 = ~n_19889 & ~n_19890;
assign n_19892 =  x_1131 &  n_6430;
assign n_19893 = ~x_1131 & ~n_6430;
assign n_19894 = ~n_19892 & ~n_19893;
assign n_19895 =  x_1130 &  n_6463;
assign n_19896 = ~x_1130 & ~n_6463;
assign n_19897 = ~n_19895 & ~n_19896;
assign n_19898 =  x_1129 &  n_6496;
assign n_19899 = ~x_1129 & ~n_6496;
assign n_19900 = ~n_19898 & ~n_19899;
assign n_19901 =  x_1128 &  n_6529;
assign n_19902 = ~x_1128 & ~n_6529;
assign n_19903 = ~n_19901 & ~n_19902;
assign n_19904 =  x_1127 &  n_6562;
assign n_19905 = ~x_1127 & ~n_6562;
assign n_19906 = ~n_19904 & ~n_19905;
assign n_19907 =  x_1126 &  n_6595;
assign n_19908 = ~x_1126 & ~n_6595;
assign n_19909 = ~n_19907 & ~n_19908;
assign n_19910 =  x_1125 &  n_6628;
assign n_19911 = ~x_1125 & ~n_6628;
assign n_19912 = ~n_19910 & ~n_19911;
assign n_19913 =  x_1124 &  n_6665;
assign n_19914 = ~x_1124 & ~n_6665;
assign n_19915 = ~n_19913 & ~n_19914;
assign n_19916 =  x_1123 &  n_6695;
assign n_19917 = ~x_1123 & ~n_6695;
assign n_19918 = ~n_19916 & ~n_19917;
assign n_19919 =  x_1122 &  n_6728;
assign n_19920 = ~x_1122 & ~n_6728;
assign n_19921 = ~n_19919 & ~n_19920;
assign n_19922 =  x_1121 &  n_6761;
assign n_19923 = ~x_1121 & ~n_6761;
assign n_19924 = ~n_19922 & ~n_19923;
assign n_19925 =  x_1120 &  n_6794;
assign n_19926 = ~x_1120 & ~n_6794;
assign n_19927 = ~n_19925 & ~n_19926;
assign n_19928 =  x_1119 &  n_6827;
assign n_19929 = ~x_1119 & ~n_6827;
assign n_19930 = ~n_19928 & ~n_19929;
assign n_19931 =  x_1118 &  n_6860;
assign n_19932 = ~x_1118 & ~n_6860;
assign n_19933 = ~n_19931 & ~n_19932;
assign n_19934 =  x_1117 &  n_6893;
assign n_19935 = ~x_1117 & ~n_6893;
assign n_19936 = ~n_19934 & ~n_19935;
assign n_19937 =  x_1116 &  n_6926;
assign n_19938 = ~x_1116 & ~n_6926;
assign n_19939 = ~n_19937 & ~n_19938;
assign n_19940 =  x_1115 &  n_6960;
assign n_19941 = ~x_1115 & ~n_6960;
assign n_19942 = ~n_19940 & ~n_19941;
assign n_19943 =  x_1114 &  n_6993;
assign n_19944 = ~x_1114 & ~n_6993;
assign n_19945 = ~n_19943 & ~n_19944;
assign n_19946 =  x_1113 &  n_7026;
assign n_19947 = ~x_1113 & ~n_7026;
assign n_19948 = ~n_19946 & ~n_19947;
assign n_19949 =  x_1112 &  n_7059;
assign n_19950 = ~x_1112 & ~n_7059;
assign n_19951 = ~n_19949 & ~n_19950;
assign n_19952 =  x_1111 &  n_7092;
assign n_19953 = ~x_1111 & ~n_7092;
assign n_19954 = ~n_19952 & ~n_19953;
assign n_19955 =  x_1110 &  n_7125;
assign n_19956 = ~x_1110 & ~n_7125;
assign n_19957 = ~n_19955 & ~n_19956;
assign n_19958 =  x_1109 &  n_7158;
assign n_19959 = ~x_1109 & ~n_7158;
assign n_19960 = ~n_19958 & ~n_19959;
assign n_19961 =  x_1108 &  n_7195;
assign n_19962 = ~x_1108 & ~n_7195;
assign n_19963 = ~n_19961 & ~n_19962;
assign n_19964 =  x_1107 &  n_7225;
assign n_19965 = ~x_1107 & ~n_7225;
assign n_19966 = ~n_19964 & ~n_19965;
assign n_19967 =  x_1106 &  n_7258;
assign n_19968 = ~x_1106 & ~n_7258;
assign n_19969 = ~n_19967 & ~n_19968;
assign n_19970 =  x_1105 &  n_7291;
assign n_19971 = ~x_1105 & ~n_7291;
assign n_19972 = ~n_19970 & ~n_19971;
assign n_19973 =  x_1104 &  n_7324;
assign n_19974 = ~x_1104 & ~n_7324;
assign n_19975 = ~n_19973 & ~n_19974;
assign n_19976 =  x_1103 &  n_7357;
assign n_19977 = ~x_1103 & ~n_7357;
assign n_19978 = ~n_19976 & ~n_19977;
assign n_19979 =  x_1102 &  n_7390;
assign n_19980 = ~x_1102 & ~n_7390;
assign n_19981 = ~n_19979 & ~n_19980;
assign n_19982 =  x_1101 &  n_7423;
assign n_19983 = ~x_1101 & ~n_7423;
assign n_19984 = ~n_19982 & ~n_19983;
assign n_19985 =  x_1100 &  n_7456;
assign n_19986 = ~x_1100 & ~n_7456;
assign n_19987 = ~n_19985 & ~n_19986;
assign n_19988 =  x_1099 &  n_7490;
assign n_19989 = ~x_1099 & ~n_7490;
assign n_19990 = ~n_19988 & ~n_19989;
assign n_19991 =  x_1098 &  n_7523;
assign n_19992 = ~x_1098 & ~n_7523;
assign n_19993 = ~n_19991 & ~n_19992;
assign n_19994 =  x_1097 &  n_7556;
assign n_19995 = ~x_1097 & ~n_7556;
assign n_19996 = ~n_19994 & ~n_19995;
assign n_19997 =  x_1096 &  n_7589;
assign n_19998 = ~x_1096 & ~n_7589;
assign n_19999 = ~n_19997 & ~n_19998;
assign n_20000 =  x_1095 &  n_7622;
assign n_20001 = ~x_1095 & ~n_7622;
assign n_20002 = ~n_20000 & ~n_20001;
assign n_20003 =  x_1094 &  n_7655;
assign n_20004 = ~x_1094 & ~n_7655;
assign n_20005 = ~n_20003 & ~n_20004;
assign n_20006 =  x_1093 &  n_7688;
assign n_20007 = ~x_1093 & ~n_7688;
assign n_20008 = ~n_20006 & ~n_20007;
assign n_20009 =  x_1092 &  n_7725;
assign n_20010 = ~x_1092 & ~n_7725;
assign n_20011 = ~n_20009 & ~n_20010;
assign n_20012 =  x_1091 &  n_7755;
assign n_20013 = ~x_1091 & ~n_7755;
assign n_20014 = ~n_20012 & ~n_20013;
assign n_20015 =  x_1090 &  n_7788;
assign n_20016 = ~x_1090 & ~n_7788;
assign n_20017 = ~n_20015 & ~n_20016;
assign n_20018 =  x_1089 &  n_7821;
assign n_20019 = ~x_1089 & ~n_7821;
assign n_20020 = ~n_20018 & ~n_20019;
assign n_20021 =  x_1088 &  n_7854;
assign n_20022 = ~x_1088 & ~n_7854;
assign n_20023 = ~n_20021 & ~n_20022;
assign n_20024 =  x_1087 &  n_7887;
assign n_20025 = ~x_1087 & ~n_7887;
assign n_20026 = ~n_20024 & ~n_20025;
assign n_20027 =  x_1086 &  n_7920;
assign n_20028 = ~x_1086 & ~n_7920;
assign n_20029 = ~n_20027 & ~n_20028;
assign n_20030 =  x_1085 &  n_7953;
assign n_20031 = ~x_1085 & ~n_7953;
assign n_20032 = ~n_20030 & ~n_20031;
assign n_20033 =  x_1084 &  n_7986;
assign n_20034 = ~x_1084 & ~n_7986;
assign n_20035 = ~n_20033 & ~n_20034;
assign n_20036 =  x_1083 & ~n_17789;
assign n_20037 =  x_1732 &  x_1779;
assign n_20038 =  n_17789 &  n_20037;
assign n_20039 = ~n_20036 & ~n_20038;
assign n_20040 =  x_1083 & ~n_20039;
assign n_20041 = ~x_1083 &  n_20039;
assign n_20042 = ~n_20040 & ~n_20041;
assign n_20043 =  x_1082 & ~n_17807;
assign n_20044 =  n_17807 &  n_20037;
assign n_20045 = ~n_20043 & ~n_20044;
assign n_20046 =  x_1082 & ~n_20045;
assign n_20047 = ~x_1082 &  n_20045;
assign n_20048 = ~n_20046 & ~n_20047;
assign n_20049 =  x_1081 & ~n_17815;
assign n_20050 =  n_17815 &  n_20037;
assign n_20051 = ~n_20049 & ~n_20050;
assign n_20052 =  x_1081 & ~n_20051;
assign n_20053 = ~x_1081 &  n_20051;
assign n_20054 = ~n_20052 & ~n_20053;
assign n_20055 =  x_1080 & ~n_17823;
assign n_20056 =  n_17823 &  n_20037;
assign n_20057 = ~n_20055 & ~n_20056;
assign n_20058 =  x_1080 & ~n_20057;
assign n_20059 = ~x_1080 &  n_20057;
assign n_20060 = ~n_20058 & ~n_20059;
assign n_20061 =  x_1079 & ~n_17830;
assign n_20062 =  n_17830 &  n_20037;
assign n_20063 = ~n_20061 & ~n_20062;
assign n_20064 =  x_1079 & ~n_20063;
assign n_20065 = ~x_1079 &  n_20063;
assign n_20066 = ~n_20064 & ~n_20065;
assign n_20067 =  x_1078 & ~n_17837;
assign n_20068 =  n_17837 &  n_20037;
assign n_20069 = ~n_20067 & ~n_20068;
assign n_20070 =  x_1078 & ~n_20069;
assign n_20071 = ~x_1078 &  n_20069;
assign n_20072 = ~n_20070 & ~n_20071;
assign n_20073 =  x_1077 & ~n_17844;
assign n_20074 =  n_17844 &  n_20037;
assign n_20075 = ~n_20073 & ~n_20074;
assign n_20076 =  x_1077 & ~n_20075;
assign n_20077 = ~x_1077 &  n_20075;
assign n_20078 = ~n_20076 & ~n_20077;
assign n_20079 =  x_1076 & ~n_17851;
assign n_20080 =  n_17851 &  n_20037;
assign n_20081 = ~n_20079 & ~n_20080;
assign n_20082 =  x_1076 & ~n_20081;
assign n_20083 = ~x_1076 &  n_20081;
assign n_20084 = ~n_20082 & ~n_20083;
assign n_20085 =  x_1075 &  n_8020;
assign n_20086 = ~x_1075 & ~n_8020;
assign n_20087 = ~n_20085 & ~n_20086;
assign n_20088 =  x_1074 & ~n_17789;
assign n_20089 =  x_1732 &  x_1778;
assign n_20090 =  n_17789 &  n_20089;
assign n_20091 = ~n_20088 & ~n_20090;
assign n_20092 =  x_1074 & ~n_20091;
assign n_20093 = ~x_1074 &  n_20091;
assign n_20094 = ~n_20092 & ~n_20093;
assign n_20095 =  x_1073 & ~n_17807;
assign n_20096 =  n_17807 &  n_20089;
assign n_20097 = ~n_20095 & ~n_20096;
assign n_20098 =  x_1073 & ~n_20097;
assign n_20099 = ~x_1073 &  n_20097;
assign n_20100 = ~n_20098 & ~n_20099;
assign n_20101 =  x_1072 & ~n_17815;
assign n_20102 =  n_17815 &  n_20089;
assign n_20103 = ~n_20101 & ~n_20102;
assign n_20104 =  x_1072 & ~n_20103;
assign n_20105 = ~x_1072 &  n_20103;
assign n_20106 = ~n_20104 & ~n_20105;
assign n_20107 =  x_1071 & ~n_17823;
assign n_20108 =  n_17823 &  n_20089;
assign n_20109 = ~n_20107 & ~n_20108;
assign n_20110 =  x_1071 & ~n_20109;
assign n_20111 = ~x_1071 &  n_20109;
assign n_20112 = ~n_20110 & ~n_20111;
assign n_20113 =  x_1070 & ~n_17830;
assign n_20114 =  n_17830 &  n_20089;
assign n_20115 = ~n_20113 & ~n_20114;
assign n_20116 =  x_1070 & ~n_20115;
assign n_20117 = ~x_1070 &  n_20115;
assign n_20118 = ~n_20116 & ~n_20117;
assign n_20119 =  x_1069 & ~n_17837;
assign n_20120 =  n_17837 &  n_20089;
assign n_20121 = ~n_20119 & ~n_20120;
assign n_20122 =  x_1069 & ~n_20121;
assign n_20123 = ~x_1069 &  n_20121;
assign n_20124 = ~n_20122 & ~n_20123;
assign n_20125 =  x_1068 & ~n_17844;
assign n_20126 =  n_17844 &  n_20089;
assign n_20127 = ~n_20125 & ~n_20126;
assign n_20128 =  x_1068 & ~n_20127;
assign n_20129 = ~x_1068 &  n_20127;
assign n_20130 = ~n_20128 & ~n_20129;
assign n_20131 =  x_1067 & ~n_17851;
assign n_20132 =  n_17851 &  n_20089;
assign n_20133 = ~n_20131 & ~n_20132;
assign n_20134 =  x_1067 & ~n_20133;
assign n_20135 = ~x_1067 &  n_20133;
assign n_20136 = ~n_20134 & ~n_20135;
assign n_20137 =  x_1066 &  n_8053;
assign n_20138 = ~x_1066 & ~n_8053;
assign n_20139 = ~n_20137 & ~n_20138;
assign n_20140 =  x_1065 & ~n_17789;
assign n_20141 =  x_1732 &  x_1777;
assign n_20142 =  n_17789 &  n_20141;
assign n_20143 = ~n_20140 & ~n_20142;
assign n_20144 =  x_1065 & ~n_20143;
assign n_20145 = ~x_1065 &  n_20143;
assign n_20146 = ~n_20144 & ~n_20145;
assign n_20147 =  x_1064 & ~n_17807;
assign n_20148 =  n_17807 &  n_20141;
assign n_20149 = ~n_20147 & ~n_20148;
assign n_20150 =  x_1064 & ~n_20149;
assign n_20151 = ~x_1064 &  n_20149;
assign n_20152 = ~n_20150 & ~n_20151;
assign n_20153 =  x_1063 & ~n_17815;
assign n_20154 =  n_17815 &  n_20141;
assign n_20155 = ~n_20153 & ~n_20154;
assign n_20156 =  x_1063 & ~n_20155;
assign n_20157 = ~x_1063 &  n_20155;
assign n_20158 = ~n_20156 & ~n_20157;
assign n_20159 =  x_1062 & ~n_17823;
assign n_20160 =  n_17823 &  n_20141;
assign n_20161 = ~n_20159 & ~n_20160;
assign n_20162 =  x_1062 & ~n_20161;
assign n_20163 = ~x_1062 &  n_20161;
assign n_20164 = ~n_20162 & ~n_20163;
assign n_20165 =  x_1061 & ~n_17830;
assign n_20166 =  n_17830 &  n_20141;
assign n_20167 = ~n_20165 & ~n_20166;
assign n_20168 =  x_1061 & ~n_20167;
assign n_20169 = ~x_1061 &  n_20167;
assign n_20170 = ~n_20168 & ~n_20169;
assign n_20171 =  x_1060 & ~n_17837;
assign n_20172 =  n_17837 &  n_20141;
assign n_20173 = ~n_20171 & ~n_20172;
assign n_20174 =  x_1060 & ~n_20173;
assign n_20175 = ~x_1060 &  n_20173;
assign n_20176 = ~n_20174 & ~n_20175;
assign n_20177 =  x_1059 & ~n_17844;
assign n_20178 =  n_17844 &  n_20141;
assign n_20179 = ~n_20177 & ~n_20178;
assign n_20180 =  x_1059 & ~n_20179;
assign n_20181 = ~x_1059 &  n_20179;
assign n_20182 = ~n_20180 & ~n_20181;
assign n_20183 =  x_1058 & ~n_17851;
assign n_20184 =  n_17851 &  n_20141;
assign n_20185 = ~n_20183 & ~n_20184;
assign n_20186 =  x_1058 & ~n_20185;
assign n_20187 = ~x_1058 &  n_20185;
assign n_20188 = ~n_20186 & ~n_20187;
assign n_20189 =  x_1057 &  n_8086;
assign n_20190 = ~x_1057 & ~n_8086;
assign n_20191 = ~n_20189 & ~n_20190;
assign n_20192 =  x_1056 & ~n_17789;
assign n_20193 =  x_1732 &  x_1776;
assign n_20194 =  n_17789 &  n_20193;
assign n_20195 = ~n_20192 & ~n_20194;
assign n_20196 =  x_1056 & ~n_20195;
assign n_20197 = ~x_1056 &  n_20195;
assign n_20198 = ~n_20196 & ~n_20197;
assign n_20199 =  x_1055 & ~n_17807;
assign n_20200 =  n_17807 &  n_20193;
assign n_20201 = ~n_20199 & ~n_20200;
assign n_20202 =  x_1055 & ~n_20201;
assign n_20203 = ~x_1055 &  n_20201;
assign n_20204 = ~n_20202 & ~n_20203;
assign n_20205 =  x_1054 & ~n_17815;
assign n_20206 =  n_17815 &  n_20193;
assign n_20207 = ~n_20205 & ~n_20206;
assign n_20208 =  x_1054 & ~n_20207;
assign n_20209 = ~x_1054 &  n_20207;
assign n_20210 = ~n_20208 & ~n_20209;
assign n_20211 =  x_1053 & ~n_17823;
assign n_20212 =  n_17823 &  n_20193;
assign n_20213 = ~n_20211 & ~n_20212;
assign n_20214 =  x_1053 & ~n_20213;
assign n_20215 = ~x_1053 &  n_20213;
assign n_20216 = ~n_20214 & ~n_20215;
assign n_20217 =  x_1052 & ~n_17830;
assign n_20218 =  n_17830 &  n_20193;
assign n_20219 = ~n_20217 & ~n_20218;
assign n_20220 =  x_1052 & ~n_20219;
assign n_20221 = ~x_1052 &  n_20219;
assign n_20222 = ~n_20220 & ~n_20221;
assign n_20223 =  x_1051 & ~n_17837;
assign n_20224 =  n_17837 &  n_20193;
assign n_20225 = ~n_20223 & ~n_20224;
assign n_20226 =  x_1051 & ~n_20225;
assign n_20227 = ~x_1051 &  n_20225;
assign n_20228 = ~n_20226 & ~n_20227;
assign n_20229 =  x_1050 & ~n_17844;
assign n_20230 =  n_17844 &  n_20193;
assign n_20231 = ~n_20229 & ~n_20230;
assign n_20232 =  x_1050 & ~n_20231;
assign n_20233 = ~x_1050 &  n_20231;
assign n_20234 = ~n_20232 & ~n_20233;
assign n_20235 =  x_1049 & ~n_17851;
assign n_20236 =  n_17851 &  n_20193;
assign n_20237 = ~n_20235 & ~n_20236;
assign n_20238 =  x_1049 & ~n_20237;
assign n_20239 = ~x_1049 &  n_20237;
assign n_20240 = ~n_20238 & ~n_20239;
assign n_20241 =  x_1048 &  n_8119;
assign n_20242 = ~x_1048 & ~n_8119;
assign n_20243 = ~n_20241 & ~n_20242;
assign n_20244 =  x_1047 & ~n_17789;
assign n_20245 =  x_1732 &  x_1775;
assign n_20246 =  n_17789 &  n_20245;
assign n_20247 = ~n_20244 & ~n_20246;
assign n_20248 =  x_1047 & ~n_20247;
assign n_20249 = ~x_1047 &  n_20247;
assign n_20250 = ~n_20248 & ~n_20249;
assign n_20251 =  x_1046 & ~n_17807;
assign n_20252 =  n_17807 &  n_20245;
assign n_20253 = ~n_20251 & ~n_20252;
assign n_20254 =  x_1046 & ~n_20253;
assign n_20255 = ~x_1046 &  n_20253;
assign n_20256 = ~n_20254 & ~n_20255;
assign n_20257 =  x_1045 & ~n_17815;
assign n_20258 =  n_17815 &  n_20245;
assign n_20259 = ~n_20257 & ~n_20258;
assign n_20260 =  x_1045 & ~n_20259;
assign n_20261 = ~x_1045 &  n_20259;
assign n_20262 = ~n_20260 & ~n_20261;
assign n_20263 =  x_1044 & ~n_17823;
assign n_20264 =  n_17823 &  n_20245;
assign n_20265 = ~n_20263 & ~n_20264;
assign n_20266 =  x_1044 & ~n_20265;
assign n_20267 = ~x_1044 &  n_20265;
assign n_20268 = ~n_20266 & ~n_20267;
assign n_20269 =  x_1043 & ~n_17830;
assign n_20270 =  n_17830 &  n_20245;
assign n_20271 = ~n_20269 & ~n_20270;
assign n_20272 =  x_1043 & ~n_20271;
assign n_20273 = ~x_1043 &  n_20271;
assign n_20274 = ~n_20272 & ~n_20273;
assign n_20275 =  x_1042 & ~n_17837;
assign n_20276 =  n_17837 &  n_20245;
assign n_20277 = ~n_20275 & ~n_20276;
assign n_20278 =  x_1042 & ~n_20277;
assign n_20279 = ~x_1042 &  n_20277;
assign n_20280 = ~n_20278 & ~n_20279;
assign n_20281 =  x_1041 & ~n_17844;
assign n_20282 =  n_17844 &  n_20245;
assign n_20283 = ~n_20281 & ~n_20282;
assign n_20284 =  x_1041 & ~n_20283;
assign n_20285 = ~x_1041 &  n_20283;
assign n_20286 = ~n_20284 & ~n_20285;
assign n_20287 =  x_1040 & ~n_17851;
assign n_20288 =  n_17851 &  n_20245;
assign n_20289 = ~n_20287 & ~n_20288;
assign n_20290 =  x_1040 & ~n_20289;
assign n_20291 = ~x_1040 &  n_20289;
assign n_20292 = ~n_20290 & ~n_20291;
assign n_20293 =  x_1039 &  n_8152;
assign n_20294 = ~x_1039 & ~n_8152;
assign n_20295 = ~n_20293 & ~n_20294;
assign n_20296 =  x_1038 & ~n_17789;
assign n_20297 =  x_1732 &  x_1774;
assign n_20298 =  n_17789 &  n_20297;
assign n_20299 = ~n_20296 & ~n_20298;
assign n_20300 =  x_1038 & ~n_20299;
assign n_20301 = ~x_1038 &  n_20299;
assign n_20302 = ~n_20300 & ~n_20301;
assign n_20303 =  x_1037 & ~n_17807;
assign n_20304 =  n_17807 &  n_20297;
assign n_20305 = ~n_20303 & ~n_20304;
assign n_20306 =  x_1037 & ~n_20305;
assign n_20307 = ~x_1037 &  n_20305;
assign n_20308 = ~n_20306 & ~n_20307;
assign n_20309 =  x_1036 & ~n_17815;
assign n_20310 =  n_17815 &  n_20297;
assign n_20311 = ~n_20309 & ~n_20310;
assign n_20312 =  x_1036 & ~n_20311;
assign n_20313 = ~x_1036 &  n_20311;
assign n_20314 = ~n_20312 & ~n_20313;
assign n_20315 =  x_1035 & ~n_17823;
assign n_20316 =  n_17823 &  n_20297;
assign n_20317 = ~n_20315 & ~n_20316;
assign n_20318 =  x_1035 & ~n_20317;
assign n_20319 = ~x_1035 &  n_20317;
assign n_20320 = ~n_20318 & ~n_20319;
assign n_20321 =  x_1034 & ~n_17830;
assign n_20322 =  n_17830 &  n_20297;
assign n_20323 = ~n_20321 & ~n_20322;
assign n_20324 =  x_1034 & ~n_20323;
assign n_20325 = ~x_1034 &  n_20323;
assign n_20326 = ~n_20324 & ~n_20325;
assign n_20327 =  x_1033 & ~n_17837;
assign n_20328 =  n_17837 &  n_20297;
assign n_20329 = ~n_20327 & ~n_20328;
assign n_20330 =  x_1033 & ~n_20329;
assign n_20331 = ~x_1033 &  n_20329;
assign n_20332 = ~n_20330 & ~n_20331;
assign n_20333 =  x_1032 & ~n_17844;
assign n_20334 =  n_17844 &  n_20297;
assign n_20335 = ~n_20333 & ~n_20334;
assign n_20336 =  x_1032 & ~n_20335;
assign n_20337 = ~x_1032 &  n_20335;
assign n_20338 = ~n_20336 & ~n_20337;
assign n_20339 =  x_1031 & ~n_17851;
assign n_20340 =  n_17851 &  n_20297;
assign n_20341 = ~n_20339 & ~n_20340;
assign n_20342 =  x_1031 & ~n_20341;
assign n_20343 = ~x_1031 &  n_20341;
assign n_20344 = ~n_20342 & ~n_20343;
assign n_20345 =  x_1030 &  n_8185;
assign n_20346 = ~x_1030 & ~n_8185;
assign n_20347 = ~n_20345 & ~n_20346;
assign n_20348 =  x_1029 & ~n_17789;
assign n_20349 =  x_1732 &  x_1773;
assign n_20350 =  n_17789 &  n_20349;
assign n_20351 = ~n_20348 & ~n_20350;
assign n_20352 =  x_1029 & ~n_20351;
assign n_20353 = ~x_1029 &  n_20351;
assign n_20354 = ~n_20352 & ~n_20353;
assign n_20355 =  x_1028 & ~n_17807;
assign n_20356 =  n_17807 &  n_20349;
assign n_20357 = ~n_20355 & ~n_20356;
assign n_20358 =  x_1028 & ~n_20357;
assign n_20359 = ~x_1028 &  n_20357;
assign n_20360 = ~n_20358 & ~n_20359;
assign n_20361 =  x_1027 & ~n_17815;
assign n_20362 =  n_17815 &  n_20349;
assign n_20363 = ~n_20361 & ~n_20362;
assign n_20364 =  x_1027 & ~n_20363;
assign n_20365 = ~x_1027 &  n_20363;
assign n_20366 = ~n_20364 & ~n_20365;
assign n_20367 =  x_1026 & ~n_17823;
assign n_20368 =  n_17823 &  n_20349;
assign n_20369 = ~n_20367 & ~n_20368;
assign n_20370 =  x_1026 & ~n_20369;
assign n_20371 = ~x_1026 &  n_20369;
assign n_20372 = ~n_20370 & ~n_20371;
assign n_20373 =  x_1025 & ~n_17830;
assign n_20374 =  n_17830 &  n_20349;
assign n_20375 = ~n_20373 & ~n_20374;
assign n_20376 =  x_1025 & ~n_20375;
assign n_20377 = ~x_1025 &  n_20375;
assign n_20378 = ~n_20376 & ~n_20377;
assign n_20379 =  x_1024 & ~n_17837;
assign n_20380 =  n_17837 &  n_20349;
assign n_20381 = ~n_20379 & ~n_20380;
assign n_20382 =  x_1024 & ~n_20381;
assign n_20383 = ~x_1024 &  n_20381;
assign n_20384 = ~n_20382 & ~n_20383;
assign n_20385 =  x_1023 & ~n_17844;
assign n_20386 =  n_17844 &  n_20349;
assign n_20387 = ~n_20385 & ~n_20386;
assign n_20388 =  x_1023 & ~n_20387;
assign n_20389 = ~x_1023 &  n_20387;
assign n_20390 = ~n_20388 & ~n_20389;
assign n_20391 =  x_1022 & ~n_17851;
assign n_20392 =  n_17851 &  n_20349;
assign n_20393 = ~n_20391 & ~n_20392;
assign n_20394 =  x_1022 & ~n_20393;
assign n_20395 = ~x_1022 &  n_20393;
assign n_20396 = ~n_20394 & ~n_20395;
assign n_20397 =  x_1021 & ~n_17789;
assign n_20398 =  x_1732 &  x_1772;
assign n_20399 =  n_17789 &  n_20398;
assign n_20400 = ~n_20397 & ~n_20399;
assign n_20401 =  x_1021 & ~n_20400;
assign n_20402 = ~x_1021 &  n_20400;
assign n_20403 = ~n_20401 & ~n_20402;
assign n_20404 =  x_1020 & ~n_17807;
assign n_20405 =  n_17807 &  n_20398;
assign n_20406 = ~n_20404 & ~n_20405;
assign n_20407 =  x_1020 & ~n_20406;
assign n_20408 = ~x_1020 &  n_20406;
assign n_20409 = ~n_20407 & ~n_20408;
assign n_20410 =  x_1019 & ~n_17815;
assign n_20411 =  n_17815 &  n_20398;
assign n_20412 = ~n_20410 & ~n_20411;
assign n_20413 =  x_1019 & ~n_20412;
assign n_20414 = ~x_1019 &  n_20412;
assign n_20415 = ~n_20413 & ~n_20414;
assign n_20416 =  x_1018 & ~n_17823;
assign n_20417 =  n_17823 &  n_20398;
assign n_20418 = ~n_20416 & ~n_20417;
assign n_20419 =  x_1018 & ~n_20418;
assign n_20420 = ~x_1018 &  n_20418;
assign n_20421 = ~n_20419 & ~n_20420;
assign n_20422 =  x_1017 & ~n_17830;
assign n_20423 =  n_17830 &  n_20398;
assign n_20424 = ~n_20422 & ~n_20423;
assign n_20425 =  x_1017 & ~n_20424;
assign n_20426 = ~x_1017 &  n_20424;
assign n_20427 = ~n_20425 & ~n_20426;
assign n_20428 =  x_1016 & ~n_17837;
assign n_20429 =  n_17837 &  n_20398;
assign n_20430 = ~n_20428 & ~n_20429;
assign n_20431 =  x_1016 & ~n_20430;
assign n_20432 = ~x_1016 &  n_20430;
assign n_20433 = ~n_20431 & ~n_20432;
assign n_20434 =  x_1015 & ~n_17844;
assign n_20435 =  n_17844 &  n_20398;
assign n_20436 = ~n_20434 & ~n_20435;
assign n_20437 =  x_1015 & ~n_20436;
assign n_20438 = ~x_1015 &  n_20436;
assign n_20439 = ~n_20437 & ~n_20438;
assign n_20440 =  x_1014 & ~n_17851;
assign n_20441 =  n_17851 &  n_20398;
assign n_20442 = ~n_20440 & ~n_20441;
assign n_20443 =  x_1014 & ~n_20442;
assign n_20444 = ~x_1014 &  n_20442;
assign n_20445 = ~n_20443 & ~n_20444;
assign n_20446 = ~x_1013 & ~x_1618;
assign n_20447 =  x_1618 & ~x_1812;
assign n_20448 = ~n_20446 & ~n_20447;
assign n_20449 =  x_1013 &  n_20448;
assign n_20450 = ~x_1013 & ~n_20448;
assign n_20451 = ~n_20449 & ~n_20450;
assign n_20452 = ~x_1012 & ~x_1618;
assign n_20453 =  x_1618 & ~x_1845;
assign n_20454 = ~n_20452 & ~n_20453;
assign n_20455 =  x_1012 &  n_20454;
assign n_20456 = ~x_1012 & ~n_20454;
assign n_20457 = ~n_20455 & ~n_20456;
assign n_20458 = ~x_1011 & ~x_1618;
assign n_20459 =  x_1618 & ~x_1811;
assign n_20460 = ~n_20458 & ~n_20459;
assign n_20461 =  x_1011 &  n_20460;
assign n_20462 = ~x_1011 & ~n_20460;
assign n_20463 = ~n_20461 & ~n_20462;
assign n_20464 = ~x_1010 & ~x_1618;
assign n_20465 =  x_1618 & ~x_1844;
assign n_20466 = ~n_20464 & ~n_20465;
assign n_20467 =  x_1010 &  n_20466;
assign n_20468 = ~x_1010 & ~n_20466;
assign n_20469 = ~n_20467 & ~n_20468;
assign n_20470 = ~x_1009 & ~x_1618;
assign n_20471 =  x_1618 & ~x_1810;
assign n_20472 = ~n_20470 & ~n_20471;
assign n_20473 =  x_1009 &  n_20472;
assign n_20474 = ~x_1009 & ~n_20472;
assign n_20475 = ~n_20473 & ~n_20474;
assign n_20476 = ~x_1008 & ~x_1618;
assign n_20477 =  x_1618 & ~x_1843;
assign n_20478 = ~n_20476 & ~n_20477;
assign n_20479 =  x_1008 &  n_20478;
assign n_20480 = ~x_1008 & ~n_20478;
assign n_20481 = ~n_20479 & ~n_20480;
assign n_20482 = ~x_1007 & ~x_1618;
assign n_20483 =  x_1618 & ~x_1809;
assign n_20484 = ~n_20482 & ~n_20483;
assign n_20485 =  x_1007 &  n_20484;
assign n_20486 = ~x_1007 & ~n_20484;
assign n_20487 = ~n_20485 & ~n_20486;
assign n_20488 = ~x_1006 & ~x_1618;
assign n_20489 =  x_1618 & ~x_1842;
assign n_20490 = ~n_20488 & ~n_20489;
assign n_20491 =  x_1006 &  n_20490;
assign n_20492 = ~x_1006 & ~n_20490;
assign n_20493 = ~n_20491 & ~n_20492;
assign n_20494 = ~x_1005 & ~x_1618;
assign n_20495 =  x_1618 & ~x_1808;
assign n_20496 = ~n_20494 & ~n_20495;
assign n_20497 =  x_1005 &  n_20496;
assign n_20498 = ~x_1005 & ~n_20496;
assign n_20499 = ~n_20497 & ~n_20498;
assign n_20500 = ~x_1004 & ~x_1618;
assign n_20501 =  x_1618 & ~x_1841;
assign n_20502 = ~n_20500 & ~n_20501;
assign n_20503 =  x_1004 &  n_20502;
assign n_20504 = ~x_1004 & ~n_20502;
assign n_20505 = ~n_20503 & ~n_20504;
assign n_20506 = ~x_1003 & ~x_1618;
assign n_20507 =  x_1618 & ~x_1807;
assign n_20508 = ~n_20506 & ~n_20507;
assign n_20509 =  x_1003 &  n_20508;
assign n_20510 = ~x_1003 & ~n_20508;
assign n_20511 = ~n_20509 & ~n_20510;
assign n_20512 = ~x_1002 & ~x_1618;
assign n_20513 =  x_1618 & ~x_1840;
assign n_20514 = ~n_20512 & ~n_20513;
assign n_20515 =  x_1002 &  n_20514;
assign n_20516 = ~x_1002 & ~n_20514;
assign n_20517 = ~n_20515 & ~n_20516;
assign n_20518 = ~x_1001 & ~x_1618;
assign n_20519 =  x_1618 & ~x_1806;
assign n_20520 = ~n_20518 & ~n_20519;
assign n_20521 =  x_1001 &  n_20520;
assign n_20522 = ~x_1001 & ~n_20520;
assign n_20523 = ~n_20521 & ~n_20522;
assign n_20524 = ~x_1000 & ~x_1618;
assign n_20525 =  x_1618 & ~x_1839;
assign n_20526 = ~n_20524 & ~n_20525;
assign n_20527 =  x_1000 &  n_20526;
assign n_20528 = ~x_1000 & ~n_20526;
assign n_20529 = ~n_20527 & ~n_20528;
assign n_20530 = ~x_999 & ~x_1618;
assign n_20531 =  x_1618 & ~x_1805;
assign n_20532 = ~n_20530 & ~n_20531;
assign n_20533 =  x_999 &  n_20532;
assign n_20534 = ~x_999 & ~n_20532;
assign n_20535 = ~n_20533 & ~n_20534;
assign n_20536 = ~x_998 & ~x_1618;
assign n_20537 =  x_1618 & ~x_1838;
assign n_20538 = ~n_20536 & ~n_20537;
assign n_20539 =  x_998 &  n_20538;
assign n_20540 = ~x_998 & ~n_20538;
assign n_20541 = ~n_20539 & ~n_20540;
assign n_20542 = ~x_997 & ~x_1618;
assign n_20543 =  x_1618 & ~x_1804;
assign n_20544 = ~n_20542 & ~n_20543;
assign n_20545 =  x_997 &  n_20544;
assign n_20546 = ~x_997 & ~n_20544;
assign n_20547 = ~n_20545 & ~n_20546;
assign n_20548 = ~x_996 & ~x_1618;
assign n_20549 =  x_1618 & ~x_1837;
assign n_20550 = ~n_20548 & ~n_20549;
assign n_20551 =  x_996 &  n_20550;
assign n_20552 = ~x_996 & ~n_20550;
assign n_20553 = ~n_20551 & ~n_20552;
assign n_20554 = ~x_995 & ~x_1618;
assign n_20555 =  x_1618 & ~x_1803;
assign n_20556 = ~n_20554 & ~n_20555;
assign n_20557 =  x_995 &  n_20556;
assign n_20558 = ~x_995 & ~n_20556;
assign n_20559 = ~n_20557 & ~n_20558;
assign n_20560 = ~x_994 & ~x_1618;
assign n_20561 =  x_1618 & ~x_1836;
assign n_20562 = ~n_20560 & ~n_20561;
assign n_20563 =  x_994 &  n_20562;
assign n_20564 = ~x_994 & ~n_20562;
assign n_20565 = ~n_20563 & ~n_20564;
assign n_20566 = ~x_993 & ~x_1618;
assign n_20567 =  x_1618 & ~x_1802;
assign n_20568 = ~n_20566 & ~n_20567;
assign n_20569 =  x_993 &  n_20568;
assign n_20570 = ~x_993 & ~n_20568;
assign n_20571 = ~n_20569 & ~n_20570;
assign n_20572 = ~x_992 & ~x_1618;
assign n_20573 =  x_1618 & ~x_1835;
assign n_20574 = ~n_20572 & ~n_20573;
assign n_20575 =  x_992 &  n_20574;
assign n_20576 = ~x_992 & ~n_20574;
assign n_20577 = ~n_20575 & ~n_20576;
assign n_20578 = ~x_991 & ~x_1618;
assign n_20579 =  x_1618 & ~x_1801;
assign n_20580 = ~n_20578 & ~n_20579;
assign n_20581 =  x_991 &  n_20580;
assign n_20582 = ~x_991 & ~n_20580;
assign n_20583 = ~n_20581 & ~n_20582;
assign n_20584 = ~x_990 & ~x_1618;
assign n_20585 =  x_1618 & ~x_1834;
assign n_20586 = ~n_20584 & ~n_20585;
assign n_20587 =  x_990 &  n_20586;
assign n_20588 = ~x_990 & ~n_20586;
assign n_20589 = ~n_20587 & ~n_20588;
assign n_20590 = ~x_989 & ~x_1618;
assign n_20591 =  x_1618 & ~x_1800;
assign n_20592 = ~n_20590 & ~n_20591;
assign n_20593 =  x_989 &  n_20592;
assign n_20594 = ~x_989 & ~n_20592;
assign n_20595 = ~n_20593 & ~n_20594;
assign n_20596 = ~x_988 & ~x_1618;
assign n_20597 =  x_1618 & ~x_1833;
assign n_20598 = ~n_20596 & ~n_20597;
assign n_20599 =  x_988 &  n_20598;
assign n_20600 = ~x_988 & ~n_20598;
assign n_20601 = ~n_20599 & ~n_20600;
assign n_20602 = ~x_987 & ~x_1618;
assign n_20603 =  x_1618 & ~x_1799;
assign n_20604 = ~n_20602 & ~n_20603;
assign n_20605 =  x_987 &  n_20604;
assign n_20606 = ~x_987 & ~n_20604;
assign n_20607 = ~n_20605 & ~n_20606;
assign n_20608 = ~x_986 & ~x_1618;
assign n_20609 =  x_1618 & ~x_1832;
assign n_20610 = ~n_20608 & ~n_20609;
assign n_20611 =  x_986 &  n_20610;
assign n_20612 = ~x_986 & ~n_20610;
assign n_20613 = ~n_20611 & ~n_20612;
assign n_20614 = ~x_985 & ~x_1618;
assign n_20615 =  x_1618 & ~x_1798;
assign n_20616 = ~n_20614 & ~n_20615;
assign n_20617 =  x_985 &  n_20616;
assign n_20618 = ~x_985 & ~n_20616;
assign n_20619 = ~n_20617 & ~n_20618;
assign n_20620 = ~x_984 & ~x_1618;
assign n_20621 =  x_1618 & ~x_1831;
assign n_20622 = ~n_20620 & ~n_20621;
assign n_20623 =  x_984 &  n_20622;
assign n_20624 = ~x_984 & ~n_20622;
assign n_20625 = ~n_20623 & ~n_20624;
assign n_20626 = ~x_983 & ~x_1618;
assign n_20627 =  x_1618 & ~x_1797;
assign n_20628 = ~n_20626 & ~n_20627;
assign n_20629 =  x_983 &  n_20628;
assign n_20630 = ~x_983 & ~n_20628;
assign n_20631 = ~n_20629 & ~n_20630;
assign n_20632 = ~x_982 & ~x_1618;
assign n_20633 =  x_1618 & ~x_1830;
assign n_20634 = ~n_20632 & ~n_20633;
assign n_20635 =  x_982 &  n_20634;
assign n_20636 = ~x_982 & ~n_20634;
assign n_20637 = ~n_20635 & ~n_20636;
assign n_20638 = ~x_981 & ~x_1618;
assign n_20639 =  x_1618 & ~x_1796;
assign n_20640 = ~n_20638 & ~n_20639;
assign n_20641 =  x_981 &  n_20640;
assign n_20642 = ~x_981 & ~n_20640;
assign n_20643 = ~n_20641 & ~n_20642;
assign n_20644 = ~x_980 & ~x_1618;
assign n_20645 =  x_1618 & ~x_1829;
assign n_20646 = ~n_20644 & ~n_20645;
assign n_20647 =  x_980 &  n_20646;
assign n_20648 = ~x_980 & ~n_20646;
assign n_20649 = ~n_20647 & ~n_20648;
assign n_20650 = ~x_979 & ~x_1618;
assign n_20651 =  x_1618 & ~x_1795;
assign n_20652 = ~n_20650 & ~n_20651;
assign n_20653 =  x_979 &  n_20652;
assign n_20654 = ~x_979 & ~n_20652;
assign n_20655 = ~n_20653 & ~n_20654;
assign n_20656 = ~x_978 & ~x_1618;
assign n_20657 =  x_1618 & ~x_1828;
assign n_20658 = ~n_20656 & ~n_20657;
assign n_20659 =  x_978 &  n_20658;
assign n_20660 = ~x_978 & ~n_20658;
assign n_20661 = ~n_20659 & ~n_20660;
assign n_20662 = ~x_977 & ~x_1618;
assign n_20663 =  x_1618 & ~x_1794;
assign n_20664 = ~n_20662 & ~n_20663;
assign n_20665 =  x_977 &  n_20664;
assign n_20666 = ~x_977 & ~n_20664;
assign n_20667 = ~n_20665 & ~n_20666;
assign n_20668 = ~x_976 & ~x_1618;
assign n_20669 =  x_1618 & ~x_1827;
assign n_20670 = ~n_20668 & ~n_20669;
assign n_20671 =  x_976 &  n_20670;
assign n_20672 = ~x_976 & ~n_20670;
assign n_20673 = ~n_20671 & ~n_20672;
assign n_20674 = ~x_975 & ~x_1618;
assign n_20675 =  x_1618 & ~x_1793;
assign n_20676 = ~n_20674 & ~n_20675;
assign n_20677 =  x_975 &  n_20676;
assign n_20678 = ~x_975 & ~n_20676;
assign n_20679 = ~n_20677 & ~n_20678;
assign n_20680 = ~x_974 & ~x_1618;
assign n_20681 =  x_1618 & ~x_1826;
assign n_20682 = ~n_20680 & ~n_20681;
assign n_20683 =  x_974 &  n_20682;
assign n_20684 = ~x_974 & ~n_20682;
assign n_20685 = ~n_20683 & ~n_20684;
assign n_20686 = ~x_973 & ~x_1618;
assign n_20687 =  x_1618 & ~x_1792;
assign n_20688 = ~n_20686 & ~n_20687;
assign n_20689 =  x_973 &  n_20688;
assign n_20690 = ~x_973 & ~n_20688;
assign n_20691 = ~n_20689 & ~n_20690;
assign n_20692 = ~x_972 & ~x_1618;
assign n_20693 =  x_1618 & ~x_1825;
assign n_20694 = ~n_20692 & ~n_20693;
assign n_20695 =  x_972 &  n_20694;
assign n_20696 = ~x_972 & ~n_20694;
assign n_20697 = ~n_20695 & ~n_20696;
assign n_20698 = ~x_971 & ~x_1618;
assign n_20699 =  x_1618 & ~x_1791;
assign n_20700 = ~n_20698 & ~n_20699;
assign n_20701 =  x_971 &  n_20700;
assign n_20702 = ~x_971 & ~n_20700;
assign n_20703 = ~n_20701 & ~n_20702;
assign n_20704 = ~x_970 & ~x_1618;
assign n_20705 =  x_1618 & ~x_1824;
assign n_20706 = ~n_20704 & ~n_20705;
assign n_20707 =  x_970 &  n_20706;
assign n_20708 = ~x_970 & ~n_20706;
assign n_20709 = ~n_20707 & ~n_20708;
assign n_20710 = ~x_969 & ~x_1618;
assign n_20711 =  x_1618 & ~x_1790;
assign n_20712 = ~n_20710 & ~n_20711;
assign n_20713 =  x_969 &  n_20712;
assign n_20714 = ~x_969 & ~n_20712;
assign n_20715 = ~n_20713 & ~n_20714;
assign n_20716 = ~x_968 & ~x_1618;
assign n_20717 =  x_1618 & ~x_1823;
assign n_20718 = ~n_20716 & ~n_20717;
assign n_20719 =  x_968 &  n_20718;
assign n_20720 = ~x_968 & ~n_20718;
assign n_20721 = ~n_20719 & ~n_20720;
assign n_20722 = ~x_967 & ~x_1618;
assign n_20723 =  x_1618 & ~x_1789;
assign n_20724 = ~n_20722 & ~n_20723;
assign n_20725 =  x_967 &  n_20724;
assign n_20726 = ~x_967 & ~n_20724;
assign n_20727 = ~n_20725 & ~n_20726;
assign n_20728 = ~x_966 & ~x_1618;
assign n_20729 =  x_1618 & ~x_1822;
assign n_20730 = ~n_20728 & ~n_20729;
assign n_20731 =  x_966 &  n_20730;
assign n_20732 = ~x_966 & ~n_20730;
assign n_20733 = ~n_20731 & ~n_20732;
assign n_20734 = ~x_965 & ~x_1618;
assign n_20735 =  x_1618 & ~x_1788;
assign n_20736 = ~n_20734 & ~n_20735;
assign n_20737 =  x_965 &  n_20736;
assign n_20738 = ~x_965 & ~n_20736;
assign n_20739 = ~n_20737 & ~n_20738;
assign n_20740 = ~x_964 & ~x_1618;
assign n_20741 =  x_1618 & ~x_1821;
assign n_20742 = ~n_20740 & ~n_20741;
assign n_20743 =  x_964 &  n_20742;
assign n_20744 = ~x_964 & ~n_20742;
assign n_20745 = ~n_20743 & ~n_20744;
assign n_20746 = ~x_963 & ~x_1618;
assign n_20747 =  x_1618 & ~x_1787;
assign n_20748 = ~n_20746 & ~n_20747;
assign n_20749 =  x_963 &  n_20748;
assign n_20750 = ~x_963 & ~n_20748;
assign n_20751 = ~n_20749 & ~n_20750;
assign n_20752 = ~x_962 & ~x_1618;
assign n_20753 =  x_1618 & ~x_1820;
assign n_20754 = ~n_20752 & ~n_20753;
assign n_20755 =  x_962 &  n_20754;
assign n_20756 = ~x_962 & ~n_20754;
assign n_20757 = ~n_20755 & ~n_20756;
assign n_20758 = ~x_961 & ~x_1618;
assign n_20759 =  x_1618 & ~x_1786;
assign n_20760 = ~n_20758 & ~n_20759;
assign n_20761 =  x_961 &  n_20760;
assign n_20762 = ~x_961 & ~n_20760;
assign n_20763 = ~n_20761 & ~n_20762;
assign n_20764 = ~x_960 & ~x_1618;
assign n_20765 =  x_1618 & ~x_1819;
assign n_20766 = ~n_20764 & ~n_20765;
assign n_20767 =  x_960 &  n_20766;
assign n_20768 = ~x_960 & ~n_20766;
assign n_20769 = ~n_20767 & ~n_20768;
assign n_20770 = ~x_959 & ~x_1618;
assign n_20771 =  x_1618 & ~x_1785;
assign n_20772 = ~n_20770 & ~n_20771;
assign n_20773 =  x_959 &  n_20772;
assign n_20774 = ~x_959 & ~n_20772;
assign n_20775 = ~n_20773 & ~n_20774;
assign n_20776 = ~x_958 & ~x_1618;
assign n_20777 =  x_1618 & ~x_1818;
assign n_20778 = ~n_20776 & ~n_20777;
assign n_20779 =  x_958 &  n_20778;
assign n_20780 = ~x_958 & ~n_20778;
assign n_20781 = ~n_20779 & ~n_20780;
assign n_20782 = ~x_957 & ~x_1618;
assign n_20783 =  x_1618 & ~x_1784;
assign n_20784 = ~n_20782 & ~n_20783;
assign n_20785 =  x_957 &  n_20784;
assign n_20786 = ~x_957 & ~n_20784;
assign n_20787 = ~n_20785 & ~n_20786;
assign n_20788 = ~x_956 & ~x_1618;
assign n_20789 =  x_1618 & ~x_1817;
assign n_20790 = ~n_20788 & ~n_20789;
assign n_20791 =  x_956 &  n_20790;
assign n_20792 = ~x_956 & ~n_20790;
assign n_20793 = ~n_20791 & ~n_20792;
assign n_20794 = ~x_955 & ~x_1618;
assign n_20795 =  x_1618 & ~x_1783;
assign n_20796 = ~n_20794 & ~n_20795;
assign n_20797 =  x_955 &  n_20796;
assign n_20798 = ~x_955 & ~n_20796;
assign n_20799 = ~n_20797 & ~n_20798;
assign n_20800 = ~x_954 & ~x_1618;
assign n_20801 =  x_1618 & ~x_1816;
assign n_20802 = ~n_20800 & ~n_20801;
assign n_20803 =  x_954 &  n_20802;
assign n_20804 = ~x_954 & ~n_20802;
assign n_20805 = ~n_20803 & ~n_20804;
assign n_20806 = ~x_953 & ~x_1618;
assign n_20807 =  x_1618 & ~x_1782;
assign n_20808 = ~n_20806 & ~n_20807;
assign n_20809 =  x_953 &  n_20808;
assign n_20810 = ~x_953 & ~n_20808;
assign n_20811 = ~n_20809 & ~n_20810;
assign n_20812 = ~x_952 & ~x_1618;
assign n_20813 =  x_1618 & ~x_1815;
assign n_20814 = ~n_20812 & ~n_20813;
assign n_20815 =  x_952 &  n_20814;
assign n_20816 = ~x_952 & ~n_20814;
assign n_20817 = ~n_20815 & ~n_20816;
assign n_20818 = ~x_951 & ~x_1618;
assign n_20819 =  x_1618 & ~x_1781;
assign n_20820 = ~n_20818 & ~n_20819;
assign n_20821 =  x_951 &  n_20820;
assign n_20822 = ~x_951 & ~n_20820;
assign n_20823 = ~n_20821 & ~n_20822;
assign n_20824 = ~x_950 & ~x_1618;
assign n_20825 =  x_1618 & ~x_1814;
assign n_20826 = ~n_20824 & ~n_20825;
assign n_20827 =  x_950 &  n_20826;
assign n_20828 = ~x_950 & ~n_20826;
assign n_20829 = ~n_20827 & ~n_20828;
assign n_20830 = ~x_949 & ~x_1618;
assign n_20831 =  x_1618 & ~x_1780;
assign n_20832 = ~n_20830 & ~n_20831;
assign n_20833 =  x_949 &  n_20832;
assign n_20834 = ~x_949 & ~n_20832;
assign n_20835 = ~n_20833 & ~n_20834;
assign n_20836 = ~x_948 & ~x_1618;
assign n_20837 =  x_1618 & ~x_1813;
assign n_20838 = ~n_20836 & ~n_20837;
assign n_20839 =  x_948 &  n_20838;
assign n_20840 = ~x_948 & ~n_20838;
assign n_20841 = ~n_20839 & ~n_20840;
assign n_20842 =  x_947 & ~n_17789;
assign n_20843 =  x_1732 & ~x_1737;
assign n_20844 =  n_17789 &  n_20843;
assign n_20845 = ~n_20842 & ~n_20844;
assign n_20846 =  x_947 & ~n_20845;
assign n_20847 = ~x_947 &  n_20845;
assign n_20848 = ~n_20846 & ~n_20847;
assign n_20849 =  x_946 & ~n_17807;
assign n_20850 =  n_17807 &  n_20843;
assign n_20851 = ~n_20849 & ~n_20850;
assign n_20852 =  x_946 & ~n_20851;
assign n_20853 = ~x_946 &  n_20851;
assign n_20854 = ~n_20852 & ~n_20853;
assign n_20855 =  x_945 & ~n_17815;
assign n_20856 =  n_17815 &  n_20843;
assign n_20857 = ~n_20855 & ~n_20856;
assign n_20858 =  x_945 & ~n_20857;
assign n_20859 = ~x_945 &  n_20857;
assign n_20860 = ~n_20858 & ~n_20859;
assign n_20861 =  x_944 & ~n_17823;
assign n_20862 =  n_17823 &  n_20843;
assign n_20863 = ~n_20861 & ~n_20862;
assign n_20864 =  x_944 & ~n_20863;
assign n_20865 = ~x_944 &  n_20863;
assign n_20866 = ~n_20864 & ~n_20865;
assign n_20867 =  x_943 & ~n_17830;
assign n_20868 =  n_17830 &  n_20843;
assign n_20869 = ~n_20867 & ~n_20868;
assign n_20870 =  x_943 & ~n_20869;
assign n_20871 = ~x_943 &  n_20869;
assign n_20872 = ~n_20870 & ~n_20871;
assign n_20873 =  x_942 & ~n_17837;
assign n_20874 =  n_17837 &  n_20843;
assign n_20875 = ~n_20873 & ~n_20874;
assign n_20876 =  x_942 & ~n_20875;
assign n_20877 = ~x_942 &  n_20875;
assign n_20878 = ~n_20876 & ~n_20877;
assign n_20879 =  x_941 & ~n_17844;
assign n_20880 =  n_17844 &  n_20843;
assign n_20881 = ~n_20879 & ~n_20880;
assign n_20882 =  x_941 & ~n_20881;
assign n_20883 = ~x_941 &  n_20881;
assign n_20884 = ~n_20882 & ~n_20883;
assign n_20885 =  x_940 & ~n_17851;
assign n_20886 =  n_17851 &  n_20843;
assign n_20887 = ~n_20885 & ~n_20886;
assign n_20888 =  x_940 & ~n_20887;
assign n_20889 = ~x_940 &  n_20887;
assign n_20890 = ~n_20888 & ~n_20889;
assign n_20891 =  x_939 & ~n_17789;
assign n_20892 =  x_1732 & ~x_1741;
assign n_20893 =  n_17789 &  n_20892;
assign n_20894 = ~n_20891 & ~n_20893;
assign n_20895 =  x_939 & ~n_20894;
assign n_20896 = ~x_939 &  n_20894;
assign n_20897 = ~n_20895 & ~n_20896;
assign n_20898 =  x_938 & ~n_17807;
assign n_20899 =  n_17807 &  n_20892;
assign n_20900 = ~n_20898 & ~n_20899;
assign n_20901 =  x_938 & ~n_20900;
assign n_20902 = ~x_938 &  n_20900;
assign n_20903 = ~n_20901 & ~n_20902;
assign n_20904 =  x_937 & ~n_17815;
assign n_20905 =  n_17815 &  n_20892;
assign n_20906 = ~n_20904 & ~n_20905;
assign n_20907 =  x_937 & ~n_20906;
assign n_20908 = ~x_937 &  n_20906;
assign n_20909 = ~n_20907 & ~n_20908;
assign n_20910 =  x_936 & ~n_17823;
assign n_20911 =  n_17823 &  n_20892;
assign n_20912 = ~n_20910 & ~n_20911;
assign n_20913 =  x_936 & ~n_20912;
assign n_20914 = ~x_936 &  n_20912;
assign n_20915 = ~n_20913 & ~n_20914;
assign n_20916 =  x_935 & ~n_17830;
assign n_20917 =  n_17830 &  n_20892;
assign n_20918 = ~n_20916 & ~n_20917;
assign n_20919 =  x_935 & ~n_20918;
assign n_20920 = ~x_935 &  n_20918;
assign n_20921 = ~n_20919 & ~n_20920;
assign n_20922 =  x_934 & ~n_17837;
assign n_20923 =  n_17837 &  n_20892;
assign n_20924 = ~n_20922 & ~n_20923;
assign n_20925 =  x_934 & ~n_20924;
assign n_20926 = ~x_934 &  n_20924;
assign n_20927 = ~n_20925 & ~n_20926;
assign n_20928 =  x_933 & ~n_17844;
assign n_20929 =  n_17844 &  n_20892;
assign n_20930 = ~n_20928 & ~n_20929;
assign n_20931 =  x_933 & ~n_20930;
assign n_20932 = ~x_933 &  n_20930;
assign n_20933 = ~n_20931 & ~n_20932;
assign n_20934 =  x_932 & ~n_17851;
assign n_20935 =  n_17851 &  n_20892;
assign n_20936 = ~n_20934 & ~n_20935;
assign n_20937 =  x_932 & ~n_20936;
assign n_20938 = ~x_932 &  n_20936;
assign n_20939 = ~n_20937 & ~n_20938;
assign n_20940 =  x_931 & ~n_17789;
assign n_20941 =  x_1732 &  x_1742;
assign n_20942 =  n_17789 &  n_20941;
assign n_20943 = ~n_20940 & ~n_20942;
assign n_20944 =  x_931 & ~n_20943;
assign n_20945 = ~x_931 &  n_20943;
assign n_20946 = ~n_20944 & ~n_20945;
assign n_20947 =  x_930 & ~n_17807;
assign n_20948 =  n_17807 &  n_20941;
assign n_20949 = ~n_20947 & ~n_20948;
assign n_20950 =  x_930 & ~n_20949;
assign n_20951 = ~x_930 &  n_20949;
assign n_20952 = ~n_20950 & ~n_20951;
assign n_20953 =  x_929 & ~n_17815;
assign n_20954 =  n_17815 &  n_20941;
assign n_20955 = ~n_20953 & ~n_20954;
assign n_20956 =  x_929 & ~n_20955;
assign n_20957 = ~x_929 &  n_20955;
assign n_20958 = ~n_20956 & ~n_20957;
assign n_20959 =  x_928 & ~n_17823;
assign n_20960 =  n_17823 &  n_20941;
assign n_20961 = ~n_20959 & ~n_20960;
assign n_20962 =  x_928 & ~n_20961;
assign n_20963 = ~x_928 &  n_20961;
assign n_20964 = ~n_20962 & ~n_20963;
assign n_20965 =  x_927 & ~n_17830;
assign n_20966 =  n_17830 &  n_20941;
assign n_20967 = ~n_20965 & ~n_20966;
assign n_20968 =  x_927 & ~n_20967;
assign n_20969 = ~x_927 &  n_20967;
assign n_20970 = ~n_20968 & ~n_20969;
assign n_20971 =  x_926 & ~n_17837;
assign n_20972 =  n_17837 &  n_20941;
assign n_20973 = ~n_20971 & ~n_20972;
assign n_20974 =  x_926 & ~n_20973;
assign n_20975 = ~x_926 &  n_20973;
assign n_20976 = ~n_20974 & ~n_20975;
assign n_20977 =  x_925 & ~n_17844;
assign n_20978 =  n_17844 &  n_20941;
assign n_20979 = ~n_20977 & ~n_20978;
assign n_20980 =  x_925 & ~n_20979;
assign n_20981 = ~x_925 &  n_20979;
assign n_20982 = ~n_20980 & ~n_20981;
assign n_20983 =  x_924 & ~n_17851;
assign n_20984 =  n_17851 &  n_20941;
assign n_20985 = ~n_20983 & ~n_20984;
assign n_20986 =  x_924 & ~n_20985;
assign n_20987 = ~x_924 &  n_20985;
assign n_20988 = ~n_20986 & ~n_20987;
assign n_20989 =  x_923 & ~n_17789;
assign n_20990 =  x_1732 &  x_1740;
assign n_20991 =  n_17789 &  n_20990;
assign n_20992 = ~n_20989 & ~n_20991;
assign n_20993 =  x_923 & ~n_20992;
assign n_20994 = ~x_923 &  n_20992;
assign n_20995 = ~n_20993 & ~n_20994;
assign n_20996 =  x_922 & ~n_17807;
assign n_20997 =  n_17807 &  n_20990;
assign n_20998 = ~n_20996 & ~n_20997;
assign n_20999 =  x_922 & ~n_20998;
assign n_21000 = ~x_922 &  n_20998;
assign n_21001 = ~n_20999 & ~n_21000;
assign n_21002 =  x_921 & ~n_17815;
assign n_21003 =  n_17815 &  n_20990;
assign n_21004 = ~n_21002 & ~n_21003;
assign n_21005 =  x_921 & ~n_21004;
assign n_21006 = ~x_921 &  n_21004;
assign n_21007 = ~n_21005 & ~n_21006;
assign n_21008 =  x_920 & ~n_17823;
assign n_21009 =  n_17823 &  n_20990;
assign n_21010 = ~n_21008 & ~n_21009;
assign n_21011 =  x_920 & ~n_21010;
assign n_21012 = ~x_920 &  n_21010;
assign n_21013 = ~n_21011 & ~n_21012;
assign n_21014 =  x_919 & ~n_17830;
assign n_21015 =  n_17830 &  n_20990;
assign n_21016 = ~n_21014 & ~n_21015;
assign n_21017 =  x_919 & ~n_21016;
assign n_21018 = ~x_919 &  n_21016;
assign n_21019 = ~n_21017 & ~n_21018;
assign n_21020 =  x_918 & ~n_17837;
assign n_21021 =  n_17837 &  n_20990;
assign n_21022 = ~n_21020 & ~n_21021;
assign n_21023 =  x_918 & ~n_21022;
assign n_21024 = ~x_918 &  n_21022;
assign n_21025 = ~n_21023 & ~n_21024;
assign n_21026 =  x_917 & ~n_17844;
assign n_21027 =  n_17844 &  n_20990;
assign n_21028 = ~n_21026 & ~n_21027;
assign n_21029 =  x_917 & ~n_21028;
assign n_21030 = ~x_917 &  n_21028;
assign n_21031 = ~n_21029 & ~n_21030;
assign n_21032 =  x_916 & ~n_17851;
assign n_21033 =  n_17851 &  n_20990;
assign n_21034 = ~n_21032 & ~n_21033;
assign n_21035 =  x_916 & ~n_21034;
assign n_21036 = ~x_916 &  n_21034;
assign n_21037 = ~n_21035 & ~n_21036;
assign n_21038 =  x_915 & ~n_17789;
assign n_21039 =  x_1732 & ~x_1739;
assign n_21040 =  n_17789 &  n_21039;
assign n_21041 = ~n_21038 & ~n_21040;
assign n_21042 =  x_915 & ~n_21041;
assign n_21043 = ~x_915 &  n_21041;
assign n_21044 = ~n_21042 & ~n_21043;
assign n_21045 =  x_914 & ~n_17807;
assign n_21046 =  n_17807 &  n_21039;
assign n_21047 = ~n_21045 & ~n_21046;
assign n_21048 =  x_914 & ~n_21047;
assign n_21049 = ~x_914 &  n_21047;
assign n_21050 = ~n_21048 & ~n_21049;
assign n_21051 =  x_913 & ~n_17815;
assign n_21052 =  n_17815 &  n_21039;
assign n_21053 = ~n_21051 & ~n_21052;
assign n_21054 =  x_913 & ~n_21053;
assign n_21055 = ~x_913 &  n_21053;
assign n_21056 = ~n_21054 & ~n_21055;
assign n_21057 =  x_912 & ~n_17823;
assign n_21058 =  n_17823 &  n_21039;
assign n_21059 = ~n_21057 & ~n_21058;
assign n_21060 =  x_912 & ~n_21059;
assign n_21061 = ~x_912 &  n_21059;
assign n_21062 = ~n_21060 & ~n_21061;
assign n_21063 =  x_911 & ~n_17830;
assign n_21064 =  n_17830 &  n_21039;
assign n_21065 = ~n_21063 & ~n_21064;
assign n_21066 =  x_911 & ~n_21065;
assign n_21067 = ~x_911 &  n_21065;
assign n_21068 = ~n_21066 & ~n_21067;
assign n_21069 =  x_910 & ~n_17837;
assign n_21070 =  n_17837 &  n_21039;
assign n_21071 = ~n_21069 & ~n_21070;
assign n_21072 =  x_910 & ~n_21071;
assign n_21073 = ~x_910 &  n_21071;
assign n_21074 = ~n_21072 & ~n_21073;
assign n_21075 =  x_909 & ~n_17844;
assign n_21076 =  n_17844 &  n_21039;
assign n_21077 = ~n_21075 & ~n_21076;
assign n_21078 =  x_909 & ~n_21077;
assign n_21079 = ~x_909 &  n_21077;
assign n_21080 = ~n_21078 & ~n_21079;
assign n_21081 =  x_908 & ~n_17851;
assign n_21082 =  n_17851 &  n_21039;
assign n_21083 = ~n_21081 & ~n_21082;
assign n_21084 =  x_908 & ~n_21083;
assign n_21085 = ~x_908 &  n_21083;
assign n_21086 = ~n_21084 & ~n_21085;
assign n_21087 =  x_907 & ~n_17789;
assign n_21088 =  x_1732 &  x_1743;
assign n_21089 =  n_17789 &  n_21088;
assign n_21090 = ~n_21087 & ~n_21089;
assign n_21091 =  x_907 & ~n_21090;
assign n_21092 = ~x_907 &  n_21090;
assign n_21093 = ~n_21091 & ~n_21092;
assign n_21094 =  x_906 & ~n_17807;
assign n_21095 =  n_17807 &  n_21088;
assign n_21096 = ~n_21094 & ~n_21095;
assign n_21097 =  x_906 & ~n_21096;
assign n_21098 = ~x_906 &  n_21096;
assign n_21099 = ~n_21097 & ~n_21098;
assign n_21100 =  x_905 & ~n_17815;
assign n_21101 =  n_17815 &  n_21088;
assign n_21102 = ~n_21100 & ~n_21101;
assign n_21103 =  x_905 & ~n_21102;
assign n_21104 = ~x_905 &  n_21102;
assign n_21105 = ~n_21103 & ~n_21104;
assign n_21106 =  x_904 & ~n_17823;
assign n_21107 =  n_17823 &  n_21088;
assign n_21108 = ~n_21106 & ~n_21107;
assign n_21109 =  x_904 & ~n_21108;
assign n_21110 = ~x_904 &  n_21108;
assign n_21111 = ~n_21109 & ~n_21110;
assign n_21112 =  x_903 & ~n_17830;
assign n_21113 =  n_17830 &  n_21088;
assign n_21114 = ~n_21112 & ~n_21113;
assign n_21115 =  x_903 & ~n_21114;
assign n_21116 = ~x_903 &  n_21114;
assign n_21117 = ~n_21115 & ~n_21116;
assign n_21118 =  x_902 & ~n_17837;
assign n_21119 =  n_17837 &  n_21088;
assign n_21120 = ~n_21118 & ~n_21119;
assign n_21121 =  x_902 & ~n_21120;
assign n_21122 = ~x_902 &  n_21120;
assign n_21123 = ~n_21121 & ~n_21122;
assign n_21124 =  x_901 & ~n_17844;
assign n_21125 =  n_17844 &  n_21088;
assign n_21126 = ~n_21124 & ~n_21125;
assign n_21127 =  x_901 & ~n_21126;
assign n_21128 = ~x_901 &  n_21126;
assign n_21129 = ~n_21127 & ~n_21128;
assign n_21130 =  x_900 & ~n_17851;
assign n_21131 =  n_17851 &  n_21088;
assign n_21132 = ~n_21130 & ~n_21131;
assign n_21133 =  x_900 & ~n_21132;
assign n_21134 = ~x_900 &  n_21132;
assign n_21135 = ~n_21133 & ~n_21134;
assign n_21136 =  x_899 & ~n_17789;
assign n_21137 =  x_1732 & ~x_1738;
assign n_21138 =  n_17789 &  n_21137;
assign n_21139 = ~n_21136 & ~n_21138;
assign n_21140 =  x_899 & ~n_21139;
assign n_21141 = ~x_899 &  n_21139;
assign n_21142 = ~n_21140 & ~n_21141;
assign n_21143 =  x_898 & ~n_17807;
assign n_21144 =  n_17807 &  n_21137;
assign n_21145 = ~n_21143 & ~n_21144;
assign n_21146 =  x_898 & ~n_21145;
assign n_21147 = ~x_898 &  n_21145;
assign n_21148 = ~n_21146 & ~n_21147;
assign n_21149 =  x_897 & ~n_17815;
assign n_21150 =  n_17815 &  n_21137;
assign n_21151 = ~n_21149 & ~n_21150;
assign n_21152 =  x_897 & ~n_21151;
assign n_21153 = ~x_897 &  n_21151;
assign n_21154 = ~n_21152 & ~n_21153;
assign n_21155 =  x_896 & ~n_17823;
assign n_21156 =  n_17823 &  n_21137;
assign n_21157 = ~n_21155 & ~n_21156;
assign n_21158 =  x_896 & ~n_21157;
assign n_21159 = ~x_896 &  n_21157;
assign n_21160 = ~n_21158 & ~n_21159;
assign n_21161 =  x_895 & ~n_17830;
assign n_21162 =  n_17830 &  n_21137;
assign n_21163 = ~n_21161 & ~n_21162;
assign n_21164 =  x_895 & ~n_21163;
assign n_21165 = ~x_895 &  n_21163;
assign n_21166 = ~n_21164 & ~n_21165;
assign n_21167 =  x_894 & ~n_17837;
assign n_21168 =  n_17837 &  n_21137;
assign n_21169 = ~n_21167 & ~n_21168;
assign n_21170 =  x_894 & ~n_21169;
assign n_21171 = ~x_894 &  n_21169;
assign n_21172 = ~n_21170 & ~n_21171;
assign n_21173 =  x_893 & ~n_17844;
assign n_21174 =  n_17844 &  n_21137;
assign n_21175 = ~n_21173 & ~n_21174;
assign n_21176 =  x_893 & ~n_21175;
assign n_21177 = ~x_893 &  n_21175;
assign n_21178 = ~n_21176 & ~n_21177;
assign n_21179 =  x_892 & ~n_17851;
assign n_21180 =  n_17851 &  n_21137;
assign n_21181 = ~n_21179 & ~n_21180;
assign n_21182 =  x_892 & ~n_21181;
assign n_21183 = ~x_892 &  n_21181;
assign n_21184 = ~n_21182 & ~n_21183;
assign n_21185 =  x_891 & ~n_17789;
assign n_21186 =  x_1732 &  x_1744;
assign n_21187 =  n_21186 &  n_17789;
assign n_21188 = ~n_21185 & ~n_21187;
assign n_21189 =  x_891 & ~n_21188;
assign n_21190 = ~x_891 &  n_21188;
assign n_21191 = ~n_21189 & ~n_21190;
assign n_21192 =  x_890 & ~n_17807;
assign n_21193 =  n_21186 &  n_17807;
assign n_21194 = ~n_21192 & ~n_21193;
assign n_21195 =  x_890 & ~n_21194;
assign n_21196 = ~x_890 &  n_21194;
assign n_21197 = ~n_21195 & ~n_21196;
assign n_21198 =  x_889 & ~n_17815;
assign n_21199 =  n_21186 &  n_17815;
assign n_21200 = ~n_21198 & ~n_21199;
assign n_21201 =  x_889 & ~n_21200;
assign n_21202 = ~x_889 &  n_21200;
assign n_21203 = ~n_21201 & ~n_21202;
assign n_21204 =  x_888 & ~n_17823;
assign n_21205 =  n_17823 &  n_21186;
assign n_21206 = ~n_21204 & ~n_21205;
assign n_21207 =  x_888 & ~n_21206;
assign n_21208 = ~x_888 &  n_21206;
assign n_21209 = ~n_21207 & ~n_21208;
assign n_21210 =  x_887 & ~n_17830;
assign n_21211 =  n_21186 &  n_17830;
assign n_21212 = ~n_21210 & ~n_21211;
assign n_21213 =  x_887 & ~n_21212;
assign n_21214 = ~x_887 &  n_21212;
assign n_21215 = ~n_21213 & ~n_21214;
assign n_21216 =  x_886 & ~n_17837;
assign n_21217 =  n_21186 &  n_17837;
assign n_21218 = ~n_21216 & ~n_21217;
assign n_21219 =  x_886 & ~n_21218;
assign n_21220 = ~x_886 &  n_21218;
assign n_21221 = ~n_21219 & ~n_21220;
assign n_21222 =  x_885 & ~n_17844;
assign n_21223 =  n_21186 &  n_17844;
assign n_21224 = ~n_21222 & ~n_21223;
assign n_21225 =  x_885 & ~n_21224;
assign n_21226 = ~x_885 &  n_21224;
assign n_21227 = ~n_21225 & ~n_21226;
assign n_21228 =  x_884 & ~n_17851;
assign n_21229 =  n_17851 &  n_21186;
assign n_21230 = ~n_21228 & ~n_21229;
assign n_21231 =  x_884 & ~n_21230;
assign n_21232 = ~x_884 &  n_21230;
assign n_21233 = ~n_21231 & ~n_21232;
assign n_21234 =  x_883 & ~n_17822;
assign n_21235 = ~n_17823 & ~n_21234;
assign n_21236 =  x_883 & ~n_21235;
assign n_21237 = ~x_883 &  n_21235;
assign n_21238 = ~n_21236 & ~n_21237;
assign n_21239 = ~x_882 & ~n_17805;
assign n_21240 = ~n_17822 & ~n_21239;
assign n_21241 =  x_882 &  n_21240;
assign n_21242 = ~x_882 & ~n_21240;
assign n_21243 = ~n_21241 & ~n_21242;
assign n_21244 =  x_881 & ~x_1732;
assign n_21245 = ~n_17787 & ~n_21244;
assign n_21246 =  x_881 & ~n_21245;
assign n_21247 = ~x_881 &  n_21245;
assign n_21248 = ~n_21246 & ~n_21247;
assign n_21249 = ~x_1588 & ~x_1589;
assign n_21250 = ~x_1590 & ~x_1591;
assign n_21251 =  n_21249 &  n_21250;
assign n_21252 = ~x_1584 & ~x_1585;
assign n_21253 = ~x_1586 & ~x_1587;
assign n_21254 =  n_21252 &  n_21253;
assign n_21255 = ~x_1580 & ~x_1581;
assign n_21256 = ~x_1582 & ~x_1583;
assign n_21257 =  n_21255 &  n_21256;
assign n_21258 =  n_21254 &  n_21257;
assign n_21259 =  n_21251 &  n_21258;
assign n_21260 = ~x_1568 & ~x_1569;
assign n_21261 = ~x_1570 & ~x_1571;
assign n_21262 =  n_21260 &  n_21261;
assign n_21263 = ~x_1564 & ~x_1565;
assign n_21264 = ~x_1566 & ~x_1567;
assign n_21265 =  n_21263 &  n_21264;
assign n_21266 =  n_21262 &  n_21265;
assign n_21267 = ~x_1576 & ~x_1577;
assign n_21268 = ~x_1578 & ~x_1579;
assign n_21269 =  n_21267 &  n_21268;
assign n_21270 = ~x_1572 & ~x_1573;
assign n_21271 = ~x_1574 & ~x_1575;
assign n_21272 =  n_21270 &  n_21271;
assign n_21273 =  n_21269 &  n_21272;
assign n_21274 =  n_21266 &  n_21273;
assign n_21275 =  n_21259 &  n_21274;
assign n_21276 =  x_1563 & ~x_1592;
assign n_21277 =  n_21275 &  n_21276;
assign n_21278 =  n_17121 &  n_21277;
assign n_21279 = ~x_1594 &  x_1596;
assign n_21280 =  n_21278 &  n_21279;
assign n_21281 = ~n_3266 & ~n_21280;
assign n_21282 =  x_880 &  n_21281;
assign n_21283 =  x_434 & ~n_3266;
assign n_21284 =  n_21280 &  n_21283;
assign n_21285 = ~n_21282 & ~n_21284;
assign n_21286 =  x_880 & ~n_21285;
assign n_21287 = ~x_880 &  n_21285;
assign n_21288 = ~n_21286 & ~n_21287;
assign n_21289 = ~x_1563 &  n_21275;
assign n_21290 =  n_17129 &  n_21289;
assign n_21291 =  x_1593 &  n_21290;
assign n_21292 =  n_21279 &  n_21291;
assign n_21293 = ~n_3266 & ~n_21292;
assign n_21294 =  x_879 &  n_21293;
assign n_21295 =  n_21292 &  n_21283;
assign n_21296 = ~n_21294 & ~n_21295;
assign n_21297 =  x_879 & ~n_21296;
assign n_21298 = ~x_879 &  n_21296;
assign n_21299 = ~n_21297 & ~n_21298;
assign n_21300 = ~n_17129 &  n_21289;
assign n_21301 = ~n_17121 &  n_21300;
assign n_21302 =  n_21301 &  n_21279;
assign n_21303 = ~n_3266 & ~n_21302;
assign n_21304 =  x_878 &  n_21303;
assign n_21305 =  n_21302 &  n_21283;
assign n_21306 = ~n_21304 & ~n_21305;
assign n_21307 =  x_878 & ~n_21306;
assign n_21308 = ~x_878 &  n_21306;
assign n_21309 = ~n_21307 & ~n_21308;
assign n_21310 =  x_1595 &  n_21301;
assign n_21311 = ~n_3266 & ~n_21310;
assign n_21312 =  x_877 &  n_21311;
assign n_21313 =  n_21310 &  n_21283;
assign n_21314 = ~n_21312 & ~n_21313;
assign n_21315 =  x_877 & ~n_21314;
assign n_21316 = ~x_877 &  n_21314;
assign n_21317 = ~n_21315 & ~n_21316;
assign n_21318 =  x_1595 &  n_21291;
assign n_21319 = ~n_3266 & ~n_21318;
assign n_21320 =  x_876 &  n_21319;
assign n_21321 =  n_21318 &  n_21283;
assign n_21322 = ~n_21320 & ~n_21321;
assign n_21323 =  x_876 & ~n_21322;
assign n_21324 = ~x_876 &  n_21322;
assign n_21325 = ~n_21323 & ~n_21324;
assign n_21326 = ~x_1593 &  n_21290;
assign n_21327 =  n_21279 &  n_21326;
assign n_21328 = ~n_3266 & ~n_21327;
assign n_21329 =  x_875 &  n_21328;
assign n_21330 =  n_21327 &  n_21283;
assign n_21331 = ~n_21329 & ~n_21330;
assign n_21332 =  x_875 & ~n_21331;
assign n_21333 = ~x_875 &  n_21331;
assign n_21334 = ~n_21332 & ~n_21333;
assign n_21335 =  n_17121 &  n_21300;
assign n_21336 =  n_21279 &  n_21335;
assign n_21337 = ~n_3266 & ~n_21336;
assign n_21338 =  x_874 &  n_21337;
assign n_21339 =  n_21336 &  n_21283;
assign n_21340 = ~n_21338 & ~n_21339;
assign n_21341 =  x_874 & ~n_21340;
assign n_21342 = ~x_874 &  n_21340;
assign n_21343 = ~n_21341 & ~n_21342;
assign n_21344 =  x_1595 &  n_21326;
assign n_21345 = ~n_3266 & ~n_21344;
assign n_21346 =  x_873 &  n_21345;
assign n_21347 =  n_21344 &  n_21283;
assign n_21348 = ~n_21346 & ~n_21347;
assign n_21349 =  x_873 & ~n_21348;
assign n_21350 = ~x_873 &  n_21348;
assign n_21351 = ~n_21349 & ~n_21350;
assign n_21352 =  x_1595 &  n_21335;
assign n_21353 = ~n_3266 & ~n_21352;
assign n_21354 =  x_872 &  n_21353;
assign n_21355 =  n_21352 &  n_21283;
assign n_21356 = ~n_21354 & ~n_21355;
assign n_21357 =  x_872 & ~n_21356;
assign n_21358 = ~x_872 &  n_21356;
assign n_21359 = ~n_21357 & ~n_21358;
assign n_21360 = ~x_1593 &  n_21277;
assign n_21361 =  x_1595 &  n_21360;
assign n_21362 = ~n_3266 & ~n_21361;
assign n_21363 =  x_871 &  n_21362;
assign n_21364 =  n_21361 &  n_21283;
assign n_21365 = ~n_21363 & ~n_21364;
assign n_21366 =  x_871 & ~n_21365;
assign n_21367 = ~x_871 &  n_21365;
assign n_21368 = ~n_21366 & ~n_21367;
assign n_21369 =  x_1595 &  n_21278;
assign n_21370 = ~n_3266 & ~n_21369;
assign n_21371 =  x_870 &  n_21370;
assign n_21372 =  n_21369 &  n_21283;
assign n_21373 = ~n_21371 & ~n_21372;
assign n_21374 =  x_870 & ~n_21373;
assign n_21375 = ~x_870 &  n_21373;
assign n_21376 = ~n_21374 & ~n_21375;
assign n_21377 =  n_21279 &  n_21360;
assign n_21378 = ~n_3266 & ~n_21377;
assign n_21379 =  x_869 &  n_21378;
assign n_21380 =  n_21377 &  n_21283;
assign n_21381 = ~n_21379 & ~n_21380;
assign n_21382 =  x_869 & ~n_21381;
assign n_21383 = ~x_869 &  n_21381;
assign n_21384 = ~n_21382 & ~n_21383;
assign n_21385 =  x_868 &  n_21328;
assign n_21386 =  x_433 & ~n_3266;
assign n_21387 =  n_21327 &  n_21386;
assign n_21388 = ~n_21385 & ~n_21387;
assign n_21389 =  x_868 & ~n_21388;
assign n_21390 = ~x_868 &  n_21388;
assign n_21391 = ~n_21389 & ~n_21390;
assign n_21392 =  x_867 &  n_21281;
assign n_21393 =  n_21280 &  n_21386;
assign n_21394 = ~n_21392 & ~n_21393;
assign n_21395 =  x_867 & ~n_21394;
assign n_21396 = ~x_867 &  n_21394;
assign n_21397 = ~n_21395 & ~n_21396;
assign n_21398 =  x_866 &  n_21337;
assign n_21399 =  n_21336 &  n_21386;
assign n_21400 = ~n_21398 & ~n_21399;
assign n_21401 =  x_866 & ~n_21400;
assign n_21402 = ~x_866 &  n_21400;
assign n_21403 = ~n_21401 & ~n_21402;
assign n_21404 =  x_865 &  n_21353;
assign n_21405 =  n_21352 &  n_21386;
assign n_21406 = ~n_21404 & ~n_21405;
assign n_21407 =  x_865 & ~n_21406;
assign n_21408 = ~x_865 &  n_21406;
assign n_21409 = ~n_21407 & ~n_21408;
assign n_21410 =  x_864 &  n_21311;
assign n_21411 =  n_21310 &  n_21386;
assign n_21412 = ~n_21410 & ~n_21411;
assign n_21413 =  x_864 & ~n_21412;
assign n_21414 = ~x_864 &  n_21412;
assign n_21415 = ~n_21413 & ~n_21414;
assign n_21416 =  x_863 &  n_21362;
assign n_21417 =  n_21361 &  n_21386;
assign n_21418 = ~n_21416 & ~n_21417;
assign n_21419 =  x_863 & ~n_21418;
assign n_21420 = ~x_863 &  n_21418;
assign n_21421 = ~n_21419 & ~n_21420;
assign n_21422 =  x_862 &  n_21303;
assign n_21423 =  n_21302 &  n_21386;
assign n_21424 = ~n_21422 & ~n_21423;
assign n_21425 =  x_862 & ~n_21424;
assign n_21426 = ~x_862 &  n_21424;
assign n_21427 = ~n_21425 & ~n_21426;
assign n_21428 =  x_861 &  n_21345;
assign n_21429 =  n_21344 &  n_21386;
assign n_21430 = ~n_21428 & ~n_21429;
assign n_21431 =  x_861 & ~n_21430;
assign n_21432 = ~x_861 &  n_21430;
assign n_21433 = ~n_21431 & ~n_21432;
assign n_21434 =  x_860 &  n_21319;
assign n_21435 =  n_21318 &  n_21386;
assign n_21436 = ~n_21434 & ~n_21435;
assign n_21437 =  x_860 & ~n_21436;
assign n_21438 = ~x_860 &  n_21436;
assign n_21439 = ~n_21437 & ~n_21438;
assign n_21440 =  x_859 &  n_21378;
assign n_21441 =  n_21377 &  n_21386;
assign n_21442 = ~n_21440 & ~n_21441;
assign n_21443 =  x_859 & ~n_21442;
assign n_21444 = ~x_859 &  n_21442;
assign n_21445 = ~n_21443 & ~n_21444;
assign n_21446 =  x_858 &  n_21370;
assign n_21447 =  n_21369 &  n_21386;
assign n_21448 = ~n_21446 & ~n_21447;
assign n_21449 =  x_858 & ~n_21448;
assign n_21450 = ~x_858 &  n_21448;
assign n_21451 = ~n_21449 & ~n_21450;
assign n_21452 =  x_857 &  n_21293;
assign n_21453 =  n_21292 &  n_21386;
assign n_21454 = ~n_21452 & ~n_21453;
assign n_21455 =  x_857 & ~n_21454;
assign n_21456 = ~x_857 &  n_21454;
assign n_21457 = ~n_21455 & ~n_21456;
assign n_21458 =  x_856 &  n_21370;
assign n_21459 =  x_432 & ~n_3266;
assign n_21460 =  n_21369 &  n_21459;
assign n_21461 = ~n_21458 & ~n_21460;
assign n_21462 =  x_856 & ~n_21461;
assign n_21463 = ~x_856 &  n_21461;
assign n_21464 = ~n_21462 & ~n_21463;
assign n_21465 =  x_855 &  n_21378;
assign n_21466 =  n_21377 &  n_21459;
assign n_21467 = ~n_21465 & ~n_21466;
assign n_21468 =  x_855 & ~n_21467;
assign n_21469 = ~x_855 &  n_21467;
assign n_21470 = ~n_21468 & ~n_21469;
assign n_21471 =  x_854 &  n_21328;
assign n_21472 =  n_21327 &  n_21459;
assign n_21473 = ~n_21471 & ~n_21472;
assign n_21474 =  x_854 & ~n_21473;
assign n_21475 = ~x_854 &  n_21473;
assign n_21476 = ~n_21474 & ~n_21475;
assign n_21477 =  x_853 &  n_21311;
assign n_21478 =  n_21310 &  n_21459;
assign n_21479 = ~n_21477 & ~n_21478;
assign n_21480 =  x_853 & ~n_21479;
assign n_21481 = ~x_853 &  n_21479;
assign n_21482 = ~n_21480 & ~n_21481;
assign n_21483 =  x_852 &  n_21319;
assign n_21484 =  n_21318 &  n_21459;
assign n_21485 = ~n_21483 & ~n_21484;
assign n_21486 =  x_852 & ~n_21485;
assign n_21487 = ~x_852 &  n_21485;
assign n_21488 = ~n_21486 & ~n_21487;
assign n_21489 =  x_851 &  n_21337;
assign n_21490 =  n_21336 &  n_21459;
assign n_21491 = ~n_21489 & ~n_21490;
assign n_21492 =  x_851 & ~n_21491;
assign n_21493 = ~x_851 &  n_21491;
assign n_21494 = ~n_21492 & ~n_21493;
assign n_21495 =  x_850 &  n_21281;
assign n_21496 =  n_21280 &  n_21459;
assign n_21497 = ~n_21495 & ~n_21496;
assign n_21498 =  x_850 & ~n_21497;
assign n_21499 = ~x_850 &  n_21497;
assign n_21500 = ~n_21498 & ~n_21499;
assign n_21501 =  x_849 &  n_21362;
assign n_21502 =  n_21361 &  n_21459;
assign n_21503 = ~n_21501 & ~n_21502;
assign n_21504 =  x_849 & ~n_21503;
assign n_21505 = ~x_849 &  n_21503;
assign n_21506 = ~n_21504 & ~n_21505;
assign n_21507 =  x_848 &  n_21293;
assign n_21508 =  n_21292 &  n_21459;
assign n_21509 = ~n_21507 & ~n_21508;
assign n_21510 =  x_848 & ~n_21509;
assign n_21511 = ~x_848 &  n_21509;
assign n_21512 = ~n_21510 & ~n_21511;
assign n_21513 =  x_847 &  n_21303;
assign n_21514 =  n_21302 &  n_21459;
assign n_21515 = ~n_21513 & ~n_21514;
assign n_21516 =  x_847 & ~n_21515;
assign n_21517 = ~x_847 &  n_21515;
assign n_21518 = ~n_21516 & ~n_21517;
assign n_21519 =  x_846 &  n_21345;
assign n_21520 =  n_21344 &  n_21459;
assign n_21521 = ~n_21519 & ~n_21520;
assign n_21522 =  x_846 & ~n_21521;
assign n_21523 = ~x_846 &  n_21521;
assign n_21524 = ~n_21522 & ~n_21523;
assign n_21525 =  x_845 &  n_21353;
assign n_21526 =  n_21352 &  n_21459;
assign n_21527 = ~n_21525 & ~n_21526;
assign n_21528 =  x_845 & ~n_21527;
assign n_21529 = ~x_845 &  n_21527;
assign n_21530 = ~n_21528 & ~n_21529;
assign n_21531 =  x_844 &  n_21378;
assign n_21532 =  x_431 & ~n_3266;
assign n_21533 =  n_21377 &  n_21532;
assign n_21534 = ~n_21531 & ~n_21533;
assign n_21535 =  x_844 & ~n_21534;
assign n_21536 = ~x_844 &  n_21534;
assign n_21537 = ~n_21535 & ~n_21536;
assign n_21538 =  x_843 &  n_21303;
assign n_21539 =  n_21302 &  n_21532;
assign n_21540 = ~n_21538 & ~n_21539;
assign n_21541 =  x_843 & ~n_21540;
assign n_21542 = ~x_843 &  n_21540;
assign n_21543 = ~n_21541 & ~n_21542;
assign n_21544 =  x_842 &  n_21319;
assign n_21545 =  n_21318 &  n_21532;
assign n_21546 = ~n_21544 & ~n_21545;
assign n_21547 =  x_842 & ~n_21546;
assign n_21548 = ~x_842 &  n_21546;
assign n_21549 = ~n_21547 & ~n_21548;
assign n_21550 =  x_841 &  n_21293;
assign n_21551 =  n_21292 &  n_21532;
assign n_21552 = ~n_21550 & ~n_21551;
assign n_21553 =  x_841 & ~n_21552;
assign n_21554 = ~x_841 &  n_21552;
assign n_21555 = ~n_21553 & ~n_21554;
assign n_21556 =  x_840 &  n_21337;
assign n_21557 =  n_21336 &  n_21532;
assign n_21558 = ~n_21556 & ~n_21557;
assign n_21559 =  x_840 & ~n_21558;
assign n_21560 = ~x_840 &  n_21558;
assign n_21561 = ~n_21559 & ~n_21560;
assign n_21562 =  x_839 &  n_21370;
assign n_21563 =  n_21369 &  n_21532;
assign n_21564 = ~n_21562 & ~n_21563;
assign n_21565 =  x_839 & ~n_21564;
assign n_21566 = ~x_839 &  n_21564;
assign n_21567 = ~n_21565 & ~n_21566;
assign n_21568 =  x_838 &  n_21281;
assign n_21569 =  n_21280 &  n_21532;
assign n_21570 = ~n_21568 & ~n_21569;
assign n_21571 =  x_838 & ~n_21570;
assign n_21572 = ~x_838 &  n_21570;
assign n_21573 = ~n_21571 & ~n_21572;
assign n_21574 =  x_837 &  n_21353;
assign n_21575 =  n_21352 &  n_21532;
assign n_21576 = ~n_21574 & ~n_21575;
assign n_21577 =  x_837 & ~n_21576;
assign n_21578 = ~x_837 &  n_21576;
assign n_21579 = ~n_21577 & ~n_21578;
assign n_21580 =  x_836 &  n_21311;
assign n_21581 =  n_21310 &  n_21532;
assign n_21582 = ~n_21580 & ~n_21581;
assign n_21583 =  x_836 & ~n_21582;
assign n_21584 = ~x_836 &  n_21582;
assign n_21585 = ~n_21583 & ~n_21584;
assign n_21586 =  x_835 &  n_21328;
assign n_21587 =  n_21327 &  n_21532;
assign n_21588 = ~n_21586 & ~n_21587;
assign n_21589 =  x_835 & ~n_21588;
assign n_21590 = ~x_835 &  n_21588;
assign n_21591 = ~n_21589 & ~n_21590;
assign n_21592 =  x_834 &  n_21345;
assign n_21593 =  n_21344 &  n_21532;
assign n_21594 = ~n_21592 & ~n_21593;
assign n_21595 =  x_834 & ~n_21594;
assign n_21596 = ~x_834 &  n_21594;
assign n_21597 = ~n_21595 & ~n_21596;
assign n_21598 =  x_833 &  n_21362;
assign n_21599 =  n_21361 &  n_21532;
assign n_21600 = ~n_21598 & ~n_21599;
assign n_21601 =  x_833 & ~n_21600;
assign n_21602 = ~x_833 &  n_21600;
assign n_21603 = ~n_21601 & ~n_21602;
assign n_21604 =  x_832 &  n_21319;
assign n_21605 =  x_430 & ~n_3266;
assign n_21606 =  n_21318 &  n_21605;
assign n_21607 = ~n_21604 & ~n_21606;
assign n_21608 =  x_832 & ~n_21607;
assign n_21609 = ~x_832 &  n_21607;
assign n_21610 = ~n_21608 & ~n_21609;
assign n_21611 =  x_831 &  n_21328;
assign n_21612 =  n_21327 &  n_21605;
assign n_21613 = ~n_21611 & ~n_21612;
assign n_21614 =  x_831 & ~n_21613;
assign n_21615 = ~x_831 &  n_21613;
assign n_21616 = ~n_21614 & ~n_21615;
assign n_21617 =  x_830 &  n_21362;
assign n_21618 =  n_21361 &  n_21605;
assign n_21619 = ~n_21617 & ~n_21618;
assign n_21620 =  x_830 & ~n_21619;
assign n_21621 = ~x_830 &  n_21619;
assign n_21622 = ~n_21620 & ~n_21621;
assign n_21623 =  x_829 &  n_21311;
assign n_21624 =  n_21310 &  n_21605;
assign n_21625 = ~n_21623 & ~n_21624;
assign n_21626 =  x_829 & ~n_21625;
assign n_21627 = ~x_829 &  n_21625;
assign n_21628 = ~n_21626 & ~n_21627;
assign n_21629 =  x_828 &  n_21353;
assign n_21630 =  n_21352 &  n_21605;
assign n_21631 = ~n_21629 & ~n_21630;
assign n_21632 =  x_828 & ~n_21631;
assign n_21633 = ~x_828 &  n_21631;
assign n_21634 = ~n_21632 & ~n_21633;
assign n_21635 =  x_827 &  n_21337;
assign n_21636 =  n_21336 &  n_21605;
assign n_21637 = ~n_21635 & ~n_21636;
assign n_21638 =  x_827 & ~n_21637;
assign n_21639 = ~x_827 &  n_21637;
assign n_21640 = ~n_21638 & ~n_21639;
assign n_21641 =  x_826 &  n_21378;
assign n_21642 =  n_21377 &  n_21605;
assign n_21643 = ~n_21641 & ~n_21642;
assign n_21644 =  x_826 & ~n_21643;
assign n_21645 = ~x_826 &  n_21643;
assign n_21646 = ~n_21644 & ~n_21645;
assign n_21647 =  x_825 &  n_21293;
assign n_21648 =  n_21292 &  n_21605;
assign n_21649 = ~n_21647 & ~n_21648;
assign n_21650 =  x_825 & ~n_21649;
assign n_21651 = ~x_825 &  n_21649;
assign n_21652 = ~n_21650 & ~n_21651;
assign n_21653 =  x_824 &  n_21345;
assign n_21654 =  n_21344 &  n_21605;
assign n_21655 = ~n_21653 & ~n_21654;
assign n_21656 =  x_824 & ~n_21655;
assign n_21657 = ~x_824 &  n_21655;
assign n_21658 = ~n_21656 & ~n_21657;
assign n_21659 =  x_823 &  n_21281;
assign n_21660 =  n_21280 &  n_21605;
assign n_21661 = ~n_21659 & ~n_21660;
assign n_21662 =  x_823 & ~n_21661;
assign n_21663 = ~x_823 &  n_21661;
assign n_21664 = ~n_21662 & ~n_21663;
assign n_21665 =  x_822 &  n_21370;
assign n_21666 =  n_21369 &  n_21605;
assign n_21667 = ~n_21665 & ~n_21666;
assign n_21668 =  x_822 & ~n_21667;
assign n_21669 = ~x_822 &  n_21667;
assign n_21670 = ~n_21668 & ~n_21669;
assign n_21671 =  x_821 &  n_21303;
assign n_21672 =  n_21302 &  n_21605;
assign n_21673 = ~n_21671 & ~n_21672;
assign n_21674 =  x_821 & ~n_21673;
assign n_21675 = ~x_821 &  n_21673;
assign n_21676 = ~n_21674 & ~n_21675;
assign n_21677 =  x_820 &  n_21293;
assign n_21678 =  x_429 & ~n_3266;
assign n_21679 =  n_21292 &  n_21678;
assign n_21680 = ~n_21677 & ~n_21679;
assign n_21681 =  x_820 & ~n_21680;
assign n_21682 = ~x_820 &  n_21680;
assign n_21683 = ~n_21681 & ~n_21682;
assign n_21684 =  x_819 &  n_21328;
assign n_21685 =  n_21327 &  n_21678;
assign n_21686 = ~n_21684 & ~n_21685;
assign n_21687 =  x_819 & ~n_21686;
assign n_21688 = ~x_819 &  n_21686;
assign n_21689 = ~n_21687 & ~n_21688;
assign n_21690 =  x_818 &  n_21370;
assign n_21691 =  n_21369 &  n_21678;
assign n_21692 = ~n_21690 & ~n_21691;
assign n_21693 =  x_818 & ~n_21692;
assign n_21694 = ~x_818 &  n_21692;
assign n_21695 = ~n_21693 & ~n_21694;
assign n_21696 =  x_817 &  n_21281;
assign n_21697 =  n_21280 &  n_21678;
assign n_21698 = ~n_21696 & ~n_21697;
assign n_21699 =  x_817 & ~n_21698;
assign n_21700 = ~x_817 &  n_21698;
assign n_21701 = ~n_21699 & ~n_21700;
assign n_21702 =  x_816 &  n_21378;
assign n_21703 =  n_21377 &  n_21678;
assign n_21704 = ~n_21702 & ~n_21703;
assign n_21705 =  x_816 & ~n_21704;
assign n_21706 = ~x_816 &  n_21704;
assign n_21707 = ~n_21705 & ~n_21706;
assign n_21708 =  x_815 &  n_21337;
assign n_21709 =  n_21336 &  n_21678;
assign n_21710 = ~n_21708 & ~n_21709;
assign n_21711 =  x_815 & ~n_21710;
assign n_21712 = ~x_815 &  n_21710;
assign n_21713 = ~n_21711 & ~n_21712;
assign n_21714 =  x_814 &  n_21345;
assign n_21715 =  n_21344 &  n_21678;
assign n_21716 = ~n_21714 & ~n_21715;
assign n_21717 =  x_814 & ~n_21716;
assign n_21718 = ~x_814 &  n_21716;
assign n_21719 = ~n_21717 & ~n_21718;
assign n_21720 =  x_813 &  n_21353;
assign n_21721 =  n_21352 &  n_21678;
assign n_21722 = ~n_21720 & ~n_21721;
assign n_21723 =  x_813 & ~n_21722;
assign n_21724 = ~x_813 &  n_21722;
assign n_21725 = ~n_21723 & ~n_21724;
assign n_21726 =  x_812 &  n_21303;
assign n_21727 =  n_21302 &  n_21678;
assign n_21728 = ~n_21726 & ~n_21727;
assign n_21729 =  x_812 & ~n_21728;
assign n_21730 = ~x_812 &  n_21728;
assign n_21731 = ~n_21729 & ~n_21730;
assign n_21732 =  x_811 &  n_21319;
assign n_21733 =  n_21318 &  n_21678;
assign n_21734 = ~n_21732 & ~n_21733;
assign n_21735 =  x_811 & ~n_21734;
assign n_21736 = ~x_811 &  n_21734;
assign n_21737 = ~n_21735 & ~n_21736;
assign n_21738 =  x_810 &  n_21311;
assign n_21739 =  n_21310 &  n_21678;
assign n_21740 = ~n_21738 & ~n_21739;
assign n_21741 =  x_810 & ~n_21740;
assign n_21742 = ~x_810 &  n_21740;
assign n_21743 = ~n_21741 & ~n_21742;
assign n_21744 =  x_809 &  n_21362;
assign n_21745 =  n_21361 &  n_21678;
assign n_21746 = ~n_21744 & ~n_21745;
assign n_21747 =  x_809 & ~n_21746;
assign n_21748 = ~x_809 &  n_21746;
assign n_21749 = ~n_21747 & ~n_21748;
assign n_21750 =  x_808 &  n_21328;
assign n_21751 =  x_428 & ~n_3266;
assign n_21752 =  n_21327 &  n_21751;
assign n_21753 = ~n_21750 & ~n_21752;
assign n_21754 =  x_808 & ~n_21753;
assign n_21755 = ~x_808 &  n_21753;
assign n_21756 = ~n_21754 & ~n_21755;
assign n_21757 =  x_807 &  n_21303;
assign n_21758 =  n_21302 &  n_21751;
assign n_21759 = ~n_21757 & ~n_21758;
assign n_21760 =  x_807 & ~n_21759;
assign n_21761 = ~x_807 &  n_21759;
assign n_21762 = ~n_21760 & ~n_21761;
assign n_21763 =  x_806 &  n_21370;
assign n_21764 =  n_21369 &  n_21751;
assign n_21765 = ~n_21763 & ~n_21764;
assign n_21766 =  x_806 & ~n_21765;
assign n_21767 = ~x_806 &  n_21765;
assign n_21768 = ~n_21766 & ~n_21767;
assign n_21769 =  x_805 &  n_21362;
assign n_21770 =  n_21361 &  n_21751;
assign n_21771 = ~n_21769 & ~n_21770;
assign n_21772 =  x_805 & ~n_21771;
assign n_21773 = ~x_805 &  n_21771;
assign n_21774 = ~n_21772 & ~n_21773;
assign n_21775 =  x_804 &  n_21378;
assign n_21776 =  n_21377 &  n_21751;
assign n_21777 = ~n_21775 & ~n_21776;
assign n_21778 =  x_804 & ~n_21777;
assign n_21779 = ~x_804 &  n_21777;
assign n_21780 = ~n_21778 & ~n_21779;
assign n_21781 =  x_803 &  n_21311;
assign n_21782 =  n_21310 &  n_21751;
assign n_21783 = ~n_21781 & ~n_21782;
assign n_21784 =  x_803 & ~n_21783;
assign n_21785 = ~x_803 &  n_21783;
assign n_21786 = ~n_21784 & ~n_21785;
assign n_21787 =  x_802 &  n_21345;
assign n_21788 =  n_21344 &  n_21751;
assign n_21789 = ~n_21787 & ~n_21788;
assign n_21790 =  x_802 & ~n_21789;
assign n_21791 = ~x_802 &  n_21789;
assign n_21792 = ~n_21790 & ~n_21791;
assign n_21793 =  x_801 &  n_21293;
assign n_21794 =  n_21292 &  n_21751;
assign n_21795 = ~n_21793 & ~n_21794;
assign n_21796 =  x_801 & ~n_21795;
assign n_21797 = ~x_801 &  n_21795;
assign n_21798 = ~n_21796 & ~n_21797;
assign n_21799 =  x_800 &  n_21337;
assign n_21800 =  n_21336 &  n_21751;
assign n_21801 = ~n_21799 & ~n_21800;
assign n_21802 =  x_800 & ~n_21801;
assign n_21803 = ~x_800 &  n_21801;
assign n_21804 = ~n_21802 & ~n_21803;
assign n_21805 =  x_799 &  n_21353;
assign n_21806 =  n_21352 &  n_21751;
assign n_21807 = ~n_21805 & ~n_21806;
assign n_21808 =  x_799 & ~n_21807;
assign n_21809 = ~x_799 &  n_21807;
assign n_21810 = ~n_21808 & ~n_21809;
assign n_21811 =  x_798 &  n_21319;
assign n_21812 =  n_21318 &  n_21751;
assign n_21813 = ~n_21811 & ~n_21812;
assign n_21814 =  x_798 & ~n_21813;
assign n_21815 = ~x_798 &  n_21813;
assign n_21816 = ~n_21814 & ~n_21815;
assign n_21817 =  x_797 &  n_21281;
assign n_21818 =  n_21280 &  n_21751;
assign n_21819 = ~n_21817 & ~n_21818;
assign n_21820 =  x_797 & ~n_21819;
assign n_21821 = ~x_797 &  n_21819;
assign n_21822 = ~n_21820 & ~n_21821;
assign n_21823 =  x_796 &  n_21362;
assign n_21824 =  x_427 & ~n_3266;
assign n_21825 =  n_21361 &  n_21824;
assign n_21826 = ~n_21823 & ~n_21825;
assign n_21827 =  x_796 & ~n_21826;
assign n_21828 = ~x_796 &  n_21826;
assign n_21829 = ~n_21827 & ~n_21828;
assign n_21830 =  x_795 &  n_21281;
assign n_21831 =  n_21280 &  n_21824;
assign n_21832 = ~n_21830 & ~n_21831;
assign n_21833 =  x_795 & ~n_21832;
assign n_21834 = ~x_795 &  n_21832;
assign n_21835 = ~n_21833 & ~n_21834;
assign n_21836 =  x_794 &  n_21328;
assign n_21837 =  n_21327 &  n_21824;
assign n_21838 = ~n_21836 & ~n_21837;
assign n_21839 =  x_794 & ~n_21838;
assign n_21840 = ~x_794 &  n_21838;
assign n_21841 = ~n_21839 & ~n_21840;
assign n_21842 =  x_793 &  n_21353;
assign n_21843 =  n_21352 &  n_21824;
assign n_21844 = ~n_21842 & ~n_21843;
assign n_21845 =  x_793 & ~n_21844;
assign n_21846 = ~x_793 &  n_21844;
assign n_21847 = ~n_21845 & ~n_21846;
assign n_21848 =  x_792 &  n_21293;
assign n_21849 =  n_21292 &  n_21824;
assign n_21850 = ~n_21848 & ~n_21849;
assign n_21851 =  x_792 & ~n_21850;
assign n_21852 = ~x_792 &  n_21850;
assign n_21853 = ~n_21851 & ~n_21852;
assign n_21854 =  x_791 &  n_21370;
assign n_21855 =  n_21369 &  n_21824;
assign n_21856 = ~n_21854 & ~n_21855;
assign n_21857 =  x_791 & ~n_21856;
assign n_21858 = ~x_791 &  n_21856;
assign n_21859 = ~n_21857 & ~n_21858;
assign n_21860 =  x_790 &  n_21303;
assign n_21861 =  n_21302 &  n_21824;
assign n_21862 = ~n_21860 & ~n_21861;
assign n_21863 =  x_790 & ~n_21862;
assign n_21864 = ~x_790 &  n_21862;
assign n_21865 = ~n_21863 & ~n_21864;
assign n_21866 =  x_789 &  n_21345;
assign n_21867 =  n_21344 &  n_21824;
assign n_21868 = ~n_21866 & ~n_21867;
assign n_21869 =  x_789 & ~n_21868;
assign n_21870 = ~x_789 &  n_21868;
assign n_21871 = ~n_21869 & ~n_21870;
assign n_21872 =  x_788 &  n_21337;
assign n_21873 =  n_21336 &  n_21824;
assign n_21874 = ~n_21872 & ~n_21873;
assign n_21875 =  x_788 & ~n_21874;
assign n_21876 = ~x_788 &  n_21874;
assign n_21877 = ~n_21875 & ~n_21876;
assign n_21878 =  x_787 &  n_21311;
assign n_21879 =  n_21310 &  n_21824;
assign n_21880 = ~n_21878 & ~n_21879;
assign n_21881 =  x_787 & ~n_21880;
assign n_21882 = ~x_787 &  n_21880;
assign n_21883 = ~n_21881 & ~n_21882;
assign n_21884 =  x_786 &  n_21378;
assign n_21885 =  n_21377 &  n_21824;
assign n_21886 = ~n_21884 & ~n_21885;
assign n_21887 =  x_786 & ~n_21886;
assign n_21888 = ~x_786 &  n_21886;
assign n_21889 = ~n_21887 & ~n_21888;
assign n_21890 =  x_785 &  n_21319;
assign n_21891 =  n_21318 &  n_21824;
assign n_21892 = ~n_21890 & ~n_21891;
assign n_21893 =  x_785 & ~n_21892;
assign n_21894 = ~x_785 &  n_21892;
assign n_21895 = ~n_21893 & ~n_21894;
assign n_21896 =  x_784 &  n_21281;
assign n_21897 =  x_426 & ~n_3266;
assign n_21898 =  n_21280 &  n_21897;
assign n_21899 = ~n_21896 & ~n_21898;
assign n_21900 =  x_784 & ~n_21899;
assign n_21901 = ~x_784 &  n_21899;
assign n_21902 = ~n_21900 & ~n_21901;
assign n_21903 =  x_783 &  n_21293;
assign n_21904 =  n_21292 &  n_21897;
assign n_21905 = ~n_21903 & ~n_21904;
assign n_21906 =  x_783 & ~n_21905;
assign n_21907 = ~x_783 &  n_21905;
assign n_21908 = ~n_21906 & ~n_21907;
assign n_21909 =  x_782 &  n_21319;
assign n_21910 =  n_21318 &  n_21897;
assign n_21911 = ~n_21909 & ~n_21910;
assign n_21912 =  x_782 & ~n_21911;
assign n_21913 = ~x_782 &  n_21911;
assign n_21914 = ~n_21912 & ~n_21913;
assign n_21915 =  x_781 &  n_21303;
assign n_21916 =  n_21302 &  n_21897;
assign n_21917 = ~n_21915 & ~n_21916;
assign n_21918 =  x_781 & ~n_21917;
assign n_21919 = ~x_781 &  n_21917;
assign n_21920 = ~n_21918 & ~n_21919;
assign n_21921 =  x_780 &  n_21311;
assign n_21922 =  n_21310 &  n_21897;
assign n_21923 = ~n_21921 & ~n_21922;
assign n_21924 =  x_780 & ~n_21923;
assign n_21925 = ~x_780 &  n_21923;
assign n_21926 = ~n_21924 & ~n_21925;
assign n_21927 =  x_779 &  n_21328;
assign n_21928 =  n_21327 &  n_21897;
assign n_21929 = ~n_21927 & ~n_21928;
assign n_21930 =  x_779 & ~n_21929;
assign n_21931 = ~x_779 &  n_21929;
assign n_21932 = ~n_21930 & ~n_21931;
assign n_21933 =  x_778 &  n_21337;
assign n_21934 =  n_21336 &  n_21897;
assign n_21935 = ~n_21933 & ~n_21934;
assign n_21936 =  x_778 & ~n_21935;
assign n_21937 = ~x_778 &  n_21935;
assign n_21938 = ~n_21936 & ~n_21937;
assign n_21939 =  x_777 &  n_21345;
assign n_21940 =  n_21344 &  n_21897;
assign n_21941 = ~n_21939 & ~n_21940;
assign n_21942 =  x_777 & ~n_21941;
assign n_21943 = ~x_777 &  n_21941;
assign n_21944 = ~n_21942 & ~n_21943;
assign n_21945 =  x_776 &  n_21353;
assign n_21946 =  n_21352 &  n_21897;
assign n_21947 = ~n_21945 & ~n_21946;
assign n_21948 =  x_776 & ~n_21947;
assign n_21949 = ~x_776 &  n_21947;
assign n_21950 = ~n_21948 & ~n_21949;
assign n_21951 =  x_775 &  n_21362;
assign n_21952 =  n_21361 &  n_21897;
assign n_21953 = ~n_21951 & ~n_21952;
assign n_21954 =  x_775 & ~n_21953;
assign n_21955 = ~x_775 &  n_21953;
assign n_21956 = ~n_21954 & ~n_21955;
assign n_21957 =  x_774 &  n_21370;
assign n_21958 =  n_21369 &  n_21897;
assign n_21959 = ~n_21957 & ~n_21958;
assign n_21960 =  x_774 & ~n_21959;
assign n_21961 = ~x_774 &  n_21959;
assign n_21962 = ~n_21960 & ~n_21961;
assign n_21963 =  x_773 &  n_21378;
assign n_21964 =  n_21377 &  n_21897;
assign n_21965 = ~n_21963 & ~n_21964;
assign n_21966 =  x_773 & ~n_21965;
assign n_21967 = ~x_773 &  n_21965;
assign n_21968 = ~n_21966 & ~n_21967;
assign n_21969 =  x_772 &  n_21337;
assign n_21970 =  x_425 & ~n_3266;
assign n_21971 =  n_21336 &  n_21970;
assign n_21972 = ~n_21969 & ~n_21971;
assign n_21973 =  x_772 & ~n_21972;
assign n_21974 = ~x_772 &  n_21972;
assign n_21975 = ~n_21973 & ~n_21974;
assign n_21976 =  x_771 &  n_21378;
assign n_21977 =  n_21377 &  n_21970;
assign n_21978 = ~n_21976 & ~n_21977;
assign n_21979 =  x_771 & ~n_21978;
assign n_21980 = ~x_771 &  n_21978;
assign n_21981 = ~n_21979 & ~n_21980;
assign n_21982 =  x_770 &  n_21353;
assign n_21983 =  n_21352 &  n_21970;
assign n_21984 = ~n_21982 & ~n_21983;
assign n_21985 =  x_770 & ~n_21984;
assign n_21986 = ~x_770 &  n_21984;
assign n_21987 = ~n_21985 & ~n_21986;
assign n_21988 =  x_769 &  n_21303;
assign n_21989 =  n_21302 &  n_21970;
assign n_21990 = ~n_21988 & ~n_21989;
assign n_21991 =  x_769 & ~n_21990;
assign n_21992 = ~x_769 &  n_21990;
assign n_21993 = ~n_21991 & ~n_21992;
assign n_21994 =  x_768 &  n_21328;
assign n_21995 =  n_21327 &  n_21970;
assign n_21996 = ~n_21994 & ~n_21995;
assign n_21997 =  x_768 & ~n_21996;
assign n_21998 = ~x_768 &  n_21996;
assign n_21999 = ~n_21997 & ~n_21998;
assign n_22000 =  x_767 &  n_21281;
assign n_22001 =  n_21280 &  n_21970;
assign n_22002 = ~n_22000 & ~n_22001;
assign n_22003 =  x_767 & ~n_22002;
assign n_22004 = ~x_767 &  n_22002;
assign n_22005 = ~n_22003 & ~n_22004;
assign n_22006 =  x_766 &  n_21293;
assign n_22007 =  n_21292 &  n_21970;
assign n_22008 = ~n_22006 & ~n_22007;
assign n_22009 =  x_766 & ~n_22008;
assign n_22010 = ~x_766 &  n_22008;
assign n_22011 = ~n_22009 & ~n_22010;
assign n_22012 =  x_765 &  n_21345;
assign n_22013 =  n_21344 &  n_21970;
assign n_22014 = ~n_22012 & ~n_22013;
assign n_22015 =  x_765 & ~n_22014;
assign n_22016 = ~x_765 &  n_22014;
assign n_22017 = ~n_22015 & ~n_22016;
assign n_22018 =  x_764 &  n_21319;
assign n_22019 =  n_21318 &  n_21970;
assign n_22020 = ~n_22018 & ~n_22019;
assign n_22021 =  x_764 & ~n_22020;
assign n_22022 = ~x_764 &  n_22020;
assign n_22023 = ~n_22021 & ~n_22022;
assign n_22024 =  x_763 &  n_21362;
assign n_22025 =  n_21361 &  n_21970;
assign n_22026 = ~n_22024 & ~n_22025;
assign n_22027 =  x_763 & ~n_22026;
assign n_22028 = ~x_763 &  n_22026;
assign n_22029 = ~n_22027 & ~n_22028;
assign n_22030 =  x_762 &  n_21370;
assign n_22031 =  n_21369 &  n_21970;
assign n_22032 = ~n_22030 & ~n_22031;
assign n_22033 =  x_762 & ~n_22032;
assign n_22034 = ~x_762 &  n_22032;
assign n_22035 = ~n_22033 & ~n_22034;
assign n_22036 =  x_761 &  n_21311;
assign n_22037 =  n_21310 &  n_21970;
assign n_22038 = ~n_22036 & ~n_22037;
assign n_22039 =  x_761 & ~n_22038;
assign n_22040 = ~x_761 &  n_22038;
assign n_22041 = ~n_22039 & ~n_22040;
assign n_22042 =  x_760 &  n_21328;
assign n_22043 =  x_424 & ~n_3266;
assign n_22044 =  n_21327 &  n_22043;
assign n_22045 = ~n_22042 & ~n_22044;
assign n_22046 =  x_760 & ~n_22045;
assign n_22047 = ~x_760 &  n_22045;
assign n_22048 = ~n_22046 & ~n_22047;
assign n_22049 =  x_759 &  n_21293;
assign n_22050 =  n_21292 &  n_22043;
assign n_22051 = ~n_22049 & ~n_22050;
assign n_22052 =  x_759 & ~n_22051;
assign n_22053 = ~x_759 &  n_22051;
assign n_22054 = ~n_22052 & ~n_22053;
assign n_22055 =  x_758 &  n_21362;
assign n_22056 =  n_21361 &  n_22043;
assign n_22057 = ~n_22055 & ~n_22056;
assign n_22058 =  x_758 & ~n_22057;
assign n_22059 = ~x_758 &  n_22057;
assign n_22060 = ~n_22058 & ~n_22059;
assign n_22061 =  x_757 &  n_21353;
assign n_22062 =  n_21352 &  n_22043;
assign n_22063 = ~n_22061 & ~n_22062;
assign n_22064 =  x_757 & ~n_22063;
assign n_22065 = ~x_757 &  n_22063;
assign n_22066 = ~n_22064 & ~n_22065;
assign n_22067 =  x_756 &  n_21303;
assign n_22068 =  n_21302 &  n_22043;
assign n_22069 = ~n_22067 & ~n_22068;
assign n_22070 =  x_756 & ~n_22069;
assign n_22071 = ~x_756 &  n_22069;
assign n_22072 = ~n_22070 & ~n_22071;
assign n_22073 =  x_755 &  n_21281;
assign n_22074 =  n_21280 &  n_22043;
assign n_22075 = ~n_22073 & ~n_22074;
assign n_22076 =  x_755 & ~n_22075;
assign n_22077 = ~x_755 &  n_22075;
assign n_22078 = ~n_22076 & ~n_22077;
assign n_22079 =  x_754 &  n_21378;
assign n_22080 =  n_21377 &  n_22043;
assign n_22081 = ~n_22079 & ~n_22080;
assign n_22082 =  x_754 & ~n_22081;
assign n_22083 = ~x_754 &  n_22081;
assign n_22084 = ~n_22082 & ~n_22083;
assign n_22085 =  x_753 &  n_21319;
assign n_22086 =  n_21318 &  n_22043;
assign n_22087 = ~n_22085 & ~n_22086;
assign n_22088 =  x_753 & ~n_22087;
assign n_22089 = ~x_753 &  n_22087;
assign n_22090 = ~n_22088 & ~n_22089;
assign n_22091 =  x_752 &  n_21311;
assign n_22092 =  n_21310 &  n_22043;
assign n_22093 = ~n_22091 & ~n_22092;
assign n_22094 =  x_752 & ~n_22093;
assign n_22095 = ~x_752 &  n_22093;
assign n_22096 = ~n_22094 & ~n_22095;
assign n_22097 =  x_751 &  n_21345;
assign n_22098 =  n_21344 &  n_22043;
assign n_22099 = ~n_22097 & ~n_22098;
assign n_22100 =  x_751 & ~n_22099;
assign n_22101 = ~x_751 &  n_22099;
assign n_22102 = ~n_22100 & ~n_22101;
assign n_22103 =  x_750 &  n_21337;
assign n_22104 =  n_21336 &  n_22043;
assign n_22105 = ~n_22103 & ~n_22104;
assign n_22106 =  x_750 & ~n_22105;
assign n_22107 = ~x_750 &  n_22105;
assign n_22108 = ~n_22106 & ~n_22107;
assign n_22109 =  x_749 &  n_21370;
assign n_22110 =  n_21369 &  n_22043;
assign n_22111 = ~n_22109 & ~n_22110;
assign n_22112 =  x_749 & ~n_22111;
assign n_22113 = ~x_749 &  n_22111;
assign n_22114 = ~n_22112 & ~n_22113;
assign n_22115 =  x_748 &  n_21281;
assign n_22116 =  x_423 & ~n_3266;
assign n_22117 =  n_21280 &  n_22116;
assign n_22118 = ~n_22115 & ~n_22117;
assign n_22119 =  x_748 & ~n_22118;
assign n_22120 = ~x_748 &  n_22118;
assign n_22121 = ~n_22119 & ~n_22120;
assign n_22122 =  x_747 &  n_21303;
assign n_22123 =  n_21302 &  n_22116;
assign n_22124 = ~n_22122 & ~n_22123;
assign n_22125 =  x_747 & ~n_22124;
assign n_22126 = ~x_747 &  n_22124;
assign n_22127 = ~n_22125 & ~n_22126;
assign n_22128 =  x_746 &  n_21328;
assign n_22129 =  n_21327 &  n_22116;
assign n_22130 = ~n_22128 & ~n_22129;
assign n_22131 =  x_746 & ~n_22130;
assign n_22132 = ~x_746 &  n_22130;
assign n_22133 = ~n_22131 & ~n_22132;
assign n_22134 =  x_745 &  n_21337;
assign n_22135 =  n_21336 &  n_22116;
assign n_22136 = ~n_22134 & ~n_22135;
assign n_22137 =  x_745 & ~n_22136;
assign n_22138 = ~x_745 &  n_22136;
assign n_22139 = ~n_22137 & ~n_22138;
assign n_22140 =  x_744 &  n_21370;
assign n_22141 =  n_21369 &  n_22116;
assign n_22142 = ~n_22140 & ~n_22141;
assign n_22143 =  x_744 & ~n_22142;
assign n_22144 = ~x_744 &  n_22142;
assign n_22145 = ~n_22143 & ~n_22144;
assign n_22146 =  x_743 &  n_21319;
assign n_22147 =  n_21318 &  n_22116;
assign n_22148 = ~n_22146 & ~n_22147;
assign n_22149 =  x_743 & ~n_22148;
assign n_22150 = ~x_743 &  n_22148;
assign n_22151 = ~n_22149 & ~n_22150;
assign n_22152 =  x_742 &  n_21311;
assign n_22153 =  n_21310 &  n_22116;
assign n_22154 = ~n_22152 & ~n_22153;
assign n_22155 =  x_742 & ~n_22154;
assign n_22156 = ~x_742 &  n_22154;
assign n_22157 = ~n_22155 & ~n_22156;
assign n_22158 =  x_741 &  n_21293;
assign n_22159 =  n_21292 &  n_22116;
assign n_22160 = ~n_22158 & ~n_22159;
assign n_22161 =  x_741 & ~n_22160;
assign n_22162 = ~x_741 &  n_22160;
assign n_22163 = ~n_22161 & ~n_22162;
assign n_22164 =  x_740 &  n_21345;
assign n_22165 =  n_21344 &  n_22116;
assign n_22166 = ~n_22164 & ~n_22165;
assign n_22167 =  x_740 & ~n_22166;
assign n_22168 = ~x_740 &  n_22166;
assign n_22169 = ~n_22167 & ~n_22168;
assign n_22170 =  x_739 &  n_21378;
assign n_22171 =  n_21377 &  n_22116;
assign n_22172 = ~n_22170 & ~n_22171;
assign n_22173 =  x_739 & ~n_22172;
assign n_22174 = ~x_739 &  n_22172;
assign n_22175 = ~n_22173 & ~n_22174;
assign n_22176 =  x_738 &  n_21362;
assign n_22177 =  n_21361 &  n_22116;
assign n_22178 = ~n_22176 & ~n_22177;
assign n_22179 =  x_738 & ~n_22178;
assign n_22180 = ~x_738 &  n_22178;
assign n_22181 = ~n_22179 & ~n_22180;
assign n_22182 =  x_737 &  n_21353;
assign n_22183 =  n_21352 &  n_22116;
assign n_22184 = ~n_22182 & ~n_22183;
assign n_22185 =  x_737 & ~n_22184;
assign n_22186 = ~x_737 &  n_22184;
assign n_22187 = ~n_22185 & ~n_22186;
assign n_22188 =  x_736 &  n_21303;
assign n_22189 =  x_422 & ~n_3266;
assign n_22190 =  n_21302 &  n_22189;
assign n_22191 = ~n_22188 & ~n_22190;
assign n_22192 =  x_736 & ~n_22191;
assign n_22193 = ~x_736 &  n_22191;
assign n_22194 = ~n_22192 & ~n_22193;
assign n_22195 =  x_735 &  n_21311;
assign n_22196 =  n_21310 &  n_22189;
assign n_22197 = ~n_22195 & ~n_22196;
assign n_22198 =  x_735 & ~n_22197;
assign n_22199 = ~x_735 &  n_22197;
assign n_22200 = ~n_22198 & ~n_22199;
assign n_22201 =  x_734 &  n_21378;
assign n_22202 =  n_21377 &  n_22189;
assign n_22203 = ~n_22201 & ~n_22202;
assign n_22204 =  x_734 & ~n_22203;
assign n_22205 = ~x_734 &  n_22203;
assign n_22206 = ~n_22204 & ~n_22205;
assign n_22207 =  x_733 &  n_21337;
assign n_22208 =  n_21336 &  n_22189;
assign n_22209 = ~n_22207 & ~n_22208;
assign n_22210 =  x_733 & ~n_22209;
assign n_22211 = ~x_733 &  n_22209;
assign n_22212 = ~n_22210 & ~n_22211;
assign n_22213 =  x_732 &  n_21345;
assign n_22214 =  n_21344 &  n_22189;
assign n_22215 = ~n_22213 & ~n_22214;
assign n_22216 =  x_732 & ~n_22215;
assign n_22217 = ~x_732 &  n_22215;
assign n_22218 = ~n_22216 & ~n_22217;
assign n_22219 =  x_731 &  n_21362;
assign n_22220 =  n_21361 &  n_22189;
assign n_22221 = ~n_22219 & ~n_22220;
assign n_22222 =  x_731 & ~n_22221;
assign n_22223 = ~x_731 &  n_22221;
assign n_22224 = ~n_22222 & ~n_22223;
assign n_22225 =  x_730 &  n_21281;
assign n_22226 =  n_21280 &  n_22189;
assign n_22227 = ~n_22225 & ~n_22226;
assign n_22228 =  x_730 & ~n_22227;
assign n_22229 = ~x_730 &  n_22227;
assign n_22230 = ~n_22228 & ~n_22229;
assign n_22231 =  x_729 &  n_21370;
assign n_22232 =  n_21369 &  n_22189;
assign n_22233 = ~n_22231 & ~n_22232;
assign n_22234 =  x_729 & ~n_22233;
assign n_22235 = ~x_729 &  n_22233;
assign n_22236 = ~n_22234 & ~n_22235;
assign n_22237 =  x_728 &  n_21328;
assign n_22238 =  n_21327 &  n_22189;
assign n_22239 = ~n_22237 & ~n_22238;
assign n_22240 =  x_728 & ~n_22239;
assign n_22241 = ~x_728 &  n_22239;
assign n_22242 = ~n_22240 & ~n_22241;
assign n_22243 =  x_727 &  n_21319;
assign n_22244 =  n_21318 &  n_22189;
assign n_22245 = ~n_22243 & ~n_22244;
assign n_22246 =  x_727 & ~n_22245;
assign n_22247 = ~x_727 &  n_22245;
assign n_22248 = ~n_22246 & ~n_22247;
assign n_22249 =  x_726 &  n_21293;
assign n_22250 =  n_21292 &  n_22189;
assign n_22251 = ~n_22249 & ~n_22250;
assign n_22252 =  x_726 & ~n_22251;
assign n_22253 = ~x_726 &  n_22251;
assign n_22254 = ~n_22252 & ~n_22253;
assign n_22255 =  x_725 &  n_21353;
assign n_22256 =  n_21352 &  n_22189;
assign n_22257 = ~n_22255 & ~n_22256;
assign n_22258 =  x_725 & ~n_22257;
assign n_22259 = ~x_725 &  n_22257;
assign n_22260 = ~n_22258 & ~n_22259;
assign n_22261 =  x_724 &  n_21378;
assign n_22262 =  x_421 & ~n_3266;
assign n_22263 =  n_21377 &  n_22262;
assign n_22264 = ~n_22261 & ~n_22263;
assign n_22265 =  x_724 & ~n_22264;
assign n_22266 = ~x_724 &  n_22264;
assign n_22267 = ~n_22265 & ~n_22266;
assign n_22268 =  x_723 &  n_21337;
assign n_22269 =  n_21336 &  n_22262;
assign n_22270 = ~n_22268 & ~n_22269;
assign n_22271 =  x_723 & ~n_22270;
assign n_22272 = ~x_723 &  n_22270;
assign n_22273 = ~n_22271 & ~n_22272;
assign n_22274 =  x_722 &  n_21328;
assign n_22275 =  n_21327 &  n_22262;
assign n_22276 = ~n_22274 & ~n_22275;
assign n_22277 =  x_722 & ~n_22276;
assign n_22278 = ~x_722 &  n_22276;
assign n_22279 = ~n_22277 & ~n_22278;
assign n_22280 =  x_721 &  n_21303;
assign n_22281 =  n_21302 &  n_22262;
assign n_22282 = ~n_22280 & ~n_22281;
assign n_22283 =  x_721 & ~n_22282;
assign n_22284 = ~x_721 &  n_22282;
assign n_22285 = ~n_22283 & ~n_22284;
assign n_22286 =  x_720 &  n_21362;
assign n_22287 =  n_21361 &  n_22262;
assign n_22288 = ~n_22286 & ~n_22287;
assign n_22289 =  x_720 & ~n_22288;
assign n_22290 = ~x_720 &  n_22288;
assign n_22291 = ~n_22289 & ~n_22290;
assign n_22292 =  x_719 &  n_21293;
assign n_22293 =  n_21292 &  n_22262;
assign n_22294 = ~n_22292 & ~n_22293;
assign n_22295 =  x_719 & ~n_22294;
assign n_22296 = ~x_719 &  n_22294;
assign n_22297 = ~n_22295 & ~n_22296;
assign n_22298 =  x_718 &  n_21345;
assign n_22299 =  n_21344 &  n_22262;
assign n_22300 = ~n_22298 & ~n_22299;
assign n_22301 =  x_718 & ~n_22300;
assign n_22302 = ~x_718 &  n_22300;
assign n_22303 = ~n_22301 & ~n_22302;
assign n_22304 =  x_717 &  n_21353;
assign n_22305 =  n_21352 &  n_22262;
assign n_22306 = ~n_22304 & ~n_22305;
assign n_22307 =  x_717 & ~n_22306;
assign n_22308 = ~x_717 &  n_22306;
assign n_22309 = ~n_22307 & ~n_22308;
assign n_22310 =  x_716 &  n_21319;
assign n_22311 =  n_21318 &  n_22262;
assign n_22312 = ~n_22310 & ~n_22311;
assign n_22313 =  x_716 & ~n_22312;
assign n_22314 = ~x_716 &  n_22312;
assign n_22315 = ~n_22313 & ~n_22314;
assign n_22316 =  x_715 &  n_21370;
assign n_22317 =  n_21369 &  n_22262;
assign n_22318 = ~n_22316 & ~n_22317;
assign n_22319 =  x_715 & ~n_22318;
assign n_22320 = ~x_715 &  n_22318;
assign n_22321 = ~n_22319 & ~n_22320;
assign n_22322 =  x_714 &  n_21281;
assign n_22323 =  n_21280 &  n_22262;
assign n_22324 = ~n_22322 & ~n_22323;
assign n_22325 =  x_714 & ~n_22324;
assign n_22326 = ~x_714 &  n_22324;
assign n_22327 = ~n_22325 & ~n_22326;
assign n_22328 =  x_713 &  n_21311;
assign n_22329 =  n_21310 &  n_22262;
assign n_22330 = ~n_22328 & ~n_22329;
assign n_22331 =  x_713 & ~n_22330;
assign n_22332 = ~x_713 &  n_22330;
assign n_22333 = ~n_22331 & ~n_22332;
assign n_22334 =  x_712 &  n_21370;
assign n_22335 =  x_420 & ~n_3266;
assign n_22336 =  n_21369 &  n_22335;
assign n_22337 = ~n_22334 & ~n_22336;
assign n_22338 =  x_712 & ~n_22337;
assign n_22339 = ~x_712 &  n_22337;
assign n_22340 = ~n_22338 & ~n_22339;
assign n_22341 =  x_711 &  n_21353;
assign n_22342 =  n_21352 &  n_22335;
assign n_22343 = ~n_22341 & ~n_22342;
assign n_22344 =  x_711 & ~n_22343;
assign n_22345 = ~x_711 &  n_22343;
assign n_22346 = ~n_22344 & ~n_22345;
assign n_22347 =  x_710 &  n_21328;
assign n_22348 =  n_21327 &  n_22335;
assign n_22349 = ~n_22347 & ~n_22348;
assign n_22350 =  x_710 & ~n_22349;
assign n_22351 = ~x_710 &  n_22349;
assign n_22352 = ~n_22350 & ~n_22351;
assign n_22353 =  x_709 &  n_21378;
assign n_22354 =  n_21377 &  n_22335;
assign n_22355 = ~n_22353 & ~n_22354;
assign n_22356 =  x_709 & ~n_22355;
assign n_22357 = ~x_709 &  n_22355;
assign n_22358 = ~n_22356 & ~n_22357;
assign n_22359 =  x_708 &  n_21319;
assign n_22360 =  n_21318 &  n_22335;
assign n_22361 = ~n_22359 & ~n_22360;
assign n_22362 =  x_708 & ~n_22361;
assign n_22363 = ~x_708 &  n_22361;
assign n_22364 = ~n_22362 & ~n_22363;
assign n_22365 =  x_707 &  n_21293;
assign n_22366 =  n_21292 &  n_22335;
assign n_22367 = ~n_22365 & ~n_22366;
assign n_22368 =  x_707 & ~n_22367;
assign n_22369 = ~x_707 &  n_22367;
assign n_22370 = ~n_22368 & ~n_22369;
assign n_22371 =  x_706 &  n_21303;
assign n_22372 =  n_21302 &  n_22335;
assign n_22373 = ~n_22371 & ~n_22372;
assign n_22374 =  x_706 & ~n_22373;
assign n_22375 = ~x_706 &  n_22373;
assign n_22376 = ~n_22374 & ~n_22375;
assign n_22377 =  x_705 &  n_21337;
assign n_22378 =  n_21336 &  n_22335;
assign n_22379 = ~n_22377 & ~n_22378;
assign n_22380 =  x_705 & ~n_22379;
assign n_22381 = ~x_705 &  n_22379;
assign n_22382 = ~n_22380 & ~n_22381;
assign n_22383 =  x_704 &  n_21345;
assign n_22384 =  n_21344 &  n_22335;
assign n_22385 = ~n_22383 & ~n_22384;
assign n_22386 =  x_704 & ~n_22385;
assign n_22387 = ~x_704 &  n_22385;
assign n_22388 = ~n_22386 & ~n_22387;
assign n_22389 =  x_703 &  n_21362;
assign n_22390 =  n_21361 &  n_22335;
assign n_22391 = ~n_22389 & ~n_22390;
assign n_22392 =  x_703 & ~n_22391;
assign n_22393 = ~x_703 &  n_22391;
assign n_22394 = ~n_22392 & ~n_22393;
assign n_22395 =  x_702 &  n_21281;
assign n_22396 =  n_21280 &  n_22335;
assign n_22397 = ~n_22395 & ~n_22396;
assign n_22398 =  x_702 & ~n_22397;
assign n_22399 = ~x_702 &  n_22397;
assign n_22400 = ~n_22398 & ~n_22399;
assign n_22401 =  x_701 &  n_21311;
assign n_22402 =  n_21310 &  n_22335;
assign n_22403 = ~n_22401 & ~n_22402;
assign n_22404 =  x_701 & ~n_22403;
assign n_22405 = ~x_701 &  n_22403;
assign n_22406 = ~n_22404 & ~n_22405;
assign n_22407 =  x_700 &  n_21378;
assign n_22408 =  x_419 & ~n_3266;
assign n_22409 =  n_21377 &  n_22408;
assign n_22410 = ~n_22407 & ~n_22409;
assign n_22411 =  x_700 & ~n_22410;
assign n_22412 = ~x_700 &  n_22410;
assign n_22413 = ~n_22411 & ~n_22412;
assign n_22414 =  x_699 &  n_21362;
assign n_22415 =  n_21361 &  n_22408;
assign n_22416 = ~n_22414 & ~n_22415;
assign n_22417 =  x_699 & ~n_22416;
assign n_22418 = ~x_699 &  n_22416;
assign n_22419 = ~n_22417 & ~n_22418;
assign n_22420 =  x_698 &  n_21293;
assign n_22421 =  n_21292 &  n_22408;
assign n_22422 = ~n_22420 & ~n_22421;
assign n_22423 =  x_698 & ~n_22422;
assign n_22424 = ~x_698 &  n_22422;
assign n_22425 = ~n_22423 & ~n_22424;
assign n_22426 =  x_697 &  n_21311;
assign n_22427 =  n_21310 &  n_22408;
assign n_22428 = ~n_22426 & ~n_22427;
assign n_22429 =  x_697 & ~n_22428;
assign n_22430 = ~x_697 &  n_22428;
assign n_22431 = ~n_22429 & ~n_22430;
assign n_22432 =  x_696 &  n_21337;
assign n_22433 =  n_21336 &  n_22408;
assign n_22434 = ~n_22432 & ~n_22433;
assign n_22435 =  x_696 & ~n_22434;
assign n_22436 = ~x_696 &  n_22434;
assign n_22437 = ~n_22435 & ~n_22436;
assign n_22438 =  x_695 &  n_21328;
assign n_22439 =  n_21327 &  n_22408;
assign n_22440 = ~n_22438 & ~n_22439;
assign n_22441 =  x_695 & ~n_22440;
assign n_22442 = ~x_695 &  n_22440;
assign n_22443 = ~n_22441 & ~n_22442;
assign n_22444 =  x_694 &  n_21345;
assign n_22445 =  n_21344 &  n_22408;
assign n_22446 = ~n_22444 & ~n_22445;
assign n_22447 =  x_694 & ~n_22446;
assign n_22448 = ~x_694 &  n_22446;
assign n_22449 = ~n_22447 & ~n_22448;
assign n_22450 =  x_693 &  n_21319;
assign n_22451 =  n_21318 &  n_22408;
assign n_22452 = ~n_22450 & ~n_22451;
assign n_22453 =  x_693 & ~n_22452;
assign n_22454 = ~x_693 &  n_22452;
assign n_22455 = ~n_22453 & ~n_22454;
assign n_22456 =  x_692 &  n_21303;
assign n_22457 =  n_21302 &  n_22408;
assign n_22458 = ~n_22456 & ~n_22457;
assign n_22459 =  x_692 & ~n_22458;
assign n_22460 = ~x_692 &  n_22458;
assign n_22461 = ~n_22459 & ~n_22460;
assign n_22462 =  x_691 &  n_21353;
assign n_22463 =  n_21352 &  n_22408;
assign n_22464 = ~n_22462 & ~n_22463;
assign n_22465 =  x_691 & ~n_22464;
assign n_22466 = ~x_691 &  n_22464;
assign n_22467 = ~n_22465 & ~n_22466;
assign n_22468 =  x_690 &  n_21370;
assign n_22469 =  n_21369 &  n_22408;
assign n_22470 = ~n_22468 & ~n_22469;
assign n_22471 =  x_690 & ~n_22470;
assign n_22472 = ~x_690 &  n_22470;
assign n_22473 = ~n_22471 & ~n_22472;
assign n_22474 =  x_689 &  n_21281;
assign n_22475 =  n_21280 &  n_22408;
assign n_22476 = ~n_22474 & ~n_22475;
assign n_22477 =  x_689 & ~n_22476;
assign n_22478 = ~x_689 &  n_22476;
assign n_22479 = ~n_22477 & ~n_22478;
assign n_22480 =  x_688 &  n_21281;
assign n_22481 =  x_418 & ~n_3266;
assign n_22482 =  n_21280 &  n_22481;
assign n_22483 = ~n_22480 & ~n_22482;
assign n_22484 =  x_688 & ~n_22483;
assign n_22485 = ~x_688 &  n_22483;
assign n_22486 = ~n_22484 & ~n_22485;
assign n_22487 =  x_687 &  n_21378;
assign n_22488 =  n_21377 &  n_22481;
assign n_22489 = ~n_22487 & ~n_22488;
assign n_22490 =  x_687 & ~n_22489;
assign n_22491 = ~x_687 &  n_22489;
assign n_22492 = ~n_22490 & ~n_22491;
assign n_22493 =  x_686 &  n_21353;
assign n_22494 =  n_21352 &  n_22481;
assign n_22495 = ~n_22493 & ~n_22494;
assign n_22496 =  x_686 & ~n_22495;
assign n_22497 = ~x_686 &  n_22495;
assign n_22498 = ~n_22496 & ~n_22497;
assign n_22499 =  x_685 &  n_21319;
assign n_22500 =  n_21318 &  n_22481;
assign n_22501 = ~n_22499 & ~n_22500;
assign n_22502 =  x_685 & ~n_22501;
assign n_22503 = ~x_685 &  n_22501;
assign n_22504 = ~n_22502 & ~n_22503;
assign n_22505 =  x_684 &  n_21303;
assign n_22506 =  n_21302 &  n_22481;
assign n_22507 = ~n_22505 & ~n_22506;
assign n_22508 =  x_684 & ~n_22507;
assign n_22509 = ~x_684 &  n_22507;
assign n_22510 = ~n_22508 & ~n_22509;
assign n_22511 =  x_683 &  n_21370;
assign n_22512 =  n_21369 &  n_22481;
assign n_22513 = ~n_22511 & ~n_22512;
assign n_22514 =  x_683 & ~n_22513;
assign n_22515 = ~x_683 &  n_22513;
assign n_22516 = ~n_22514 & ~n_22515;
assign n_22517 =  x_682 &  n_21337;
assign n_22518 =  n_21336 &  n_22481;
assign n_22519 = ~n_22517 & ~n_22518;
assign n_22520 =  x_682 & ~n_22519;
assign n_22521 = ~x_682 &  n_22519;
assign n_22522 = ~n_22520 & ~n_22521;
assign n_22523 =  x_681 &  n_21345;
assign n_22524 =  n_21344 &  n_22481;
assign n_22525 = ~n_22523 & ~n_22524;
assign n_22526 =  x_681 & ~n_22525;
assign n_22527 = ~x_681 &  n_22525;
assign n_22528 = ~n_22526 & ~n_22527;
assign n_22529 =  x_680 &  n_21328;
assign n_22530 =  n_21327 &  n_22481;
assign n_22531 = ~n_22529 & ~n_22530;
assign n_22532 =  x_680 & ~n_22531;
assign n_22533 = ~x_680 &  n_22531;
assign n_22534 = ~n_22532 & ~n_22533;
assign n_22535 =  x_679 &  n_21293;
assign n_22536 =  n_21292 &  n_22481;
assign n_22537 = ~n_22535 & ~n_22536;
assign n_22538 =  x_679 & ~n_22537;
assign n_22539 = ~x_679 &  n_22537;
assign n_22540 = ~n_22538 & ~n_22539;
assign n_22541 =  x_678 &  n_21362;
assign n_22542 =  n_21361 &  n_22481;
assign n_22543 = ~n_22541 & ~n_22542;
assign n_22544 =  x_678 & ~n_22543;
assign n_22545 = ~x_678 &  n_22543;
assign n_22546 = ~n_22544 & ~n_22545;
assign n_22547 =  x_677 &  n_21311;
assign n_22548 =  n_21310 &  n_22481;
assign n_22549 = ~n_22547 & ~n_22548;
assign n_22550 =  x_677 & ~n_22549;
assign n_22551 = ~x_677 &  n_22549;
assign n_22552 = ~n_22550 & ~n_22551;
assign n_22553 =  x_676 &  n_21281;
assign n_22554 =  x_417 & ~n_3266;
assign n_22555 =  n_21280 &  n_22554;
assign n_22556 = ~n_22553 & ~n_22555;
assign n_22557 =  x_676 & ~n_22556;
assign n_22558 = ~x_676 &  n_22556;
assign n_22559 = ~n_22557 & ~n_22558;
assign n_22560 =  x_675 &  n_21378;
assign n_22561 =  n_21377 &  n_22554;
assign n_22562 = ~n_22560 & ~n_22561;
assign n_22563 =  x_675 & ~n_22562;
assign n_22564 = ~x_675 &  n_22562;
assign n_22565 = ~n_22563 & ~n_22564;
assign n_22566 =  x_674 &  n_21293;
assign n_22567 =  n_21292 &  n_22554;
assign n_22568 = ~n_22566 & ~n_22567;
assign n_22569 =  x_674 & ~n_22568;
assign n_22570 = ~x_674 &  n_22568;
assign n_22571 = ~n_22569 & ~n_22570;
assign n_22572 =  x_673 &  n_21311;
assign n_22573 =  n_21310 &  n_22554;
assign n_22574 = ~n_22572 & ~n_22573;
assign n_22575 =  x_673 & ~n_22574;
assign n_22576 = ~x_673 &  n_22574;
assign n_22577 = ~n_22575 & ~n_22576;
assign n_22578 =  x_672 &  n_21303;
assign n_22579 =  n_21302 &  n_22554;
assign n_22580 = ~n_22578 & ~n_22579;
assign n_22581 =  x_672 & ~n_22580;
assign n_22582 = ~x_672 &  n_22580;
assign n_22583 = ~n_22581 & ~n_22582;
assign n_22584 =  x_671 &  n_21328;
assign n_22585 =  n_21327 &  n_22554;
assign n_22586 = ~n_22584 & ~n_22585;
assign n_22587 =  x_671 & ~n_22586;
assign n_22588 = ~x_671 &  n_22586;
assign n_22589 = ~n_22587 & ~n_22588;
assign n_22590 =  x_670 &  n_21353;
assign n_22591 =  n_21352 &  n_22554;
assign n_22592 = ~n_22590 & ~n_22591;
assign n_22593 =  x_670 & ~n_22592;
assign n_22594 = ~x_670 &  n_22592;
assign n_22595 = ~n_22593 & ~n_22594;
assign n_22596 =  x_669 &  n_21337;
assign n_22597 =  n_21336 &  n_22554;
assign n_22598 = ~n_22596 & ~n_22597;
assign n_22599 =  x_669 & ~n_22598;
assign n_22600 = ~x_669 &  n_22598;
assign n_22601 = ~n_22599 & ~n_22600;
assign n_22602 =  x_668 &  n_21319;
assign n_22603 =  n_21318 &  n_22554;
assign n_22604 = ~n_22602 & ~n_22603;
assign n_22605 =  x_668 & ~n_22604;
assign n_22606 = ~x_668 &  n_22604;
assign n_22607 = ~n_22605 & ~n_22606;
assign n_22608 =  x_667 &  n_21370;
assign n_22609 =  n_21369 &  n_22554;
assign n_22610 = ~n_22608 & ~n_22609;
assign n_22611 =  x_667 & ~n_22610;
assign n_22612 = ~x_667 &  n_22610;
assign n_22613 = ~n_22611 & ~n_22612;
assign n_22614 =  x_666 &  n_21345;
assign n_22615 =  n_21344 &  n_22554;
assign n_22616 = ~n_22614 & ~n_22615;
assign n_22617 =  x_666 & ~n_22616;
assign n_22618 = ~x_666 &  n_22616;
assign n_22619 = ~n_22617 & ~n_22618;
assign n_22620 =  x_665 &  n_21362;
assign n_22621 =  n_21361 &  n_22554;
assign n_22622 = ~n_22620 & ~n_22621;
assign n_22623 =  x_665 & ~n_22622;
assign n_22624 = ~x_665 &  n_22622;
assign n_22625 = ~n_22623 & ~n_22624;
assign n_22626 =  x_664 &  n_21328;
assign n_22627 =  x_416 & ~n_3266;
assign n_22628 =  n_21327 &  n_22627;
assign n_22629 = ~n_22626 & ~n_22628;
assign n_22630 =  x_664 & ~n_22629;
assign n_22631 = ~x_664 &  n_22629;
assign n_22632 = ~n_22630 & ~n_22631;
assign n_22633 =  x_663 &  n_21319;
assign n_22634 =  n_21318 &  n_22627;
assign n_22635 = ~n_22633 & ~n_22634;
assign n_22636 =  x_663 & ~n_22635;
assign n_22637 = ~x_663 &  n_22635;
assign n_22638 = ~n_22636 & ~n_22637;
assign n_22639 =  x_662 &  n_21378;
assign n_22640 =  n_21377 &  n_22627;
assign n_22641 = ~n_22639 & ~n_22640;
assign n_22642 =  x_662 & ~n_22641;
assign n_22643 = ~x_662 &  n_22641;
assign n_22644 = ~n_22642 & ~n_22643;
assign n_22645 =  x_661 &  n_21311;
assign n_22646 =  n_21310 &  n_22627;
assign n_22647 = ~n_22645 & ~n_22646;
assign n_22648 =  x_661 & ~n_22647;
assign n_22649 = ~x_661 &  n_22647;
assign n_22650 = ~n_22648 & ~n_22649;
assign n_22651 =  x_660 &  n_21345;
assign n_22652 =  n_21344 &  n_22627;
assign n_22653 = ~n_22651 & ~n_22652;
assign n_22654 =  x_660 & ~n_22653;
assign n_22655 = ~x_660 &  n_22653;
assign n_22656 = ~n_22654 & ~n_22655;
assign n_22657 =  x_659 &  n_21353;
assign n_22658 =  n_21352 &  n_22627;
assign n_22659 = ~n_22657 & ~n_22658;
assign n_22660 =  x_659 & ~n_22659;
assign n_22661 = ~x_659 &  n_22659;
assign n_22662 = ~n_22660 & ~n_22661;
assign n_22663 =  x_658 &  n_21370;
assign n_22664 =  n_21369 &  n_22627;
assign n_22665 = ~n_22663 & ~n_22664;
assign n_22666 =  x_658 & ~n_22665;
assign n_22667 = ~x_658 &  n_22665;
assign n_22668 = ~n_22666 & ~n_22667;
assign n_22669 =  x_657 &  n_21303;
assign n_22670 =  n_21302 &  n_22627;
assign n_22671 = ~n_22669 & ~n_22670;
assign n_22672 =  x_657 & ~n_22671;
assign n_22673 = ~x_657 &  n_22671;
assign n_22674 = ~n_22672 & ~n_22673;
assign n_22675 =  x_656 &  n_21293;
assign n_22676 =  n_21292 &  n_22627;
assign n_22677 = ~n_22675 & ~n_22676;
assign n_22678 =  x_656 & ~n_22677;
assign n_22679 = ~x_656 &  n_22677;
assign n_22680 = ~n_22678 & ~n_22679;
assign n_22681 =  x_655 &  n_21362;
assign n_22682 =  n_21361 &  n_22627;
assign n_22683 = ~n_22681 & ~n_22682;
assign n_22684 =  x_655 & ~n_22683;
assign n_22685 = ~x_655 &  n_22683;
assign n_22686 = ~n_22684 & ~n_22685;
assign n_22687 =  x_654 &  n_21281;
assign n_22688 =  n_21280 &  n_22627;
assign n_22689 = ~n_22687 & ~n_22688;
assign n_22690 =  x_654 & ~n_22689;
assign n_22691 = ~x_654 &  n_22689;
assign n_22692 = ~n_22690 & ~n_22691;
assign n_22693 =  x_653 &  n_21337;
assign n_22694 =  n_21336 &  n_22627;
assign n_22695 = ~n_22693 & ~n_22694;
assign n_22696 =  x_653 & ~n_22695;
assign n_22697 = ~x_653 &  n_22695;
assign n_22698 = ~n_22696 & ~n_22697;
assign n_22699 =  x_652 &  n_21311;
assign n_22700 =  x_415 & ~n_3266;
assign n_22701 =  n_21310 &  n_22700;
assign n_22702 = ~n_22699 & ~n_22701;
assign n_22703 =  x_652 & ~n_22702;
assign n_22704 = ~x_652 &  n_22702;
assign n_22705 = ~n_22703 & ~n_22704;
assign n_22706 =  x_651 &  n_21328;
assign n_22707 =  n_21327 &  n_22700;
assign n_22708 = ~n_22706 & ~n_22707;
assign n_22709 =  x_651 & ~n_22708;
assign n_22710 = ~x_651 &  n_22708;
assign n_22711 = ~n_22709 & ~n_22710;
assign n_22712 =  x_650 &  n_21378;
assign n_22713 =  n_21377 &  n_22700;
assign n_22714 = ~n_22712 & ~n_22713;
assign n_22715 =  x_650 & ~n_22714;
assign n_22716 = ~x_650 &  n_22714;
assign n_22717 = ~n_22715 & ~n_22716;
assign n_22718 =  x_649 &  n_21281;
assign n_22719 =  n_21280 &  n_22700;
assign n_22720 = ~n_22718 & ~n_22719;
assign n_22721 =  x_649 & ~n_22720;
assign n_22722 = ~x_649 &  n_22720;
assign n_22723 = ~n_22721 & ~n_22722;
assign n_22724 =  x_648 &  n_21362;
assign n_22725 =  n_21361 &  n_22700;
assign n_22726 = ~n_22724 & ~n_22725;
assign n_22727 =  x_648 & ~n_22726;
assign n_22728 = ~x_648 &  n_22726;
assign n_22729 = ~n_22727 & ~n_22728;
assign n_22730 =  x_647 &  n_21353;
assign n_22731 =  n_21352 &  n_22700;
assign n_22732 = ~n_22730 & ~n_22731;
assign n_22733 =  x_647 & ~n_22732;
assign n_22734 = ~x_647 &  n_22732;
assign n_22735 = ~n_22733 & ~n_22734;
assign n_22736 =  x_646 &  n_21293;
assign n_22737 =  n_21292 &  n_22700;
assign n_22738 = ~n_22736 & ~n_22737;
assign n_22739 =  x_646 & ~n_22738;
assign n_22740 = ~x_646 &  n_22738;
assign n_22741 = ~n_22739 & ~n_22740;
assign n_22742 =  x_645 &  n_21337;
assign n_22743 =  n_21336 &  n_22700;
assign n_22744 = ~n_22742 & ~n_22743;
assign n_22745 =  x_645 & ~n_22744;
assign n_22746 = ~x_645 &  n_22744;
assign n_22747 = ~n_22745 & ~n_22746;
assign n_22748 =  x_644 &  n_21303;
assign n_22749 =  n_21302 &  n_22700;
assign n_22750 = ~n_22748 & ~n_22749;
assign n_22751 =  x_644 & ~n_22750;
assign n_22752 = ~x_644 &  n_22750;
assign n_22753 = ~n_22751 & ~n_22752;
assign n_22754 =  x_643 &  n_21345;
assign n_22755 =  n_21344 &  n_22700;
assign n_22756 = ~n_22754 & ~n_22755;
assign n_22757 =  x_643 & ~n_22756;
assign n_22758 = ~x_643 &  n_22756;
assign n_22759 = ~n_22757 & ~n_22758;
assign n_22760 =  x_642 &  n_21319;
assign n_22761 =  n_21318 &  n_22700;
assign n_22762 = ~n_22760 & ~n_22761;
assign n_22763 =  x_642 & ~n_22762;
assign n_22764 = ~x_642 &  n_22762;
assign n_22765 = ~n_22763 & ~n_22764;
assign n_22766 =  x_641 &  n_21370;
assign n_22767 =  n_21369 &  n_22700;
assign n_22768 = ~n_22766 & ~n_22767;
assign n_22769 =  x_641 & ~n_22768;
assign n_22770 = ~x_641 &  n_22768;
assign n_22771 = ~n_22769 & ~n_22770;
assign n_22772 =  x_640 &  n_21303;
assign n_22773 =  x_414 & ~n_3266;
assign n_22774 =  n_21302 &  n_22773;
assign n_22775 = ~n_22772 & ~n_22774;
assign n_22776 =  x_640 & ~n_22775;
assign n_22777 = ~x_640 &  n_22775;
assign n_22778 = ~n_22776 & ~n_22777;
assign n_22779 =  x_639 &  n_21345;
assign n_22780 =  n_21344 &  n_22773;
assign n_22781 = ~n_22779 & ~n_22780;
assign n_22782 =  x_639 & ~n_22781;
assign n_22783 = ~x_639 &  n_22781;
assign n_22784 = ~n_22782 & ~n_22783;
assign n_22785 =  x_638 &  n_21370;
assign n_22786 =  n_21369 &  n_22773;
assign n_22787 = ~n_22785 & ~n_22786;
assign n_22788 =  x_638 & ~n_22787;
assign n_22789 = ~x_638 &  n_22787;
assign n_22790 = ~n_22788 & ~n_22789;
assign n_22791 =  x_637 &  n_21353;
assign n_22792 =  n_21352 &  n_22773;
assign n_22793 = ~n_22791 & ~n_22792;
assign n_22794 =  x_637 & ~n_22793;
assign n_22795 = ~x_637 &  n_22793;
assign n_22796 = ~n_22794 & ~n_22795;
assign n_22797 =  x_636 &  n_21311;
assign n_22798 =  n_21310 &  n_22773;
assign n_22799 = ~n_22797 & ~n_22798;
assign n_22800 =  x_636 & ~n_22799;
assign n_22801 = ~x_636 &  n_22799;
assign n_22802 = ~n_22800 & ~n_22801;
assign n_22803 =  x_635 &  n_21328;
assign n_22804 =  n_21327 &  n_22773;
assign n_22805 = ~n_22803 & ~n_22804;
assign n_22806 =  x_635 & ~n_22805;
assign n_22807 = ~x_635 &  n_22805;
assign n_22808 = ~n_22806 & ~n_22807;
assign n_22809 =  x_634 &  n_21378;
assign n_22810 =  n_21377 &  n_22773;
assign n_22811 = ~n_22809 & ~n_22810;
assign n_22812 =  x_634 & ~n_22811;
assign n_22813 = ~x_634 &  n_22811;
assign n_22814 = ~n_22812 & ~n_22813;
assign n_22815 =  x_633 &  n_21293;
assign n_22816 =  n_21292 &  n_22773;
assign n_22817 = ~n_22815 & ~n_22816;
assign n_22818 =  x_633 & ~n_22817;
assign n_22819 = ~x_633 &  n_22817;
assign n_22820 = ~n_22818 & ~n_22819;
assign n_22821 =  x_632 &  n_21319;
assign n_22822 =  n_21318 &  n_22773;
assign n_22823 = ~n_22821 & ~n_22822;
assign n_22824 =  x_632 & ~n_22823;
assign n_22825 = ~x_632 &  n_22823;
assign n_22826 = ~n_22824 & ~n_22825;
assign n_22827 =  x_631 &  n_21362;
assign n_22828 =  n_21361 &  n_22773;
assign n_22829 = ~n_22827 & ~n_22828;
assign n_22830 =  x_631 & ~n_22829;
assign n_22831 = ~x_631 &  n_22829;
assign n_22832 = ~n_22830 & ~n_22831;
assign n_22833 =  x_630 &  n_21281;
assign n_22834 =  n_21280 &  n_22773;
assign n_22835 = ~n_22833 & ~n_22834;
assign n_22836 =  x_630 & ~n_22835;
assign n_22837 = ~x_630 &  n_22835;
assign n_22838 = ~n_22836 & ~n_22837;
assign n_22839 =  x_629 &  n_21337;
assign n_22840 =  n_21336 &  n_22773;
assign n_22841 = ~n_22839 & ~n_22840;
assign n_22842 =  x_629 & ~n_22841;
assign n_22843 = ~x_629 &  n_22841;
assign n_22844 = ~n_22842 & ~n_22843;
assign n_22845 =  x_628 &  n_21378;
assign n_22846 =  x_413 & ~n_3266;
assign n_22847 =  n_21377 &  n_22846;
assign n_22848 = ~n_22845 & ~n_22847;
assign n_22849 =  x_628 & ~n_22848;
assign n_22850 = ~x_628 &  n_22848;
assign n_22851 = ~n_22849 & ~n_22850;
assign n_22852 =  x_627 &  n_21362;
assign n_22853 =  n_21361 &  n_22846;
assign n_22854 = ~n_22852 & ~n_22853;
assign n_22855 =  x_627 & ~n_22854;
assign n_22856 = ~x_627 &  n_22854;
assign n_22857 = ~n_22855 & ~n_22856;
assign n_22858 =  x_626 &  n_21311;
assign n_22859 =  n_21310 &  n_22846;
assign n_22860 = ~n_22858 & ~n_22859;
assign n_22861 =  x_626 & ~n_22860;
assign n_22862 = ~x_626 &  n_22860;
assign n_22863 = ~n_22861 & ~n_22862;
assign n_22864 =  x_625 &  n_21303;
assign n_22865 =  n_21302 &  n_22846;
assign n_22866 = ~n_22864 & ~n_22865;
assign n_22867 =  x_625 & ~n_22866;
assign n_22868 = ~x_625 &  n_22866;
assign n_22869 = ~n_22867 & ~n_22868;
assign n_22870 =  x_624 &  n_21345;
assign n_22871 =  n_21344 &  n_22846;
assign n_22872 = ~n_22870 & ~n_22871;
assign n_22873 =  x_624 & ~n_22872;
assign n_22874 = ~x_624 &  n_22872;
assign n_22875 = ~n_22873 & ~n_22874;
assign n_22876 =  x_623 &  n_21293;
assign n_22877 =  n_21292 &  n_22846;
assign n_22878 = ~n_22876 & ~n_22877;
assign n_22879 =  x_623 & ~n_22878;
assign n_22880 = ~x_623 &  n_22878;
assign n_22881 = ~n_22879 & ~n_22880;
assign n_22882 =  x_622 &  n_21319;
assign n_22883 =  n_21318 &  n_22846;
assign n_22884 = ~n_22882 & ~n_22883;
assign n_22885 =  x_622 & ~n_22884;
assign n_22886 = ~x_622 &  n_22884;
assign n_22887 = ~n_22885 & ~n_22886;
assign n_22888 =  x_621 &  n_21353;
assign n_22889 =  n_21352 &  n_22846;
assign n_22890 = ~n_22888 & ~n_22889;
assign n_22891 =  x_621 & ~n_22890;
assign n_22892 = ~x_621 &  n_22890;
assign n_22893 = ~n_22891 & ~n_22892;
assign n_22894 =  x_620 &  n_21370;
assign n_22895 =  n_21369 &  n_22846;
assign n_22896 = ~n_22894 & ~n_22895;
assign n_22897 =  x_620 & ~n_22896;
assign n_22898 = ~x_620 &  n_22896;
assign n_22899 = ~n_22897 & ~n_22898;
assign n_22900 =  x_619 &  n_21281;
assign n_22901 =  n_21280 &  n_22846;
assign n_22902 = ~n_22900 & ~n_22901;
assign n_22903 =  x_619 & ~n_22902;
assign n_22904 = ~x_619 &  n_22902;
assign n_22905 = ~n_22903 & ~n_22904;
assign n_22906 =  x_618 &  n_21328;
assign n_22907 =  n_21327 &  n_22846;
assign n_22908 = ~n_22906 & ~n_22907;
assign n_22909 =  x_618 & ~n_22908;
assign n_22910 = ~x_618 &  n_22908;
assign n_22911 = ~n_22909 & ~n_22910;
assign n_22912 =  x_617 &  n_21337;
assign n_22913 =  n_21336 &  n_22846;
assign n_22914 = ~n_22912 & ~n_22913;
assign n_22915 =  x_617 & ~n_22914;
assign n_22916 = ~x_617 &  n_22914;
assign n_22917 = ~n_22915 & ~n_22916;
assign n_22918 =  x_616 &  n_21362;
assign n_22919 =  x_412 & ~n_3266;
assign n_22920 =  n_21361 &  n_22919;
assign n_22921 = ~n_22918 & ~n_22920;
assign n_22922 =  x_616 & ~n_22921;
assign n_22923 = ~x_616 &  n_22921;
assign n_22924 = ~n_22922 & ~n_22923;
assign n_22925 =  x_615 &  n_21328;
assign n_22926 =  n_21327 &  n_22919;
assign n_22927 = ~n_22925 & ~n_22926;
assign n_22928 =  x_615 & ~n_22927;
assign n_22929 = ~x_615 &  n_22927;
assign n_22930 = ~n_22928 & ~n_22929;
assign n_22931 =  x_614 &  n_21353;
assign n_22932 =  n_21352 &  n_22919;
assign n_22933 = ~n_22931 & ~n_22932;
assign n_22934 =  x_614 & ~n_22933;
assign n_22935 = ~x_614 &  n_22933;
assign n_22936 = ~n_22934 & ~n_22935;
assign n_22937 =  x_613 &  n_21293;
assign n_22938 =  n_21292 &  n_22919;
assign n_22939 = ~n_22937 & ~n_22938;
assign n_22940 =  x_613 & ~n_22939;
assign n_22941 = ~x_613 &  n_22939;
assign n_22942 = ~n_22940 & ~n_22941;
assign n_22943 =  x_612 &  n_21319;
assign n_22944 =  n_21318 &  n_22919;
assign n_22945 = ~n_22943 & ~n_22944;
assign n_22946 =  x_612 & ~n_22945;
assign n_22947 = ~x_612 &  n_22945;
assign n_22948 = ~n_22946 & ~n_22947;
assign n_22949 =  x_611 &  n_21337;
assign n_22950 =  n_21336 &  n_22919;
assign n_22951 = ~n_22949 & ~n_22950;
assign n_22952 =  x_611 & ~n_22951;
assign n_22953 = ~x_611 &  n_22951;
assign n_22954 = ~n_22952 & ~n_22953;
assign n_22955 =  x_610 &  n_21345;
assign n_22956 =  n_21344 &  n_22919;
assign n_22957 = ~n_22955 & ~n_22956;
assign n_22958 =  x_610 & ~n_22957;
assign n_22959 = ~x_610 &  n_22957;
assign n_22960 = ~n_22958 & ~n_22959;
assign n_22961 =  x_609 &  n_21311;
assign n_22962 =  n_21310 &  n_22919;
assign n_22963 = ~n_22961 & ~n_22962;
assign n_22964 =  x_609 & ~n_22963;
assign n_22965 = ~x_609 &  n_22963;
assign n_22966 = ~n_22964 & ~n_22965;
assign n_22967 =  x_608 &  n_21378;
assign n_22968 =  n_21377 &  n_22919;
assign n_22969 = ~n_22967 & ~n_22968;
assign n_22970 =  x_608 & ~n_22969;
assign n_22971 = ~x_608 &  n_22969;
assign n_22972 = ~n_22970 & ~n_22971;
assign n_22973 =  x_607 &  n_21281;
assign n_22974 =  n_21280 &  n_22919;
assign n_22975 = ~n_22973 & ~n_22974;
assign n_22976 =  x_607 & ~n_22975;
assign n_22977 = ~x_607 &  n_22975;
assign n_22978 = ~n_22976 & ~n_22977;
assign n_22979 =  x_606 &  n_21303;
assign n_22980 =  n_21302 &  n_22919;
assign n_22981 = ~n_22979 & ~n_22980;
assign n_22982 =  x_606 & ~n_22981;
assign n_22983 = ~x_606 &  n_22981;
assign n_22984 = ~n_22982 & ~n_22983;
assign n_22985 =  x_605 &  n_21370;
assign n_22986 =  n_21369 &  n_22919;
assign n_22987 = ~n_22985 & ~n_22986;
assign n_22988 =  x_605 & ~n_22987;
assign n_22989 = ~x_605 &  n_22987;
assign n_22990 = ~n_22988 & ~n_22989;
assign n_22991 =  x_604 &  n_21337;
assign n_22992 =  x_411 & ~n_3266;
assign n_22993 =  n_21336 &  n_22992;
assign n_22994 = ~n_22991 & ~n_22993;
assign n_22995 =  x_604 & ~n_22994;
assign n_22996 = ~x_604 &  n_22994;
assign n_22997 = ~n_22995 & ~n_22996;
assign n_22998 =  x_603 &  n_21293;
assign n_22999 =  n_21292 &  n_22992;
assign n_23000 = ~n_22998 & ~n_22999;
assign n_23001 =  x_603 & ~n_23000;
assign n_23002 = ~x_603 &  n_23000;
assign n_23003 = ~n_23001 & ~n_23002;
assign n_23004 =  x_602 &  n_21345;
assign n_23005 =  n_21344 &  n_22992;
assign n_23006 = ~n_23004 & ~n_23005;
assign n_23007 =  x_602 & ~n_23006;
assign n_23008 = ~x_602 &  n_23006;
assign n_23009 = ~n_23007 & ~n_23008;
assign n_23010 =  x_601 &  n_21370;
assign n_23011 =  n_21369 &  n_22992;
assign n_23012 = ~n_23010 & ~n_23011;
assign n_23013 =  x_601 & ~n_23012;
assign n_23014 = ~x_601 &  n_23012;
assign n_23015 = ~n_23013 & ~n_23014;
assign n_23016 =  x_600 &  n_21303;
assign n_23017 =  n_21302 &  n_22992;
assign n_23018 = ~n_23016 & ~n_23017;
assign n_23019 =  x_600 & ~n_23018;
assign n_23020 = ~x_600 &  n_23018;
assign n_23021 = ~n_23019 & ~n_23020;
assign n_23022 =  x_599 &  n_21319;
assign n_23023 =  n_21318 &  n_22992;
assign n_23024 = ~n_23022 & ~n_23023;
assign n_23025 =  x_599 & ~n_23024;
assign n_23026 = ~x_599 &  n_23024;
assign n_23027 = ~n_23025 & ~n_23026;
assign n_23028 =  x_598 &  n_21311;
assign n_23029 =  n_21310 &  n_22992;
assign n_23030 = ~n_23028 & ~n_23029;
assign n_23031 =  x_598 & ~n_23030;
assign n_23032 = ~x_598 &  n_23030;
assign n_23033 = ~n_23031 & ~n_23032;
assign n_23034 =  x_597 &  n_21353;
assign n_23035 =  n_21352 &  n_22992;
assign n_23036 = ~n_23034 & ~n_23035;
assign n_23037 =  x_597 & ~n_23036;
assign n_23038 = ~x_597 &  n_23036;
assign n_23039 = ~n_23037 & ~n_23038;
assign n_23040 =  x_596 &  n_21328;
assign n_23041 =  n_21327 &  n_22992;
assign n_23042 = ~n_23040 & ~n_23041;
assign n_23043 =  x_596 & ~n_23042;
assign n_23044 = ~x_596 &  n_23042;
assign n_23045 = ~n_23043 & ~n_23044;
assign n_23046 =  x_595 &  n_21378;
assign n_23047 =  n_21377 &  n_22992;
assign n_23048 = ~n_23046 & ~n_23047;
assign n_23049 =  x_595 & ~n_23048;
assign n_23050 = ~x_595 &  n_23048;
assign n_23051 = ~n_23049 & ~n_23050;
assign n_23052 =  x_594 &  n_21281;
assign n_23053 =  n_21280 &  n_22992;
assign n_23054 = ~n_23052 & ~n_23053;
assign n_23055 =  x_594 & ~n_23054;
assign n_23056 = ~x_594 &  n_23054;
assign n_23057 = ~n_23055 & ~n_23056;
assign n_23058 =  x_593 &  n_21362;
assign n_23059 =  n_21361 &  n_22992;
assign n_23060 = ~n_23058 & ~n_23059;
assign n_23061 =  x_593 & ~n_23060;
assign n_23062 = ~x_593 &  n_23060;
assign n_23063 = ~n_23061 & ~n_23062;
assign n_23064 =  x_592 &  n_21311;
assign n_23065 =  x_410 & ~n_3266;
assign n_23066 =  n_21310 &  n_23065;
assign n_23067 = ~n_23064 & ~n_23066;
assign n_23068 =  x_592 & ~n_23067;
assign n_23069 = ~x_592 &  n_23067;
assign n_23070 = ~n_23068 & ~n_23069;
assign n_23071 =  x_591 &  n_21378;
assign n_23072 =  n_21377 &  n_23065;
assign n_23073 = ~n_23071 & ~n_23072;
assign n_23074 =  x_591 & ~n_23073;
assign n_23075 = ~x_591 &  n_23073;
assign n_23076 = ~n_23074 & ~n_23075;
assign n_23077 =  x_590 &  n_21345;
assign n_23078 =  n_21344 &  n_23065;
assign n_23079 = ~n_23077 & ~n_23078;
assign n_23080 =  x_590 & ~n_23079;
assign n_23081 = ~x_590 &  n_23079;
assign n_23082 = ~n_23080 & ~n_23081;
assign n_23083 =  x_589 &  n_21337;
assign n_23084 =  n_21336 &  n_23065;
assign n_23085 = ~n_23083 & ~n_23084;
assign n_23086 =  x_589 & ~n_23085;
assign n_23087 = ~x_589 &  n_23085;
assign n_23088 = ~n_23086 & ~n_23087;
assign n_23089 =  x_588 &  n_21353;
assign n_23090 =  n_21352 &  n_23065;
assign n_23091 = ~n_23089 & ~n_23090;
assign n_23092 =  x_588 & ~n_23091;
assign n_23093 = ~x_588 &  n_23091;
assign n_23094 = ~n_23092 & ~n_23093;
assign n_23095 =  x_587 &  n_21281;
assign n_23096 =  n_21280 &  n_23065;
assign n_23097 = ~n_23095 & ~n_23096;
assign n_23098 =  x_587 & ~n_23097;
assign n_23099 = ~x_587 &  n_23097;
assign n_23100 = ~n_23098 & ~n_23099;
assign n_23101 =  x_586 &  n_21293;
assign n_23102 =  n_21292 &  n_23065;
assign n_23103 = ~n_23101 & ~n_23102;
assign n_23104 =  x_586 & ~n_23103;
assign n_23105 = ~x_586 &  n_23103;
assign n_23106 = ~n_23104 & ~n_23105;
assign n_23107 =  x_585 &  n_21328;
assign n_23108 =  n_21327 &  n_23065;
assign n_23109 = ~n_23107 & ~n_23108;
assign n_23110 =  x_585 & ~n_23109;
assign n_23111 = ~x_585 &  n_23109;
assign n_23112 = ~n_23110 & ~n_23111;
assign n_23113 =  x_584 &  n_21303;
assign n_23114 =  n_21302 &  n_23065;
assign n_23115 = ~n_23113 & ~n_23114;
assign n_23116 =  x_584 & ~n_23115;
assign n_23117 = ~x_584 &  n_23115;
assign n_23118 = ~n_23116 & ~n_23117;
assign n_23119 =  x_583 &  n_21370;
assign n_23120 =  n_21369 &  n_23065;
assign n_23121 = ~n_23119 & ~n_23120;
assign n_23122 =  x_583 & ~n_23121;
assign n_23123 = ~x_583 &  n_23121;
assign n_23124 = ~n_23122 & ~n_23123;
assign n_23125 =  x_582 &  n_21362;
assign n_23126 =  n_21361 &  n_23065;
assign n_23127 = ~n_23125 & ~n_23126;
assign n_23128 =  x_582 & ~n_23127;
assign n_23129 = ~x_582 &  n_23127;
assign n_23130 = ~n_23128 & ~n_23129;
assign n_23131 =  x_581 &  n_21319;
assign n_23132 =  n_21318 &  n_23065;
assign n_23133 = ~n_23131 & ~n_23132;
assign n_23134 =  x_581 & ~n_23133;
assign n_23135 = ~x_581 &  n_23133;
assign n_23136 = ~n_23134 & ~n_23135;
assign n_23137 =  x_580 &  n_21303;
assign n_23138 =  x_409 & ~n_3266;
assign n_23139 =  n_21302 &  n_23138;
assign n_23140 = ~n_23137 & ~n_23139;
assign n_23141 =  x_580 & ~n_23140;
assign n_23142 = ~x_580 &  n_23140;
assign n_23143 = ~n_23141 & ~n_23142;
assign n_23144 =  x_579 &  n_21345;
assign n_23145 =  n_21344 &  n_23138;
assign n_23146 = ~n_23144 & ~n_23145;
assign n_23147 =  x_579 & ~n_23146;
assign n_23148 = ~x_579 &  n_23146;
assign n_23149 = ~n_23147 & ~n_23148;
assign n_23150 =  x_578 &  n_21370;
assign n_23151 =  n_21369 &  n_23138;
assign n_23152 = ~n_23150 & ~n_23151;
assign n_23153 =  x_578 & ~n_23152;
assign n_23154 = ~x_578 &  n_23152;
assign n_23155 = ~n_23153 & ~n_23154;
assign n_23156 =  x_577 &  n_21353;
assign n_23157 =  n_21352 &  n_23138;
assign n_23158 = ~n_23156 & ~n_23157;
assign n_23159 =  x_577 & ~n_23158;
assign n_23160 = ~x_577 &  n_23158;
assign n_23161 = ~n_23159 & ~n_23160;
assign n_23162 =  x_576 &  n_21311;
assign n_23163 =  n_21310 &  n_23138;
assign n_23164 = ~n_23162 & ~n_23163;
assign n_23165 =  x_576 & ~n_23164;
assign n_23166 = ~x_576 &  n_23164;
assign n_23167 = ~n_23165 & ~n_23166;
assign n_23168 =  x_575 &  n_21328;
assign n_23169 =  n_21327 &  n_23138;
assign n_23170 = ~n_23168 & ~n_23169;
assign n_23171 =  x_575 & ~n_23170;
assign n_23172 = ~x_575 &  n_23170;
assign n_23173 = ~n_23171 & ~n_23172;
assign n_23174 =  x_574 &  n_21378;
assign n_23175 =  n_21377 &  n_23138;
assign n_23176 = ~n_23174 & ~n_23175;
assign n_23177 =  x_574 & ~n_23176;
assign n_23178 = ~x_574 &  n_23176;
assign n_23179 = ~n_23177 & ~n_23178;
assign n_23180 =  x_573 &  n_21293;
assign n_23181 =  n_21292 &  n_23138;
assign n_23182 = ~n_23180 & ~n_23181;
assign n_23183 =  x_573 & ~n_23182;
assign n_23184 = ~x_573 &  n_23182;
assign n_23185 = ~n_23183 & ~n_23184;
assign n_23186 =  x_572 &  n_21319;
assign n_23187 =  n_21318 &  n_23138;
assign n_23188 = ~n_23186 & ~n_23187;
assign n_23189 =  x_572 & ~n_23188;
assign n_23190 = ~x_572 &  n_23188;
assign n_23191 = ~n_23189 & ~n_23190;
assign n_23192 =  x_571 &  n_21362;
assign n_23193 =  n_21361 &  n_23138;
assign n_23194 = ~n_23192 & ~n_23193;
assign n_23195 =  x_571 & ~n_23194;
assign n_23196 = ~x_571 &  n_23194;
assign n_23197 = ~n_23195 & ~n_23196;
assign n_23198 =  x_570 &  n_21281;
assign n_23199 =  n_21280 &  n_23138;
assign n_23200 = ~n_23198 & ~n_23199;
assign n_23201 =  x_570 & ~n_23200;
assign n_23202 = ~x_570 &  n_23200;
assign n_23203 = ~n_23201 & ~n_23202;
assign n_23204 =  x_569 &  n_21337;
assign n_23205 =  n_21336 &  n_23138;
assign n_23206 = ~n_23204 & ~n_23205;
assign n_23207 =  x_569 & ~n_23206;
assign n_23208 = ~x_569 &  n_23206;
assign n_23209 = ~n_23207 & ~n_23208;
assign n_23210 =  x_568 &  n_21353;
assign n_23211 =  x_408 & ~n_3266;
assign n_23212 =  n_21352 &  n_23211;
assign n_23213 = ~n_23210 & ~n_23212;
assign n_23214 =  x_568 & ~n_23213;
assign n_23215 = ~x_568 &  n_23213;
assign n_23216 = ~n_23214 & ~n_23215;
assign n_23217 =  x_567 &  n_21319;
assign n_23218 =  n_21318 &  n_23211;
assign n_23219 = ~n_23217 & ~n_23218;
assign n_23220 =  x_567 & ~n_23219;
assign n_23221 = ~x_567 &  n_23219;
assign n_23222 = ~n_23220 & ~n_23221;
assign n_23223 =  x_566 &  n_21345;
assign n_23224 =  n_21344 &  n_23211;
assign n_23225 = ~n_23223 & ~n_23224;
assign n_23226 =  x_566 & ~n_23225;
assign n_23227 = ~x_566 &  n_23225;
assign n_23228 = ~n_23226 & ~n_23227;
assign n_23229 =  x_565 &  n_21328;
assign n_23230 =  n_21327 &  n_23211;
assign n_23231 = ~n_23229 & ~n_23230;
assign n_23232 =  x_565 & ~n_23231;
assign n_23233 = ~x_565 &  n_23231;
assign n_23234 = ~n_23232 & ~n_23233;
assign n_23235 =  x_564 &  n_21281;
assign n_23236 =  n_21280 &  n_23211;
assign n_23237 = ~n_23235 & ~n_23236;
assign n_23238 =  x_564 & ~n_23237;
assign n_23239 = ~x_564 &  n_23237;
assign n_23240 = ~n_23238 & ~n_23239;
assign n_23241 =  x_563 &  n_21293;
assign n_23242 =  n_21292 &  n_23211;
assign n_23243 = ~n_23241 & ~n_23242;
assign n_23244 =  x_563 & ~n_23243;
assign n_23245 = ~x_563 &  n_23243;
assign n_23246 = ~n_23244 & ~n_23245;
assign n_23247 =  x_562 &  n_21362;
assign n_23248 =  n_21361 &  n_23211;
assign n_23249 = ~n_23247 & ~n_23248;
assign n_23250 =  x_562 & ~n_23249;
assign n_23251 = ~x_562 &  n_23249;
assign n_23252 = ~n_23250 & ~n_23251;
assign n_23253 =  x_561 &  n_21378;
assign n_23254 =  n_21377 &  n_23211;
assign n_23255 = ~n_23253 & ~n_23254;
assign n_23256 =  x_561 & ~n_23255;
assign n_23257 = ~x_561 &  n_23255;
assign n_23258 = ~n_23256 & ~n_23257;
assign n_23259 =  x_560 &  n_21311;
assign n_23260 =  n_21310 &  n_23211;
assign n_23261 = ~n_23259 & ~n_23260;
assign n_23262 =  x_560 & ~n_23261;
assign n_23263 = ~x_560 &  n_23261;
assign n_23264 = ~n_23262 & ~n_23263;
assign n_23265 =  x_559 &  n_21303;
assign n_23266 =  n_21302 &  n_23211;
assign n_23267 = ~n_23265 & ~n_23266;
assign n_23268 =  x_559 & ~n_23267;
assign n_23269 = ~x_559 &  n_23267;
assign n_23270 = ~n_23268 & ~n_23269;
assign n_23271 =  x_558 &  n_21337;
assign n_23272 =  n_21336 &  n_23211;
assign n_23273 = ~n_23271 & ~n_23272;
assign n_23274 =  x_558 & ~n_23273;
assign n_23275 = ~x_558 &  n_23273;
assign n_23276 = ~n_23274 & ~n_23275;
assign n_23277 =  x_557 &  n_21370;
assign n_23278 =  n_21369 &  n_23211;
assign n_23279 = ~n_23277 & ~n_23278;
assign n_23280 =  x_557 & ~n_23279;
assign n_23281 = ~x_557 &  n_23279;
assign n_23282 = ~n_23280 & ~n_23281;
assign n_23283 =  x_556 &  n_21293;
assign n_23284 =  x_407 & ~n_3266;
assign n_23285 =  n_21292 &  n_23284;
assign n_23286 = ~n_23283 & ~n_23285;
assign n_23287 =  x_556 & ~n_23286;
assign n_23288 = ~x_556 &  n_23286;
assign n_23289 = ~n_23287 & ~n_23288;
assign n_23290 =  x_555 &  n_21353;
assign n_23291 =  n_21352 &  n_23284;
assign n_23292 = ~n_23290 & ~n_23291;
assign n_23293 =  x_555 & ~n_23292;
assign n_23294 = ~x_555 &  n_23292;
assign n_23295 = ~n_23293 & ~n_23294;
assign n_23296 =  x_554 &  n_21319;
assign n_23297 =  n_21318 &  n_23284;
assign n_23298 = ~n_23296 & ~n_23297;
assign n_23299 =  x_554 & ~n_23298;
assign n_23300 = ~x_554 &  n_23298;
assign n_23301 = ~n_23299 & ~n_23300;
assign n_23302 =  x_553 &  n_21345;
assign n_23303 =  n_21344 &  n_23284;
assign n_23304 = ~n_23302 & ~n_23303;
assign n_23305 =  x_553 & ~n_23304;
assign n_23306 = ~x_553 &  n_23304;
assign n_23307 = ~n_23305 & ~n_23306;
assign n_23308 =  x_552 &  n_21328;
assign n_23309 =  n_21327 &  n_23284;
assign n_23310 = ~n_23308 & ~n_23309;
assign n_23311 =  x_552 & ~n_23310;
assign n_23312 = ~x_552 &  n_23310;
assign n_23313 = ~n_23311 & ~n_23312;
assign n_23314 =  x_551 &  n_21281;
assign n_23315 =  n_21280 &  n_23284;
assign n_23316 = ~n_23314 & ~n_23315;
assign n_23317 =  x_551 & ~n_23316;
assign n_23318 = ~x_551 &  n_23316;
assign n_23319 = ~n_23317 & ~n_23318;
assign n_23320 =  x_550 &  n_21362;
assign n_23321 =  n_21361 &  n_23284;
assign n_23322 = ~n_23320 & ~n_23321;
assign n_23323 =  x_550 & ~n_23322;
assign n_23324 = ~x_550 &  n_23322;
assign n_23325 = ~n_23323 & ~n_23324;
assign n_23326 =  x_549 &  n_21370;
assign n_23327 =  n_21369 &  n_23284;
assign n_23328 = ~n_23326 & ~n_23327;
assign n_23329 =  x_549 & ~n_23328;
assign n_23330 = ~x_549 &  n_23328;
assign n_23331 = ~n_23329 & ~n_23330;
assign n_23332 =  x_548 &  n_21311;
assign n_23333 =  n_21310 &  n_23284;
assign n_23334 = ~n_23332 & ~n_23333;
assign n_23335 =  x_548 & ~n_23334;
assign n_23336 = ~x_548 &  n_23334;
assign n_23337 = ~n_23335 & ~n_23336;
assign n_23338 =  x_547 &  n_21303;
assign n_23339 =  n_21302 &  n_23284;
assign n_23340 = ~n_23338 & ~n_23339;
assign n_23341 =  x_547 & ~n_23340;
assign n_23342 = ~x_547 &  n_23340;
assign n_23343 = ~n_23341 & ~n_23342;
assign n_23344 =  x_546 &  n_21337;
assign n_23345 =  n_21336 &  n_23284;
assign n_23346 = ~n_23344 & ~n_23345;
assign n_23347 =  x_546 & ~n_23346;
assign n_23348 = ~x_546 &  n_23346;
assign n_23349 = ~n_23347 & ~n_23348;
assign n_23350 =  x_545 &  n_21378;
assign n_23351 =  n_21377 &  n_23284;
assign n_23352 = ~n_23350 & ~n_23351;
assign n_23353 =  x_545 & ~n_23352;
assign n_23354 = ~x_545 &  n_23352;
assign n_23355 = ~n_23353 & ~n_23354;
assign n_23356 =  x_544 &  n_21328;
assign n_23357 =  x_406 & ~n_3266;
assign n_23358 =  n_21327 &  n_23357;
assign n_23359 = ~n_23356 & ~n_23358;
assign n_23360 =  x_544 & ~n_23359;
assign n_23361 = ~x_544 &  n_23359;
assign n_23362 = ~n_23360 & ~n_23361;
assign n_23363 =  x_543 &  n_21303;
assign n_23364 =  n_21302 &  n_23357;
assign n_23365 = ~n_23363 & ~n_23364;
assign n_23366 =  x_543 & ~n_23365;
assign n_23367 = ~x_543 &  n_23365;
assign n_23368 = ~n_23366 & ~n_23367;
assign n_23369 =  x_542 &  n_21311;
assign n_23370 =  n_21310 &  n_23357;
assign n_23371 = ~n_23369 & ~n_23370;
assign n_23372 =  x_542 & ~n_23371;
assign n_23373 = ~x_542 &  n_23371;
assign n_23374 = ~n_23372 & ~n_23373;
assign n_23375 =  x_541 &  n_21345;
assign n_23376 =  n_21344 &  n_23357;
assign n_23377 = ~n_23375 & ~n_23376;
assign n_23378 =  x_541 & ~n_23377;
assign n_23379 = ~x_541 &  n_23377;
assign n_23380 = ~n_23378 & ~n_23379;
assign n_23381 =  x_540 &  n_21281;
assign n_23382 =  n_21280 &  n_23357;
assign n_23383 = ~n_23381 & ~n_23382;
assign n_23384 =  x_540 & ~n_23383;
assign n_23385 = ~x_540 &  n_23383;
assign n_23386 = ~n_23384 & ~n_23385;
assign n_23387 =  x_539 &  n_21293;
assign n_23388 =  n_21292 &  n_23357;
assign n_23389 = ~n_23387 & ~n_23388;
assign n_23390 =  x_539 & ~n_23389;
assign n_23391 = ~x_539 &  n_23389;
assign n_23392 = ~n_23390 & ~n_23391;
assign n_23393 =  x_538 &  n_21370;
assign n_23394 =  n_21369 &  n_23357;
assign n_23395 = ~n_23393 & ~n_23394;
assign n_23396 =  x_538 & ~n_23395;
assign n_23397 = ~x_538 &  n_23395;
assign n_23398 = ~n_23396 & ~n_23397;
assign n_23399 =  x_537 &  n_21362;
assign n_23400 =  n_21361 &  n_23357;
assign n_23401 = ~n_23399 & ~n_23400;
assign n_23402 =  x_537 & ~n_23401;
assign n_23403 = ~x_537 &  n_23401;
assign n_23404 = ~n_23402 & ~n_23403;
assign n_23405 =  x_536 &  n_21337;
assign n_23406 =  n_21336 &  n_23357;
assign n_23407 = ~n_23405 & ~n_23406;
assign n_23408 =  x_536 & ~n_23407;
assign n_23409 = ~x_536 &  n_23407;
assign n_23410 = ~n_23408 & ~n_23409;
assign n_23411 =  x_535 &  n_21319;
assign n_23412 =  n_21318 &  n_23357;
assign n_23413 = ~n_23411 & ~n_23412;
assign n_23414 =  x_535 & ~n_23413;
assign n_23415 = ~x_535 &  n_23413;
assign n_23416 = ~n_23414 & ~n_23415;
assign n_23417 =  x_534 &  n_21353;
assign n_23418 =  n_21352 &  n_23357;
assign n_23419 = ~n_23417 & ~n_23418;
assign n_23420 =  x_534 & ~n_23419;
assign n_23421 = ~x_534 &  n_23419;
assign n_23422 = ~n_23420 & ~n_23421;
assign n_23423 =  x_533 &  n_21378;
assign n_23424 =  n_21377 &  n_23357;
assign n_23425 = ~n_23423 & ~n_23424;
assign n_23426 =  x_533 & ~n_23425;
assign n_23427 = ~x_533 &  n_23425;
assign n_23428 = ~n_23426 & ~n_23427;
assign n_23429 =  x_532 &  n_21370;
assign n_23430 =  x_405 & ~n_3266;
assign n_23431 =  n_21369 &  n_23430;
assign n_23432 = ~n_23429 & ~n_23431;
assign n_23433 =  x_532 & ~n_23432;
assign n_23434 = ~x_532 &  n_23432;
assign n_23435 = ~n_23433 & ~n_23434;
assign n_23436 =  x_531 &  n_21378;
assign n_23437 =  n_21377 &  n_23430;
assign n_23438 = ~n_23436 & ~n_23437;
assign n_23439 =  x_531 & ~n_23438;
assign n_23440 = ~x_531 &  n_23438;
assign n_23441 = ~n_23439 & ~n_23440;
assign n_23442 =  x_530 &  n_21319;
assign n_23443 =  n_21318 &  n_23430;
assign n_23444 = ~n_23442 & ~n_23443;
assign n_23445 =  x_530 & ~n_23444;
assign n_23446 = ~x_530 &  n_23444;
assign n_23447 = ~n_23445 & ~n_23446;
assign n_23448 =  x_529 &  n_21353;
assign n_23449 =  n_21352 &  n_23430;
assign n_23450 = ~n_23448 & ~n_23449;
assign n_23451 =  x_529 & ~n_23450;
assign n_23452 = ~x_529 &  n_23450;
assign n_23453 = ~n_23451 & ~n_23452;
assign n_23454 =  x_528 &  n_21293;
assign n_23455 =  n_21292 &  n_23430;
assign n_23456 = ~n_23454 & ~n_23455;
assign n_23457 =  x_528 & ~n_23456;
assign n_23458 = ~x_528 &  n_23456;
assign n_23459 = ~n_23457 & ~n_23458;
assign n_23460 =  x_527 &  n_21328;
assign n_23461 =  n_21327 &  n_23430;
assign n_23462 = ~n_23460 & ~n_23461;
assign n_23463 =  x_527 & ~n_23462;
assign n_23464 = ~x_527 &  n_23462;
assign n_23465 = ~n_23463 & ~n_23464;
assign n_23466 =  x_526 &  n_21311;
assign n_23467 =  n_21310 &  n_23430;
assign n_23468 = ~n_23466 & ~n_23467;
assign n_23469 =  x_526 & ~n_23468;
assign n_23470 = ~x_526 &  n_23468;
assign n_23471 = ~n_23469 & ~n_23470;
assign n_23472 =  x_525 &  n_21337;
assign n_23473 =  n_21336 &  n_23430;
assign n_23474 = ~n_23472 & ~n_23473;
assign n_23475 =  x_525 & ~n_23474;
assign n_23476 = ~x_525 &  n_23474;
assign n_23477 = ~n_23475 & ~n_23476;
assign n_23478 =  x_524 &  n_21345;
assign n_23479 =  n_21344 &  n_23430;
assign n_23480 = ~n_23478 & ~n_23479;
assign n_23481 =  x_524 & ~n_23480;
assign n_23482 = ~x_524 &  n_23480;
assign n_23483 = ~n_23481 & ~n_23482;
assign n_23484 =  x_523 &  n_21303;
assign n_23485 =  n_21302 &  n_23430;
assign n_23486 = ~n_23484 & ~n_23485;
assign n_23487 =  x_523 & ~n_23486;
assign n_23488 = ~x_523 &  n_23486;
assign n_23489 = ~n_23487 & ~n_23488;
assign n_23490 =  x_522 &  n_21362;
assign n_23491 =  n_21361 &  n_23430;
assign n_23492 = ~n_23490 & ~n_23491;
assign n_23493 =  x_522 & ~n_23492;
assign n_23494 = ~x_522 &  n_23492;
assign n_23495 = ~n_23493 & ~n_23494;
assign n_23496 =  x_521 &  n_21281;
assign n_23497 =  n_21280 &  n_23430;
assign n_23498 = ~n_23496 & ~n_23497;
assign n_23499 =  x_521 & ~n_23498;
assign n_23500 = ~x_521 &  n_23498;
assign n_23501 = ~n_23499 & ~n_23500;
assign n_23502 =  x_520 &  n_21281;
assign n_23503 =  x_404 & ~n_3266;
assign n_23504 =  n_21280 &  n_23503;
assign n_23505 = ~n_23502 & ~n_23504;
assign n_23506 =  x_520 & ~n_23505;
assign n_23507 = ~x_520 &  n_23505;
assign n_23508 = ~n_23506 & ~n_23507;
assign n_23509 =  x_519 &  n_21353;
assign n_23510 =  n_21352 &  n_23503;
assign n_23511 = ~n_23509 & ~n_23510;
assign n_23512 =  x_519 & ~n_23511;
assign n_23513 = ~x_519 &  n_23511;
assign n_23514 = ~n_23512 & ~n_23513;
assign n_23515 =  x_518 &  n_21311;
assign n_23516 =  n_21310 &  n_23503;
assign n_23517 = ~n_23515 & ~n_23516;
assign n_23518 =  x_518 & ~n_23517;
assign n_23519 = ~x_518 &  n_23517;
assign n_23520 = ~n_23518 & ~n_23519;
assign n_23521 =  x_517 &  n_21328;
assign n_23522 =  n_21327 &  n_23503;
assign n_23523 = ~n_23521 & ~n_23522;
assign n_23524 =  x_517 & ~n_23523;
assign n_23525 = ~x_517 &  n_23523;
assign n_23526 = ~n_23524 & ~n_23525;
assign n_23527 =  x_516 &  n_21370;
assign n_23528 =  n_21369 &  n_23503;
assign n_23529 = ~n_23527 & ~n_23528;
assign n_23530 =  x_516 & ~n_23529;
assign n_23531 = ~x_516 &  n_23529;
assign n_23532 = ~n_23530 & ~n_23531;
assign n_23533 =  x_515 &  n_21319;
assign n_23534 =  n_21318 &  n_23503;
assign n_23535 = ~n_23533 & ~n_23534;
assign n_23536 =  x_515 & ~n_23535;
assign n_23537 = ~x_515 &  n_23535;
assign n_23538 = ~n_23536 & ~n_23537;
assign n_23539 =  x_514 &  n_21293;
assign n_23540 =  n_21292 &  n_23503;
assign n_23541 = ~n_23539 & ~n_23540;
assign n_23542 =  x_514 & ~n_23541;
assign n_23543 = ~x_514 &  n_23541;
assign n_23544 = ~n_23542 & ~n_23543;
assign n_23545 =  x_513 &  n_21303;
assign n_23546 =  n_21302 &  n_23503;
assign n_23547 = ~n_23545 & ~n_23546;
assign n_23548 =  x_513 & ~n_23547;
assign n_23549 = ~x_513 &  n_23547;
assign n_23550 = ~n_23548 & ~n_23549;
assign n_23551 =  x_512 &  n_21345;
assign n_23552 =  n_21344 &  n_23503;
assign n_23553 = ~n_23551 & ~n_23552;
assign n_23554 =  x_512 & ~n_23553;
assign n_23555 = ~x_512 &  n_23553;
assign n_23556 = ~n_23554 & ~n_23555;
assign n_23557 =  x_511 &  n_21378;
assign n_23558 =  n_21377 &  n_23503;
assign n_23559 = ~n_23557 & ~n_23558;
assign n_23560 =  x_511 & ~n_23559;
assign n_23561 = ~x_511 &  n_23559;
assign n_23562 = ~n_23560 & ~n_23561;
assign n_23563 =  x_510 &  n_21362;
assign n_23564 =  n_21361 &  n_23503;
assign n_23565 = ~n_23563 & ~n_23564;
assign n_23566 =  x_510 & ~n_23565;
assign n_23567 = ~x_510 &  n_23565;
assign n_23568 = ~n_23566 & ~n_23567;
assign n_23569 =  x_509 &  n_21337;
assign n_23570 =  n_21336 &  n_23503;
assign n_23571 = ~n_23569 & ~n_23570;
assign n_23572 =  x_509 & ~n_23571;
assign n_23573 = ~x_509 &  n_23571;
assign n_23574 = ~n_23572 & ~n_23573;
assign n_23575 =  x_508 &  n_21281;
assign n_23576 =  x_403 & ~n_3266;
assign n_23577 =  n_21280 &  n_23576;
assign n_23578 = ~n_23575 & ~n_23577;
assign n_23579 =  x_508 & ~n_23578;
assign n_23580 = ~x_508 &  n_23578;
assign n_23581 = ~n_23579 & ~n_23580;
assign n_23582 =  x_507 &  n_21311;
assign n_23583 =  n_21310 &  n_23576;
assign n_23584 = ~n_23582 & ~n_23583;
assign n_23585 =  x_507 & ~n_23584;
assign n_23586 = ~x_507 &  n_23584;
assign n_23587 = ~n_23585 & ~n_23586;
assign n_23588 =  x_506 &  n_21303;
assign n_23589 =  n_21302 &  n_23576;
assign n_23590 = ~n_23588 & ~n_23589;
assign n_23591 =  x_506 & ~n_23590;
assign n_23592 = ~x_506 &  n_23590;
assign n_23593 = ~n_23591 & ~n_23592;
assign n_23594 =  x_505 &  n_21370;
assign n_23595 =  n_21369 &  n_23576;
assign n_23596 = ~n_23594 & ~n_23595;
assign n_23597 =  x_505 & ~n_23596;
assign n_23598 = ~x_505 &  n_23596;
assign n_23599 = ~n_23597 & ~n_23598;
assign n_23600 =  x_504 &  n_21345;
assign n_23601 =  n_21344 &  n_23576;
assign n_23602 = ~n_23600 & ~n_23601;
assign n_23603 =  x_504 & ~n_23602;
assign n_23604 = ~x_504 &  n_23602;
assign n_23605 = ~n_23603 & ~n_23604;
assign n_23606 =  x_503 &  n_21353;
assign n_23607 =  n_21352 &  n_23576;
assign n_23608 = ~n_23606 & ~n_23607;
assign n_23609 =  x_503 & ~n_23608;
assign n_23610 = ~x_503 &  n_23608;
assign n_23611 = ~n_23609 & ~n_23610;
assign n_23612 =  x_502 &  n_21378;
assign n_23613 =  n_21377 &  n_23576;
assign n_23614 = ~n_23612 & ~n_23613;
assign n_23615 =  x_502 & ~n_23614;
assign n_23616 = ~x_502 &  n_23614;
assign n_23617 = ~n_23615 & ~n_23616;
assign n_23618 =  x_501 &  n_21293;
assign n_23619 =  n_21292 &  n_23576;
assign n_23620 = ~n_23618 & ~n_23619;
assign n_23621 =  x_501 & ~n_23620;
assign n_23622 = ~x_501 &  n_23620;
assign n_23623 = ~n_23621 & ~n_23622;
assign n_23624 =  x_500 &  n_21319;
assign n_23625 =  n_21318 &  n_23576;
assign n_23626 = ~n_23624 & ~n_23625;
assign n_23627 =  x_500 & ~n_23626;
assign n_23628 = ~x_500 &  n_23626;
assign n_23629 = ~n_23627 & ~n_23628;
assign n_23630 =  x_499 &  n_21328;
assign n_23631 =  n_21327 &  n_23576;
assign n_23632 = ~n_23630 & ~n_23631;
assign n_23633 =  x_499 & ~n_23632;
assign n_23634 = ~x_499 &  n_23632;
assign n_23635 = ~n_23633 & ~n_23634;
assign n_23636 =  x_498 &  n_21337;
assign n_23637 =  n_21336 &  n_23576;
assign n_23638 = ~n_23636 & ~n_23637;
assign n_23639 =  x_498 & ~n_23638;
assign n_23640 = ~x_498 &  n_23638;
assign n_23641 = ~n_23639 & ~n_23640;
assign n_23642 =  x_497 &  n_21362;
assign n_23643 =  n_21361 &  n_23576;
assign n_23644 = ~n_23642 & ~n_23643;
assign n_23645 =  x_497 & ~n_23644;
assign n_23646 = ~x_497 &  n_23644;
assign n_23647 = ~n_23645 & ~n_23646;
assign n_23648 =  x_496 &  n_21362;
assign n_23649 =  x_402 & ~n_3266;
assign n_23650 =  n_23649 &  n_21361;
assign n_23651 = ~n_23648 & ~n_23650;
assign n_23652 =  x_496 & ~n_23651;
assign n_23653 = ~x_496 &  n_23651;
assign n_23654 = ~n_23652 & ~n_23653;
assign n_23655 =  x_495 &  n_21319;
assign n_23656 =  n_23649 &  n_21318;
assign n_23657 = ~n_23655 & ~n_23656;
assign n_23658 =  x_495 & ~n_23657;
assign n_23659 = ~x_495 &  n_23657;
assign n_23660 = ~n_23658 & ~n_23659;
assign n_23661 =  x_494 &  n_21353;
assign n_23662 =  n_23649 &  n_21352;
assign n_23663 = ~n_23661 & ~n_23662;
assign n_23664 =  x_494 & ~n_23663;
assign n_23665 = ~x_494 &  n_23663;
assign n_23666 = ~n_23664 & ~n_23665;
assign n_23667 =  x_493 &  n_21293;
assign n_23668 =  n_23649 &  n_21292;
assign n_23669 = ~n_23667 & ~n_23668;
assign n_23670 =  x_493 & ~n_23669;
assign n_23671 = ~x_493 &  n_23669;
assign n_23672 = ~n_23670 & ~n_23671;
assign n_23673 =  x_492 &  n_21378;
assign n_23674 =  n_23649 &  n_21377;
assign n_23675 = ~n_23673 & ~n_23674;
assign n_23676 =  x_492 & ~n_23675;
assign n_23677 = ~x_492 &  n_23675;
assign n_23678 = ~n_23676 & ~n_23677;
assign n_23679 =  x_491 &  n_21328;
assign n_23680 =  n_23649 &  n_21327;
assign n_23681 = ~n_23679 & ~n_23680;
assign n_23682 =  x_491 & ~n_23681;
assign n_23683 = ~x_491 &  n_23681;
assign n_23684 = ~n_23682 & ~n_23683;
assign n_23685 =  x_490 &  n_21337;
assign n_23686 =  n_23649 &  n_21336;
assign n_23687 = ~n_23685 & ~n_23686;
assign n_23688 =  x_490 & ~n_23687;
assign n_23689 = ~x_490 &  n_23687;
assign n_23690 = ~n_23688 & ~n_23689;
assign n_23691 =  x_489 &  n_21345;
assign n_23692 =  n_23649 &  n_21344;
assign n_23693 = ~n_23691 & ~n_23692;
assign n_23694 =  x_489 & ~n_23693;
assign n_23695 = ~x_489 &  n_23693;
assign n_23696 = ~n_23694 & ~n_23695;
assign n_23697 =  x_488 &  n_21303;
assign n_23698 =  n_23649 &  n_21302;
assign n_23699 = ~n_23697 & ~n_23698;
assign n_23700 =  x_488 & ~n_23699;
assign n_23701 = ~x_488 &  n_23699;
assign n_23702 = ~n_23700 & ~n_23701;
assign n_23703 =  x_487 &  n_21281;
assign n_23704 =  n_23649 &  n_21280;
assign n_23705 = ~n_23703 & ~n_23704;
assign n_23706 =  x_487 & ~n_23705;
assign n_23707 = ~x_487 &  n_23705;
assign n_23708 = ~n_23706 & ~n_23707;
assign n_23709 =  x_486 &  n_21370;
assign n_23710 =  n_23649 &  n_21369;
assign n_23711 = ~n_23709 & ~n_23710;
assign n_23712 =  x_486 & ~n_23711;
assign n_23713 = ~x_486 &  n_23711;
assign n_23714 = ~n_23712 & ~n_23713;
assign n_23715 =  x_2399 &  n_12630;
assign n_23716 =  x_455 &  n_23715;
assign n_23717 =  n_23716 &  n_12631;
assign n_23718 =  x_457 &  n_23717;
assign n_23719 =  x_458 &  n_23718;
assign n_23720 =  x_459 &  n_23719;
assign n_23721 =  x_460 &  n_23720;
assign n_23722 =  x_461 &  n_23721;
assign n_23723 =  x_462 &  n_23722;
assign n_23724 =  x_463 &  n_23723;
assign n_23725 =  x_464 &  n_23724;
assign n_23726 =  x_465 &  n_23725;
assign n_23727 =  x_466 &  n_23726;
assign n_23728 =  x_467 &  n_23727;
assign n_23729 =  x_468 &  n_23728;
assign n_23730 =  x_469 &  n_23729;
assign n_23731 =  x_470 &  n_23730;
assign n_23732 =  x_471 &  n_23731;
assign n_23733 =  x_472 &  n_23732;
assign n_23734 =  x_473 &  n_23733;
assign n_23735 =  x_474 &  n_23734;
assign n_23736 =  x_475 &  n_23735;
assign n_23737 =  x_476 &  n_23736;
assign n_23738 =  x_477 &  n_23737;
assign n_23739 =  x_478 &  n_23738;
assign n_23740 =  x_479 &  n_23739;
assign n_23741 =  x_480 &  n_23740;
assign n_23742 =  x_481 &  n_23741;
assign n_23743 =  x_482 &  n_23742;
assign n_23744 =  x_483 &  n_23743;
assign n_23745 =  x_484 &  n_23744;
assign n_23746 =  x_485 &  n_23745;
assign n_23747 = ~x_485 & ~n_23745;
assign n_23748 = ~n_1192 & ~n_23747;
assign n_23749 = ~n_23746 &  n_23748;
assign n_23750 =  x_485 &  n_23749;
assign n_23751 = ~x_485 & ~n_23749;
assign n_23752 = ~n_23750 & ~n_23751;
assign n_23753 = ~x_484 & ~n_23744;
assign n_23754 = ~n_1192 & ~n_23745;
assign n_23755 = ~n_23753 &  n_23754;
assign n_23756 =  x_484 &  n_23755;
assign n_23757 = ~x_484 & ~n_23755;
assign n_23758 = ~n_23756 & ~n_23757;
assign n_23759 = ~x_483 & ~n_23743;
assign n_23760 = ~n_1192 & ~n_23744;
assign n_23761 = ~n_23759 &  n_23760;
assign n_23762 =  x_483 &  n_23761;
assign n_23763 = ~x_483 & ~n_23761;
assign n_23764 = ~n_23762 & ~n_23763;
assign n_23765 = ~x_482 & ~n_23742;
assign n_23766 = ~n_1192 & ~n_23743;
assign n_23767 = ~n_23765 &  n_23766;
assign n_23768 =  x_482 &  n_23767;
assign n_23769 = ~x_482 & ~n_23767;
assign n_23770 = ~n_23768 & ~n_23769;
assign n_23771 = ~x_481 & ~n_23741;
assign n_23772 = ~n_1192 & ~n_23742;
assign n_23773 = ~n_23771 &  n_23772;
assign n_23774 =  x_481 &  n_23773;
assign n_23775 = ~x_481 & ~n_23773;
assign n_23776 = ~n_23774 & ~n_23775;
assign n_23777 = ~x_480 & ~n_23740;
assign n_23778 = ~n_1192 & ~n_23741;
assign n_23779 = ~n_23777 &  n_23778;
assign n_23780 =  x_480 &  n_23779;
assign n_23781 = ~x_480 & ~n_23779;
assign n_23782 = ~n_23780 & ~n_23781;
assign n_23783 = ~x_479 & ~n_23739;
assign n_23784 = ~n_1192 & ~n_23740;
assign n_23785 = ~n_23783 &  n_23784;
assign n_23786 =  x_479 &  n_23785;
assign n_23787 = ~x_479 & ~n_23785;
assign n_23788 = ~n_23786 & ~n_23787;
assign n_23789 = ~x_478 & ~n_23738;
assign n_23790 = ~n_1192 & ~n_23739;
assign n_23791 = ~n_23789 &  n_23790;
assign n_23792 =  x_478 &  n_23791;
assign n_23793 = ~x_478 & ~n_23791;
assign n_23794 = ~n_23792 & ~n_23793;
assign n_23795 = ~x_477 & ~n_23737;
assign n_23796 = ~n_1192 & ~n_23738;
assign n_23797 = ~n_23795 &  n_23796;
assign n_23798 =  x_477 &  n_23797;
assign n_23799 = ~x_477 & ~n_23797;
assign n_23800 = ~n_23798 & ~n_23799;
assign n_23801 = ~x_476 & ~n_23736;
assign n_23802 = ~n_1192 & ~n_23737;
assign n_23803 = ~n_23801 &  n_23802;
assign n_23804 =  x_476 &  n_23803;
assign n_23805 = ~x_476 & ~n_23803;
assign n_23806 = ~n_23804 & ~n_23805;
assign n_23807 = ~x_475 & ~n_23735;
assign n_23808 = ~n_1192 & ~n_23736;
assign n_23809 = ~n_23807 &  n_23808;
assign n_23810 =  x_475 &  n_23809;
assign n_23811 = ~x_475 & ~n_23809;
assign n_23812 = ~n_23810 & ~n_23811;
assign n_23813 = ~x_474 & ~n_23734;
assign n_23814 = ~n_1192 & ~n_23735;
assign n_23815 = ~n_23813 &  n_23814;
assign n_23816 =  x_474 &  n_23815;
assign n_23817 = ~x_474 & ~n_23815;
assign n_23818 = ~n_23816 & ~n_23817;
assign n_23819 = ~x_473 & ~n_23733;
assign n_23820 = ~n_1192 & ~n_23734;
assign n_23821 = ~n_23819 &  n_23820;
assign n_23822 =  x_473 &  n_23821;
assign n_23823 = ~x_473 & ~n_23821;
assign n_23824 = ~n_23822 & ~n_23823;
assign n_23825 = ~x_472 & ~n_23732;
assign n_23826 = ~n_1192 & ~n_23733;
assign n_23827 = ~n_23825 &  n_23826;
assign n_23828 =  x_472 &  n_23827;
assign n_23829 = ~x_472 & ~n_23827;
assign n_23830 = ~n_23828 & ~n_23829;
assign n_23831 = ~x_471 & ~n_23731;
assign n_23832 = ~n_1192 & ~n_23732;
assign n_23833 = ~n_23831 &  n_23832;
assign n_23834 =  x_471 &  n_23833;
assign n_23835 = ~x_471 & ~n_23833;
assign n_23836 = ~n_23834 & ~n_23835;
assign n_23837 = ~x_470 & ~n_23730;
assign n_23838 = ~n_1192 & ~n_23731;
assign n_23839 = ~n_23837 &  n_23838;
assign n_23840 =  x_470 &  n_23839;
assign n_23841 = ~x_470 & ~n_23839;
assign n_23842 = ~n_23840 & ~n_23841;
assign n_23843 = ~x_469 & ~n_23729;
assign n_23844 = ~n_1192 & ~n_23730;
assign n_23845 = ~n_23843 &  n_23844;
assign n_23846 =  x_469 &  n_23845;
assign n_23847 = ~x_469 & ~n_23845;
assign n_23848 = ~n_23846 & ~n_23847;
assign n_23849 = ~x_468 & ~n_23728;
assign n_23850 = ~n_1192 & ~n_23729;
assign n_23851 = ~n_23849 &  n_23850;
assign n_23852 =  x_468 &  n_23851;
assign n_23853 = ~x_468 & ~n_23851;
assign n_23854 = ~n_23852 & ~n_23853;
assign n_23855 = ~x_467 & ~n_23727;
assign n_23856 = ~n_1192 & ~n_23728;
assign n_23857 = ~n_23855 &  n_23856;
assign n_23858 =  x_467 &  n_23857;
assign n_23859 = ~x_467 & ~n_23857;
assign n_23860 = ~n_23858 & ~n_23859;
assign n_23861 = ~x_466 & ~n_23726;
assign n_23862 = ~n_1192 & ~n_23727;
assign n_23863 = ~n_23861 &  n_23862;
assign n_23864 =  x_466 &  n_23863;
assign n_23865 = ~x_466 & ~n_23863;
assign n_23866 = ~n_23864 & ~n_23865;
assign n_23867 = ~x_465 & ~n_23725;
assign n_23868 = ~n_1192 & ~n_23726;
assign n_23869 = ~n_23867 &  n_23868;
assign n_23870 =  x_465 &  n_23869;
assign n_23871 = ~x_465 & ~n_23869;
assign n_23872 = ~n_23870 & ~n_23871;
assign n_23873 = ~x_464 & ~n_23724;
assign n_23874 = ~n_1192 & ~n_23725;
assign n_23875 = ~n_23873 &  n_23874;
assign n_23876 =  x_464 &  n_23875;
assign n_23877 = ~x_464 & ~n_23875;
assign n_23878 = ~n_23876 & ~n_23877;
assign n_23879 = ~x_463 & ~n_23723;
assign n_23880 = ~n_1192 & ~n_23724;
assign n_23881 = ~n_23879 &  n_23880;
assign n_23882 =  x_463 &  n_23881;
assign n_23883 = ~x_463 & ~n_23881;
assign n_23884 = ~n_23882 & ~n_23883;
assign n_23885 = ~x_462 & ~n_23722;
assign n_23886 = ~n_1192 & ~n_23723;
assign n_23887 = ~n_23885 &  n_23886;
assign n_23888 =  x_462 &  n_23887;
assign n_23889 = ~x_462 & ~n_23887;
assign n_23890 = ~n_23888 & ~n_23889;
assign n_23891 = ~x_461 & ~n_23721;
assign n_23892 = ~n_1192 & ~n_23722;
assign n_23893 = ~n_23891 &  n_23892;
assign n_23894 =  x_461 &  n_23893;
assign n_23895 = ~x_461 & ~n_23893;
assign n_23896 = ~n_23894 & ~n_23895;
assign n_23897 = ~x_460 & ~n_23720;
assign n_23898 = ~n_1192 & ~n_23721;
assign n_23899 = ~n_23897 &  n_23898;
assign n_23900 =  x_460 &  n_23899;
assign n_23901 = ~x_460 & ~n_23899;
assign n_23902 = ~n_23900 & ~n_23901;
assign n_23903 = ~x_459 & ~n_23719;
assign n_23904 = ~n_1192 & ~n_23720;
assign n_23905 = ~n_23903 &  n_23904;
assign n_23906 =  x_459 &  n_23905;
assign n_23907 = ~x_459 & ~n_23905;
assign n_23908 = ~n_23906 & ~n_23907;
assign n_23909 = ~x_458 & ~n_23718;
assign n_23910 = ~n_1192 & ~n_23719;
assign n_23911 = ~n_23909 &  n_23910;
assign n_23912 =  x_458 &  n_23911;
assign n_23913 = ~x_458 & ~n_23911;
assign n_23914 = ~n_23912 & ~n_23913;
assign n_23915 = ~x_457 & ~n_23717;
assign n_23916 = ~n_1192 & ~n_23718;
assign n_23917 = ~n_23915 &  n_23916;
assign n_23918 =  x_457 &  n_23917;
assign n_23919 = ~x_457 & ~n_23917;
assign n_23920 = ~n_23918 & ~n_23919;
assign n_23921 = ~n_23716 & ~n_12631;
assign n_23922 = ~n_23921 & ~n_23717;
assign n_23923 =  x_456 &  n_23922;
assign n_23924 = ~x_456 & ~n_23922;
assign n_23925 = ~n_23923 & ~n_23924;
assign n_23926 = ~n_23715 & ~n_12679;
assign n_23927 = ~n_23926 & ~n_23716;
assign n_23928 =  x_455 &  n_23927;
assign n_23929 = ~x_455 & ~n_23927;
assign n_23930 = ~n_23928 & ~n_23929;
assign n_23931 = ~x_2399 & ~n_12630;
assign n_23932 = ~n_23715 & ~n_23931;
assign n_23933 =  x_454 &  n_23932;
assign n_23934 = ~x_454 & ~n_23932;
assign n_23935 = ~n_23933 & ~n_23934;
assign n_23936 =  x_453 &  n_21311;
assign n_23937 =  n_21310 &  n_23649;
assign n_23938 = ~n_23936 & ~n_23937;
assign n_23939 =  x_453 & ~n_23938;
assign n_23940 = ~x_453 &  n_23938;
assign n_23941 = ~n_23939 & ~n_23940;
assign n_23942 =  x_452 & ~n_3266;
assign n_23943 = ~x_452 &  n_3266;
assign n_23944 = ~n_23942 & ~n_23943;
assign n_23945 =  x_451 &  n_6111;
assign n_23946 = ~x_451 & ~n_6111;
assign n_23947 = ~n_23945 & ~n_23946;
assign n_23948 = ~x_1078 &  n_5;
assign n_23949 = ~x_1082 &  n_13;
assign n_23950 = ~n_23948 & ~n_23949;
assign n_23951 = ~x_1080 &  n_11;
assign n_23952 = ~x_1076 &  n_8;
assign n_23953 = ~n_23951 & ~n_23952;
assign n_23954 =  n_23950 &  n_23953;
assign n_23955 = ~x_1081 &  n_32;
assign n_23956 = ~x_1083 &  n_26;
assign n_23957 = ~n_23955 & ~n_23956;
assign n_23958 = ~x_1077 &  n_30;
assign n_23959 = ~x_1079 &  n_24;
assign n_23960 = ~n_23958 & ~n_23959;
assign n_23961 =  n_23957 &  n_23960;
assign n_23962 =  n_23954 &  n_23961;
assign n_23963 =  x_450 &  n_23962;
assign n_23964 = ~x_450 & ~n_23962;
assign n_23965 = ~n_23963 & ~n_23964;
assign n_23966 = ~x_1058 &  n_8;
assign n_23967 = ~x_1060 &  n_5;
assign n_23968 = ~n_23966 & ~n_23967;
assign n_23969 = ~x_1062 &  n_11;
assign n_23970 = ~x_1064 &  n_13;
assign n_23971 = ~n_23969 & ~n_23970;
assign n_23972 =  n_23968 &  n_23971;
assign n_23973 = ~x_1065 &  n_26;
assign n_23974 = ~x_1061 &  n_24;
assign n_23975 = ~n_23973 & ~n_23974;
assign n_23976 = ~x_1059 &  n_30;
assign n_23977 = ~x_1063 &  n_32;
assign n_23978 = ~n_23976 & ~n_23977;
assign n_23979 =  n_23975 &  n_23978;
assign n_23980 =  n_23972 &  n_23979;
assign n_23981 =  x_449 &  n_23980;
assign n_23982 = ~x_449 & ~n_23980;
assign n_23983 = ~n_23981 & ~n_23982;
assign n_23984 = ~x_1046 &  n_13;
assign n_23985 = ~x_1044 &  n_11;
assign n_23986 = ~n_23984 & ~n_23985;
assign n_23987 = ~x_1040 &  n_8;
assign n_23988 = ~x_1042 &  n_5;
assign n_23989 = ~n_23987 & ~n_23988;
assign n_23990 =  n_23986 &  n_23989;
assign n_23991 = ~x_1041 &  n_30;
assign n_23992 = ~x_1043 &  n_24;
assign n_23993 = ~n_23991 & ~n_23992;
assign n_23994 = ~x_1047 &  n_26;
assign n_23995 = ~x_1045 &  n_32;
assign n_23996 = ~n_23994 & ~n_23995;
assign n_23997 =  n_23993 &  n_23996;
assign n_23998 =  n_23990 &  n_23997;
assign n_23999 =  x_448 &  n_23998;
assign n_24000 = ~x_448 & ~n_23998;
assign n_24001 = ~n_23999 & ~n_24000;
assign n_24002 = ~x_1026 &  n_11;
assign n_24003 = ~x_1028 &  n_13;
assign n_24004 = ~n_24002 & ~n_24003;
assign n_24005 = ~x_1024 &  n_5;
assign n_24006 = ~x_1022 &  n_8;
assign n_24007 = ~n_24005 & ~n_24006;
assign n_24008 =  n_24004 &  n_24007;
assign n_24009 = ~x_1023 &  n_30;
assign n_24010 = ~x_1027 &  n_32;
assign n_24011 = ~n_24009 & ~n_24010;
assign n_24012 = ~x_1025 &  n_24;
assign n_24013 = ~x_1029 &  n_26;
assign n_24014 = ~n_24012 & ~n_24013;
assign n_24015 =  n_24011 &  n_24014;
assign n_24016 =  n_24008 &  n_24015;
assign n_24017 =  x_447 &  n_24016;
assign n_24018 = ~x_447 & ~n_24016;
assign n_24019 = ~n_24017 & ~n_24018;
assign n_24020 = ~x_1069 &  n_5;
assign n_24021 = ~x_1071 &  n_11;
assign n_24022 = ~n_24020 & ~n_24021;
assign n_24023 = ~x_1073 &  n_13;
assign n_24024 = ~x_1067 &  n_8;
assign n_24025 = ~n_24023 & ~n_24024;
assign n_24026 =  n_24022 &  n_24025;
assign n_24027 = ~x_1068 &  n_30;
assign n_24028 = ~x_1074 &  n_26;
assign n_24029 = ~n_24027 & ~n_24028;
assign n_24030 = ~x_1070 &  n_24;
assign n_24031 = ~x_1072 &  n_32;
assign n_24032 = ~n_24030 & ~n_24031;
assign n_24033 =  n_24029 &  n_24032;
assign n_24034 =  n_24026 &  n_24033;
assign n_24035 =  x_446 &  n_24034;
assign n_24036 = ~x_446 & ~n_24034;
assign n_24037 = ~n_24035 & ~n_24036;
assign n_24038 = ~x_1051 &  n_5;
assign n_24039 = ~x_1055 &  n_13;
assign n_24040 = ~n_24038 & ~n_24039;
assign n_24041 = ~x_1049 &  n_8;
assign n_24042 = ~x_1053 &  n_11;
assign n_24043 = ~n_24041 & ~n_24042;
assign n_24044 =  n_24040 &  n_24043;
assign n_24045 = ~x_1054 &  n_32;
assign n_24046 = ~x_1050 &  n_30;
assign n_24047 = ~n_24045 & ~n_24046;
assign n_24048 = ~x_1052 &  n_24;
assign n_24049 = ~x_1056 &  n_26;
assign n_24050 = ~n_24048 & ~n_24049;
assign n_24051 =  n_24047 &  n_24050;
assign n_24052 =  n_24044 &  n_24051;
assign n_24053 =  x_445 &  n_24052;
assign n_24054 = ~x_445 & ~n_24052;
assign n_24055 = ~n_24053 & ~n_24054;
assign n_24056 = ~x_1035 &  n_11;
assign n_24057 = ~x_1033 &  n_5;
assign n_24058 = ~n_24056 & ~n_24057;
assign n_24059 = ~x_1031 &  n_8;
assign n_24060 = ~x_1037 &  n_13;
assign n_24061 = ~n_24059 & ~n_24060;
assign n_24062 =  n_24058 &  n_24061;
assign n_24063 = ~x_1032 &  n_30;
assign n_24064 = ~x_1036 &  n_32;
assign n_24065 = ~n_24063 & ~n_24064;
assign n_24066 = ~x_1034 &  n_24;
assign n_24067 = ~x_1038 &  n_26;
assign n_24068 = ~n_24066 & ~n_24067;
assign n_24069 =  n_24065 &  n_24068;
assign n_24070 =  n_24062 &  n_24069;
assign n_24071 =  x_444 &  n_24070;
assign n_24072 = ~x_444 & ~n_24070;
assign n_24073 = ~n_24071 & ~n_24072;
assign n_24074 = ~x_1016 &  n_5;
assign n_24075 = ~x_1018 &  n_11;
assign n_24076 = ~n_24074 & ~n_24075;
assign n_24077 = ~x_1014 &  n_8;
assign n_24078 = ~x_1020 &  n_13;
assign n_24079 = ~n_24077 & ~n_24078;
assign n_24080 =  n_24076 &  n_24079;
assign n_24081 = ~x_1019 &  n_32;
assign n_24082 = ~x_1017 &  n_24;
assign n_24083 = ~n_24081 & ~n_24082;
assign n_24084 = ~x_1015 &  n_30;
assign n_24085 = ~x_1021 &  n_26;
assign n_24086 = ~n_24084 & ~n_24085;
assign n_24087 =  n_24083 &  n_24086;
assign n_24088 =  n_24080 &  n_24087;
assign n_24089 =  x_443 &  n_24088;
assign n_24090 = ~x_443 & ~n_24088;
assign n_24091 = ~n_24089 & ~n_24090;
assign n_24092 = ~x_940 &  n_8;
assign n_24093 = ~x_944 &  n_11;
assign n_24094 = ~n_24092 & ~n_24093;
assign n_24095 = ~x_946 &  n_13;
assign n_24096 = ~x_942 &  n_5;
assign n_24097 = ~n_24095 & ~n_24096;
assign n_24098 =  n_24094 &  n_24097;
assign n_24099 = ~x_943 &  n_24;
assign n_24100 = ~x_941 &  n_30;
assign n_24101 = ~n_24099 & ~n_24100;
assign n_24102 = ~x_945 &  n_32;
assign n_24103 = ~x_947 &  n_26;
assign n_24104 = ~n_24102 & ~n_24103;
assign n_24105 =  n_24101 &  n_24104;
assign n_24106 =  n_24098 &  n_24105;
assign n_24107 =  x_442 &  n_24106;
assign n_24108 = ~x_442 & ~n_24106;
assign n_24109 = ~n_24107 & ~n_24108;
assign n_24110 = ~x_934 &  n_5;
assign n_24111 = ~x_938 &  n_13;
assign n_24112 = ~n_24110 & ~n_24111;
assign n_24113 = ~x_932 &  n_8;
assign n_24114 = ~x_936 &  n_11;
assign n_24115 = ~n_24113 & ~n_24114;
assign n_24116 =  n_24112 &  n_24115;
assign n_24117 = ~x_937 &  n_32;
assign n_24118 = ~x_933 &  n_30;
assign n_24119 = ~n_24117 & ~n_24118;
assign n_24120 = ~x_935 &  n_24;
assign n_24121 = ~x_939 &  n_26;
assign n_24122 = ~n_24120 & ~n_24121;
assign n_24123 =  n_24119 &  n_24122;
assign n_24124 =  n_24116 &  n_24123;
assign n_24125 =  x_441 &  n_24124;
assign n_24126 = ~x_441 & ~n_24124;
assign n_24127 = ~n_24125 & ~n_24126;
assign n_24128 = ~x_924 &  n_8;
assign n_24129 = ~x_930 &  n_13;
assign n_24130 = ~n_24128 & ~n_24129;
assign n_24131 = ~x_926 &  n_5;
assign n_24132 = ~x_928 &  n_11;
assign n_24133 = ~n_24131 & ~n_24132;
assign n_24134 =  n_24130 &  n_24133;
assign n_24135 = ~x_925 &  n_30;
assign n_24136 = ~x_931 &  n_26;
assign n_24137 = ~n_24135 & ~n_24136;
assign n_24138 = ~x_929 &  n_32;
assign n_24139 = ~x_927 &  n_24;
assign n_24140 = ~n_24138 & ~n_24139;
assign n_24141 =  n_24137 &  n_24140;
assign n_24142 =  n_24134 &  n_24141;
assign n_24143 =  x_440 &  n_24142;
assign n_24144 = ~x_440 & ~n_24142;
assign n_24145 = ~n_24143 & ~n_24144;
assign n_24146 = ~x_916 &  n_8;
assign n_24147 = ~x_920 &  n_11;
assign n_24148 = ~n_24146 & ~n_24147;
assign n_24149 = ~x_922 &  n_13;
assign n_24150 = ~x_918 &  n_5;
assign n_24151 = ~n_24149 & ~n_24150;
assign n_24152 =  n_24148 &  n_24151;
assign n_24153 = ~x_921 &  n_32;
assign n_24154 = ~x_919 &  n_24;
assign n_24155 = ~n_24153 & ~n_24154;
assign n_24156 = ~x_917 &  n_30;
assign n_24157 = ~x_923 &  n_26;
assign n_24158 = ~n_24156 & ~n_24157;
assign n_24159 =  n_24155 &  n_24158;
assign n_24160 =  n_24152 &  n_24159;
assign n_24161 =  x_439 &  n_24160;
assign n_24162 = ~x_439 & ~n_24160;
assign n_24163 = ~n_24161 & ~n_24162;
assign n_24164 = ~x_910 &  n_5;
assign n_24165 = ~x_914 &  n_13;
assign n_24166 = ~n_24164 & ~n_24165;
assign n_24167 = ~x_912 &  n_11;
assign n_24168 = ~x_908 &  n_8;
assign n_24169 = ~n_24167 & ~n_24168;
assign n_24170 =  n_24166 &  n_24169;
assign n_24171 = ~x_909 &  n_30;
assign n_24172 = ~x_913 &  n_32;
assign n_24173 = ~n_24171 & ~n_24172;
assign n_24174 = ~x_915 &  n_26;
assign n_24175 = ~x_911 &  n_24;
assign n_24176 = ~n_24174 & ~n_24175;
assign n_24177 =  n_24173 &  n_24176;
assign n_24178 =  n_24170 &  n_24177;
assign n_24179 =  x_438 &  n_24178;
assign n_24180 = ~x_438 & ~n_24178;
assign n_24181 = ~n_24179 & ~n_24180;
assign n_24182 = ~x_904 &  n_11;
assign n_24183 = ~x_902 &  n_5;
assign n_24184 = ~n_24182 & ~n_24183;
assign n_24185 = ~x_906 &  n_13;
assign n_24186 = ~x_900 &  n_8;
assign n_24187 = ~n_24185 & ~n_24186;
assign n_24188 =  n_24184 &  n_24187;
assign n_24189 = ~x_905 &  n_32;
assign n_24190 = ~x_907 &  n_26;
assign n_24191 = ~n_24189 & ~n_24190;
assign n_24192 = ~x_903 &  n_24;
assign n_24193 = ~x_901 &  n_30;
assign n_24194 = ~n_24192 & ~n_24193;
assign n_24195 =  n_24191 &  n_24194;
assign n_24196 =  n_24188 &  n_24195;
assign n_24197 =  x_437 &  n_24196;
assign n_24198 = ~x_437 & ~n_24196;
assign n_24199 = ~n_24197 & ~n_24198;
assign n_24200 = ~x_898 &  n_13;
assign n_24201 = ~x_894 &  n_5;
assign n_24202 = ~n_24200 & ~n_24201;
assign n_24203 = ~x_892 &  n_8;
assign n_24204 = ~x_896 &  n_11;
assign n_24205 = ~n_24203 & ~n_24204;
assign n_24206 =  n_24202 &  n_24205;
assign n_24207 = ~x_895 &  n_24;
assign n_24208 = ~x_897 &  n_32;
assign n_24209 = ~n_24207 & ~n_24208;
assign n_24210 = ~x_893 &  n_30;
assign n_24211 = ~x_899 &  n_26;
assign n_24212 = ~n_24210 & ~n_24211;
assign n_24213 =  n_24209 &  n_24212;
assign n_24214 =  n_24206 &  n_24213;
assign n_24215 =  x_436 &  n_24214;
assign n_24216 = ~x_436 & ~n_24214;
assign n_24217 = ~n_24215 & ~n_24216;
assign n_24218 = ~x_886 &  n_5;
assign n_24219 = ~x_890 &  n_13;
assign n_24220 = ~n_24218 & ~n_24219;
assign n_24221 = ~x_888 &  n_11;
assign n_24222 = ~x_884 &  n_8;
assign n_24223 = ~n_24221 & ~n_24222;
assign n_24224 =  n_24220 &  n_24223;
assign n_24225 = ~x_889 &  n_32;
assign n_24226 = ~x_887 &  n_24;
assign n_24227 = ~n_24225 & ~n_24226;
assign n_24228 = ~x_885 &  n_30;
assign n_24229 = ~x_891 &  n_26;
assign n_24230 = ~n_24228 & ~n_24229;
assign n_24231 =  n_24227 &  n_24230;
assign n_24232 =  n_24224 &  n_24231;
assign n_24233 =  x_435 &  n_24232;
assign n_24234 = ~x_435 & ~n_24232;
assign n_24235 = ~n_24233 & ~n_24234;
assign n_24236 = ~x_1464 &  n_13;
assign n_24237 = ~x_1462 &  n_11;
assign n_24238 = ~n_24236 & ~n_24237;
assign n_24239 = ~x_1460 &  n_5;
assign n_24240 = ~x_1458 &  n_8;
assign n_24241 = ~n_24239 & ~n_24240;
assign n_24242 =  n_24238 &  n_24241;
assign n_24243 = ~x_1463 &  n_32;
assign n_24244 = ~x_1465 &  n_26;
assign n_24245 = ~n_24243 & ~n_24244;
assign n_24246 = ~x_1459 &  n_30;
assign n_24247 = ~x_1461 &  n_24;
assign n_24248 = ~n_24246 & ~n_24247;
assign n_24249 =  n_24245 &  n_24248;
assign n_24250 =  n_24242 &  n_24249;
assign n_24251 =  x_434 &  n_24250;
assign n_24252 = ~x_434 & ~n_24250;
assign n_24253 = ~n_24251 & ~n_24252;
assign n_24254 = ~x_1450 &  n_8;
assign n_24255 = ~x_1452 &  n_5;
assign n_24256 = ~n_24254 & ~n_24255;
assign n_24257 = ~x_1456 &  n_13;
assign n_24258 = ~x_1454 &  n_11;
assign n_24259 = ~n_24257 & ~n_24258;
assign n_24260 =  n_24256 &  n_24259;
assign n_24261 = ~x_1457 &  n_26;
assign n_24262 = ~x_1455 &  n_32;
assign n_24263 = ~n_24261 & ~n_24262;
assign n_24264 = ~x_1451 &  n_30;
assign n_24265 = ~x_1453 &  n_24;
assign n_24266 = ~n_24264 & ~n_24265;
assign n_24267 =  n_24263 &  n_24266;
assign n_24268 =  n_24260 &  n_24267;
assign n_24269 =  x_433 &  n_24268;
assign n_24270 = ~x_433 & ~n_24268;
assign n_24271 = ~n_24269 & ~n_24270;
assign n_24272 = ~x_1442 &  n_8;
assign n_24273 = ~x_1444 &  n_5;
assign n_24274 = ~n_24272 & ~n_24273;
assign n_24275 = ~x_1448 &  n_13;
assign n_24276 = ~x_1446 &  n_11;
assign n_24277 = ~n_24275 & ~n_24276;
assign n_24278 =  n_24274 &  n_24277;
assign n_24279 = ~x_1447 &  n_32;
assign n_24280 = ~x_1445 &  n_24;
assign n_24281 = ~n_24279 & ~n_24280;
assign n_24282 = ~x_1449 &  n_26;
assign n_24283 = ~x_1443 &  n_30;
assign n_24284 = ~n_24282 & ~n_24283;
assign n_24285 =  n_24281 &  n_24284;
assign n_24286 =  n_24278 &  n_24285;
assign n_24287 =  x_432 &  n_24286;
assign n_24288 = ~x_432 & ~n_24286;
assign n_24289 = ~n_24287 & ~n_24288;
assign n_24290 = ~x_1436 &  n_5;
assign n_24291 = ~x_1438 &  n_11;
assign n_24292 = ~n_24290 & ~n_24291;
assign n_24293 = ~x_1434 &  n_8;
assign n_24294 = ~x_1440 &  n_13;
assign n_24295 = ~n_24293 & ~n_24294;
assign n_24296 =  n_24292 &  n_24295;
assign n_24297 = ~x_1439 &  n_32;
assign n_24298 = ~x_1437 &  n_24;
assign n_24299 = ~n_24297 & ~n_24298;
assign n_24300 = ~x_1441 &  n_26;
assign n_24301 = ~x_1435 &  n_30;
assign n_24302 = ~n_24300 & ~n_24301;
assign n_24303 =  n_24299 &  n_24302;
assign n_24304 =  n_24296 &  n_24303;
assign n_24305 =  x_431 &  n_24304;
assign n_24306 = ~x_431 & ~n_24304;
assign n_24307 = ~n_24305 & ~n_24306;
assign n_24308 = ~x_1428 &  n_5;
assign n_24309 = ~x_1426 &  n_8;
assign n_24310 = ~n_24308 & ~n_24309;
assign n_24311 = ~x_1432 &  n_13;
assign n_24312 = ~x_1430 &  n_11;
assign n_24313 = ~n_24311 & ~n_24312;
assign n_24314 =  n_24310 &  n_24313;
assign n_24315 = ~x_1427 &  n_30;
assign n_24316 = ~x_1429 &  n_24;
assign n_24317 = ~n_24315 & ~n_24316;
assign n_24318 = ~x_1431 &  n_32;
assign n_24319 = ~x_1433 &  n_26;
assign n_24320 = ~n_24318 & ~n_24319;
assign n_24321 =  n_24317 &  n_24320;
assign n_24322 =  n_24314 &  n_24321;
assign n_24323 =  x_430 &  n_24322;
assign n_24324 = ~x_430 & ~n_24322;
assign n_24325 = ~n_24323 & ~n_24324;
assign n_24326 = ~x_1420 &  n_5;
assign n_24327 = ~x_1422 &  n_11;
assign n_24328 = ~n_24326 & ~n_24327;
assign n_24329 = ~x_1418 &  n_8;
assign n_24330 = ~x_1424 &  n_13;
assign n_24331 = ~n_24329 & ~n_24330;
assign n_24332 =  n_24328 &  n_24331;
assign n_24333 = ~x_1419 &  n_30;
assign n_24334 = ~x_1425 &  n_26;
assign n_24335 = ~n_24333 & ~n_24334;
assign n_24336 = ~x_1423 &  n_32;
assign n_24337 = ~x_1421 &  n_24;
assign n_24338 = ~n_24336 & ~n_24337;
assign n_24339 =  n_24335 &  n_24338;
assign n_24340 =  n_24332 &  n_24339;
assign n_24341 =  x_429 &  n_24340;
assign n_24342 = ~x_429 & ~n_24340;
assign n_24343 = ~n_24341 & ~n_24342;
assign n_24344 = ~x_1414 &  n_11;
assign n_24345 = ~x_1412 &  n_5;
assign n_24346 = ~n_24344 & ~n_24345;
assign n_24347 = ~x_1416 &  n_13;
assign n_24348 = ~x_1410 &  n_8;
assign n_24349 = ~n_24347 & ~n_24348;
assign n_24350 =  n_24346 &  n_24349;
assign n_24351 = ~x_1413 &  n_24;
assign n_24352 = ~x_1411 &  n_30;
assign n_24353 = ~n_24351 & ~n_24352;
assign n_24354 = ~x_1415 &  n_32;
assign n_24355 = ~x_1417 &  n_26;
assign n_24356 = ~n_24354 & ~n_24355;
assign n_24357 =  n_24353 &  n_24356;
assign n_24358 =  n_24350 &  n_24357;
assign n_24359 =  x_428 &  n_24358;
assign n_24360 = ~x_428 & ~n_24358;
assign n_24361 = ~n_24359 & ~n_24360;
assign n_24362 = ~x_1408 &  n_13;
assign n_24363 = ~x_1406 &  n_11;
assign n_24364 = ~n_24362 & ~n_24363;
assign n_24365 = ~x_1404 &  n_5;
assign n_24366 = ~x_1402 &  n_8;
assign n_24367 = ~n_24365 & ~n_24366;
assign n_24368 =  n_24364 &  n_24367;
assign n_24369 = ~x_1403 &  n_30;
assign n_24370 = ~x_1405 &  n_24;
assign n_24371 = ~n_24369 & ~n_24370;
assign n_24372 = ~x_1409 &  n_26;
assign n_24373 = ~x_1407 &  n_32;
assign n_24374 = ~n_24372 & ~n_24373;
assign n_24375 =  n_24371 &  n_24374;
assign n_24376 =  n_24368 &  n_24375;
assign n_24377 =  x_427 &  n_24376;
assign n_24378 = ~x_427 & ~n_24376;
assign n_24379 = ~n_24377 & ~n_24378;
assign n_24380 = ~x_1392 &  n_13;
assign n_24381 = ~x_1388 &  n_5;
assign n_24382 = ~n_24380 & ~n_24381;
assign n_24383 = ~x_1390 &  n_11;
assign n_24384 = ~x_1386 &  n_8;
assign n_24385 = ~n_24383 & ~n_24384;
assign n_24386 =  n_24382 &  n_24385;
assign n_24387 = ~x_1387 &  n_30;
assign n_24388 = ~x_1393 &  n_26;
assign n_24389 = ~n_24387 & ~n_24388;
assign n_24390 = ~x_1391 &  n_32;
assign n_24391 = ~x_1389 &  n_24;
assign n_24392 = ~n_24390 & ~n_24391;
assign n_24393 =  n_24389 &  n_24392;
assign n_24394 =  n_24386 &  n_24393;
assign n_24395 =  x_425 &  n_24394;
assign n_24396 = ~x_425 & ~n_24394;
assign n_24397 = ~n_24395 & ~n_24396;
assign n_24398 = ~x_1400 &  n_13;
assign n_24399 = ~x_1396 &  n_5;
assign n_24400 = ~n_24398 & ~n_24399;
assign n_24401 = ~x_1398 &  n_11;
assign n_24402 = ~x_1394 &  n_8;
assign n_24403 = ~n_24401 & ~n_24402;
assign n_24404 =  n_24400 &  n_24403;
assign n_24405 = ~x_1399 &  n_32;
assign n_24406 = ~x_1401 &  n_26;
assign n_24407 = ~n_24405 & ~n_24406;
assign n_24408 = ~x_1395 &  n_30;
assign n_24409 = ~x_1397 &  n_24;
assign n_24410 = ~n_24408 & ~n_24409;
assign n_24411 =  n_24407 &  n_24410;
assign n_24412 =  n_24404 &  n_24411;
assign n_24413 =  x_426 &  n_24412;
assign n_24414 = ~x_426 & ~n_24412;
assign n_24415 = ~n_24413 & ~n_24414;
assign n_24416 = ~n_24397 & ~n_24415;
assign n_24417 = ~n_24379 &  n_24416;
assign n_24418 = ~n_24361 &  n_24417;
assign n_24419 = ~n_24343 &  n_24418;
assign n_24420 = ~n_24325 &  n_24419;
assign n_24421 = ~n_24307 &  n_24420;
assign n_24422 = ~n_24289 &  n_24421;
assign n_24423 = ~n_24271 &  n_24422;
assign n_24424 = ~n_24253 &  n_24423;
assign n_24425 = ~n_24235 &  n_24424;
assign n_24426 = ~n_24217 &  n_24425;
assign n_24427 = ~n_24199 &  n_24426;
assign n_24428 = ~n_24181 &  n_24427;
assign n_24429 = ~n_24163 &  n_24428;
assign n_24430 = ~n_24145 &  n_24429;
assign n_24431 = ~n_24127 &  n_24430;
assign n_24432 = ~n_24109 &  n_24431;
assign n_24433 = ~n_24091 &  n_24432;
assign n_24434 = ~n_24073 &  n_24433;
assign n_24435 = ~n_24055 &  n_24434;
assign n_24436 = ~n_24037 &  n_24435;
assign n_24437 = ~n_24019 &  n_24436;
assign n_24438 = ~n_24001 &  n_24437;
assign n_24439 = ~n_23983 &  n_24438;
assign n_24440 = ~n_23965 &  n_24439;
assign n_24441 = ~n_23947 &  n_24440;
assign n_24442 = ~n_23944 &  n_24441;
assign n_24443 = ~n_23941 &  n_24442;
assign n_24444 = ~n_23935 &  n_24443;
assign n_24445 = ~n_23930 &  n_24444;
assign n_24446 = ~n_23925 &  n_24445;
assign n_24447 = ~n_23920 &  n_24446;
assign n_24448 = ~n_23914 &  n_24447;
assign n_24449 = ~n_23908 &  n_24448;
assign n_24450 = ~n_23902 &  n_24449;
assign n_24451 = ~n_23896 &  n_24450;
assign n_24452 = ~n_23890 &  n_24451;
assign n_24453 = ~n_23884 &  n_24452;
assign n_24454 = ~n_23878 &  n_24453;
assign n_24455 = ~n_23872 &  n_24454;
assign n_24456 = ~n_23866 &  n_24455;
assign n_24457 = ~n_23860 &  n_24456;
assign n_24458 = ~n_23854 &  n_24457;
assign n_24459 = ~n_23848 &  n_24458;
assign n_24460 = ~n_23842 &  n_24459;
assign n_24461 = ~n_23836 &  n_24460;
assign n_24462 = ~n_23830 &  n_24461;
assign n_24463 = ~n_23824 &  n_24462;
assign n_24464 = ~n_23818 &  n_24463;
assign n_24465 = ~n_23812 &  n_24464;
assign n_24466 = ~n_23806 &  n_24465;
assign n_24467 = ~n_23800 &  n_24466;
assign n_24468 = ~n_23794 &  n_24467;
assign n_24469 = ~n_23788 &  n_24468;
assign n_24470 = ~n_23782 &  n_24469;
assign n_24471 = ~n_23776 &  n_24470;
assign n_24472 = ~n_23770 &  n_24471;
assign n_24473 = ~n_23764 &  n_24472;
assign n_24474 = ~n_23758 &  n_24473;
assign n_24475 = ~n_23752 &  n_24474;
assign n_24476 = ~n_23714 &  n_24475;
assign n_24477 = ~n_23708 &  n_24476;
assign n_24478 = ~n_23702 &  n_24477;
assign n_24479 = ~n_23696 &  n_24478;
assign n_24480 = ~n_23690 &  n_24479;
assign n_24481 = ~n_23684 &  n_24480;
assign n_24482 = ~n_23678 &  n_24481;
assign n_24483 = ~n_23672 &  n_24482;
assign n_24484 = ~n_23666 &  n_24483;
assign n_24485 = ~n_23660 &  n_24484;
assign n_24486 = ~n_23654 &  n_24485;
assign n_24487 = ~n_23647 &  n_24486;
assign n_24488 = ~n_23641 &  n_24487;
assign n_24489 = ~n_23635 &  n_24488;
assign n_24490 = ~n_23629 &  n_24489;
assign n_24491 = ~n_23623 &  n_24490;
assign n_24492 = ~n_23617 &  n_24491;
assign n_24493 = ~n_23611 &  n_24492;
assign n_24494 = ~n_23605 &  n_24493;
assign n_24495 = ~n_23599 &  n_24494;
assign n_24496 = ~n_23593 &  n_24495;
assign n_24497 = ~n_23587 &  n_24496;
assign n_24498 = ~n_23581 &  n_24497;
assign n_24499 = ~n_23574 &  n_24498;
assign n_24500 = ~n_23568 &  n_24499;
assign n_24501 = ~n_23562 &  n_24500;
assign n_24502 = ~n_23556 &  n_24501;
assign n_24503 = ~n_23550 &  n_24502;
assign n_24504 = ~n_23544 &  n_24503;
assign n_24505 = ~n_23538 &  n_24504;
assign n_24506 = ~n_23532 &  n_24505;
assign n_24507 = ~n_23526 &  n_24506;
assign n_24508 = ~n_23520 &  n_24507;
assign n_24509 = ~n_23514 &  n_24508;
assign n_24510 = ~n_23508 &  n_24509;
assign n_24511 = ~n_23501 &  n_24510;
assign n_24512 = ~n_23495 &  n_24511;
assign n_24513 = ~n_23489 &  n_24512;
assign n_24514 = ~n_23483 &  n_24513;
assign n_24515 = ~n_23477 &  n_24514;
assign n_24516 = ~n_23471 &  n_24515;
assign n_24517 = ~n_23465 &  n_24516;
assign n_24518 = ~n_23459 &  n_24517;
assign n_24519 = ~n_23453 &  n_24518;
assign n_24520 = ~n_23447 &  n_24519;
assign n_24521 = ~n_23441 &  n_24520;
assign n_24522 = ~n_23435 &  n_24521;
assign n_24523 = ~n_23428 &  n_24522;
assign n_24524 = ~n_23422 &  n_24523;
assign n_24525 = ~n_23416 &  n_24524;
assign n_24526 = ~n_23410 &  n_24525;
assign n_24527 = ~n_23404 &  n_24526;
assign n_24528 = ~n_23398 &  n_24527;
assign n_24529 = ~n_23392 &  n_24528;
assign n_24530 = ~n_23386 &  n_24529;
assign n_24531 = ~n_23380 &  n_24530;
assign n_24532 = ~n_23374 &  n_24531;
assign n_24533 = ~n_23368 &  n_24532;
assign n_24534 = ~n_23362 &  n_24533;
assign n_24535 = ~n_23355 &  n_24534;
assign n_24536 = ~n_23349 &  n_24535;
assign n_24537 = ~n_23343 &  n_24536;
assign n_24538 = ~n_23337 &  n_24537;
assign n_24539 = ~n_23331 &  n_24538;
assign n_24540 = ~n_23325 &  n_24539;
assign n_24541 = ~n_23319 &  n_24540;
assign n_24542 = ~n_23313 &  n_24541;
assign n_24543 = ~n_23307 &  n_24542;
assign n_24544 = ~n_23301 &  n_24543;
assign n_24545 = ~n_23295 &  n_24544;
assign n_24546 = ~n_23289 &  n_24545;
assign n_24547 = ~n_23282 &  n_24546;
assign n_24548 = ~n_23276 &  n_24547;
assign n_24549 = ~n_23270 &  n_24548;
assign n_24550 = ~n_23264 &  n_24549;
assign n_24551 = ~n_23258 &  n_24550;
assign n_24552 = ~n_23252 &  n_24551;
assign n_24553 = ~n_23246 &  n_24552;
assign n_24554 = ~n_23240 &  n_24553;
assign n_24555 = ~n_23234 &  n_24554;
assign n_24556 = ~n_23228 &  n_24555;
assign n_24557 = ~n_23222 &  n_24556;
assign n_24558 = ~n_23216 &  n_24557;
assign n_24559 = ~n_23209 &  n_24558;
assign n_24560 = ~n_23203 &  n_24559;
assign n_24561 = ~n_23197 &  n_24560;
assign n_24562 = ~n_23191 &  n_24561;
assign n_24563 = ~n_23185 &  n_24562;
assign n_24564 = ~n_23179 &  n_24563;
assign n_24565 = ~n_23173 &  n_24564;
assign n_24566 = ~n_23167 &  n_24565;
assign n_24567 = ~n_23161 &  n_24566;
assign n_24568 = ~n_23155 &  n_24567;
assign n_24569 = ~n_23149 &  n_24568;
assign n_24570 = ~n_23143 &  n_24569;
assign n_24571 = ~n_23136 &  n_24570;
assign n_24572 = ~n_23130 &  n_24571;
assign n_24573 = ~n_23124 &  n_24572;
assign n_24574 = ~n_23118 &  n_24573;
assign n_24575 = ~n_23112 &  n_24574;
assign n_24576 = ~n_23106 &  n_24575;
assign n_24577 = ~n_23100 &  n_24576;
assign n_24578 = ~n_23094 &  n_24577;
assign n_24579 = ~n_23088 &  n_24578;
assign n_24580 = ~n_23082 &  n_24579;
assign n_24581 = ~n_23076 &  n_24580;
assign n_24582 = ~n_23070 &  n_24581;
assign n_24583 = ~n_23063 &  n_24582;
assign n_24584 = ~n_23057 &  n_24583;
assign n_24585 = ~n_23051 &  n_24584;
assign n_24586 = ~n_23045 &  n_24585;
assign n_24587 = ~n_23039 &  n_24586;
assign n_24588 = ~n_23033 &  n_24587;
assign n_24589 = ~n_23027 &  n_24588;
assign n_24590 = ~n_23021 &  n_24589;
assign n_24591 = ~n_23015 &  n_24590;
assign n_24592 = ~n_23009 &  n_24591;
assign n_24593 = ~n_23003 &  n_24592;
assign n_24594 = ~n_22997 &  n_24593;
assign n_24595 = ~n_22990 &  n_24594;
assign n_24596 = ~n_22984 &  n_24595;
assign n_24597 = ~n_22978 &  n_24596;
assign n_24598 = ~n_22972 &  n_24597;
assign n_24599 = ~n_22966 &  n_24598;
assign n_24600 = ~n_22960 &  n_24599;
assign n_24601 = ~n_22954 &  n_24600;
assign n_24602 = ~n_22948 &  n_24601;
assign n_24603 = ~n_22942 &  n_24602;
assign n_24604 = ~n_22936 &  n_24603;
assign n_24605 = ~n_22930 &  n_24604;
assign n_24606 = ~n_22924 &  n_24605;
assign n_24607 = ~n_22917 &  n_24606;
assign n_24608 = ~n_22911 &  n_24607;
assign n_24609 = ~n_22905 &  n_24608;
assign n_24610 = ~n_22899 &  n_24609;
assign n_24611 = ~n_22893 &  n_24610;
assign n_24612 = ~n_22887 &  n_24611;
assign n_24613 = ~n_22881 &  n_24612;
assign n_24614 = ~n_22875 &  n_24613;
assign n_24615 = ~n_22869 &  n_24614;
assign n_24616 = ~n_22863 &  n_24615;
assign n_24617 = ~n_22857 &  n_24616;
assign n_24618 = ~n_22851 &  n_24617;
assign n_24619 = ~n_22844 &  n_24618;
assign n_24620 = ~n_22838 &  n_24619;
assign n_24621 = ~n_22832 &  n_24620;
assign n_24622 = ~n_22826 &  n_24621;
assign n_24623 = ~n_22820 &  n_24622;
assign n_24624 = ~n_22814 &  n_24623;
assign n_24625 = ~n_22808 &  n_24624;
assign n_24626 = ~n_22802 &  n_24625;
assign n_24627 = ~n_22796 &  n_24626;
assign n_24628 = ~n_22790 &  n_24627;
assign n_24629 = ~n_22784 &  n_24628;
assign n_24630 = ~n_22778 &  n_24629;
assign n_24631 = ~n_22771 &  n_24630;
assign n_24632 = ~n_22765 &  n_24631;
assign n_24633 = ~n_22759 &  n_24632;
assign n_24634 = ~n_22753 &  n_24633;
assign n_24635 = ~n_22747 &  n_24634;
assign n_24636 = ~n_22741 &  n_24635;
assign n_24637 = ~n_22735 &  n_24636;
assign n_24638 = ~n_22729 &  n_24637;
assign n_24639 = ~n_22723 &  n_24638;
assign n_24640 = ~n_22717 &  n_24639;
assign n_24641 = ~n_22711 &  n_24640;
assign n_24642 = ~n_22705 &  n_24641;
assign n_24643 = ~n_22698 &  n_24642;
assign n_24644 = ~n_22692 &  n_24643;
assign n_24645 = ~n_22686 &  n_24644;
assign n_24646 = ~n_22680 &  n_24645;
assign n_24647 = ~n_22674 &  n_24646;
assign n_24648 = ~n_22668 &  n_24647;
assign n_24649 = ~n_22662 &  n_24648;
assign n_24650 = ~n_22656 &  n_24649;
assign n_24651 = ~n_22650 &  n_24650;
assign n_24652 = ~n_22644 &  n_24651;
assign n_24653 = ~n_22638 &  n_24652;
assign n_24654 = ~n_22632 &  n_24653;
assign n_24655 = ~n_22625 &  n_24654;
assign n_24656 = ~n_22619 &  n_24655;
assign n_24657 = ~n_22613 &  n_24656;
assign n_24658 = ~n_22607 &  n_24657;
assign n_24659 = ~n_22601 &  n_24658;
assign n_24660 = ~n_22595 &  n_24659;
assign n_24661 = ~n_22589 &  n_24660;
assign n_24662 = ~n_22583 &  n_24661;
assign n_24663 = ~n_22577 &  n_24662;
assign n_24664 = ~n_22571 &  n_24663;
assign n_24665 = ~n_22565 &  n_24664;
assign n_24666 = ~n_22559 &  n_24665;
assign n_24667 = ~n_22552 &  n_24666;
assign n_24668 = ~n_22546 &  n_24667;
assign n_24669 = ~n_22540 &  n_24668;
assign n_24670 = ~n_22534 &  n_24669;
assign n_24671 = ~n_22528 &  n_24670;
assign n_24672 = ~n_22522 &  n_24671;
assign n_24673 = ~n_22516 &  n_24672;
assign n_24674 = ~n_22510 &  n_24673;
assign n_24675 = ~n_22504 &  n_24674;
assign n_24676 = ~n_22498 &  n_24675;
assign n_24677 = ~n_22492 &  n_24676;
assign n_24678 = ~n_22486 &  n_24677;
assign n_24679 = ~n_22479 &  n_24678;
assign n_24680 = ~n_22473 &  n_24679;
assign n_24681 = ~n_22467 &  n_24680;
assign n_24682 = ~n_22461 &  n_24681;
assign n_24683 = ~n_22455 &  n_24682;
assign n_24684 = ~n_22449 &  n_24683;
assign n_24685 = ~n_22443 &  n_24684;
assign n_24686 = ~n_22437 &  n_24685;
assign n_24687 = ~n_22431 &  n_24686;
assign n_24688 = ~n_22425 &  n_24687;
assign n_24689 = ~n_22419 &  n_24688;
assign n_24690 = ~n_22413 &  n_24689;
assign n_24691 = ~n_22406 &  n_24690;
assign n_24692 = ~n_22400 &  n_24691;
assign n_24693 = ~n_22394 &  n_24692;
assign n_24694 = ~n_22388 &  n_24693;
assign n_24695 = ~n_22382 &  n_24694;
assign n_24696 = ~n_22376 &  n_24695;
assign n_24697 = ~n_22370 &  n_24696;
assign n_24698 = ~n_22364 &  n_24697;
assign n_24699 = ~n_22358 &  n_24698;
assign n_24700 = ~n_22352 &  n_24699;
assign n_24701 = ~n_22346 &  n_24700;
assign n_24702 = ~n_22340 &  n_24701;
assign n_24703 = ~n_22333 &  n_24702;
assign n_24704 = ~n_22327 &  n_24703;
assign n_24705 = ~n_22321 &  n_24704;
assign n_24706 = ~n_22315 &  n_24705;
assign n_24707 = ~n_22309 &  n_24706;
assign n_24708 = ~n_22303 &  n_24707;
assign n_24709 = ~n_22297 &  n_24708;
assign n_24710 = ~n_22291 &  n_24709;
assign n_24711 = ~n_22285 &  n_24710;
assign n_24712 = ~n_22279 &  n_24711;
assign n_24713 = ~n_22273 &  n_24712;
assign n_24714 = ~n_22267 &  n_24713;
assign n_24715 = ~n_22260 &  n_24714;
assign n_24716 = ~n_22254 &  n_24715;
assign n_24717 = ~n_22248 &  n_24716;
assign n_24718 = ~n_22242 &  n_24717;
assign n_24719 = ~n_22236 &  n_24718;
assign n_24720 = ~n_22230 &  n_24719;
assign n_24721 = ~n_22224 &  n_24720;
assign n_24722 = ~n_22218 &  n_24721;
assign n_24723 = ~n_22212 &  n_24722;
assign n_24724 = ~n_22206 &  n_24723;
assign n_24725 = ~n_22200 &  n_24724;
assign n_24726 = ~n_22194 &  n_24725;
assign n_24727 = ~n_22187 &  n_24726;
assign n_24728 = ~n_22181 &  n_24727;
assign n_24729 = ~n_22175 &  n_24728;
assign n_24730 = ~n_22169 &  n_24729;
assign n_24731 = ~n_22163 &  n_24730;
assign n_24732 = ~n_22157 &  n_24731;
assign n_24733 = ~n_22151 &  n_24732;
assign n_24734 = ~n_22145 &  n_24733;
assign n_24735 = ~n_22139 &  n_24734;
assign n_24736 = ~n_22133 &  n_24735;
assign n_24737 = ~n_22127 &  n_24736;
assign n_24738 = ~n_22121 &  n_24737;
assign n_24739 = ~n_22114 &  n_24738;
assign n_24740 = ~n_22108 &  n_24739;
assign n_24741 = ~n_22102 &  n_24740;
assign n_24742 = ~n_22096 &  n_24741;
assign n_24743 = ~n_22090 &  n_24742;
assign n_24744 = ~n_22084 &  n_24743;
assign n_24745 = ~n_22078 &  n_24744;
assign n_24746 = ~n_22072 &  n_24745;
assign n_24747 = ~n_22066 &  n_24746;
assign n_24748 = ~n_22060 &  n_24747;
assign n_24749 = ~n_22054 &  n_24748;
assign n_24750 = ~n_22048 &  n_24749;
assign n_24751 = ~n_22041 &  n_24750;
assign n_24752 = ~n_22035 &  n_24751;
assign n_24753 = ~n_22029 &  n_24752;
assign n_24754 = ~n_22023 &  n_24753;
assign n_24755 = ~n_22017 &  n_24754;
assign n_24756 = ~n_22011 &  n_24755;
assign n_24757 = ~n_22005 &  n_24756;
assign n_24758 = ~n_21999 &  n_24757;
assign n_24759 = ~n_21993 &  n_24758;
assign n_24760 = ~n_21987 &  n_24759;
assign n_24761 = ~n_21981 &  n_24760;
assign n_24762 = ~n_21975 &  n_24761;
assign n_24763 = ~n_21968 &  n_24762;
assign n_24764 = ~n_21962 &  n_24763;
assign n_24765 = ~n_21956 &  n_24764;
assign n_24766 = ~n_21950 &  n_24765;
assign n_24767 = ~n_21944 &  n_24766;
assign n_24768 = ~n_21938 &  n_24767;
assign n_24769 = ~n_21932 &  n_24768;
assign n_24770 = ~n_21926 &  n_24769;
assign n_24771 = ~n_21920 &  n_24770;
assign n_24772 = ~n_21914 &  n_24771;
assign n_24773 = ~n_21908 &  n_24772;
assign n_24774 = ~n_21902 &  n_24773;
assign n_24775 = ~n_21895 &  n_24774;
assign n_24776 = ~n_21889 &  n_24775;
assign n_24777 = ~n_21883 &  n_24776;
assign n_24778 = ~n_21877 &  n_24777;
assign n_24779 = ~n_21871 &  n_24778;
assign n_24780 = ~n_21865 &  n_24779;
assign n_24781 = ~n_21859 &  n_24780;
assign n_24782 = ~n_21853 &  n_24781;
assign n_24783 = ~n_21847 &  n_24782;
assign n_24784 = ~n_21841 &  n_24783;
assign n_24785 = ~n_21835 &  n_24784;
assign n_24786 = ~n_21829 &  n_24785;
assign n_24787 = ~n_21822 &  n_24786;
assign n_24788 = ~n_21816 &  n_24787;
assign n_24789 = ~n_21810 &  n_24788;
assign n_24790 = ~n_21804 &  n_24789;
assign n_24791 = ~n_21798 &  n_24790;
assign n_24792 = ~n_21792 &  n_24791;
assign n_24793 = ~n_21786 &  n_24792;
assign n_24794 = ~n_21780 &  n_24793;
assign n_24795 = ~n_21774 &  n_24794;
assign n_24796 = ~n_21768 &  n_24795;
assign n_24797 = ~n_21762 &  n_24796;
assign n_24798 = ~n_21756 &  n_24797;
assign n_24799 = ~n_21749 &  n_24798;
assign n_24800 = ~n_21743 &  n_24799;
assign n_24801 = ~n_21737 &  n_24800;
assign n_24802 = ~n_21731 &  n_24801;
assign n_24803 = ~n_21725 &  n_24802;
assign n_24804 = ~n_21719 &  n_24803;
assign n_24805 = ~n_21713 &  n_24804;
assign n_24806 = ~n_21707 &  n_24805;
assign n_24807 = ~n_21701 &  n_24806;
assign n_24808 = ~n_21695 &  n_24807;
assign n_24809 = ~n_21689 &  n_24808;
assign n_24810 = ~n_21683 &  n_24809;
assign n_24811 = ~n_21676 &  n_24810;
assign n_24812 = ~n_21670 &  n_24811;
assign n_24813 = ~n_21664 &  n_24812;
assign n_24814 = ~n_21658 &  n_24813;
assign n_24815 = ~n_21652 &  n_24814;
assign n_24816 = ~n_21646 &  n_24815;
assign n_24817 = ~n_21640 &  n_24816;
assign n_24818 = ~n_21634 &  n_24817;
assign n_24819 = ~n_21628 &  n_24818;
assign n_24820 = ~n_21622 &  n_24819;
assign n_24821 = ~n_21616 &  n_24820;
assign n_24822 = ~n_21610 &  n_24821;
assign n_24823 = ~n_21603 &  n_24822;
assign n_24824 = ~n_21597 &  n_24823;
assign n_24825 = ~n_21591 &  n_24824;
assign n_24826 = ~n_21585 &  n_24825;
assign n_24827 = ~n_21579 &  n_24826;
assign n_24828 = ~n_21573 &  n_24827;
assign n_24829 = ~n_21567 &  n_24828;
assign n_24830 = ~n_21561 &  n_24829;
assign n_24831 = ~n_21555 &  n_24830;
assign n_24832 = ~n_21549 &  n_24831;
assign n_24833 = ~n_21543 &  n_24832;
assign n_24834 = ~n_21537 &  n_24833;
assign n_24835 = ~n_21530 &  n_24834;
assign n_24836 = ~n_21524 &  n_24835;
assign n_24837 = ~n_21518 &  n_24836;
assign n_24838 = ~n_21512 &  n_24837;
assign n_24839 = ~n_21506 &  n_24838;
assign n_24840 = ~n_21500 &  n_24839;
assign n_24841 = ~n_21494 &  n_24840;
assign n_24842 = ~n_21488 &  n_24841;
assign n_24843 = ~n_21482 &  n_24842;
assign n_24844 = ~n_21476 &  n_24843;
assign n_24845 = ~n_21470 &  n_24844;
assign n_24846 = ~n_21464 &  n_24845;
assign n_24847 = ~n_21457 &  n_24846;
assign n_24848 = ~n_21451 &  n_24847;
assign n_24849 = ~n_21445 &  n_24848;
assign n_24850 = ~n_21439 &  n_24849;
assign n_24851 = ~n_21433 &  n_24850;
assign n_24852 = ~n_21427 &  n_24851;
assign n_24853 = ~n_21421 &  n_24852;
assign n_24854 = ~n_21415 &  n_24853;
assign n_24855 = ~n_21409 &  n_24854;
assign n_24856 = ~n_21403 &  n_24855;
assign n_24857 = ~n_21397 &  n_24856;
assign n_24858 = ~n_21391 &  n_24857;
assign n_24859 = ~n_21384 &  n_24858;
assign n_24860 = ~n_21376 &  n_24859;
assign n_24861 = ~n_21368 &  n_24860;
assign n_24862 = ~n_21359 &  n_24861;
assign n_24863 = ~n_21351 &  n_24862;
assign n_24864 = ~n_21343 &  n_24863;
assign n_24865 = ~n_21334 &  n_24864;
assign n_24866 = ~n_21325 &  n_24865;
assign n_24867 = ~n_21317 &  n_24866;
assign n_24868 = ~n_21309 &  n_24867;
assign n_24869 = ~n_21299 &  n_24868;
assign n_24870 = ~n_21288 &  n_24869;
assign n_24871 = ~n_21248 &  n_24870;
assign n_24872 = ~n_21243 &  n_24871;
assign n_24873 = ~n_21238 &  n_24872;
assign n_24874 = ~n_21233 &  n_24873;
assign n_24875 = ~n_21227 &  n_24874;
assign n_24876 = ~n_21221 &  n_24875;
assign n_24877 = ~n_21215 &  n_24876;
assign n_24878 = ~n_21209 &  n_24877;
assign n_24879 = ~n_21203 &  n_24878;
assign n_24880 = ~n_21197 &  n_24879;
assign n_24881 = ~n_21191 &  n_24880;
assign n_24882 = ~n_21184 &  n_24881;
assign n_24883 = ~n_21178 &  n_24882;
assign n_24884 = ~n_21172 &  n_24883;
assign n_24885 = ~n_21166 &  n_24884;
assign n_24886 = ~n_21160 &  n_24885;
assign n_24887 = ~n_21154 &  n_24886;
assign n_24888 = ~n_21148 &  n_24887;
assign n_24889 = ~n_21142 &  n_24888;
assign n_24890 = ~n_21135 &  n_24889;
assign n_24891 = ~n_21129 &  n_24890;
assign n_24892 = ~n_21123 &  n_24891;
assign n_24893 = ~n_21117 &  n_24892;
assign n_24894 = ~n_21111 &  n_24893;
assign n_24895 = ~n_21105 &  n_24894;
assign n_24896 = ~n_21099 &  n_24895;
assign n_24897 = ~n_21093 &  n_24896;
assign n_24898 = ~n_21086 &  n_24897;
assign n_24899 = ~n_21080 &  n_24898;
assign n_24900 = ~n_21074 &  n_24899;
assign n_24901 = ~n_21068 &  n_24900;
assign n_24902 = ~n_21062 &  n_24901;
assign n_24903 = ~n_21056 &  n_24902;
assign n_24904 = ~n_21050 &  n_24903;
assign n_24905 = ~n_21044 &  n_24904;
assign n_24906 = ~n_21037 &  n_24905;
assign n_24907 = ~n_21031 &  n_24906;
assign n_24908 = ~n_21025 &  n_24907;
assign n_24909 = ~n_21019 &  n_24908;
assign n_24910 = ~n_21013 &  n_24909;
assign n_24911 = ~n_21007 &  n_24910;
assign n_24912 = ~n_21001 &  n_24911;
assign n_24913 = ~n_20995 &  n_24912;
assign n_24914 = ~n_20988 &  n_24913;
assign n_24915 = ~n_20982 &  n_24914;
assign n_24916 = ~n_20976 &  n_24915;
assign n_24917 = ~n_20970 &  n_24916;
assign n_24918 = ~n_20964 &  n_24917;
assign n_24919 = ~n_20958 &  n_24918;
assign n_24920 = ~n_20952 &  n_24919;
assign n_24921 = ~n_20946 &  n_24920;
assign n_24922 = ~n_20939 &  n_24921;
assign n_24923 = ~n_20933 &  n_24922;
assign n_24924 = ~n_20927 &  n_24923;
assign n_24925 = ~n_20921 &  n_24924;
assign n_24926 = ~n_20915 &  n_24925;
assign n_24927 = ~n_20909 &  n_24926;
assign n_24928 = ~n_20903 &  n_24927;
assign n_24929 = ~n_20897 &  n_24928;
assign n_24930 = ~n_20890 &  n_24929;
assign n_24931 = ~n_20884 &  n_24930;
assign n_24932 = ~n_20878 &  n_24931;
assign n_24933 = ~n_20872 &  n_24932;
assign n_24934 = ~n_20866 &  n_24933;
assign n_24935 = ~n_20860 &  n_24934;
assign n_24936 = ~n_20854 &  n_24935;
assign n_24937 = ~n_20848 &  n_24936;
assign n_24938 = ~n_20841 &  n_24937;
assign n_24939 = ~n_20835 &  n_24938;
assign n_24940 = ~n_20829 &  n_24939;
assign n_24941 = ~n_20823 &  n_24940;
assign n_24942 = ~n_20817 &  n_24941;
assign n_24943 = ~n_20811 &  n_24942;
assign n_24944 = ~n_20805 &  n_24943;
assign n_24945 = ~n_20799 &  n_24944;
assign n_24946 = ~n_20793 &  n_24945;
assign n_24947 = ~n_20787 &  n_24946;
assign n_24948 = ~n_20781 &  n_24947;
assign n_24949 = ~n_20775 &  n_24948;
assign n_24950 = ~n_20769 &  n_24949;
assign n_24951 = ~n_20763 &  n_24950;
assign n_24952 = ~n_20757 &  n_24951;
assign n_24953 = ~n_20751 &  n_24952;
assign n_24954 = ~n_20745 &  n_24953;
assign n_24955 = ~n_20739 &  n_24954;
assign n_24956 = ~n_20733 &  n_24955;
assign n_24957 = ~n_20727 &  n_24956;
assign n_24958 = ~n_20721 &  n_24957;
assign n_24959 = ~n_20715 &  n_24958;
assign n_24960 = ~n_20709 &  n_24959;
assign n_24961 = ~n_20703 &  n_24960;
assign n_24962 = ~n_20697 &  n_24961;
assign n_24963 = ~n_20691 &  n_24962;
assign n_24964 = ~n_20685 &  n_24963;
assign n_24965 = ~n_20679 &  n_24964;
assign n_24966 = ~n_20673 &  n_24965;
assign n_24967 = ~n_20667 &  n_24966;
assign n_24968 = ~n_20661 &  n_24967;
assign n_24969 = ~n_20655 &  n_24968;
assign n_24970 = ~n_20649 &  n_24969;
assign n_24971 = ~n_20643 &  n_24970;
assign n_24972 = ~n_20637 &  n_24971;
assign n_24973 = ~n_20631 &  n_24972;
assign n_24974 = ~n_20625 &  n_24973;
assign n_24975 = ~n_20619 &  n_24974;
assign n_24976 = ~n_20613 &  n_24975;
assign n_24977 = ~n_20607 &  n_24976;
assign n_24978 = ~n_20601 &  n_24977;
assign n_24979 = ~n_20595 &  n_24978;
assign n_24980 = ~n_20589 &  n_24979;
assign n_24981 = ~n_20583 &  n_24980;
assign n_24982 = ~n_20577 &  n_24981;
assign n_24983 = ~n_20571 &  n_24982;
assign n_24984 = ~n_20565 &  n_24983;
assign n_24985 = ~n_20559 &  n_24984;
assign n_24986 = ~n_20553 &  n_24985;
assign n_24987 = ~n_20547 &  n_24986;
assign n_24988 = ~n_20541 &  n_24987;
assign n_24989 = ~n_20535 &  n_24988;
assign n_24990 = ~n_20529 &  n_24989;
assign n_24991 = ~n_20523 &  n_24990;
assign n_24992 = ~n_20517 &  n_24991;
assign n_24993 = ~n_20511 &  n_24992;
assign n_24994 = ~n_20505 &  n_24993;
assign n_24995 = ~n_20499 &  n_24994;
assign n_24996 = ~n_20493 &  n_24995;
assign n_24997 = ~n_20487 &  n_24996;
assign n_24998 = ~n_20481 &  n_24997;
assign n_24999 = ~n_20475 &  n_24998;
assign n_25000 = ~n_20469 &  n_24999;
assign n_25001 = ~n_20463 &  n_25000;
assign n_25002 = ~n_20457 &  n_25001;
assign n_25003 = ~n_20451 &  n_25002;
assign n_25004 = ~n_20445 &  n_25003;
assign n_25005 = ~n_20439 &  n_25004;
assign n_25006 = ~n_20433 &  n_25005;
assign n_25007 = ~n_20427 &  n_25006;
assign n_25008 = ~n_20421 &  n_25007;
assign n_25009 = ~n_20415 &  n_25008;
assign n_25010 = ~n_20409 &  n_25009;
assign n_25011 = ~n_20403 &  n_25010;
assign n_25012 = ~n_20396 &  n_25011;
assign n_25013 = ~n_20390 &  n_25012;
assign n_25014 = ~n_20384 &  n_25013;
assign n_25015 = ~n_20378 &  n_25014;
assign n_25016 = ~n_20372 &  n_25015;
assign n_25017 = ~n_20366 &  n_25016;
assign n_25018 = ~n_20360 &  n_25017;
assign n_25019 = ~n_20354 &  n_25018;
assign n_25020 = ~n_20347 &  n_25019;
assign n_25021 = ~n_20344 &  n_25020;
assign n_25022 = ~n_20338 &  n_25021;
assign n_25023 = ~n_20332 &  n_25022;
assign n_25024 = ~n_20326 &  n_25023;
assign n_25025 = ~n_20320 &  n_25024;
assign n_25026 = ~n_20314 &  n_25025;
assign n_25027 = ~n_20308 &  n_25026;
assign n_25028 = ~n_20302 &  n_25027;
assign n_25029 = ~n_20295 &  n_25028;
assign n_25030 = ~n_20292 &  n_25029;
assign n_25031 = ~n_20286 &  n_25030;
assign n_25032 = ~n_20280 &  n_25031;
assign n_25033 = ~n_20274 &  n_25032;
assign n_25034 = ~n_20268 &  n_25033;
assign n_25035 = ~n_20262 &  n_25034;
assign n_25036 = ~n_20256 &  n_25035;
assign n_25037 = ~n_20250 &  n_25036;
assign n_25038 = ~n_20243 &  n_25037;
assign n_25039 = ~n_20240 &  n_25038;
assign n_25040 = ~n_20234 &  n_25039;
assign n_25041 = ~n_20228 &  n_25040;
assign n_25042 = ~n_20222 &  n_25041;
assign n_25043 = ~n_20216 &  n_25042;
assign n_25044 = ~n_20210 &  n_25043;
assign n_25045 = ~n_20204 &  n_25044;
assign n_25046 = ~n_20198 &  n_25045;
assign n_25047 = ~n_20191 &  n_25046;
assign n_25048 = ~n_20188 &  n_25047;
assign n_25049 = ~n_20182 &  n_25048;
assign n_25050 = ~n_20176 &  n_25049;
assign n_25051 = ~n_20170 &  n_25050;
assign n_25052 = ~n_20164 &  n_25051;
assign n_25053 = ~n_20158 &  n_25052;
assign n_25054 = ~n_20152 &  n_25053;
assign n_25055 = ~n_20146 &  n_25054;
assign n_25056 = ~n_20139 &  n_25055;
assign n_25057 = ~n_20136 &  n_25056;
assign n_25058 = ~n_20130 &  n_25057;
assign n_25059 = ~n_20124 &  n_25058;
assign n_25060 = ~n_20118 &  n_25059;
assign n_25061 = ~n_20112 &  n_25060;
assign n_25062 = ~n_20106 &  n_25061;
assign n_25063 = ~n_20100 &  n_25062;
assign n_25064 = ~n_20094 &  n_25063;
assign n_25065 = ~n_20087 &  n_25064;
assign n_25066 = ~n_20084 &  n_25065;
assign n_25067 = ~n_20078 &  n_25066;
assign n_25068 = ~n_20072 &  n_25067;
assign n_25069 = ~n_20066 &  n_25068;
assign n_25070 = ~n_20060 &  n_25069;
assign n_25071 = ~n_20054 &  n_25070;
assign n_25072 = ~n_20048 &  n_25071;
assign n_25073 = ~n_20042 &  n_25072;
assign n_25074 = ~n_20035 &  n_25073;
assign n_25075 = ~n_20032 &  n_25074;
assign n_25076 = ~n_20029 &  n_25075;
assign n_25077 = ~n_20026 &  n_25076;
assign n_25078 = ~n_20023 &  n_25077;
assign n_25079 = ~n_20020 &  n_25078;
assign n_25080 = ~n_20017 &  n_25079;
assign n_25081 = ~n_20014 &  n_25080;
assign n_25082 = ~n_20011 &  n_25081;
assign n_25083 = ~n_20008 &  n_25082;
assign n_25084 = ~n_20005 &  n_25083;
assign n_25085 = ~n_20002 &  n_25084;
assign n_25086 = ~n_19999 &  n_25085;
assign n_25087 = ~n_19996 &  n_25086;
assign n_25088 = ~n_19993 &  n_25087;
assign n_25089 = ~n_19990 &  n_25088;
assign n_25090 = ~n_19987 &  n_25089;
assign n_25091 = ~n_19984 &  n_25090;
assign n_25092 = ~n_19981 &  n_25091;
assign n_25093 = ~n_19978 &  n_25092;
assign n_25094 = ~n_19975 &  n_25093;
assign n_25095 = ~n_19972 &  n_25094;
assign n_25096 = ~n_19969 &  n_25095;
assign n_25097 = ~n_19966 &  n_25096;
assign n_25098 = ~n_19963 &  n_25097;
assign n_25099 = ~n_19960 &  n_25098;
assign n_25100 = ~n_19957 &  n_25099;
assign n_25101 = ~n_19954 &  n_25100;
assign n_25102 = ~n_19951 &  n_25101;
assign n_25103 = ~n_19948 &  n_25102;
assign n_25104 = ~n_19945 &  n_25103;
assign n_25105 = ~n_19942 &  n_25104;
assign n_25106 = ~n_19939 &  n_25105;
assign n_25107 = ~n_19936 &  n_25106;
assign n_25108 = ~n_19933 &  n_25107;
assign n_25109 = ~n_19930 &  n_25108;
assign n_25110 = ~n_19927 &  n_25109;
assign n_25111 = ~n_19924 &  n_25110;
assign n_25112 = ~n_19921 &  n_25111;
assign n_25113 = ~n_19918 &  n_25112;
assign n_25114 = ~n_19915 &  n_25113;
assign n_25115 = ~n_19912 &  n_25114;
assign n_25116 = ~n_19909 &  n_25115;
assign n_25117 = ~n_19906 &  n_25116;
assign n_25118 = ~n_19903 &  n_25117;
assign n_25119 = ~n_19900 &  n_25118;
assign n_25120 = ~n_19897 &  n_25119;
assign n_25121 = ~n_19894 &  n_25120;
assign n_25122 = ~n_19891 &  n_25121;
assign n_25123 = ~n_19888 &  n_25122;
assign n_25124 = ~n_19885 &  n_25123;
assign n_25125 = ~n_19882 &  n_25124;
assign n_25126 = ~n_19879 &  n_25125;
assign n_25127 = ~n_19876 &  n_25126;
assign n_25128 = ~n_19873 &  n_25127;
assign n_25129 = ~n_19870 &  n_25128;
assign n_25130 = ~n_19867 &  n_25129;
assign n_25131 = ~n_19864 &  n_25130;
assign n_25132 = ~n_19861 &  n_25131;
assign n_25133 = ~n_19858 &  n_25132;
assign n_25134 = ~n_19855 &  n_25133;
assign n_25135 = ~n_19852 &  n_25134;
assign n_25136 = ~n_19849 &  n_25135;
assign n_25137 = ~n_19846 &  n_25136;
assign n_25138 = ~n_19843 &  n_25137;
assign n_25139 = ~n_19840 &  n_25138;
assign n_25140 = ~n_19837 &  n_25139;
assign n_25141 = ~n_19834 &  n_25140;
assign n_25142 = ~n_19831 &  n_25141;
assign n_25143 = ~n_19828 &  n_25142;
assign n_25144 = ~n_19825 &  n_25143;
assign n_25145 = ~n_19822 &  n_25144;
assign n_25146 = ~n_19819 &  n_25145;
assign n_25147 = ~n_19816 &  n_25146;
assign n_25148 = ~n_19813 &  n_25147;
assign n_25149 = ~n_19810 &  n_25148;
assign n_25150 = ~n_19807 &  n_25149;
assign n_25151 = ~n_19804 &  n_25150;
assign n_25152 = ~n_19801 &  n_25151;
assign n_25153 = ~n_19798 &  n_25152;
assign n_25154 = ~n_19795 &  n_25153;
assign n_25155 = ~n_19792 &  n_25154;
assign n_25156 = ~n_19789 &  n_25155;
assign n_25157 = ~n_19786 &  n_25156;
assign n_25158 = ~n_19783 &  n_25157;
assign n_25159 = ~n_19780 &  n_25158;
assign n_25160 = ~n_19777 &  n_25159;
assign n_25161 = ~n_19774 &  n_25160;
assign n_25162 = ~n_19771 &  n_25161;
assign n_25163 = ~n_19768 &  n_25162;
assign n_25164 = ~n_19765 &  n_25163;
assign n_25165 = ~n_19762 &  n_25164;
assign n_25166 = ~n_19759 &  n_25165;
assign n_25167 = ~n_19756 &  n_25166;
assign n_25168 = ~n_19753 &  n_25167;
assign n_25169 = ~n_19750 &  n_25168;
assign n_25170 = ~n_19747 &  n_25169;
assign n_25171 = ~n_19744 &  n_25170;
assign n_25172 = ~n_19741 &  n_25171;
assign n_25173 = ~n_19738 &  n_25172;
assign n_25174 = ~n_19735 &  n_25173;
assign n_25175 = ~n_19732 &  n_25174;
assign n_25176 = ~n_19729 &  n_25175;
assign n_25177 = ~n_19726 &  n_25176;
assign n_25178 = ~n_19723 &  n_25177;
assign n_25179 = ~n_19720 &  n_25178;
assign n_25180 = ~n_19717 &  n_25179;
assign n_25181 = ~n_19714 &  n_25180;
assign n_25182 = ~n_19711 &  n_25181;
assign n_25183 = ~n_19708 &  n_25182;
assign n_25184 = ~n_19705 &  n_25183;
assign n_25185 = ~n_19702 &  n_25184;
assign n_25186 = ~n_19699 &  n_25185;
assign n_25187 = ~n_19696 &  n_25186;
assign n_25188 = ~n_19693 &  n_25187;
assign n_25189 = ~n_19690 &  n_25188;
assign n_25190 = ~n_19687 &  n_25189;
assign n_25191 = ~n_19684 &  n_25190;
assign n_25192 = ~n_19681 &  n_25191;
assign n_25193 = ~n_19675 &  n_25192;
assign n_25194 = ~n_19669 &  n_25193;
assign n_25195 = ~n_19663 &  n_25194;
assign n_25196 = ~n_19657 &  n_25195;
assign n_25197 = ~n_19651 &  n_25196;
assign n_25198 = ~n_19645 &  n_25197;
assign n_25199 = ~n_19639 &  n_25198;
assign n_25200 = ~n_19624 &  n_25199;
assign n_25201 = ~n_19618 &  n_25200;
assign n_25202 = ~n_19612 &  n_25201;
assign n_25203 = ~n_19606 &  n_25202;
assign n_25204 = ~n_19600 &  n_25203;
assign n_25205 = ~n_19594 &  n_25204;
assign n_25206 = ~n_19588 &  n_25205;
assign n_25207 = ~n_19582 &  n_25206;
assign n_25208 = ~n_19567 &  n_25207;
assign n_25209 = ~n_19561 &  n_25208;
assign n_25210 = ~n_19555 &  n_25209;
assign n_25211 = ~n_19549 &  n_25210;
assign n_25212 = ~n_19543 &  n_25211;
assign n_25213 = ~n_19537 &  n_25212;
assign n_25214 = ~n_19531 &  n_25213;
assign n_25215 = ~n_19525 &  n_25214;
assign n_25216 = ~n_19510 &  n_25215;
assign n_25217 = ~n_19504 &  n_25216;
assign n_25218 = ~n_19498 &  n_25217;
assign n_25219 = ~n_19492 &  n_25218;
assign n_25220 = ~n_19486 &  n_25219;
assign n_25221 = ~n_19480 &  n_25220;
assign n_25222 = ~n_19474 &  n_25221;
assign n_25223 = ~n_19468 &  n_25222;
assign n_25224 = ~n_19453 &  n_25223;
assign n_25225 = ~n_19447 &  n_25224;
assign n_25226 = ~n_19441 &  n_25225;
assign n_25227 = ~n_19435 &  n_25226;
assign n_25228 = ~n_19429 &  n_25227;
assign n_25229 = ~n_19423 &  n_25228;
assign n_25230 = ~n_19417 &  n_25229;
assign n_25231 = ~n_19411 &  n_25230;
assign n_25232 = ~n_19396 &  n_25231;
assign n_25233 = ~n_19390 &  n_25232;
assign n_25234 = ~n_19384 &  n_25233;
assign n_25235 = ~n_19378 &  n_25234;
assign n_25236 = ~n_19372 &  n_25235;
assign n_25237 = ~n_19366 &  n_25236;
assign n_25238 = ~n_19360 &  n_25237;
assign n_25239 = ~n_19354 &  n_25238;
assign n_25240 = ~n_19339 &  n_25239;
assign n_25241 = ~n_19333 &  n_25240;
assign n_25242 = ~n_19327 &  n_25241;
assign n_25243 = ~n_19321 &  n_25242;
assign n_25244 = ~n_19315 &  n_25243;
assign n_25245 = ~n_19309 &  n_25244;
assign n_25246 = ~n_19303 &  n_25245;
assign n_25247 = ~n_19297 &  n_25246;
assign n_25248 = ~n_19282 &  n_25247;
assign n_25249 = ~n_19276 &  n_25248;
assign n_25250 = ~n_19270 &  n_25249;
assign n_25251 = ~n_19264 &  n_25250;
assign n_25252 = ~n_19258 &  n_25251;
assign n_25253 = ~n_19252 &  n_25252;
assign n_25254 = ~n_19246 &  n_25253;
assign n_25255 = ~n_19240 &  n_25254;
assign n_25256 = ~n_19225 &  n_25255;
assign n_25257 = ~n_19219 &  n_25256;
assign n_25258 = ~n_19213 &  n_25257;
assign n_25259 = ~n_19207 &  n_25258;
assign n_25260 = ~n_19201 &  n_25259;
assign n_25261 = ~n_19195 &  n_25260;
assign n_25262 = ~n_19189 &  n_25261;
assign n_25263 = ~n_19183 &  n_25262;
assign n_25264 = ~n_19168 &  n_25263;
assign n_25265 = ~n_19162 &  n_25264;
assign n_25266 = ~n_19156 &  n_25265;
assign n_25267 = ~n_19150 &  n_25266;
assign n_25268 = ~n_19144 &  n_25267;
assign n_25269 = ~n_19138 &  n_25268;
assign n_25270 = ~n_19132 &  n_25269;
assign n_25271 = ~n_19126 &  n_25270;
assign n_25272 = ~n_19111 &  n_25271;
assign n_25273 = ~n_19105 &  n_25272;
assign n_25274 = ~n_19099 &  n_25273;
assign n_25275 = ~n_19093 &  n_25274;
assign n_25276 = ~n_19087 &  n_25275;
assign n_25277 = ~n_19081 &  n_25276;
assign n_25278 = ~n_19075 &  n_25277;
assign n_25279 = ~n_19069 &  n_25278;
assign n_25280 = ~n_19054 &  n_25279;
assign n_25281 = ~n_19048 &  n_25280;
assign n_25282 = ~n_19042 &  n_25281;
assign n_25283 = ~n_19036 &  n_25282;
assign n_25284 = ~n_19030 &  n_25283;
assign n_25285 = ~n_19024 &  n_25284;
assign n_25286 = ~n_19018 &  n_25285;
assign n_25287 = ~n_19012 &  n_25286;
assign n_25288 = ~n_18997 &  n_25287;
assign n_25289 = ~n_18991 &  n_25288;
assign n_25290 = ~n_18985 &  n_25289;
assign n_25291 = ~n_18979 &  n_25290;
assign n_25292 = ~n_18973 &  n_25291;
assign n_25293 = ~n_18967 &  n_25292;
assign n_25294 = ~n_18961 &  n_25293;
assign n_25295 = ~n_18955 &  n_25294;
assign n_25296 = ~n_18940 &  n_25295;
assign n_25297 = ~n_18934 &  n_25296;
assign n_25298 = ~n_18928 &  n_25297;
assign n_25299 = ~n_18922 &  n_25298;
assign n_25300 = ~n_18916 &  n_25299;
assign n_25301 = ~n_18910 &  n_25300;
assign n_25302 = ~n_18904 &  n_25301;
assign n_25303 = ~n_18898 &  n_25302;
assign n_25304 = ~n_18883 &  n_25303;
assign n_25305 = ~n_18877 &  n_25304;
assign n_25306 = ~n_18871 &  n_25305;
assign n_25307 = ~n_18865 &  n_25306;
assign n_25308 = ~n_18859 &  n_25307;
assign n_25309 = ~n_18853 &  n_25308;
assign n_25310 = ~n_18847 &  n_25309;
assign n_25311 = ~n_18841 &  n_25310;
assign n_25312 = ~n_18826 &  n_25311;
assign n_25313 = ~n_18820 &  n_25312;
assign n_25314 = ~n_18814 &  n_25313;
assign n_25315 = ~n_18808 &  n_25314;
assign n_25316 = ~n_18802 &  n_25315;
assign n_25317 = ~n_18796 &  n_25316;
assign n_25318 = ~n_18790 &  n_25317;
assign n_25319 = ~n_18784 &  n_25318;
assign n_25320 = ~n_18769 &  n_25319;
assign n_25321 = ~n_18763 &  n_25320;
assign n_25322 = ~n_18757 &  n_25321;
assign n_25323 = ~n_18751 &  n_25322;
assign n_25324 = ~n_18745 &  n_25323;
assign n_25325 = ~n_18739 &  n_25324;
assign n_25326 = ~n_18733 &  n_25325;
assign n_25327 = ~n_18727 &  n_25326;
assign n_25328 = ~n_18712 &  n_25327;
assign n_25329 = ~n_18706 &  n_25328;
assign n_25330 = ~n_18700 &  n_25329;
assign n_25331 = ~n_18694 &  n_25330;
assign n_25332 = ~n_18688 &  n_25331;
assign n_25333 = ~n_18682 &  n_25332;
assign n_25334 = ~n_18676 &  n_25333;
assign n_25335 = ~n_18670 &  n_25334;
assign n_25336 = ~n_18655 &  n_25335;
assign n_25337 = ~n_18649 &  n_25336;
assign n_25338 = ~n_18643 &  n_25337;
assign n_25339 = ~n_18637 &  n_25338;
assign n_25340 = ~n_18631 &  n_25339;
assign n_25341 = ~n_18625 &  n_25340;
assign n_25342 = ~n_18619 &  n_25341;
assign n_25343 = ~n_18613 &  n_25342;
assign n_25344 = ~n_18598 &  n_25343;
assign n_25345 = ~n_18592 &  n_25344;
assign n_25346 = ~n_18586 &  n_25345;
assign n_25347 = ~n_18580 &  n_25346;
assign n_25348 = ~n_18574 &  n_25347;
assign n_25349 = ~n_18568 &  n_25348;
assign n_25350 = ~n_18562 &  n_25349;
assign n_25351 = ~n_18556 &  n_25350;
assign n_25352 = ~n_18541 &  n_25351;
assign n_25353 = ~n_18535 &  n_25352;
assign n_25354 = ~n_18529 &  n_25353;
assign n_25355 = ~n_18523 &  n_25354;
assign n_25356 = ~n_18517 &  n_25355;
assign n_25357 = ~n_18511 &  n_25356;
assign n_25358 = ~n_18505 &  n_25357;
assign n_25359 = ~n_18499 &  n_25358;
assign n_25360 = ~n_18484 &  n_25359;
assign n_25361 = ~n_18478 &  n_25360;
assign n_25362 = ~n_18472 &  n_25361;
assign n_25363 = ~n_18466 &  n_25362;
assign n_25364 = ~n_18460 &  n_25363;
assign n_25365 = ~n_18454 &  n_25364;
assign n_25366 = ~n_18448 &  n_25365;
assign n_25367 = ~n_18442 &  n_25366;
assign n_25368 = ~n_18427 &  n_25367;
assign n_25369 = ~n_18421 &  n_25368;
assign n_25370 = ~n_18415 &  n_25369;
assign n_25371 = ~n_18409 &  n_25370;
assign n_25372 = ~n_18403 &  n_25371;
assign n_25373 = ~n_18397 &  n_25372;
assign n_25374 = ~n_18391 &  n_25373;
assign n_25375 = ~n_18385 &  n_25374;
assign n_25376 = ~n_18370 &  n_25375;
assign n_25377 = ~n_18364 &  n_25376;
assign n_25378 = ~n_18358 &  n_25377;
assign n_25379 = ~n_18352 &  n_25378;
assign n_25380 = ~n_18346 &  n_25379;
assign n_25381 = ~n_18340 &  n_25380;
assign n_25382 = ~n_18334 &  n_25381;
assign n_25383 = ~n_18328 &  n_25382;
assign n_25384 = ~n_18313 &  n_25383;
assign n_25385 = ~n_18307 &  n_25384;
assign n_25386 = ~n_18301 &  n_25385;
assign n_25387 = ~n_18295 &  n_25386;
assign n_25388 = ~n_18289 &  n_25387;
assign n_25389 = ~n_18283 &  n_25388;
assign n_25390 = ~n_18277 &  n_25389;
assign n_25391 = ~n_18271 &  n_25390;
assign n_25392 = ~n_18256 &  n_25391;
assign n_25393 = ~n_18250 &  n_25392;
assign n_25394 = ~n_18244 &  n_25393;
assign n_25395 = ~n_18238 &  n_25394;
assign n_25396 = ~n_18232 &  n_25395;
assign n_25397 = ~n_18226 &  n_25396;
assign n_25398 = ~n_18220 &  n_25397;
assign n_25399 = ~n_18214 &  n_25398;
assign n_25400 = ~n_18199 &  n_25399;
assign n_25401 = ~n_18193 &  n_25400;
assign n_25402 = ~n_18187 &  n_25401;
assign n_25403 = ~n_18181 &  n_25402;
assign n_25404 = ~n_18175 &  n_25403;
assign n_25405 = ~n_18169 &  n_25404;
assign n_25406 = ~n_18163 &  n_25405;
assign n_25407 = ~n_18157 &  n_25406;
assign n_25408 = ~n_18142 &  n_25407;
assign n_25409 = ~n_18136 &  n_25408;
assign n_25410 = ~n_18130 &  n_25409;
assign n_25411 = ~n_18124 &  n_25410;
assign n_25412 = ~n_18118 &  n_25411;
assign n_25413 = ~n_18112 &  n_25412;
assign n_25414 = ~n_18106 &  n_25413;
assign n_25415 = ~n_18100 &  n_25414;
assign n_25416 = ~n_18085 &  n_25415;
assign n_25417 = ~n_18079 &  n_25416;
assign n_25418 = ~n_18073 &  n_25417;
assign n_25419 = ~n_18067 &  n_25418;
assign n_25420 = ~n_18061 &  n_25419;
assign n_25421 = ~n_18055 &  n_25420;
assign n_25422 = ~n_18049 &  n_25421;
assign n_25423 = ~n_18043 &  n_25422;
assign n_25424 = ~n_18028 &  n_25423;
assign n_25425 = ~n_18022 &  n_25424;
assign n_25426 = ~n_18016 &  n_25425;
assign n_25427 = ~n_18010 &  n_25426;
assign n_25428 = ~n_18004 &  n_25427;
assign n_25429 = ~n_17998 &  n_25428;
assign n_25430 = ~n_17992 &  n_25429;
assign n_25431 = ~n_17986 &  n_25430;
assign n_25432 = ~n_17971 &  n_25431;
assign n_25433 = ~n_17965 &  n_25432;
assign n_25434 = ~n_17959 &  n_25433;
assign n_25435 = ~n_17953 &  n_25434;
assign n_25436 = ~n_17947 &  n_25435;
assign n_25437 = ~n_17941 &  n_25436;
assign n_25438 = ~n_17935 &  n_25437;
assign n_25439 = ~n_17929 &  n_25438;
assign n_25440 = ~n_17914 &  n_25439;
assign n_25441 = ~n_17908 &  n_25440;
assign n_25442 = ~n_17902 &  n_25441;
assign n_25443 = ~n_17896 &  n_25442;
assign n_25444 = ~n_17890 &  n_25443;
assign n_25445 = ~n_17884 &  n_25444;
assign n_25446 = ~n_17878 &  n_25445;
assign n_25447 = ~n_17872 &  n_25446;
assign n_25448 = ~n_17857 &  n_25447;
assign n_25449 = ~n_17850 &  n_25448;
assign n_25450 = ~n_17843 &  n_25449;
assign n_25451 = ~n_17836 &  n_25450;
assign n_25452 = ~n_17829 &  n_25451;
assign n_25453 = ~n_17821 &  n_25452;
assign n_25454 = ~n_17813 &  n_25453;
assign n_25455 = ~n_17804 &  n_25454;
assign n_25456 = ~n_17786 &  n_25455;
assign n_25457 = ~n_17784 &  n_25456;
assign n_25458 = ~n_17782 &  n_25457;
assign n_25459 = ~n_17779 &  n_25458;
assign n_25460 = ~n_17776 &  n_25459;
assign n_25461 = ~n_17774 &  n_25460;
assign n_25462 = ~n_17771 &  n_25461;
assign n_25463 = ~n_17768 &  n_25462;
assign n_25464 = ~n_17762 &  n_25463;
assign n_25465 = ~n_17756 &  n_25464;
assign n_25466 = ~n_17750 &  n_25465;
assign n_25467 = ~n_17744 &  n_25466;
assign n_25468 = ~n_17738 &  n_25467;
assign n_25469 = ~n_17732 &  n_25468;
assign n_25470 = ~n_17726 &  n_25469;
assign n_25471 = ~n_17720 &  n_25470;
assign n_25472 = ~n_17716 &  n_25471;
assign n_25473 = ~n_17710 &  n_25472;
assign n_25474 = ~n_17704 &  n_25473;
assign n_25475 = ~n_17698 &  n_25474;
assign n_25476 = ~n_17686 &  n_25475;
assign n_25477 = ~n_17683 &  n_25476;
assign n_25478 = ~n_17679 &  n_25477;
assign n_25479 = ~n_17675 &  n_25478;
assign n_25480 = ~n_17668 &  n_25479;
assign n_25481 = ~n_17663 &  n_25480;
assign n_25482 = ~n_17657 &  n_25481;
assign n_25483 = ~n_17652 &  n_25482;
assign n_25484 = ~n_17647 &  n_25483;
assign n_25485 = ~n_17642 &  n_25484;
assign n_25486 = ~n_17639 &  n_25485;
assign n_25487 = ~n_17636 &  n_25486;
assign n_25488 = ~n_17632 &  n_25487;
assign n_25489 = ~n_17626 &  n_25488;
assign n_25490 = ~n_17623 &  n_25489;
assign n_25491 = ~n_17620 &  n_25490;
assign n_25492 = ~n_17615 &  n_25491;
assign n_25493 = ~n_17610 &  n_25492;
assign n_25494 = ~n_17605 &  n_25493;
assign n_25495 = ~n_17600 &  n_25494;
assign n_25496 = ~n_17595 &  n_25495;
assign n_25497 = ~n_17590 &  n_25496;
assign n_25498 = ~n_17585 &  n_25497;
assign n_25499 = ~n_17580 &  n_25498;
assign n_25500 = ~n_17575 &  n_25499;
assign n_25501 = ~n_17570 &  n_25500;
assign n_25502 = ~n_17565 &  n_25501;
assign n_25503 = ~n_17560 &  n_25502;
assign n_25504 = ~n_17555 &  n_25503;
assign n_25505 = ~n_17550 &  n_25504;
assign n_25506 = ~n_17545 &  n_25505;
assign n_25507 = ~n_17540 &  n_25506;
assign n_25508 = ~n_17535 &  n_25507;
assign n_25509 = ~n_17530 &  n_25508;
assign n_25510 = ~n_17525 &  n_25509;
assign n_25511 = ~n_17520 &  n_25510;
assign n_25512 = ~n_17515 &  n_25511;
assign n_25513 = ~n_17510 &  n_25512;
assign n_25514 = ~n_17505 &  n_25513;
assign n_25515 = ~n_17500 &  n_25514;
assign n_25516 = ~n_17495 &  n_25515;
assign n_25517 = ~n_17490 &  n_25516;
assign n_25518 = ~n_17485 &  n_25517;
assign n_25519 = ~n_17480 &  n_25518;
assign n_25520 = ~n_17475 &  n_25519;
assign n_25521 = ~n_17470 &  n_25520;
assign n_25522 = ~n_17467 &  n_25521;
assign n_25523 = ~n_17464 &  n_25522;
assign n_25524 = ~n_17461 &  n_25523;
assign n_25525 = ~n_17458 &  n_25524;
assign n_25526 = ~n_17455 &  n_25525;
assign n_25527 = ~n_17452 &  n_25526;
assign n_25528 = ~n_17449 &  n_25527;
assign n_25529 = ~n_17446 &  n_25528;
assign n_25530 = ~n_17443 &  n_25529;
assign n_25531 = ~n_17440 &  n_25530;
assign n_25532 = ~n_17437 &  n_25531;
assign n_25533 = ~n_17434 &  n_25532;
assign n_25534 = ~n_17431 &  n_25533;
assign n_25535 = ~n_17428 &  n_25534;
assign n_25536 = ~n_17425 &  n_25535;
assign n_25537 = ~n_17422 &  n_25536;
assign n_25538 = ~n_17419 &  n_25537;
assign n_25539 = ~n_17416 &  n_25538;
assign n_25540 = ~n_17413 &  n_25539;
assign n_25541 = ~n_17410 &  n_25540;
assign n_25542 = ~n_17407 &  n_25541;
assign n_25543 = ~n_17404 &  n_25542;
assign n_25544 = ~n_17401 &  n_25543;
assign n_25545 = ~n_17398 &  n_25544;
assign n_25546 = ~n_17395 &  n_25545;
assign n_25547 = ~n_17392 &  n_25546;
assign n_25548 = ~n_17389 &  n_25547;
assign n_25549 = ~n_17384 &  n_25548;
assign n_25550 = ~n_17347 &  n_25549;
assign n_25551 = ~n_17344 &  n_25550;
assign n_25552 = ~n_17341 &  n_25551;
assign n_25553 = ~n_17337 &  n_25552;
assign n_25554 = ~n_17331 &  n_25553;
assign n_25555 = ~n_17324 &  n_25554;
assign n_25556 = ~n_17317 &  n_25555;
assign n_25557 = ~n_17310 &  n_25556;
assign n_25558 = ~n_17303 &  n_25557;
assign n_25559 = ~n_17296 &  n_25558;
assign n_25560 = ~n_17289 &  n_25559;
assign n_25561 = ~n_17282 &  n_25560;
assign n_25562 = ~n_17275 &  n_25561;
assign n_25563 = ~n_17268 &  n_25562;
assign n_25564 = ~n_17261 &  n_25563;
assign n_25565 = ~n_17254 &  n_25564;
assign n_25566 = ~n_17247 &  n_25565;
assign n_25567 = ~n_17240 &  n_25566;
assign n_25568 = ~n_17233 &  n_25567;
assign n_25569 = ~n_17226 &  n_25568;
assign n_25570 = ~n_17219 &  n_25569;
assign n_25571 = ~n_17212 &  n_25570;
assign n_25572 = ~n_17205 &  n_25571;
assign n_25573 = ~n_17198 &  n_25572;
assign n_25574 = ~n_17191 &  n_25573;
assign n_25575 = ~n_17184 &  n_25574;
assign n_25576 = ~n_17177 &  n_25575;
assign n_25577 = ~n_17170 &  n_25576;
assign n_25578 = ~n_17163 &  n_25577;
assign n_25579 = ~n_17156 &  n_25578;
assign n_25580 = ~n_17149 &  n_25579;
assign n_25581 = ~n_17142 &  n_25580;
assign n_25582 = ~n_17134 &  n_25581;
assign n_25583 = ~n_17127 &  n_25582;
assign n_25584 = ~n_17120 &  n_25583;
assign n_25585 = ~n_17117 &  n_25584;
assign n_25586 = ~n_17107 &  n_25585;
assign n_25587 = ~n_17104 &  n_25586;
assign n_25588 = ~n_17099 &  n_25587;
assign n_25589 = ~n_17092 &  n_25588;
assign n_25590 = ~n_17082 &  n_25589;
assign n_25591 = ~n_17077 &  n_25590;
assign n_25592 = ~n_17056 &  n_25591;
assign n_25593 = ~n_17050 &  n_25592;
assign n_25594 = ~n_17044 &  n_25593;
assign n_25595 = ~n_17038 &  n_25594;
assign n_25596 = ~n_17032 &  n_25595;
assign n_25597 = ~n_17026 &  n_25596;
assign n_25598 = ~n_17020 &  n_25597;
assign n_25599 = ~n_17014 &  n_25598;
assign n_25600 = ~n_17008 &  n_25599;
assign n_25601 = ~n_17002 &  n_25600;
assign n_25602 = ~n_16996 &  n_25601;
assign n_25603 = ~n_16990 &  n_25602;
assign n_25604 = ~n_16984 &  n_25603;
assign n_25605 = ~n_16978 &  n_25604;
assign n_25606 = ~n_16972 &  n_25605;
assign n_25607 = ~n_16966 &  n_25606;
assign n_25608 = ~n_16960 &  n_25607;
assign n_25609 = ~n_16957 &  n_25608;
assign n_25610 = ~n_16951 &  n_25609;
assign n_25611 = ~n_16945 &  n_25610;
assign n_25612 = ~n_16939 &  n_25611;
assign n_25613 = ~n_16933 &  n_25612;
assign n_25614 = ~n_16927 &  n_25613;
assign n_25615 = ~n_16921 &  n_25614;
assign n_25616 = ~n_16915 &  n_25615;
assign n_25617 = ~n_16909 &  n_25616;
assign n_25618 = ~n_16903 &  n_25617;
assign n_25619 = ~n_16897 &  n_25618;
assign n_25620 = ~n_16891 &  n_25619;
assign n_25621 = ~n_16885 &  n_25620;
assign n_25622 = ~n_16879 &  n_25621;
assign n_25623 = ~n_16873 &  n_25622;
assign n_25624 = ~n_16867 &  n_25623;
assign n_25625 = ~n_16861 &  n_25624;
assign n_25626 = ~n_16855 &  n_25625;
assign n_25627 = ~n_16849 &  n_25626;
assign n_25628 = ~n_16843 &  n_25627;
assign n_25629 = ~n_16837 &  n_25628;
assign n_25630 = ~n_16831 &  n_25629;
assign n_25631 = ~n_16825 &  n_25630;
assign n_25632 = ~n_16819 &  n_25631;
assign n_25633 = ~n_16813 &  n_25632;
assign n_25634 = ~n_16807 &  n_25633;
assign n_25635 = ~n_16801 &  n_25634;
assign n_25636 = ~n_16795 &  n_25635;
assign n_25637 = ~n_16789 &  n_25636;
assign n_25638 = ~n_16783 &  n_25637;
assign n_25639 = ~n_16777 &  n_25638;
assign n_25640 = ~n_16771 &  n_25639;
assign n_25641 = ~n_16765 &  n_25640;
assign n_25642 = ~n_16758 &  n_25641;
assign n_25643 = ~n_16755 &  n_25642;
assign n_25644 = ~n_16749 &  n_25643;
assign n_25645 = ~n_16743 &  n_25644;
assign n_25646 = ~n_16737 &  n_25645;
assign n_25647 = ~n_16731 &  n_25646;
assign n_25648 = ~n_16725 &  n_25647;
assign n_25649 = ~n_16719 &  n_25648;
assign n_25650 = ~n_16713 &  n_25649;
assign n_25651 = ~n_16707 &  n_25650;
assign n_25652 = ~n_16701 &  n_25651;
assign n_25653 = ~n_16695 &  n_25652;
assign n_25654 = ~n_16689 &  n_25653;
assign n_25655 = ~n_16683 &  n_25654;
assign n_25656 = ~n_16677 &  n_25655;
assign n_25657 = ~n_16671 &  n_25656;
assign n_25658 = ~n_16665 &  n_25657;
assign n_25659 = ~n_16659 &  n_25658;
assign n_25660 = ~n_16653 &  n_25659;
assign n_25661 = ~n_16647 &  n_25660;
assign n_25662 = ~n_16641 &  n_25661;
assign n_25663 = ~n_16635 &  n_25662;
assign n_25664 = ~n_16629 &  n_25663;
assign n_25665 = ~n_16623 &  n_25664;
assign n_25666 = ~n_16617 &  n_25665;
assign n_25667 = ~n_16611 &  n_25666;
assign n_25668 = ~n_16605 &  n_25667;
assign n_25669 = ~n_16599 &  n_25668;
assign n_25670 = ~n_16593 &  n_25669;
assign n_25671 = ~n_16587 &  n_25670;
assign n_25672 = ~n_16581 &  n_25671;
assign n_25673 = ~n_16575 &  n_25672;
assign n_25674 = ~n_16569 &  n_25673;
assign n_25675 = ~n_16563 &  n_25674;
assign n_25676 = ~n_16557 &  n_25675;
assign n_25677 = ~n_16551 &  n_25676;
assign n_25678 = ~n_16545 &  n_25677;
assign n_25679 = ~n_16539 &  n_25678;
assign n_25680 = ~n_16533 &  n_25679;
assign n_25681 = ~n_16527 &  n_25680;
assign n_25682 = ~n_16521 &  n_25681;
assign n_25683 = ~n_16515 &  n_25682;
assign n_25684 = ~n_16509 &  n_25683;
assign n_25685 = ~n_16503 &  n_25684;
assign n_25686 = ~n_16497 &  n_25685;
assign n_25687 = ~n_16491 &  n_25686;
assign n_25688 = ~n_16485 &  n_25687;
assign n_25689 = ~n_16479 &  n_25688;
assign n_25690 = ~n_16473 &  n_25689;
assign n_25691 = ~n_16467 &  n_25690;
assign n_25692 = ~n_16461 &  n_25691;
assign n_25693 = ~n_16455 &  n_25692;
assign n_25694 = ~n_16449 &  n_25693;
assign n_25695 = ~n_16443 &  n_25694;
assign n_25696 = ~n_16437 &  n_25695;
assign n_25697 = ~n_16431 &  n_25696;
assign n_25698 = ~n_16425 &  n_25697;
assign n_25699 = ~n_16419 &  n_25698;
assign n_25700 = ~n_16413 &  n_25699;
assign n_25701 = ~n_16407 &  n_25700;
assign n_25702 = ~n_16401 &  n_25701;
assign n_25703 = ~n_16395 &  n_25702;
assign n_25704 = ~n_16389 &  n_25703;
assign n_25705 = ~n_16383 &  n_25704;
assign n_25706 = ~n_16377 &  n_25705;
assign n_25707 = ~n_16371 &  n_25706;
assign n_25708 = ~n_16365 &  n_25707;
assign n_25709 = ~n_16361 &  n_25708;
assign n_25710 = ~n_16357 &  n_25709;
assign n_25711 = ~n_16352 &  n_25710;
assign n_25712 = ~n_16332 &  n_25711;
assign n_25713 = ~n_16304 &  n_25712;
assign n_25714 = ~n_16293 &  n_25713;
assign n_25715 = ~n_16262 &  n_25714;
assign n_25716 = ~n_16259 &  n_25715;
assign n_25717 = ~n_16243 &  n_25716;
assign n_25718 = ~n_16218 &  n_25717;
assign n_25719 = ~n_16150 &  n_25718;
assign n_25720 = ~n_16123 &  n_25719;
assign n_25721 = ~n_16120 &  n_25720;
assign n_25722 = ~n_16117 &  n_25721;
assign n_25723 = ~n_16114 &  n_25722;
assign n_25724 = ~n_16109 &  n_25723;
assign n_25725 = ~n_16106 &  n_25724;
assign n_25726 = ~n_16098 &  n_25725;
assign n_25727 = ~n_16094 &  n_25726;
assign n_25728 = ~n_16089 &  n_25727;
assign n_25729 = ~n_16084 &  n_25728;
assign n_25730 = ~n_16078 &  n_25729;
assign n_25731 = ~n_16072 &  n_25730;
assign n_25732 = ~n_16066 &  n_25731;
assign n_25733 = ~n_16060 &  n_25732;
assign n_25734 = ~n_16054 &  n_25733;
assign n_25735 = ~n_16048 &  n_25734;
assign n_25736 = ~n_16045 &  n_25735;
assign n_25737 = ~n_16042 &  n_25736;
assign n_25738 = ~n_16039 &  n_25737;
assign n_25739 = ~n_16036 &  n_25738;
assign n_25740 = ~n_16033 &  n_25739;
assign n_25741 = ~n_16029 &  n_25740;
assign n_25742 = ~n_16019 &  n_25741;
assign n_25743 = ~n_16013 &  n_25742;
assign n_25744 = ~n_16010 &  n_25743;
assign n_25745 = ~n_16007 &  n_25744;
assign n_25746 = ~n_16004 &  n_25745;
assign n_25747 = ~n_16001 &  n_25746;
assign n_25748 = ~n_15998 &  n_25747;
assign n_25749 = ~n_15995 &  n_25748;
assign n_25750 = ~n_15992 &  n_25749;
assign n_25751 = ~n_15989 &  n_25750;
assign n_25752 = ~n_15986 &  n_25751;
assign n_25753 = ~n_15983 &  n_25752;
assign n_25754 = ~n_15980 &  n_25753;
assign n_25755 = ~n_15962 &  n_25754;
assign n_25756 = ~n_15954 &  n_25755;
assign n_25757 = ~n_15940 &  n_25756;
assign n_25758 = ~n_15936 &  n_25757;
assign n_25759 = ~n_15927 &  n_25758;
assign n_25760 = ~n_15909 &  n_25759;
assign n_25761 = ~n_15901 &  n_25760;
assign n_25762 = ~n_15888 &  n_25761;
assign n_25763 = ~n_15882 &  n_25762;
assign n_25764 = ~n_15876 &  n_25763;
assign n_25765 = ~n_15870 &  n_25764;
assign n_25766 = ~n_15864 &  n_25765;
assign n_25767 = ~n_15858 &  n_25766;
assign n_25768 = ~n_15852 &  n_25767;
assign n_25769 = ~n_15846 &  n_25768;
assign n_25770 = ~n_15840 &  n_25769;
assign n_25771 = ~n_15834 &  n_25770;
assign n_25772 = ~n_15828 &  n_25771;
assign n_25773 = ~n_15822 &  n_25772;
assign n_25774 = ~n_15816 &  n_25773;
assign n_25775 = ~n_15810 &  n_25774;
assign n_25776 = ~n_15804 &  n_25775;
assign n_25777 = ~n_15798 &  n_25776;
assign n_25778 = ~n_15792 &  n_25777;
assign n_25779 = ~n_15786 &  n_25778;
assign n_25780 = ~n_15780 &  n_25779;
assign n_25781 = ~n_15774 &  n_25780;
assign n_25782 = ~n_15768 &  n_25781;
assign n_25783 = ~n_15762 &  n_25782;
assign n_25784 = ~n_15756 &  n_25783;
assign n_25785 = ~n_15750 &  n_25784;
assign n_25786 = ~n_15744 &  n_25785;
assign n_25787 = ~n_15738 &  n_25786;
assign n_25788 = ~n_15732 &  n_25787;
assign n_25789 = ~n_15726 &  n_25788;
assign n_25790 = ~n_15720 &  n_25789;
assign n_25791 = ~n_15714 &  n_25790;
assign n_25792 = ~n_15708 &  n_25791;
assign n_25793 = ~n_15702 &  n_25792;
assign n_25794 = ~n_15696 &  n_25793;
assign n_25795 = ~n_15690 &  n_25794;
assign n_25796 = ~n_15684 &  n_25795;
assign n_25797 = ~n_15678 &  n_25796;
assign n_25798 = ~n_15672 &  n_25797;
assign n_25799 = ~n_15666 &  n_25798;
assign n_25800 = ~n_15660 &  n_25799;
assign n_25801 = ~n_15654 &  n_25800;
assign n_25802 = ~n_15648 &  n_25801;
assign n_25803 = ~n_15642 &  n_25802;
assign n_25804 = ~n_15637 &  n_25803;
assign n_25805 = ~n_15631 &  n_25804;
assign n_25806 = ~n_15625 &  n_25805;
assign n_25807 = ~n_15619 &  n_25806;
assign n_25808 = ~n_15613 &  n_25807;
assign n_25809 = ~n_15607 &  n_25808;
assign n_25810 = ~n_15601 &  n_25809;
assign n_25811 = ~n_15595 &  n_25810;
assign n_25812 = ~n_15589 &  n_25811;
assign n_25813 = ~n_15583 &  n_25812;
assign n_25814 = ~n_15577 &  n_25813;
assign n_25815 = ~n_15571 &  n_25814;
assign n_25816 = ~n_15565 &  n_25815;
assign n_25817 = ~n_15559 &  n_25816;
assign n_25818 = ~n_15553 &  n_25817;
assign n_25819 = ~n_15547 &  n_25818;
assign n_25820 = ~n_15541 &  n_25819;
assign n_25821 = ~n_15535 &  n_25820;
assign n_25822 = ~n_15529 &  n_25821;
assign n_25823 = ~n_15523 &  n_25822;
assign n_25824 = ~n_15517 &  n_25823;
assign n_25825 = ~n_15511 &  n_25824;
assign n_25826 = ~n_15505 &  n_25825;
assign n_25827 = ~n_15499 &  n_25826;
assign n_25828 = ~n_15493 &  n_25827;
assign n_25829 = ~n_15487 &  n_25828;
assign n_25830 = ~n_15481 &  n_25829;
assign n_25831 = ~n_15475 &  n_25830;
assign n_25832 = ~n_15469 &  n_25831;
assign n_25833 = ~n_15463 &  n_25832;
assign n_25834 = ~n_15457 &  n_25833;
assign n_25835 = ~n_15451 &  n_25834;
assign n_25836 = ~n_15445 &  n_25835;
assign n_25837 = ~n_15439 &  n_25836;
assign n_25838 = ~n_15433 &  n_25837;
assign n_25839 = ~n_15427 &  n_25838;
assign n_25840 = ~n_15421 &  n_25839;
assign n_25841 = ~n_15415 &  n_25840;
assign n_25842 = ~n_15409 &  n_25841;
assign n_25843 = ~n_15403 &  n_25842;
assign n_25844 = ~n_15396 &  n_25843;
assign n_25845 = ~n_15390 &  n_25844;
assign n_25846 = ~n_15384 &  n_25845;
assign n_25847 = ~n_15378 &  n_25846;
assign n_25848 = ~n_15372 &  n_25847;
assign n_25849 = ~n_15366 &  n_25848;
assign n_25850 = ~n_15360 &  n_25849;
assign n_25851 = ~n_15354 &  n_25850;
assign n_25852 = ~n_15347 &  n_25851;
assign n_25853 = ~n_15341 &  n_25852;
assign n_25854 = ~n_15335 &  n_25853;
assign n_25855 = ~n_15329 &  n_25854;
assign n_25856 = ~n_15323 &  n_25855;
assign n_25857 = ~n_15317 &  n_25856;
assign n_25858 = ~n_15311 &  n_25857;
assign n_25859 = ~n_15305 &  n_25858;
assign n_25860 = ~n_15299 &  n_25859;
assign n_25861 = ~n_15293 &  n_25860;
assign n_25862 = ~n_15286 &  n_25861;
assign n_25863 = ~n_15280 &  n_25862;
assign n_25864 = ~n_15274 &  n_25863;
assign n_25865 = ~n_15268 &  n_25864;
assign n_25866 = ~n_15262 &  n_25865;
assign n_25867 = ~n_15256 &  n_25866;
assign n_25868 = ~n_15250 &  n_25867;
assign n_25869 = ~n_15244 &  n_25868;
assign n_25870 = ~n_15238 &  n_25869;
assign n_25871 = ~n_15231 &  n_25870;
assign n_25872 = ~n_15225 &  n_25871;
assign n_25873 = ~n_15219 &  n_25872;
assign n_25874 = ~n_15213 &  n_25873;
assign n_25875 = ~n_15207 &  n_25874;
assign n_25876 = ~n_15201 &  n_25875;
assign n_25877 = ~n_15195 &  n_25876;
assign n_25878 = ~n_15189 &  n_25877;
assign n_25879 = ~n_15183 &  n_25878;
assign n_25880 = ~n_15177 &  n_25879;
assign n_25881 = ~n_15171 &  n_25880;
assign n_25882 = ~n_15165 &  n_25881;
assign n_25883 = ~n_15159 &  n_25882;
assign n_25884 = ~n_15153 &  n_25883;
assign n_25885 = ~n_15147 &  n_25884;
assign n_25886 = ~n_15141 &  n_25885;
assign n_25887 = ~n_15135 &  n_25886;
assign n_25888 = ~n_15129 &  n_25887;
assign n_25889 = ~n_15122 &  n_25888;
assign n_25890 = ~n_15116 &  n_25889;
assign n_25891 = ~n_15110 &  n_25890;
assign n_25892 = ~n_15104 &  n_25891;
assign n_25893 = ~n_15098 &  n_25892;
assign n_25894 = ~n_15092 &  n_25893;
assign n_25895 = ~n_15086 &  n_25894;
assign n_25896 = ~n_15080 &  n_25895;
assign n_25897 = ~n_15073 &  n_25896;
assign n_25898 = ~n_15067 &  n_25897;
assign n_25899 = ~n_15061 &  n_25898;
assign n_25900 = ~n_15055 &  n_25899;
assign n_25901 = ~n_15049 &  n_25900;
assign n_25902 = ~n_15043 &  n_25901;
assign n_25903 = ~n_15037 &  n_25902;
assign n_25904 = ~n_15031 &  n_25903;
assign n_25905 = ~n_15024 &  n_25904;
assign n_25906 = ~n_15018 &  n_25905;
assign n_25907 = ~n_15012 &  n_25906;
assign n_25908 = ~n_15006 &  n_25907;
assign n_25909 = ~n_15000 &  n_25908;
assign n_25910 = ~n_14994 &  n_25909;
assign n_25911 = ~n_14988 &  n_25910;
assign n_25912 = ~n_14982 &  n_25911;
assign n_25913 = ~n_14975 &  n_25912;
assign n_25914 = ~n_14969 &  n_25913;
assign n_25915 = ~n_14963 &  n_25914;
assign n_25916 = ~n_14957 &  n_25915;
assign n_25917 = ~n_14951 &  n_25916;
assign n_25918 = ~n_14945 &  n_25917;
assign n_25919 = ~n_14939 &  n_25918;
assign n_25920 = ~n_14933 &  n_25919;
assign n_25921 = ~n_14926 &  n_25920;
assign n_25922 = ~n_14920 &  n_25921;
assign n_25923 = ~n_14914 &  n_25922;
assign n_25924 = ~n_14908 &  n_25923;
assign n_25925 = ~n_14902 &  n_25924;
assign n_25926 = ~n_14896 &  n_25925;
assign n_25927 = ~n_14890 &  n_25926;
assign n_25928 = ~n_14884 &  n_25927;
assign n_25929 = ~n_14877 &  n_25928;
assign n_25930 = ~n_14871 &  n_25929;
assign n_25931 = ~n_14865 &  n_25930;
assign n_25932 = ~n_14859 &  n_25931;
assign n_25933 = ~n_14853 &  n_25932;
assign n_25934 = ~n_14847 &  n_25933;
assign n_25935 = ~n_14841 &  n_25934;
assign n_25936 = ~n_14835 &  n_25935;
assign n_25937 = ~n_14828 &  n_25936;
assign n_25938 = ~n_14822 &  n_25937;
assign n_25939 = ~n_14816 &  n_25938;
assign n_25940 = ~n_14810 &  n_25939;
assign n_25941 = ~n_14804 &  n_25940;
assign n_25942 = ~n_14798 &  n_25941;
assign n_25943 = ~n_14792 &  n_25942;
assign n_25944 = ~n_14786 &  n_25943;
assign n_25945 = ~n_14779 &  n_25944;
assign n_25946 = ~n_14773 &  n_25945;
assign n_25947 = ~n_14767 &  n_25946;
assign n_25948 = ~n_14761 &  n_25947;
assign n_25949 = ~n_14755 &  n_25948;
assign n_25950 = ~n_14749 &  n_25949;
assign n_25951 = ~n_14743 &  n_25950;
assign n_25952 = ~n_14737 &  n_25951;
assign n_25953 = ~n_14730 &  n_25952;
assign n_25954 = ~n_14724 &  n_25953;
assign n_25955 = ~n_14718 &  n_25954;
assign n_25956 = ~n_14712 &  n_25955;
assign n_25957 = ~n_14706 &  n_25956;
assign n_25958 = ~n_14700 &  n_25957;
assign n_25959 = ~n_14694 &  n_25958;
assign n_25960 = ~n_14688 &  n_25959;
assign n_25961 = ~n_14681 &  n_25960;
assign n_25962 = ~n_14675 &  n_25961;
assign n_25963 = ~n_14669 &  n_25962;
assign n_25964 = ~n_14663 &  n_25963;
assign n_25965 = ~n_14657 &  n_25964;
assign n_25966 = ~n_14651 &  n_25965;
assign n_25967 = ~n_14645 &  n_25966;
assign n_25968 = ~n_14639 &  n_25967;
assign n_25969 = ~n_14632 &  n_25968;
assign n_25970 = ~n_14626 &  n_25969;
assign n_25971 = ~n_14620 &  n_25970;
assign n_25972 = ~n_14614 &  n_25971;
assign n_25973 = ~n_14608 &  n_25972;
assign n_25974 = ~n_14602 &  n_25973;
assign n_25975 = ~n_14596 &  n_25974;
assign n_25976 = ~n_14590 &  n_25975;
assign n_25977 = ~n_14583 &  n_25976;
assign n_25978 = ~n_14577 &  n_25977;
assign n_25979 = ~n_14571 &  n_25978;
assign n_25980 = ~n_14565 &  n_25979;
assign n_25981 = ~n_14559 &  n_25980;
assign n_25982 = ~n_14553 &  n_25981;
assign n_25983 = ~n_14547 &  n_25982;
assign n_25984 = ~n_14541 &  n_25983;
assign n_25985 = ~n_14534 &  n_25984;
assign n_25986 = ~n_14528 &  n_25985;
assign n_25987 = ~n_14522 &  n_25986;
assign n_25988 = ~n_14516 &  n_25987;
assign n_25989 = ~n_14510 &  n_25988;
assign n_25990 = ~n_14504 &  n_25989;
assign n_25991 = ~n_14498 &  n_25990;
assign n_25992 = ~n_14492 &  n_25991;
assign n_25993 = ~n_14485 &  n_25992;
assign n_25994 = ~n_14479 &  n_25993;
assign n_25995 = ~n_14473 &  n_25994;
assign n_25996 = ~n_14467 &  n_25995;
assign n_25997 = ~n_14461 &  n_25996;
assign n_25998 = ~n_14455 &  n_25997;
assign n_25999 = ~n_14449 &  n_25998;
assign n_26000 = ~n_14443 &  n_25999;
assign n_26001 = ~n_14436 &  n_26000;
assign n_26002 = ~n_14430 &  n_26001;
assign n_26003 = ~n_14424 &  n_26002;
assign n_26004 = ~n_14418 &  n_26003;
assign n_26005 = ~n_14412 &  n_26004;
assign n_26006 = ~n_14406 &  n_26005;
assign n_26007 = ~n_14400 &  n_26006;
assign n_26008 = ~n_14394 &  n_26007;
assign n_26009 = ~n_14387 &  n_26008;
assign n_26010 = ~n_14381 &  n_26009;
assign n_26011 = ~n_14375 &  n_26010;
assign n_26012 = ~n_14369 &  n_26011;
assign n_26013 = ~n_14363 &  n_26012;
assign n_26014 = ~n_14357 &  n_26013;
assign n_26015 = ~n_14351 &  n_26014;
assign n_26016 = ~n_14345 &  n_26015;
assign n_26017 = ~n_14338 &  n_26016;
assign n_26018 = ~n_14332 &  n_26017;
assign n_26019 = ~n_14326 &  n_26018;
assign n_26020 = ~n_14320 &  n_26019;
assign n_26021 = ~n_14314 &  n_26020;
assign n_26022 = ~n_14308 &  n_26021;
assign n_26023 = ~n_14302 &  n_26022;
assign n_26024 = ~n_14296 &  n_26023;
assign n_26025 = ~n_14289 &  n_26024;
assign n_26026 = ~n_14283 &  n_26025;
assign n_26027 = ~n_14277 &  n_26026;
assign n_26028 = ~n_14271 &  n_26027;
assign n_26029 = ~n_14265 &  n_26028;
assign n_26030 = ~n_14259 &  n_26029;
assign n_26031 = ~n_14253 &  n_26030;
assign n_26032 = ~n_14247 &  n_26031;
assign n_26033 = ~n_14240 &  n_26032;
assign n_26034 = ~n_14234 &  n_26033;
assign n_26035 = ~n_14228 &  n_26034;
assign n_26036 = ~n_14222 &  n_26035;
assign n_26037 = ~n_14216 &  n_26036;
assign n_26038 = ~n_14210 &  n_26037;
assign n_26039 = ~n_14204 &  n_26038;
assign n_26040 = ~n_14198 &  n_26039;
assign n_26041 = ~n_14191 &  n_26040;
assign n_26042 = ~n_14185 &  n_26041;
assign n_26043 = ~n_14179 &  n_26042;
assign n_26044 = ~n_14173 &  n_26043;
assign n_26045 = ~n_14167 &  n_26044;
assign n_26046 = ~n_14161 &  n_26045;
assign n_26047 = ~n_14155 &  n_26046;
assign n_26048 = ~n_14149 &  n_26047;
assign n_26049 = ~n_14142 &  n_26048;
assign n_26050 = ~n_14136 &  n_26049;
assign n_26051 = ~n_14130 &  n_26050;
assign n_26052 = ~n_14124 &  n_26051;
assign n_26053 = ~n_14118 &  n_26052;
assign n_26054 = ~n_14112 &  n_26053;
assign n_26055 = ~n_14106 &  n_26054;
assign n_26056 = ~n_14100 &  n_26055;
assign n_26057 = ~n_14093 &  n_26056;
assign n_26058 = ~n_14087 &  n_26057;
assign n_26059 = ~n_14081 &  n_26058;
assign n_26060 = ~n_14075 &  n_26059;
assign n_26061 = ~n_14069 &  n_26060;
assign n_26062 = ~n_14063 &  n_26061;
assign n_26063 = ~n_14057 &  n_26062;
assign n_26064 = ~n_14051 &  n_26063;
assign n_26065 = ~n_14044 &  n_26064;
assign n_26066 = ~n_14038 &  n_26065;
assign n_26067 = ~n_14032 &  n_26066;
assign n_26068 = ~n_14026 &  n_26067;
assign n_26069 = ~n_14020 &  n_26068;
assign n_26070 = ~n_14014 &  n_26069;
assign n_26071 = ~n_14008 &  n_26070;
assign n_26072 = ~n_14002 &  n_26071;
assign n_26073 = ~n_13995 &  n_26072;
assign n_26074 = ~n_13989 &  n_26073;
assign n_26075 = ~n_13983 &  n_26074;
assign n_26076 = ~n_13977 &  n_26075;
assign n_26077 = ~n_13971 &  n_26076;
assign n_26078 = ~n_13965 &  n_26077;
assign n_26079 = ~n_13959 &  n_26078;
assign n_26080 = ~n_13953 &  n_26079;
assign n_26081 = ~n_13946 &  n_26080;
assign n_26082 = ~n_13940 &  n_26081;
assign n_26083 = ~n_13934 &  n_26082;
assign n_26084 = ~n_13928 &  n_26083;
assign n_26085 = ~n_13922 &  n_26084;
assign n_26086 = ~n_13916 &  n_26085;
assign n_26087 = ~n_13910 &  n_26086;
assign n_26088 = ~n_13904 &  n_26087;
assign n_26089 = ~n_13898 &  n_26088;
assign n_26090 = ~n_13892 &  n_26089;
assign n_26091 = ~n_13886 &  n_26090;
assign n_26092 = ~n_13880 &  n_26091;
assign n_26093 = ~n_13874 &  n_26092;
assign n_26094 = ~n_13868 &  n_26093;
assign n_26095 = ~n_13862 &  n_26094;
assign n_26096 = ~n_13856 &  n_26095;
assign n_26097 = ~n_13850 &  n_26096;
assign n_26098 = ~n_13844 &  n_26097;
assign n_26099 = ~n_13838 &  n_26098;
assign n_26100 = ~n_13832 &  n_26099;
assign n_26101 = ~n_13826 &  n_26100;
assign n_26102 = ~n_13820 &  n_26101;
assign n_26103 = ~n_13814 &  n_26102;
assign n_26104 = ~n_13808 &  n_26103;
assign n_26105 = ~n_13802 &  n_26104;
assign n_26106 = ~n_13796 &  n_26105;
assign n_26107 = ~n_13790 &  n_26106;
assign n_26108 = ~n_13784 &  n_26107;
assign n_26109 = ~n_13778 &  n_26108;
assign n_26110 = ~n_13772 &  n_26109;
assign n_26111 = ~n_13766 &  n_26110;
assign n_26112 = ~n_13760 &  n_26111;
assign n_26113 = ~n_13754 &  n_26112;
assign n_26114 = ~n_13748 &  n_26113;
assign n_26115 = ~n_13740 &  n_26114;
assign n_26116 = ~n_13708 &  n_26115;
assign n_26117 = ~n_13676 &  n_26116;
assign n_26118 = ~n_13644 &  n_26117;
assign n_26119 = ~n_13612 &  n_26118;
assign n_26120 = ~n_13580 &  n_26119;
assign n_26121 = ~n_13548 &  n_26120;
assign n_26122 = ~n_13516 &  n_26121;
assign n_26123 = ~n_13484 &  n_26122;
assign n_26124 = ~n_13452 &  n_26123;
assign n_26125 = ~n_13420 &  n_26124;
assign n_26126 = ~n_13388 &  n_26125;
assign n_26127 = ~n_13356 &  n_26126;
assign n_26128 = ~n_13324 &  n_26127;
assign n_26129 = ~n_13292 &  n_26128;
assign n_26130 = ~n_13260 &  n_26129;
assign n_26131 = ~n_13228 &  n_26130;
assign n_26132 = ~n_13196 &  n_26131;
assign n_26133 = ~n_13164 &  n_26132;
assign n_26134 = ~n_13132 &  n_26133;
assign n_26135 = ~n_13100 &  n_26134;
assign n_26136 = ~n_13068 &  n_26135;
assign n_26137 = ~n_13036 &  n_26136;
assign n_26138 = ~n_13004 &  n_26137;
assign n_26139 = ~n_12972 &  n_26138;
assign n_26140 = ~n_12940 &  n_26139;
assign n_26141 = ~n_12908 &  n_26140;
assign n_26142 = ~n_12876 &  n_26141;
assign n_26143 = ~n_12844 &  n_26142;
assign n_26144 = ~n_12812 &  n_26143;
assign n_26145 = ~n_12780 &  n_26144;
assign n_26146 = ~n_12748 &  n_26145;
assign n_26147 = ~n_12716 &  n_26146;
assign n_26148 = ~n_12626 &  n_26147;
assign n_26149 = ~n_12623 &  n_26148;
assign n_26150 = ~n_12621 &  n_26149;
assign n_26151 = ~n_12618 &  n_26150;
assign n_26152 = ~n_12615 &  n_26151;
assign n_26153 = ~n_12612 &  n_26152;
assign n_26154 = ~n_12609 &  n_26153;
assign n_26155 = ~n_12606 &  n_26154;
assign n_26156 = ~n_12509 &  n_26155;
assign n_26157 = ~n_12506 &  n_26156;
assign n_26158 = ~n_12503 &  n_26157;
assign n_26159 = ~n_12500 &  n_26158;
assign n_26160 = ~n_12497 &  n_26159;
assign n_26161 = ~n_12494 &  n_26160;
assign n_26162 = ~n_12491 &  n_26161;
assign n_26163 = ~n_12486 &  n_26162;
assign n_26164 = ~n_12482 &  n_26163;
assign n_26165 = ~n_12479 &  n_26164;
assign n_26166 = ~n_12473 &  n_26165;
assign n_26167 = ~n_12464 &  n_26166;
assign n_26168 = ~n_12457 &  n_26167;
assign n_26169 = ~n_12451 &  n_26168;
assign n_26170 = ~n_12444 &  n_26169;
assign n_26171 = ~n_12438 &  n_26170;
assign n_26172 = ~n_12423 &  n_26171;
assign n_26173 = ~n_12420 &  n_26172;
assign n_26174 = ~n_12417 &  n_26173;
assign n_26175 = ~n_12411 &  n_26174;
assign n_26176 = ~n_12405 &  n_26175;
assign n_26177 = ~n_12399 &  n_26176;
assign n_26178 = ~n_12393 &  n_26177;
assign n_26179 = ~n_12386 &  n_26178;
assign n_26180 = ~n_12380 &  n_26179;
assign n_26181 = ~n_12374 &  n_26180;
assign n_26182 = ~n_12368 &  n_26181;
assign n_26183 = ~n_12362 &  n_26182;
assign n_26184 = ~n_12355 &  n_26183;
assign n_26185 = ~n_12349 &  n_26184;
assign n_26186 = ~n_12343 &  n_26185;
assign n_26187 = ~n_12337 &  n_26186;
assign n_26188 = ~n_12330 &  n_26187;
assign n_26189 = ~n_12324 &  n_26188;
assign n_26190 = ~n_12318 &  n_26189;
assign n_26191 = ~n_12312 &  n_26190;
assign n_26192 = ~n_12306 &  n_26191;
assign n_26193 = ~n_12300 &  n_26192;
assign n_26194 = ~n_12293 &  n_26193;
assign n_26195 = ~n_12287 &  n_26194;
assign n_26196 = ~n_12281 &  n_26195;
assign n_26197 = ~n_12275 &  n_26196;
assign n_26198 = ~n_12269 &  n_26197;
assign n_26199 = ~n_12261 &  n_26198;
assign n_26200 = ~n_12257 &  n_26199;
assign n_26201 = ~n_12253 &  n_26200;
assign n_26202 = ~n_12243 &  n_26201;
assign n_26203 = ~n_12237 &  n_26202;
assign n_26204 = ~n_12226 &  n_26203;
assign n_26205 = ~n_12212 &  n_26204;
assign n_26206 = ~n_12199 &  n_26205;
assign n_26207 = ~n_12168 &  n_26206;
assign n_26208 = ~n_12164 &  n_26207;
assign n_26209 = ~n_12159 &  n_26208;
assign n_26210 = ~n_12154 &  n_26209;
assign n_26211 = ~n_12149 &  n_26210;
assign n_26212 = ~n_12144 &  n_26211;
assign n_26213 = ~n_12139 &  n_26212;
assign n_26214 = ~n_12134 &  n_26213;
assign n_26215 = ~n_12129 &  n_26214;
assign n_26216 = ~n_12124 &  n_26215;
assign n_26217 = ~n_12119 &  n_26216;
assign n_26218 = ~n_12114 &  n_26217;
assign n_26219 = ~n_12109 &  n_26218;
assign n_26220 = ~n_12104 &  n_26219;
assign n_26221 = ~n_12099 &  n_26220;
assign n_26222 = ~n_12094 &  n_26221;
assign n_26223 = ~n_12089 &  n_26222;
assign n_26224 = ~n_12084 &  n_26223;
assign n_26225 = ~n_12079 &  n_26224;
assign n_26226 = ~n_12074 &  n_26225;
assign n_26227 = ~n_12069 &  n_26226;
assign n_26228 = ~n_12064 &  n_26227;
assign n_26229 = ~n_12059 &  n_26228;
assign n_26230 = ~n_12054 &  n_26229;
assign n_26231 = ~n_12049 &  n_26230;
assign n_26232 = ~n_12044 &  n_26231;
assign n_26233 = ~n_12039 &  n_26232;
assign n_26234 = ~n_12034 &  n_26233;
assign n_26235 = ~n_12029 &  n_26234;
assign n_26236 = ~n_12024 &  n_26235;
assign n_26237 = ~n_12019 &  n_26236;
assign n_26238 = ~n_12016 &  n_26237;
assign n_26239 = ~n_11980 &  n_26238;
assign n_26240 = ~n_11975 &  n_26239;
assign n_26241 = ~n_11970 &  n_26240;
assign n_26242 = ~n_11964 &  n_26241;
assign n_26243 = ~n_11958 &  n_26242;
assign n_26244 = ~n_11953 &  n_26243;
assign n_26245 = ~n_11943 &  n_26244;
assign n_26246 = ~n_11933 &  n_26245;
assign n_26247 = ~n_11923 &  n_26246;
assign n_26248 = ~n_11917 &  n_26247;
assign n_26249 = ~n_11899 &  n_26248;
assign n_26250 = ~n_11894 &  n_26249;
assign n_26251 = ~n_11884 &  n_26250;
assign n_26252 = ~n_11874 &  n_26251;
assign n_26253 = ~n_11864 &  n_26252;
assign n_26254 = ~n_11858 &  n_26253;
assign n_26255 = ~n_11840 &  n_26254;
assign n_26256 = ~n_11834 &  n_26255;
assign n_26257 = ~n_11829 &  n_26256;
assign n_26258 = ~n_11824 &  n_26257;
assign n_26259 = ~n_11819 &  n_26258;
assign n_26260 = ~n_11809 &  n_26259;
assign n_26261 = ~n_11800 &  n_26260;
assign n_26262 = ~n_11790 &  n_26261;
assign n_26263 = ~n_11784 &  n_26262;
assign n_26264 = ~n_11770 &  n_26263;
assign n_26265 = ~n_11765 &  n_26264;
assign n_26266 = ~n_11760 &  n_26265;
assign n_26267 = ~n_11755 &  n_26266;
assign n_26268 = ~n_11746 &  n_26267;
assign n_26269 = ~n_11741 &  n_26268;
assign n_26270 = ~n_11736 &  n_26269;
assign n_26271 = ~n_11731 &  n_26270;
assign n_26272 = ~n_11726 &  n_26271;
assign n_26273 = ~n_11720 &  n_26272;
assign n_26274 = ~n_11714 &  n_26273;
assign n_26275 = ~n_11708 &  n_26274;
assign n_26276 = ~n_11702 &  n_26275;
assign n_26277 = ~n_11696 &  n_26276;
assign n_26278 = ~n_11690 &  n_26277;
assign n_26279 = ~n_11684 &  n_26278;
assign n_26280 = ~n_11678 &  n_26279;
assign n_26281 = ~n_11672 &  n_26280;
assign n_26282 = ~n_11666 &  n_26281;
assign n_26283 = ~n_11660 &  n_26282;
assign n_26284 = ~n_11654 &  n_26283;
assign n_26285 = ~n_11648 &  n_26284;
assign n_26286 = ~n_11642 &  n_26285;
assign n_26287 = ~n_11636 &  n_26286;
assign n_26288 = ~n_11630 &  n_26287;
assign n_26289 = ~n_11624 &  n_26288;
assign n_26290 = ~n_11618 &  n_26289;
assign n_26291 = ~n_11612 &  n_26290;
assign n_26292 = ~n_11606 &  n_26291;
assign n_26293 = ~n_11600 &  n_26292;
assign n_26294 = ~n_11594 &  n_26293;
assign n_26295 = ~n_11588 &  n_26294;
assign n_26296 = ~n_11582 &  n_26295;
assign n_26297 = ~n_11576 &  n_26296;
assign n_26298 = ~n_11570 &  n_26297;
assign n_26299 = ~n_11564 &  n_26298;
assign n_26300 = ~n_11558 &  n_26299;
assign n_26301 = ~n_11552 &  n_26300;
assign n_26302 = ~n_11546 &  n_26301;
assign n_26303 = ~n_11540 &  n_26302;
assign n_26304 = ~n_11534 &  n_26303;
assign n_26305 = ~n_11528 &  n_26304;
assign n_26306 = ~n_11522 &  n_26305;
assign n_26307 = ~n_11516 &  n_26306;
assign n_26308 = ~n_11510 &  n_26307;
assign n_26309 = ~n_11504 &  n_26308;
assign n_26310 = ~n_11498 &  n_26309;
assign n_26311 = ~n_11492 &  n_26310;
assign n_26312 = ~n_11486 &  n_26311;
assign n_26313 = ~n_11480 &  n_26312;
assign n_26314 = ~n_11474 &  n_26313;
assign n_26315 = ~n_11468 &  n_26314;
assign n_26316 = ~n_11462 &  n_26315;
assign n_26317 = ~n_11456 &  n_26316;
assign n_26318 = ~n_11450 &  n_26317;
assign n_26319 = ~n_11444 &  n_26318;
assign n_26320 = ~n_11438 &  n_26319;
assign n_26321 = ~n_11432 &  n_26320;
assign n_26322 = ~n_11426 &  n_26321;
assign n_26323 = ~n_11420 &  n_26322;
assign n_26324 = ~n_11414 &  n_26323;
assign n_26325 = ~n_11408 &  n_26324;
assign n_26326 = ~n_11402 &  n_26325;
assign n_26327 = ~n_11396 &  n_26326;
assign n_26328 = ~n_11390 &  n_26327;
assign n_26329 = ~n_11384 &  n_26328;
assign n_26330 = ~n_11378 &  n_26329;
assign n_26331 = ~n_11372 &  n_26330;
assign n_26332 = ~n_11366 &  n_26331;
assign n_26333 = ~n_11360 &  n_26332;
assign n_26334 = ~n_11354 &  n_26333;
assign n_26335 = ~n_11348 &  n_26334;
assign n_26336 = ~n_11342 &  n_26335;
assign n_26337 = ~n_11336 &  n_26336;
assign n_26338 = ~n_11330 &  n_26337;
assign n_26339 = ~n_11324 &  n_26338;
assign n_26340 = ~n_11318 &  n_26339;
assign n_26341 = ~n_11312 &  n_26340;
assign n_26342 = ~n_11306 &  n_26341;
assign n_26343 = ~n_11300 &  n_26342;
assign n_26344 = ~n_11294 &  n_26343;
assign n_26345 = ~n_11288 &  n_26344;
assign n_26346 = ~n_11282 &  n_26345;
assign n_26347 = ~n_11276 &  n_26346;
assign n_26348 = ~n_11270 &  n_26347;
assign n_26349 = ~n_11264 &  n_26348;
assign n_26350 = ~n_11258 &  n_26349;
assign n_26351 = ~n_11252 &  n_26350;
assign n_26352 = ~n_11246 &  n_26351;
assign n_26353 = ~n_11240 &  n_26352;
assign n_26354 = ~n_11234 &  n_26353;
assign n_26355 = ~n_11228 &  n_26354;
assign n_26356 = ~n_11222 &  n_26355;
assign n_26357 = ~n_11216 &  n_26356;
assign n_26358 = ~n_11210 &  n_26357;
assign n_26359 = ~n_11204 &  n_26358;
assign n_26360 = ~n_11198 &  n_26359;
assign n_26361 = ~n_11192 &  n_26360;
assign n_26362 = ~n_11186 &  n_26361;
assign n_26363 = ~n_11180 &  n_26362;
assign n_26364 = ~n_11174 &  n_26363;
assign n_26365 = ~n_11168 &  n_26364;
assign n_26366 = ~n_11162 &  n_26365;
assign n_26367 = ~n_11156 &  n_26366;
assign n_26368 = ~n_11150 &  n_26367;
assign n_26369 = ~n_11144 &  n_26368;
assign n_26370 = ~n_11138 &  n_26369;
assign n_26371 = ~n_11132 &  n_26370;
assign n_26372 = ~n_11126 &  n_26371;
assign n_26373 = ~n_11120 &  n_26372;
assign n_26374 = ~n_11114 &  n_26373;
assign n_26375 = ~n_11108 &  n_26374;
assign n_26376 = ~n_11102 &  n_26375;
assign n_26377 = ~n_11096 &  n_26376;
assign n_26378 = ~n_11090 &  n_26377;
assign n_26379 = ~n_11084 &  n_26378;
assign n_26380 = ~n_11078 &  n_26379;
assign n_26381 = ~n_11072 &  n_26380;
assign n_26382 = ~n_11066 &  n_26381;
assign n_26383 = ~n_11060 &  n_26382;
assign n_26384 = ~n_11054 &  n_26383;
assign n_26385 = ~n_11048 &  n_26384;
assign n_26386 = ~n_11042 &  n_26385;
assign n_26387 = ~n_11036 &  n_26386;
assign n_26388 = ~n_11030 &  n_26387;
assign n_26389 = ~n_11024 &  n_26388;
assign n_26390 = ~n_11018 &  n_26389;
assign n_26391 = ~n_11012 &  n_26390;
assign n_26392 = ~n_11006 &  n_26391;
assign n_26393 = ~n_11000 &  n_26392;
assign n_26394 = ~n_10994 &  n_26393;
assign n_26395 = ~n_10988 &  n_26394;
assign n_26396 = ~n_10982 &  n_26395;
assign n_26397 = ~n_10976 &  n_26396;
assign n_26398 = ~n_10970 &  n_26397;
assign n_26399 = ~n_10964 &  n_26398;
assign n_26400 = ~n_10958 &  n_26399;
assign n_26401 = ~n_10952 &  n_26400;
assign n_26402 = ~n_10946 &  n_26401;
assign n_26403 = ~n_10940 &  n_26402;
assign n_26404 = ~n_10934 &  n_26403;
assign n_26405 = ~n_10928 &  n_26404;
assign n_26406 = ~n_10922 &  n_26405;
assign n_26407 = ~n_10916 &  n_26406;
assign n_26408 = ~n_10910 &  n_26407;
assign n_26409 = ~n_10904 &  n_26408;
assign n_26410 = ~n_10898 &  n_26409;
assign n_26411 = ~n_10892 &  n_26410;
assign n_26412 = ~n_10886 &  n_26411;
assign n_26413 = ~n_10880 &  n_26412;
assign n_26414 = ~n_10874 &  n_26413;
assign n_26415 = ~n_10868 &  n_26414;
assign n_26416 = ~n_10862 &  n_26415;
assign n_26417 = ~n_10856 &  n_26416;
assign n_26418 = ~n_10850 &  n_26417;
assign n_26419 = ~n_10844 &  n_26418;
assign n_26420 = ~n_10838 &  n_26419;
assign n_26421 = ~n_10832 &  n_26420;
assign n_26422 = ~n_10826 &  n_26421;
assign n_26423 = ~n_10820 &  n_26422;
assign n_26424 = ~n_10814 &  n_26423;
assign n_26425 = ~n_10808 &  n_26424;
assign n_26426 = ~n_10802 &  n_26425;
assign n_26427 = ~n_10796 &  n_26426;
assign n_26428 = ~n_10790 &  n_26427;
assign n_26429 = ~n_10784 &  n_26428;
assign n_26430 = ~n_10778 &  n_26429;
assign n_26431 = ~n_10772 &  n_26430;
assign n_26432 = ~n_10766 &  n_26431;
assign n_26433 = ~n_10760 &  n_26432;
assign n_26434 = ~n_10754 &  n_26433;
assign n_26435 = ~n_10748 &  n_26434;
assign n_26436 = ~n_10742 &  n_26435;
assign n_26437 = ~n_10736 &  n_26436;
assign n_26438 = ~n_10730 &  n_26437;
assign n_26439 = ~n_10724 &  n_26438;
assign n_26440 = ~n_10718 &  n_26439;
assign n_26441 = ~n_10712 &  n_26440;
assign n_26442 = ~n_10706 &  n_26441;
assign n_26443 = ~n_10700 &  n_26442;
assign n_26444 = ~n_10694 &  n_26443;
assign n_26445 = ~n_10688 &  n_26444;
assign n_26446 = ~n_10682 &  n_26445;
assign n_26447 = ~n_10676 &  n_26446;
assign n_26448 = ~n_10670 &  n_26447;
assign n_26449 = ~n_10664 &  n_26448;
assign n_26450 = ~n_10658 &  n_26449;
assign n_26451 = ~n_10652 &  n_26450;
assign n_26452 = ~n_10646 &  n_26451;
assign n_26453 = ~n_10640 &  n_26452;
assign n_26454 = ~n_10634 &  n_26453;
assign n_26455 = ~n_10628 &  n_26454;
assign n_26456 = ~n_10622 &  n_26455;
assign n_26457 = ~n_10616 &  n_26456;
assign n_26458 = ~n_10610 &  n_26457;
assign n_26459 = ~n_10604 &  n_26458;
assign n_26460 = ~n_10598 &  n_26459;
assign n_26461 = ~n_10592 &  n_26460;
assign n_26462 = ~n_10586 &  n_26461;
assign n_26463 = ~n_10580 &  n_26462;
assign n_26464 = ~n_10574 &  n_26463;
assign n_26465 = ~n_10568 &  n_26464;
assign n_26466 = ~n_10562 &  n_26465;
assign n_26467 = ~n_10556 &  n_26466;
assign n_26468 = ~n_10550 &  n_26467;
assign n_26469 = ~n_10544 &  n_26468;
assign n_26470 = ~n_10538 &  n_26469;
assign n_26471 = ~n_10532 &  n_26470;
assign n_26472 = ~n_10526 &  n_26471;
assign n_26473 = ~n_10520 &  n_26472;
assign n_26474 = ~n_10514 &  n_26473;
assign n_26475 = ~n_10508 &  n_26474;
assign n_26476 = ~n_10502 &  n_26475;
assign n_26477 = ~n_10496 &  n_26476;
assign n_26478 = ~n_10490 &  n_26477;
assign n_26479 = ~n_10484 &  n_26478;
assign n_26480 = ~n_10478 &  n_26479;
assign n_26481 = ~n_10472 &  n_26480;
assign n_26482 = ~n_10466 &  n_26481;
assign n_26483 = ~n_10460 &  n_26482;
assign n_26484 = ~n_10454 &  n_26483;
assign n_26485 = ~n_10448 &  n_26484;
assign n_26486 = ~n_10442 &  n_26485;
assign n_26487 = ~n_10436 &  n_26486;
assign n_26488 = ~n_10430 &  n_26487;
assign n_26489 = ~n_10424 &  n_26488;
assign n_26490 = ~n_10418 &  n_26489;
assign n_26491 = ~n_10412 &  n_26490;
assign n_26492 = ~n_10406 &  n_26491;
assign n_26493 = ~n_10400 &  n_26492;
assign n_26494 = ~n_10394 &  n_26493;
assign n_26495 = ~n_10388 &  n_26494;
assign n_26496 = ~n_10382 &  n_26495;
assign n_26497 = ~n_10376 &  n_26496;
assign n_26498 = ~n_10370 &  n_26497;
assign n_26499 = ~n_10364 &  n_26498;
assign n_26500 = ~n_10358 &  n_26499;
assign n_26501 = ~n_10352 &  n_26500;
assign n_26502 = ~n_10346 &  n_26501;
assign n_26503 = ~n_10340 &  n_26502;
assign n_26504 = ~n_10334 &  n_26503;
assign n_26505 = ~n_10328 &  n_26504;
assign n_26506 = ~n_10322 &  n_26505;
assign n_26507 = ~n_10316 &  n_26506;
assign n_26508 = ~n_10310 &  n_26507;
assign n_26509 = ~n_10304 &  n_26508;
assign n_26510 = ~n_10298 &  n_26509;
assign n_26511 = ~n_10292 &  n_26510;
assign n_26512 = ~n_10286 &  n_26511;
assign n_26513 = ~n_10280 &  n_26512;
assign n_26514 = ~n_10274 &  n_26513;
assign n_26515 = ~n_10268 &  n_26514;
assign n_26516 = ~n_10262 &  n_26515;
assign n_26517 = ~n_10256 &  n_26516;
assign n_26518 = ~n_10250 &  n_26517;
assign n_26519 = ~n_10244 &  n_26518;
assign n_26520 = ~n_10238 &  n_26519;
assign n_26521 = ~n_10232 &  n_26520;
assign n_26522 = ~n_10226 &  n_26521;
assign n_26523 = ~n_10220 &  n_26522;
assign n_26524 = ~n_10214 &  n_26523;
assign n_26525 = ~n_10208 &  n_26524;
assign n_26526 = ~n_10202 &  n_26525;
assign n_26527 = ~n_10196 &  n_26526;
assign n_26528 = ~n_10190 &  n_26527;
assign n_26529 = ~n_10184 &  n_26528;
assign n_26530 = ~n_10178 &  n_26529;
assign n_26531 = ~n_10172 &  n_26530;
assign n_26532 = ~n_10166 &  n_26531;
assign n_26533 = ~n_10160 &  n_26532;
assign n_26534 = ~n_10154 &  n_26533;
assign n_26535 = ~n_10148 &  n_26534;
assign n_26536 = ~n_10142 &  n_26535;
assign n_26537 = ~n_10136 &  n_26536;
assign n_26538 = ~n_10130 &  n_26537;
assign n_26539 = ~n_10124 &  n_26538;
assign n_26540 = ~n_10118 &  n_26539;
assign n_26541 = ~n_10112 &  n_26540;
assign n_26542 = ~n_10106 &  n_26541;
assign n_26543 = ~n_10100 &  n_26542;
assign n_26544 = ~n_10094 &  n_26543;
assign n_26545 = ~n_10088 &  n_26544;
assign n_26546 = ~n_10082 &  n_26545;
assign n_26547 = ~n_10076 &  n_26546;
assign n_26548 = ~n_10070 &  n_26547;
assign n_26549 = ~n_10064 &  n_26548;
assign n_26550 = ~n_10058 &  n_26549;
assign n_26551 = ~n_10052 &  n_26550;
assign n_26552 = ~n_10046 &  n_26551;
assign n_26553 = ~n_10040 &  n_26552;
assign n_26554 = ~n_10034 &  n_26553;
assign n_26555 = ~n_10028 &  n_26554;
assign n_26556 = ~n_10022 &  n_26555;
assign n_26557 = ~n_10016 &  n_26556;
assign n_26558 = ~n_10010 &  n_26557;
assign n_26559 = ~n_10004 &  n_26558;
assign n_26560 = ~n_9998 &  n_26559;
assign n_26561 = ~n_9992 &  n_26560;
assign n_26562 = ~n_9986 &  n_26561;
assign n_26563 = ~n_9980 &  n_26562;
assign n_26564 = ~n_9974 &  n_26563;
assign n_26565 = ~n_9968 &  n_26564;
assign n_26566 = ~n_9962 &  n_26565;
assign n_26567 = ~n_9956 &  n_26566;
assign n_26568 = ~n_9950 &  n_26567;
assign n_26569 = ~n_9944 &  n_26568;
assign n_26570 = ~n_9938 &  n_26569;
assign n_26571 = ~n_9932 &  n_26570;
assign n_26572 = ~n_9926 &  n_26571;
assign n_26573 = ~n_9920 &  n_26572;
assign n_26574 = ~n_9914 &  n_26573;
assign n_26575 = ~n_9908 &  n_26574;
assign n_26576 = ~n_9902 &  n_26575;
assign n_26577 = ~n_9896 &  n_26576;
assign n_26578 = ~n_9890 &  n_26577;
assign n_26579 = ~n_9884 &  n_26578;
assign n_26580 = ~n_9878 &  n_26579;
assign n_26581 = ~n_9872 &  n_26580;
assign n_26582 = ~n_9866 &  n_26581;
assign n_26583 = ~n_9860 &  n_26582;
assign n_26584 = ~n_9854 &  n_26583;
assign n_26585 = ~n_9848 &  n_26584;
assign n_26586 = ~n_9842 &  n_26585;
assign n_26587 = ~n_9836 &  n_26586;
assign n_26588 = ~n_9830 &  n_26587;
assign n_26589 = ~n_9824 &  n_26588;
assign n_26590 = ~n_9818 &  n_26589;
assign n_26591 = ~n_9812 &  n_26590;
assign n_26592 = ~n_9806 &  n_26591;
assign n_26593 = ~n_9800 &  n_26592;
assign n_26594 = ~n_9794 &  n_26593;
assign n_26595 = ~n_9788 &  n_26594;
assign n_26596 = ~n_9782 &  n_26595;
assign n_26597 = ~n_9776 &  n_26596;
assign n_26598 = ~n_9770 &  n_26597;
assign n_26599 = ~n_9764 &  n_26598;
assign n_26600 = ~n_9758 &  n_26599;
assign n_26601 = ~n_9752 &  n_26600;
assign n_26602 = ~n_9746 &  n_26601;
assign n_26603 = ~n_9740 &  n_26602;
assign n_26604 = ~n_9734 &  n_26603;
assign n_26605 = ~n_9728 &  n_26604;
assign n_26606 = ~n_9722 &  n_26605;
assign n_26607 = ~n_9716 &  n_26606;
assign n_26608 = ~n_9710 &  n_26607;
assign n_26609 = ~n_9704 &  n_26608;
assign n_26610 = ~n_9698 &  n_26609;
assign n_26611 = ~n_9692 &  n_26610;
assign n_26612 = ~n_9686 &  n_26611;
assign n_26613 = ~n_9680 &  n_26612;
assign n_26614 = ~n_9674 &  n_26613;
assign n_26615 = ~n_9668 &  n_26614;
assign n_26616 = ~n_9662 &  n_26615;
assign n_26617 = ~n_9656 &  n_26616;
assign n_26618 = ~n_9650 &  n_26617;
assign n_26619 = ~n_9644 &  n_26618;
assign n_26620 = ~n_9638 &  n_26619;
assign n_26621 = ~n_9632 &  n_26620;
assign n_26622 = ~n_9626 &  n_26621;
assign n_26623 = ~n_9620 &  n_26622;
assign n_26624 = ~n_9614 &  n_26623;
assign n_26625 = ~n_9608 &  n_26624;
assign n_26626 = ~n_9602 &  n_26625;
assign n_26627 = ~n_9596 &  n_26626;
assign n_26628 = ~n_9590 &  n_26627;
assign n_26629 = ~n_9584 &  n_26628;
assign n_26630 = ~n_9578 &  n_26629;
assign n_26631 = ~n_9572 &  n_26630;
assign n_26632 = ~n_9566 &  n_26631;
assign n_26633 = ~n_9560 &  n_26632;
assign n_26634 = ~n_9554 &  n_26633;
assign n_26635 = ~n_9548 &  n_26634;
assign n_26636 = ~n_9542 &  n_26635;
assign n_26637 = ~n_9536 &  n_26636;
assign n_26638 = ~n_9530 &  n_26637;
assign n_26639 = ~n_9524 &  n_26638;
assign n_26640 = ~n_9518 &  n_26639;
assign n_26641 = ~n_9512 &  n_26640;
assign n_26642 = ~n_9506 &  n_26641;
assign n_26643 = ~n_9500 &  n_26642;
assign n_26644 = ~n_9494 &  n_26643;
assign n_26645 = ~n_9488 &  n_26644;
assign n_26646 = ~n_9482 &  n_26645;
assign n_26647 = ~n_9476 &  n_26646;
assign n_26648 = ~n_9470 &  n_26647;
assign n_26649 = ~n_9464 &  n_26648;
assign n_26650 = ~n_9458 &  n_26649;
assign n_26651 = ~n_9452 &  n_26650;
assign n_26652 = ~n_9446 &  n_26651;
assign n_26653 = ~n_9440 &  n_26652;
assign n_26654 = ~n_9434 &  n_26653;
assign n_26655 = ~n_9428 &  n_26654;
assign n_26656 = ~n_9422 &  n_26655;
assign n_26657 = ~n_9416 &  n_26656;
assign n_26658 = ~n_9410 &  n_26657;
assign n_26659 = ~n_9404 &  n_26658;
assign n_26660 = ~n_9398 &  n_26659;
assign n_26661 = ~n_9392 &  n_26660;
assign n_26662 = ~n_9386 &  n_26661;
assign n_26663 = ~n_9380 &  n_26662;
assign n_26664 = ~n_9374 &  n_26663;
assign n_26665 = ~n_9368 &  n_26664;
assign n_26666 = ~n_9362 &  n_26665;
assign n_26667 = ~n_9356 &  n_26666;
assign n_26668 = ~n_9350 &  n_26667;
assign n_26669 = ~n_9344 &  n_26668;
assign n_26670 = ~n_9338 &  n_26669;
assign n_26671 = ~n_9332 &  n_26670;
assign n_26672 = ~n_9326 &  n_26671;
assign n_26673 = ~n_9320 &  n_26672;
assign n_26674 = ~n_9314 &  n_26673;
assign n_26675 = ~n_9308 &  n_26674;
assign n_26676 = ~n_9302 &  n_26675;
assign n_26677 = ~n_9296 &  n_26676;
assign n_26678 = ~n_9290 &  n_26677;
assign n_26679 = ~n_9284 &  n_26678;
assign n_26680 = ~n_9278 &  n_26679;
assign n_26681 = ~n_9272 &  n_26680;
assign n_26682 = ~n_9266 &  n_26681;
assign n_26683 = ~n_9260 &  n_26682;
assign n_26684 = ~n_9254 &  n_26683;
assign n_26685 = ~n_9248 &  n_26684;
assign n_26686 = ~n_9242 &  n_26685;
assign n_26687 = ~n_9236 &  n_26686;
assign n_26688 = ~n_9230 &  n_26687;
assign n_26689 = ~n_9224 &  n_26688;
assign n_26690 = ~n_9218 &  n_26689;
assign n_26691 = ~n_9212 &  n_26690;
assign n_26692 = ~n_9206 &  n_26691;
assign n_26693 = ~n_9200 &  n_26692;
assign n_26694 = ~n_9194 &  n_26693;
assign n_26695 = ~n_9188 &  n_26694;
assign n_26696 = ~n_9182 &  n_26695;
assign n_26697 = ~n_9176 &  n_26696;
assign n_26698 = ~n_9170 &  n_26697;
assign n_26699 = ~n_9164 &  n_26698;
assign n_26700 = ~n_9158 &  n_26699;
assign n_26701 = ~n_9152 &  n_26700;
assign n_26702 = ~n_9146 &  n_26701;
assign n_26703 = ~n_9140 &  n_26702;
assign n_26704 = ~n_9134 &  n_26703;
assign n_26705 = ~n_9128 &  n_26704;
assign n_26706 = ~n_9122 &  n_26705;
assign n_26707 = ~n_9116 &  n_26706;
assign n_26708 = ~n_9110 &  n_26707;
assign n_26709 = ~n_9104 &  n_26708;
assign n_26710 = ~n_9098 &  n_26709;
assign n_26711 = ~n_9092 &  n_26710;
assign n_26712 = ~n_9086 &  n_26711;
assign n_26713 = ~n_9080 &  n_26712;
assign n_26714 = ~n_9074 &  n_26713;
assign n_26715 = ~n_9068 &  n_26714;
assign n_26716 = ~n_9062 &  n_26715;
assign n_26717 = ~n_9056 &  n_26716;
assign n_26718 = ~n_9050 &  n_26717;
assign n_26719 = ~n_9044 &  n_26718;
assign n_26720 = ~n_9038 &  n_26719;
assign n_26721 = ~n_9032 &  n_26720;
assign n_26722 = ~n_9026 &  n_26721;
assign n_26723 = ~n_9020 &  n_26722;
assign n_26724 = ~n_9014 &  n_26723;
assign n_26725 = ~n_9008 &  n_26724;
assign n_26726 = ~n_9002 &  n_26725;
assign n_26727 = ~n_8996 &  n_26726;
assign n_26728 = ~n_8990 &  n_26727;
assign n_26729 = ~n_8984 &  n_26728;
assign n_26730 = ~n_8978 &  n_26729;
assign n_26731 = ~n_8972 &  n_26730;
assign n_26732 = ~n_8966 &  n_26731;
assign n_26733 = ~n_8960 &  n_26732;
assign n_26734 = ~n_8954 &  n_26733;
assign n_26735 = ~n_8948 &  n_26734;
assign n_26736 = ~n_8942 &  n_26735;
assign n_26737 = ~n_8936 &  n_26736;
assign n_26738 = ~n_8930 &  n_26737;
assign n_26739 = ~n_8924 &  n_26738;
assign n_26740 = ~n_8918 &  n_26739;
assign n_26741 = ~n_8912 &  n_26740;
assign n_26742 = ~n_8906 &  n_26741;
assign n_26743 = ~n_8900 &  n_26742;
assign n_26744 = ~n_8894 &  n_26743;
assign n_26745 = ~n_8888 &  n_26744;
assign n_26746 = ~n_8882 &  n_26745;
assign n_26747 = ~n_8876 &  n_26746;
assign n_26748 = ~n_8870 &  n_26747;
assign n_26749 = ~n_8864 &  n_26748;
assign n_26750 = ~n_8858 &  n_26749;
assign n_26751 = ~n_8852 &  n_26750;
assign n_26752 = ~n_8846 &  n_26751;
assign n_26753 = ~n_8840 &  n_26752;
assign n_26754 = ~n_8834 &  n_26753;
assign n_26755 = ~n_8828 &  n_26754;
assign n_26756 = ~n_8822 &  n_26755;
assign n_26757 = ~n_8816 &  n_26756;
assign n_26758 = ~n_8810 &  n_26757;
assign n_26759 = ~n_8804 &  n_26758;
assign n_26760 = ~n_8798 &  n_26759;
assign n_26761 = ~n_8792 &  n_26760;
assign n_26762 = ~n_8786 &  n_26761;
assign n_26763 = ~n_8780 &  n_26762;
assign n_26764 = ~n_8774 &  n_26763;
assign n_26765 = ~n_8768 &  n_26764;
assign n_26766 = ~n_8762 &  n_26765;
assign n_26767 = ~n_8756 &  n_26766;
assign n_26768 = ~n_8750 &  n_26767;
assign n_26769 = ~n_8742 &  n_26768;
assign n_26770 = ~n_8735 &  n_26769;
assign n_26771 = ~n_8727 &  n_26770;
assign n_26772 = ~n_8720 &  n_26771;
assign n_26773 = ~n_8712 &  n_26772;
assign n_26774 = ~n_8705 &  n_26773;
assign n_26775 = ~n_8697 &  n_26774;
assign n_26776 = ~n_8690 &  n_26775;
assign n_26777 = ~n_8682 &  n_26776;
assign n_26778 = ~n_8675 &  n_26777;
assign n_26779 = ~n_8667 &  n_26778;
assign n_26780 = ~n_8660 &  n_26779;
assign n_26781 = ~n_8651 &  n_26780;
assign n_26782 = ~n_8644 &  n_26781;
assign n_26783 = ~n_8635 &  n_26782;
assign n_26784 = ~n_8621 &  n_26783;
assign n_26785 = ~n_8616 &  n_26784;
assign n_26786 = ~n_8610 &  n_26785;
assign n_26787 = ~n_8604 &  n_26786;
assign n_26788 = ~n_8599 &  n_26787;
assign n_26789 = ~n_8593 &  n_26788;
assign n_26790 = ~n_8588 &  n_26789;
assign n_26791 = ~n_8582 &  n_26790;
assign n_26792 = ~n_8577 &  n_26791;
assign n_26793 = ~n_8572 &  n_26792;
assign n_26794 = ~n_8567 &  n_26793;
assign n_26795 = ~n_8562 &  n_26794;
assign n_26796 = ~n_8557 &  n_26795;
assign n_26797 = ~n_8552 &  n_26796;
assign n_26798 = ~n_8547 &  n_26797;
assign n_26799 = ~n_8542 &  n_26798;
assign n_26800 = ~n_8537 &  n_26799;
assign n_26801 = ~n_8532 &  n_26800;
assign n_26802 = ~n_8527 &  n_26801;
assign n_26803 = ~n_8522 &  n_26802;
assign n_26804 = ~n_8517 &  n_26803;
assign n_26805 = ~n_8512 &  n_26804;
assign n_26806 = ~n_8507 &  n_26805;
assign n_26807 = ~n_8502 &  n_26806;
assign n_26808 = ~n_8497 &  n_26807;
assign n_26809 = ~n_8492 &  n_26808;
assign n_26810 = ~n_8487 &  n_26809;
assign n_26811 = ~n_8482 &  n_26810;
assign n_26812 = ~n_8477 &  n_26811;
assign n_26813 = ~n_8472 &  n_26812;
assign n_26814 = ~n_8467 &  n_26813;
assign n_26815 = ~n_8462 &  n_26814;
assign n_26816 = ~n_8457 &  n_26815;
assign n_26817 = ~n_8452 &  n_26816;
assign n_26818 = ~n_8447 &  n_26817;
assign n_26819 = ~n_8442 &  n_26818;
assign n_26820 = ~n_8437 &  n_26819;
assign n_26821 = ~n_8434 &  n_26820;
assign n_26822 = ~n_8400 &  n_26821;
assign n_26823 = ~n_8396 &  n_26822;
assign n_26824 = ~n_8390 &  n_26823;
assign n_26825 = ~n_8387 &  n_26824;
assign n_26826 = ~n_8384 &  n_26825;
assign n_26827 = ~n_8381 &  n_26826;
assign n_26828 = ~n_8378 &  n_26827;
assign n_26829 = ~n_8375 &  n_26828;
assign n_26830 = ~n_8372 &  n_26829;
assign n_26831 = ~n_8369 &  n_26830;
assign n_26832 = ~n_8366 &  n_26831;
assign n_26833 = ~n_8363 &  n_26832;
assign n_26834 = ~n_8360 &  n_26833;
assign n_26835 = ~n_8357 &  n_26834;
assign n_26836 = ~n_8354 &  n_26835;
assign n_26837 = ~n_8351 &  n_26836;
assign n_26838 = ~n_8348 &  n_26837;
assign n_26839 = ~n_8345 &  n_26838;
assign n_26840 = ~n_8342 &  n_26839;
assign n_26841 = ~n_8339 &  n_26840;
assign n_26842 = ~n_8336 &  n_26841;
assign n_26843 = ~n_8333 &  n_26842;
assign n_26844 = ~n_8330 &  n_26843;
assign n_26845 = ~n_8327 &  n_26844;
assign n_26846 = ~n_8324 &  n_26845;
assign n_26847 = ~n_8321 &  n_26846;
assign n_26848 = ~n_8318 &  n_26847;
assign n_26849 = ~n_8315 &  n_26848;
assign n_26850 = ~n_8312 &  n_26849;
assign n_26851 = ~n_8309 &  n_26850;
assign n_26852 = ~n_8306 &  n_26851;
assign n_26853 = ~n_8303 &  n_26852;
assign n_26854 = ~n_8300 &  n_26853;
assign n_26855 = ~n_8297 &  n_26854;
assign n_26856 = ~n_8294 &  n_26855;
assign n_26857 = ~n_8289 &  n_26856;
assign n_26858 = ~n_8284 &  n_26857;
assign n_26859 = ~n_8278 &  n_26858;
assign n_26860 = ~n_8275 &  n_26859;
assign n_26861 = ~n_8269 &  n_26860;
assign n_26862 = ~n_8263 &  n_26861;
assign n_26863 = ~n_8257 &  n_26862;
assign n_26864 = ~n_8251 &  n_26863;
assign n_26865 = ~n_8245 &  n_26864;
assign n_26866 = ~n_8239 &  n_26865;
assign n_26867 = ~n_8233 &  n_26866;
assign n_26868 = ~n_8227 &  n_26867;
assign n_26869 = ~n_8222 &  n_26868;
assign n_26870 = ~n_8217 &  n_26869;
assign n_26871 = ~n_8213 &  n_26870;
assign n_26872 = ~n_8209 &  n_26871;
assign n_26873 = ~n_8205 &  n_26872;
assign n_26874 = ~n_8202 &  n_26873;
assign n_26875 = ~n_8199 &  n_26874;
assign n_26876 = ~n_8166 &  n_26875;
assign n_26877 = ~n_8133 &  n_26876;
assign n_26878 = ~n_8100 &  n_26877;
assign n_26879 = ~n_8067 &  n_26878;
assign n_26880 = ~n_8034 &  n_26879;
assign n_26881 = ~n_8001 &  n_26880;
assign n_26882 = ~n_7997 &  n_26881;
assign n_26883 = ~n_7967 &  n_26882;
assign n_26884 = ~n_7934 &  n_26883;
assign n_26885 = ~n_7901 &  n_26884;
assign n_26886 = ~n_7868 &  n_26885;
assign n_26887 = ~n_7835 &  n_26886;
assign n_26888 = ~n_7802 &  n_26887;
assign n_26889 = ~n_7769 &  n_26888;
assign n_26890 = ~n_7736 &  n_26889;
assign n_26891 = ~n_7732 &  n_26890;
assign n_26892 = ~n_7702 &  n_26891;
assign n_26893 = ~n_7669 &  n_26892;
assign n_26894 = ~n_7636 &  n_26893;
assign n_26895 = ~n_7603 &  n_26894;
assign n_26896 = ~n_7570 &  n_26895;
assign n_26897 = ~n_7537 &  n_26896;
assign n_26898 = ~n_7504 &  n_26897;
assign n_26899 = ~n_7471 &  n_26898;
assign n_26900 = ~n_7467 &  n_26899;
assign n_26901 = ~n_7437 &  n_26900;
assign n_26902 = ~n_7404 &  n_26901;
assign n_26903 = ~n_7371 &  n_26902;
assign n_26904 = ~n_7338 &  n_26903;
assign n_26905 = ~n_7305 &  n_26904;
assign n_26906 = ~n_7272 &  n_26905;
assign n_26907 = ~n_7239 &  n_26906;
assign n_26908 = ~n_7206 &  n_26907;
assign n_26909 = ~n_7202 &  n_26908;
assign n_26910 = ~n_7172 &  n_26909;
assign n_26911 = ~n_7139 &  n_26910;
assign n_26912 = ~n_7106 &  n_26911;
assign n_26913 = ~n_7073 &  n_26912;
assign n_26914 = ~n_7040 &  n_26913;
assign n_26915 = ~n_7007 &  n_26914;
assign n_26916 = ~n_6974 &  n_26915;
assign n_26917 = ~n_6941 &  n_26916;
assign n_26918 = ~n_6937 &  n_26917;
assign n_26919 = ~n_6907 &  n_26918;
assign n_26920 = ~n_6874 &  n_26919;
assign n_26921 = ~n_6841 &  n_26920;
assign n_26922 = ~n_6808 &  n_26921;
assign n_26923 = ~n_6775 &  n_26922;
assign n_26924 = ~n_6742 &  n_26923;
assign n_26925 = ~n_6709 &  n_26924;
assign n_26926 = ~n_6676 &  n_26925;
assign n_26927 = ~n_6672 &  n_26926;
assign n_26928 = ~n_6642 &  n_26927;
assign n_26929 = ~n_6609 &  n_26928;
assign n_26930 = ~n_6576 &  n_26929;
assign n_26931 = ~n_6543 &  n_26930;
assign n_26932 = ~n_6510 &  n_26931;
assign n_26933 = ~n_6477 &  n_26932;
assign n_26934 = ~n_6444 &  n_26933;
assign n_26935 = ~n_6411 &  n_26934;
assign n_26936 = ~n_6407 &  n_26935;
assign n_26937 = ~n_6377 &  n_26936;
assign n_26938 = ~n_6344 &  n_26937;
assign n_26939 = ~n_6311 &  n_26938;
assign n_26940 = ~n_6278 &  n_26939;
assign n_26941 = ~n_6245 &  n_26940;
assign n_26942 = ~n_6212 &  n_26941;
assign n_26943 = ~n_6179 &  n_26942;
assign n_26944 = ~n_6141 &  n_26943;
assign n_26945 = ~n_6108 &  n_26944;
assign n_26946 = ~n_4367 &  n_26945;
assign n_26947 = ~n_4345 &  n_26946;
assign n_26948 = ~n_4301 &  n_26947;
assign n_26949 = ~n_3987 &  n_26948;
assign n_26950 = ~n_3983 &  n_26949;
assign n_26951 = ~n_3945 &  n_26950;
assign n_26952 = ~n_3725 &  n_26951;
assign n_26953 = ~n_3712 &  n_26952;
assign n_26954 = ~n_3553 &  n_26953;
assign n_26955 =  x_295 &  n_26954;
assign n_26956 = ~n_3516 &  n_26955;
assign n_26957 = ~n_3510 &  n_26956;
assign n_26958 = ~n_3504 &  n_26957;
assign n_26959 = ~n_3498 &  n_26958;
assign n_26960 = ~n_3492 &  n_26959;
assign n_26961 = ~n_3486 &  n_26960;
assign n_26962 = ~n_3479 &  n_26961;
assign n_26963 = ~n_3473 &  n_26962;
assign n_26964 = ~n_3467 &  n_26963;
assign n_26965 = ~n_3461 &  n_26964;
assign n_26966 = ~n_3455 &  n_26965;
assign n_26967 = ~n_3449 &  n_26966;
assign n_26968 = ~n_3443 &  n_26967;
assign n_26969 = ~n_3437 &  n_26968;
assign n_26970 = ~n_3431 &  n_26969;
assign n_26971 = ~n_3424 &  n_26970;
assign n_26972 = ~n_3418 &  n_26971;
assign n_26973 = ~n_3412 &  n_26972;
assign n_26974 = ~n_3406 &  n_26973;
assign n_26975 = ~n_3400 &  n_26974;
assign n_26976 = ~n_3394 &  n_26975;
assign n_26977 = ~n_3388 &  n_26976;
assign n_26978 = ~n_3382 &  n_26977;
assign n_26979 = ~n_3376 &  n_26978;
assign n_26980 = ~n_3369 &  n_26979;
assign n_26981 = ~n_3363 &  n_26980;
assign n_26982 = ~n_3357 &  n_26981;
assign n_26983 = ~n_3351 &  n_26982;
assign n_26984 = ~n_3345 &  n_26983;
assign n_26985 = ~n_3339 &  n_26984;
assign n_26986 = ~n_3333 &  n_26985;
assign n_26987 = ~n_3327 &  n_26986;
assign n_26988 = ~n_3321 &  n_26987;
assign n_26989 = ~n_3314 &  n_26988;
assign n_26990 = ~n_3239 &  n_26989;
assign n_26991 = ~n_3233 &  n_26990;
assign n_26992 = ~n_3227 &  n_26991;
assign n_26993 = ~n_3221 &  n_26992;
assign n_26994 = ~n_3215 &  n_26993;
assign n_26995 = ~n_3209 &  n_26994;
assign n_26996 = ~n_3203 &  n_26995;
assign n_26997 = ~n_3197 &  n_26996;
assign n_26998 = ~n_3190 &  n_26997;
assign n_26999 = ~n_3184 &  n_26998;
assign n_27000 = ~n_3178 &  n_26999;
assign n_27001 = ~n_3172 &  n_27000;
assign n_27002 = ~n_3166 &  n_27001;
assign n_27003 = ~n_3160 &  n_27002;
assign n_27004 = ~n_3154 &  n_27003;
assign n_27005 = ~n_3148 &  n_27004;
assign n_27006 = ~n_3141 &  n_27005;
assign n_27007 = ~n_3135 &  n_27006;
assign n_27008 = ~n_3129 &  n_27007;
assign n_27009 = ~n_3123 &  n_27008;
assign n_27010 = ~n_3117 &  n_27009;
assign n_27011 = ~n_3111 &  n_27010;
assign n_27012 = ~n_3105 &  n_27011;
assign n_27013 = ~n_3099 &  n_27012;
assign n_27014 = ~n_3092 &  n_27013;
assign n_27015 = ~n_3086 &  n_27014;
assign n_27016 = ~n_3080 &  n_27015;
assign n_27017 = ~n_3074 &  n_27016;
assign n_27018 = ~n_3068 &  n_27017;
assign n_27019 = ~n_3062 &  n_27018;
assign n_27020 = ~n_3056 &  n_27019;
assign n_27021 = ~n_3050 &  n_27020;
assign n_27022 = ~n_3043 &  n_27021;
assign n_27023 = ~n_3037 &  n_27022;
assign n_27024 = ~n_3031 &  n_27023;
assign n_27025 = ~n_3025 &  n_27024;
assign n_27026 = ~n_3019 &  n_27025;
assign n_27027 = ~n_3013 &  n_27026;
assign n_27028 = ~n_3007 &  n_27027;
assign n_27029 = ~n_3001 &  n_27028;
assign n_27030 = ~n_2994 &  n_27029;
assign n_27031 = ~n_2988 &  n_27030;
assign n_27032 = ~n_2982 &  n_27031;
assign n_27033 = ~n_2976 &  n_27032;
assign n_27034 = ~n_2970 &  n_27033;
assign n_27035 = ~n_2964 &  n_27034;
assign n_27036 = ~n_2958 &  n_27035;
assign n_27037 = ~n_2952 &  n_27036;
assign n_27038 = ~n_2945 &  n_27037;
assign n_27039 = ~n_2939 &  n_27038;
assign n_27040 = ~n_2933 &  n_27039;
assign n_27041 = ~n_2927 &  n_27040;
assign n_27042 = ~n_2921 &  n_27041;
assign n_27043 = ~n_2915 &  n_27042;
assign n_27044 = ~n_2909 &  n_27043;
assign n_27045 = ~n_2903 &  n_27044;
assign n_27046 = ~n_2896 &  n_27045;
assign n_27047 = ~n_2890 &  n_27046;
assign n_27048 = ~n_2884 &  n_27047;
assign n_27049 = ~n_2878 &  n_27048;
assign n_27050 = ~n_2872 &  n_27049;
assign n_27051 = ~n_2866 &  n_27050;
assign n_27052 = ~n_2860 &  n_27051;
assign n_27053 = ~n_2854 &  n_27052;
assign n_27054 = ~n_2847 &  n_27053;
assign n_27055 = ~n_2841 &  n_27054;
assign n_27056 = ~n_2835 &  n_27055;
assign n_27057 = ~n_2829 &  n_27056;
assign n_27058 = ~n_2823 &  n_27057;
assign n_27059 = ~n_2817 &  n_27058;
assign n_27060 = ~n_2811 &  n_27059;
assign n_27061 = ~n_2805 &  n_27060;
assign n_27062 = ~n_2798 &  n_27061;
assign n_27063 = ~n_2792 &  n_27062;
assign n_27064 = ~n_2786 &  n_27063;
assign n_27065 = ~n_2780 &  n_27064;
assign n_27066 = ~n_2774 &  n_27065;
assign n_27067 = ~n_2768 &  n_27066;
assign n_27068 = ~n_2762 &  n_27067;
assign n_27069 = ~n_2756 &  n_27068;
assign n_27070 = ~n_2749 &  n_27069;
assign n_27071 = ~n_2743 &  n_27070;
assign n_27072 = ~n_2737 &  n_27071;
assign n_27073 = ~n_2731 &  n_27072;
assign n_27074 = ~n_2725 &  n_27073;
assign n_27075 = ~n_2719 &  n_27074;
assign n_27076 = ~n_2713 &  n_27075;
assign n_27077 = ~n_2707 &  n_27076;
assign n_27078 = ~n_2700 &  n_27077;
assign n_27079 = ~n_2694 &  n_27078;
assign n_27080 = ~n_2688 &  n_27079;
assign n_27081 = ~n_2682 &  n_27080;
assign n_27082 = ~n_2676 &  n_27081;
assign n_27083 = ~n_2670 &  n_27082;
assign n_27084 = ~n_2664 &  n_27083;
assign n_27085 = ~n_2658 &  n_27084;
assign n_27086 = ~n_2651 &  n_27085;
assign n_27087 = ~n_2645 &  n_27086;
assign n_27088 = ~n_2639 &  n_27087;
assign n_27089 = ~n_2633 &  n_27088;
assign n_27090 = ~n_2627 &  n_27089;
assign n_27091 = ~n_2621 &  n_27090;
assign n_27092 = ~n_2615 &  n_27091;
assign n_27093 = ~n_2609 &  n_27092;
assign n_27094 = ~n_2602 &  n_27093;
assign n_27095 = ~n_2596 &  n_27094;
assign n_27096 = ~n_2590 &  n_27095;
assign n_27097 = ~n_2584 &  n_27096;
assign n_27098 = ~n_2578 &  n_27097;
assign n_27099 = ~n_2572 &  n_27098;
assign n_27100 = ~n_2566 &  n_27099;
assign n_27101 = ~n_2560 &  n_27100;
assign n_27102 = ~n_2553 &  n_27101;
assign n_27103 = ~n_2547 &  n_27102;
assign n_27104 = ~n_2541 &  n_27103;
assign n_27105 = ~n_2535 &  n_27104;
assign n_27106 = ~n_2529 &  n_27105;
assign n_27107 = ~n_2523 &  n_27106;
assign n_27108 = ~n_2517 &  n_27107;
assign n_27109 = ~n_2511 &  n_27108;
assign n_27110 = ~n_2504 &  n_27109;
assign n_27111 = ~n_2498 &  n_27110;
assign n_27112 = ~n_2492 &  n_27111;
assign n_27113 = ~n_2486 &  n_27112;
assign n_27114 = ~n_2480 &  n_27113;
assign n_27115 = ~n_2474 &  n_27114;
assign n_27116 = ~n_2468 &  n_27115;
assign n_27117 = ~n_2462 &  n_27116;
assign n_27118 = ~n_2455 &  n_27117;
assign n_27119 = ~n_2449 &  n_27118;
assign n_27120 = ~n_2443 &  n_27119;
assign n_27121 = ~n_2437 &  n_27120;
assign n_27122 = ~n_2431 &  n_27121;
assign n_27123 = ~n_2425 &  n_27122;
assign n_27124 = ~n_2419 &  n_27123;
assign n_27125 = ~n_2413 &  n_27124;
assign n_27126 = ~n_2406 &  n_27125;
assign n_27127 = ~n_2400 &  n_27126;
assign n_27128 = ~n_2394 &  n_27127;
assign n_27129 = ~n_2388 &  n_27128;
assign n_27130 = ~n_2382 &  n_27129;
assign n_27131 = ~n_2376 &  n_27130;
assign n_27132 = ~n_2370 &  n_27131;
assign n_27133 = ~n_2364 &  n_27132;
assign n_27134 = ~n_2357 &  n_27133;
assign n_27135 = ~n_2351 &  n_27134;
assign n_27136 = ~n_2345 &  n_27135;
assign n_27137 = ~n_2339 &  n_27136;
assign n_27138 = ~n_2333 &  n_27137;
assign n_27139 = ~n_2327 &  n_27138;
assign n_27140 = ~n_2321 &  n_27139;
assign n_27141 = ~n_2315 &  n_27140;
assign n_27142 = ~n_2308 &  n_27141;
assign n_27143 = ~n_2302 &  n_27142;
assign n_27144 = ~n_2296 &  n_27143;
assign n_27145 = ~n_2290 &  n_27144;
assign n_27146 = ~n_2284 &  n_27145;
assign n_27147 = ~n_2278 &  n_27146;
assign n_27148 = ~n_2272 &  n_27147;
assign n_27149 = ~n_2266 &  n_27148;
assign n_27150 = ~n_2259 &  n_27149;
assign n_27151 = ~n_2253 &  n_27150;
assign n_27152 = ~n_2247 &  n_27151;
assign n_27153 = ~n_2241 &  n_27152;
assign n_27154 = ~n_2235 &  n_27153;
assign n_27155 = ~n_2229 &  n_27154;
assign n_27156 = ~n_2223 &  n_27155;
assign n_27157 = ~n_2217 &  n_27156;
assign n_27158 = ~n_2210 &  n_27157;
assign n_27159 = ~n_2204 &  n_27158;
assign n_27160 = ~n_2198 &  n_27159;
assign n_27161 = ~n_2192 &  n_27160;
assign n_27162 = ~n_2186 &  n_27161;
assign n_27163 = ~n_2180 &  n_27162;
assign n_27164 = ~n_2174 &  n_27163;
assign n_27165 = ~n_2168 &  n_27164;
assign n_27166 = ~n_2161 &  n_27165;
assign n_27167 = ~n_2155 &  n_27166;
assign n_27168 = ~n_2149 &  n_27167;
assign n_27169 = ~n_2143 &  n_27168;
assign n_27170 = ~n_2137 &  n_27169;
assign n_27171 = ~n_2131 &  n_27170;
assign n_27172 = ~n_2125 &  n_27171;
assign n_27173 = ~n_2119 &  n_27172;
assign n_27174 = ~n_2112 &  n_27173;
assign n_27175 = ~n_2106 &  n_27174;
assign n_27176 = ~n_2100 &  n_27175;
assign n_27177 = ~n_2094 &  n_27176;
assign n_27178 = ~n_2088 &  n_27177;
assign n_27179 = ~n_2082 &  n_27178;
assign n_27180 = ~n_2076 &  n_27179;
assign n_27181 = ~n_2070 &  n_27180;
assign n_27182 = ~n_2063 &  n_27181;
assign n_27183 = ~n_2057 &  n_27182;
assign n_27184 = ~n_2051 &  n_27183;
assign n_27185 = ~n_2045 &  n_27184;
assign n_27186 = ~n_2039 &  n_27185;
assign n_27187 = ~n_2033 &  n_27186;
assign n_27188 = ~n_2027 &  n_27187;
assign n_27189 = ~n_2021 &  n_27188;
assign n_27190 = ~n_2014 &  n_27189;
assign n_27191 = ~n_2008 &  n_27190;
assign n_27192 = ~n_2002 &  n_27191;
assign n_27193 = ~n_1996 &  n_27192;
assign n_27194 = ~n_1990 &  n_27193;
assign n_27195 = ~n_1984 &  n_27194;
assign n_27196 = ~n_1978 &  n_27195;
assign n_27197 = ~n_1972 &  n_27196;
assign n_27198 = ~n_1965 &  n_27197;
assign n_27199 = ~n_1959 &  n_27198;
assign n_27200 = ~n_1953 &  n_27199;
assign n_27201 = ~n_1947 &  n_27200;
assign n_27202 = ~n_1941 &  n_27201;
assign n_27203 = ~n_1935 &  n_27202;
assign n_27204 = ~n_1929 &  n_27203;
assign n_27205 = ~n_1923 &  n_27204;
assign n_27206 = ~n_1916 &  n_27205;
assign n_27207 = ~n_1910 &  n_27206;
assign n_27208 = ~n_1904 &  n_27207;
assign n_27209 = ~n_1898 &  n_27208;
assign n_27210 = ~n_1892 &  n_27209;
assign n_27211 = ~n_1886 &  n_27210;
assign n_27212 = ~n_1880 &  n_27211;
assign n_27213 = ~n_1874 &  n_27212;
assign n_27214 = ~n_1867 &  n_27213;
assign n_27215 = ~n_1861 &  n_27214;
assign n_27216 = ~n_1855 &  n_27215;
assign n_27217 = ~n_1849 &  n_27216;
assign n_27218 = ~n_1843 &  n_27217;
assign n_27219 = ~n_1837 &  n_27218;
assign n_27220 = ~n_1831 &  n_27219;
assign n_27221 = ~n_1825 &  n_27220;
assign n_27222 = ~n_1818 &  n_27221;
assign n_27223 = ~n_1812 &  n_27222;
assign n_27224 = ~n_1805 &  n_27223;
assign n_27225 = ~n_1798 &  n_27224;
assign n_27226 = ~n_1791 &  n_27225;
assign n_27227 = ~n_1784 &  n_27226;
assign n_27228 = ~n_1776 &  n_27227;
assign n_27229 = ~n_1768 &  n_27228;
assign n_27230 = ~n_1758 &  n_27229;
assign n_27231 = ~n_1747 &  n_27230;
assign n_27232 = ~n_1744 &  n_27231;
assign n_27233 = ~n_1738 &  n_27232;
assign n_27234 = ~n_1735 &  n_27233;
assign n_27235 = ~n_1730 &  n_27234;
assign n_27236 = ~n_1727 &  n_27235;
assign n_27237 = ~n_1722 &  n_27236;
assign n_27238 = ~n_1711 &  n_27237;
assign n_27239 = ~n_1705 &  n_27238;
assign n_27240 = ~n_1699 &  n_27239;
assign n_27241 = ~n_1693 &  n_27240;
assign n_27242 = ~n_1687 &  n_27241;
assign n_27243 = ~n_1681 &  n_27242;
assign n_27244 = ~n_1675 &  n_27243;
assign n_27245 = ~n_1669 &  n_27244;
assign n_27246 = ~n_1663 &  n_27245;
assign n_27247 = ~n_1657 &  n_27246;
assign n_27248 = ~n_1651 &  n_27247;
assign n_27249 = ~n_1645 &  n_27248;
assign n_27250 = ~n_1639 &  n_27249;
assign n_27251 = ~n_1633 &  n_27250;
assign n_27252 = ~n_1627 &  n_27251;
assign n_27253 = ~n_1621 &  n_27252;
assign n_27254 = ~n_1615 &  n_27253;
assign n_27255 = ~n_1609 &  n_27254;
assign n_27256 = ~n_1603 &  n_27255;
assign n_27257 = ~n_1597 &  n_27256;
assign n_27258 = ~n_1591 &  n_27257;
assign n_27259 = ~n_1585 &  n_27258;
assign n_27260 = ~n_1579 &  n_27259;
assign n_27261 = ~n_1573 &  n_27260;
assign n_27262 = ~n_1567 &  n_27261;
assign n_27263 = ~n_1561 &  n_27262;
assign n_27264 = ~n_1555 &  n_27263;
assign n_27265 = ~n_1549 &  n_27264;
assign n_27266 = ~n_1543 &  n_27265;
assign n_27267 = ~n_1537 &  n_27266;
assign n_27268 = ~n_1531 &  n_27267;
assign n_27269 = ~n_1521 &  n_27268;
assign n_27270 = ~n_1518 &  n_27269;
assign n_27271 = ~n_1515 &  n_27270;
assign n_27272 = ~n_1512 &  n_27271;
assign n_27273 = ~n_1496 &  n_27272;
assign n_27274 = ~n_1490 &  n_27273;
assign n_27275 = ~n_1484 &  n_27274;
assign n_27276 = ~n_1478 &  n_27275;
assign n_27277 = ~n_1472 &  n_27276;
assign n_27278 = ~n_1466 &  n_27277;
assign n_27279 = ~n_1460 &  n_27278;
assign n_27280 = ~n_1454 &  n_27279;
assign n_27281 = ~n_1448 &  n_27280;
assign n_27282 = ~n_1442 &  n_27281;
assign n_27283 = ~n_1436 &  n_27282;
assign n_27284 = ~n_1430 &  n_27283;
assign n_27285 = ~n_1424 &  n_27284;
assign n_27286 = ~n_1418 &  n_27285;
assign n_27287 = ~n_1412 &  n_27286;
assign n_27288 = ~n_1406 &  n_27287;
assign n_27289 = ~n_1400 &  n_27288;
assign n_27290 = ~n_1394 &  n_27289;
assign n_27291 = ~n_1388 &  n_27290;
assign n_27292 = ~n_1382 &  n_27291;
assign n_27293 = ~n_1376 &  n_27292;
assign n_27294 = ~n_1370 &  n_27293;
assign n_27295 = ~n_1364 &  n_27294;
assign n_27296 = ~n_1358 &  n_27295;
assign n_27297 = ~n_1352 &  n_27296;
assign n_27298 = ~n_1346 &  n_27297;
assign n_27299 = ~n_1340 &  n_27298;
assign n_27300 = ~n_1334 &  n_27299;
assign n_27301 = ~n_1324 &  n_27300;
assign n_27302 = ~n_1320 &  n_27301;
assign n_27303 = ~n_1317 &  n_27302;
assign n_27304 = ~n_1314 &  n_27303;
assign n_27305 = ~n_1311 &  n_27304;
assign n_27306 = ~n_1306 &  n_27305;
assign n_27307 = ~n_1303 &  n_27306;
assign n_27308 = ~n_1297 &  n_27307;
assign n_27309 = ~n_1275 &  n_27308;
assign n_27310 = ~n_1272 &  n_27309;
assign n_27311 = ~n_1269 &  n_27310;
assign n_27312 = ~n_1265 &  n_27311;
assign n_27313 = ~n_1261 &  n_27312;
assign n_27314 = ~n_1247 &  n_27313;
assign n_27315 = ~n_1244 &  n_27314;
assign n_27316 = ~n_1241 &  n_27315;
assign n_27317 = ~n_1238 &  n_27316;
assign n_27318 = ~n_1235 &  n_27317;
assign n_27319 = ~n_1232 &  n_27318;
assign n_27320 = ~n_1229 &  n_27319;
assign n_27321 = ~n_1223 &  n_27320;
assign n_27322 = ~n_1214 &  n_27321;
assign n_27323 = ~n_1207 &  n_27322;
assign n_27324 = ~n_1201 &  n_27323;
assign n_27325 = ~n_1198 &  n_27324;
assign n_27326 = ~n_1177 &  n_27325;
assign n_27327 = ~n_1169 &  n_27326;
assign n_27328 = ~n_1163 &  n_27327;
assign n_27329 = ~n_1142 &  n_27328;
assign n_27330 = ~n_1132 &  n_27329;
assign n_27331 = ~n_1125 &  n_27330;
assign n_27332 = ~n_1104 &  n_27331;
assign n_27333 = ~n_1095 &  n_27332;
assign n_27334 = ~n_1074 &  n_27333;
assign n_27335 = ~n_1065 &  n_27334;
assign n_27336 = ~n_1044 &  n_27335;
assign n_27337 = ~n_1035 &  n_27336;
assign n_27338 = ~n_1014 &  n_27337;
assign n_27339 = ~n_1005 &  n_27338;
assign n_27340 = ~n_984 &  n_27339;
assign n_27341 = ~n_975 &  n_27340;
assign n_27342 = ~n_954 &  n_27341;
assign n_27343 = ~n_945 &  n_27342;
assign n_27344 = ~n_922 &  n_27343;
assign n_27345 = ~n_912 &  n_27344;
assign n_27346 = ~n_905 &  n_27345;
assign n_27347 = ~n_899 &  n_27346;
assign n_27348 = ~n_893 &  n_27347;
assign n_27349 = ~n_887 &  n_27348;
assign n_27350 = ~n_881 &  n_27349;
assign n_27351 = ~n_875 &  n_27350;
assign n_27352 = ~n_869 &  n_27351;
assign n_27353 = ~n_863 &  n_27352;
assign n_27354 = ~n_856 &  n_27353;
assign n_27355 = ~n_850 &  n_27354;
assign n_27356 = ~n_844 &  n_27355;
assign n_27357 = ~n_838 &  n_27356;
assign n_27358 = ~n_832 &  n_27357;
assign n_27359 = ~n_826 &  n_27358;
assign n_27360 = ~n_820 &  n_27359;
assign n_27361 = ~n_814 &  n_27360;
assign n_27362 = ~n_807 &  n_27361;
assign n_27363 = ~n_801 &  n_27362;
assign n_27364 = ~n_795 &  n_27363;
assign n_27365 = ~n_789 &  n_27364;
assign n_27366 = ~n_783 &  n_27365;
assign n_27367 = ~n_777 &  n_27366;
assign n_27368 = ~n_771 &  n_27367;
assign n_27369 = ~n_765 &  n_27368;
assign n_27370 = ~n_758 &  n_27369;
assign n_27371 = ~n_752 &  n_27370;
assign n_27372 = ~n_746 &  n_27371;
assign n_27373 = ~n_740 &  n_27372;
assign n_27374 = ~n_734 &  n_27373;
assign n_27375 = ~n_728 &  n_27374;
assign n_27376 = ~n_722 &  n_27375;
assign n_27377 = ~n_716 &  n_27376;
assign n_27378 = ~n_709 &  n_27377;
assign n_27379 = ~n_703 &  n_27378;
assign n_27380 = ~n_697 &  n_27379;
assign n_27381 = ~n_691 &  n_27380;
assign n_27382 = ~n_685 &  n_27381;
assign n_27383 = ~n_679 &  n_27382;
assign n_27384 = ~n_673 &  n_27383;
assign n_27385 = ~n_667 &  n_27384;
assign n_27386 = ~n_660 &  n_27385;
assign n_27387 = ~n_654 &  n_27386;
assign n_27388 = ~n_648 &  n_27387;
assign n_27389 = ~n_642 &  n_27388;
assign n_27390 = ~n_636 &  n_27389;
assign n_27391 = ~n_630 &  n_27390;
assign n_27392 = ~n_624 &  n_27391;
assign n_27393 = ~n_618 &  n_27392;
assign n_27394 = ~n_577 &  n_27393;
assign n_27395 = ~n_571 &  n_27394;
assign n_27396 = ~n_565 &  n_27395;
assign n_27397 = ~n_559 &  n_27396;
assign n_27398 = ~n_553 &  n_27397;
assign n_27399 = ~n_547 &  n_27398;
assign n_27400 = ~n_541 &  n_27399;
assign n_27401 = ~n_530 &  n_27400;
assign n_27402 = ~n_527 &  n_27401;
assign n_27403 = ~n_522 &  n_27402;
assign n_27404 = ~n_519 &  n_27403;
assign n_27405 = ~n_516 &  n_27404;
assign n_27406 = ~n_513 &  n_27405;
assign n_27407 = ~n_435 &  n_27406;
assign n_27408 = ~n_417 &  n_27407;
assign n_27409 = ~n_399 &  n_27408;
assign n_27410 = ~n_381 &  n_27409;
assign n_27411 = ~n_363 &  n_27410;
assign n_27412 = ~n_345 &  n_27411;
assign n_27413 = ~n_327 &  n_27412;
assign n_27414 = ~n_309 &  n_27413;
assign n_27415 = ~n_291 &  n_27414;
assign n_27416 = ~n_273 &  n_27415;
assign n_27417 = ~n_255 &  n_27416;
assign n_27418 = ~n_237 &  n_27417;
assign n_27419 = ~n_219 &  n_27418;
assign n_27420 = ~n_201 &  n_27419;
assign n_27421 = ~n_183 &  n_27420;
assign n_27422 = ~n_165 &  n_27421;
assign n_27423 = ~n_147 &  n_27422;
assign n_27424 = ~n_129 &  n_27423;
assign n_27425 = ~n_111 &  n_27424;
assign n_27426 = ~n_93 &  n_27425;
assign n_27427 = ~n_75 &  n_27426;
assign n_27428 = ~n_57 &  n_27427;
assign n_27429 = ~n_39 &  n_27428;
assign o_1 = ~n_27429;
endmodule

