module formula(v_185,v_186,v_187,v_188,v_189,v_190,v_191,v_192,v_193,v_194,v_195,v_196,v_197,v_198,v_199,v_200,v_201,v_202,v_203,v_204,v_205,v_206,v_207,v_208,v_209,v_210,v_211,v_212,v_213,v_214,v_215,v_216,v_217,v_218,v_219,v_220,v_221,v_222,v_223,v_224,v_225,v_226,v_227,v_228,v_229,v_230,v_231,v_232,v_233,v_234,v_235,v_236,v_237,v_238,v_239,v_240,v_241,v_242,v_243,v_244,v_245,v_246,v_247,v_248,v_184,v_249,v_250,v_251,v_252,v_253,v_254,v_255,v_256,v_257,v_258,v_259,v_260,v_261,v_262,v_263,v_264,v_265,v_266,v_267,v_268,v_269,v_270,v_271,v_272,v_273,v_274,v_275,v_276,v_277,v_278,v_7,v_8,v_9,v_10,v_11,v_12,v_13,v_14,v_15,v_16,v_17,v_18,v_19,v_20,v_21,v_22,v_23,v_24,v_25,v_26,v_27,v_28,v_29,v_30,v_31,v_32,v_33,v_34,v_35,v_36,v_37,v_38,v_39,v_40,v_41,v_42,v_43,v_44,v_45,v_46,v_47,v_48,v_49,v_50,v_51,v_52,v_53,v_54,v_55,v_56,v_57,v_60,v_61,v_64,v_69,v_70,o_1);
	input v_185;
	input v_186;
	input v_187;
	input v_188;
	input v_189;
	input v_190;
	input v_191;
	input v_192;
	input v_193;
	input v_194;
	input v_195;
	input v_196;
	input v_197;
	input v_198;
	input v_199;
	input v_200;
	input v_201;
	input v_202;
	input v_203;
	input v_204;
	input v_205;
	input v_206;
	input v_207;
	input v_208;
	input v_209;
	input v_210;
	input v_211;
	input v_212;
	input v_213;
	input v_214;
	input v_215;
	input v_216;
	input v_217;
	input v_218;
	input v_219;
	input v_220;
	input v_221;
	input v_222;
	input v_223;
	input v_224;
	input v_225;
	input v_226;
	input v_227;
	input v_228;
	input v_229;
	input v_230;
	input v_231;
	input v_232;
	input v_233;
	input v_234;
	input v_235;
	input v_236;
	input v_237;
	input v_238;
	input v_239;
	input v_240;
	input v_241;
	input v_242;
	input v_243;
	input v_244;
	input v_245;
	input v_246;
	input v_247;
	input v_248;
	input v_184;
	input v_249;
	input v_250;
	input v_251;
	input v_252;
	input v_253;
	input v_254;
	input v_255;
	input v_256;
	input v_257;
	input v_258;
	input v_259;
	input v_260;
	input v_261;
	input v_262;
	input v_263;
	input v_264;
	input v_265;
	input v_266;
	input v_267;
	input v_268;
	input v_269;
	input v_270;
	input v_271;
	input v_272;
	input v_273;
	input v_274;
	input v_275;
	input v_276;
	input v_277;
	input v_278;
	input v_7;
	input v_8;
	input v_9;
	input v_10;
	input v_11;
	input v_12;
	input v_13;
	input v_14;
	input v_15;
	input v_16;
	input v_17;
	input v_18;
	input v_19;
	input v_20;
	input v_21;
	input v_22;
	input v_23;
	input v_24;
	input v_25;
	input v_26;
	input v_27;
	input v_28;
	input v_29;
	input v_30;
	input v_31;
	input v_32;
	input v_33;
	input v_34;
	input v_35;
	input v_36;
	input v_37;
	input v_38;
	input v_39;
	input v_40;
	input v_41;
	input v_42;
	input v_43;
	input v_44;
	input v_45;
	input v_46;
	input v_47;
	input v_48;
	input v_49;
	input v_50;
	input v_51;
	input v_52;
	input v_53;
	input v_54;
	input v_55;
	input v_56;
	input v_57;
	input v_60;
	input v_61;
	input v_64;
	input v_69;
	input v_70;
	wire v_1;
	wire v_2;
	wire v_3;
	wire v_4;
	wire v_5;
	wire v_6;
	wire v_58;
	wire v_59;
	wire v_62;
	wire v_63;
	wire v_65;
	wire v_66;
	wire v_67;
	wire v_68;
	wire v_71;
	wire v_72;
	wire v_73;
	wire v_74;
	wire v_75;
	wire v_76;
	wire v_77;
	wire v_78;
	wire v_79;
	wire v_80;
	wire v_81;
	wire v_82;
	wire v_83;
	wire v_84;
	wire v_85;
	wire v_86;
	wire v_87;
	wire v_88;
	wire v_89;
	wire v_90;
	wire v_91;
	wire v_92;
	wire v_93;
	wire v_94;
	wire v_95;
	wire v_96;
	wire v_97;
	wire v_98;
	wire v_99;
	wire v_100;
	wire v_101;
	wire v_102;
	wire v_103;
	wire v_104;
	wire v_105;
	wire v_106;
	wire v_107;
	wire v_108;
	wire v_109;
	wire v_110;
	wire v_111;
	wire v_112;
	wire v_113;
	wire v_114;
	wire v_115;
	wire v_116;
	wire v_117;
	wire v_118;
	wire v_119;
	wire v_120;
	wire v_121;
	wire v_122;
	wire v_123;
	wire v_124;
	wire v_125;
	wire v_126;
	wire v_127;
	wire v_128;
	wire v_129;
	wire v_130;
	wire v_131;
	wire v_132;
	wire v_133;
	wire v_134;
	wire v_135;
	wire v_136;
	wire v_137;
	wire v_138;
	wire v_139;
	wire v_140;
	wire v_141;
	wire v_142;
	wire v_143;
	wire v_144;
	wire v_145;
	wire v_146;
	wire v_147;
	wire v_148;
	wire v_149;
	wire v_150;
	wire v_151;
	wire v_152;
	wire v_153;
	wire v_154;
	wire v_155;
	wire v_156;
	wire v_157;
	wire v_158;
	wire v_159;
	wire v_160;
	wire v_161;
	wire v_162;
	wire v_163;
	wire v_164;
	wire v_165;
	wire v_166;
	wire v_167;
	wire v_168;
	wire v_169;
	wire v_170;
	wire v_171;
	wire v_172;
	wire v_173;
	wire v_174;
	wire v_175;
	wire v_176;
	wire v_177;
	wire v_178;
	wire v_179;
	wire v_180;
	wire v_181;
	wire v_182;
	wire v_183;
	wire v_279;
	wire x_1;
	wire x_2;
	wire x_3;
	wire x_4;
	wire x_5;
	wire x_6;
	wire x_7;
	wire x_8;
	wire x_9;
	wire x_10;
	wire x_11;
	wire x_12;
	wire x_13;
	wire x_14;
	wire x_15;
	wire x_16;
	wire x_17;
	wire x_18;
	wire x_19;
	wire x_20;
	wire x_21;
	wire x_22;
	wire x_23;
	wire x_24;
	wire x_25;
	wire x_26;
	wire x_27;
	wire x_28;
	wire x_29;
	wire x_30;
	wire x_31;
	wire x_32;
	wire x_33;
	wire x_34;
	wire x_35;
	wire x_36;
	wire x_37;
	wire x_38;
	wire x_39;
	wire x_40;
	wire x_41;
	wire x_42;
	wire x_43;
	wire x_44;
	wire x_45;
	wire x_46;
	wire x_47;
	wire x_48;
	wire x_49;
	wire x_50;
	wire x_51;
	wire x_52;
	wire x_53;
	wire x_54;
	wire x_55;
	wire x_56;
	wire x_57;
	wire x_58;
	wire x_59;
	wire x_60;
	wire x_61;
	wire x_62;
	wire x_63;
	wire x_64;
	wire x_65;
	wire x_66;
	wire x_67;
	wire x_68;
	wire x_69;
	wire x_70;
	wire x_71;
	wire x_72;
	wire x_73;
	wire x_74;
	wire x_75;
	wire x_76;
	wire x_77;
	wire x_78;
	wire x_79;
	wire x_80;
	wire x_81;
	wire x_82;
	wire x_83;
	wire x_84;
	wire x_85;
	wire x_86;
	wire x_87;
	wire x_88;
	wire x_89;
	wire x_90;
	wire x_91;
	wire x_92;
	wire x_93;
	wire x_94;
	wire x_95;
	wire x_96;
	wire x_97;
	wire x_98;
	wire x_99;
	wire x_100;
	wire x_101;
	wire x_102;
	wire x_103;
	wire x_104;
	wire x_105;
	wire x_106;
	wire x_107;
	wire x_108;
	wire x_109;
	wire x_110;
	wire x_111;
	wire x_112;
	wire x_113;
	wire x_114;
	wire x_115;
	wire x_116;
	wire x_117;
	wire x_118;
	wire x_119;
	wire x_120;
	wire x_121;
	wire x_122;
	wire x_123;
	wire x_124;
	wire x_125;
	wire x_126;
	wire x_127;
	wire x_128;
	wire x_129;
	wire x_130;
	wire x_131;
	wire x_132;
	wire x_133;
	wire x_134;
	wire x_135;
	wire x_136;
	wire x_137;
	wire x_138;
	wire x_139;
	wire x_140;
	wire x_141;
	wire x_142;
	wire x_143;
	wire x_144;
	wire x_145;
	wire x_146;
	wire x_147;
	wire x_148;
	wire x_149;
	wire x_150;
	wire x_151;
	wire x_152;
	wire x_153;
	wire x_154;
	wire x_155;
	wire x_156;
	wire x_157;
	wire x_158;
	wire x_159;
	wire x_160;
	wire x_161;
	wire x_162;
	wire x_163;
	wire x_164;
	wire x_165;
	wire x_166;
	wire x_167;
	wire x_168;
	wire x_169;
	wire x_170;
	wire x_171;
	wire x_172;
	wire x_173;
	wire x_174;
	wire x_175;
	wire x_176;
	wire x_177;
	wire x_178;
	wire x_179;
	wire x_180;
	wire x_181;
	wire x_182;
	wire x_183;
	wire x_184;
	wire x_185;
	wire x_186;
	wire x_187;
	wire x_188;
	wire x_189;
	wire x_190;
	wire x_191;
	wire x_192;
	wire x_193;
	wire x_194;
	wire x_195;
	wire x_196;
	wire x_197;
	wire x_198;
	wire x_199;
	wire x_200;
	wire x_201;
	wire x_202;
	wire x_203;
	wire x_204;
	wire x_205;
	wire x_206;
	wire x_207;
	wire x_208;
	wire x_209;
	wire x_210;
	wire x_211;
	wire x_212;
	wire x_213;
	wire x_214;
	wire x_215;
	wire x_216;
	wire x_217;
	wire x_218;
	wire x_219;
	wire x_220;
	wire x_221;
	wire x_222;
	wire x_223;
	wire x_224;
	wire x_225;
	wire x_226;
	wire x_227;
	wire x_228;
	wire x_229;
	wire x_230;
	wire x_231;
	wire x_232;
	wire x_233;
	wire x_234;
	wire x_235;
	wire x_236;
	wire x_237;
	wire x_238;
	wire x_239;
	wire x_240;
	wire x_241;
	wire x_242;
	wire x_243;
	wire x_244;
	wire x_245;
	wire x_246;
	wire x_247;
	wire x_248;
	wire x_249;
	wire x_250;
	wire x_251;
	wire x_252;
	wire x_253;
	wire x_254;
	wire x_255;
	wire x_256;
	wire x_257;
	wire x_258;
	wire x_259;
	wire x_260;
	wire x_261;
	wire x_262;
	wire x_263;
	wire x_264;
	wire x_265;
	wire x_266;
	wire x_267;
	wire x_268;
	wire x_269;
	wire x_270;
	wire x_271;
	wire x_272;
	wire x_273;
	wire x_274;
	wire x_275;
	wire x_276;
	wire x_277;
	wire x_278;
	wire x_279;
	wire x_280;
	wire x_281;
	wire x_282;
	wire x_283;
	wire x_284;
	wire x_285;
	wire x_286;
	wire x_287;
	wire x_288;
	wire x_289;
	wire x_290;
	wire x_291;
	wire x_292;
	wire x_293;
	wire x_294;
	wire x_295;
	wire x_296;
	wire x_297;
	wire x_298;
	wire x_299;
	wire x_300;
	wire x_301;
	wire x_302;
	wire x_303;
	wire x_304;
	wire x_305;
	wire x_306;
	wire x_307;
	wire x_308;
	wire x_309;
	wire x_310;
	wire x_311;
	wire x_312;
	wire x_313;
	wire x_314;
	wire x_315;
	wire x_316;
	wire x_317;
	wire x_318;
	wire x_319;
	wire x_320;
	wire x_321;
	wire x_322;
	wire x_323;
	wire x_324;
	wire x_325;
	wire x_326;
	wire x_327;
	wire x_328;
	wire x_329;
	wire x_330;
	wire x_331;
	wire x_332;
	wire x_333;
	wire x_334;
	wire x_335;
	wire x_336;
	wire x_337;
	wire x_338;
	wire x_339;
	wire x_340;
	wire x_341;
	wire x_342;
	wire x_343;
	wire x_344;
	wire x_345;
	wire x_346;
	wire x_347;
	wire x_348;
	wire x_349;
	wire x_350;
	wire x_351;
	wire x_352;
	wire x_353;
	wire x_354;
	wire x_355;
	wire x_356;
	wire x_357;
	wire x_358;
	wire x_359;
	wire x_360;
	wire x_361;
	wire x_362;
	wire x_363;
	wire x_364;
	wire x_365;
	wire x_366;
	wire x_367;
	wire x_368;
	wire x_369;
	wire x_370;
	wire x_371;
	wire x_372;
	wire x_373;
	wire x_374;
	wire x_375;
	wire x_376;
	wire x_377;
	wire x_378;
	wire x_379;
	wire x_380;
	wire x_381;
	wire x_382;
	wire x_383;
	wire x_384;
	wire x_385;
	wire x_386;
	wire x_387;
	wire x_388;
	wire x_389;
	wire x_390;
	wire x_391;
	wire x_392;
	wire x_393;
	wire x_394;
	wire x_395;
	wire x_396;
	wire x_397;
	wire x_398;
	wire x_399;
	wire x_400;
	wire x_401;
	wire x_402;
	wire x_403;
	wire x_404;
	wire x_405;
	wire x_406;
	wire x_407;
	wire x_408;
	wire x_409;
	wire x_410;
	wire x_411;
	wire x_412;
	wire x_413;
	wire x_414;
	wire x_415;
	wire x_416;
	wire x_417;
	wire x_418;
	wire x_419;
	wire x_420;
	wire x_421;
	wire x_422;
	wire x_423;
	wire x_424;
	wire x_425;
	wire x_426;
	wire x_427;
	wire x_428;
	wire x_429;
	wire x_430;
	wire x_431;
	wire x_432;
	wire x_433;
	wire x_434;
	wire x_435;
	wire x_436;
	wire x_437;
	wire x_438;
	wire x_439;
	wire x_440;
	wire x_441;
	wire x_442;
	wire x_443;
	wire x_444;
	wire x_445;
	wire x_446;
	wire x_447;
	wire x_448;
	wire x_449;
	wire x_450;
	wire x_451;
	wire x_452;
	wire x_453;
	wire x_454;
	wire x_455;
	wire x_456;
	wire x_457;
	wire x_458;
	wire x_459;
	wire x_460;
	wire x_461;
	wire x_462;
	wire x_463;
	wire x_464;
	wire x_465;
	wire x_466;
	wire x_467;
	wire x_468;
	wire x_469;
	wire x_470;
	wire x_471;
	wire x_472;
	wire x_473;
	wire x_474;
	wire x_475;
	wire x_476;
	wire x_477;
	wire x_478;
	wire x_479;
	wire x_480;
	wire x_481;
	wire x_482;
	wire x_483;
	wire x_484;
	wire x_485;
	wire x_486;
	wire x_487;
	wire x_488;
	wire x_489;
	wire x_490;
	wire x_491;
	wire x_492;
	wire x_493;
	wire x_494;
	wire x_495;
	wire x_496;
	wire x_497;
	wire x_498;
	wire x_499;
	wire x_500;
	wire x_501;
	wire x_502;
	wire x_503;
	wire x_504;
	wire x_505;
	wire x_506;
	wire x_507;
	wire x_508;
	wire x_509;
	wire x_510;
	wire x_511;
	wire x_512;
	wire x_513;
	wire x_514;
	wire x_515;
	wire x_516;
	wire x_517;
	wire x_518;
	wire x_519;
	wire x_520;
	wire x_521;
	wire x_522;
	wire x_523;
	wire x_524;
	wire x_525;
	wire x_526;
	wire x_527;
	wire x_528;
	wire x_529;
	wire x_530;
	wire x_531;
	wire x_532;
	wire x_533;
	wire x_534;
	wire x_535;
	wire x_536;
	wire x_537;
	wire x_538;
	wire x_539;
	wire x_540;
	wire x_541;
	wire x_542;
	wire x_543;
	wire x_544;
	wire x_545;
	wire x_546;
	wire x_547;
	wire x_548;
	wire x_549;
	wire x_550;
	wire x_551;
	wire x_552;
	wire x_553;
	wire x_554;
	wire x_555;
	wire x_556;
	wire x_557;
	wire x_558;
	wire x_559;
	wire x_560;
	wire x_561;
	wire x_562;
	wire x_563;
	wire x_564;
	wire x_565;
	wire x_566;
	wire x_567;
	wire x_568;
	wire x_569;
	wire x_570;
	wire x_571;
	wire x_572;
	wire x_573;
	wire x_574;
	wire x_575;
	wire x_576;
	wire x_577;
	wire x_578;
	wire x_579;
	wire x_580;
	wire x_581;
	wire x_582;
	wire x_583;
	wire x_584;
	wire x_585;
	wire x_586;
	wire x_587;
	wire x_588;
	wire x_589;
	wire x_590;
	wire x_591;
	wire x_592;
	wire x_593;
	wire x_594;
	wire x_595;
	wire x_596;
	wire x_597;
	wire x_598;
	wire x_599;
	wire x_600;
	wire x_601;
	wire x_602;
	wire x_603;
	wire x_604;
	wire x_605;
	wire x_606;
	wire x_607;
	wire x_608;
	wire x_609;
	wire x_610;
	wire x_611;
	wire x_612;
	wire x_613;
	wire x_614;
	wire x_615;
	wire x_616;
	wire x_617;
	wire x_618;
	wire x_619;
	wire x_620;
	wire x_621;
	wire x_622;
	wire x_623;
	wire x_624;
	wire x_625;
	wire x_626;
	wire x_627;
	wire x_628;
	wire x_629;
	wire x_630;
	wire x_631;
	wire x_632;
	wire x_633;
	wire x_634;
	wire x_635;
	wire x_636;
	wire x_637;
	wire x_638;
	wire x_639;
	wire x_640;
	wire x_641;
	wire x_642;
	wire x_643;
	wire x_644;
	wire x_645;
	wire x_646;
	wire x_647;
	wire x_648;
	wire x_649;
	wire x_650;
	wire x_651;
	wire x_652;
	wire x_653;
	wire x_654;
	wire x_655;
	wire x_656;
	wire x_657;
	wire x_658;
	wire x_659;
	wire x_660;
	wire x_661;
	wire x_662;
	wire x_663;
	wire x_664;
	wire x_665;
	wire x_666;
	wire x_667;
	wire x_668;
	wire x_669;
	wire x_670;
	wire x_671;
	wire x_672;
	wire x_673;
	wire x_674;
	wire x_675;
	wire x_676;
	wire x_677;
	wire x_678;
	wire x_679;
	wire x_680;
	wire x_681;
	wire x_682;
	wire x_683;
	wire x_684;
	wire x_685;
	wire x_686;
	wire x_687;
	wire x_688;
	wire x_689;
	wire x_690;
	wire x_691;
	wire x_692;
	wire x_693;
	wire x_694;
	wire x_695;
	wire x_696;
	wire x_697;
	wire x_698;
	wire x_699;
	wire x_700;
	wire x_701;
	wire x_702;
	wire x_703;
	wire x_704;
	wire x_705;
	wire x_706;
	wire x_707;
	wire x_708;
	wire x_709;
	wire x_710;
	wire x_711;
	wire x_712;
	wire x_713;
	wire x_714;
	wire x_715;
	wire x_716;
	wire x_717;
	wire x_718;
	wire x_719;
	wire x_720;
	wire x_721;
	wire x_722;
	wire x_723;
	wire x_724;
	wire x_725;
	wire x_726;
	wire x_727;
	wire x_728;
	wire x_729;
	wire x_730;
	wire x_731;
	wire x_732;
	wire x_733;
	wire x_734;
	wire x_735;
	wire x_736;
	wire x_737;
	wire x_738;
	wire x_739;
	wire x_740;
	wire x_741;
	wire x_742;
	wire x_743;
	wire x_744;
	wire x_745;
	wire x_746;
	wire x_747;
	wire x_748;
	wire x_749;
	wire x_750;
	wire x_751;
	wire x_752;
	wire x_753;
	output o_1;
	assign v_65 = (v_241 ^ v_242) ;
	assign v_165 = v_277 ;
	assign v_66 = (v_237 ^ v_238) ;
	assign v_159 = v_275 ;
	assign v_168 = (v_245 & v_246) ;
	assign v_167 = v_278 ;
	assign v_162 = v_276 ;
	assign v_156 = v_274 ;
	assign v_153 = v_273 ;
	assign v_149 = v_272 ;
	assign v_146 = v_271 ;
	assign v_143 = v_270 ;
	assign v_139 = v_269 ;
	assign v_136 = v_268 ;
	assign v_133 = v_267 ;
	assign v_129 = v_266 ;
	assign v_126 = v_265 ;
	assign v_123 = v_264 ;
	assign v_119 = v_263 ;
	assign v_116 = v_262 ;
	assign v_113 = v_261 ;
	assign v_109 = v_260 ;
	assign v_106 = v_259 ;
	assign v_102 = v_258 ;
	assign v_99 = v_257 ;
	assign v_95 = v_256 ;
	assign v_92 = v_255 ;
	assign v_88 = v_254 ;
	assign v_85 = v_253 ;
	assign v_81 = v_252 ;
	assign v_78 = v_251 ;
	assign v_74 = v_250 ;
	assign v_71 = ~v_69 ;
	assign v_6 = v_249 ;
	assign v_63 = (v_165 ^ ~v_65) ;
	assign v_59 = (v_159 ^ ~v_66) ;
	assign v_169 = (v_167 ^ v_168) ;
	assign v_163 = (v_162 ^ ~v_61) ;
	assign v_157 = (v_156 ^ ~v_57) ;
	assign v_154 = (v_153 ^ ~v_55) ;
	assign v_150 = (v_149 ^ ~v_53) ;
	assign v_147 = (v_146 ^ ~v_51) ;
	assign v_144 = (v_143 ^ ~v_49) ;
	assign v_140 = (v_139 ^ ~v_47) ;
	assign v_137 = (v_136 ^ ~v_45) ;
	assign v_134 = (v_133 ^ ~v_43) ;
	assign v_130 = (v_129 ^ ~v_41) ;
	assign v_127 = (v_126 ^ ~v_39) ;
	assign v_124 = (v_123 ^ ~v_37) ;
	assign v_120 = (v_119 ^ ~v_35) ;
	assign v_117 = (v_116 ^ ~v_33) ;
	assign v_114 = (v_113 ^ ~v_31) ;
	assign v_110 = (v_109 ^ ~v_29) ;
	assign v_107 = (v_106 ^ ~v_27) ;
	assign v_103 = (v_102 ^ ~v_25) ;
	assign v_100 = (v_99 ^ ~v_23) ;
	assign v_96 = (v_95 ^ ~v_21) ;
	assign v_93 = (v_92 ^ ~v_19) ;
	assign v_89 = (v_88 ^ ~v_17) ;
	assign v_86 = (v_85 ^ ~v_15) ;
	assign v_82 = (v_81 ^ ~v_13) ;
	assign v_79 = (v_78 ^ ~v_11) ;
	assign v_75 = (v_74 ^ ~v_9) ;
	assign v_72 = (v_71 ^ v_184) ;
	assign v_67 = (v_6 ^ ~v_7) ;
	assign v_62 = (~v_63 & v_65) ;
	assign v_58 = (~v_59 & v_66) ;
	assign x_377 = ((~v_169 | v_243) | v_244) ;
	assign x_376 = ((~v_169 | ~v_243) | ~v_244) ;
	assign x_374 = ((v_169 | v_243) | ~v_244) ;
	assign x_373 = ((~v_163 | v_239) | v_240) ;
	assign x_371 = ((v_163 | ~v_239) | v_240) ;
	assign x_370 = ((v_163 | v_239) | ~v_240) ;
	assign x_368 = ((~v_157 | ~v_235) | ~v_236) ;
	assign x_367 = ((v_157 | ~v_235) | v_236) ;
	assign x_365 = ((~v_154 | v_233) | v_234) ;
	assign x_364 = ((~v_154 | ~v_233) | ~v_234) ;
	assign x_362 = ((v_154 | v_233) | ~v_234) ;
	assign x_361 = ((~v_150 | v_231) | v_232) ;
	assign x_359 = ((v_150 | ~v_231) | v_232) ;
	assign x_358 = ((v_150 | v_231) | ~v_232) ;
	assign x_356 = ((~v_147 | ~v_229) | ~v_230) ;
	assign x_355 = ((v_147 | ~v_229) | v_230) ;
	assign x_353 = ((~v_144 | v_227) | v_228) ;
	assign x_352 = ((~v_144 | ~v_227) | ~v_228) ;
	assign x_350 = ((v_144 | v_227) | ~v_228) ;
	assign x_349 = ((~v_140 | v_225) | v_226) ;
	assign x_347 = ((v_140 | ~v_225) | v_226) ;
	assign x_346 = ((v_140 | v_225) | ~v_226) ;
	assign x_344 = ((~v_137 | ~v_223) | ~v_224) ;
	assign x_343 = ((v_137 | ~v_223) | v_224) ;
	assign x_341 = ((~v_134 | v_221) | v_222) ;
	assign x_340 = ((~v_134 | ~v_221) | ~v_222) ;
	assign x_338 = ((v_134 | v_221) | ~v_222) ;
	assign x_337 = ((~v_130 | v_219) | v_220) ;
	assign x_335 = ((v_130 | ~v_219) | v_220) ;
	assign x_334 = ((v_130 | v_219) | ~v_220) ;
	assign x_332 = ((~v_127 | ~v_217) | ~v_218) ;
	assign x_331 = ((v_127 | ~v_217) | v_218) ;
	assign x_329 = ((~v_124 | v_215) | v_216) ;
	assign x_328 = ((~v_124 | ~v_215) | ~v_216) ;
	assign x_326 = ((v_124 | v_215) | ~v_216) ;
	assign x_325 = ((~v_120 | v_213) | v_214) ;
	assign x_323 = ((v_120 | ~v_213) | v_214) ;
	assign x_322 = ((v_120 | v_213) | ~v_214) ;
	assign x_320 = ((~v_117 | ~v_211) | ~v_212) ;
	assign x_319 = ((v_117 | ~v_211) | v_212) ;
	assign x_317 = ((~v_114 | v_209) | v_210) ;
	assign x_316 = ((~v_114 | ~v_209) | ~v_210) ;
	assign x_314 = ((v_114 | v_209) | ~v_210) ;
	assign x_313 = ((~v_110 | v_207) | v_208) ;
	assign x_311 = ((v_110 | ~v_207) | v_208) ;
	assign x_310 = ((v_110 | v_207) | ~v_208) ;
	assign x_308 = ((~v_107 | ~v_205) | ~v_206) ;
	assign x_307 = ((v_107 | ~v_205) | v_206) ;
	assign x_305 = ((~v_103 | v_203) | v_204) ;
	assign x_304 = ((~v_103 | ~v_203) | ~v_204) ;
	assign x_302 = ((v_103 | v_203) | ~v_204) ;
	assign x_301 = ((~v_100 | v_201) | v_202) ;
	assign x_299 = ((v_100 | ~v_201) | v_202) ;
	assign x_298 = ((v_100 | v_201) | ~v_202) ;
	assign x_296 = ((~v_96 | ~v_199) | ~v_200) ;
	assign x_295 = ((v_96 | ~v_199) | v_200) ;
	assign x_293 = ((~v_93 | v_197) | v_198) ;
	assign x_292 = ((~v_93 | ~v_197) | ~v_198) ;
	assign x_290 = ((v_93 | v_197) | ~v_198) ;
	assign x_289 = ((~v_89 | v_195) | v_196) ;
	assign x_287 = ((v_89 | ~v_195) | v_196) ;
	assign x_286 = ((v_89 | v_195) | ~v_196) ;
	assign x_282 = ((v_86 | v_193) | ~v_194) ;
	assign x_281 = ((~v_82 | v_191) | v_192) ;
	assign x_279 = ((v_82 | ~v_191) | v_192) ;
	assign x_278 = ((v_82 | v_191) | ~v_192) ;
	assign x_276 = ((~v_79 | ~v_189) | ~v_190) ;
	assign x_275 = ((v_79 | ~v_189) | v_190) ;
	assign x_273 = ((~v_75 | v_187) | v_188) ;
	assign x_272 = ((~v_75 | ~v_187) | ~v_188) ;
	assign x_270 = ((v_75 | v_187) | ~v_188) ;
	assign x_269 = ((~v_72 | v_247) | v_248) ;
	assign x_267 = ((v_72 | ~v_247) | v_248) ;
	assign x_266 = ((v_72 | v_247) | ~v_248) ;
	assign x_264 = ((~v_70 | v_185) | v_186) ;
	assign x_263 = (~v_70 | ~v_7) ;
	assign x_261 = (((v_70 | v_185) | ~v_186) | v_7) ;
	assign x_260 = ((~v_69 | ~v_185) | ~v_186) ;
	assign x_258 = ((v_69 | v_186) | v_70) ;
	assign x_257 = ((v_69 | v_185) | v_70) ;
	assign x_255 = ((~v_67 | ~v_185) | ~v_186) ;
	assign x_254 = ((v_67 | ~v_185) | v_186) ;
	assign x_252 = ((~v_64 | ~v_243) | ~v_244) ;
	assign x_251 = (~v_64 | v_245) ;
	assign x_249 = (~v_64 | v_246) ;
	assign x_248 = ((((v_64 | ~v_243) | v_244) | ~v_245) | ~v_246) ;
	assign x_246 = ((~v_63 | ~v_243) | ~v_244) ;
	assign x_245 = (~v_63 | ~v_64) ;
	assign x_243 = ((v_63 | v_243) | v_64) ;
	assign x_242 = ((~v_61 | ~v_241) | ~v_242) ;
	assign x_240 = ((v_61 | v_242) | v_62) ;
	assign x_239 = ((v_61 | v_241) | v_62) ;
	assign x_235 = (((v_60 | ~v_239) | v_240) | v_61) ;
	assign x_234 = (((v_60 | v_239) | ~v_240) | v_61) ;
	assign x_232 = (~v_59 | ~v_60) ;
	assign x_231 = ((v_59 | v_240) | v_60) ;
	assign x_229 = ((~v_57 | ~v_237) | ~v_238) ;
	assign x_228 = (~v_57 | ~v_58) ;
	assign x_226 = ((v_57 | v_237) | v_58) ;
	assign x_225 = ((~v_56 | ~v_235) | ~v_236) ;
	assign x_223 = (~v_56 | ~v_57) ;
	assign x_222 = (((v_56 | ~v_235) | v_236) | v_57) ;
	assign x_220 = ((~v_55 | ~v_235) | ~v_236) ;
	assign x_219 = (~v_55 | ~v_56) ;
	assign x_217 = ((v_55 | v_235) | v_56) ;
	assign x_216 = ((~v_54 | ~v_233) | ~v_234) ;
	assign x_214 = (~v_54 | ~v_55) ;
	assign x_213 = (((v_54 | ~v_233) | v_234) | v_55) ;
	assign x_211 = ((~v_53 | ~v_233) | ~v_234) ;
	assign x_210 = (~v_53 | ~v_54) ;
	assign x_208 = ((v_53 | v_233) | v_54) ;
	assign x_207 = ((~v_52 | ~v_231) | ~v_232) ;
	assign x_205 = (~v_52 | ~v_53) ;
	assign x_204 = (((v_52 | ~v_231) | v_232) | v_53) ;
	assign x_202 = ((~v_51 | ~v_231) | ~v_232) ;
	assign x_201 = (~v_51 | ~v_52) ;
	assign x_199 = ((v_51 | v_231) | v_52) ;
	assign x_198 = ((~v_50 | ~v_229) | ~v_230) ;
	assign x_196 = (~v_50 | ~v_51) ;
	assign x_195 = (((v_50 | ~v_229) | v_230) | v_51) ;
	assign x_193 = ((~v_49 | ~v_229) | ~v_230) ;
	assign x_192 = (~v_49 | ~v_50) ;
	assign x_188 = ((~v_48 | v_227) | v_228) ;
	assign x_187 = (~v_48 | ~v_49) ;
	assign x_185 = (((v_48 | v_227) | ~v_228) | v_49) ;
	assign x_184 = ((~v_47 | ~v_227) | ~v_228) ;
	assign x_182 = ((v_47 | v_228) | v_48) ;
	assign x_181 = ((v_47 | v_227) | v_48) ;
	assign x_179 = ((~v_46 | v_225) | v_226) ;
	assign x_178 = (~v_46 | ~v_47) ;
	assign x_176 = (((v_46 | v_225) | ~v_226) | v_47) ;
	assign x_175 = ((~v_45 | ~v_225) | ~v_226) ;
	assign x_173 = ((v_45 | v_226) | v_46) ;
	assign x_172 = ((v_45 | v_225) | v_46) ;
	assign x_170 = ((~v_44 | v_223) | v_224) ;
	assign x_169 = (~v_44 | ~v_45) ;
	assign x_167 = (((v_44 | v_223) | ~v_224) | v_45) ;
	assign x_166 = ((~v_43 | ~v_223) | ~v_224) ;
	assign x_164 = ((v_43 | v_224) | v_44) ;
	assign x_163 = ((v_43 | v_223) | v_44) ;
	assign x_161 = ((~v_42 | v_221) | v_222) ;
	assign x_160 = (~v_42 | ~v_43) ;
	assign x_158 = (((v_42 | v_221) | ~v_222) | v_43) ;
	assign x_157 = ((~v_41 | ~v_221) | ~v_222) ;
	assign x_155 = ((v_41 | v_222) | v_42) ;
	assign x_154 = ((v_41 | v_221) | v_42) ;
	assign x_152 = ((~v_40 | v_219) | v_220) ;
	assign x_151 = (~v_40 | ~v_41) ;
	assign x_149 = (((v_40 | v_219) | ~v_220) | v_41) ;
	assign x_148 = ((~v_39 | ~v_219) | ~v_220) ;
	assign x_146 = ((v_39 | v_220) | v_40) ;
	assign x_145 = ((v_39 | v_219) | v_40) ;
	assign x_141 = (((v_38 | ~v_217) | v_218) | v_39) ;
	assign x_140 = (((v_38 | v_217) | ~v_218) | v_39) ;
	assign x_138 = (~v_37 | ~v_38) ;
	assign x_137 = ((v_37 | v_218) | v_38) ;
	assign x_135 = ((~v_36 | ~v_215) | ~v_216) ;
	assign x_134 = ((~v_36 | v_215) | v_216) ;
	assign x_132 = (((v_36 | ~v_215) | v_216) | v_37) ;
	assign x_131 = (((v_36 | v_215) | ~v_216) | v_37) ;
	assign x_129 = (~v_35 | ~v_36) ;
	assign x_128 = ((v_35 | v_216) | v_36) ;
	assign x_126 = ((~v_34 | ~v_213) | ~v_214) ;
	assign x_125 = ((~v_34 | v_213) | v_214) ;
	assign x_123 = (((v_34 | ~v_213) | v_214) | v_35) ;
	assign x_122 = (((v_34 | v_213) | ~v_214) | v_35) ;
	assign x_120 = (~v_33 | ~v_34) ;
	assign x_119 = ((v_33 | v_214) | v_34) ;
	assign x_117 = ((~v_32 | ~v_211) | ~v_212) ;
	assign x_116 = ((~v_32 | v_211) | v_212) ;
	assign x_114 = (((v_32 | ~v_211) | v_212) | v_33) ;
	assign x_113 = (((v_32 | v_211) | ~v_212) | v_33) ;
	assign x_111 = (~v_31 | ~v_32) ;
	assign x_110 = ((v_31 | v_212) | v_32) ;
	assign x_108 = ((~v_30 | ~v_209) | ~v_210) ;
	assign x_107 = ((~v_30 | v_209) | v_210) ;
	assign x_105 = (((v_30 | ~v_209) | v_210) | v_31) ;
	assign x_104 = (((v_30 | v_209) | ~v_210) | v_31) ;
	assign x_102 = (~v_29 | ~v_30) ;
	assign x_101 = ((v_29 | v_210) | v_30) ;
	assign x_99 = ((~v_28 | ~v_207) | ~v_208) ;
	assign x_98 = ((~v_28 | v_207) | v_208) ;
	assign x_94 = ((~v_27 | ~v_207) | ~v_208) ;
	assign x_93 = (~v_27 | ~v_28) ;
	assign x_91 = ((v_27 | v_207) | v_28) ;
	assign x_90 = ((~v_26 | ~v_205) | ~v_206) ;
	assign x_88 = (~v_26 | ~v_27) ;
	assign x_87 = (((v_26 | ~v_205) | v_206) | v_27) ;
	assign x_85 = ((~v_25 | ~v_205) | ~v_206) ;
	assign x_84 = (~v_25 | ~v_26) ;
	assign x_82 = ((v_25 | v_205) | v_26) ;
	assign x_81 = ((~v_24 | ~v_203) | ~v_204) ;
	assign x_79 = (~v_24 | ~v_25) ;
	assign x_78 = (((v_24 | ~v_203) | v_204) | v_25) ;
	assign x_76 = ((~v_23 | ~v_203) | ~v_204) ;
	assign x_75 = (~v_23 | ~v_24) ;
	assign x_73 = ((v_23 | v_203) | v_24) ;
	assign x_72 = ((~v_22 | ~v_201) | ~v_202) ;
	assign x_70 = (~v_22 | ~v_23) ;
	assign x_69 = (((v_22 | ~v_201) | v_202) | v_23) ;
	assign x_67 = ((~v_21 | ~v_201) | ~v_202) ;
	assign x_66 = (~v_21 | ~v_22) ;
	assign x_64 = ((v_21 | v_201) | v_22) ;
	assign x_63 = ((~v_20 | ~v_199) | ~v_200) ;
	assign x_61 = (~v_20 | ~v_21) ;
	assign x_60 = (((v_20 | ~v_199) | v_200) | v_21) ;
	assign x_58 = ((~v_19 | ~v_199) | ~v_200) ;
	assign x_57 = (~v_19 | ~v_20) ;
	assign x_55 = ((v_19 | v_199) | v_20) ;
	assign x_54 = ((~v_18 | ~v_197) | ~v_198) ;
	assign x_52 = (~v_18 | ~v_19) ;
	assign x_51 = (((v_18 | ~v_197) | v_198) | v_19) ;
	assign x_47 = ((v_17 | v_198) | v_18) ;
	assign x_46 = ((v_17 | v_197) | v_18) ;
	assign x_44 = ((~v_16 | v_195) | v_196) ;
	assign x_43 = (~v_16 | ~v_17) ;
	assign x_41 = (((v_16 | v_195) | ~v_196) | v_17) ;
	assign x_40 = ((~v_15 | ~v_195) | ~v_196) ;
	assign x_38 = ((v_15 | v_196) | v_16) ;
	assign x_37 = ((v_15 | v_195) | v_16) ;
	assign x_35 = ((~v_14 | v_193) | v_194) ;
	assign x_34 = (~v_14 | ~v_15) ;
	assign x_32 = (((v_14 | v_193) | ~v_194) | v_15) ;
	assign x_31 = ((~v_13 | ~v_193) | ~v_194) ;
	assign x_29 = ((v_13 | v_194) | v_14) ;
	assign x_28 = ((v_13 | v_193) | v_14) ;
	assign x_26 = ((~v_12 | v_191) | v_192) ;
	assign x_25 = (~v_12 | ~v_13) ;
	assign x_23 = (((v_12 | v_191) | ~v_192) | v_13) ;
	assign x_22 = ((~v_11 | ~v_191) | ~v_192) ;
	assign x_20 = ((v_11 | v_192) | v_12) ;
	assign x_19 = ((v_11 | v_191) | v_12) ;
	assign x_17 = ((~v_10 | v_189) | v_190) ;
	assign x_16 = (~v_10 | ~v_11) ;
	assign x_14 = (((v_10 | v_189) | ~v_190) | v_11) ;
	assign x_13 = ((~v_9 | ~v_189) | ~v_190) ;
	assign x_11 = ((v_9 | v_190) | v_10) ;
	assign x_10 = ((v_9 | v_189) | v_10) ;
	assign x_8 = ((~v_8 | v_187) | v_188) ;
	assign x_7 = (~v_8 | ~v_9) ;
	assign x_5 = (((v_8 | v_187) | ~v_188) | v_9) ;
	assign x_4 = ((~v_7 | ~v_187) | ~v_188) ;
	assign x_745 = (x_376 & x_377) ;
	assign x_375 = ((v_169 | ~v_243) | v_244) ;
	assign x_743 = (x_373 & x_374) ;
	assign x_372 = ((~v_163 | ~v_239) | ~v_240) ;
	assign x_740 = (x_370 & x_371) ;
	assign x_369 = ((~v_157 | v_235) | v_236) ;
	assign x_738 = (x_367 & x_368) ;
	assign x_366 = ((v_157 | v_235) | ~v_236) ;
	assign x_734 = (x_364 & x_365) ;
	assign x_363 = ((v_154 | ~v_233) | v_234) ;
	assign x_732 = (x_361 & x_362) ;
	assign x_360 = ((~v_150 | ~v_231) | ~v_232) ;
	assign x_729 = (x_358 & x_359) ;
	assign x_357 = ((~v_147 | v_229) | v_230) ;
	assign x_727 = (x_355 & x_356) ;
	assign x_354 = ((v_147 | v_229) | ~v_230) ;
	assign x_722 = (x_352 & x_353) ;
	assign x_351 = ((v_144 | ~v_227) | v_228) ;
	assign x_720 = (x_349 & x_350) ;
	assign x_348 = ((~v_140 | ~v_225) | ~v_226) ;
	assign x_717 = (x_346 & x_347) ;
	assign x_345 = ((~v_137 | v_223) | v_224) ;
	assign x_715 = (x_343 & x_344) ;
	assign x_342 = ((v_137 | v_223) | ~v_224) ;
	assign x_711 = (x_340 & x_341) ;
	assign x_339 = ((v_134 | ~v_221) | v_222) ;
	assign x_709 = (x_337 & x_338) ;
	assign x_336 = ((~v_130 | ~v_219) | ~v_220) ;
	assign x_706 = (x_334 & x_335) ;
	assign x_333 = ((~v_127 | v_217) | v_218) ;
	assign x_704 = (x_331 & x_332) ;
	assign x_330 = ((v_127 | v_217) | ~v_218) ;
	assign x_698 = (x_328 & x_329) ;
	assign x_327 = ((v_124 | ~v_215) | v_216) ;
	assign x_696 = (x_325 & x_326) ;
	assign x_324 = ((~v_120 | ~v_213) | ~v_214) ;
	assign x_693 = (x_322 & x_323) ;
	assign x_321 = ((~v_117 | v_211) | v_212) ;
	assign x_691 = (x_319 & x_320) ;
	assign x_318 = ((v_117 | v_211) | ~v_212) ;
	assign x_687 = (x_316 & x_317) ;
	assign x_315 = ((v_114 | ~v_209) | v_210) ;
	assign x_685 = (x_313 & x_314) ;
	assign x_312 = ((~v_110 | ~v_207) | ~v_208) ;
	assign x_682 = (x_310 & x_311) ;
	assign x_309 = ((~v_107 | v_205) | v_206) ;
	assign x_680 = (x_307 & x_308) ;
	assign x_306 = ((v_107 | v_205) | ~v_206) ;
	assign x_675 = (x_304 & x_305) ;
	assign x_303 = ((v_103 | ~v_203) | v_204) ;
	assign x_673 = (x_301 & x_302) ;
	assign x_300 = ((~v_100 | ~v_201) | ~v_202) ;
	assign x_670 = (x_298 & x_299) ;
	assign x_297 = ((~v_96 | v_199) | v_200) ;
	assign x_668 = (x_295 & x_296) ;
	assign x_294 = ((v_96 | v_199) | ~v_200) ;
	assign x_664 = (x_292 & x_293) ;
	assign x_291 = ((v_93 | ~v_197) | v_198) ;
	assign x_662 = (x_289 & x_290) ;
	assign x_288 = ((~v_89 | ~v_195) | ~v_196) ;
	assign x_659 = (x_286 & x_287) ;
	assign x_285 = ((~v_86 | v_193) | v_194) ;
	assign x_284 = ((~v_86 | ~v_193) | ~v_194) ;
	assign x_283 = ((v_86 | ~v_193) | v_194) ;
	assign x_651 = (x_281 & x_282) ;
	assign x_280 = ((~v_82 | ~v_191) | ~v_192) ;
	assign x_649 = (x_278 & x_279) ;
	assign x_277 = ((~v_79 | v_189) | v_190) ;
	assign x_646 = (x_275 & x_276) ;
	assign x_274 = ((v_79 | v_189) | ~v_190) ;
	assign x_644 = (x_272 & x_273) ;
	assign x_271 = ((v_75 | ~v_187) | v_188) ;
	assign x_640 = (x_269 & x_270) ;
	assign x_268 = ((~v_72 | ~v_247) | ~v_248) ;
	assign x_638 = (x_266 & x_267) ;
	assign x_265 = ((~v_70 | ~v_185) | ~v_186) ;
	assign x_635 = (x_263 & x_264) ;
	assign x_262 = (((v_70 | ~v_185) | v_186) | v_7) ;
	assign x_633 = (x_260 & x_261) ;
	assign x_259 = (~v_69 | ~v_70) ;
	assign x_628 = (x_257 & x_258) ;
	assign x_256 = ((~v_67 | v_185) | v_186) ;
	assign x_626 = (x_254 & x_255) ;
	assign x_253 = ((v_67 | v_185) | ~v_186) ;
	assign x_623 = (x_251 & x_252) ;
	assign x_250 = ((~v_64 | v_243) | v_244) ;
	assign x_621 = (x_248 & x_249) ;
	assign x_247 = ((((v_64 | v_243) | ~v_244) | ~v_245) | ~v_246) ;
	assign x_617 = (x_245 & x_246) ;
	assign x_244 = ((v_63 | v_244) | v_64) ;
	assign x_615 = (x_242 & x_243) ;
	assign x_241 = (~v_61 | ~v_62) ;
	assign x_612 = (x_239 & x_240) ;
	assign x_238 = ((~v_60 | ~v_239) | ~v_240) ;
	assign x_237 = ((~v_60 | v_239) | v_240) ;
	assign x_236 = (~v_60 | ~v_61) ;
	assign x_605 = (x_234 & x_235) ;
	assign x_233 = ((~v_59 | ~v_239) | ~v_240) ;
	assign x_603 = (x_231 & x_232) ;
	assign x_230 = ((v_59 | v_239) | v_60) ;
	assign x_600 = (x_228 & x_229) ;
	assign x_227 = ((v_57 | v_238) | v_58) ;
	assign x_598 = (x_225 & x_226) ;
	assign x_224 = ((~v_56 | v_235) | v_236) ;
	assign x_594 = (x_222 & x_223) ;
	assign x_221 = (((v_56 | v_235) | ~v_236) | v_57) ;
	assign x_592 = (x_219 & x_220) ;
	assign x_218 = ((v_55 | v_236) | v_56) ;
	assign x_589 = (x_216 & x_217) ;
	assign x_215 = ((~v_54 | v_233) | v_234) ;
	assign x_587 = (x_213 & x_214) ;
	assign x_212 = (((v_54 | v_233) | ~v_234) | v_55) ;
	assign x_582 = (x_210 & x_211) ;
	assign x_209 = ((v_53 | v_234) | v_54) ;
	assign x_580 = (x_207 & x_208) ;
	assign x_206 = ((~v_52 | v_231) | v_232) ;
	assign x_577 = (x_204 & x_205) ;
	assign x_203 = (((v_52 | v_231) | ~v_232) | v_53) ;
	assign x_575 = (x_201 & x_202) ;
	assign x_200 = ((v_51 | v_232) | v_52) ;
	assign x_571 = (x_198 & x_199) ;
	assign x_197 = ((~v_50 | v_229) | v_230) ;
	assign x_569 = (x_195 & x_196) ;
	assign x_194 = (((v_50 | v_229) | ~v_230) | v_51) ;
	assign x_566 = (x_192 & x_193) ;
	assign x_191 = ((v_49 | v_230) | v_50) ;
	assign x_190 = ((v_49 | v_229) | v_50) ;
	assign x_189 = ((~v_48 | ~v_227) | ~v_228) ;
	assign x_557 = (x_187 & x_188) ;
	assign x_186 = (((v_48 | ~v_227) | v_228) | v_49) ;
	assign x_555 = (x_184 & x_185) ;
	assign x_183 = (~v_47 | ~v_48) ;
	assign x_552 = (x_181 & x_182) ;
	assign x_180 = ((~v_46 | ~v_225) | ~v_226) ;
	assign x_550 = (x_178 & x_179) ;
	assign x_177 = (((v_46 | ~v_225) | v_226) | v_47) ;
	assign x_546 = (x_175 & x_176) ;
	assign x_174 = (~v_45 | ~v_46) ;
	assign x_544 = (x_172 & x_173) ;
	assign x_171 = ((~v_44 | ~v_223) | ~v_224) ;
	assign x_541 = (x_169 & x_170) ;
	assign x_168 = (((v_44 | ~v_223) | v_224) | v_45) ;
	assign x_539 = (x_166 & x_167) ;
	assign x_165 = (~v_43 | ~v_44) ;
	assign x_534 = (x_163 & x_164) ;
	assign x_162 = ((~v_42 | ~v_221) | ~v_222) ;
	assign x_532 = (x_160 & x_161) ;
	assign x_159 = (((v_42 | ~v_221) | v_222) | v_43) ;
	assign x_529 = (x_157 & x_158) ;
	assign x_156 = (~v_41 | ~v_42) ;
	assign x_527 = (x_154 & x_155) ;
	assign x_153 = ((~v_40 | ~v_219) | ~v_220) ;
	assign x_523 = (x_151 & x_152) ;
	assign x_150 = (((v_40 | ~v_219) | v_220) | v_41) ;
	assign x_521 = (x_148 & x_149) ;
	assign x_147 = (~v_39 | ~v_40) ;
	assign x_518 = (x_145 & x_146) ;
	assign x_144 = ((~v_38 | ~v_217) | ~v_218) ;
	assign x_143 = ((~v_38 | v_217) | v_218) ;
	assign x_142 = (~v_38 | ~v_39) ;
	assign x_511 = (x_140 & x_141) ;
	assign x_139 = ((~v_37 | ~v_217) | ~v_218) ;
	assign x_509 = (x_137 & x_138) ;
	assign x_136 = ((v_37 | v_217) | v_38) ;
	assign x_506 = (x_134 & x_135) ;
	assign x_133 = (~v_36 | ~v_37) ;
	assign x_504 = (x_131 & x_132) ;
	assign x_130 = ((~v_35 | ~v_215) | ~v_216) ;
	assign x_500 = (x_128 & x_129) ;
	assign x_127 = ((v_35 | v_215) | v_36) ;
	assign x_498 = (x_125 & x_126) ;
	assign x_124 = (~v_34 | ~v_35) ;
	assign x_495 = (x_122 & x_123) ;
	assign x_121 = ((~v_33 | ~v_213) | ~v_214) ;
	assign x_493 = (x_119 & x_120) ;
	assign x_118 = ((v_33 | v_213) | v_34) ;
	assign x_488 = (x_116 & x_117) ;
	assign x_115 = (~v_32 | ~v_33) ;
	assign x_486 = (x_113 & x_114) ;
	assign x_112 = ((~v_31 | ~v_211) | ~v_212) ;
	assign x_483 = (x_110 & x_111) ;
	assign x_109 = ((v_31 | v_211) | v_32) ;
	assign x_481 = (x_107 & x_108) ;
	assign x_106 = (~v_30 | ~v_31) ;
	assign x_477 = (x_104 & x_105) ;
	assign x_103 = ((~v_29 | ~v_209) | ~v_210) ;
	assign x_475 = (x_101 & x_102) ;
	assign x_100 = ((v_29 | v_209) | v_30) ;
	assign x_472 = (x_98 & x_99) ;
	assign x_97 = (~v_28 | ~v_29) ;
	assign x_96 = (((v_28 | ~v_207) | v_208) | v_29) ;
	assign x_95 = (((v_28 | v_207) | ~v_208) | v_29) ;
	assign x_464 = (x_93 & x_94) ;
	assign x_92 = ((v_27 | v_208) | v_28) ;
	assign x_462 = (x_90 & x_91) ;
	assign x_89 = ((~v_26 | v_205) | v_206) ;
	assign x_459 = (x_87 & x_88) ;
	assign x_86 = (((v_26 | v_205) | ~v_206) | v_27) ;
	assign x_457 = (x_84 & x_85) ;
	assign x_83 = ((v_25 | v_206) | v_26) ;
	assign x_453 = (x_81 & x_82) ;
	assign x_80 = ((~v_24 | v_203) | v_204) ;
	assign x_451 = (x_78 & x_79) ;
	assign x_77 = (((v_24 | v_203) | ~v_204) | v_25) ;
	assign x_448 = (x_75 & x_76) ;
	assign x_74 = ((v_23 | v_204) | v_24) ;
	assign x_446 = (x_72 & x_73) ;
	assign x_71 = ((~v_22 | v_201) | v_202) ;
	assign x_441 = (x_69 & x_70) ;
	assign x_68 = (((v_22 | v_201) | ~v_202) | v_23) ;
	assign x_439 = (x_66 & x_67) ;
	assign x_65 = ((v_21 | v_202) | v_22) ;
	assign x_436 = (x_63 & x_64) ;
	assign x_62 = ((~v_20 | v_199) | v_200) ;
	assign x_434 = (x_60 & x_61) ;
	assign x_59 = (((v_20 | v_199) | ~v_200) | v_21) ;
	assign x_430 = (x_57 & x_58) ;
	assign x_56 = ((v_19 | v_200) | v_20) ;
	assign x_428 = (x_54 & x_55) ;
	assign x_53 = ((~v_18 | v_197) | v_198) ;
	assign x_425 = (x_51 & x_52) ;
	assign x_50 = (((v_18 | v_197) | ~v_198) | v_19) ;
	assign x_49 = ((~v_17 | ~v_197) | ~v_198) ;
	assign x_48 = (~v_17 | ~v_18) ;
	assign x_418 = (x_46 & x_47) ;
	assign x_45 = ((~v_16 | ~v_195) | ~v_196) ;
	assign x_416 = (x_43 & x_44) ;
	assign x_42 = (((v_16 | ~v_195) | v_196) | v_17) ;
	assign x_413 = (x_40 & x_41) ;
	assign x_39 = (~v_15 | ~v_16) ;
	assign x_411 = (x_37 & x_38) ;
	assign x_36 = ((~v_14 | ~v_193) | ~v_194) ;
	assign x_407 = (x_34 & x_35) ;
	assign x_33 = (((v_14 | ~v_193) | v_194) | v_15) ;
	assign x_405 = (x_31 & x_32) ;
	assign x_30 = (~v_13 | ~v_14) ;
	assign x_402 = (x_28 & x_29) ;
	assign x_27 = ((~v_12 | ~v_191) | ~v_192) ;
	assign x_400 = (x_25 & x_26) ;
	assign x_24 = (((v_12 | ~v_191) | v_192) | v_13) ;
	assign x_395 = (x_22 & x_23) ;
	assign x_21 = (~v_11 | ~v_12) ;
	assign x_393 = (x_19 & x_20) ;
	assign x_18 = ((~v_10 | ~v_189) | ~v_190) ;
	assign x_390 = (x_16 & x_17) ;
	assign x_15 = (((v_10 | ~v_189) | v_190) | v_11) ;
	assign x_388 = (x_13 & x_14) ;
	assign x_12 = (~v_9 | ~v_10) ;
	assign x_384 = (x_10 & x_11) ;
	assign x_9 = ((~v_8 | ~v_187) | ~v_188) ;
	assign x_382 = (x_7 & x_8) ;
	assign x_6 = (((v_8 | ~v_187) | v_188) | v_9) ;
	assign x_379 = (x_4 & x_5) ;
	assign x_3 = (~v_7 | ~v_8) ;
	assign x_2 = ((v_7 | v_188) | v_8) ;
	assign x_1 = ((v_7 | v_187) | v_8) ;
	assign x_746 = (x_375 & x_745) ;
	assign x_744 = (x_372 & x_743) ;
	assign x_741 = (x_369 & x_740) ;
	assign x_739 = (x_366 & x_738) ;
	assign x_735 = (x_363 & x_734) ;
	assign x_733 = (x_360 & x_732) ;
	assign x_730 = (x_357 & x_729) ;
	assign x_728 = (x_354 & x_727) ;
	assign x_723 = (x_351 & x_722) ;
	assign x_721 = (x_348 & x_720) ;
	assign x_718 = (x_345 & x_717) ;
	assign x_716 = (x_342 & x_715) ;
	assign x_712 = (x_339 & x_711) ;
	assign x_710 = (x_336 & x_709) ;
	assign x_707 = (x_333 & x_706) ;
	assign x_705 = (x_330 & x_704) ;
	assign x_699 = (x_327 & x_698) ;
	assign x_697 = (x_324 & x_696) ;
	assign x_694 = (x_321 & x_693) ;
	assign x_692 = (x_318 & x_691) ;
	assign x_688 = (x_315 & x_687) ;
	assign x_686 = (x_312 & x_685) ;
	assign x_683 = (x_309 & x_682) ;
	assign x_681 = (x_306 & x_680) ;
	assign x_676 = (x_303 & x_675) ;
	assign x_674 = (x_300 & x_673) ;
	assign x_671 = (x_297 & x_670) ;
	assign x_669 = (x_294 & x_668) ;
	assign x_665 = (x_291 & x_664) ;
	assign x_663 = (x_288 & x_662) ;
	assign x_660 = (x_285 & x_659) ;
	assign x_658 = (x_283 & x_284) ;
	assign x_652 = (x_280 & x_651) ;
	assign x_650 = (x_277 & x_649) ;
	assign x_647 = (x_274 & x_646) ;
	assign x_645 = (x_271 & x_644) ;
	assign x_641 = (x_268 & x_640) ;
	assign x_639 = (x_265 & x_638) ;
	assign x_636 = (x_262 & x_635) ;
	assign x_634 = (x_259 & x_633) ;
	assign x_629 = (x_256 & x_628) ;
	assign x_627 = (x_253 & x_626) ;
	assign x_624 = (x_250 & x_623) ;
	assign x_622 = (x_247 & x_621) ;
	assign x_618 = (x_244 & x_617) ;
	assign x_616 = (x_241 & x_615) ;
	assign x_613 = (x_238 & x_612) ;
	assign x_611 = (x_236 & x_237) ;
	assign x_606 = (x_233 & x_605) ;
	assign x_604 = (x_230 & x_603) ;
	assign x_601 = (x_227 & x_600) ;
	assign x_599 = (x_224 & x_598) ;
	assign x_595 = (x_221 & x_594) ;
	assign x_593 = (x_218 & x_592) ;
	assign x_590 = (x_215 & x_589) ;
	assign x_588 = (x_212 & x_587) ;
	assign x_583 = (x_209 & x_582) ;
	assign x_581 = (x_206 & x_580) ;
	assign x_578 = (x_203 & x_577) ;
	assign x_576 = (x_200 & x_575) ;
	assign x_572 = (x_197 & x_571) ;
	assign x_570 = (x_194 & x_569) ;
	assign x_567 = (x_191 & x_566) ;
	assign x_565 = (x_189 & x_190) ;
	assign x_558 = (x_186 & x_557) ;
	assign x_556 = (x_183 & x_555) ;
	assign x_553 = (x_180 & x_552) ;
	assign x_551 = (x_177 & x_550) ;
	assign x_547 = (x_174 & x_546) ;
	assign x_545 = (x_171 & x_544) ;
	assign x_542 = (x_168 & x_541) ;
	assign x_540 = (x_165 & x_539) ;
	assign x_535 = (x_162 & x_534) ;
	assign x_533 = (x_159 & x_532) ;
	assign x_530 = (x_156 & x_529) ;
	assign x_528 = (x_153 & x_527) ;
	assign x_524 = (x_150 & x_523) ;
	assign x_522 = (x_147 & x_521) ;
	assign x_519 = (x_144 & x_518) ;
	assign x_517 = (x_142 & x_143) ;
	assign x_512 = (x_139 & x_511) ;
	assign x_510 = (x_136 & x_509) ;
	assign x_507 = (x_133 & x_506) ;
	assign x_505 = (x_130 & x_504) ;
	assign x_501 = (x_127 & x_500) ;
	assign x_499 = (x_124 & x_498) ;
	assign x_496 = (x_121 & x_495) ;
	assign x_494 = (x_118 & x_493) ;
	assign x_489 = (x_115 & x_488) ;
	assign x_487 = (x_112 & x_486) ;
	assign x_484 = (x_109 & x_483) ;
	assign x_482 = (x_106 & x_481) ;
	assign x_478 = (x_103 & x_477) ;
	assign x_476 = (x_100 & x_475) ;
	assign x_473 = (x_97 & x_472) ;
	assign x_471 = (x_95 & x_96) ;
	assign x_465 = (x_92 & x_464) ;
	assign x_463 = (x_89 & x_462) ;
	assign x_460 = (x_86 & x_459) ;
	assign x_458 = (x_83 & x_457) ;
	assign x_454 = (x_80 & x_453) ;
	assign x_452 = (x_77 & x_451) ;
	assign x_449 = (x_74 & x_448) ;
	assign x_447 = (x_71 & x_446) ;
	assign x_442 = (x_68 & x_441) ;
	assign x_440 = (x_65 & x_439) ;
	assign x_437 = (x_62 & x_436) ;
	assign x_435 = (x_59 & x_434) ;
	assign x_431 = (x_56 & x_430) ;
	assign x_429 = (x_53 & x_428) ;
	assign x_426 = (x_50 & x_425) ;
	assign x_424 = (x_48 & x_49) ;
	assign x_419 = (x_45 & x_418) ;
	assign x_417 = (x_42 & x_416) ;
	assign x_414 = (x_39 & x_413) ;
	assign x_412 = (x_36 & x_411) ;
	assign x_408 = (x_33 & x_407) ;
	assign x_406 = (x_30 & x_405) ;
	assign x_403 = (x_27 & x_402) ;
	assign x_401 = (x_24 & x_400) ;
	assign x_396 = (x_21 & x_395) ;
	assign x_394 = (x_18 & x_393) ;
	assign x_391 = (x_15 & x_390) ;
	assign x_389 = (x_12 & x_388) ;
	assign x_385 = (x_9 & x_384) ;
	assign x_383 = (x_6 & x_382) ;
	assign x_380 = (x_3 & x_379) ;
	assign x_378 = (x_1 & x_2) ;
	assign x_747 = (x_744 & x_746) ;
	assign x_742 = (x_739 & x_741) ;
	assign x_736 = (x_733 & x_735) ;
	assign x_731 = (x_728 & x_730) ;
	assign x_724 = (x_721 & x_723) ;
	assign x_719 = (x_716 & x_718) ;
	assign x_713 = (x_710 & x_712) ;
	assign x_708 = (x_705 & x_707) ;
	assign x_700 = (x_697 & x_699) ;
	assign x_695 = (x_692 & x_694) ;
	assign x_689 = (x_686 & x_688) ;
	assign x_684 = (x_681 & x_683) ;
	assign x_677 = (x_674 & x_676) ;
	assign x_672 = (x_669 & x_671) ;
	assign x_666 = (x_663 & x_665) ;
	assign x_661 = (x_658 & x_660) ;
	assign x_653 = (x_650 & x_652) ;
	assign x_648 = (x_645 & x_647) ;
	assign x_642 = (x_639 & x_641) ;
	assign x_637 = (x_634 & x_636) ;
	assign x_630 = (x_627 & x_629) ;
	assign x_625 = (x_622 & x_624) ;
	assign x_619 = (x_616 & x_618) ;
	assign x_614 = (x_611 & x_613) ;
	assign x_607 = (x_604 & x_606) ;
	assign x_602 = (x_599 & x_601) ;
	assign x_596 = (x_593 & x_595) ;
	assign x_591 = (x_588 & x_590) ;
	assign x_584 = (x_581 & x_583) ;
	assign x_579 = (x_576 & x_578) ;
	assign x_573 = (x_570 & x_572) ;
	assign x_568 = (x_565 & x_567) ;
	assign x_559 = (x_556 & x_558) ;
	assign x_554 = (x_551 & x_553) ;
	assign x_548 = (x_545 & x_547) ;
	assign x_543 = (x_540 & x_542) ;
	assign x_536 = (x_533 & x_535) ;
	assign x_531 = (x_528 & x_530) ;
	assign x_525 = (x_522 & x_524) ;
	assign x_520 = (x_517 & x_519) ;
	assign x_513 = (x_510 & x_512) ;
	assign x_508 = (x_505 & x_507) ;
	assign x_502 = (x_499 & x_501) ;
	assign x_497 = (x_494 & x_496) ;
	assign x_490 = (x_487 & x_489) ;
	assign x_485 = (x_482 & x_484) ;
	assign x_479 = (x_476 & x_478) ;
	assign x_474 = (x_471 & x_473) ;
	assign x_466 = (x_463 & x_465) ;
	assign x_461 = (x_458 & x_460) ;
	assign x_455 = (x_452 & x_454) ;
	assign x_450 = (x_447 & x_449) ;
	assign x_443 = (x_440 & x_442) ;
	assign x_438 = (x_435 & x_437) ;
	assign x_432 = (x_429 & x_431) ;
	assign x_427 = (x_424 & x_426) ;
	assign x_420 = (x_417 & x_419) ;
	assign x_415 = (x_412 & x_414) ;
	assign x_409 = (x_406 & x_408) ;
	assign x_404 = (x_401 & x_403) ;
	assign x_397 = (x_394 & x_396) ;
	assign x_392 = (x_389 & x_391) ;
	assign x_386 = (x_383 & x_385) ;
	assign x_381 = (x_378 & x_380) ;
	assign x_748 = (x_742 & x_747) ;
	assign x_737 = (x_731 & x_736) ;
	assign x_725 = (x_719 & x_724) ;
	assign x_714 = (x_708 & x_713) ;
	assign x_701 = (x_695 & x_700) ;
	assign x_690 = (x_684 & x_689) ;
	assign x_678 = (x_672 & x_677) ;
	assign x_667 = (x_661 & x_666) ;
	assign x_654 = (x_648 & x_653) ;
	assign x_643 = (x_637 & x_642) ;
	assign x_631 = (x_625 & x_630) ;
	assign x_620 = (x_614 & x_619) ;
	assign x_608 = (x_602 & x_607) ;
	assign x_597 = (x_591 & x_596) ;
	assign x_585 = (x_579 & x_584) ;
	assign x_574 = (x_568 & x_573) ;
	assign x_560 = (x_554 & x_559) ;
	assign x_549 = (x_543 & x_548) ;
	assign x_537 = (x_531 & x_536) ;
	assign x_526 = (x_520 & x_525) ;
	assign x_514 = (x_508 & x_513) ;
	assign x_503 = (x_497 & x_502) ;
	assign x_491 = (x_485 & x_490) ;
	assign x_480 = (x_474 & x_479) ;
	assign x_467 = (x_461 & x_466) ;
	assign x_456 = (x_450 & x_455) ;
	assign x_444 = (x_438 & x_443) ;
	assign x_433 = (x_427 & x_432) ;
	assign x_421 = (x_415 & x_420) ;
	assign x_410 = (x_404 & x_409) ;
	assign x_398 = (x_392 & x_397) ;
	assign x_387 = (x_381 & x_386) ;
	assign x_749 = (x_737 & x_748) ;
	assign x_726 = (x_714 & x_725) ;
	assign x_702 = (x_690 & x_701) ;
	assign x_679 = (x_667 & x_678) ;
	assign x_655 = (x_643 & x_654) ;
	assign x_632 = (x_620 & x_631) ;
	assign x_609 = (x_597 & x_608) ;
	assign x_586 = (x_574 & x_585) ;
	assign x_561 = (x_549 & x_560) ;
	assign x_538 = (x_526 & x_537) ;
	assign x_515 = (x_503 & x_514) ;
	assign x_492 = (x_480 & x_491) ;
	assign x_468 = (x_456 & x_467) ;
	assign x_445 = (x_433 & x_444) ;
	assign x_422 = (x_410 & x_421) ;
	assign x_399 = (x_387 & x_398) ;
	assign x_750 = (x_726 & x_749) ;
	assign x_703 = (x_679 & x_702) ;
	assign x_656 = (x_632 & x_655) ;
	assign x_610 = (x_586 & x_609) ;
	assign x_562 = (x_538 & x_561) ;
	assign x_516 = (x_492 & x_515) ;
	assign x_469 = (x_445 & x_468) ;
	assign x_423 = (x_399 & x_422) ;
	assign x_751 = (x_703 & x_750) ;
	assign x_657 = (x_610 & x_656) ;
	assign x_563 = (x_516 & x_562) ;
	assign x_470 = (x_423 & x_469) ;
	assign x_752 = (x_657 & x_751) ;
	assign x_564 = (x_470 & x_563) ;
	assign x_753 = (x_564 & x_752) ;
	assign v_279 = 1 ;
	assign v_183 = 1 ;
	assign v_182 = 1 ;
	assign v_181 = 1 ;
	assign v_180 = 1 ;
	assign v_179 = 1 ;
	assign v_178 = 1 ;
	assign v_177 = 1 ;
	assign v_176 = 1 ;
	assign v_175 = 1 ;
	assign v_174 = 1 ;
	assign v_173 = 1 ;
	assign v_172 = 1 ;
	assign v_171 = 1 ;
	assign v_170 = 1 ;
	assign v_166 = 0 ;
	assign v_164 = 0 ;
	assign v_161 = 0 ;
	assign v_160 = 1 ;
	assign v_158 = 0 ;
	assign v_155 = 0 ;
	assign v_152 = 0 ;
	assign v_151 = 1 ;
	assign v_148 = 0 ;
	assign v_145 = 0 ;
	assign v_142 = 0 ;
	assign v_141 = 1 ;
	assign v_138 = 0 ;
	assign v_135 = 0 ;
	assign v_132 = 0 ;
	assign v_131 = 1 ;
	assign v_128 = 0 ;
	assign v_125 = 0 ;
	assign v_122 = 0 ;
	assign v_121 = 1 ;
	assign v_118 = 0 ;
	assign v_115 = 0 ;
	assign v_112 = 0 ;
	assign v_111 = 1 ;
	assign v_108 = 0 ;
	assign v_105 = 0 ;
	assign v_104 = 1 ;
	assign v_101 = 0 ;
	assign v_98 = 0 ;
	assign v_97 = 1 ;
	assign v_94 = 0 ;
	assign v_91 = 0 ;
	assign v_90 = 1 ;
	assign v_87 = 0 ;
	assign v_84 = 0 ;
	assign v_83 = 1 ;
	assign v_80 = 0 ;
	assign v_77 = 0 ;
	assign v_76 = 1 ;
	assign v_73 = 0 ;
	assign v_68 = 0 ;
	assign v_5 = 0 ;
	assign v_4 = 1 ;
	assign v_3 = 1 ;
	assign v_2 = 1 ;
	assign v_1 = 0 ;
	assign o_1 = x_753 ;
endmodule
