// skolem function for order file variables
// Generated using findDep.cpp 
module formula (v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_15, v_20, v_22, v_24, v_25, v_26, v_29, v_31, v_33, v_34, v_36, v_38, v_40, v_41, v_43, v_45, v_47, v_49, v_51, v_53, v_55, v_58, v_59, v_66, v_68, v_72, v_76, v_78, v_80, v_84, v_91, v_96, v_101, v_107, v_108, v_112, v_115, v_116, v_125, v_131, v_132, v_136, v_139, v_140, v_329, v_330, v_331, v_332, v_333, v_334, v_335, v_336, v_337, v_338, v_342, v_347, v_349, v_351, v_352, v_353, v_356, v_358, v_360, v_361, v_363, v_365, v_367, v_368, v_370, v_372, v_374, v_376, v_378, v_380, v_382, v_385, v_386, v_393, v_395, v_399, v_403, v_405, v_407, v_411, v_418, v_423, v_428, v_434, v_435, v_439, v_442, v_443, v_452, v_458, v_459, v_463, v_466, v_467, o_1);
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_15;
input v_20;
input v_22;
input v_24;
input v_25;
input v_26;
input v_29;
input v_31;
input v_33;
input v_34;
input v_36;
input v_38;
input v_40;
input v_41;
input v_43;
input v_45;
input v_47;
input v_49;
input v_51;
input v_53;
input v_55;
input v_58;
input v_59;
input v_66;
input v_68;
input v_72;
input v_76;
input v_78;
input v_80;
input v_84;
input v_91;
input v_96;
input v_101;
input v_107;
input v_108;
input v_112;
input v_115;
input v_116;
input v_125;
input v_131;
input v_132;
input v_136;
input v_139;
input v_140;
input v_329;
input v_330;
input v_331;
input v_332;
input v_333;
input v_334;
input v_335;
input v_336;
input v_337;
input v_338;
input v_342;
input v_347;
input v_349;
input v_351;
input v_352;
input v_353;
input v_356;
input v_358;
input v_360;
input v_361;
input v_363;
input v_365;
input v_367;
input v_368;
input v_370;
input v_372;
input v_374;
input v_376;
input v_378;
input v_380;
input v_382;
input v_385;
input v_386;
input v_393;
input v_395;
input v_399;
input v_403;
input v_405;
input v_407;
input v_411;
input v_418;
input v_423;
input v_428;
input v_434;
input v_435;
input v_439;
input v_442;
input v_443;
input v_452;
input v_458;
input v_459;
input v_463;
input v_466;
input v_467;
output o_1;
wire v_1;
wire v_12;
wire v_13;
wire v_14;
wire v_16;
wire v_17;
wire v_18;
wire v_19;
wire v_21;
wire v_23;
wire v_27;
wire v_28;
wire v_30;
wire v_32;
wire v_35;
wire v_37;
wire v_39;
wire v_42;
wire v_44;
wire v_46;
wire v_48;
wire v_50;
wire v_52;
wire v_54;
wire v_56;
wire v_57;
wire v_60;
wire v_61;
wire v_62;
wire v_63;
wire v_64;
wire v_65;
wire v_67;
wire v_69;
wire v_70;
wire v_71;
wire v_73;
wire v_74;
wire v_75;
wire v_77;
wire v_79;
wire v_81;
wire v_82;
wire v_83;
wire v_85;
wire v_86;
wire v_87;
wire v_88;
wire v_89;
wire v_90;
wire v_92;
wire v_93;
wire v_94;
wire v_95;
wire v_97;
wire v_98;
wire v_99;
wire v_100;
wire v_102;
wire v_103;
wire v_104;
wire v_105;
wire v_106;
wire v_109;
wire v_110;
wire v_111;
wire v_113;
wire v_114;
wire v_117;
wire v_118;
wire v_119;
wire v_120;
wire v_121;
wire v_122;
wire v_123;
wire v_124;
wire v_126;
wire v_127;
wire v_128;
wire v_129;
wire v_130;
wire v_133;
wire v_134;
wire v_135;
wire v_137;
wire v_138;
wire v_141;
wire v_142;
wire v_143;
wire v_144;
wire v_145;
wire v_146;
wire v_147;
wire v_148;
wire v_149;
wire v_150;
wire v_151;
wire v_152;
wire v_153;
wire v_154;
wire v_155;
wire v_156;
wire v_157;
wire v_158;
wire v_159;
wire v_160;
wire v_161;
wire v_162;
wire v_163;
wire v_164;
wire v_165;
wire v_166;
wire v_167;
wire v_168;
wire v_169;
wire v_170;
wire v_171;
wire v_172;
wire v_173;
wire v_174;
wire v_175;
wire v_176;
wire v_177;
wire v_178;
wire v_179;
wire v_180;
wire v_181;
wire v_182;
wire v_183;
wire v_184;
wire v_185;
wire v_186;
wire v_187;
wire v_188;
wire v_189;
wire v_190;
wire v_191;
wire v_192;
wire v_193;
wire v_194;
wire v_195;
wire v_196;
wire v_197;
wire v_198;
wire v_199;
wire v_200;
wire v_201;
wire v_202;
wire v_203;
wire v_204;
wire v_205;
wire v_206;
wire v_207;
wire v_208;
wire v_209;
wire v_210;
wire v_211;
wire v_212;
wire v_213;
wire v_214;
wire v_215;
wire v_216;
wire v_217;
wire v_218;
wire v_219;
wire v_220;
wire v_221;
wire v_222;
wire v_223;
wire v_224;
wire v_225;
wire v_226;
wire v_227;
wire v_228;
wire v_229;
wire v_230;
wire v_231;
wire v_232;
wire v_233;
wire v_234;
wire v_235;
wire v_236;
wire v_237;
wire v_238;
wire v_239;
wire v_240;
wire v_241;
wire v_242;
wire v_243;
wire v_244;
wire v_245;
wire v_246;
wire v_247;
wire v_248;
wire v_249;
wire v_250;
wire v_251;
wire v_252;
wire v_253;
wire v_254;
wire v_255;
wire v_256;
wire v_257;
wire v_258;
wire v_259;
wire v_260;
wire v_261;
wire v_262;
wire v_263;
wire v_264;
wire v_265;
wire v_266;
wire v_267;
wire v_268;
wire v_269;
wire v_270;
wire v_271;
wire v_272;
wire v_273;
wire v_274;
wire v_275;
wire v_276;
wire v_277;
wire v_278;
wire v_279;
wire v_280;
wire v_281;
wire v_282;
wire v_283;
wire v_284;
wire v_285;
wire v_286;
wire v_287;
wire v_288;
wire v_289;
wire v_290;
wire v_291;
wire v_292;
wire v_293;
wire v_294;
wire v_295;
wire v_296;
wire v_297;
wire v_298;
wire v_299;
wire v_300;
wire v_301;
wire v_302;
wire v_303;
wire v_304;
wire v_305;
wire v_306;
wire v_307;
wire v_308;
wire v_309;
wire v_310;
wire v_311;
wire v_312;
wire v_313;
wire v_314;
wire v_315;
wire v_316;
wire v_317;
wire v_318;
wire v_319;
wire v_320;
wire v_321;
wire v_322;
wire v_323;
wire v_324;
wire v_325;
wire v_326;
wire v_327;
wire v_328;
wire v_339;
wire v_340;
wire v_341;
wire v_343;
wire v_344;
wire v_345;
wire v_346;
wire v_348;
wire v_350;
wire v_354;
wire v_355;
wire v_357;
wire v_359;
wire v_362;
wire v_364;
wire v_366;
wire v_369;
wire v_371;
wire v_373;
wire v_375;
wire v_377;
wire v_379;
wire v_381;
wire v_383;
wire v_384;
wire v_387;
wire v_388;
wire v_389;
wire v_390;
wire v_391;
wire v_392;
wire v_394;
wire v_396;
wire v_397;
wire v_398;
wire v_400;
wire v_401;
wire v_402;
wire v_404;
wire v_406;
wire v_408;
wire v_409;
wire v_410;
wire v_412;
wire v_413;
wire v_414;
wire v_415;
wire v_416;
wire v_417;
wire v_419;
wire v_420;
wire v_421;
wire v_422;
wire v_424;
wire v_425;
wire v_426;
wire v_427;
wire v_429;
wire v_430;
wire v_431;
wire v_432;
wire v_433;
wire v_436;
wire v_437;
wire v_438;
wire v_440;
wire v_441;
wire v_444;
wire v_445;
wire v_446;
wire v_447;
wire v_448;
wire v_449;
wire v_450;
wire v_451;
wire v_453;
wire v_454;
wire v_455;
wire v_456;
wire v_457;
wire v_460;
wire v_461;
wire v_462;
wire v_464;
wire v_465;
wire v_468;
wire v_469;
wire v_470;
wire v_471;
wire v_472;
wire v_473;
wire v_474;
wire v_475;
wire v_476;
wire v_477;
wire v_478;
wire v_479;
wire v_480;
wire v_481;
wire v_482;
wire v_483;
wire v_484;
wire v_485;
wire v_486;
wire v_487;
wire v_488;
wire v_489;
wire v_490;
wire v_491;
wire v_492;
wire v_493;
wire v_494;
wire v_495;
wire v_496;
wire v_497;
wire v_498;
wire v_499;
wire v_500;
wire v_501;
wire v_502;
wire v_503;
wire v_504;
wire v_505;
wire v_506;
wire v_507;
wire v_508;
wire v_509;
wire v_510;
wire v_511;
wire v_512;
wire v_513;
wire v_514;
wire v_515;
wire v_516;
wire v_517;
wire v_518;
wire v_519;
wire v_520;
wire v_521;
wire v_522;
wire v_523;
wire v_524;
wire v_525;
wire v_526;
wire v_527;
wire v_528;
wire v_529;
wire v_530;
wire v_531;
wire v_532;
wire v_533;
wire v_534;
wire v_535;
wire v_536;
wire v_537;
wire v_538;
wire v_539;
wire v_540;
wire v_541;
wire v_542;
wire v_543;
wire v_544;
wire v_545;
wire v_546;
wire v_547;
wire v_548;
wire v_549;
wire v_550;
wire v_551;
wire v_552;
wire v_553;
wire v_554;
wire v_555;
wire v_556;
wire v_557;
wire v_558;
wire v_559;
wire v_560;
wire v_561;
wire v_562;
wire v_563;
wire v_564;
wire v_565;
wire v_566;
wire v_567;
wire v_568;
wire v_569;
wire v_570;
wire v_571;
wire v_572;
wire v_573;
wire v_574;
wire v_575;
wire v_576;
wire v_577;
wire v_578;
wire v_579;
wire v_580;
wire v_581;
wire v_582;
wire v_583;
wire v_584;
wire v_585;
wire v_586;
wire v_587;
wire v_588;
wire v_589;
wire v_590;
wire v_591;
wire v_592;
wire v_593;
wire v_594;
wire v_595;
wire v_596;
wire v_597;
wire v_598;
wire v_599;
wire v_600;
wire v_601;
wire v_602;
wire v_603;
wire v_604;
wire v_605;
wire v_606;
wire v_607;
wire v_608;
wire v_609;
wire v_610;
wire v_611;
wire v_612;
wire v_613;
wire v_614;
wire v_615;
wire v_616;
wire v_617;
wire v_618;
wire v_619;
wire v_620;
wire v_621;
wire v_622;
wire v_623;
wire v_624;
wire v_625;
wire v_626;
wire v_627;
wire v_628;
wire v_629;
wire v_630;
wire v_631;
wire v_632;
wire v_633;
wire v_634;
wire v_635;
wire v_636;
wire v_637;
wire v_638;
wire v_639;
wire v_640;
wire v_641;
wire v_642;
wire v_643;
wire v_644;
wire v_645;
wire v_646;
wire v_647;
wire v_648;
wire v_649;
wire v_650;
wire v_651;
wire v_652;
wire v_653;
wire v_654;
wire v_655;
wire v_656;
wire v_657;
wire v_658;
wire v_659;
wire v_660;
wire v_661;
wire v_662;
wire v_663;
wire v_664;
wire v_665;
wire v_666;
wire v_667;
wire v_668;
wire v_669;
wire v_670;
wire v_671;
wire v_672;
wire v_673;
wire v_674;
wire v_675;
wire v_676;
wire v_677;
wire v_678;
wire v_679;
wire v_680;
wire v_681;
wire v_682;
wire v_683;
wire v_684;
wire v_685;
wire v_686;
wire v_687;
wire v_688;
wire v_689;
wire v_690;
wire v_691;
wire v_692;
wire v_693;
wire v_694;
wire v_695;
wire v_696;
wire v_697;
wire v_698;
wire v_699;
wire v_700;
wire x_1;
assign v_1 = 1;
assign v_16 = 1;
assign v_21 = 1;
assign v_23 = 1;
assign v_30 = 1;
assign v_35 = 1;
assign v_54 = 1;
assign v_77 = 1;
assign v_81 = 1;
assign v_92 = 1;
assign v_97 = 1;
assign v_102 = 1;
assign v_113 = 1;
assign v_117 = 1;
assign v_126 = 1;
assign v_137 = 1;
assign v_141 = 1;
assign v_149 = 1;
assign v_240 = 1;
assign v_343 = 1;
assign v_348 = 1;
assign v_350 = 1;
assign v_357 = 1;
assign v_362 = 1;
assign v_381 = 1;
assign v_404 = 1;
assign v_408 = 1;
assign v_419 = 1;
assign v_424 = 1;
assign v_429 = 1;
assign v_440 = 1;
assign v_444 = 1;
assign v_453 = 1;
assign v_464 = 1;
assign v_468 = 1;
assign v_476 = 1;
assign v_567 = 1;
assign v_12 = v_10 & v_11;
assign v_13 = v_10 & ~v_11;
assign v_17 = v_9 & v_14;
assign v_18 = ~v_9 & v_14;
assign v_27 = v_25 & ~v_26;
assign v_32 = v_31;
assign v_37 = ~v_36;
assign v_39 = v_36 & v_38;
assign v_42 = v_36 & ~v_38 & v_40 & v_41;
assign v_44 = v_36 & ~v_38 & v_40 & ~v_41 & ~v_43;
assign v_46 = v_36 & ~v_38 & ~v_40 & ~v_45;
assign v_48 = v_36 & ~v_38 & ~v_40 & v_45 & v_47;
assign v_50 = v_659 & v_660;
assign v_52 = v_661 & v_662;
assign v_56 = v_663 & v_664;
assign v_57 = v_665 & v_666;
assign v_60 = v_58 & v_59;
assign v_61 = v_58 & ~v_59;
assign v_63 = v_667 & v_668;
assign v_65 = ~v_31 & ~v_33 & v_64;
assign v_67 = ~v_31 & v_33 & ~v_66;
assign v_69 = ~v_31 & v_33 & v_66 & ~v_68;
assign v_70 = ~v_31 & v_33 & v_66 & v_68;
assign v_73 = v_71 & v_72;
assign v_74 = v_71 & ~v_72;
assign v_79 = v_24 & v_28 & v_75 & v_78;
assign v_82 = v_24 & v_28 & v_75 & ~v_78;
assign v_85 = v_83 & v_84;
assign v_86 = v_83 & ~v_84;
assign v_88 = v_8 & v_19 & v_87;
assign v_89 = ~v_8 & v_19;
assign v_93 = v_7 & v_90;
assign v_94 = ~v_7 & v_90;
assign v_98 = v_6 & v_95;
assign v_99 = ~v_6 & v_95;
assign v_103 = v_5 & v_100;
assign v_104 = ~v_5 & v_100;
assign v_106 = v_4 & v_105;
assign v_109 = v_108 & v_100;
assign v_110 = ~v_108 & v_100;
assign v_114 = v_107 & v_111;
assign v_118 = v_115 & v_111;
assign v_119 = ~v_115 & v_111;
assign v_121 = ~v_107 & v_120;
assign v_123 = ~v_4 & v_122;
assign v_127 = v_3 & v_124;
assign v_128 = ~v_3 & v_124;
assign v_130 = v_2 & v_129;
assign v_133 = v_132 & v_124;
assign v_134 = ~v_132 & v_124;
assign v_138 = v_131 & v_135;
assign v_142 = v_139 & v_135;
assign v_143 = ~v_139 & v_135;
assign v_145 = ~v_131 & v_144;
assign v_147 = ~v_2 & v_146;
assign v_150 = v_9;
assign v_152 = v_151 & ~v_24;
assign v_153 = v_151 & v_31;
assign v_154 = v_151 & ~v_31 & v_33 & v_66 & ~v_68;
assign v_155 = v_151 & ~v_31 & v_33 & v_66 & v_68;
assign v_156 = v_151 & ~v_31 & v_33 & ~v_66;
assign v_157 = v_151 & v_34;
assign v_158 = v_151 & ~v_34;
assign v_161 = v_159 & v_160;
assign v_162 = v_669 & v_670;
assign v_164 = v_159 & v_163;
assign v_166 = v_165 & ~v_31 & ~v_33 & v_64;
assign v_168 = v_167 & v_71 & v_72;
assign v_169 = v_167 & v_71 & ~v_72;
assign v_171 = v_170 & v_24 & v_28 & v_75 & v_78;
assign v_172 = v_170 & v_24 & v_28 & v_75 & ~v_78;
assign v_175 = v_173 & v_174;
assign v_177 = v_8 & v_176;
assign v_178 = ~v_8 & v_151;
assign v_180 = v_179 & ~v_91;
assign v_181 = v_179 & v_91;
assign v_183 = v_7 & v_182;
assign v_184 = ~v_7 & v_179;
assign v_186 = v_185 & ~v_96;
assign v_187 = v_185 & v_96;
assign v_189 = v_6 & v_188;
assign v_190 = ~v_6 & v_185;
assign v_192 = v_191 & ~v_101;
assign v_193 = v_191 & v_101;
assign v_195 = v_5 & v_194;
assign v_196 = ~v_5 & v_191;
assign v_198 = v_4 & v_197;
assign v_199 = v_108 & v_194;
assign v_200 = ~v_108 & v_191;
assign v_202 = v_201 & ~v_112;
assign v_203 = v_201 & v_112;
assign v_205 = v_107 & v_204;
assign v_206 = v_201 & ~v_116;
assign v_207 = v_201 & v_116;
assign v_209 = v_115 & v_208;
assign v_210 = ~v_115 & v_201;
assign v_212 = ~v_107 & v_211;
assign v_214 = ~v_4 & v_213;
assign v_216 = v_215 & ~v_125;
assign v_217 = v_215 & v_125;
assign v_219 = v_3 & v_218;
assign v_220 = ~v_3 & v_215;
assign v_222 = v_2 & v_221;
assign v_223 = v_132 & v_218;
assign v_224 = ~v_132 & v_215;
assign v_226 = v_225 & ~v_136;
assign v_227 = v_225 & v_136;
assign v_229 = v_131 & v_228;
assign v_230 = v_225 & ~v_140;
assign v_231 = v_225 & v_140;
assign v_233 = v_139 & v_232;
assign v_234 = ~v_139 & v_225;
assign v_236 = ~v_131 & v_235;
assign v_238 = ~v_2 & v_237;
assign v_241 = v_9;
assign v_243 = v_242 & ~v_24;
assign v_244 = v_242 & v_31;
assign v_245 = v_242 & ~v_31 & v_33 & v_66 & ~v_68;
assign v_246 = v_242 & ~v_31 & v_33 & v_66 & v_68;
assign v_247 = v_242 & ~v_31 & v_33 & ~v_66;
assign v_248 = v_242 & v_34;
assign v_249 = v_242 & ~v_34;
assign v_252 = v_250 & v_251;
assign v_253 = v_671 & v_672;
assign v_254 = v_250 & v_163;
assign v_256 = v_255 & ~v_31 & ~v_33 & v_64;
assign v_258 = v_257 & v_71 & v_72;
assign v_259 = v_257 & v_71 & ~v_72;
assign v_261 = v_260 & v_24 & v_28 & v_75 & v_78;
assign v_262 = v_260 & v_24 & v_28 & v_75 & ~v_78;
assign v_264 = v_263 & v_174;
assign v_266 = v_8 & v_265;
assign v_267 = ~v_8 & v_242;
assign v_269 = v_268 & ~v_91;
assign v_270 = v_268 & v_91;
assign v_272 = v_7 & v_271;
assign v_273 = ~v_7 & v_268;
assign v_275 = v_274 & ~v_96;
assign v_276 = v_274 & v_96;
assign v_278 = v_6 & v_277;
assign v_279 = ~v_6 & v_274;
assign v_281 = v_280 & ~v_101;
assign v_282 = v_280 & v_101;
assign v_284 = v_5 & v_283;
assign v_285 = ~v_5 & v_280;
assign v_287 = v_4 & v_286;
assign v_288 = v_108 & v_283;
assign v_289 = ~v_108 & v_280;
assign v_291 = v_290 & ~v_112;
assign v_292 = v_290 & v_112;
assign v_294 = v_107 & v_293;
assign v_295 = v_290 & ~v_116;
assign v_296 = v_290 & v_116;
assign v_298 = v_115 & v_297;
assign v_299 = ~v_115 & v_290;
assign v_301 = ~v_107 & v_300;
assign v_303 = ~v_4 & v_302;
assign v_305 = v_304 & ~v_125;
assign v_306 = v_304 & v_125;
assign v_308 = v_3 & v_307;
assign v_309 = ~v_3 & v_304;
assign v_311 = v_2 & v_310;
assign v_312 = v_132 & v_307;
assign v_313 = ~v_132 & v_304;
assign v_315 = v_314 & ~v_136;
assign v_316 = v_314 & v_136;
assign v_318 = v_131 & v_317;
assign v_319 = v_314 & ~v_140;
assign v_320 = v_314 & v_140;
assign v_322 = v_139 & v_321;
assign v_323 = ~v_139 & v_314;
assign v_325 = ~v_131 & v_324;
assign v_327 = ~v_2 & v_326;
assign v_339 = v_337 & v_338;
assign v_340 = v_337 & ~v_338;
assign v_344 = v_336 & v_341;
assign v_345 = ~v_336 & v_341;
assign v_354 = v_352 & ~v_353;
assign v_359 = v_358;
assign v_364 = ~v_363;
assign v_366 = v_363 & v_365;
assign v_369 = v_363 & ~v_365 & v_367 & v_368;
assign v_371 = v_363 & ~v_365 & v_367 & ~v_368 & ~v_370;
assign v_373 = v_363 & ~v_365 & ~v_367 & ~v_372;
assign v_375 = v_363 & ~v_365 & ~v_367 & v_372 & v_374;
assign v_377 = v_673 & v_674;
assign v_379 = v_675 & v_676;
assign v_383 = v_677 & v_678;
assign v_384 = v_679 & v_680;
assign v_387 = v_385 & v_386;
assign v_388 = v_385 & ~v_386;
assign v_390 = v_681 & v_682;
assign v_392 = ~v_358 & ~v_360 & v_391;
assign v_394 = ~v_358 & v_360 & ~v_393;
assign v_396 = ~v_358 & v_360 & v_393 & ~v_395;
assign v_397 = ~v_358 & v_360 & v_393 & v_395;
assign v_400 = v_398 & v_399;
assign v_401 = v_398 & ~v_399;
assign v_406 = v_351 & v_355 & v_402 & v_405;
assign v_409 = v_351 & v_355 & v_402 & ~v_405;
assign v_412 = v_410 & v_411;
assign v_413 = v_410 & ~v_411;
assign v_415 = v_335 & v_346 & v_414;
assign v_416 = ~v_335 & v_346;
assign v_420 = v_334 & v_417;
assign v_421 = ~v_334 & v_417;
assign v_425 = v_333 & v_422;
assign v_426 = ~v_333 & v_422;
assign v_430 = v_332 & v_427;
assign v_431 = ~v_332 & v_427;
assign v_433 = v_331 & v_432;
assign v_436 = v_435 & v_427;
assign v_437 = ~v_435 & v_427;
assign v_441 = v_434 & v_438;
assign v_445 = v_442 & v_438;
assign v_446 = ~v_442 & v_438;
assign v_448 = ~v_434 & v_447;
assign v_450 = ~v_331 & v_449;
assign v_454 = v_330 & v_451;
assign v_455 = ~v_330 & v_451;
assign v_457 = v_329 & v_456;
assign v_460 = v_459 & v_451;
assign v_461 = ~v_459 & v_451;
assign v_465 = v_458 & v_462;
assign v_469 = v_466 & v_462;
assign v_470 = ~v_466 & v_462;
assign v_472 = ~v_458 & v_471;
assign v_474 = ~v_329 & v_473;
assign v_477 = v_336;
assign v_479 = v_478 & ~v_351;
assign v_480 = v_478 & v_358;
assign v_481 = v_478 & ~v_358 & v_360 & v_393 & ~v_395;
assign v_482 = v_478 & ~v_358 & v_360 & v_393 & v_395;
assign v_483 = v_478 & ~v_358 & v_360 & ~v_393;
assign v_484 = v_478 & v_361;
assign v_485 = v_478 & ~v_361;
assign v_488 = v_486 & v_487;
assign v_489 = v_683 & v_684;
assign v_491 = v_486 & v_490;
assign v_493 = v_492 & ~v_358 & ~v_360 & v_391;
assign v_495 = v_494 & v_398 & v_399;
assign v_496 = v_494 & v_398 & ~v_399;
assign v_498 = v_497 & v_351 & v_355 & v_402 & v_405;
assign v_499 = v_497 & v_351 & v_355 & v_402 & ~v_405;
assign v_502 = v_500 & v_501;
assign v_504 = v_335 & v_503;
assign v_505 = ~v_335 & v_478;
assign v_507 = v_506 & ~v_418;
assign v_508 = v_506 & v_418;
assign v_510 = v_334 & v_509;
assign v_511 = ~v_334 & v_506;
assign v_513 = v_512 & ~v_423;
assign v_514 = v_512 & v_423;
assign v_516 = v_333 & v_515;
assign v_517 = ~v_333 & v_512;
assign v_519 = v_518 & ~v_428;
assign v_520 = v_518 & v_428;
assign v_522 = v_332 & v_521;
assign v_523 = ~v_332 & v_518;
assign v_525 = v_331 & v_524;
assign v_526 = v_435 & v_521;
assign v_527 = ~v_435 & v_518;
assign v_529 = v_528 & ~v_439;
assign v_530 = v_528 & v_439;
assign v_532 = v_434 & v_531;
assign v_533 = v_528 & ~v_443;
assign v_534 = v_528 & v_443;
assign v_536 = v_442 & v_535;
assign v_537 = ~v_442 & v_528;
assign v_539 = ~v_434 & v_538;
assign v_541 = ~v_331 & v_540;
assign v_543 = v_542 & ~v_452;
assign v_544 = v_542 & v_452;
assign v_546 = v_330 & v_545;
assign v_547 = ~v_330 & v_542;
assign v_549 = v_329 & v_548;
assign v_550 = v_459 & v_545;
assign v_551 = ~v_459 & v_542;
assign v_553 = v_552 & ~v_463;
assign v_554 = v_552 & v_463;
assign v_556 = v_458 & v_555;
assign v_557 = v_552 & ~v_467;
assign v_558 = v_552 & v_467;
assign v_560 = v_466 & v_559;
assign v_561 = ~v_466 & v_552;
assign v_563 = ~v_458 & v_562;
assign v_565 = ~v_329 & v_564;
assign v_568 = v_336;
assign v_570 = v_569 & ~v_351;
assign v_571 = v_569 & v_358;
assign v_572 = v_569 & ~v_358 & v_360 & v_393 & ~v_395;
assign v_573 = v_569 & ~v_358 & v_360 & v_393 & v_395;
assign v_574 = v_569 & ~v_358 & v_360 & ~v_393;
assign v_575 = v_569 & v_361;
assign v_576 = v_569 & ~v_361;
assign v_579 = v_577 & v_578;
assign v_580 = v_685 & v_686;
assign v_581 = v_577 & v_490;
assign v_583 = v_582 & ~v_358 & ~v_360 & v_391;
assign v_585 = v_584 & v_398 & v_399;
assign v_586 = v_584 & v_398 & ~v_399;
assign v_588 = v_587 & v_351 & v_355 & v_402 & v_405;
assign v_589 = v_587 & v_351 & v_355 & v_402 & ~v_405;
assign v_591 = v_590 & v_501;
assign v_593 = v_335 & v_592;
assign v_594 = ~v_335 & v_569;
assign v_596 = v_595 & ~v_418;
assign v_597 = v_595 & v_418;
assign v_599 = v_334 & v_598;
assign v_600 = ~v_334 & v_595;
assign v_602 = v_601 & ~v_423;
assign v_603 = v_601 & v_423;
assign v_605 = v_333 & v_604;
assign v_606 = ~v_333 & v_601;
assign v_608 = v_607 & ~v_428;
assign v_609 = v_607 & v_428;
assign v_611 = v_332 & v_610;
assign v_612 = ~v_332 & v_607;
assign v_614 = v_331 & v_613;
assign v_615 = v_435 & v_610;
assign v_616 = ~v_435 & v_607;
assign v_618 = v_617 & ~v_439;
assign v_619 = v_617 & v_439;
assign v_621 = v_434 & v_620;
assign v_622 = v_617 & ~v_443;
assign v_623 = v_617 & v_443;
assign v_625 = v_442 & v_624;
assign v_626 = ~v_442 & v_617;
assign v_628 = ~v_434 & v_627;
assign v_630 = ~v_331 & v_629;
assign v_632 = v_631 & ~v_452;
assign v_633 = v_631 & v_452;
assign v_635 = v_330 & v_634;
assign v_636 = ~v_330 & v_631;
assign v_638 = v_329 & v_637;
assign v_639 = v_459 & v_634;
assign v_640 = ~v_459 & v_631;
assign v_642 = v_641 & ~v_463;
assign v_643 = v_641 & v_463;
assign v_645 = v_458 & v_644;
assign v_646 = v_641 & ~v_467;
assign v_647 = v_641 & v_467;
assign v_649 = v_466 & v_648;
assign v_650 = ~v_466 & v_641;
assign v_652 = ~v_458 & v_651;
assign v_654 = ~v_329 & v_653;
assign v_658 = ~v_656 & ~v_657 & v_475;
assign v_659 = v_36 & ~v_38 & v_40 & ~v_41 & v_43;
assign v_660 = v_49;
assign v_661 = v_36 & ~v_38 & v_40 & ~v_41 & v_43;
assign v_662 = ~v_49 & v_51;
assign v_663 = v_36 & ~v_38 & ~v_40 & v_45 & ~v_47;
assign v_664 = v_55;
assign v_665 = v_36 & ~v_38 & ~v_40 & v_45 & ~v_47;
assign v_666 = ~v_55;
assign v_667 = v_36 & ~v_38 & v_40 & ~v_41 & v_43;
assign v_668 = ~v_49 & ~v_51 & v_62;
assign v_669 = v_159 & v_36 & ~v_38 & v_40 & ~v_41;
assign v_670 = v_43 & ~v_49 & ~v_51 & v_62;
assign v_671 = v_250 & v_36 & ~v_38 & v_40 & ~v_41;
assign v_672 = v_43 & ~v_49 & ~v_51 & v_62;
assign v_673 = v_363 & ~v_365 & v_367 & ~v_368 & v_370;
assign v_674 = v_376;
assign v_675 = v_363 & ~v_365 & v_367 & ~v_368 & v_370;
assign v_676 = ~v_376 & v_378;
assign v_677 = v_363 & ~v_365 & ~v_367 & v_372 & ~v_374;
assign v_678 = v_382;
assign v_679 = v_363 & ~v_365 & ~v_367 & v_372 & ~v_374;
assign v_680 = ~v_382;
assign v_681 = v_363 & ~v_365 & v_367 & ~v_368 & v_370;
assign v_682 = ~v_376 & ~v_378 & v_389;
assign v_683 = v_486 & v_363 & ~v_365 & v_367 & ~v_368;
assign v_684 = v_370 & ~v_376 & ~v_378 & v_389;
assign v_685 = v_577 & v_363 & ~v_365 & v_367 & ~v_368;
assign v_686 = v_370 & ~v_376 & ~v_378 & v_389;
assign v_14 = ~v_10 | v_12 | v_13;
assign v_19 = v_17 | v_18;
assign v_28 = ~v_25 | v_27;
assign v_62 = ~v_58 | v_60 | v_61;
assign v_64 = v_687 | v_688 | v_689;
assign v_71 = v_65 | v_67 | v_69 | v_70;
assign v_75 = v_32 | v_73 | v_74;
assign v_83 = v_79 | v_82;
assign v_87 = ~v_24 | v_85 | v_86;
assign v_90 = v_88 | v_89;
assign v_95 = v_93 | v_94;
assign v_100 = v_98 | v_99;
assign v_105 = v_103 | v_104;
assign v_111 = v_109 | v_110;
assign v_120 = v_118 | v_119;
assign v_122 = v_114 | v_121;
assign v_124 = v_106 | v_123;
assign v_129 = v_127 | v_128;
assign v_135 = v_133 | v_134;
assign v_144 = v_142 | v_143;
assign v_146 = v_138 | v_145;
assign v_148 = v_130 | v_147;
assign v_151 = v_150 | ~v_9;
assign v_159 = v_157 | v_158;
assign v_160 = v_690 | v_691;
assign v_163 = v_56 | v_57;
assign v_165 = v_161 | v_162 | v_164;
assign v_167 = v_154 | v_155 | v_156 | v_166;
assign v_170 = v_153 | v_168 | v_169;
assign v_173 = v_171 | v_172;
assign v_174 = v_85 | v_86;
assign v_176 = v_152 | v_175;
assign v_179 = v_177 | v_178;
assign v_182 = v_180 | v_181;
assign v_185 = v_183 | v_184;
assign v_188 = v_186 | v_187;
assign v_191 = v_189 | v_190;
assign v_194 = v_192 | v_193;
assign v_197 = v_195 | v_196;
assign v_201 = v_199 | v_200;
assign v_204 = v_202 | v_203;
assign v_208 = v_206 | v_207;
assign v_211 = v_209 | v_210;
assign v_213 = v_205 | v_212;
assign v_215 = v_198 | v_214;
assign v_218 = v_216 | v_217;
assign v_221 = v_219 | v_220;
assign v_225 = v_223 | v_224;
assign v_228 = v_226 | v_227;
assign v_232 = v_230 | v_231;
assign v_235 = v_233 | v_234;
assign v_237 = v_229 | v_236;
assign v_239 = v_222 | v_238;
assign v_242 = v_241 | ~v_9;
assign v_250 = v_248 | v_249;
assign v_251 = v_692 | v_693;
assign v_255 = v_252 | v_253 | v_254;
assign v_257 = v_245 | v_246 | v_247 | v_256;
assign v_260 = v_244 | v_258 | v_259;
assign v_263 = v_261 | v_262;
assign v_265 = v_243 | v_264;
assign v_268 = v_266 | v_267;
assign v_271 = v_269 | v_270;
assign v_274 = v_272 | v_273;
assign v_277 = v_275 | v_276;
assign v_280 = v_278 | v_279;
assign v_283 = v_281 | v_282;
assign v_286 = v_284 | v_285;
assign v_290 = v_288 | v_289;
assign v_293 = v_291 | v_292;
assign v_297 = v_295 | v_296;
assign v_300 = v_298 | v_299;
assign v_302 = v_294 | v_301;
assign v_304 = v_287 | v_303;
assign v_307 = v_305 | v_306;
assign v_310 = v_308 | v_309;
assign v_314 = v_312 | v_313;
assign v_317 = v_315 | v_316;
assign v_321 = v_319 | v_320;
assign v_324 = v_322 | v_323;
assign v_326 = v_318 | v_325;
assign v_328 = v_311 | v_327;
assign v_341 = ~v_337 | v_339 | v_340;
assign v_346 = v_344 | v_345;
assign v_355 = ~v_352 | v_354;
assign v_389 = ~v_385 | v_387 | v_388;
assign v_391 = v_694 | v_695 | v_696;
assign v_398 = v_392 | v_394 | v_396 | v_397;
assign v_402 = v_359 | v_400 | v_401;
assign v_410 = v_406 | v_409;
assign v_414 = ~v_351 | v_412 | v_413;
assign v_417 = v_415 | v_416;
assign v_422 = v_420 | v_421;
assign v_427 = v_425 | v_426;
assign v_432 = v_430 | v_431;
assign v_438 = v_436 | v_437;
assign v_447 = v_445 | v_446;
assign v_449 = v_441 | v_448;
assign v_451 = v_433 | v_450;
assign v_456 = v_454 | v_455;
assign v_462 = v_460 | v_461;
assign v_471 = v_469 | v_470;
assign v_473 = v_465 | v_472;
assign v_475 = v_457 | v_474;
assign v_478 = v_477 | ~v_336;
assign v_486 = v_484 | v_485;
assign v_487 = v_697 | v_698;
assign v_490 = v_383 | v_384;
assign v_492 = v_488 | v_489 | v_491;
assign v_494 = v_481 | v_482 | v_483 | v_493;
assign v_497 = v_480 | v_495 | v_496;
assign v_500 = v_498 | v_499;
assign v_501 = v_412 | v_413;
assign v_503 = v_479 | v_502;
assign v_506 = v_504 | v_505;
assign v_509 = v_507 | v_508;
assign v_512 = v_510 | v_511;
assign v_515 = v_513 | v_514;
assign v_518 = v_516 | v_517;
assign v_521 = v_519 | v_520;
assign v_524 = v_522 | v_523;
assign v_528 = v_526 | v_527;
assign v_531 = v_529 | v_530;
assign v_535 = v_533 | v_534;
assign v_538 = v_536 | v_537;
assign v_540 = v_532 | v_539;
assign v_542 = v_525 | v_541;
assign v_545 = v_543 | v_544;
assign v_548 = v_546 | v_547;
assign v_552 = v_550 | v_551;
assign v_555 = v_553 | v_554;
assign v_559 = v_557 | v_558;
assign v_562 = v_560 | v_561;
assign v_564 = v_556 | v_563;
assign v_566 = v_549 | v_565;
assign v_569 = v_568 | ~v_336;
assign v_577 = v_575 | v_576;
assign v_578 = v_699 | v_700;
assign v_582 = v_579 | v_580 | v_581;
assign v_584 = v_572 | v_573 | v_574 | v_583;
assign v_587 = v_571 | v_585 | v_586;
assign v_590 = v_588 | v_589;
assign v_592 = v_570 | v_591;
assign v_595 = v_593 | v_594;
assign v_598 = v_596 | v_597;
assign v_601 = v_599 | v_600;
assign v_604 = v_602 | v_603;
assign v_607 = v_605 | v_606;
assign v_610 = v_608 | v_609;
assign v_613 = v_611 | v_612;
assign v_617 = v_615 | v_616;
assign v_620 = v_618 | v_619;
assign v_624 = v_622 | v_623;
assign v_627 = v_625 | v_626;
assign v_629 = v_621 | v_628;
assign v_631 = v_614 | v_630;
assign v_634 = v_632 | v_633;
assign v_637 = v_635 | v_636;
assign v_641 = v_639 | v_640;
assign v_644 = v_642 | v_643;
assign v_648 = v_646 | v_647;
assign v_651 = v_649 | v_650;
assign v_653 = v_645 | v_652;
assign v_655 = v_638 | v_654;
assign v_687 = v_37 | v_39 | v_42 | v_44 | v_46;
assign v_688 = v_48 | v_50 | v_52 | v_56 | v_57;
assign v_689 = v_63;
assign v_690 = v_37 | v_39 | v_42 | v_44 | v_46;
assign v_691 = v_48 | v_50 | v_52;
assign v_692 = v_37 | v_39 | v_42 | v_44 | v_46;
assign v_693 = v_48 | v_50 | v_52;
assign v_694 = v_364 | v_366 | v_369 | v_371 | v_373;
assign v_695 = v_375 | v_377 | v_379 | v_383 | v_384;
assign v_696 = v_390;
assign v_697 = v_364 | v_366 | v_369 | v_371 | v_373;
assign v_698 = v_375 | v_377 | v_379;
assign v_699 = v_364 | v_366 | v_369 | v_371 | v_373;
assign v_700 = v_375 | v_377 | v_379;
assign v_656 = ~v_566 ^ ~v_239;
assign v_657 = ~v_655 ^ ~v_328;
assign x_1 = ~v_148 | v_658;
assign o_1 = x_1;
endmodule
