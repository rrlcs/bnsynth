// skolem function for order file variables
// Generated using findDep.cpp 
module formula (v_131, v_144, v_1128, v_1138, v_1148, v_224, v_237, v_250, v_711, v_1018, v_1028, v_1038, v_816, v_185, v_198, v_211, v_4, v_3, v_98, v_111, v_124, v_141, v_8, v_13, v_182, v_195, v_208, v_221, v_234, v_247, v_6, v_9, v_2, v_362, v_381, v_394, v_407, v_420, v_433, v_446, v_467, v_482, v_503, v_576, v_560, v_558, v_511, v_505, v_518, v_1, v_17, v_42, v_39, v_721, v_715, v_734, v_728, v_741, v_530, v_10, v_11, v_15, v_21, v_525, v_527, v_539, v_765, v_759, v_772, v_452, v_470, v_485, v_23, v_66, v_65, v_68, v_88, v_101, v_114, v_998, v_1008, v_556, v_77, v_277, v_371, v_384, v_397, v_410, v_423, v_436, v_566, v_265, v_71, v_70, v_73, v_75, v_271, v_62, v_63, v_97, v_110, v_123, v_140, v_153, v_170, v_181, v_194, v_207, v_220, v_233, v_246, v_259, v_335, v_350, v_361, v_380, v_393, v_406, v_419, v_432, v_445, v_466, v_481, v_496, v_499, v_502, v_634, v_649, v_658, v_667, v_676, v_949, v_972, v_985, v_996, v_1006, v_1016, v_1026, v_1036, v_1046, v_1049, v_1056, v_1069, v_1082, v_1095, v_1108, v_1117, v_1126, v_1136, v_1146, v_1156, v_1165, v_1174, v_1183, o_1);
input v_131;
input v_144;
input v_1128;
input v_1138;
input v_1148;
input v_224;
input v_237;
input v_250;
input v_711;
input v_1018;
input v_1028;
input v_1038;
input v_816;
input v_185;
input v_198;
input v_211;
input v_4;
input v_3;
input v_98;
input v_111;
input v_124;
input v_141;
input v_8;
input v_13;
input v_182;
input v_195;
input v_208;
input v_221;
input v_234;
input v_247;
input v_6;
input v_9;
input v_2;
input v_362;
input v_381;
input v_394;
input v_407;
input v_420;
input v_433;
input v_446;
input v_467;
input v_482;
input v_503;
input v_576;
input v_560;
input v_558;
input v_511;
input v_505;
input v_518;
input v_1;
input v_17;
input v_42;
input v_39;
input v_721;
input v_715;
input v_734;
input v_728;
input v_741;
input v_530;
input v_10;
input v_11;
input v_15;
input v_21;
input v_525;
input v_527;
input v_539;
input v_765;
input v_759;
input v_772;
input v_452;
input v_470;
input v_485;
input v_23;
input v_66;
input v_65;
input v_68;
input v_88;
input v_101;
input v_114;
input v_998;
input v_1008;
input v_556;
input v_77;
input v_277;
input v_371;
input v_384;
input v_397;
input v_410;
input v_423;
input v_436;
input v_566;
input v_265;
input v_71;
input v_70;
input v_73;
input v_75;
input v_271;
input v_62;
input v_63;
input v_97;
input v_110;
input v_123;
input v_140;
input v_153;
input v_170;
input v_181;
input v_194;
input v_207;
input v_220;
input v_233;
input v_246;
input v_259;
input v_335;
input v_350;
input v_361;
input v_380;
input v_393;
input v_406;
input v_419;
input v_432;
input v_445;
input v_466;
input v_481;
input v_496;
input v_499;
input v_502;
input v_634;
input v_649;
input v_658;
input v_667;
input v_676;
input v_949;
input v_972;
input v_985;
input v_996;
input v_1006;
input v_1016;
input v_1026;
input v_1036;
input v_1046;
input v_1049;
input v_1056;
input v_1069;
input v_1082;
input v_1095;
input v_1108;
input v_1117;
input v_1126;
input v_1136;
input v_1146;
input v_1156;
input v_1165;
input v_1174;
input v_1183;
output o_1;
wire v_5;
wire v_7;
wire v_12;
wire v_14;
wire v_16;
wire v_18;
wire v_19;
wire v_20;
wire v_22;
wire v_24;
wire v_25;
wire v_26;
wire v_27;
wire v_28;
wire v_29;
wire v_30;
wire v_31;
wire v_32;
wire v_33;
wire v_34;
wire v_35;
wire v_36;
wire v_37;
wire v_38;
wire v_40;
wire v_41;
wire v_43;
wire v_44;
wire v_45;
wire v_46;
wire v_47;
wire v_48;
wire v_49;
wire v_50;
wire v_51;
wire v_52;
wire v_53;
wire v_54;
wire v_55;
wire v_56;
wire v_57;
wire v_58;
wire v_59;
wire v_60;
wire v_61;
wire v_64;
wire v_67;
wire v_69;
wire v_72;
wire v_74;
wire v_76;
wire v_78;
wire v_79;
wire v_80;
wire v_81;
wire v_82;
wire v_83;
wire v_84;
wire v_85;
wire v_86;
wire v_87;
wire v_89;
wire v_90;
wire v_91;
wire v_92;
wire v_93;
wire v_94;
wire v_95;
wire v_96;
wire v_99;
wire v_100;
wire v_102;
wire v_103;
wire v_104;
wire v_105;
wire v_106;
wire v_107;
wire v_108;
wire v_109;
wire v_112;
wire v_113;
wire v_115;
wire v_116;
wire v_117;
wire v_118;
wire v_119;
wire v_120;
wire v_121;
wire v_122;
wire v_125;
wire v_126;
wire v_127;
wire v_128;
wire v_129;
wire v_130;
wire v_132;
wire v_133;
wire v_134;
wire v_135;
wire v_136;
wire v_137;
wire v_138;
wire v_139;
wire v_142;
wire v_143;
wire v_145;
wire v_146;
wire v_147;
wire v_148;
wire v_149;
wire v_150;
wire v_151;
wire v_152;
wire v_154;
wire v_155;
wire v_156;
wire v_157;
wire v_158;
wire v_159;
wire v_160;
wire v_161;
wire v_162;
wire v_163;
wire v_164;
wire v_165;
wire v_166;
wire v_167;
wire v_168;
wire v_169;
wire v_171;
wire v_172;
wire v_173;
wire v_174;
wire v_175;
wire v_176;
wire v_177;
wire v_178;
wire v_179;
wire v_180;
wire v_183;
wire v_184;
wire v_186;
wire v_187;
wire v_188;
wire v_189;
wire v_190;
wire v_191;
wire v_192;
wire v_193;
wire v_196;
wire v_197;
wire v_199;
wire v_200;
wire v_201;
wire v_202;
wire v_203;
wire v_204;
wire v_205;
wire v_206;
wire v_209;
wire v_210;
wire v_212;
wire v_213;
wire v_214;
wire v_215;
wire v_216;
wire v_217;
wire v_218;
wire v_219;
wire v_222;
wire v_223;
wire v_225;
wire v_226;
wire v_227;
wire v_228;
wire v_229;
wire v_230;
wire v_231;
wire v_232;
wire v_235;
wire v_236;
wire v_238;
wire v_239;
wire v_240;
wire v_241;
wire v_242;
wire v_243;
wire v_244;
wire v_245;
wire v_248;
wire v_249;
wire v_251;
wire v_252;
wire v_253;
wire v_254;
wire v_255;
wire v_256;
wire v_257;
wire v_258;
wire v_260;
wire v_261;
wire v_262;
wire v_263;
wire v_264;
wire v_266;
wire v_267;
wire v_268;
wire v_269;
wire v_270;
wire v_272;
wire v_273;
wire v_274;
wire v_275;
wire v_276;
wire v_278;
wire v_279;
wire v_280;
wire v_281;
wire v_282;
wire v_283;
wire v_284;
wire v_285;
wire v_286;
wire v_287;
wire v_288;
wire v_289;
wire v_290;
wire v_291;
wire v_292;
wire v_293;
wire v_294;
wire v_295;
wire v_296;
wire v_297;
wire v_298;
wire v_299;
wire v_300;
wire v_301;
wire v_302;
wire v_303;
wire v_304;
wire v_305;
wire v_306;
wire v_307;
wire v_308;
wire v_309;
wire v_310;
wire v_311;
wire v_312;
wire v_313;
wire v_314;
wire v_315;
wire v_316;
wire v_317;
wire v_318;
wire v_319;
wire v_320;
wire v_321;
wire v_322;
wire v_323;
wire v_324;
wire v_325;
wire v_326;
wire v_327;
wire v_328;
wire v_329;
wire v_330;
wire v_331;
wire v_332;
wire v_333;
wire v_334;
wire v_336;
wire v_337;
wire v_338;
wire v_339;
wire v_340;
wire v_341;
wire v_342;
wire v_343;
wire v_344;
wire v_345;
wire v_346;
wire v_347;
wire v_348;
wire v_349;
wire v_351;
wire v_352;
wire v_353;
wire v_354;
wire v_355;
wire v_356;
wire v_357;
wire v_358;
wire v_359;
wire v_360;
wire v_363;
wire v_364;
wire v_365;
wire v_366;
wire v_367;
wire v_368;
wire v_369;
wire v_370;
wire v_372;
wire v_373;
wire v_374;
wire v_375;
wire v_376;
wire v_377;
wire v_378;
wire v_379;
wire v_382;
wire v_383;
wire v_385;
wire v_386;
wire v_387;
wire v_388;
wire v_389;
wire v_390;
wire v_391;
wire v_392;
wire v_395;
wire v_396;
wire v_398;
wire v_399;
wire v_400;
wire v_401;
wire v_402;
wire v_403;
wire v_404;
wire v_405;
wire v_408;
wire v_409;
wire v_411;
wire v_412;
wire v_413;
wire v_414;
wire v_415;
wire v_416;
wire v_417;
wire v_418;
wire v_421;
wire v_422;
wire v_424;
wire v_425;
wire v_426;
wire v_427;
wire v_428;
wire v_429;
wire v_430;
wire v_431;
wire v_434;
wire v_435;
wire v_437;
wire v_438;
wire v_439;
wire v_440;
wire v_441;
wire v_442;
wire v_443;
wire v_444;
wire v_447;
wire v_448;
wire v_449;
wire v_450;
wire v_451;
wire v_453;
wire v_454;
wire v_455;
wire v_456;
wire v_457;
wire v_458;
wire v_459;
wire v_460;
wire v_461;
wire v_462;
wire v_463;
wire v_464;
wire v_465;
wire v_468;
wire v_469;
wire v_471;
wire v_472;
wire v_473;
wire v_474;
wire v_475;
wire v_476;
wire v_477;
wire v_478;
wire v_479;
wire v_480;
wire v_483;
wire v_484;
wire v_486;
wire v_487;
wire v_488;
wire v_489;
wire v_490;
wire v_491;
wire v_492;
wire v_493;
wire v_494;
wire v_495;
wire v_497;
wire v_498;
wire v_500;
wire v_501;
wire v_504;
wire v_506;
wire v_507;
wire v_508;
wire v_509;
wire v_510;
wire v_512;
wire v_513;
wire v_514;
wire v_515;
wire v_516;
wire v_517;
wire v_519;
wire v_520;
wire v_521;
wire v_522;
wire v_523;
wire v_524;
wire v_526;
wire v_528;
wire v_529;
wire v_531;
wire v_532;
wire v_533;
wire v_534;
wire v_535;
wire v_536;
wire v_537;
wire v_538;
wire v_540;
wire v_541;
wire v_542;
wire v_543;
wire v_544;
wire v_545;
wire v_546;
wire v_547;
wire v_548;
wire v_549;
wire v_550;
wire v_551;
wire v_552;
wire v_553;
wire v_554;
wire v_555;
wire v_557;
wire v_559;
wire v_561;
wire v_562;
wire v_563;
wire v_564;
wire v_565;
wire v_567;
wire v_568;
wire v_569;
wire v_570;
wire v_571;
wire v_572;
wire v_573;
wire v_574;
wire v_575;
wire v_577;
wire v_578;
wire v_579;
wire v_580;
wire v_581;
wire v_582;
wire v_583;
wire v_584;
wire v_585;
wire v_586;
wire v_587;
wire v_588;
wire v_589;
wire v_590;
wire v_591;
wire v_592;
wire v_593;
wire v_594;
wire v_595;
wire v_596;
wire v_597;
wire v_598;
wire v_599;
wire v_600;
wire v_601;
wire v_602;
wire v_603;
wire v_604;
wire v_605;
wire v_606;
wire v_607;
wire v_608;
wire v_609;
wire v_610;
wire v_611;
wire v_612;
wire v_613;
wire v_614;
wire v_615;
wire v_616;
wire v_617;
wire v_618;
wire v_619;
wire v_620;
wire v_621;
wire v_622;
wire v_623;
wire v_624;
wire v_625;
wire v_626;
wire v_627;
wire v_628;
wire v_629;
wire v_630;
wire v_631;
wire v_632;
wire v_633;
wire v_635;
wire v_636;
wire v_637;
wire v_638;
wire v_639;
wire v_640;
wire v_641;
wire v_642;
wire v_643;
wire v_644;
wire v_645;
wire v_646;
wire v_647;
wire v_648;
wire v_650;
wire v_651;
wire v_652;
wire v_653;
wire v_654;
wire v_655;
wire v_656;
wire v_657;
wire v_659;
wire v_660;
wire v_661;
wire v_662;
wire v_663;
wire v_664;
wire v_665;
wire v_666;
wire v_668;
wire v_669;
wire v_670;
wire v_671;
wire v_672;
wire v_673;
wire v_674;
wire v_675;
wire v_677;
wire v_678;
wire v_679;
wire v_680;
wire v_681;
wire v_682;
wire v_683;
wire v_684;
wire v_685;
wire v_686;
wire v_687;
wire v_688;
wire v_689;
wire v_690;
wire v_691;
wire v_692;
wire v_693;
wire v_694;
wire v_695;
wire v_696;
wire v_697;
wire v_698;
wire v_699;
wire v_700;
wire v_701;
wire v_702;
wire v_703;
wire v_704;
wire v_705;
wire v_706;
wire v_707;
wire v_708;
wire v_709;
wire v_710;
wire v_712;
wire v_713;
wire v_714;
wire v_716;
wire v_717;
wire v_718;
wire v_719;
wire v_720;
wire v_722;
wire v_723;
wire v_724;
wire v_725;
wire v_726;
wire v_727;
wire v_729;
wire v_730;
wire v_731;
wire v_732;
wire v_733;
wire v_735;
wire v_736;
wire v_737;
wire v_738;
wire v_739;
wire v_740;
wire v_742;
wire v_743;
wire v_744;
wire v_745;
wire v_746;
wire v_747;
wire v_748;
wire v_749;
wire v_750;
wire v_751;
wire v_752;
wire v_753;
wire v_754;
wire v_755;
wire v_756;
wire v_757;
wire v_758;
wire v_760;
wire v_761;
wire v_762;
wire v_763;
wire v_764;
wire v_766;
wire v_767;
wire v_768;
wire v_769;
wire v_770;
wire v_771;
wire v_773;
wire v_774;
wire v_775;
wire v_776;
wire v_777;
wire v_778;
wire v_779;
wire v_780;
wire v_781;
wire v_782;
wire v_783;
wire v_784;
wire v_785;
wire v_786;
wire v_787;
wire v_788;
wire v_789;
wire v_790;
wire v_791;
wire v_792;
wire v_793;
wire v_794;
wire v_795;
wire v_796;
wire v_797;
wire v_798;
wire v_799;
wire v_800;
wire v_801;
wire v_802;
wire v_803;
wire v_804;
wire v_805;
wire v_806;
wire v_807;
wire v_808;
wire v_809;
wire v_810;
wire v_811;
wire v_812;
wire v_813;
wire v_814;
wire v_815;
wire v_817;
wire v_818;
wire v_819;
wire v_820;
wire v_821;
wire v_822;
wire v_823;
wire v_824;
wire v_825;
wire v_826;
wire v_827;
wire v_828;
wire v_829;
wire v_830;
wire v_831;
wire v_832;
wire v_833;
wire v_834;
wire v_835;
wire v_836;
wire v_837;
wire v_838;
wire v_839;
wire v_840;
wire v_841;
wire v_842;
wire v_843;
wire v_844;
wire v_845;
wire v_846;
wire v_847;
wire v_848;
wire v_849;
wire v_850;
wire v_851;
wire v_852;
wire v_853;
wire v_854;
wire v_855;
wire v_856;
wire v_857;
wire v_858;
wire v_859;
wire v_860;
wire v_861;
wire v_862;
wire v_863;
wire v_864;
wire v_865;
wire v_866;
wire v_867;
wire v_868;
wire v_869;
wire v_870;
wire v_871;
wire v_872;
wire v_873;
wire v_874;
wire v_875;
wire v_876;
wire v_877;
wire v_878;
wire v_879;
wire v_880;
wire v_881;
wire v_882;
wire v_883;
wire v_884;
wire v_885;
wire v_886;
wire v_887;
wire v_888;
wire v_889;
wire v_890;
wire v_891;
wire v_892;
wire v_893;
wire v_894;
wire v_895;
wire v_896;
wire v_897;
wire v_898;
wire v_899;
wire v_900;
wire v_901;
wire v_902;
wire v_903;
wire v_904;
wire v_905;
wire v_906;
wire v_907;
wire v_908;
wire v_909;
wire v_910;
wire v_911;
wire v_912;
wire v_913;
wire v_914;
wire v_915;
wire v_916;
wire v_917;
wire v_918;
wire v_919;
wire v_920;
wire v_921;
wire v_922;
wire v_923;
wire v_924;
wire v_925;
wire v_926;
wire v_927;
wire v_928;
wire v_929;
wire v_930;
wire v_931;
wire v_932;
wire v_933;
wire v_934;
wire v_935;
wire v_936;
wire v_937;
wire v_938;
wire v_939;
wire v_940;
wire v_941;
wire v_942;
wire v_943;
wire v_944;
wire v_945;
wire v_946;
wire v_947;
wire v_948;
wire v_950;
wire v_951;
wire v_952;
wire v_953;
wire v_954;
wire v_955;
wire v_956;
wire v_957;
wire v_958;
wire v_959;
wire v_960;
wire v_961;
wire v_962;
wire v_963;
wire v_964;
wire v_965;
wire v_966;
wire v_967;
wire v_968;
wire v_969;
wire v_970;
wire v_971;
wire v_973;
wire v_974;
wire v_975;
wire v_976;
wire v_977;
wire v_978;
wire v_979;
wire v_980;
wire v_981;
wire v_982;
wire v_983;
wire v_984;
wire v_986;
wire v_987;
wire v_988;
wire v_989;
wire v_990;
wire v_991;
wire v_992;
wire v_993;
wire v_994;
wire v_995;
wire v_997;
wire v_999;
wire v_1000;
wire v_1001;
wire v_1002;
wire v_1003;
wire v_1004;
wire v_1005;
wire v_1007;
wire v_1009;
wire v_1010;
wire v_1011;
wire v_1012;
wire v_1013;
wire v_1014;
wire v_1015;
wire v_1017;
wire v_1019;
wire v_1020;
wire v_1021;
wire v_1022;
wire v_1023;
wire v_1024;
wire v_1025;
wire v_1027;
wire v_1029;
wire v_1030;
wire v_1031;
wire v_1032;
wire v_1033;
wire v_1034;
wire v_1035;
wire v_1037;
wire v_1039;
wire v_1040;
wire v_1041;
wire v_1042;
wire v_1043;
wire v_1044;
wire v_1045;
wire v_1047;
wire v_1048;
wire v_1050;
wire v_1051;
wire v_1052;
wire v_1053;
wire v_1054;
wire v_1055;
wire v_1057;
wire v_1058;
wire v_1059;
wire v_1060;
wire v_1061;
wire v_1062;
wire v_1063;
wire v_1064;
wire v_1065;
wire v_1066;
wire v_1067;
wire v_1068;
wire v_1070;
wire v_1071;
wire v_1072;
wire v_1073;
wire v_1074;
wire v_1075;
wire v_1076;
wire v_1077;
wire v_1078;
wire v_1079;
wire v_1080;
wire v_1081;
wire v_1083;
wire v_1084;
wire v_1085;
wire v_1086;
wire v_1087;
wire v_1088;
wire v_1089;
wire v_1090;
wire v_1091;
wire v_1092;
wire v_1093;
wire v_1094;
wire v_1096;
wire v_1097;
wire v_1098;
wire v_1099;
wire v_1100;
wire v_1101;
wire v_1102;
wire v_1103;
wire v_1104;
wire v_1105;
wire v_1106;
wire v_1107;
wire v_1109;
wire v_1110;
wire v_1111;
wire v_1112;
wire v_1113;
wire v_1114;
wire v_1115;
wire v_1116;
wire v_1118;
wire v_1119;
wire v_1120;
wire v_1121;
wire v_1122;
wire v_1123;
wire v_1124;
wire v_1125;
wire v_1127;
wire v_1129;
wire v_1130;
wire v_1131;
wire v_1132;
wire v_1133;
wire v_1134;
wire v_1135;
wire v_1137;
wire v_1139;
wire v_1140;
wire v_1141;
wire v_1142;
wire v_1143;
wire v_1144;
wire v_1145;
wire v_1147;
wire v_1149;
wire v_1150;
wire v_1151;
wire v_1152;
wire v_1153;
wire v_1154;
wire v_1155;
wire v_1157;
wire v_1158;
wire v_1159;
wire v_1160;
wire v_1161;
wire v_1162;
wire v_1163;
wire v_1164;
wire v_1166;
wire v_1167;
wire v_1168;
wire v_1169;
wire v_1170;
wire v_1171;
wire v_1172;
wire v_1173;
wire v_1175;
wire v_1176;
wire v_1177;
wire v_1178;
wire v_1179;
wire v_1180;
wire v_1181;
wire v_1182;
wire v_1184;
wire v_1185;
wire v_1186;
wire v_1187;
wire v_1188;
wire v_1189;
wire v_1190;
wire v_1191;
wire v_1192;
wire v_1193;
wire v_1194;
wire v_1195;
wire v_1196;
wire v_1197;
wire v_1198;
wire v_1199;
wire v_1200;
wire v_1201;
wire v_1202;
wire v_1203;
wire v_1204;
wire v_1205;
wire v_1206;
wire v_1207;
wire v_1208;
wire v_1209;
wire v_1210;
wire v_1211;
wire v_1212;
wire v_1213;
wire v_1214;
wire v_1215;
wire v_1216;
wire v_1217;
wire v_1218;
wire v_1219;
wire v_1220;
wire v_1221;
wire v_1222;
wire v_1223;
wire v_1224;
wire v_1225;
wire v_1226;
wire v_1227;
wire v_1228;
wire v_1229;
wire v_1230;
wire v_1231;
wire v_1232;
wire v_1233;
wire v_1234;
wire v_1235;
wire v_1236;
wire v_1237;
wire v_1238;
wire v_1239;
wire v_1240;
wire v_1241;
wire v_1242;
wire v_1243;
wire v_1244;
wire v_1245;
wire v_1246;
wire v_1247;
wire v_1248;
wire v_1249;
wire v_1250;
wire v_1251;
wire v_1252;
wire v_1253;
wire v_1254;
wire v_1255;
wire v_1256;
wire v_1257;
wire v_1258;
wire v_1259;
wire v_1260;
wire v_1261;
wire v_1262;
wire v_1263;
wire v_1264;
wire v_1265;
wire v_1266;
wire v_1267;
wire v_1268;
wire v_1269;
wire v_1270;
wire v_1271;
wire v_1272;
wire v_1273;
wire v_1274;
wire v_1275;
wire v_1276;
wire v_1277;
wire v_1278;
wire v_1279;
wire v_1280;
wire v_1281;
wire v_1282;
wire v_1283;
wire v_1284;
wire v_1285;
wire v_1286;
wire v_1287;
wire v_1288;
wire v_1289;
wire v_1290;
wire v_1291;
wire v_1292;
wire v_1293;
wire v_1294;
wire v_1295;
wire v_1296;
wire v_1297;
wire v_1298;
wire v_1299;
wire v_1300;
wire v_1301;
wire v_1302;
wire v_1303;
wire v_1304;
wire v_1305;
wire v_1306;
wire v_1307;
wire v_1308;
wire v_1309;
wire v_1310;
wire v_1311;
wire v_1312;
wire v_1313;
wire v_1314;
wire v_1315;
wire v_1316;
wire v_1317;
wire v_1318;
wire v_1319;
wire v_1320;
wire v_1321;
wire v_1322;
wire v_1323;
wire v_1324;
wire v_1325;
wire v_1326;
wire v_1327;
wire v_1328;
wire x_1;
assign v_1242 = 1;
assign v_5 = ~v_1 & ~v_2 & v_3 & v_4;
assign v_7 = ~v_1 & v_4 & v_6;
assign v_12 = v_1243 & v_1244;
assign v_14 = v_1245 & v_1246;
assign v_16 = v_1247 & v_1248;
assign v_18 = v_2 & v_4 & ~v_17;
assign v_19 = ~v_1 & v_2 & v_4 & ~v_15;
assign v_20 = ~v_1 & v_4 & ~v_15 & v_17;
assign v_22 = ~v_1 & v_4 & v_21;
assign v_24 = v_23;
assign v_25 = ~v_1 & v_4 & v_9 & v_17;
assign v_26 = ~v_1 & v_4 & v_9 & v_10 & v_15;
assign v_27 = v_3 & v_4 & ~v_17;
assign v_28 = v_4 & v_6 & ~v_17;
assign v_29 = v_4 & ~v_17 & v_21;
assign v_30 = v_4 & v_9 & v_15 & v_17;
assign v_31 = v_4 & v_10 & ~v_13 & v_15 & ~v_17;
assign v_32 = v_4 & ~v_8 & v_10 & v_15 & ~v_17;
assign v_33 = v_4 & ~v_9 & v_15 & ~v_17;
assign v_34 = v_1 & ~v_2 & v_4 & v_10 & v_17;
assign v_35 = v_1 & ~v_2 & v_4 & ~v_9 & v_15;
assign v_36 = v_1 & v_2 & v_4 & v_10 & ~v_11;
assign v_37 = v_1 & v_2 & v_4 & ~v_10 & v_11;
assign v_38 = v_2 & v_4 & v_10 & ~v_15;
assign v_40 = v_4 & v_39;
assign v_41 = v_1249 & v_1250;
assign v_43 = v_4 & v_42;
assign v_44 = ~v_1 & v_3 & v_4 & ~v_10;
assign v_45 = ~v_1 & v_3 & v_4 & ~v_11;
assign v_46 = v_3 & v_4 & ~v_10 & v_15;
assign v_47 = v_1 & v_4 & ~v_9 & ~v_10 & v_15;
assign v_48 = v_4 & v_6 & v_10;
assign v_49 = v_4 & v_10 & v_21;
assign v_50 = v_2 & v_4 & ~v_10 & v_11 & ~v_13;
assign v_51 = v_2 & v_4 & ~v_8 & ~v_10 & v_11;
assign v_52 = ~v_2 & v_4 & v_11 & ~v_13 & v_17;
assign v_53 = ~v_2 & v_4 & ~v_8 & v_11 & v_17;
assign v_54 = v_1251 & v_1252;
assign v_55 = v_4 & v_9 & v_11 & v_15;
assign v_56 = v_1253 & v_1254;
assign v_57 = v_1255 & v_1256;
assign v_58 = v_1257 & v_1258;
assign v_59 = v_1259 & v_1260;
assign v_60 = v_1 & ~v_2 & v_4 & v_11 & v_17;
assign v_64 = v_3 & v_4;
assign v_80 = v_64 & v_79;
assign v_81 = v_65 & ~v_66;
assign v_82 = ~v_68 & v_81;
assign v_83 = ~v_70 & ~v_71;
assign v_84 = ~v_73 & v_83;
assign v_85 = ~v_75 & v_84;
assign v_86 = v_77 & v_85;
assign v_87 = v_82 & v_86;
assign v_89 = v_87 & v_88;
assign v_95 = v_93 & v_94;
assign v_99 = v_4 & v_98;
assign v_100 = v_79 & v_99;
assign v_102 = v_87 & v_101;
assign v_108 = v_106 & v_107;
assign v_112 = v_4 & v_111;
assign v_113 = v_79 & v_112;
assign v_115 = v_87 & v_114;
assign v_121 = v_119 & v_120;
assign v_125 = v_4 & v_124;
assign v_128 = v_125 & v_127;
assign v_129 = v_73 & v_83;
assign v_130 = ~v_75 & v_129;
assign v_132 = v_130 & v_131;
assign v_138 = v_136 & v_137;
assign v_142 = v_4 & v_141;
assign v_143 = v_127 & v_142;
assign v_145 = v_130 & v_144;
assign v_151 = v_149 & v_150;
assign v_154 = v_4 & v_8;
assign v_158 = v_154 & v_157;
assign v_159 = ~v_65 & v_66;
assign v_160 = ~v_68 & v_159;
assign v_161 = v_86 & v_160;
assign v_162 = v_88 & v_161;
assign v_168 = v_166 & v_167;
assign v_171 = v_4 & v_13;
assign v_172 = v_157 & v_171;
assign v_173 = v_101 & v_161;
assign v_179 = v_177 & v_178;
assign v_183 = v_4 & v_182;
assign v_184 = v_127 & v_183;
assign v_186 = v_130 & v_185;
assign v_192 = v_190 & v_191;
assign v_196 = v_4 & v_195;
assign v_197 = v_127 & v_196;
assign v_199 = v_130 & v_198;
assign v_205 = v_203 & v_204;
assign v_209 = v_4 & v_208;
assign v_210 = v_127 & v_209;
assign v_212 = v_130 & v_211;
assign v_218 = v_216 & v_217;
assign v_222 = v_4 & v_221;
assign v_223 = v_127 & v_222;
assign v_225 = v_130 & v_224;
assign v_231 = v_229 & v_230;
assign v_235 = v_4 & v_234;
assign v_236 = v_127 & v_235;
assign v_238 = v_130 & v_237;
assign v_244 = v_242 & v_243;
assign v_248 = v_4 & v_247;
assign v_249 = v_127 & v_248;
assign v_251 = v_130 & v_250;
assign v_257 = v_255 & v_256;
assign v_260 = v_4 & v_9;
assign v_263 = v_2 & v_4;
assign v_268 = v_4 & v_6;
assign v_273 = v_266 & v_272;
assign v_279 = v_273 & v_278;
assign v_288 = v_268 & v_287;
assign v_289 = v_283 & v_288;
assign v_290 = v_64 & v_99;
assign v_291 = v_112 & v_290;
assign v_292 = v_154 & v_171;
assign v_293 = v_261 & v_267;
assign v_294 = v_275 & v_293;
assign v_295 = ~v_70 & v_71;
assign v_296 = ~v_73 & v_295;
assign v_297 = v_75 & v_296;
assign v_298 = v_294 & v_297;
assign v_299 = v_292 & v_298;
assign v_300 = v_291 & v_299;
assign v_302 = v_154 & v_176;
assign v_303 = v_298 & v_302;
assign v_306 = v_267 & v_268;
assign v_307 = v_275 & v_306;
assign v_308 = v_265 & v_307;
assign v_309 = v_260 & v_261;
assign v_310 = v_275 & v_309;
assign v_311 = v_271 & v_310;
assign v_313 = v_263 & v_293;
assign v_314 = v_277 & v_313;
assign v_316 = v_297 & v_315;
assign v_317 = v_277 & v_297;
assign v_318 = v_260 & v_268;
assign v_319 = v_275 & v_318;
assign v_320 = v_317 & v_319;
assign v_330 = v_322 & v_329;
assign v_333 = v_330 & v_332;
assign v_336 = v_165 & v_171;
assign v_337 = v_298 & v_336;
assign v_339 = v_260 & v_283;
assign v_340 = v_287 & v_339;
assign v_345 = v_329 & v_344;
assign v_348 = v_345 & v_347;
assign v_352 = v_263 & v_351;
assign v_354 = v_345 & v_353;
assign v_356 = v_293 & v_317;
assign v_358 = v_328 & v_357;
assign v_363 = v_4 & v_362;
assign v_367 = v_363 & v_366;
assign v_368 = v_70 & ~v_71;
assign v_369 = ~v_73 & v_368;
assign v_370 = ~v_75 & v_369;
assign v_372 = v_370 & v_371;
assign v_378 = v_376 & v_377;
assign v_382 = v_4 & v_381;
assign v_383 = v_366 & v_382;
assign v_385 = v_370 & v_384;
assign v_391 = v_389 & v_390;
assign v_395 = v_4 & v_394;
assign v_396 = v_366 & v_395;
assign v_398 = v_370 & v_397;
assign v_404 = v_402 & v_403;
assign v_408 = v_4 & v_407;
assign v_409 = v_366 & v_408;
assign v_411 = v_370 & v_410;
assign v_417 = v_415 & v_416;
assign v_421 = v_4 & v_420;
assign v_422 = v_366 & v_421;
assign v_424 = v_370 & v_423;
assign v_430 = v_428 & v_429;
assign v_434 = v_4 & v_433;
assign v_435 = v_366 & v_434;
assign v_437 = v_370 & v_436;
assign v_443 = v_441 & v_442;
assign v_447 = v_4 & v_446;
assign v_451 = v_447 & v_450;
assign v_453 = v_4 & v_452;
assign v_454 = v_65 & v_66;
assign v_455 = ~v_68 & v_454;
assign v_456 = v_86 & v_455;
assign v_457 = v_453 & v_456;
assign v_464 = v_461 & v_463;
assign v_468 = v_4 & v_467;
assign v_469 = v_450 & v_468;
assign v_471 = v_4 & v_470;
assign v_472 = v_456 & v_471;
assign v_479 = v_476 & v_478;
assign v_483 = v_4 & v_482;
assign v_484 = v_450 & v_483;
assign v_486 = v_4 & v_485;
assign v_487 = v_456 & v_486;
assign v_494 = v_491 & v_493;
assign v_504 = v_4 & v_503;
assign v_508 = v_4 & v_505;
assign v_510 = v_507 & v_509;
assign v_514 = v_4 & v_511;
assign v_516 = v_513 & v_515;
assign v_517 = v_510 & v_516;
assign v_521 = v_4 & v_518;
assign v_523 = v_520 & v_522;
assign v_524 = v_517 & v_523;
assign v_528 = v_4 & v_527;
assign v_529 = v_526 & v_528;
assign v_532 = v_529 & v_531;
assign v_533 = v_4 & v_530;
assign v_534 = v_4 & v_525;
assign v_536 = v_534 & v_535;
assign v_537 = v_533 & v_536;
assign v_541 = v_538 & v_540;
assign v_544 = v_542 & v_543;
assign v_547 = v_545 & v_546;
assign v_548 = v_544 & v_547;
assign v_551 = v_549 & v_550;
assign v_552 = v_548 & v_551;
assign v_553 = v_541 & v_552;
assign v_554 = v_524 & v_553;
assign v_555 = v_504 & v_554;
assign v_557 = v_555 & v_556;
assign v_559 = v_4 & v_558;
assign v_562 = v_559 & v_561;
assign v_563 = v_557 & v_562;
assign v_568 = v_4 & v_560;
assign v_569 = v_567 & v_568;
assign v_575 = v_570 & v_574;
assign v_577 = v_4 & v_576;
assign v_579 = v_568 & v_578;
assign v_580 = ~v_65 & ~v_66;
assign v_581 = ~v_68 & v_580;
assign v_582 = ~v_77 & v_85;
assign v_583 = v_581 & v_582;
assign v_584 = v_579 & v_583;
assign v_588 = v_427 & v_508;
assign v_589 = v_421 & v_506;
assign v_591 = v_414 & v_514;
assign v_592 = v_408 & v_512;
assign v_595 = v_440 & v_521;
assign v_596 = v_434 & v_519;
assign v_603 = v_600 & v_602;
assign v_604 = v_4 & v_539;
assign v_606 = v_99 & v_388;
assign v_607 = v_105 & v_382;
assign v_609 = v_64 & v_375;
assign v_610 = v_92 & v_363;
assign v_613 = v_112 & v_401;
assign v_614 = v_118 & v_395;
assign v_623 = v_559 & v_568;
assign v_624 = v_566 & v_623;
assign v_626 = v_622 & v_625;
assign v_629 = v_88 & v_628;
assign v_632 = v_627 & v_631;
assign v_635 = v_567 & v_623;
assign v_637 = v_574 & v_636;
assign v_639 = v_583 & v_638;
assign v_643 = v_621 & v_642;
assign v_645 = v_564 & v_578;
assign v_647 = v_644 & v_646;
assign v_650 = v_79 & v_514;
assign v_651 = v_64 & v_87;
assign v_656 = v_654 & v_655;
assign v_659 = v_79 & v_508;
assign v_660 = v_87 & v_99;
assign v_665 = v_663 & v_664;
assign v_668 = v_79 & v_521;
assign v_669 = v_87 & v_112;
assign v_674 = v_672 & v_673;
assign v_677 = v_70 & v_71;
assign v_678 = v_73 & v_677;
assign v_679 = ~v_75 & v_678;
assign v_682 = v_680 & v_681;
assign v_684 = v_682 & v_683;
assign v_685 = v_4 & v_39;
assign v_686 = v_684 & v_685;
assign v_687 = v_679 & v_686;
assign v_688 = v_73 & v_368;
assign v_689 = ~v_75 & v_688;
assign v_690 = v_4 & v_17;
assign v_691 = v_1 & v_4;
assign v_692 = v_690 & v_691;
assign v_693 = v_4 & v_42;
assign v_694 = v_692 & v_693;
assign v_696 = v_694 & v_695;
assign v_697 = v_689 & v_696;
assign v_699 = v_73 & v_295;
assign v_700 = ~v_75 & v_699;
assign v_701 = v_681 & v_690;
assign v_702 = v_693 & v_701;
assign v_703 = v_695 & v_702;
assign v_704 = v_700 & v_703;
assign v_714 = v_706 & v_713;
assign v_716 = v_4 & v_715;
assign v_720 = v_717 & v_719;
assign v_722 = v_4 & v_721;
assign v_726 = v_723 & v_725;
assign v_727 = v_720 & v_726;
assign v_731 = v_4 & v_728;
assign v_733 = v_730 & v_732;
assign v_737 = v_4 & v_734;
assign v_739 = v_736 & v_738;
assign v_740 = v_733 & v_739;
assign v_744 = v_4 & v_741;
assign v_746 = v_743 & v_745;
assign v_747 = v_740 & v_746;
assign v_750 = v_748 & v_749;
assign v_753 = v_751 & v_752;
assign v_754 = v_750 & v_753;
assign v_757 = v_755 & v_756;
assign v_758 = v_754 & v_757;
assign v_762 = v_4 & v_759;
assign v_764 = v_761 & v_763;
assign v_768 = v_4 & v_765;
assign v_770 = v_767 & v_769;
assign v_771 = v_764 & v_770;
assign v_775 = v_4 & v_772;
assign v_777 = v_774 & v_776;
assign v_778 = v_771 & v_777;
assign v_781 = v_779 & v_780;
assign v_784 = v_782 & v_783;
assign v_785 = v_781 & v_784;
assign v_788 = v_786 & v_787;
assign v_789 = v_785 & v_788;
assign v_790 = v_778 & v_789;
assign v_791 = v_758 & v_790;
assign v_792 = v_747 & v_791;
assign v_793 = v_727 & v_792;
assign v_794 = v_533 & v_793;
assign v_797 = v_714 & v_796;
assign v_798 = v_682 & v_693;
assign v_799 = v_695 & v_798;
assign v_800 = v_624 & v_799;
assign v_801 = ~v_711 & v_800;
assign v_802 = v_297 & v_801;
assign v_804 = v_531 & v_793;
assign v_811 = v_803 & v_810;
assign v_818 = v_811 & v_817;
assign v_819 = v_683 & v_701;
assign v_820 = v_695 & v_819;
assign v_821 = v_314 & v_820;
assign v_822 = v_297 & v_821;
assign v_828 = v_823 & v_827;
assign v_829 = ~v_73 & v_677;
assign v_830 = ~v_75 & v_829;
assign v_831 = v_684 & v_695;
assign v_832 = v_830 & v_831;
assign v_846 = v_840 & v_845;
assign v_853 = v_846 & v_852;
assign v_854 = v_681 & v_853;
assign v_855 = v_680 & v_691;
assign v_856 = v_693 & v_855;
assign v_857 = v_695 & v_856;
assign v_858 = v_624 & v_857;
assign v_859 = v_711 & v_858;
assign v_860 = v_297 & v_859;
assign v_862 = v_142 & v_718;
assign v_863 = v_148 & v_716;
assign v_865 = v_125 & v_724;
assign v_866 = v_135 & v_722;
assign v_869 = v_506 & v_731;
assign v_870 = v_508 & v_729;
assign v_872 = v_512 & v_737;
assign v_873 = v_514 & v_735;
assign v_876 = v_519 & v_744;
assign v_877 = v_521 & v_742;
assign v_880 = v_105 & v_196;
assign v_881 = v_99 & v_202;
assign v_883 = v_92 & v_183;
assign v_884 = v_64 & v_189;
assign v_887 = v_118 & v_209;
assign v_888 = v_112 & v_215;
assign v_891 = v_475 & v_762;
assign v_892 = v_468 & v_760;
assign v_894 = v_460 & v_768;
assign v_895 = v_447 & v_766;
assign v_898 = v_490 & v_775;
assign v_899 = v_483 & v_773;
assign v_902 = v_235 & v_477;
assign v_903 = v_241 & v_471;
assign v_905 = v_222 & v_462;
assign v_906 = v_228 & v_453;
assign v_909 = v_248 & v_492;
assign v_910 = v_254 & v_486;
assign v_918 = v_858 & v_917;
assign v_919 = v_297 & v_918;
assign v_923 = v_920 & v_922;
assign v_925 = v_800 & v_924;
assign v_926 = v_297 & v_925;
assign v_928 = v_683 & v_692;
assign v_929 = v_695 & v_928;
assign v_930 = v_130 & v_929;
assign v_931 = ~v_816 & v_930;
assign v_937 = v_932 & v_936;
assign v_938 = v_683 & v_855;
assign v_939 = v_695 & v_938;
assign v_940 = v_311 & v_939;
assign v_941 = v_297 & v_940;
assign v_947 = v_942 & v_946;
assign v_950 = v_297 & v_800;
assign v_951 = v_75 & v_84;
assign v_952 = v_685 & v_938;
assign v_953 = v_951 & v_952;
assign v_958 = v_815 & v_957;
assign v_965 = v_680 & v_964;
assign v_966 = v_853 & v_965;
assign v_967 = v_796 & v_966;
assign v_968 = v_961 & v_967;
assign v_970 = v_827 & v_969;
assign v_974 = v_693 & v_853;
assign v_975 = v_973 & v_974;
assign v_976 = v_810 & v_975;
assign v_979 = v_297 & v_858;
assign v_983 = v_815 & v_982;
assign v_986 = v_685 & v_964;
assign v_987 = v_853 & v_986;
assign v_993 = v_973 & v_992;
assign v_994 = v_810 & v_993;
assign v_997 = v_366 & v_722;
assign v_999 = v_370 & v_998;
assign v_1004 = v_1002 & v_1003;
assign v_1007 = v_366 & v_716;
assign v_1009 = v_370 & v_1008;
assign v_1014 = v_1012 & v_1013;
assign v_1017 = v_127 & v_737;
assign v_1019 = v_130 & v_1018;
assign v_1024 = v_1022 & v_1023;
assign v_1027 = v_127 & v_731;
assign v_1029 = v_130 & v_1028;
assign v_1034 = v_1032 & v_1033;
assign v_1037 = v_127 & v_744;
assign v_1039 = v_130 & v_1038;
assign v_1044 = v_1042 & v_1043;
assign v_1051 = v_814 & v_1050;
assign v_1053 = v_4 & v_10;
assign v_1059 = v_4 & v_11;
assign v_1061 = v_1058 & v_1060;
assign v_1062 = v_814 & v_1061;
assign v_1064 = v_1053 & v_1059;
assign v_1065 = v_1050 & v_1057;
assign v_1070 = v_4 & v_15;
assign v_1074 = v_1071 & v_1073;
assign v_1075 = v_814 & v_1074;
assign v_1077 = v_1058 & v_1072;
assign v_1078 = v_1064 & v_1070;
assign v_1083 = v_4 & v_21;
assign v_1084 = v_1073 & v_1083;
assign v_1086 = v_1078 & v_1085;
assign v_1088 = v_814 & v_1087;
assign v_1092 = v_1090 & v_1091;
assign v_1098 = v_534 & v_1097;
assign v_1099 = v_68 & v_454;
assign v_1100 = v_86 & v_1099;
assign v_1101 = v_88 & v_1100;
assign v_1106 = v_1104 & v_1105;
assign v_1109 = v_528 & v_1097;
assign v_1110 = v_101 & v_1100;
assign v_1115 = v_1113 & v_1114;
assign v_1118 = v_604 & v_1097;
assign v_1119 = v_114 & v_1100;
assign v_1124 = v_1122 & v_1123;
assign v_1127 = v_127 & v_768;
assign v_1129 = v_130 & v_1128;
assign v_1134 = v_1132 & v_1133;
assign v_1137 = v_127 & v_762;
assign v_1139 = v_130 & v_1138;
assign v_1144 = v_1142 & v_1143;
assign v_1147 = v_127 & v_775;
assign v_1149 = v_130 & v_1148;
assign v_1154 = v_1152 & v_1153;
assign v_1157 = v_450 & v_453;
assign v_1158 = v_88 & v_456;
assign v_1163 = v_1161 & v_1162;
assign v_1166 = v_450 & v_471;
assign v_1167 = v_101 & v_456;
assign v_1172 = v_1170 & v_1171;
assign v_1175 = v_450 & v_486;
assign v_1176 = v_114 & v_456;
assign v_1181 = v_1179 & v_1180;
assign v_1185 = v_75 & v_1184;
assign v_1187 = v_1083 & v_1186;
assign v_1190 = ~v_70 & ~v_73;
assign v_1192 = v_1065 & v_1072;
assign v_1194 = v_1191 & v_1193;
assign v_1205 = ~v_1183;
assign v_1240 = v_1270 & v_1271;
assign v_1241 = v_1295 & v_1296 & v_1297 & v_1298 & v_1299;
assign v_1243 = ~v_1 & v_4 & ~v_8 & v_9 & ~v_10;
assign v_1244 = ~v_11;
assign v_1245 = ~v_1 & v_4 & v_9 & ~v_10 & ~v_11;
assign v_1246 = ~v_13;
assign v_1247 = ~v_1 & v_4 & v_9 & ~v_10 & ~v_11;
assign v_1248 = ~v_15;
assign v_1249 = v_4 & v_9 & ~v_10 & ~v_11 & ~v_15;
assign v_1250 = ~v_17;
assign v_1251 = ~v_1 & ~v_2 & v_4 & ~v_9 & v_10;
assign v_1252 = v_11;
assign v_1253 = ~v_1 & v_4 & v_8 & ~v_9 & v_11;
assign v_1254 = ~v_17;
assign v_1255 = ~v_1 & v_4 & ~v_9 & v_11 & ~v_13;
assign v_1256 = ~v_17;
assign v_1257 = ~v_2 & v_4 & v_8 & ~v_9 & v_10;
assign v_1258 = v_11;
assign v_1259 = ~v_2 & v_4 & ~v_9 & v_10 & v_11;
assign v_1260 = ~v_13;
assign v_1261 = v_1196 & v_1197 & v_1198 & v_1199 & v_1200;
assign v_1262 = v_1201 & v_1202 & v_1203 & v_1204 & v_1205;
assign v_1263 = v_1206 & v_1207 & v_1208 & v_1209 & v_1210;
assign v_1264 = v_1211 & v_1212 & v_1213 & v_1214 & v_1215;
assign v_1265 = v_1216 & v_1217 & v_1218 & v_1219 & v_1220;
assign v_1266 = v_1221 & v_1222 & v_1223 & v_1224 & v_1225;
assign v_1267 = v_1226 & v_1227 & v_1228 & v_1229 & v_1230;
assign v_1268 = v_1231 & v_1232 & v_1233 & v_1234 & v_1235;
assign v_1269 = v_1236 & v_1237 & v_1238 & v_1239;
assign v_1270 = v_1261 & v_1262 & v_1263 & v_1264 & v_1265;
assign v_1271 = v_1266 & v_1267 & v_1268 & v_1269;
assign v_1272 = v_62 & v_91 & v_96 & v_104 & v_109;
assign v_1273 = v_117 & v_122 & v_134 & v_139 & v_147;
assign v_1274 = v_152 & v_164 & v_169 & v_175 & v_180;
assign v_1275 = v_188 & v_193 & v_201 & v_206 & v_214;
assign v_1276 = v_219 & v_227 & v_232 & v_240 & v_245;
assign v_1277 = v_253 & v_258 & v_305 & v_334 & v_342;
assign v_1278 = v_349 & v_355 & v_360 & v_374 & v_379;
assign v_1279 = v_387 & v_392 & v_400 & v_405 & v_413;
assign v_1280 = v_418 & v_426 & v_431 & v_439 & v_444;
assign v_1281 = v_459 & v_465 & v_474 & v_480 & v_489;
assign v_1282 = v_495 & v_497 & v_498 & v_500 & v_501;
assign v_1283 = v_586 & v_633 & v_641 & v_648 & v_653;
assign v_1284 = v_657 & v_662 & v_666 & v_671 & v_675;
assign v_1285 = v_834 & v_948 & v_960 & v_971 & v_978;
assign v_1286 = v_984 & v_990 & v_995 & v_1001 & v_1005;
assign v_1287 = v_1011 & v_1015 & v_1021 & v_1025 & v_1031;
assign v_1288 = v_1035 & v_1041 & v_1045 & v_1047 & v_1048;
assign v_1289 = v_1052 & v_1055 & v_1063 & v_1068 & v_1076;
assign v_1290 = v_1081 & v_1089 & v_1094 & v_1103 & v_1107;
assign v_1291 = v_1112 & v_1116 & v_1121 & v_1125 & v_1131;
assign v_1292 = v_1135 & v_1141 & v_1145 & v_1151 & v_1155;
assign v_1293 = v_1160 & v_1164 & v_1169 & v_1173 & v_1178;
assign v_1294 = v_1182 & v_1189 & v_1195 & v_1240;
assign v_1295 = v_1272 & v_1273 & v_1274 & v_1275 & v_1276;
assign v_1296 = v_1277 & v_1278 & v_1279 & v_1280 & v_1281;
assign v_1297 = v_1282 & v_1283 & v_1284 & v_1285 & v_1286;
assign v_1298 = v_1287 & v_1288 & v_1289 & v_1290 & v_1291;
assign v_1299 = v_1292 & v_1293 & v_1294;
assign v_61 = v_1309 | v_1310;
assign v_67 = ~v_65 | v_66;
assign v_69 = v_67 | v_68;
assign v_72 = v_70 | v_71;
assign v_74 = v_72 | v_73;
assign v_76 = v_74 | v_75;
assign v_78 = v_76 | ~v_77;
assign v_79 = v_69 | v_78;
assign v_90 = v_80 | v_89;
assign v_91 = ~v_63 | v_90;
assign v_92 = ~v_3 | ~v_4;
assign v_93 = v_87 | v_92;
assign v_94 = v_79 | ~v_88;
assign v_96 = v_63 | v_95;
assign v_103 = v_100 | v_102;
assign v_104 = ~v_97 | v_103;
assign v_105 = ~v_4 | ~v_98;
assign v_106 = v_87 | v_105;
assign v_107 = v_79 | ~v_101;
assign v_109 = v_97 | v_108;
assign v_116 = v_113 | v_115;
assign v_117 = ~v_110 | v_116;
assign v_118 = ~v_4 | ~v_111;
assign v_119 = v_87 | v_118;
assign v_120 = v_79 | ~v_114;
assign v_122 = v_110 | v_121;
assign v_126 = v_72 | ~v_73;
assign v_127 = v_75 | v_126;
assign v_133 = v_128 | v_132;
assign v_134 = ~v_123 | v_133;
assign v_135 = ~v_4 | ~v_124;
assign v_136 = v_130 | v_135;
assign v_137 = v_127 | ~v_131;
assign v_139 = v_123 | v_138;
assign v_146 = v_143 | v_145;
assign v_147 = ~v_140 | v_146;
assign v_148 = ~v_4 | ~v_141;
assign v_149 = v_130 | v_148;
assign v_150 = v_127 | ~v_144;
assign v_152 = v_140 | v_151;
assign v_155 = v_65 | ~v_66;
assign v_156 = v_68 | v_155;
assign v_157 = v_78 | v_156;
assign v_163 = v_158 | v_162;
assign v_164 = ~v_153 | v_163;
assign v_165 = ~v_4 | ~v_8;
assign v_166 = v_161 | v_165;
assign v_167 = ~v_88 | v_157;
assign v_169 = v_153 | v_168;
assign v_174 = v_172 | v_173;
assign v_175 = ~v_170 | v_174;
assign v_176 = ~v_4 | ~v_13;
assign v_177 = v_161 | v_176;
assign v_178 = ~v_101 | v_157;
assign v_180 = v_170 | v_179;
assign v_187 = v_184 | v_186;
assign v_188 = ~v_181 | v_187;
assign v_189 = ~v_4 | ~v_182;
assign v_190 = v_130 | v_189;
assign v_191 = v_127 | ~v_185;
assign v_193 = v_181 | v_192;
assign v_200 = v_197 | v_199;
assign v_201 = ~v_194 | v_200;
assign v_202 = ~v_4 | ~v_195;
assign v_203 = v_130 | v_202;
assign v_204 = v_127 | ~v_198;
assign v_206 = v_194 | v_205;
assign v_213 = v_210 | v_212;
assign v_214 = ~v_207 | v_213;
assign v_215 = ~v_4 | ~v_208;
assign v_216 = v_130 | v_215;
assign v_217 = v_127 | ~v_211;
assign v_219 = v_207 | v_218;
assign v_226 = v_223 | v_225;
assign v_227 = ~v_220 | v_226;
assign v_228 = ~v_4 | ~v_221;
assign v_229 = v_130 | v_228;
assign v_230 = v_127 | ~v_224;
assign v_232 = v_220 | v_231;
assign v_239 = v_236 | v_238;
assign v_240 = ~v_233 | v_239;
assign v_241 = ~v_4 | ~v_234;
assign v_242 = v_130 | v_241;
assign v_243 = v_127 | ~v_237;
assign v_245 = v_233 | v_244;
assign v_252 = v_249 | v_251;
assign v_253 = ~v_246 | v_252;
assign v_254 = ~v_4 | ~v_247;
assign v_255 = v_130 | v_254;
assign v_256 = v_127 | ~v_250;
assign v_258 = v_246 | v_257;
assign v_261 = ~v_4 | ~v_6;
assign v_262 = v_260 | v_261;
assign v_264 = v_262 | v_263;
assign v_266 = v_264 | ~v_265;
assign v_267 = ~v_4 | ~v_9;
assign v_269 = v_267 | v_268;
assign v_270 = v_263 | v_269;
assign v_272 = v_270 | ~v_271;
assign v_274 = v_260 | v_268;
assign v_275 = ~v_2 | ~v_4;
assign v_276 = v_274 | v_275;
assign v_278 = v_276 | ~v_277;
assign v_280 = v_70 | ~v_71;
assign v_281 = v_73 | v_280;
assign v_282 = ~v_75 | v_281;
assign v_283 = v_279 | v_282;
assign v_284 = ~v_277 | v_282;
assign v_285 = v_261 | v_267;
assign v_286 = v_263 | v_285;
assign v_287 = v_284 | v_286;
assign v_301 = v_289 | v_300;
assign v_304 = v_301 | v_303;
assign v_305 = ~v_259 | v_304;
assign v_312 = v_308 | v_311;
assign v_315 = v_312 | v_314;
assign v_321 = v_261 | v_320;
assign v_322 = v_316 | v_321;
assign v_323 = v_92 | v_105;
assign v_324 = v_118 | v_323;
assign v_325 = v_165 | v_176;
assign v_326 = v_263 | v_274;
assign v_327 = v_282 | v_326;
assign v_328 = v_325 | v_327;
assign v_329 = v_324 | v_328;
assign v_331 = v_165 | v_171;
assign v_332 = v_327 | v_331;
assign v_334 = v_259 | v_333;
assign v_338 = v_300 | v_337;
assign v_341 = v_338 | v_340;
assign v_342 = ~v_335 | v_341;
assign v_343 = v_154 | v_176;
assign v_344 = v_327 | v_343;
assign v_346 = v_267 | v_316;
assign v_347 = v_320 | v_346;
assign v_349 = v_335 | v_348;
assign v_351 = v_274 | v_284;
assign v_353 = v_299 | v_352;
assign v_355 = ~v_350 | v_354;
assign v_357 = v_275 | v_356;
assign v_359 = v_338 | v_358;
assign v_360 = v_350 | v_359;
assign v_364 = ~v_70 | v_71;
assign v_365 = v_73 | v_364;
assign v_366 = v_75 | v_365;
assign v_373 = v_367 | v_372;
assign v_374 = ~v_361 | v_373;
assign v_375 = ~v_4 | ~v_362;
assign v_376 = v_370 | v_375;
assign v_377 = v_366 | ~v_371;
assign v_379 = v_361 | v_378;
assign v_386 = v_383 | v_385;
assign v_387 = ~v_380 | v_386;
assign v_388 = ~v_4 | ~v_381;
assign v_389 = v_370 | v_388;
assign v_390 = v_366 | ~v_384;
assign v_392 = v_380 | v_391;
assign v_399 = v_396 | v_398;
assign v_400 = ~v_393 | v_399;
assign v_401 = ~v_4 | ~v_394;
assign v_402 = v_370 | v_401;
assign v_403 = v_366 | ~v_397;
assign v_405 = v_393 | v_404;
assign v_412 = v_409 | v_411;
assign v_413 = ~v_406 | v_412;
assign v_414 = ~v_4 | ~v_407;
assign v_415 = v_370 | v_414;
assign v_416 = v_366 | ~v_410;
assign v_418 = v_406 | v_417;
assign v_425 = v_422 | v_424;
assign v_426 = ~v_419 | v_425;
assign v_427 = ~v_4 | ~v_420;
assign v_428 = v_370 | v_427;
assign v_429 = v_366 | ~v_423;
assign v_431 = v_419 | v_430;
assign v_438 = v_435 | v_437;
assign v_439 = ~v_432 | v_438;
assign v_440 = ~v_4 | ~v_433;
assign v_441 = v_370 | v_440;
assign v_442 = v_366 | ~v_436;
assign v_444 = v_432 | v_443;
assign v_448 = ~v_65 | ~v_66;
assign v_449 = v_68 | v_448;
assign v_450 = v_78 | v_449;
assign v_458 = v_451 | v_457;
assign v_459 = ~v_445 | v_458;
assign v_460 = ~v_4 | ~v_446;
assign v_461 = v_456 | v_460;
assign v_462 = ~v_4 | ~v_452;
assign v_463 = v_450 | v_462;
assign v_465 = v_445 | v_464;
assign v_473 = v_469 | v_472;
assign v_474 = ~v_466 | v_473;
assign v_475 = ~v_4 | ~v_467;
assign v_476 = v_456 | v_475;
assign v_477 = ~v_4 | ~v_470;
assign v_478 = v_450 | v_477;
assign v_480 = v_466 | v_479;
assign v_488 = v_484 | v_487;
assign v_489 = ~v_481 | v_488;
assign v_490 = ~v_4 | ~v_482;
assign v_491 = v_456 | v_490;
assign v_492 = ~v_4 | ~v_485;
assign v_493 = v_450 | v_492;
assign v_495 = v_481 | v_494;
assign v_497 = v_114 | ~v_496;
assign v_498 = ~v_114 | v_496;
assign v_500 = v_88 | ~v_499;
assign v_501 = ~v_88 | v_499;
assign v_506 = ~v_4 | ~v_505;
assign v_507 = v_421 | v_506;
assign v_509 = v_427 | v_508;
assign v_512 = ~v_4 | ~v_511;
assign v_513 = v_408 | v_512;
assign v_515 = v_414 | v_514;
assign v_519 = ~v_4 | ~v_518;
assign v_520 = v_434 | v_519;
assign v_522 = v_440 | v_521;
assign v_526 = ~v_4 | ~v_525;
assign v_531 = ~v_4 | ~v_530;
assign v_535 = ~v_4 | ~v_527;
assign v_538 = v_532 | v_537;
assign v_540 = ~v_4 | ~v_539;
assign v_542 = v_105 | v_382;
assign v_543 = v_99 | v_388;
assign v_545 = v_92 | v_363;
assign v_546 = v_64 | v_375;
assign v_549 = v_118 | v_395;
assign v_550 = v_112 | v_401;
assign v_561 = ~v_4 | ~v_560;
assign v_564 = ~v_4 | ~v_558;
assign v_565 = v_561 | v_564;
assign v_567 = v_565 | ~v_566;
assign v_570 = v_563 | v_569;
assign v_571 = v_65 | v_66;
assign v_572 = v_68 | v_571;
assign v_573 = v_76 | v_77;
assign v_574 = v_572 | v_573;
assign v_578 = ~v_88 | v_577;
assign v_585 = v_575 | v_584;
assign v_586 = ~v_502 | v_585;
assign v_587 = ~v_4 | ~v_503;
assign v_590 = v_588 | v_589;
assign v_593 = v_591 | v_592;
assign v_594 = v_590 | v_593;
assign v_597 = v_595 | v_596;
assign v_598 = v_594 | v_597;
assign v_599 = v_534 | v_535;
assign v_600 = v_533 | v_599;
assign v_601 = v_526 | v_528;
assign v_602 = v_531 | v_601;
assign v_605 = v_603 | v_604;
assign v_608 = v_606 | v_607;
assign v_611 = v_609 | v_610;
assign v_612 = v_608 | v_611;
assign v_615 = v_613 | v_614;
assign v_616 = v_612 | v_615;
assign v_617 = v_605 | v_616;
assign v_618 = v_598 | v_617;
assign v_619 = v_587 | v_618;
assign v_620 = ~v_556 | v_619;
assign v_621 = v_564 | v_568;
assign v_622 = v_620 | v_621;
assign v_625 = v_561 | v_624;
assign v_627 = v_583 | v_626;
assign v_628 = ~v_4 | ~v_576;
assign v_630 = v_561 | v_629;
assign v_631 = v_574 | v_630;
assign v_633 = v_502 | v_632;
assign v_636 = v_562 | v_635;
assign v_638 = v_559 | v_629;
assign v_640 = v_637 | v_639;
assign v_641 = ~v_634 | v_640;
assign v_642 = v_565 | v_624;
assign v_644 = v_583 | v_643;
assign v_646 = v_574 | v_645;
assign v_648 = v_634 | v_647;
assign v_652 = v_650 | v_651;
assign v_653 = ~v_649 | v_652;
assign v_654 = v_87 | v_512;
assign v_655 = v_79 | v_92;
assign v_657 = v_649 | v_656;
assign v_661 = v_659 | v_660;
assign v_662 = ~v_658 | v_661;
assign v_663 = v_87 | v_506;
assign v_664 = v_79 | v_105;
assign v_666 = v_658 | v_665;
assign v_670 = v_668 | v_669;
assign v_671 = ~v_667 | v_670;
assign v_672 = v_87 | v_519;
assign v_673 = v_79 | v_118;
assign v_675 = v_667 | v_674;
assign v_680 = ~v_4 | ~v_17;
assign v_681 = ~v_1 | ~v_4;
assign v_683 = ~v_4 | ~v_42;
assign v_695 = ~v_4 | ~v_39;
assign v_698 = v_687 | v_697;
assign v_705 = v_698 | v_704;
assign v_706 = v_691 | v_705;
assign v_707 = v_681 | v_690;
assign v_708 = v_683 | v_707;
assign v_709 = v_685 | v_708;
assign v_710 = v_567 | v_709;
assign v_712 = v_710 | ~v_711;
assign v_713 = v_282 | v_712;
assign v_717 = v_148 | v_716;
assign v_718 = ~v_4 | ~v_715;
assign v_719 = v_142 | v_718;
assign v_723 = v_135 | v_722;
assign v_724 = ~v_4 | ~v_721;
assign v_725 = v_125 | v_724;
assign v_729 = ~v_4 | ~v_728;
assign v_730 = v_508 | v_729;
assign v_732 = v_506 | v_731;
assign v_735 = ~v_4 | ~v_734;
assign v_736 = v_514 | v_735;
assign v_738 = v_512 | v_737;
assign v_742 = ~v_4 | ~v_741;
assign v_743 = v_521 | v_742;
assign v_745 = v_519 | v_744;
assign v_748 = v_99 | v_202;
assign v_749 = v_105 | v_196;
assign v_751 = v_64 | v_189;
assign v_752 = v_92 | v_183;
assign v_755 = v_112 | v_215;
assign v_756 = v_118 | v_209;
assign v_760 = ~v_4 | ~v_759;
assign v_761 = v_468 | v_760;
assign v_763 = v_475 | v_762;
assign v_766 = ~v_4 | ~v_765;
assign v_767 = v_447 | v_766;
assign v_769 = v_460 | v_768;
assign v_773 = ~v_4 | ~v_772;
assign v_774 = v_483 | v_773;
assign v_776 = v_490 | v_775;
assign v_779 = v_241 | v_471;
assign v_780 = v_235 | v_477;
assign v_782 = v_228 | v_453;
assign v_783 = v_222 | v_462;
assign v_786 = v_254 | v_486;
assign v_787 = v_248 | v_492;
assign v_795 = v_710 | v_794;
assign v_796 = v_282 | v_795;
assign v_803 = v_797 | v_802;
assign v_805 = v_690 | v_691;
assign v_806 = v_683 | v_805;
assign v_807 = v_685 | v_806;
assign v_808 = v_567 | v_807;
assign v_809 = v_804 | v_808;
assign v_810 = v_282 | v_809;
assign v_812 = v_680 | v_681;
assign v_813 = v_693 | v_812;
assign v_814 = v_685 | v_813;
assign v_815 = v_127 | v_814;
assign v_817 = v_815 | v_816;
assign v_823 = v_818 | v_822;
assign v_824 = v_693 | v_707;
assign v_825 = v_685 | v_824;
assign v_826 = v_272 | v_825;
assign v_827 = v_282 | v_826;
assign v_833 = v_828 | v_832;
assign v_834 = ~v_676 | v_833;
assign v_835 = ~v_70 | ~v_71;
assign v_836 = ~v_73 | v_835;
assign v_837 = v_75 | v_836;
assign v_838 = v_693 | v_805;
assign v_839 = v_695 | v_838;
assign v_840 = v_837 | v_839;
assign v_841 = ~v_73 | v_364;
assign v_842 = v_75 | v_841;
assign v_843 = v_683 | v_812;
assign v_844 = v_685 | v_843;
assign v_845 = v_842 | v_844;
assign v_847 = ~v_73 | v_280;
assign v_848 = v_75 | v_847;
assign v_849 = v_680 | v_691;
assign v_850 = v_683 | v_849;
assign v_851 = v_685 | v_850;
assign v_852 = v_848 | v_851;
assign v_861 = v_854 | v_860;
assign v_864 = v_862 | v_863;
assign v_867 = v_865 | v_866;
assign v_868 = v_864 | v_867;
assign v_871 = v_869 | v_870;
assign v_874 = v_872 | v_873;
assign v_875 = v_871 | v_874;
assign v_878 = v_876 | v_877;
assign v_879 = v_875 | v_878;
assign v_882 = v_880 | v_881;
assign v_885 = v_883 | v_884;
assign v_886 = v_882 | v_885;
assign v_889 = v_887 | v_888;
assign v_890 = v_886 | v_889;
assign v_893 = v_891 | v_892;
assign v_896 = v_894 | v_895;
assign v_897 = v_893 | v_896;
assign v_900 = v_898 | v_899;
assign v_901 = v_897 | v_900;
assign v_904 = v_902 | v_903;
assign v_907 = v_905 | v_906;
assign v_908 = v_904 | v_907;
assign v_911 = v_909 | v_910;
assign v_912 = v_908 | v_911;
assign v_913 = v_901 | v_912;
assign v_914 = v_890 | v_913;
assign v_915 = v_879 | v_914;
assign v_916 = v_868 | v_915;
assign v_917 = v_531 | v_916;
assign v_920 = v_861 | v_919;
assign v_921 = v_711 | v_808;
assign v_922 = v_282 | v_921;
assign v_924 = v_533 | v_916;
assign v_927 = v_923 | v_926;
assign v_932 = v_927 | v_931;
assign v_933 = v_693 | v_849;
assign v_934 = v_685 | v_933;
assign v_935 = v_278 | v_934;
assign v_936 = v_282 | v_935;
assign v_942 = v_937 | v_941;
assign v_943 = v_73 | v_835;
assign v_944 = v_75 | v_943;
assign v_945 = v_685 | v_838;
assign v_946 = v_944 | v_945;
assign v_948 = v_676 | v_947;
assign v_954 = v_690 | v_953;
assign v_955 = v_705 | v_954;
assign v_956 = v_919 | v_955;
assign v_957 = v_950 | v_956;
assign v_959 = v_941 | v_958;
assign v_960 = ~v_949 | v_959;
assign v_961 = v_282 | v_808;
assign v_962 = v_74 | ~v_75;
assign v_963 = v_695 | v_824;
assign v_964 = v_962 | v_963;
assign v_969 = v_930 | v_968;
assign v_971 = v_949 | v_970;
assign v_973 = v_282 | v_710;
assign v_977 = v_930 | v_976;
assign v_978 = ~v_972 | v_977;
assign v_980 = v_683 | v_705;
assign v_981 = v_979 | v_980;
assign v_982 = v_926 | v_981;
assign v_984 = v_972 | v_983;
assign v_988 = v_979 | v_987;
assign v_989 = v_926 | v_988;
assign v_990 = ~v_985 | v_989;
assign v_991 = v_695 | v_953;
assign v_992 = v_705 | v_991;
assign v_995 = v_985 | v_994;
assign v_1000 = v_997 | v_999;
assign v_1001 = ~v_996 | v_1000;
assign v_1002 = v_370 | v_724;
assign v_1003 = v_366 | ~v_998;
assign v_1005 = v_996 | v_1004;
assign v_1010 = v_1007 | v_1009;
assign v_1011 = ~v_1006 | v_1010;
assign v_1012 = v_370 | v_718;
assign v_1013 = v_366 | ~v_1008;
assign v_1015 = v_1006 | v_1014;
assign v_1020 = v_1017 | v_1019;
assign v_1021 = ~v_1016 | v_1020;
assign v_1022 = v_130 | v_735;
assign v_1023 = v_127 | ~v_1018;
assign v_1025 = v_1016 | v_1024;
assign v_1030 = v_1027 | v_1029;
assign v_1031 = ~v_1026 | v_1030;
assign v_1032 = v_130 | v_729;
assign v_1033 = v_127 | ~v_1028;
assign v_1035 = v_1026 | v_1034;
assign v_1040 = v_1037 | v_1039;
assign v_1041 = ~v_1036 | v_1040;
assign v_1042 = v_130 | v_742;
assign v_1043 = v_127 | ~v_1038;
assign v_1045 = v_1036 | v_1044;
assign v_1047 = v_101 | ~v_1046;
assign v_1048 = ~v_101 | v_1046;
assign v_1050 = ~v_4 | ~v_10;
assign v_1052 = ~v_1049 | v_1051;
assign v_1054 = v_929 | v_1053;
assign v_1055 = v_1049 | v_1054;
assign v_1057 = ~v_4 | ~v_11;
assign v_1058 = v_1050 | v_1057;
assign v_1060 = v_1053 | v_1059;
assign v_1063 = ~v_1056 | v_1062;
assign v_1066 = v_1064 | v_1065;
assign v_1067 = v_929 | v_1066;
assign v_1068 = v_1056 | v_1067;
assign v_1071 = v_1064 | v_1070;
assign v_1072 = ~v_4 | ~v_15;
assign v_1073 = v_1058 | v_1072;
assign v_1076 = ~v_1069 | v_1075;
assign v_1079 = v_1077 | v_1078;
assign v_1080 = v_929 | v_1079;
assign v_1081 = v_1069 | v_1080;
assign v_1085 = ~v_4 | ~v_21;
assign v_1087 = v_1084 | v_1086;
assign v_1089 = ~v_1082 | v_1088;
assign v_1090 = v_1078 | v_1085;
assign v_1091 = v_1073 | v_1083;
assign v_1093 = v_929 | v_1092;
assign v_1094 = v_1082 | v_1093;
assign v_1096 = ~v_68 | v_448;
assign v_1097 = v_78 | v_1096;
assign v_1102 = v_1098 | v_1101;
assign v_1103 = ~v_1095 | v_1102;
assign v_1104 = v_526 | v_1100;
assign v_1105 = ~v_88 | v_1097;
assign v_1107 = v_1095 | v_1106;
assign v_1111 = v_1109 | v_1110;
assign v_1112 = ~v_1108 | v_1111;
assign v_1113 = v_535 | v_1100;
assign v_1114 = ~v_101 | v_1097;
assign v_1116 = v_1108 | v_1115;
assign v_1120 = v_1118 | v_1119;
assign v_1121 = ~v_1117 | v_1120;
assign v_1122 = v_540 | v_1100;
assign v_1123 = ~v_114 | v_1097;
assign v_1125 = v_1117 | v_1124;
assign v_1130 = v_1127 | v_1129;
assign v_1131 = ~v_1126 | v_1130;
assign v_1132 = v_130 | v_766;
assign v_1133 = v_127 | ~v_1128;
assign v_1135 = v_1126 | v_1134;
assign v_1140 = v_1137 | v_1139;
assign v_1141 = ~v_1136 | v_1140;
assign v_1142 = v_130 | v_760;
assign v_1143 = v_127 | ~v_1138;
assign v_1145 = v_1136 | v_1144;
assign v_1150 = v_1147 | v_1149;
assign v_1151 = ~v_1146 | v_1150;
assign v_1152 = v_130 | v_773;
assign v_1153 = v_127 | ~v_1148;
assign v_1155 = v_1146 | v_1154;
assign v_1159 = v_1157 | v_1158;
assign v_1160 = ~v_1156 | v_1159;
assign v_1161 = v_456 | v_462;
assign v_1162 = ~v_88 | v_450;
assign v_1164 = v_1156 | v_1163;
assign v_1168 = v_1166 | v_1167;
assign v_1169 = ~v_1165 | v_1168;
assign v_1170 = v_456 | v_477;
assign v_1171 = ~v_101 | v_450;
assign v_1173 = v_1165 | v_1172;
assign v_1177 = v_1175 | v_1176;
assign v_1178 = ~v_1174 | v_1177;
assign v_1179 = v_456 | v_492;
assign v_1180 = ~v_114 | v_450;
assign v_1182 = v_1174 | v_1181;
assign v_1184 = v_70 | v_73;
assign v_1186 = v_1060 | v_1070;
assign v_1188 = v_1185 | v_1187;
assign v_1189 = ~v_1183 | v_1188;
assign v_1191 = ~v_75 | v_1190;
assign v_1193 = v_1085 | v_1192;
assign v_1195 = v_1183 | v_1194;
assign v_1196 = ~v_62 | ~v_63 | v_350 | v_676;
assign v_1197 = ~v_62 | ~v_259 | v_676;
assign v_1198 = v_1311 | v_1312;
assign v_1199 = v_1313 | v_1314;
assign v_1200 = v_1315 | v_1316;
assign v_1201 = ~v_62 | ~v_350 | v_949;
assign v_1202 = ~v_62 | ~v_350 | v_676 | v_1069;
assign v_1203 = ~v_62 | v_676 | ~v_949 | v_1069;
assign v_1204 = ~v_62 | v_676 | ~v_1082;
assign v_1206 = ~v_62 | ~v_335 | v_676 | ~v_949;
assign v_1207 = ~v_62 | ~v_335 | v_676 | ~v_1049 | ~v_1069;
assign v_1208 = ~v_62 | ~v_63 | v_949;
assign v_1209 = ~v_62 | ~v_259 | v_949;
assign v_1210 = ~v_62 | v_949 | ~v_1082;
assign v_1211 = ~v_62 | ~v_335 | ~v_949 | ~v_1069;
assign v_1212 = ~v_62 | v_170 | v_949 | ~v_1049 | ~v_1069;
assign v_1213 = ~v_62 | v_153 | v_949 | ~v_1049 | ~v_1069;
assign v_1214 = ~v_62 | v_335 | v_949 | ~v_1069;
assign v_1215 = ~v_62 | v_350 | ~v_676 | ~v_949 | ~v_1049;
assign v_1216 = ~v_62 | v_335 | v_350 | ~v_676 | ~v_1069;
assign v_1217 = ~v_62 | ~v_350 | ~v_676 | ~v_1049 | v_1056;
assign v_1218 = ~v_62 | ~v_350 | ~v_676 | v_1049 | ~v_1056;
assign v_1219 = ~v_62 | ~v_350 | ~v_1049 | v_1069;
assign v_1220 = ~v_62 | ~v_985;
assign v_1221 = v_1317 | v_1318;
assign v_1222 = ~v_62 | ~v_972;
assign v_1223 = ~v_62 | ~v_63 | v_676 | v_1049;
assign v_1224 = ~v_62 | ~v_63 | v_676 | v_1056;
assign v_1225 = ~v_62 | ~v_63 | v_1049 | ~v_1069;
assign v_1226 = ~v_62 | v_335 | ~v_676 | v_1049 | ~v_1069;
assign v_1227 = ~v_62 | ~v_259 | ~v_1049;
assign v_1228 = ~v_62 | ~v_1049 | ~v_1082;
assign v_1229 = ~v_62 | v_170 | ~v_350 | v_1049 | ~v_1056;
assign v_1230 = ~v_62 | v_153 | ~v_350 | v_1049 | ~v_1056;
assign v_1231 = ~v_62 | v_170 | v_350 | ~v_949 | ~v_1056;
assign v_1232 = ~v_62 | v_153 | v_350 | ~v_949 | ~v_1056;
assign v_1233 = v_1319 | v_1320;
assign v_1234 = ~v_62 | ~v_335 | ~v_1056 | ~v_1069;
assign v_1235 = v_1321 | v_1322;
assign v_1236 = v_1323 | v_1324;
assign v_1237 = v_1325 | v_1326;
assign v_1238 = v_1327 | v_1328;
assign v_1239 = ~v_62 | v_350 | ~v_676 | ~v_949 | ~v_1056;
assign v_1300 = v_5 | v_7 | v_12 | v_14 | v_16;
assign v_1301 = v_18 | v_19 | v_20 | v_22 | v_24;
assign v_1302 = v_25 | v_26 | v_27 | v_28 | v_29;
assign v_1303 = v_30 | v_31 | v_32 | v_33 | v_34;
assign v_1304 = v_35 | v_36 | v_37 | v_38 | v_40;
assign v_1305 = v_41 | v_43 | v_44 | v_45 | v_46;
assign v_1306 = v_47 | v_48 | v_49 | v_50 | v_51;
assign v_1307 = v_52 | v_53 | v_54 | v_55 | v_56;
assign v_1308 = v_57 | v_58 | v_59 | v_60;
assign v_1309 = v_1300 | v_1301 | v_1302 | v_1303 | v_1304;
assign v_1310 = v_1305 | v_1306 | v_1307 | v_1308;
assign v_1311 = ~v_62 | v_153 | ~v_335 | v_676 | v_1049;
assign v_1312 = v_1056;
assign v_1313 = ~v_62 | v_170 | ~v_335 | v_676 | v_1049;
assign v_1314 = v_1056;
assign v_1315 = ~v_62 | ~v_335 | v_676 | v_1049 | v_1056;
assign v_1316 = v_1069;
assign v_1317 = ~v_62 | ~v_335 | v_949 | v_1049 | v_1056;
assign v_1318 = v_1069;
assign v_1319 = ~v_62 | v_335 | v_350 | v_676 | ~v_1049;
assign v_1320 = ~v_1056;
assign v_1321 = ~v_62 | ~v_153 | v_335 | v_676 | v_949;
assign v_1322 = ~v_1056;
assign v_1323 = ~v_62 | v_170 | v_335 | v_676 | v_949;
assign v_1324 = ~v_1056;
assign v_1325 = ~v_62 | ~v_153 | v_335 | v_350 | ~v_1049;
assign v_1326 = ~v_1056;
assign v_1327 = ~v_62 | v_170 | v_335 | v_350 | ~v_1049;
assign v_1328 = ~v_1056;
assign x_1 = v_61 | v_1241;
assign o_1 = x_1;
endmodule
